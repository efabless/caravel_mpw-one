* SPICE NETLIST
***************************************

.SUBCKT MN g s d b
.ENDS
***************************************
.SUBCKT MP g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT condiodeHvPsub pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20nativevhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT n20nativevhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT p20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_3 VNB VPB VGND VPWR
** N=20 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=0.59 W=0.55 AD=0.143 AS=0.143 PD=1.62 PS=1.62 NRD=0 NRS=0 m=1 r=0.932203 sa=295000 sb=295000 a=0.3245 p=2.28 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=0.59 W=0.87 AD=0.2262 AS=0.2262 PD=2.26 PS=2.26 NRD=0 NRS=0 m=1 r=1.47458 sa=295000 sb=295000 a=0.5133 p=2.92 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT ICV_1 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 1 0 $X=-190 $Y=-2960
X1 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_2 1 2
** N=2 EP=2 IP=4 FDC=8
*.SEEDPROM
X0 1 2 ICV_1 $T=0 -5440 0 0 $X=-190 $Y=-8400
X1 1 2 ICV_1 $T=0 0 0 0 $X=-190 $Y=-2960
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__fill_1
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VNB VPB VGND VPWR
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__fill_2
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VNB VPB VGND VPWR
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_4 VNB VPB VGND VPWR
** N=20 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=1.05 W=0.55 AD=0.143 AS=0.143 PD=1.62 PS=1.62 NRD=0 NRS=0 m=1 r=0.52381 sa=525000 sb=525000 a=0.5775 p=3.2 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=1.05 W=0.87 AD=0.2262 AS=0.2262 PD=2.26 PS=2.26 NRD=0 NRS=0 m=1 r=0.828571 sa=525000 sb=525000 a=0.9135 p=3.84 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT ICV_3 1 2
** N=2 EP=2 IP=8 FDC=2
*.SEEDPROM
X1 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_6 VNB VPB VGND VPWR
** N=22 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=1.97 W=0.55 AD=0.143 AS=0.143 PD=1.62 PS=1.62 NRD=0 NRS=0 m=1 r=0.279188 sa=984999 sb=984999 a=1.0835 p=5.04 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=1.97 W=0.87 AD=0.2262 AS=0.2262 PD=2.26 PS=2.26 NRD=0 NRS=0 m=1 r=0.441624 sa=984999 sb=984999 a=1.7139 p=5.68 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT ICV_4 1 2
** N=2 EP=2 IP=8 FDC=2
*.SEEDPROM
X1 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_8 VNB VPB VGND VPWR
** N=24 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=2.89 W=0.55 AD=0.143 AS=0.143 PD=1.62 PS=1.62 NRD=0 NRS=0 m=1 r=0.190311 sa=1.445e+06 sb=1.445e+06 a=1.5895 p=6.88 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=2.89 W=0.87 AD=0.2262 AS=0.2262 PD=2.26 PS=2.26 NRD=0 NRS=0 m=1 r=0.301038 sa=1.445e+06 sb=1.445e+06 a=2.5143 p=7.52 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__decap_12 VNB VPB VGND VPWR
** N=26 EP=4 IP=0 FDC=2
*.SEEDPROM
M0 VGND VPWR VGND VNB nshort L=4.73 W=0.55 AD=0.143 AS=0.143 PD=1.62 PS=1.62 NRD=0 NRS=0 m=1 r=0.116279 sa=2.365e+06 sb=2.365e+06 a=2.6015 p=10.56 mult=1 $X=395 $Y=235 $D=9
M1 VPWR VGND VPWR VPB phighvt L=4.73 W=0.87 AD=0.2262 AS=0.2262 PD=2.26 PS=2.26 NRD=0 NRS=0 m=1 r=0.183932 sa=2.365e+06 sb=2.365e+06 a=4.1151 p=11.2 mult=1 $X=395 $Y=1615 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__clkbuf_8 VNB VPB A VPWR X VGND
** N=149 EP=6 IP=0 FDC=20
*.SEEDPROM
M0 7 A VGND VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75004.1 a=0.063 p=1.14 mult=1 $X=400 $Y=235 $D=9
M1 VGND A 7 VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75000.6 sb=75003.6 a=0.063 p=1.14 mult=1 $X=830 $Y=235 $D=9
M2 X 7 VGND VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75001.1 sb=75003.2 a=0.063 p=1.14 mult=1 $X=1260 $Y=235 $D=9
M3 VGND 7 X VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75001.5 sb=75002.8 a=0.063 p=1.14 mult=1 $X=1690 $Y=235 $D=9
M4 X 7 VGND VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75001.9 sb=75002.3 a=0.063 p=1.14 mult=1 $X=2120 $Y=235 $D=9
M5 VGND 7 X VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75002.3 sb=75001.9 a=0.063 p=1.14 mult=1 $X=2550 $Y=235 $D=9
M6 X 7 VGND VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75002.8 sb=75001.5 a=0.063 p=1.14 mult=1 $X=2980 $Y=235 $D=9
M7 VGND 7 X VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75003.2 sb=75001.1 a=0.063 p=1.14 mult=1 $X=3410 $Y=235 $D=9
M8 X 7 VGND VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75003.6 sb=75000.6 a=0.063 p=1.14 mult=1 $X=3840 $Y=235 $D=9
M9 VGND 7 X VNB nshort L=0.15 W=0.42 AD=0.1134 AS=0.0588 PD=1.38 PS=0.7 NRD=1.428 NRS=0 m=1 r=2.8 sa=75004.1 sb=75000.2 a=0.063 p=1.14 mult=1 $X=4270 $Y=235 $D=9
M10 7 A VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=6.66667 sa=75000.2 sb=75004.1 a=0.15 p=2.3 mult=1 $X=400 $Y=1485 $D=89
M11 VPWR A 7 VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75000.6 sb=75003.6 a=0.15 p=2.3 mult=1 $X=830 $Y=1485 $D=89
M12 X 7 VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75001 sb=75003.2 a=0.15 p=2.3 mult=1 $X=1260 $Y=1485 $D=89
M13 VPWR 7 X VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75001.5 sb=75002.8 a=0.15 p=2.3 mult=1 $X=1690 $Y=1485 $D=89
M14 X 7 VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75001.9 sb=75002.3 a=0.15 p=2.3 mult=1 $X=2120 $Y=1485 $D=89
M15 VPWR 7 X VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75002.3 sb=75001.9 a=0.15 p=2.3 mult=1 $X=2550 $Y=1485 $D=89
M16 X 7 VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75002.8 sb=75001.5 a=0.15 p=2.3 mult=1 $X=2980 $Y=1485 $D=89
M17 VPWR 7 X VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75003.2 sb=75001 a=0.15 p=2.3 mult=1 $X=3410 $Y=1485 $D=89
M18 X 7 VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75003.6 sb=75000.6 a=0.15 p=2.3 mult=1 $X=3840 $Y=1485 $D=89
M19 VPWR 7 X VPB phighvt L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75004.1 sb=75000.2 a=0.15 p=2.3 mult=1 $X=4270 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__ebufn_2 VNB VPB A TE_B VPWR Z VGND
** N=72 EP=7 IP=0 FDC=12
*.SEEDPROM
M0 VGND A 9 VNB nshort L=0.15 W=0.42 AD=0.07875 AS=0.1092 PD=0.795 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75000.7 a=0.063 p=1.14 mult=1 $X=395 $Y=235 $D=9
M1 8 TE_B VGND VNB nshort L=0.15 W=0.42 AD=0.1092 AS=0.07875 PD=1.36 PS=0.795 NRD=0 NRS=28.56 m=1 r=2.8 sa=75000.7 sb=75000.2 a=0.063 p=1.14 mult=1 $X=920 $Y=235 $D=9
M2 VGND 8 11 VNB nshort L=0.15 W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 m=1 r=4.33333 sa=75000.2 sb=75001.6 a=0.0975 p=1.6 mult=1 $X=2220 $Y=235 $D=9
M3 11 8 VGND VNB nshort L=0.15 W=0.65 AD=0.125125 AS=0.08775 PD=1.035 PS=0.92 NRD=9.228 NRS=0 m=1 r=4.33333 sa=75000.6 sb=75001.1 a=0.0975 p=1.6 mult=1 $X=2640 $Y=235 $D=9
M4 Z 9 11 VNB nshort L=0.15 W=0.65 AD=0.08775 AS=0.125125 PD=0.92 PS=1.035 NRD=0 NRS=10.152 m=1 r=4.33333 sa=75001.1 sb=75000.6 a=0.0975 p=1.6 mult=1 $X=3175 $Y=235 $D=9
M5 11 9 Z VNB nshort L=0.15 W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75001.6 sb=75000.2 a=0.0975 p=1.6 mult=1 $X=3595 $Y=235 $D=9
M6 VPWR A 9 VPB phighvt L=0.15 W=0.64 AD=0.12 AS=0.1664 PD=1.015 PS=1.8 NRD=15.3857 NRS=0 m=1 r=4.26667 sa=75000.2 sb=75000.7 a=0.096 p=1.58 mult=1 $X=395 $Y=1845 $D=89
M7 8 TE_B VPWR VPB phighvt L=0.15 W=0.64 AD=0.1664 AS=0.12 PD=1.8 PS=1.015 NRD=0 NRS=13.8491 m=1 r=4.26667 sa=75000.7 sb=75000.2 a=0.096 p=1.58 mult=1 $X=920 $Y=1845 $D=89
M8 VPWR TE_B 10 VPB phighvt L=0.15 W=0.94 AD=0.1269 AS=0.2444 PD=1.21 PS=2.4 NRD=0 NRS=0 m=1 r=6.26667 sa=75000.2 sb=75001.9 a=0.141 p=2.18 mult=1 $X=1860 $Y=1545 $D=89
M9 10 TE_B VPWR VPB phighvt L=0.15 W=0.94 AD=0.358799 AS=0.1269 PD=1.69103 PS=1.21 NRD=11.5245 NRS=0 m=1 r=6.26667 sa=75000.6 sb=75001.5 a=0.141 p=2.18 mult=1 $X=2280 $Y=1545 $D=89
M10 Z 9 10 VPB phighvt L=0.15 W=1 AD=0.135 AS=0.381701 PD=1.27 PS=1.79897 NRD=0 NRS=13.7703 m=1 r=6.66667 sa=75001.4 sb=75000.6 a=0.15 p=2.3 mult=1 $X=3175 $Y=1485 $D=89
M11 10 9 Z VPB phighvt L=0.15 W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75001.9 sb=75000.2 a=0.15 p=2.3 mult=1 $X=3595 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__tapvpwrvgnd_1
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VGND VPWR
.ENDS
***************************************
.SUBCKT ICV_5 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=12
*.SEEDPROM
X0 1 2 3 4 2 5 1 sky130_fd_sc_hd__ebufn_2 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_7
** N=2 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_8
** N=2 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_9 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=5520 0 0 0 $X=5330 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_10 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_11 1 2
** N=2 EP=2 IP=8 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=5520 0 0 0 $X=5330 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_12 1 2
** N=2 EP=2 IP=6 FDC=6
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=11040 0 0 0 $X=10850 $Y=-240
X1 1 2 ICV_11 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__dfxtp_1 VNB VPB CLK D VPWR Q VGND
** N=142 EP=7 IP=0 FDC=24
*.SEEDPROM
M0 VGND CLK 8 VNB nshort L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75000.6 a=0.063 p=1.14 mult=1 $X=395 $Y=235 $D=9
M1 9 8 VGND VNB nshort L=0.15 W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 m=1 r=2.8 sa=75000.6 sb=75000.2 a=0.063 p=1.14 mult=1 $X=815 $Y=235 $D=9
M2 14 D VGND VNB nshort L=0.15 W=0.42 AD=0.0875538 AS=0.1092 PD=0.893846 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75003.3 a=0.063 p=1.14 mult=1 $X=1755 $Y=235 $D=9
M3 11 8 14 VNB nshort L=0.15 W=0.36 AD=0.0621 AS=0.0750462 PD=0.705 PS=0.766154 NRD=0 NRS=43.332 m=1 r=2.4 sa=75000.7 sb=75003.3 a=0.054 p=1.02 mult=1 $X=2315 $Y=235 $D=9
M4 17 9 11 VNB nshort L=0.15 W=0.36 AD=0.0642462 AS=0.0621 PD=0.706154 PS=0.705 NRD=41.148 NRS=23.328 m=1 r=2.4 sa=75001.2 sb=75002.8 a=0.054 p=1.02 mult=1 $X=2810 $Y=235 $D=9
M5 VGND 10 17 VNB nshort L=0.15 W=0.42 AD=0.0958472 AS=0.0749538 PD=0.859811 PS=0.823846 NRD=0 NRS=35.268 m=1 r=2.8 sa=75001.5 sb=75002.1 a=0.063 p=1.14 mult=1 $X=3305 $Y=235 $D=9
M6 10 11 VGND VNB nshort L=0.15 W=0.64 AD=0.126592 AS=0.146053 PD=1.2736 PS=1.31019 NRD=0 NRS=30.936 m=1 r=4.26667 sa=75001.4 sb=75001 a=0.096 p=1.58 mult=1 $X=3900 $Y=235 $D=9
M7 13 9 10 VNB nshort L=0.15 W=0.36 AD=0.0684 AS=0.071208 PD=0.74 PS=0.7164 NRD=3.324 NRS=24.996 m=1 r=2.4 sa=75002.8 sb=75001.2 a=0.054 p=1.02 mult=1 $X=4405 $Y=235 $D=9
M8 18 8 13 VNB nshort L=0.15 W=0.36 AD=0.0609231 AS=0.0684 PD=0.687692 PS=0.74 NRD=38.076 NRS=30 m=1 r=2.4 sa=75003.4 sb=75000.7 a=0.054 p=1.02 mult=1 $X=4935 $Y=235 $D=9
M9 VGND 12 18 VNB nshort L=0.15 W=0.42 AD=0.1092 AS=0.0710769 PD=1.36 PS=0.802308 NRD=0 NRS=32.628 m=1 r=2.8 sa=75003.3 sb=75000.2 a=0.063 p=1.14 mult=1 $X=5410 $Y=235 $D=9
M10 VGND 13 12 VNB nshort L=0.15 W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 m=1 r=4.33333 sa=75000.2 sb=75000.6 a=0.0975 p=1.6 mult=1 $X=6355 $Y=235 $D=9
M11 Q 12 VGND VNB nshort L=0.15 W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75000.6 sb=75000.2 a=0.0975 p=1.6 mult=1 $X=6775 $Y=235 $D=9
M12 VPWR CLK 8 VPB phighvt L=0.15 W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 m=1 r=4.26667 sa=75000.2 sb=75000.6 a=0.096 p=1.58 mult=1 $X=395 $Y=1815 $D=89
M13 9 8 VPWR VPB phighvt L=0.15 W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 m=1 r=4.26667 sa=75000.6 sb=75000.2 a=0.096 p=1.58 mult=1 $X=815 $Y=1815 $D=89
M14 14 D VPWR VPB phighvt L=0.15 W=0.42 AD=0.05775 AS=0.1092 PD=0.695 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75003.7 a=0.063 p=1.14 mult=1 $X=1755 $Y=2065 $D=89
M15 11 9 14 VPB phighvt L=0.15 W=0.42 AD=0.06825 AS=0.05775 PD=0.745 PS=0.695 NRD=14.0658 NRS=0 m=1 r=2.8 sa=75000.6 sb=75003.3 a=0.063 p=1.14 mult=1 $X=2180 $Y=2065 $D=89
M16 15 8 11 VPB phighvt L=0.15 W=0.42 AD=0.07665 AS=0.06825 PD=0.785 PS=0.745 NRD=59.7895 NRS=7.0329 m=1 r=2.8 sa=75001.1 sb=75002.8 a=0.063 p=1.14 mult=1 $X=2655 $Y=2065 $D=89
M17 VPWR 10 15 VPB phighvt L=0.15 W=0.42 AD=0.128423 AS=0.07665 PD=0.904615 PS=0.785 NRD=111.384 NRS=59.7895 m=1 r=2.8 sa=75001.6 sb=75002.3 a=0.063 p=1.14 mult=1 $X=3170 $Y=2065 $D=89
M18 10 11 VPWR VPB phighvt L=0.15 W=0.75 AD=0.140385 AS=0.229327 PD=1.37821 PS=1.61538 NRD=0 NRS=0 m=1 r=5 sa=75001.4 sb=75001 a=0.1125 p=1.8 mult=1 $X=3830 $Y=1735 $D=89
M19 13 8 10 VPB phighvt L=0.15 W=0.42 AD=0.0567 AS=0.0786154 PD=0.69 PS=0.771795 NRD=0 NRS=23.443 m=1 r=2.8 sa=75002.7 sb=75001.2 a=0.063 p=1.14 mult=1 $X=4305 $Y=2065 $D=89
M20 16 9 13 VPB phighvt L=0.15 W=0.42 AD=0.0882 AS=0.0567 PD=0.84 PS=0.69 NRD=72.693 NRS=0 m=1 r=2.8 sa=75003.2 sb=75000.8 a=0.063 p=1.14 mult=1 $X=4725 $Y=2065 $D=89
M21 VPWR 12 16 VPB phighvt L=0.15 W=0.42 AD=0.1113 AS=0.0882 PD=1.37 PS=0.84 NRD=0 NRS=72.693 m=1 r=2.8 sa=75003.7 sb=75000.2 a=0.063 p=1.14 mult=1 $X=5295 $Y=2065 $D=89
M22 VPWR 13 12 VPB phighvt L=0.15 W=1 AD=0.135 AS=0.27 PD=1.27 PS=2.54 NRD=0 NRS=0.9653 m=1 r=6.66667 sa=75000.2 sb=75000.6 a=0.15 p=2.3 mult=1 $X=6345 $Y=1485 $D=89
M23 Q 12 VPWR VPB phighvt L=0.15 W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75000.6 sb=75000.2 a=0.15 p=2.3 mult=1 $X=6765 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_13 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=14 FDC=36
*.SEEDPROM
X0 1 2 3 4 2 5 1 sky130_fd_sc_hd__ebufn_2 $T=7360 0 0 0 $X=7170 $Y=-240
X1 1 2 6 7 2 8 1 sky130_fd_sc_hd__dfxtp_1 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_14 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=36
*.SEEDPROM
X1 1 2 6 7 8 3 4 5 ICV_13 $T=920 0 0 0 $X=730 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_15 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=15 FDC=48
*.SEEDPROM
X0 1 2 3 4 2 5 1 sky130_fd_sc_hd__ebufn_2 $T=11500 0 0 0 $X=11310 $Y=-240
X1 1 2 9 10 11 6 7 8 ICV_13 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=36
*.SEEDPROM
X1 1 2 6 7 8 3 4 5 ICV_13 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_17 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=38
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 6 7 8 3 4 5 ICV_13 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_18
** N=2 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_19 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=38
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 6 7 8 3 4 5 ICV_13 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_20 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=24
*.SEEDPROM
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__dfxtp_1 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_21 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=26
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 3 4 5 ICV_20 $T=2760 0 0 0 $X=2570 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_22 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=10 FDC=38
*.SEEDPROM
X0 1 2 ICV_3 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 6 7 8 3 4 5 ICV_13 $T=2300 0 0 0 $X=2110 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_23 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_24 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__inv_1 VNB VPB A VPWR Y VGND
** N=25 EP=6 IP=0 FDC=2
*.SEEDPROM
M0 Y A VGND VNB nshort L=0.15 W=0.65 AD=0.169 AS=0.169 PD=1.82 PS=1.82 NRD=0 NRS=0 m=1 r=4.33333 sa=75000.2 sb=75000.2 a=0.0975 p=1.6 mult=1 $X=600 $Y=235 $D=9
M1 Y A VPWR VPB phighvt L=0.15 W=1 AD=0.26 AS=0.26 PD=2.52 PS=2.52 NRD=0 NRS=0 m=1 r=6.66667 sa=75000.2 sb=75000.2 a=0.15 p=2.3 mult=1 $X=600 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_25 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_26 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=12
*.SEEDPROM
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__ebufn_2 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_27 1 2 3 4 5 6 7
** N=7 EP=7 IP=13 FDC=26
*.SEEDPROM
X0 1 2 3 4 2 5 1 sky130_fd_sc_hd__dfxtp_1 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 6 2 7 1 sky130_fd_sc_hd__inv_1 $T=7360 0 0 0 $X=7170 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_28 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=26
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__dfxtp_1 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_29 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=26
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 3 4 5 ICV_20 $T=1840 0 0 0 $X=1650 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_30 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=14 FDC=24
*.SEEDPROM
X0 1 2 3 4 2 5 1 sky130_fd_sc_hd__ebufn_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 6 7 2 8 1 sky130_fd_sc_hd__ebufn_2 $T=4140 0 0 0 $X=3950 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__and2_1 VNB VPB A B VPWR X VGND
** N=37 EP=7 IP=0 FDC=6
*.SEEDPROM
M0 9 A 8 VNB nshort L=0.15 W=0.42 AD=0.0567 AS=0.1176 PD=0.69 PS=1.4 NRD=22.848 NRS=0 m=1 r=2.8 sa=75000.2 sb=75001.2 a=0.063 p=1.14 mult=1 $X=575 $Y=375 $D=9
M1 VGND B 9 VNB nshort L=0.15 W=0.42 AD=0.0877682 AS=0.0567 PD=0.816449 PS=0.69 NRD=34.284 NRS=22.848 m=1 r=2.8 sa=75000.6 sb=75000.7 a=0.063 p=1.14 mult=1 $X=995 $Y=375 $D=9
M2 X 8 VGND VNB nshort L=0.15 W=0.65 AD=0.182 AS=0.135832 PD=1.86 PS=1.26355 NRD=0 NRS=0 m=1 r=4.33333 sa=75000.8 sb=75000.2 a=0.0975 p=1.6 mult=1 $X=1535 $Y=235 $D=9
M3 8 A VPWR VPB phighvt L=0.15 W=0.42 AD=0.0567 AS=0.1176 PD=0.69 PS=1.4 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75001.4 a=0.063 p=1.14 mult=1 $X=575 $Y=1855 $D=89
M4 VPWR B 8 VPB phighvt L=0.15 W=0.42 AD=0.0985225 AS=0.0567 PD=0.822254 PS=0.69 NRD=55.1009 NRS=0 m=1 r=2.8 sa=75000.6 sb=75000.9 a=0.063 p=1.14 mult=1 $X=995 $Y=1855 $D=89
M5 X 8 VPWR VPB phighvt L=0.15 W=1 AD=0.475 AS=0.234577 PD=2.95 PS=1.95775 NRD=18.715 NRS=0 m=1 r=6.66667 sa=75000.6 sb=75000.4 a=0.15 p=2.3 mult=1 $X=1535 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_31 1 2
** N=2 EP=2 IP=4 FDC=2
*.SEEDPROM
X0 1 2 ICV_3 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__dlclkp_1 VNB VPB CLK GATE VPWR GCLK VGND
** N=111 EP=7 IP=0 FDC=20
*.SEEDPROM
M0 VGND CLK 9 VNB nshort L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75000.6 a=0.063 p=1.14 mult=1 $X=395 $Y=235 $D=9
M1 8 9 VGND VNB nshort L=0.15 W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 m=1 r=2.8 sa=75000.6 sb=75000.2 a=0.063 p=1.14 mult=1 $X=815 $Y=235 $D=9
M2 15 GATE VGND VNB nshort L=0.15 W=0.42 AD=0.117125 AS=0.1281 PD=1.085 PS=1.45 NRD=63.96 NRS=11.424 m=1 r=2.8 sa=75000.2 sb=75000.6 a=0.063 p=1.14 mult=1 $X=1830 $Y=595 $D=9
M3 11 9 15 VNB nshort L=0.15 W=0.42 AD=0.123615 AS=0.117125 PD=1.13037 PS=1.085 NRD=81.42 NRS=63.96 m=1 r=2.8 sa=75000.4 sb=75001.4 a=0.063 p=1.14 mult=1 $X=2380 $Y=330 $D=9
M4 16 8 11 VNB nshort L=0.15 W=0.39 AD=0.0646389 AS=0.114785 PD=0.717407 PS=1.04963 NRD=34.068 NRS=3.072 m=1 r=2.6 sa=75000.9 sb=75001.2 a=0.0585 p=1.08 mult=1 $X=3105 $Y=235 $D=9
M5 VGND 10 16 VNB nshort L=0.15 W=0.42 AD=0.0927336 AS=0.0696111 PD=0.816449 PS=0.772593 NRD=32.856 NRS=31.632 m=1 r=2.8 sa=75001.2 sb=75000.7 a=0.063 p=1.14 mult=1 $X=3580 $Y=235 $D=9
M6 10 11 VGND VNB nshort L=0.15 W=0.65 AD=0.169 AS=0.143516 PD=1.82 PS=1.26355 NRD=0 NRS=0 m=1 r=4.33333 sa=75001.2 sb=75000.2 a=0.0975 p=1.6 mult=1 $X=4120 $Y=235 $D=9
M7 17 10 12 VNB nshort L=0.15 W=0.42 AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 m=1 r=2.8 sa=75000.2 sb=75001 a=0.063 p=1.14 mult=1 $X=5060 $Y=235 $D=9
M8 VGND CLK 17 VNB nshort L=0.15 W=0.42 AD=0.0761495 AS=0.0441 PD=0.765421 PS=0.63 NRD=12.852 NRS=14.28 m=1 r=2.8 sa=75000.5 sb=75000.7 a=0.063 p=1.14 mult=1 $X=5420 $Y=235 $D=9
M9 GCLK 12 VGND VNB nshort L=0.15 W=0.65 AD=0.169 AS=0.11785 PD=1.82 PS=1.18458 NRD=0 NRS=0 m=1 r=4.33333 sa=75000.7 sb=75000.2 a=0.0975 p=1.6 mult=1 $X=5895 $Y=235 $D=9
M10 VPWR CLK 9 VPB phighvt L=0.15 W=0.64 AD=0.0864 AS=0.1664 PD=0.91 PS=1.8 NRD=0 NRS=0 m=1 r=4.26667 sa=75000.2 sb=75000.6 a=0.096 p=1.58 mult=1 $X=395 $Y=1815 $D=89
M11 8 9 VPWR VPB phighvt L=0.15 W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 m=1 r=4.26667 sa=75000.6 sb=75000.2 a=0.096 p=1.58 mult=1 $X=815 $Y=1815 $D=89
M12 13 GATE VPWR VPB phighvt L=0.15 W=0.64 AD=0.115623 AS=0.1664 PD=1.16528 PS=1.8 NRD=38.6711 NRS=0 m=1 r=4.26667 sa=75000.2 sb=75001.1 a=0.096 p=1.58 mult=1 $X=1755 $Y=1845 $D=89
M13 11 8 13 VPB phighvt L=0.15 W=0.42 AD=0.0987 AS=0.0758774 PD=0.89 PS=0.764717 NRD=56.2829 NRS=58.9227 m=1 r=2.8 sa=75000.7 sb=75001.2 a=0.063 p=1.14 mult=1 $X=2230 $Y=2065 $D=89
M14 14 9 11 VPB phighvt L=0.15 W=0.42 AD=0.0441 AS=0.0987 PD=0.63 PS=0.89 NRD=23.443 NRS=32.8202 m=1 r=2.8 sa=75001.3 sb=75000.5 a=0.063 p=1.14 mult=1 $X=2850 $Y=2065 $D=89
M15 VPWR 10 14 VPB phighvt L=0.15 W=0.42 AD=0.1092 AS=0.0441 PD=1.36 PS=0.63 NRD=0 NRS=23.443 m=1 r=2.8 sa=75001.6 sb=75000.2 a=0.063 p=1.14 mult=1 $X=3210 $Y=2065 $D=89
M16 VPWR 11 10 VPB phighvt L=0.15 W=1 AD=0.181707 AS=0.27 PD=1.61585 PS=2.54 NRD=1.9503 NRS=0 m=1 r=6.66667 sa=75000.2 sb=75001.3 a=0.15 p=2.3 mult=1 $X=4160 $Y=1485 $D=89
M17 12 10 VPWR VPB phighvt L=0.15 W=0.64 AD=0.2032 AS=0.116293 PD=1.275 PS=1.03415 NRD=75.4116 NRS=10.7562 m=1 r=4.26667 sa=75000.7 sb=75001.4 a=0.096 p=1.58 mult=1 $X=4635 $Y=1845 $D=89
M18 VPWR CLK 12 VPB phighvt L=0.15 W=0.64 AD=0.116293 AS=0.2032 PD=1.03415 PS=1.275 NRD=15.3857 NRS=33.8446 m=1 r=4.26667 sa=75001.5 sb=75000.7 a=0.096 p=1.58 mult=1 $X=5420 $Y=1845 $D=89
M19 GCLK 12 VPWR VPB phighvt L=0.15 W=1 AD=0.26 AS=0.181707 PD=2.52 PS=1.61585 NRD=0 NRS=0 m=1 r=6.66667 sa=75001.3 sb=75000.2 a=0.15 p=2.3 mult=1 $X=5895 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_32 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_33 1 2
** N=2 EP=2 IP=4 FDC=6
*.SEEDPROM
X0 1 2 ICV_10 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 ICV_11 $T=3220 0 0 0 $X=3030 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_34 1 2
** N=2 EP=2 IP=4 FDC=12
*.SEEDPROM
X0 1 2 ICV_33 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 ICV_33 $T=14260 0 0 0 $X=14070 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_35 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=24
*.SEEDPROM
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__dfxtp_1 $T=920 0 0 0 $X=730 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_36 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=26
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__dfxtp_1 $T=2760 0 0 0 $X=2570 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_37 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=24
*.SEEDPROM
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__dfxtp_1 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_38 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=14 FDC=48
*.SEEDPROM
X0 1 2 3 4 2 5 1 sky130_fd_sc_hd__dfxtp_1 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 6 7 2 8 1 sky130_fd_sc_hd__dfxtp_1 $T=7360 0 0 0 $X=7170 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_39 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=12
*.SEEDPROM
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__ebufn_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_40 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=14
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=4140 0 0 0 $X=3950 $Y=-240
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__ebufn_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_41 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=26
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=7360 0 0 0 $X=7170 $Y=-240
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__dfxtp_1 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_42 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=24
*.SEEDPROM
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__dfxtp_1 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_43 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=26
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=7360 0 0 0 $X=7170 $Y=-240
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__dfxtp_1 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_44 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=24
*.SEEDPROM
X1 1 2 3 4 5 6 7 8 ICV_30 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_45 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=14
*.SEEDPROM
X0 1 2 ICV_3 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__ebufn_2 $T=2300 0 0 0 $X=2110 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_46 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=14 FDC=44
*.SEEDPROM
X0 1 2 3 4 2 5 1 sky130_fd_sc_hd__dfxtp_1 $T=6440 0 0 0 $X=6250 $Y=-240
X1 1 2 8 6 2 7 1 sky130_fd_sc_hd__dlclkp_1 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_47 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=26
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__dfxtp_1 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_48 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=12
*.SEEDPROM
X0 1 2 3 4 2 5 1 sky130_fd_sc_hd__ebufn_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_49 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=38
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 6 7 8 3 4 5 ICV_13 $T=2760 0 0 0 $X=2570 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_50 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=38
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 6 7 8 3 4 5 ICV_13 $T=3680 0 0 0 $X=3490 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_51 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=14 FDC=36
*.SEEDPROM
X0 1 2 3 4 2 5 1 sky130_fd_sc_hd__ebufn_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 6 7 2 8 1 sky130_fd_sc_hd__dfxtp_1 $T=4140 0 0 0 $X=3950 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_52 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=14
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=4140 0 0 0 $X=3950 $Y=-240
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__ebufn_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_53 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=14
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__ebufn_2 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_54 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__clkbuf_16 VNB VPB A VPWR X VGND
** N=276 EP=6 IP=0 FDC=40
*.SEEDPROM
M0 7 A VGND VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75008.4 a=0.063 p=1.14 mult=1 $X=400 $Y=235 $D=9
M1 VGND A 7 VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75000.6 sb=75007.9 a=0.063 p=1.14 mult=1 $X=830 $Y=235 $D=9
M2 7 A VGND VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75001.1 sb=75007.5 a=0.063 p=1.14 mult=1 $X=1260 $Y=235 $D=9
M3 VGND A 7 VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75001.5 sb=75007.1 a=0.063 p=1.14 mult=1 $X=1690 $Y=235 $D=9
M4 X 7 VGND VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75001.9 sb=75006.6 a=0.063 p=1.14 mult=1 $X=2120 $Y=235 $D=9
M5 VGND 7 X VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75002.3 sb=75006.2 a=0.063 p=1.14 mult=1 $X=2550 $Y=235 $D=9
M6 X 7 VGND VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75002.8 sb=75005.8 a=0.063 p=1.14 mult=1 $X=2980 $Y=235 $D=9
M7 VGND 7 X VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75003.2 sb=75005.3 a=0.063 p=1.14 mult=1 $X=3410 $Y=235 $D=9
M8 X 7 VGND VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75003.6 sb=75004.9 a=0.063 p=1.14 mult=1 $X=3840 $Y=235 $D=9
M9 VGND 7 X VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75004.1 sb=75004.5 a=0.063 p=1.14 mult=1 $X=4270 $Y=235 $D=9
M10 X 7 VGND VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75004.5 sb=75004.1 a=0.063 p=1.14 mult=1 $X=4700 $Y=235 $D=9
M11 VGND 7 X VNB nshort L=0.15 W=0.42 AD=0.05775 AS=0.0588 PD=0.695 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75004.9 sb=75003.6 a=0.063 p=1.14 mult=1 $X=5130 $Y=235 $D=9
M12 X 7 VGND VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.05775 PD=0.7 PS=0.695 NRD=0 NRS=0 m=1 r=2.8 sa=75005.3 sb=75003.2 a=0.063 p=1.14 mult=1 $X=5555 $Y=235 $D=9
M13 VGND 7 X VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75005.8 sb=75002.8 a=0.063 p=1.14 mult=1 $X=5985 $Y=235 $D=9
M14 X 7 VGND VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75006.2 sb=75002.3 a=0.063 p=1.14 mult=1 $X=6415 $Y=235 $D=9
M15 VGND 7 X VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75006.6 sb=75001.9 a=0.063 p=1.14 mult=1 $X=6845 $Y=235 $D=9
M16 X 7 VGND VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75007.1 sb=75001.5 a=0.063 p=1.14 mult=1 $X=7275 $Y=235 $D=9
M17 VGND 7 X VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75007.5 sb=75001.1 a=0.063 p=1.14 mult=1 $X=7705 $Y=235 $D=9
M18 X 7 VGND VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75007.9 sb=75000.6 a=0.063 p=1.14 mult=1 $X=8135 $Y=235 $D=9
M19 VGND 7 X VNB nshort L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75008.4 sb=75000.2 a=0.063 p=1.14 mult=1 $X=8565 $Y=235 $D=9
M20 7 A VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=6.66667 sa=75000.2 sb=75008.4 a=0.15 p=2.3 mult=1 $X=400 $Y=1485 $D=89
M21 VPWR A 7 VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75000.6 sb=75007.9 a=0.15 p=2.3 mult=1 $X=830 $Y=1485 $D=89
M22 7 A VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75001 sb=75007.5 a=0.15 p=2.3 mult=1 $X=1260 $Y=1485 $D=89
M23 VPWR A 7 VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75001.5 sb=75007.1 a=0.15 p=2.3 mult=1 $X=1690 $Y=1485 $D=89
M24 X 7 VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75001.9 sb=75006.6 a=0.15 p=2.3 mult=1 $X=2120 $Y=1485 $D=89
M25 VPWR 7 X VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75002.3 sb=75006.2 a=0.15 p=2.3 mult=1 $X=2550 $Y=1485 $D=89
M26 X 7 VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75002.8 sb=75005.8 a=0.15 p=2.3 mult=1 $X=2980 $Y=1485 $D=89
M27 VPWR 7 X VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75003.2 sb=75005.3 a=0.15 p=2.3 mult=1 $X=3410 $Y=1485 $D=89
M28 X 7 VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75003.6 sb=75004.9 a=0.15 p=2.3 mult=1 $X=3840 $Y=1485 $D=89
M29 VPWR 7 X VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75004.1 sb=75004.5 a=0.15 p=2.3 mult=1 $X=4270 $Y=1485 $D=89
M30 X 7 VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75004.5 sb=75004.1 a=0.15 p=2.3 mult=1 $X=4700 $Y=1485 $D=89
M31 VPWR 7 X VPB phighvt L=0.15 W=1 AD=0.1375 AS=0.14 PD=1.275 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75004.9 sb=75003.6 a=0.15 p=2.3 mult=1 $X=5130 $Y=1485 $D=89
M32 X 7 VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.1375 PD=1.28 PS=1.275 NRD=0 NRS=0 m=1 r=6.66667 sa=75005.3 sb=75003.2 a=0.15 p=2.3 mult=1 $X=5555 $Y=1485 $D=89
M33 VPWR 7 X VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75005.8 sb=75002.8 a=0.15 p=2.3 mult=1 $X=5985 $Y=1485 $D=89
M34 X 7 VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75006.2 sb=75002.3 a=0.15 p=2.3 mult=1 $X=6415 $Y=1485 $D=89
M35 VPWR 7 X VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75006.6 sb=75001.9 a=0.15 p=2.3 mult=1 $X=6845 $Y=1485 $D=89
M36 X 7 VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75007.1 sb=75001.5 a=0.15 p=2.3 mult=1 $X=7275 $Y=1485 $D=89
M37 VPWR 7 X VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75007.5 sb=75001 a=0.15 p=2.3 mult=1 $X=7705 $Y=1485 $D=89
M38 X 7 VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75007.9 sb=75000.6 a=0.15 p=2.3 mult=1 $X=8135 $Y=1485 $D=89
M39 VPWR 7 X VPB phighvt L=0.15 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75008.4 sb=75000.2 a=0.15 p=2.3 mult=1 $X=8565 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_55 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
** N=1765 EP=320 IP=16115 FDC=47453
X0 1 2 Dpar a=2090.87 p=1485.04 m=1 $[nwdiode] $X=5330 $Y=444665 $D=191
X1 1 2 Dpar a=2091.12 p=1484.74 m=1 $[nwdiode] $X=5330 $Y=450105 $D=191
X2 1 2 Dpar a=2090.47 p=1485.54 m=1 $[nwdiode] $X=5330 $Y=455545 $D=191
X3 1 2 Dpar a=2090.87 p=1485.04 m=1 $[nwdiode] $X=5330 $Y=460985 $D=191
X4 1 2 Dpar a=2090.95 p=1484.94 m=1 $[nwdiode] $X=5330 $Y=466425 $D=191
X5 1 2 Dpar a=2090.55 p=1485.44 m=1 $[nwdiode] $X=5330 $Y=471865 $D=191
X6 1 2 Dpar a=2090.63 p=1485.34 m=1 $[nwdiode] $X=5330 $Y=477305 $D=191
X7 1 2 Dpar a=2091.2 p=1484.64 m=1 $[nwdiode] $X=5330 $Y=482745 $D=191
X8 1 2 Dpar a=2090.47 p=1485.54 m=1 $[nwdiode] $X=5330 $Y=488185 $D=191
X9 1 2 Dpar a=2090.79 p=1485.14 m=1 $[nwdiode] $X=5330 $Y=493625 $D=191
X10 1 2 Dpar a=2091.12 p=1484.74 m=1 $[nwdiode] $X=5330 $Y=499065 $D=191
X11 1 2 Dpar a=2091.77 p=1483.94 m=1 $[nwdiode] $X=5330 $Y=504505 $D=191
X12 1 2 Dpar a=2091.77 p=1483.94 m=1 $[nwdiode] $X=5330 $Y=509945 $D=191
X13 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 443360 0 0 $X=5330 $Y=443120
X14 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 514080 1 0 $X=5330 $Y=511120
X15 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=14260 492320 1 0 $X=14070 $Y=489360
X16 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=18400 454240 1 0 $X=18210 $Y=451280
X17 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=18400 481440 1 0 $X=18210 $Y=478480
X18 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=28980 448800 0 0 $X=28790 $Y=448560
X19 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=48300 454240 1 0 $X=48110 $Y=451280
X20 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=62100 448800 0 0 $X=61910 $Y=448560
X21 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=81880 465120 1 0 $X=81690 $Y=462160
X22 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=98440 508640 1 0 $X=98250 $Y=505680
X23 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=100740 492320 0 0 $X=100550 $Y=492080
X24 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=110400 481440 0 0 $X=110210 $Y=481200
X25 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=130640 470560 1 0 $X=130450 $Y=467600
X26 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=134320 454240 0 0 $X=134130 $Y=454000
X27 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=139380 465120 0 0 $X=139190 $Y=464880
X28 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=177560 470560 1 0 $X=177370 $Y=467600
X29 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=182620 465120 1 0 $X=182430 $Y=462160
X30 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=189520 508640 0 0 $X=189330 $Y=508400
X31 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=196420 476000 1 0 $X=196230 $Y=473040
X32 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=198720 470560 0 0 $X=198530 $Y=470320
X33 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=200560 497760 0 0 $X=200370 $Y=497520
X34 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=209300 459680 1 0 $X=209110 $Y=456720
X35 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=212520 448800 1 0 $X=212330 $Y=445840
X36 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=214820 470560 1 0 $X=214630 $Y=467600
X37 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=214820 492320 1 0 $X=214630 $Y=489360
X38 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=265420 459680 1 0 $X=265230 $Y=456720
X39 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=265420 481440 1 0 $X=265230 $Y=478480
X40 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=279680 443360 0 0 $X=279490 $Y=443120
X41 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=295780 454240 0 0 $X=295590 $Y=454000
X42 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=299000 448800 1 0 $X=298810 $Y=445840
X43 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=303140 497760 0 0 $X=302950 $Y=497520
X44 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=322920 465120 1 0 $X=322730 $Y=462160
X45 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=327060 508640 1 0 $X=326870 $Y=505680
X46 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=328900 465120 1 0 $X=328710 $Y=462160
X47 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=328900 492320 1 0 $X=328710 $Y=489360
X48 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=345000 481440 1 0 $X=344810 $Y=478480
X49 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350060 497760 0 0 $X=349870 $Y=497520
X50 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=362480 514080 1 0 $X=362290 $Y=511120
X51 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=411240 486880 1 0 $X=411050 $Y=483920
X52 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=421360 454240 1 0 $X=421170 $Y=451280
X53 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=456320 454240 0 0 $X=456130 $Y=454000
X54 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=481160 492320 0 0 $X=480970 $Y=492080
X55 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=490820 514080 1 0 $X=490630 $Y=511120
X56 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=506000 486880 1 0 $X=505810 $Y=483920
X57 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=520260 443360 0 0 $X=520070 $Y=443120
X58 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=525320 497760 1 0 $X=525130 $Y=494800
X59 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=533600 476000 1 0 $X=533410 $Y=473040
X60 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=539120 508640 0 0 $X=538930 $Y=508400
X61 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=541880 465120 1 0 $X=541690 $Y=462160
X62 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=549240 486880 1 0 $X=549050 $Y=483920
X63 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=557520 486880 1 0 $X=557330 $Y=483920
X64 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=559360 443360 0 0 $X=559170 $Y=443120
X65 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=571320 470560 0 0 $X=571130 $Y=470320
X66 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=579600 465120 1 0 $X=579410 $Y=462160
X67 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=579600 486880 0 0 $X=579410 $Y=486640
X68 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=581440 497760 1 0 $X=581250 $Y=494800
X69 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=607660 476000 1 0 $X=607470 $Y=473040
X70 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=615940 492320 1 0 $X=615750 $Y=489360
X71 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=623300 443360 0 0 $X=623110 $Y=443120
X72 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=629280 459680 1 0 $X=629090 $Y=456720
X73 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=637560 459680 1 0 $X=637370 $Y=456720
X74 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=651360 486880 0 0 $X=651170 $Y=486640
X75 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=656880 476000 0 0 $X=656690 $Y=475760
X76 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=662400 508640 0 0 $X=662210 $Y=508400
X77 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=665620 508640 1 0 $X=665430 $Y=505680
X78 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=667920 448800 0 0 $X=667730 $Y=448560
X79 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=674820 470560 1 0 $X=674630 $Y=467600
X80 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=677580 448800 0 0 $X=677390 $Y=448560
X81 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=677580 492320 0 0 $X=677390 $Y=492080
X82 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=691840 508640 1 0 $X=691650 $Y=505680
X83 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=701040 459680 1 0 $X=700850 $Y=456720
X84 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=701040 476000 1 0 $X=700850 $Y=473040
X85 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=733700 465120 0 0 $X=733510 $Y=464880
X86 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=733700 481440 0 0 $X=733510 $Y=481200
X87 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=733700 497760 0 0 $X=733510 $Y=497520
X88 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=733700 503200 0 0 $X=733510 $Y=502960
X89 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 443360 1 180 $X=742710 $Y=443120
X90 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 514080 0 180 $X=742710 $Y=511120
X91 1 2 ICV_1 $T=5520 508640 1 0 $X=5330 $Y=505680
X92 1 2 ICV_1 $T=744280 448800 0 180 $X=742710 $Y=445840
X93 1 2 ICV_1 $T=744280 465120 0 180 $X=742710 $Y=462160
X94 1 2 ICV_1 $T=744280 492320 0 180 $X=742710 $Y=489360
X95 1 2 ICV_1 $T=744280 508640 0 180 $X=742710 $Y=505680
X96 1 2 ICV_2 $T=5520 448800 1 0 $X=5330 $Y=445840
X97 1 2 ICV_2 $T=5520 459680 1 0 $X=5330 $Y=456720
X98 1 2 ICV_2 $T=5520 470560 1 0 $X=5330 $Y=467600
X99 1 2 ICV_2 $T=5520 486880 1 0 $X=5330 $Y=483920
X100 1 2 ICV_2 $T=5520 497760 1 0 $X=5330 $Y=494800
X101 1 2 ICV_2 $T=744280 454240 0 180 $X=742710 $Y=451280
X102 1 2 ICV_2 $T=744280 470560 0 180 $X=742710 $Y=467600
X103 1 2 ICV_2 $T=744280 481440 0 180 $X=742710 $Y=478480
X104 1 2 ICV_2 $T=744280 497760 0 180 $X=742710 $Y=494800
X246 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=6900 476000 1 0 $X=6710 $Y=473040
X247 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=6900 486880 1 0 $X=6710 $Y=483920
X248 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=12420 508640 0 0 $X=12230 $Y=508400
X249 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=13800 443360 0 0 $X=13610 $Y=443120
X250 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 503200 1 0 $X=17750 $Y=500240
X251 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=24380 492320 0 0 $X=24190 $Y=492080
X252 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=34040 448800 0 0 $X=33850 $Y=448560
X253 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=39560 492320 1 0 $X=39370 $Y=489360
X254 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=61640 448800 1 0 $X=61450 $Y=445840
X255 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=69920 448800 1 0 $X=69730 $Y=445840
X256 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=76360 497760 1 0 $X=76170 $Y=494800
X257 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=87860 497760 0 0 $X=87670 $Y=497520
X258 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=95220 476000 1 0 $X=95030 $Y=473040
X259 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=137080 481440 0 0 $X=136890 $Y=481200
X260 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=146280 459680 0 0 $X=146090 $Y=459440
X261 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=210680 448800 0 0 $X=210490 $Y=448560
X262 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=228160 470560 0 0 $X=227970 $Y=470320
X263 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=234600 459680 1 0 $X=234410 $Y=456720
X264 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=242420 503200 1 0 $X=242230 $Y=500240
X265 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=248860 454240 0 0 $X=248670 $Y=454000
X266 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=248860 481440 1 0 $X=248670 $Y=478480
X267 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=252080 459680 0 0 $X=251890 $Y=459440
X268 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=268180 476000 0 0 $X=267990 $Y=475760
X269 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=280140 481440 1 0 $X=279950 $Y=478480
X270 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=300840 481440 1 0 $X=300650 $Y=478480
X271 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=328900 497760 0 0 $X=328710 $Y=497520
X272 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=380880 497760 1 0 $X=380690 $Y=494800
X273 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=389160 476000 1 0 $X=388970 $Y=473040
X274 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=396520 454240 0 0 $X=396330 $Y=454000
X275 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=420440 470560 1 0 $X=420250 $Y=467600
X276 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=424580 459680 0 0 $X=424390 $Y=459440
X277 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=480700 481440 0 0 $X=480510 $Y=481200
X278 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=491740 486880 0 0 $X=491550 $Y=486640
X279 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=493580 476000 0 0 $X=493390 $Y=475760
X280 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=525320 465120 1 0 $X=525130 $Y=462160
X281 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=530380 443360 0 0 $X=530190 $Y=443120
X282 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=536820 492320 0 0 $X=536630 $Y=492080
X283 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=543260 481440 0 0 $X=543070 $Y=481200
X284 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=546480 448800 0 0 $X=546290 $Y=448560
X285 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=560740 481440 1 0 $X=560550 $Y=478480
X286 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=592940 508640 0 0 $X=592750 $Y=508400
X287 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=595240 465120 0 0 $X=595050 $Y=464880
X288 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=642620 508640 0 0 $X=642430 $Y=508400
X289 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=659180 454240 1 0 $X=658990 $Y=451280
X290 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=665620 448800 1 0 $X=665430 $Y=445840
X291 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=677120 454240 1 0 $X=676930 $Y=451280
X292 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=677120 497760 1 0 $X=676930 $Y=494800
X293 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=691380 476000 1 0 $X=691190 $Y=473040
X294 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=733240 470560 0 0 $X=733050 $Y=470320
X295 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=733240 476000 0 0 $X=733050 $Y=475760
X296 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=733240 492320 0 0 $X=733050 $Y=492080
X297 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 448800 0 0 $X=740870 $Y=448560
X298 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 454240 0 0 $X=740870 $Y=454000
X299 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 465120 0 0 $X=740870 $Y=464880
X300 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 470560 0 0 $X=740870 $Y=470320
X301 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 476000 0 0 $X=740870 $Y=475760
X302 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 481440 0 0 $X=740870 $Y=481200
X303 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 486880 0 0 $X=740870 $Y=486640
X304 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 492320 0 0 $X=740870 $Y=492080
X305 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 497760 0 0 $X=740870 $Y=497520
X306 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 503200 0 0 $X=740870 $Y=502960
X307 1 2 ICV_3 $T=16100 470560 1 0 $X=15910 $Y=467600
X308 1 2 ICV_3 $T=17480 486880 1 0 $X=17290 $Y=483920
X309 1 2 ICV_3 $T=36340 486880 1 0 $X=36150 $Y=483920
X310 1 2 ICV_3 $T=73600 459680 1 0 $X=73410 $Y=456720
X311 1 2 ICV_3 $T=73600 492320 1 0 $X=73410 $Y=489360
X312 1 2 ICV_3 $T=104420 465120 1 0 $X=104230 $Y=462160
X313 1 2 ICV_3 $T=134780 508640 0 0 $X=134590 $Y=508400
X314 1 2 ICV_3 $T=161000 448800 0 0 $X=160810 $Y=448560
X315 1 2 ICV_3 $T=195500 448800 0 0 $X=195310 $Y=448560
X316 1 2 ICV_3 $T=206080 465120 1 0 $X=205890 $Y=462160
X317 1 2 ICV_3 $T=219420 508640 0 0 $X=219230 $Y=508400
X318 1 2 ICV_3 $T=241960 465120 1 0 $X=241770 $Y=462160
X319 1 2 ICV_3 $T=255760 476000 0 0 $X=255570 $Y=475760
X320 1 2 ICV_3 $T=283820 486880 0 0 $X=283630 $Y=486640
X321 1 2 ICV_3 $T=298080 465120 1 0 $X=297890 $Y=462160
X322 1 2 ICV_3 $T=322000 476000 1 0 $X=321810 $Y=473040
X323 1 2 ICV_3 $T=344080 476000 1 0 $X=343890 $Y=473040
X324 1 2 ICV_3 $T=363860 465120 1 0 $X=363670 $Y=462160
X325 1 2 ICV_3 $T=387320 481440 0 0 $X=387130 $Y=481200
X326 1 2 ICV_3 $T=399740 481440 1 0 $X=399550 $Y=478480
X327 1 2 ICV_3 $T=406180 508640 0 0 $X=405990 $Y=508400
X328 1 2 ICV_3 $T=410320 481440 1 0 $X=410130 $Y=478480
X329 1 2 ICV_3 $T=424120 443360 0 0 $X=423930 $Y=443120
X330 1 2 ICV_3 $T=452180 492320 0 0 $X=451990 $Y=492080
X331 1 2 ICV_3 $T=459540 476000 0 0 $X=459350 $Y=475760
X332 1 2 ICV_3 $T=459540 514080 1 0 $X=459350 $Y=511120
X333 1 2 ICV_3 $T=481620 470560 1 0 $X=481430 $Y=467600
X334 1 2 ICV_3 $T=497260 486880 1 0 $X=497070 $Y=483920
X335 1 2 ICV_3 $T=523480 514080 1 0 $X=523290 $Y=511120
X336 1 2 ICV_3 $T=548780 497760 0 0 $X=548590 $Y=497520
X337 1 2 ICV_3 $T=578680 459680 1 0 $X=578490 $Y=456720
X338 1 2 ICV_3 $T=603520 481440 0 0 $X=603330 $Y=481200
X339 1 2 ICV_3 $T=606740 465120 1 0 $X=606550 $Y=462160
X340 1 2 ICV_3 $T=623300 497760 0 0 $X=623110 $Y=497520
X341 1 2 ICV_3 $T=643540 476000 0 0 $X=643350 $Y=475760
X342 1 2 ICV_3 $T=662860 465120 1 0 $X=662670 $Y=462160
X343 1 2 ICV_3 $T=665620 486880 1 0 $X=665430 $Y=483920
X344 1 2 ICV_3 $T=718980 448800 1 0 $X=718790 $Y=445840
X345 1 2 ICV_3 $T=740600 508640 0 0 $X=740410 $Y=508400
X346 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=45080 459680 1 0 $X=44890 $Y=456720
X347 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=61180 497760 1 0 $X=60990 $Y=494800
X348 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=73140 454240 1 0 $X=72950 $Y=451280
X349 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=104420 454240 1 0 $X=104230 $Y=451280
X350 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=109940 454240 0 0 $X=109750 $Y=454000
X351 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=126500 459680 0 0 $X=126310 $Y=459440
X352 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=139840 476000 1 0 $X=139650 $Y=473040
X353 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=143060 492320 0 0 $X=142870 $Y=492080
X354 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=168360 448800 1 0 $X=168170 $Y=445840
X355 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=185380 486880 1 0 $X=185190 $Y=483920
X356 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=199180 459680 0 0 $X=198990 $Y=459440
X357 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=202400 503200 0 0 $X=202210 $Y=502960
X358 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=207460 508640 0 0 $X=207270 $Y=508400
X359 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=222640 481440 0 0 $X=222450 $Y=481200
X360 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=230460 465120 0 0 $X=230270 $Y=464880
X361 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=237820 465120 0 0 $X=237630 $Y=464880
X362 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=244720 465120 0 0 $X=244530 $Y=464880
X363 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=250700 448800 0 0 $X=250510 $Y=448560
X364 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=252080 476000 1 0 $X=251890 $Y=473040
X365 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=289340 503200 1 0 $X=289150 $Y=500240
X366 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=300840 486880 1 0 $X=300650 $Y=483920
X367 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=302220 514080 1 0 $X=302030 $Y=511120
X368 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=314640 497760 0 0 $X=314450 $Y=497520
X369 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=314640 503200 0 0 $X=314450 $Y=502960
X370 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=328900 497760 1 0 $X=328710 $Y=494800
X371 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=330740 514080 1 0 $X=330550 $Y=511120
X372 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=339480 470560 0 0 $X=339290 $Y=470320
X373 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=339480 497760 0 0 $X=339290 $Y=497520
X374 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=348220 514080 1 0 $X=348030 $Y=511120
X375 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=363400 476000 1 0 $X=363210 $Y=473040
X376 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=391460 508640 0 0 $X=391270 $Y=508400
X377 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=402960 486880 0 0 $X=402770 $Y=486640
X378 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=409860 492320 1 0 $X=409670 $Y=489360
X379 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=440220 443360 0 0 $X=440030 $Y=443120
X380 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=451720 465120 0 0 $X=451530 $Y=464880
X381 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=454940 508640 0 0 $X=454750 $Y=508400
X382 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=459080 459680 0 0 $X=458890 $Y=459440
X383 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=459080 486880 0 0 $X=458890 $Y=486640
X384 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=476560 514080 1 0 $X=476370 $Y=511120
X385 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=479780 443360 0 0 $X=479590 $Y=443120
X386 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=480700 508640 1 0 $X=480510 $Y=505680
X387 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=489440 486880 1 0 $X=489250 $Y=483920
X388 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=515660 486880 1 0 $X=515470 $Y=483920
X389 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=544640 514080 1 0 $X=544450 $Y=511120
X390 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=550160 481440 1 0 $X=549970 $Y=478480
X391 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=553380 470560 1 0 $X=553190 $Y=467600
X392 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=553380 476000 1 0 $X=553190 $Y=473040
X393 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=567180 508640 0 0 $X=566990 $Y=508400
X394 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=578220 448800 1 0 $X=578030 $Y=445840
X395 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=602600 497760 1 0 $X=602410 $Y=494800
X396 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=603520 465120 0 0 $X=603330 $Y=464880
X397 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=637560 465120 1 0 $X=637370 $Y=462160
X398 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=637560 486880 1 0 $X=637370 $Y=483920
X399 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=639860 503200 0 0 $X=639670 $Y=502960
X400 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=685860 486880 0 0 $X=685670 $Y=486640
X401 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=730020 514080 1 0 $X=729830 $Y=511120
X402 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=740140 459680 1 0 $X=739950 $Y=456720
X403 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=740140 465120 1 0 $X=739950 $Y=462160
X404 1 2 ICV_4 $T=30360 492320 0 0 $X=30170 $Y=492080
X405 1 2 ICV_4 $T=34040 470560 0 0 $X=33850 $Y=470320
X406 1 2 ICV_4 $T=34040 508640 0 0 $X=33850 $Y=508400
X407 1 2 ICV_4 $T=48300 476000 1 0 $X=48110 $Y=473040
X408 1 2 ICV_4 $T=62100 443360 0 0 $X=61910 $Y=443120
X409 1 2 ICV_4 $T=76360 486880 1 0 $X=76170 $Y=483920
X410 1 2 ICV_4 $T=128800 497760 1 0 $X=128610 $Y=494800
X411 1 2 ICV_4 $T=142600 497760 0 0 $X=142410 $Y=497520
X412 1 2 ICV_4 $T=142600 503200 0 0 $X=142410 $Y=502960
X413 1 2 ICV_4 $T=144440 481440 1 0 $X=144250 $Y=478480
X414 1 2 ICV_4 $T=146280 448800 0 0 $X=146090 $Y=448560
X415 1 2 ICV_4 $T=160540 508640 1 0 $X=160350 $Y=505680
X416 1 2 ICV_4 $T=201020 454240 1 0 $X=200830 $Y=451280
X417 1 2 ICV_4 $T=202400 443360 0 0 $X=202210 $Y=443120
X418 1 2 ICV_4 $T=202400 481440 1 0 $X=202210 $Y=478480
X419 1 2 ICV_4 $T=282900 481440 0 0 $X=282710 $Y=481200
X420 1 2 ICV_4 $T=304980 448800 1 0 $X=304790 $Y=445840
X421 1 2 ICV_4 $T=310960 514080 1 0 $X=310770 $Y=511120
X422 1 2 ICV_4 $T=314640 448800 0 0 $X=314450 $Y=448560
X423 1 2 ICV_4 $T=318780 443360 0 0 $X=318590 $Y=443120
X424 1 2 ICV_4 $T=342700 454240 0 0 $X=342510 $Y=454000
X425 1 2 ICV_4 $T=465520 448800 1 0 $X=465330 $Y=445840
X426 1 2 ICV_4 $T=507380 508640 0 0 $X=507190 $Y=508400
X427 1 2 ICV_4 $T=507840 508640 1 0 $X=507650 $Y=505680
X428 1 2 ICV_4 $T=508300 503200 1 0 $X=508110 $Y=500240
X429 1 2 ICV_4 $T=535440 470560 0 0 $X=535250 $Y=470320
X430 1 2 ICV_4 $T=567180 459680 0 0 $X=566990 $Y=459440
X431 1 2 ICV_4 $T=567180 492320 0 0 $X=566990 $Y=492080
X432 1 2 ICV_4 $T=609500 481440 1 0 $X=609310 $Y=478480
X433 1 2 ICV_4 $T=618240 454240 1 0 $X=618050 $Y=451280
X434 1 2 ICV_4 $T=666540 492320 0 0 $X=666350 $Y=492080
X435 1 2 ICV_4 $T=685860 481440 0 0 $X=685670 $Y=481200
X436 1 2 ICV_4 $T=693680 454240 1 0 $X=693490 $Y=451280
X437 1 2 ICV_4 $T=695520 454240 0 0 $X=695330 $Y=454000
X438 1 2 ICV_4 $T=707480 508640 0 0 $X=707290 $Y=508400
X439 1 2 ICV_4 $T=718980 465120 0 0 $X=718790 $Y=464880
X440 1 2 ICV_4 $T=739680 443360 0 0 $X=739490 $Y=443120
X441 1 2 ICV_4 $T=739680 448800 1 0 $X=739490 $Y=445840
X442 1 2 ICV_4 $T=739680 459680 0 0 $X=739490 $Y=459440
X443 1 2 ICV_4 $T=739680 492320 1 0 $X=739490 $Y=489360
X444 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 443360 0 0 $X=6710 $Y=443120
X445 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 497760 1 0 $X=6710 $Y=494800
X446 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 497760 0 0 $X=6710 $Y=497520
X447 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=11960 465120 1 0 $X=11770 $Y=462160
X448 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=21160 454240 0 0 $X=20970 $Y=454000
X449 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=28980 503200 0 0 $X=28790 $Y=502960
X450 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=29900 465120 0 0 $X=29710 $Y=464880
X451 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=34040 503200 0 0 $X=33850 $Y=502960
X452 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=35420 503200 1 0 $X=35230 $Y=500240
X453 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=44160 465120 1 0 $X=43970 $Y=462160
X454 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=47380 448800 0 0 $X=47190 $Y=448560
X455 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=47840 481440 0 0 $X=47650 $Y=481200
X456 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=53820 503200 1 0 $X=53630 $Y=500240
X457 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=57960 476000 0 0 $X=57770 $Y=475760
X458 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=71760 492320 0 0 $X=71570 $Y=492080
X459 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=76360 476000 1 0 $X=76170 $Y=473040
X460 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=78200 508640 0 0 $X=78010 $Y=508400
X461 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=82340 503200 1 0 $X=82150 $Y=500240
X462 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=104420 459680 1 0 $X=104230 $Y=456720
X463 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=112700 508640 0 0 $X=112510 $Y=508400
X464 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=119140 465120 1 0 $X=118950 $Y=462160
X465 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=121900 454240 1 0 $X=121710 $Y=451280
X466 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=142140 508640 0 0 $X=141950 $Y=508400
X467 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=145360 465120 1 0 $X=145170 $Y=462160
X468 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=146280 470560 0 0 $X=146090 $Y=470320
X469 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=155020 508640 1 0 $X=154830 $Y=505680
X470 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=169280 465120 1 0 $X=169090 $Y=462160
X471 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=170200 465120 0 0 $X=170010 $Y=464880
X472 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=173880 470560 1 0 $X=173690 $Y=467600
X473 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=174340 459680 0 0 $X=174150 $Y=459440
X474 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=181700 443360 0 0 $X=181510 $Y=443120
X475 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=203780 470560 1 0 $X=203590 $Y=467600
X476 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=208380 476000 1 0 $X=208190 $Y=473040
X477 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=216660 481440 1 0 $X=216470 $Y=478480
X478 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=224020 470560 1 0 $X=223830 $Y=467600
X479 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=262660 481440 0 0 $X=262470 $Y=481200
X480 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=292560 486880 0 0 $X=292370 $Y=486640
X481 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=310500 470560 0 0 $X=310310 $Y=470320
X482 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=312340 470560 1 0 $X=312150 $Y=467600
X483 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=359260 481440 0 0 $X=359070 $Y=481200
X484 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=362480 465120 0 0 $X=362290 $Y=464880
X485 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=364320 503200 1 0 $X=364130 $Y=500240
X486 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=369380 508640 1 0 $X=369190 $Y=505680
X487 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=370760 508640 0 0 $X=370570 $Y=508400
X488 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=372140 514080 1 0 $X=371950 $Y=511120
X489 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=392380 476000 1 0 $X=392190 $Y=473040
X490 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=394680 470560 0 0 $X=394490 $Y=470320
X491 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=398820 459680 1 0 $X=398630 $Y=456720
X492 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=437000 508640 1 0 $X=436810 $Y=505680
X493 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=442520 503200 0 0 $X=442330 $Y=502960
X494 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=445280 508640 1 0 $X=445090 $Y=505680
X495 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=454940 470560 0 0 $X=454750 $Y=470320
X496 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=457240 481440 1 0 $X=457050 $Y=478480
X497 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=460920 508640 1 0 $X=460730 $Y=505680
X498 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=462760 508640 0 0 $X=462570 $Y=508400
X499 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=468280 459680 0 0 $X=468090 $Y=459440
X500 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=469200 486880 1 0 $X=469010 $Y=483920
X501 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=473340 465120 1 0 $X=473150 $Y=462160
X502 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=476560 492320 1 0 $X=476370 $Y=489360
X503 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=478860 508640 0 0 $X=478670 $Y=508400
X504 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=484840 459680 1 0 $X=484650 $Y=456720
X505 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=488980 481440 1 0 $X=488790 $Y=478480
X506 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=493580 470560 0 0 $X=493390 $Y=470320
X507 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=497260 503200 1 0 $X=497070 $Y=500240
X508 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=519340 492320 0 0 $X=519150 $Y=492080
X509 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=534980 486880 0 0 $X=534790 $Y=486640
X510 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=539120 443360 0 0 $X=538930 $Y=443120
X511 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=543720 503200 1 0 $X=543530 $Y=500240
X512 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=553380 497760 1 0 $X=553190 $Y=494800
X513 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=563040 448800 0 0 $X=562850 $Y=448560
X514 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=563040 503200 0 0 $X=562850 $Y=502960
X515 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=589720 459680 1 0 $X=589530 $Y=456720
X516 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=599840 514080 1 0 $X=599650 $Y=511120
X517 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=604440 503200 0 0 $X=604250 $Y=502960
X518 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=604900 503200 1 0 $X=604710 $Y=500240
X519 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=605360 508640 1 0 $X=605170 $Y=505680
X520 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=625600 492320 1 0 $X=625410 $Y=489360
X521 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=628360 508640 0 0 $X=628170 $Y=508400
X522 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=631580 481440 0 0 $X=631390 $Y=481200
X523 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=633420 492320 1 0 $X=633230 $Y=489360
X524 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=655500 503200 0 0 $X=655310 $Y=502960
X525 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=667460 454240 0 0 $X=667270 $Y=454000
X526 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=672980 476000 1 0 $X=672790 $Y=473040
X527 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=675280 476000 0 0 $X=675090 $Y=475760
X528 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=679420 497760 0 0 $X=679230 $Y=497520
X529 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=687700 465120 0 0 $X=687510 $Y=464880
X530 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=688160 486880 1 0 $X=687970 $Y=483920
X531 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=690460 503200 0 0 $X=690270 $Y=502960
X532 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=698280 492320 0 0 $X=698090 $Y=492080
X533 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=702420 503200 0 0 $X=702230 $Y=502960
X534 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=730020 497760 0 0 $X=729830 $Y=497520
X535 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=730020 503200 0 0 $X=729830 $Y=502960
X536 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=730940 486880 0 0 $X=730750 $Y=486640
X537 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=738760 514080 1 0 $X=738570 $Y=511120
X538 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 508640 0 0 $X=6710 $Y=508400
X539 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=66240 503200 0 0 $X=66050 $Y=502960
X540 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=101200 508640 0 0 $X=101010 $Y=508400
X541 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=111780 503200 0 0 $X=111590 $Y=502960
X542 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=156860 508640 0 0 $X=156670 $Y=508400
X543 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=214360 503200 0 0 $X=214170 $Y=502960
X544 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=272780 486880 1 0 $X=272590 $Y=483920
X545 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=293940 486880 1 0 $X=293750 $Y=483920
X546 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=318780 476000 0 0 $X=318590 $Y=475760
X547 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=321540 508640 1 0 $X=321350 $Y=505680
X548 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=358340 465120 1 0 $X=358150 $Y=462160
X549 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=374900 481440 1 0 $X=374710 $Y=478480
X550 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=385020 470560 0 0 $X=384830 $Y=470320
X551 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=425960 514080 1 0 $X=425770 $Y=511120
X552 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=484380 514080 1 0 $X=484190 $Y=511120
X553 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=564880 508640 1 0 $X=564690 $Y=505680
X554 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=573160 459680 1 0 $X=572970 $Y=456720
X555 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=574540 508640 1 0 $X=574350 $Y=505680
X556 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=588800 486880 0 0 $X=588610 $Y=486640
X557 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=589260 503200 0 0 $X=589070 $Y=502960
X558 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=637100 508640 0 0 $X=636910 $Y=508400
X559 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=637560 481440 1 0 $X=637370 $Y=478480
X560 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=679420 508640 0 0 $X=679230 $Y=508400
X561 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=713920 508640 1 0 $X=713730 $Y=505680
X562 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=715300 497760 1 0 $X=715110 $Y=494800
X563 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=734160 448800 1 0 $X=733970 $Y=445840
X564 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=734160 492320 1 0 $X=733970 $Y=489360
X565 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=734620 459680 1 0 $X=734430 $Y=456720
X566 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=734620 465120 1 0 $X=734430 $Y=462160
X567 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 448800 0 0 $X=735350 $Y=448560
X568 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 454240 0 0 $X=735350 $Y=454000
X569 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 486880 0 0 $X=735350 $Y=486640
X570 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=737380 486880 1 0 $X=737190 $Y=483920
X571 1 2 5 2 12 1 sky130_fd_sc_hd__clkbuf_8 $T=6900 465120 1 0 $X=6710 $Y=462160
X572 1 2 17 2 23 1 sky130_fd_sc_hd__clkbuf_8 $T=14260 508640 0 0 $X=14070 $Y=508400
X573 1 2 36 2 37 1 sky130_fd_sc_hd__clkbuf_8 $T=37260 508640 0 0 $X=37070 $Y=508400
X574 1 2 44 2 48 1 sky130_fd_sc_hd__clkbuf_8 $T=62100 508640 0 0 $X=61910 $Y=508400
X575 1 2 52 2 54 1 sky130_fd_sc_hd__clkbuf_8 $T=81880 508640 0 0 $X=81690 $Y=508400
X576 1 2 63 2 65 1 sky130_fd_sc_hd__clkbuf_8 $T=107640 508640 0 0 $X=107450 $Y=508400
X577 1 2 75 2 76 1 sky130_fd_sc_hd__clkbuf_8 $T=137080 508640 0 0 $X=136890 $Y=508400
X578 1 2 87 2 90 1 sky130_fd_sc_hd__clkbuf_8 $T=151800 508640 0 0 $X=151610 $Y=508400
X579 1 2 105 2 106 1 sky130_fd_sc_hd__clkbuf_8 $T=175260 508640 0 0 $X=175070 $Y=508400
X580 1 2 115 2 114 1 sky130_fd_sc_hd__clkbuf_8 $T=202400 508640 0 0 $X=202210 $Y=508400
X581 1 2 123 2 120 1 sky130_fd_sc_hd__clkbuf_8 $T=221720 508640 0 0 $X=221530 $Y=508400
X582 1 2 131 2 117 1 sky130_fd_sc_hd__clkbuf_8 $T=245180 508640 1 0 $X=244990 $Y=505680
X583 1 2 136 2 121 1 sky130_fd_sc_hd__clkbuf_8 $T=270020 508640 0 0 $X=269830 $Y=508400
X584 1 2 141 2 127 1 sky130_fd_sc_hd__clkbuf_8 $T=292100 503200 1 0 $X=291910 $Y=500240
X585 1 2 147 2 128 1 sky130_fd_sc_hd__clkbuf_8 $T=314180 514080 1 0 $X=313990 $Y=511120
X586 1 2 172 2 126 1 sky130_fd_sc_hd__clkbuf_8 $T=342700 508640 0 0 $X=342510 $Y=508400
X587 1 2 180 2 122 1 sky130_fd_sc_hd__clkbuf_8 $T=355120 514080 1 0 $X=354930 $Y=511120
X588 1 2 191 2 192 1 sky130_fd_sc_hd__clkbuf_8 $T=386400 508640 0 0 $X=386210 $Y=508400
X589 1 2 202 2 203 1 sky130_fd_sc_hd__clkbuf_8 $T=408480 508640 0 0 $X=408290 $Y=508400
X590 1 2 211 2 214 1 sky130_fd_sc_hd__clkbuf_8 $T=438840 508640 0 0 $X=438650 $Y=508400
X591 1 2 220 2 224 1 sky130_fd_sc_hd__clkbuf_8 $T=457700 508640 0 0 $X=457510 $Y=508400
X592 1 2 235 2 238 1 sky130_fd_sc_hd__clkbuf_8 $T=479320 514080 1 0 $X=479130 $Y=511120
X593 1 2 246 2 249 1 sky130_fd_sc_hd__clkbuf_8 $T=505080 514080 1 0 $X=504890 $Y=511120
X594 1 2 254 2 260 1 sky130_fd_sc_hd__clkbuf_8 $T=525780 514080 1 0 $X=525590 $Y=511120
X595 1 2 274 2 276 1 sky130_fd_sc_hd__clkbuf_8 $T=548780 508640 0 0 $X=548590 $Y=508400
X596 1 2 278 2 281 1 sky130_fd_sc_hd__clkbuf_8 $T=569940 508640 0 0 $X=569750 $Y=508400
X597 1 2 282 2 284 1 sky130_fd_sc_hd__clkbuf_8 $T=590640 514080 1 0 $X=590450 $Y=511120
X598 1 2 290 2 291 1 sky130_fd_sc_hd__clkbuf_8 $T=623300 508640 0 0 $X=623110 $Y=508400
X599 1 2 295 2 296 1 sky130_fd_sc_hd__clkbuf_8 $T=644460 508640 0 0 $X=644270 $Y=508400
X600 1 2 302 2 303 1 sky130_fd_sc_hd__clkbuf_8 $T=663780 508640 0 0 $X=663590 $Y=508400
X601 1 2 307 2 309 1 sky130_fd_sc_hd__clkbuf_8 $T=685400 508640 0 0 $X=685210 $Y=508400
X602 1 2 314 2 315 1 sky130_fd_sc_hd__clkbuf_8 $T=710700 508640 0 0 $X=710510 $Y=508400
X603 1 2 318 2 319 1 sky130_fd_sc_hd__clkbuf_8 $T=735540 508640 0 0 $X=735350 $Y=508400
X604 1 2 356 340 2 21 1 sky130_fd_sc_hd__ebufn_2 $T=26220 492320 0 0 $X=26030 $Y=492080
X605 1 2 366 364 2 27 1 sky130_fd_sc_hd__ebufn_2 $T=28520 465120 1 0 $X=28330 $Y=462160
X606 1 2 373 369 2 25 1 sky130_fd_sc_hd__ebufn_2 $T=35880 481440 0 0 $X=35690 $Y=481200
X607 1 2 396 369 2 21 1 sky130_fd_sc_hd__ebufn_2 $T=45540 470560 0 0 $X=45350 $Y=470320
X608 1 2 399 385 2 32 1 sky130_fd_sc_hd__ebufn_2 $T=55200 465120 0 0 $X=55010 $Y=464880
X609 1 2 409 43 2 32 1 sky130_fd_sc_hd__ebufn_2 $T=58420 454240 1 0 $X=58230 $Y=451280
X610 1 2 440 436 2 22 1 sky130_fd_sc_hd__ebufn_2 $T=71300 486880 1 0 $X=71110 $Y=483920
X611 1 2 447 448 2 30 1 sky130_fd_sc_hd__ebufn_2 $T=71760 448800 1 0 $X=71570 $Y=445840
X612 1 2 454 459 2 22 1 sky130_fd_sc_hd__ebufn_2 $T=78200 503200 1 0 $X=78010 $Y=500240
X613 1 2 460 436 2 28 1 sky130_fd_sc_hd__ebufn_2 $T=79120 481440 0 0 $X=78930 $Y=481200
X614 1 2 478 485 2 22 1 sky130_fd_sc_hd__ebufn_2 $T=90160 454240 0 0 $X=89970 $Y=454000
X615 1 2 438 364 2 20 1 sky130_fd_sc_hd__ebufn_2 $T=91540 465120 1 0 $X=91350 $Y=462160
X616 1 2 59 60 2 20 1 sky130_fd_sc_hd__ebufn_2 $T=96140 448800 1 0 $X=95950 $Y=445840
X617 1 2 507 64 2 27 1 sky130_fd_sc_hd__ebufn_2 $T=107180 454240 1 0 $X=106990 $Y=451280
X618 1 2 67 64 2 20 1 sky130_fd_sc_hd__ebufn_2 $T=113620 443360 0 0 $X=113430 $Y=443120
X619 1 2 534 513 2 25 1 sky130_fd_sc_hd__ebufn_2 $T=115000 465120 1 0 $X=114810 $Y=462160
X620 1 2 575 579 2 27 1 sky130_fd_sc_hd__ebufn_2 $T=138920 481440 0 0 $X=138730 $Y=481200
X621 1 2 583 72 2 28 1 sky130_fd_sc_hd__ebufn_2 $T=141220 454240 0 0 $X=141030 $Y=454000
X622 1 2 596 597 2 27 1 sky130_fd_sc_hd__ebufn_2 $T=149500 492320 1 0 $X=149310 $Y=489360
X623 1 2 727 704 2 25 1 sky130_fd_sc_hd__ebufn_2 $T=212520 448800 0 0 $X=212330 $Y=448560
X624 1 2 739 735 2 27 1 sky130_fd_sc_hd__ebufn_2 $T=218500 481440 0 0 $X=218310 $Y=481200
X625 1 2 740 734 2 102 1 sky130_fd_sc_hd__ebufn_2 $T=218960 465120 0 0 $X=218770 $Y=464880
X626 1 2 775 752 2 89 1 sky130_fd_sc_hd__ebufn_2 $T=236440 459680 1 0 $X=236250 $Y=456720
X627 1 2 782 781 2 92 1 sky130_fd_sc_hd__ebufn_2 $T=240580 465120 0 0 $X=240390 $Y=464880
X628 1 2 788 736 2 21 1 sky130_fd_sc_hd__ebufn_2 $T=244720 497760 1 0 $X=244530 $Y=494800
X629 1 2 803 781 2 101 1 sky130_fd_sc_hd__ebufn_2 $T=251160 486880 0 0 $X=250970 $Y=486640
X630 1 2 794 732 2 22 1 sky130_fd_sc_hd__ebufn_2 $T=251160 492320 0 0 $X=250970 $Y=492080
X631 1 2 806 133 2 102 1 sky130_fd_sc_hd__ebufn_2 $T=253460 448800 0 0 $X=253270 $Y=448560
X632 1 2 853 839 2 101 1 sky130_fd_sc_hd__ebufn_2 $T=288420 486880 0 0 $X=288230 $Y=486640
X633 1 2 857 839 2 103 1 sky130_fd_sc_hd__ebufn_2 $T=289800 486880 1 0 $X=289610 $Y=483920
X634 1 2 867 847 2 103 1 sky130_fd_sc_hd__ebufn_2 $T=300840 454240 1 0 $X=300650 $Y=451280
X635 1 2 874 876 2 92 1 sky130_fd_sc_hd__ebufn_2 $T=303600 486880 1 0 $X=303410 $Y=483920
X636 1 2 885 903 2 152 1 sky130_fd_sc_hd__ebufn_2 $T=317400 503200 0 0 $X=317210 $Y=502960
X637 1 2 939 945 2 167 1 sky130_fd_sc_hd__ebufn_2 $T=338100 465120 0 0 $X=337910 $Y=464880
X638 1 2 173 175 2 167 1 sky130_fd_sc_hd__ebufn_2 $T=342700 448800 0 0 $X=342510 $Y=448560
X639 1 2 953 925 2 167 1 sky130_fd_sc_hd__ebufn_2 $T=347760 508640 0 0 $X=347570 $Y=508400
X640 1 2 969 972 2 164 1 sky130_fd_sc_hd__ebufn_2 $T=350980 514080 1 0 $X=350790 $Y=511120
X641 1 2 973 945 2 164 1 sky130_fd_sc_hd__ebufn_2 $T=351900 465120 1 0 $X=351710 $Y=462160
X642 1 2 976 174 2 170 1 sky130_fd_sc_hd__ebufn_2 $T=354660 443360 0 0 $X=354470 $Y=443120
X643 1 2 998 1000 2 164 1 sky130_fd_sc_hd__ebufn_2 $T=366160 465120 0 0 $X=365970 $Y=464880
X644 1 2 1006 972 2 157 1 sky130_fd_sc_hd__ebufn_2 $T=368000 503200 1 0 $X=367810 $Y=500240
X645 1 2 1015 1014 2 157 1 sky130_fd_sc_hd__ebufn_2 $T=371680 476000 0 0 $X=371490 $Y=475760
X646 1 2 1028 994 2 157 1 sky130_fd_sc_hd__ebufn_2 $T=377200 492320 0 0 $X=377010 $Y=492080
X647 1 2 1035 1014 2 164 1 sky130_fd_sc_hd__ebufn_2 $T=380880 470560 0 0 $X=380690 $Y=470320
X648 1 2 1047 1046 2 170 1 sky130_fd_sc_hd__ebufn_2 $T=386860 454240 1 0 $X=386670 $Y=451280
X649 1 2 1055 1051 2 155 1 sky130_fd_sc_hd__ebufn_2 $T=390540 470560 0 0 $X=390350 $Y=470320
X650 1 2 1062 1065 2 152 1 sky130_fd_sc_hd__ebufn_2 $T=394220 497760 0 0 $X=394030 $Y=497520
X651 1 2 1063 1065 2 164 1 sky130_fd_sc_hd__ebufn_2 $T=394220 508640 0 0 $X=394030 $Y=508400
X652 1 2 1083 1065 2 155 1 sky130_fd_sc_hd__ebufn_2 $T=403420 497760 1 0 $X=403230 $Y=494800
X653 1 2 1090 1080 2 155 1 sky130_fd_sc_hd__ebufn_2 $T=405720 476000 1 0 $X=405530 $Y=473040
X654 1 2 1088 204 2 164 1 sky130_fd_sc_hd__ebufn_2 $T=419980 443360 0 0 $X=419790 $Y=443120
X655 1 2 1112 1095 2 151 1 sky130_fd_sc_hd__ebufn_2 $T=419980 486880 0 0 $X=419790 $Y=486640
X656 1 2 1139 1107 2 152 1 sky130_fd_sc_hd__ebufn_2 $T=427800 459680 1 0 $X=427610 $Y=456720
X657 1 2 1145 1142 2 164 1 sky130_fd_sc_hd__ebufn_2 $T=427800 476000 0 0 $X=427610 $Y=475760
X658 1 2 1146 1143 2 170 1 sky130_fd_sc_hd__ebufn_2 $T=427800 481440 0 0 $X=427610 $Y=481200
X659 1 2 1159 1143 2 151 1 sky130_fd_sc_hd__ebufn_2 $T=436540 481440 1 0 $X=436350 $Y=478480
X660 1 2 1160 1138 2 157 1 sky130_fd_sc_hd__ebufn_2 $T=438380 503200 0 0 $X=438190 $Y=502960
X661 1 2 1171 1142 2 167 1 sky130_fd_sc_hd__ebufn_2 $T=446660 470560 0 0 $X=446470 $Y=470320
X662 1 2 1206 1199 2 157 1 sky130_fd_sc_hd__ebufn_2 $T=458620 470560 0 0 $X=458430 $Y=470320
X663 1 2 1215 1199 2 170 1 sky130_fd_sc_hd__ebufn_2 $T=460920 481440 1 0 $X=460730 $Y=478480
X664 1 2 1227 1230 2 167 1 sky130_fd_sc_hd__ebufn_2 $T=464600 492320 1 0 $X=464410 $Y=489360
X665 1 2 1228 1216 2 167 1 sky130_fd_sc_hd__ebufn_2 $T=464600 497760 1 0 $X=464410 $Y=494800
X666 1 2 1209 1105 2 151 1 sky130_fd_sc_hd__ebufn_2 $T=469200 465120 1 0 $X=469010 $Y=462160
X667 1 2 1242 1231 2 156 1 sky130_fd_sc_hd__ebufn_2 $T=474720 508640 0 0 $X=474530 $Y=508400
X668 1 2 1254 228 2 157 1 sky130_fd_sc_hd__ebufn_2 $T=477020 465120 1 0 $X=476830 $Y=462160
X669 1 2 1259 228 2 156 1 sky130_fd_sc_hd__ebufn_2 $T=480700 459680 1 0 $X=480510 $Y=456720
X670 1 2 1279 1282 2 164 1 sky130_fd_sc_hd__ebufn_2 $T=493580 486880 0 0 $X=493390 $Y=486640
X671 1 2 1329 1293 2 156 1 sky130_fd_sc_hd__ebufn_2 $T=518420 486880 1 0 $X=518230 $Y=483920
X672 1 2 1327 1322 2 156 1 sky130_fd_sc_hd__ebufn_2 $T=519340 514080 1 0 $X=519150 $Y=511120
X673 1 2 1359 1351 2 262 1 sky130_fd_sc_hd__ebufn_2 $T=532220 443360 0 0 $X=532030 $Y=443120
X674 1 2 1363 1365 2 255 1 sky130_fd_sc_hd__ebufn_2 $T=533600 459680 1 0 $X=533410 $Y=456720
X675 1 2 1368 1371 2 266 1 sky130_fd_sc_hd__ebufn_2 $T=534520 481440 0 0 $X=534330 $Y=481200
X676 1 2 1382 1351 2 268 1 sky130_fd_sc_hd__ebufn_2 $T=548320 454240 1 0 $X=548130 $Y=451280
X677 1 2 1406 1409 2 266 1 sky130_fd_sc_hd__ebufn_2 $T=554300 459680 1 0 $X=554110 $Y=456720
X678 1 2 1407 1409 2 270 1 sky130_fd_sc_hd__ebufn_2 $T=554300 465120 1 0 $X=554110 $Y=462160
X679 1 2 1410 1412 2 264 1 sky130_fd_sc_hd__ebufn_2 $T=556140 470560 1 0 $X=555950 $Y=467600
X680 1 2 1437 1438 2 255 1 sky130_fd_sc_hd__ebufn_2 $T=570400 508640 1 0 $X=570210 $Y=505680
X681 1 2 1464 1438 2 268 1 sky130_fd_sc_hd__ebufn_2 $T=581440 503200 1 0 $X=581250 $Y=500240
X682 1 2 1468 1459 2 275 1 sky130_fd_sc_hd__ebufn_2 $T=583280 459680 1 0 $X=583090 $Y=456720
X683 1 2 1478 1476 2 275 1 sky130_fd_sc_hd__ebufn_2 $T=593400 492320 1 0 $X=593210 $Y=489360
X684 1 2 1489 1456 2 255 1 sky130_fd_sc_hd__ebufn_2 $T=595240 470560 0 0 $X=595050 $Y=470320
X685 1 2 1480 1476 2 270 1 sky130_fd_sc_hd__ebufn_2 $T=595240 486880 0 0 $X=595050 $Y=486640
X686 1 2 1479 1495 2 255 1 sky130_fd_sc_hd__ebufn_2 $T=595700 514080 1 0 $X=595510 $Y=511120
X687 1 2 1532 287 2 275 1 sky130_fd_sc_hd__ebufn_2 $T=615940 476000 1 0 $X=615750 $Y=473040
X688 1 2 1537 287 2 270 1 sky130_fd_sc_hd__ebufn_2 $T=617320 448800 1 0 $X=617130 $Y=445840
X689 1 2 1564 1556 2 266 1 sky130_fd_sc_hd__ebufn_2 $T=629280 492320 1 0 $X=629090 $Y=489360
X690 1 2 1565 287 2 262 1 sky130_fd_sc_hd__ebufn_2 $T=632500 448800 1 0 $X=632310 $Y=445840
X691 1 2 1574 1556 2 270 1 sky130_fd_sc_hd__ebufn_2 $T=632960 508640 0 0 $X=632770 $Y=508400
X692 1 2 1580 1556 2 275 1 sky130_fd_sc_hd__ebufn_2 $T=635720 503200 0 0 $X=635530 $Y=502960
X693 1 2 1628 301 2 268 1 sky130_fd_sc_hd__ebufn_2 $T=661020 454240 1 0 $X=660830 $Y=451280
X694 1 2 1645 1631 2 268 1 sky130_fd_sc_hd__ebufn_2 $T=666540 503200 1 0 $X=666350 $Y=500240
X695 1 2 1656 301 2 264 1 sky130_fd_sc_hd__ebufn_2 $T=679420 454240 0 0 $X=679230 $Y=454000
X696 1 2 1685 1658 2 270 1 sky130_fd_sc_hd__ebufn_2 $T=697820 497760 0 0 $X=697630 $Y=497520
X697 1 2 1707 1692 2 255 1 sky130_fd_sc_hd__ebufn_2 $T=702880 492320 0 0 $X=702690 $Y=492080
X698 1 2 1747 1738 2 268 1 sky130_fd_sc_hd__ebufn_2 $T=721740 497760 1 0 $X=721550 $Y=494800
X699 1 2 1757 317 2 275 1 sky130_fd_sc_hd__ebufn_2 $T=735540 443360 0 0 $X=735350 $Y=443120
X814 1 2 ICV_5 $T=47840 503200 1 0 $X=47650 $Y=500240
X815 1 2 ICV_5 $T=145820 508640 0 0 $X=145630 $Y=508400
X816 1 2 ICV_5 $T=230000 486880 0 0 $X=229810 $Y=486640
X817 1 2 ICV_5 $T=300380 492320 1 0 $X=300190 $Y=489360
X818 1 2 ICV_5 $T=304980 514080 1 0 $X=304790 $Y=511120
X819 1 2 ICV_5 $T=333500 514080 1 0 $X=333310 $Y=511120
X820 1 2 ICV_5 $T=637100 508640 1 0 $X=636910 $Y=505680
X821 1 2 ICV_5 $T=650900 476000 0 0 $X=650710 $Y=475760
X822 1 2 ICV_5 $T=732780 514080 1 0 $X=732590 $Y=511120
X823 1 2 ICV_5 $T=735080 465120 0 0 $X=734890 $Y=464880
X824 1 2 ICV_5 $T=735080 470560 0 0 $X=734890 $Y=470320
X825 1 2 ICV_5 $T=735080 476000 0 0 $X=734890 $Y=475760
X826 1 2 ICV_5 $T=735080 481440 0 0 $X=734890 $Y=481200
X827 1 2 ICV_5 $T=735080 492320 0 0 $X=734890 $Y=492080
X828 1 2 ICV_5 $T=735080 497760 0 0 $X=734890 $Y=497520
X829 1 2 ICV_5 $T=735080 503200 0 0 $X=734890 $Y=502960
X830 1 2 344 340 20 ICV_6 $T=19780 503200 1 0 $X=19590 $Y=500240
X831 1 2 400 382 28 ICV_6 $T=47840 497760 1 0 $X=47650 $Y=494800
X832 1 2 411 43 20 ICV_6 $T=61640 454240 0 0 $X=61450 $Y=454000
X833 1 2 427 364 25 ICV_6 $T=61640 459680 0 0 $X=61450 $Y=459440
X834 1 2 410 420 25 ICV_6 $T=61640 476000 0 0 $X=61450 $Y=475760
X835 1 2 422 428 22 ICV_6 $T=61640 503200 0 0 $X=61450 $Y=502960
X836 1 2 449 448 27 ICV_6 $T=75900 448800 1 0 $X=75710 $Y=445840
X837 1 2 408 364 22 ICV_6 $T=75900 465120 1 0 $X=75710 $Y=462160
X838 1 2 406 364 32 ICV_6 $T=75900 470560 1 0 $X=75710 $Y=467600
X839 1 2 482 485 30 ICV_6 $T=89700 448800 0 0 $X=89510 $Y=448560
X840 1 2 483 485 21 ICV_6 $T=89700 459680 0 0 $X=89510 $Y=459440
X841 1 2 472 470 30 ICV_6 $T=89700 476000 0 0 $X=89510 $Y=475760
X842 1 2 481 459 28 ICV_6 $T=89700 497760 0 0 $X=89510 $Y=497520
X843 1 2 517 529 25 ICV_6 $T=117760 470560 0 0 $X=117570 $Y=470320
X844 1 2 565 561 21 ICV_6 $T=132020 470560 1 0 $X=131830 $Y=467600
X845 1 2 646 616 89 ICV_6 $T=173880 465120 0 0 $X=173690 $Y=464880
X846 1 2 683 624 32 ICV_6 $T=188140 503200 1 0 $X=187950 $Y=500240
X847 1 2 708 704 20 ICV_6 $T=201940 459680 0 0 $X=201750 $Y=459440
X848 1 2 702 705 94 ICV_6 $T=201940 476000 0 0 $X=201750 $Y=475760
X849 1 2 697 705 92 ICV_6 $T=201940 481440 0 0 $X=201750 $Y=481200
X850 1 2 706 689 30 ICV_6 $T=201940 492320 0 0 $X=201750 $Y=492080
X851 1 2 709 689 21 ICV_6 $T=201940 497760 0 0 $X=201750 $Y=497520
X852 1 2 760 752 93 ICV_6 $T=230000 443360 0 0 $X=229810 $Y=443120
X853 1 2 790 769 101 ICV_6 $T=244260 481440 1 0 $X=244070 $Y=478480
X854 1 2 789 736 22 ICV_6 $T=244260 503200 1 0 $X=244070 $Y=500240
X855 1 2 816 812 89 ICV_6 $T=258060 481440 0 0 $X=257870 $Y=481200
X856 1 2 870 143 103 ICV_6 $T=300380 448800 1 0 $X=300190 $Y=445840
X857 1 2 892 143 92 ICV_6 $T=314180 443360 0 0 $X=313990 $Y=443120
X858 1 2 894 876 102 ICV_6 $T=314180 470560 0 0 $X=313990 $Y=470320
X859 1 2 893 876 96 ICV_6 $T=314180 476000 0 0 $X=313990 $Y=475760
X860 1 2 920 925 155 ICV_6 $T=328440 503200 1 0 $X=328250 $Y=500240
X861 1 2 979 958 155 ICV_6 $T=356500 470560 1 0 $X=356310 $Y=467600
X862 1 2 1003 1014 170 ICV_6 $T=370300 465120 0 0 $X=370110 $Y=464880
X863 1 2 1039 1014 155 ICV_6 $T=384560 476000 1 0 $X=384370 $Y=473040
X864 1 2 1072 1046 151 ICV_6 $T=398360 454240 0 0 $X=398170 $Y=454000
X865 1 2 1052 1051 151 ICV_6 $T=398360 465120 0 0 $X=398170 $Y=464880
X866 1 2 1066 1016 152 ICV_6 $T=398360 486880 0 0 $X=398170 $Y=486640
X867 1 2 1091 1065 170 ICV_6 $T=404800 514080 1 0 $X=404610 $Y=511120
X868 1 2 1101 204 157 ICV_6 $T=412620 448800 1 0 $X=412430 $Y=445840
X869 1 2 1140 1142 155 ICV_6 $T=426420 465120 0 0 $X=426230 $Y=464880
X870 1 2 1141 1143 152 ICV_6 $T=426420 492320 0 0 $X=426230 $Y=492080
X871 1 2 1123 1129 152 ICV_6 $T=426420 497760 0 0 $X=426230 $Y=497520
X872 1 2 1173 1176 167 ICV_6 $T=440680 459680 1 0 $X=440490 $Y=456720
X873 1 2 1157 1142 170 ICV_6 $T=440680 465120 1 0 $X=440490 $Y=462160
X874 1 2 1168 1142 151 ICV_6 $T=440680 481440 1 0 $X=440490 $Y=478480
X875 1 2 1174 1143 157 ICV_6 $T=440680 492320 1 0 $X=440490 $Y=489360
X876 1 2 1164 1138 152 ICV_6 $T=440680 503200 1 0 $X=440490 $Y=500240
X877 1 2 1158 1138 156 ICV_6 $T=440680 508640 1 0 $X=440490 $Y=505680
X878 1 2 1198 1176 157 ICV_6 $T=454480 459680 0 0 $X=454290 $Y=459440
X879 1 2 1192 1105 157 ICV_6 $T=454480 486880 0 0 $X=454290 $Y=486640
X880 1 2 1201 1205 167 ICV_6 $T=461840 514080 1 0 $X=461650 $Y=511120
X881 1 2 1222 1105 155 ICV_6 $T=468740 470560 1 0 $X=468550 $Y=467600
X882 1 2 1285 1282 152 ICV_6 $T=496800 459680 1 0 $X=496610 $Y=456720
X883 1 2 1352 1354 255 ICV_6 $T=524860 492320 1 0 $X=524670 $Y=489360
X884 1 2 1367 1365 268 ICV_6 $T=538660 465120 0 0 $X=538470 $Y=464880
X885 1 2 1372 1354 264 ICV_6 $T=538660 481440 0 0 $X=538470 $Y=481200
X886 1 2 1374 1354 266 ICV_6 $T=538660 492320 0 0 $X=538470 $Y=492080
X887 1 2 1396 1378 268 ICV_6 $T=547400 514080 1 0 $X=547210 $Y=511120
X888 1 2 1394 1371 275 ICV_6 $T=552920 486880 1 0 $X=552730 $Y=483920
X889 1 2 1427 1409 255 ICV_6 $T=566720 454240 0 0 $X=566530 $Y=454000
X890 1 2 1432 1412 268 ICV_6 $T=566720 470560 0 0 $X=566530 $Y=470320
X891 1 2 1452 1459 269 ICV_6 $T=580980 465120 1 0 $X=580790 $Y=462160
X892 1 2 1454 1459 264 ICV_6 $T=580980 470560 1 0 $X=580790 $Y=467600
X893 1 2 1462 1456 270 ICV_6 $T=580980 481440 1 0 $X=580790 $Y=478480
X894 1 2 1460 1438 270 ICV_6 $T=580980 508640 1 0 $X=580790 $Y=505680
X895 1 2 1483 1459 262 ICV_6 $T=594780 459680 0 0 $X=594590 $Y=459440
X896 1 2 1485 1495 270 ICV_6 $T=594780 508640 0 0 $X=594590 $Y=508400
X897 1 2 1509 1516 268 ICV_6 $T=609040 470560 1 0 $X=608850 $Y=467600
X898 1 2 1515 1516 264 ICV_6 $T=609040 476000 1 0 $X=608850 $Y=473040
X899 1 2 1535 1524 268 ICV_6 $T=618700 514080 1 0 $X=618510 $Y=511120
X900 1 2 1577 1556 269 ICV_6 $T=637100 497760 1 0 $X=636910 $Y=494800
X901 1 2 1611 1563 270 ICV_6 $T=650900 465120 0 0 $X=650710 $Y=464880
X902 1 2 1607 1613 262 ICV_6 $T=650900 497760 0 0 $X=650710 $Y=497520
X903 1 2 1602 1613 270 ICV_6 $T=650900 503200 0 0 $X=650710 $Y=502960
X904 1 2 1640 301 270 ICV_6 $T=665160 454240 1 0 $X=664970 $Y=451280
X905 1 2 1633 1619 268 ICV_6 $T=665160 465120 1 0 $X=664970 $Y=462160
X906 1 2 1666 301 262 ICV_6 $T=678960 443360 0 0 $X=678770 $Y=443120
X907 1 2 1660 301 255 ICV_6 $T=678960 448800 0 0 $X=678770 $Y=448560
X908 1 2 1711 1705 266 ICV_6 $T=707020 492320 0 0 $X=706830 $Y=492080
X909 1 2 1764 1733 269 ICV_6 $T=735080 459680 0 0 $X=734890 $Y=459440
X1041 1 2 ICV_9 $T=6900 492320 0 0 $X=6710 $Y=492080
X1042 1 2 ICV_9 $T=79120 503200 0 0 $X=78930 $Y=502960
X1043 1 2 ICV_9 $T=180320 508640 0 0 $X=180130 $Y=508400
X1044 1 2 ICV_9 $T=206540 508640 1 0 $X=206350 $Y=505680
X1045 1 2 ICV_9 $T=216660 508640 1 0 $X=216470 $Y=505680
X1046 1 2 ICV_9 $T=303600 486880 0 0 $X=303410 $Y=486640
X1047 1 2 ICV_9 $T=552000 514080 1 0 $X=551810 $Y=511120
X1048 1 2 ICV_9 $T=575000 508640 0 0 $X=574810 $Y=508400
X1049 1 2 ICV_9 $T=599380 508640 0 0 $X=599190 $Y=508400
X1050 1 2 ICV_9 $T=604900 514080 1 0 $X=604710 $Y=511120
X1051 1 2 ICV_9 $T=623300 514080 1 0 $X=623110 $Y=511120
X1052 1 2 ICV_9 $T=668840 508640 0 0 $X=668650 $Y=508400
X1053 1 2 ICV_9 $T=690460 508640 0 0 $X=690270 $Y=508400
X1054 1 2 ICV_9 $T=732780 503200 1 0 $X=732590 $Y=500240
X1055 1 2 ICV_9 $T=732780 508640 1 0 $X=732590 $Y=505680
X1056 1 2 ICV_9 $T=733240 454240 1 0 $X=733050 $Y=451280
X1057 1 2 ICV_9 $T=733240 470560 1 0 $X=733050 $Y=467600
X1058 1 2 ICV_9 $T=733240 481440 1 0 $X=733050 $Y=478480
X1059 1 2 ICV_9 $T=733700 476000 1 0 $X=733510 $Y=473040
X1060 1 2 ICV_10 $T=30820 459680 0 0 $X=30630 $Y=459440
X1061 1 2 ICV_10 $T=58880 443360 0 0 $X=58690 $Y=443120
X1062 1 2 ICV_10 $T=58880 486880 0 0 $X=58690 $Y=486640
X1063 1 2 ICV_10 $T=58880 508640 0 0 $X=58690 $Y=508400
X1064 1 2 ICV_10 $T=115000 448800 0 0 $X=114810 $Y=448560
X1065 1 2 ICV_10 $T=157320 486880 1 0 $X=157130 $Y=483920
X1066 1 2 ICV_10 $T=199180 508640 0 0 $X=198990 $Y=508400
X1067 1 2 ICV_10 $T=227240 448800 0 0 $X=227050 $Y=448560
X1068 1 2 ICV_10 $T=227240 497760 0 0 $X=227050 $Y=497520
X1069 1 2 ICV_10 $T=297620 481440 1 0 $X=297430 $Y=478480
X1070 1 2 ICV_10 $T=345000 514080 1 0 $X=344810 $Y=511120
X1071 1 2 ICV_10 $T=367540 486880 0 0 $X=367350 $Y=486640
X1072 1 2 ICV_10 $T=409860 476000 1 0 $X=409670 $Y=473040
X1073 1 2 ICV_10 $T=409860 497760 1 0 $X=409670 $Y=494800
X1074 1 2 ICV_10 $T=437920 476000 1 0 $X=437730 $Y=473040
X1075 1 2 ICV_10 $T=507840 503200 0 0 $X=507650 $Y=502960
X1076 1 2 ICV_10 $T=578220 454240 1 0 $X=578030 $Y=451280
X1077 1 2 ICV_10 $T=587420 514080 1 0 $X=587230 $Y=511120
X1078 1 2 ICV_10 $T=704260 508640 0 0 $X=704070 $Y=508400
X1079 1 2 ICV_10 $T=732320 508640 0 0 $X=732130 $Y=508400
X1080 1 2 ICV_11 $T=6900 503200 1 0 $X=6710 $Y=500240
X1081 1 2 ICV_11 $T=6900 503200 0 0 $X=6710 $Y=502960
X1082 1 2 ICV_11 $T=6900 508640 1 0 $X=6710 $Y=505680
X1083 1 2 ICV_11 $T=6900 514080 1 0 $X=6710 $Y=511120
X1084 1 2 ICV_11 $T=17940 503200 0 0 $X=17750 $Y=502960
X1085 1 2 ICV_11 $T=19320 508640 0 0 $X=19130 $Y=508400
X1086 1 2 ICV_11 $T=20240 508640 1 0 $X=20050 $Y=505680
X1087 1 2 ICV_11 $T=20240 514080 1 0 $X=20050 $Y=511120
X1088 1 2 ICV_11 $T=24380 503200 1 0 $X=24190 $Y=500240
X1089 1 2 ICV_11 $T=42320 503200 0 0 $X=42130 $Y=502960
X1090 1 2 ICV_11 $T=48300 508640 1 0 $X=48110 $Y=505680
X1091 1 2 ICV_11 $T=67160 508640 0 0 $X=66970 $Y=508400
X1092 1 2 ICV_11 $T=76360 508640 1 0 $X=76170 $Y=505680
X1093 1 2 ICV_11 $T=87400 508640 1 0 $X=87210 $Y=505680
X1094 1 2 ICV_11 $T=104420 508640 1 0 $X=104230 $Y=505680
X1095 1 2 ICV_11 $T=132480 508640 1 0 $X=132290 $Y=505680
X1096 1 2 ICV_11 $T=175260 508640 1 0 $X=175070 $Y=505680
X1097 1 2 ICV_11 $T=230460 508640 0 0 $X=230270 $Y=508400
X1098 1 2 ICV_11 $T=245640 503200 0 0 $X=245450 $Y=502960
X1099 1 2 ICV_11 $T=248860 497760 1 0 $X=248670 $Y=494800
X1100 1 2 ICV_11 $T=248860 503200 1 0 $X=248670 $Y=500240
X1101 1 2 ICV_11 $T=250240 508640 1 0 $X=250050 $Y=505680
X1102 1 2 ICV_11 $T=258520 497760 0 0 $X=258330 $Y=497520
X1103 1 2 ICV_11 $T=258520 503200 0 0 $X=258330 $Y=502960
X1104 1 2 ICV_11 $T=258520 508640 0 0 $X=258330 $Y=508400
X1105 1 2 ICV_11 $T=259900 497760 1 0 $X=259710 $Y=494800
X1106 1 2 ICV_11 $T=259900 503200 1 0 $X=259710 $Y=500240
X1107 1 2 ICV_11 $T=261280 508640 1 0 $X=261090 $Y=505680
X1108 1 2 ICV_11 $T=272780 492320 1 0 $X=272590 $Y=489360
X1109 1 2 ICV_11 $T=272780 497760 1 0 $X=272590 $Y=494800
X1110 1 2 ICV_11 $T=272780 508640 1 0 $X=272590 $Y=505680
X1111 1 2 ICV_11 $T=275080 508640 0 0 $X=274890 $Y=508400
X1112 1 2 ICV_11 $T=286580 503200 0 0 $X=286390 $Y=502960
X1113 1 2 ICV_11 $T=286580 508640 0 0 $X=286390 $Y=508400
X1114 1 2 ICV_11 $T=300840 503200 1 0 $X=300650 $Y=500240
X1115 1 2 ICV_11 $T=300840 508640 1 0 $X=300650 $Y=505680
X1116 1 2 ICV_11 $T=319700 514080 1 0 $X=319510 $Y=511120
X1117 1 2 ICV_11 $T=533600 514080 1 0 $X=533410 $Y=511120
X1118 1 2 ICV_11 $T=553840 508640 0 0 $X=553650 $Y=508400
X1119 1 2 ICV_11 $T=562120 514080 1 0 $X=561930 $Y=511120
X1120 1 2 ICV_11 $T=633420 514080 1 0 $X=633230 $Y=511120
X1121 1 2 ICV_11 $T=651360 508640 0 0 $X=651170 $Y=508400
X1122 1 2 ICV_11 $T=679420 503200 0 0 $X=679230 $Y=502960
X1123 1 2 ICV_11 $T=709320 503200 1 0 $X=709130 $Y=500240
X1124 1 2 ICV_11 $T=718980 497760 0 0 $X=718790 $Y=497520
X1125 1 2 ICV_11 $T=718980 503200 0 0 $X=718790 $Y=502960
X1126 1 2 ICV_11 $T=721740 503200 1 0 $X=721550 $Y=500240
X1127 1 2 ICV_11 $T=721740 508640 1 0 $X=721550 $Y=505680
X1128 1 2 ICV_12 $T=31280 508640 1 0 $X=31090 $Y=505680
X1129 1 2 ICV_12 $T=42320 508640 0 0 $X=42130 $Y=508400
X1130 1 2 ICV_12 $T=59340 508640 1 0 $X=59150 $Y=505680
X1131 1 2 ICV_12 $T=115460 508640 1 0 $X=115270 $Y=505680
X1132 1 2 ICV_12 $T=118220 508640 0 0 $X=118030 $Y=508400
X1133 1 2 ICV_12 $T=239660 497760 0 0 $X=239470 $Y=497520
X1134 1 2 ICV_12 $T=241500 508640 0 0 $X=241310 $Y=508400
X1135 1 2 ICV_12 $T=252080 492320 1 0 $X=251890 $Y=489360
X1136 1 2 ICV_12 $T=267260 486880 0 0 $X=267070 $Y=486640
X1137 1 2 ICV_12 $T=269560 492320 0 0 $X=269370 $Y=492080
X1138 1 2 ICV_12 $T=269560 497760 0 0 $X=269370 $Y=497520
X1139 1 2 ICV_12 $T=269560 503200 0 0 $X=269370 $Y=502960
X1140 1 2 ICV_12 $T=272780 503200 1 0 $X=272590 $Y=500240
X1141 1 2 ICV_12 $T=283820 492320 1 0 $X=283630 $Y=489360
X1142 1 2 ICV_12 $T=283820 497760 1 0 $X=283630 $Y=494800
X1143 1 2 ICV_12 $T=283820 508640 1 0 $X=283630 $Y=505680
X1144 1 2 ICV_12 $T=286580 492320 0 0 $X=286390 $Y=492080
X1145 1 2 ICV_12 $T=286580 497760 0 0 $X=286390 $Y=497520
X1146 1 2 ICV_12 $T=297620 503200 0 0 $X=297430 $Y=502960
X1147 1 2 ICV_12 $T=297620 508640 0 0 $X=297430 $Y=508400
X1148 1 2 ICV_12 $T=675280 508640 1 0 $X=675090 $Y=505680
X1149 1 2 ICV_12 $T=715760 508640 0 0 $X=715570 $Y=508400
X1150 1 2 ICV_12 $T=717140 481440 0 0 $X=716950 $Y=481200
X1151 1 2 ICV_12 $T=725880 497760 1 0 $X=725690 $Y=494800
X1152 1 2 328 9 2 341 1 sky130_fd_sc_hd__dfxtp_1 $T=10580 497760 1 0 $X=10390 $Y=494800
X1153 1 2 355 13 2 373 1 sky130_fd_sc_hd__dfxtp_1 $T=28980 486880 1 0 $X=28790 $Y=483920
X1154 1 2 370 24 2 399 1 sky130_fd_sc_hd__dfxtp_1 $T=41400 465120 0 0 $X=41210 $Y=464880
X1155 1 2 371 26 2 401 1 sky130_fd_sc_hd__dfxtp_1 $T=43240 486880 0 0 $X=43050 $Y=486640
X1156 1 2 407 8 2 425 1 sky130_fd_sc_hd__dfxtp_1 $T=53820 497760 0 0 $X=53630 $Y=497520
X1157 1 2 433 15 2 449 1 sky130_fd_sc_hd__dfxtp_1 $T=65780 448800 0 0 $X=65590 $Y=448560
X1158 1 2 445 24 2 456 1 sky130_fd_sc_hd__dfxtp_1 $T=71760 503200 0 0 $X=71570 $Y=502960
X1159 1 2 457 9 2 473 1 sky130_fd_sc_hd__dfxtp_1 $T=80040 476000 1 0 $X=79850 $Y=473040
X1160 1 2 445 19 2 481 1 sky130_fd_sc_hd__dfxtp_1 $T=83260 497760 1 0 $X=83070 $Y=494800
X1161 1 2 487 15 2 520 1 sky130_fd_sc_hd__dfxtp_1 $T=104420 503200 0 0 $X=104230 $Y=502960
X1162 1 2 509 24 2 527 1 sky130_fd_sc_hd__dfxtp_1 $T=105340 476000 0 0 $X=105150 $Y=475760
X1163 1 2 509 19 2 528 1 sky130_fd_sc_hd__dfxtp_1 $T=105800 481440 1 0 $X=105610 $Y=478480
X1164 1 2 511 13 2 534 1 sky130_fd_sc_hd__dfxtp_1 $T=108100 459680 1 0 $X=107910 $Y=456720
X1165 1 2 509 15 2 538 1 sky130_fd_sc_hd__dfxtp_1 $T=110400 470560 0 0 $X=110210 $Y=470320
X1166 1 2 509 7 2 542 1 sky130_fd_sc_hd__dfxtp_1 $T=115920 481440 1 0 $X=115730 $Y=478480
X1167 1 2 69 8 2 556 1 sky130_fd_sc_hd__dfxtp_1 $T=124660 448800 1 0 $X=124470 $Y=445840
X1168 1 2 547 24 2 590 1 sky130_fd_sc_hd__dfxtp_1 $T=137080 481440 1 0 $X=136890 $Y=478480
X1169 1 2 593 82 2 607 1 sky130_fd_sc_hd__dfxtp_1 $T=147660 470560 1 0 $X=147470 $Y=467600
X1170 1 2 594 86 2 622 1 sky130_fd_sc_hd__dfxtp_1 $T=149960 470560 0 0 $X=149770 $Y=470320
X1171 1 2 619 26 2 625 1 sky130_fd_sc_hd__dfxtp_1 $T=155940 492320 0 0 $X=155750 $Y=492080
X1172 1 2 635 85 2 652 1 sky130_fd_sc_hd__dfxtp_1 $T=166520 476000 0 0 $X=166330 $Y=475760
X1173 1 2 649 99 2 662 1 sky130_fd_sc_hd__dfxtp_1 $T=172960 465120 1 0 $X=172770 $Y=462160
X1174 1 2 649 86 2 673 1 sky130_fd_sc_hd__dfxtp_1 $T=178020 459680 0 0 $X=177830 $Y=459440
X1175 1 2 649 85 2 680 1 sky130_fd_sc_hd__dfxtp_1 $T=181700 448800 0 0 $X=181510 $Y=448560
X1176 1 2 665 7 2 709 1 sky130_fd_sc_hd__dfxtp_1 $T=193200 497760 0 0 $X=193010 $Y=497520
X1177 1 2 690 24 2 701 1 sky130_fd_sc_hd__dfxtp_1 $T=193660 454240 1 0 $X=193470 $Y=451280
X1178 1 2 682 98 2 703 1 sky130_fd_sc_hd__dfxtp_1 $T=195960 486880 1 0 $X=195770 $Y=483920
X1179 1 2 718 98 2 730 1 sky130_fd_sc_hd__dfxtp_1 $T=207000 470560 0 0 $X=206810 $Y=470320
X1180 1 2 718 83 2 741 1 sky130_fd_sc_hd__dfxtp_1 $T=207460 470560 1 0 $X=207270 $Y=467600
X1181 1 2 719 7 2 759 1 sky130_fd_sc_hd__dfxtp_1 $T=220340 481440 1 0 $X=220150 $Y=478480
X1182 1 2 762 97 2 787 1 sky130_fd_sc_hd__dfxtp_1 $T=235060 486880 1 0 $X=234870 $Y=483920
X1183 1 2 762 95 2 792 1 sky130_fd_sc_hd__dfxtp_1 $T=237820 470560 0 0 $X=237630 $Y=470320
X1184 1 2 798 98 2 816 1 sky130_fd_sc_hd__dfxtp_1 $T=250700 481440 0 0 $X=250510 $Y=481200
X1185 1 2 786 85 2 819 1 sky130_fd_sc_hd__dfxtp_1 $T=256680 454240 1 0 $X=256490 $Y=451280
X1186 1 2 855 99 2 873 1 sky130_fd_sc_hd__dfxtp_1 $T=296240 486880 0 0 $X=296050 $Y=486640
X1187 1 2 904 149 2 920 1 sky130_fd_sc_hd__dfxtp_1 $T=321080 503200 1 0 $X=320890 $Y=500240
X1188 1 2 895 144 2 928 1 sky130_fd_sc_hd__dfxtp_1 $T=325220 459680 0 0 $X=325030 $Y=459440
X1189 1 2 904 159 2 953 1 sky130_fd_sc_hd__dfxtp_1 $T=334880 508640 0 0 $X=334690 $Y=508400
X1190 1 2 904 161 2 951 1 sky130_fd_sc_hd__dfxtp_1 $T=336260 508640 1 0 $X=336070 $Y=505680
X1191 1 2 898 165 2 924 1 sky130_fd_sc_hd__dfxtp_1 $T=337640 481440 1 0 $X=337450 $Y=478480
X1192 1 2 968 146 2 984 1 sky130_fd_sc_hd__dfxtp_1 $T=353740 497760 0 0 $X=353550 $Y=497520
X1193 1 2 990 159 2 1011 1 sky130_fd_sc_hd__dfxtp_1 $T=362940 481440 0 0 $X=362750 $Y=481200
X1194 1 2 1019 161 2 1036 1 sky130_fd_sc_hd__dfxtp_1 $T=374440 508640 0 0 $X=374250 $Y=508400
X1195 1 2 989 165 2 1035 1 sky130_fd_sc_hd__dfxtp_1 $T=376740 470560 1 0 $X=376550 $Y=467600
X1196 1 2 1025 144 2 1042 1 sky130_fd_sc_hd__dfxtp_1 $T=377200 448800 1 0 $X=377010 $Y=445840
X1197 1 2 990 149 2 1048 1 sky130_fd_sc_hd__dfxtp_1 $T=379960 481440 0 0 $X=379770 $Y=481200
X1198 1 2 1019 165 2 1020 1 sky130_fd_sc_hd__dfxtp_1 $T=381340 503200 0 0 $X=381150 $Y=502960
X1199 1 2 1025 154 2 1068 1 sky130_fd_sc_hd__dfxtp_1 $T=391000 448800 0 0 $X=390810 $Y=448560
X1200 1 2 1034 144 2 1074 1 sky130_fd_sc_hd__dfxtp_1 $T=392380 470560 1 0 $X=392190 $Y=467600
X1201 1 2 1086 161 2 1127 1 sky130_fd_sc_hd__dfxtp_1 $T=413540 508640 0 0 $X=413350 $Y=508400
X1202 1 2 1118 159 2 1135 1 sky130_fd_sc_hd__dfxtp_1 $T=419060 481440 0 0 $X=418870 $Y=481200
X1203 1 2 1082 144 2 1139 1 sky130_fd_sc_hd__dfxtp_1 $T=420440 465120 1 0 $X=420250 $Y=462160
X1204 1 2 1130 150 2 1148 1 sky130_fd_sc_hd__dfxtp_1 $T=421820 476000 1 0 $X=421630 $Y=473040
X1205 1 2 1152 144 2 1164 1 sky130_fd_sc_hd__dfxtp_1 $T=431020 492320 0 0 $X=430830 $Y=492080
X1206 1 2 1152 146 2 1165 1 sky130_fd_sc_hd__dfxtp_1 $T=431020 497760 0 0 $X=430830 $Y=497520
X1207 1 2 1152 161 2 1167 1 sky130_fd_sc_hd__dfxtp_1 $T=431480 508640 0 0 $X=431290 $Y=508400
X1208 1 2 1180 161 2 1104 1 sky130_fd_sc_hd__dfxtp_1 $T=444820 492320 0 0 $X=444630 $Y=492080
X1209 1 2 1180 165 2 1183 1 sky130_fd_sc_hd__dfxtp_1 $T=446200 481440 0 0 $X=446010 $Y=481200
X1210 1 2 1153 146 2 1197 1 sky130_fd_sc_hd__dfxtp_1 $T=447120 454240 0 0 $X=446930 $Y=454000
X1211 1 2 1184 149 2 1200 1 sky130_fd_sc_hd__dfxtp_1 $T=447120 497760 0 0 $X=446930 $Y=497520
X1212 1 2 1184 150 2 1203 1 sky130_fd_sc_hd__dfxtp_1 $T=448960 508640 1 0 $X=448770 $Y=505680
X1213 1 2 1214 146 2 229 1 sky130_fd_sc_hd__dfxtp_1 $T=461380 459680 1 0 $X=461190 $Y=456720
X1214 1 2 1214 161 2 1235 1 sky130_fd_sc_hd__dfxtp_1 $T=461380 470560 1 0 $X=461190 $Y=467600
X1215 1 2 1213 149 2 1237 1 sky130_fd_sc_hd__dfxtp_1 $T=463220 448800 0 0 $X=463030 $Y=448560
X1216 1 2 1225 159 2 1243 1 sky130_fd_sc_hd__dfxtp_1 $T=466440 514080 1 0 $X=466250 $Y=511120
X1217 1 2 1261 165 2 1292 1 sky130_fd_sc_hd__dfxtp_1 $T=490820 503200 0 0 $X=490630 $Y=502960
X1218 1 2 1297 146 2 1317 1 sky130_fd_sc_hd__dfxtp_1 $T=500940 503200 1 0 $X=500750 $Y=500240
X1219 1 2 245 146 2 1318 1 sky130_fd_sc_hd__dfxtp_1 $T=501400 443360 0 0 $X=501210 $Y=443120
X1220 1 2 1358 257 2 1372 1 sky130_fd_sc_hd__dfxtp_1 $T=529000 497760 1 0 $X=528810 $Y=494800
X1221 1 2 1375 261 2 1396 1 sky130_fd_sc_hd__dfxtp_1 $T=544180 508640 1 0 $X=543990 $Y=505680
X1222 1 2 1386 261 2 1401 1 sky130_fd_sc_hd__dfxtp_1 $T=545560 465120 1 0 $X=545370 $Y=462160
X1223 1 2 1411 263 2 1426 1 sky130_fd_sc_hd__dfxtp_1 $T=557520 476000 0 0 $X=557330 $Y=475760
X1224 1 2 1386 256 2 1431 1 sky130_fd_sc_hd__dfxtp_1 $T=558900 459680 0 0 $X=558710 $Y=459440
X1225 1 2 1443 265 2 1453 1 sky130_fd_sc_hd__dfxtp_1 $T=572240 465120 0 0 $X=572050 $Y=464880
X1226 1 2 1446 263 2 1457 1 sky130_fd_sc_hd__dfxtp_1 $T=573620 476000 1 0 $X=573430 $Y=473040
X1227 1 2 277 258 2 1465 1 sky130_fd_sc_hd__dfxtp_1 $T=575920 454240 0 0 $X=575730 $Y=454000
X1228 1 2 1463 267 2 1478 1 sky130_fd_sc_hd__dfxtp_1 $T=583280 492320 0 0 $X=583090 $Y=492080
X1229 1 2 1446 261 2 1484 1 sky130_fd_sc_hd__dfxtp_1 $T=586500 481440 0 0 $X=586310 $Y=481200
X1230 1 2 1474 257 2 285 1 sky130_fd_sc_hd__dfxtp_1 $T=588800 448800 1 0 $X=588610 $Y=445840
X1231 1 2 1527 258 2 1545 1 sky130_fd_sc_hd__dfxtp_1 $T=613640 465120 0 0 $X=613450 $Y=464880
X1232 1 2 1527 261 2 1546 1 sky130_fd_sc_hd__dfxtp_1 $T=613640 470560 0 0 $X=613450 $Y=470320
X1233 1 2 1550 263 2 1577 1 sky130_fd_sc_hd__dfxtp_1 $T=626980 497760 1 0 $X=626790 $Y=494800
X1234 1 2 1578 258 2 1595 1 sky130_fd_sc_hd__dfxtp_1 $T=638020 470560 0 0 $X=637830 $Y=470320
X1235 1 2 1578 263 2 1599 1 sky130_fd_sc_hd__dfxtp_1 $T=643080 481440 0 0 $X=642890 $Y=481200
X1236 1 2 1576 256 2 1605 1 sky130_fd_sc_hd__dfxtp_1 $T=643540 465120 0 0 $X=643350 $Y=464880
X1237 1 2 1588 259 2 1612 1 sky130_fd_sc_hd__dfxtp_1 $T=644920 492320 1 0 $X=644730 $Y=489360
X1238 1 2 1618 261 2 1633 1 sky130_fd_sc_hd__dfxtp_1 $T=656420 470560 1 0 $X=656230 $Y=467600
X1239 1 2 300 257 2 1656 1 sky130_fd_sc_hd__dfxtp_1 $T=669760 454240 1 0 $X=669570 $Y=451280
X1240 1 2 300 258 2 1660 1 sky130_fd_sc_hd__dfxtp_1 $T=671140 454240 0 0 $X=670950 $Y=454000
X1241 1 2 1652 261 2 1671 1 sky130_fd_sc_hd__dfxtp_1 $T=673900 481440 1 0 $X=673710 $Y=478480
X1242 1 2 1668 265 2 1697 1 sky130_fd_sc_hd__dfxtp_1 $T=691380 465120 0 0 $X=691190 $Y=464880
X1243 1 2 1681 257 2 1709 1 sky130_fd_sc_hd__dfxtp_1 $T=696440 470560 0 0 $X=696250 $Y=470320
X1244 1 2 329 18 21 3 7 329 ICV_13 $T=6900 448800 1 0 $X=6710 $Y=445840
X1245 1 2 330 18 20 3 8 330 ICV_13 $T=6900 454240 1 0 $X=6710 $Y=451280
X1246 1 2 331 334 21 323 7 331 ICV_13 $T=6900 476000 0 0 $X=6710 $Y=475760
X1247 1 2 351 334 32 328 15 346 ICV_13 $T=17480 486880 0 0 $X=17290 $Y=486640
X1248 1 2 357 339 27 325 15 357 ICV_13 $T=20240 459680 1 0 $X=20050 $Y=456720
X1249 1 2 359 340 30 328 26 359 ICV_13 $T=20240 492320 1 0 $X=20050 $Y=489360
X1250 1 2 360 340 28 328 19 360 ICV_13 $T=20240 497760 1 0 $X=20050 $Y=494800
X1251 1 2 363 340 32 328 24 363 ICV_13 $T=21620 497760 0 0 $X=21430 $Y=497520
X1252 1 2 377 385 30 370 26 377 ICV_13 $T=32200 454240 1 0 $X=32010 $Y=451280
X1253 1 2 383 385 25 370 13 383 ICV_13 $T=32660 465120 1 0 $X=32470 $Y=462160
X1254 1 2 386 35 28 33 19 386 ICV_13 $T=34040 443360 0 0 $X=33850 $Y=443120
X1255 1 2 388 385 28 370 19 388 ICV_13 $T=34040 459680 0 0 $X=33850 $Y=459440
X1256 1 2 378 385 20 392 24 406 ICV_13 $T=45540 459680 0 0 $X=45350 $Y=459440
X1257 1 2 413 420 21 404 7 413 ICV_13 $T=51520 476000 1 0 $X=51330 $Y=473040
X1258 1 2 441 436 20 392 8 438 ICV_13 $T=63480 465120 1 0 $X=63290 $Y=462160
X1259 1 2 439 436 25 429 13 439 ICV_13 $T=63480 481440 1 0 $X=63290 $Y=478480
X1260 1 2 446 50 32 47 24 446 ICV_13 $T=65320 443360 0 0 $X=65130 $Y=443120
X1261 1 2 455 436 27 429 15 455 ICV_13 $T=71760 476000 0 0 $X=71570 $Y=475760
X1262 1 2 468 50 20 47 8 468 ICV_13 $T=76820 443360 0 0 $X=76630 $Y=443120
X1263 1 2 492 60 28 57 19 492 ICV_13 $T=90160 443360 0 0 $X=89970 $Y=443120
X1264 1 2 494 470 25 457 13 494 ICV_13 $T=90160 470560 0 0 $X=89970 $Y=470320
X1265 1 2 486 484 27 474 7 490 ICV_13 $T=90160 481440 0 0 $X=89970 $Y=481200
X1266 1 2 497 484 22 474 24 480 ICV_13 $T=90160 486880 0 0 $X=89970 $Y=486640
X1267 1 2 495 459 20 445 8 495 ICV_13 $T=90620 497760 1 0 $X=90430 $Y=494800
X1268 1 2 519 64 25 58 13 519 ICV_13 $T=103500 448800 0 0 $X=103310 $Y=448560
X1269 1 2 521 64 21 58 7 521 ICV_13 $T=104420 448800 1 0 $X=104230 $Y=445840
X1270 1 2 548 533 30 536 7 549 ICV_13 $T=118220 486880 0 0 $X=118030 $Y=486640
X1271 1 2 550 533 25 536 13 550 ICV_13 $T=118220 492320 0 0 $X=118030 $Y=492080
X1272 1 2 551 533 32 536 24 551 ICV_13 $T=118220 497760 0 0 $X=118030 $Y=497520
X1273 1 2 552 533 22 536 9 552 ICV_13 $T=118220 503200 0 0 $X=118030 $Y=502960
X1274 1 2 569 568 20 559 8 569 ICV_13 $T=127880 465120 0 0 $X=127690 $Y=464880
X1275 1 2 571 561 30 547 26 571 ICV_13 $T=129260 470560 0 0 $X=129070 $Y=470320
X1276 1 2 576 579 25 563 13 576 ICV_13 $T=132480 486880 1 0 $X=132290 $Y=483920
X1277 1 2 578 579 21 563 8 577 ICV_13 $T=132480 492320 1 0 $X=132290 $Y=489360
X1278 1 2 580 579 28 563 19 580 ICV_13 $T=132480 503200 1 0 $X=132290 $Y=500240
X1279 1 2 589 568 25 559 13 589 ICV_13 $T=137080 459680 1 0 $X=136890 $Y=456720
X1280 1 2 592 568 30 559 26 592 ICV_13 $T=139840 454240 1 0 $X=139650 $Y=451280
X1281 1 2 601 597 28 588 9 598 ICV_13 $T=143520 508640 1 0 $X=143330 $Y=505680
X1282 1 2 609 618 92 594 83 609 ICV_13 $T=147660 481440 1 0 $X=147470 $Y=478480
X1283 1 2 611 603 93 81 82 611 ICV_13 $T=148580 448800 1 0 $X=148390 $Y=445840
X1284 1 2 613 91 96 84 86 613 ICV_13 $T=149040 443360 0 0 $X=148850 $Y=443120
X1285 1 2 620 603 96 81 86 620 ICV_13 $T=149500 448800 0 0 $X=149310 $Y=448560
X1286 1 2 633 616 102 593 95 633 ICV_13 $T=159160 459680 0 0 $X=158970 $Y=459440
X1287 1 2 637 603 102 81 95 637 ICV_13 $T=160540 454240 1 0 $X=160350 $Y=451280
X1288 1 2 639 618 101 594 99 639 ICV_13 $T=160540 486880 1 0 $X=160350 $Y=483920
X1289 1 2 641 630 25 619 13 641 ICV_13 $T=160540 497760 1 0 $X=160350 $Y=494800
X1290 1 2 644 603 103 81 97 644 ICV_13 $T=161920 443360 0 0 $X=161730 $Y=443120
X1291 1 2 648 630 32 619 24 648 ICV_13 $T=163760 508640 1 0 $X=163570 $Y=505680
X1292 1 2 668 663 96 635 86 668 ICV_13 $T=174340 470560 0 0 $X=174150 $Y=470320
X1293 1 2 656 663 92 635 97 669 ICV_13 $T=174340 481440 0 0 $X=174150 $Y=481200
X1294 1 2 657 624 27 636 24 683 ICV_13 $T=181700 497760 0 0 $X=181510 $Y=497520
X1295 1 2 712 689 28 665 19 712 ICV_13 $T=195040 508640 1 0 $X=194850 $Y=505680
X1296 1 2 726 704 28 690 19 726 ICV_13 $T=204240 454240 1 0 $X=204050 $Y=451280
X1297 1 2 747 736 27 720 15 747 ICV_13 $T=215740 497760 0 0 $X=215550 $Y=497520
X1298 1 2 751 752 103 718 82 748 ICV_13 $T=216660 459680 1 0 $X=216470 $Y=456720
X1299 1 2 750 734 101 719 24 731 ICV_13 $T=216660 476000 1 0 $X=216470 $Y=473040
X1300 1 2 755 752 102 746 97 751 ICV_13 $T=218500 454240 0 0 $X=218310 $Y=454000
X1301 1 2 763 736 20 720 8 763 ICV_13 $T=222180 503200 1 0 $X=221990 $Y=500240
X1302 1 2 767 732 30 722 26 767 ICV_13 $T=224020 492320 1 0 $X=223830 $Y=489360
X1303 1 2 776 752 94 746 98 775 ICV_13 $T=230460 448800 0 0 $X=230270 $Y=448560
X1304 1 2 779 781 96 768 98 778 ICV_13 $T=232760 459680 0 0 $X=232570 $Y=459440
X1305 1 2 783 769 93 762 82 783 ICV_13 $T=234140 476000 0 0 $X=233950 $Y=475760
X1306 1 2 797 133 101 768 82 796 ICV_13 $T=244720 459680 1 0 $X=244530 $Y=456720
X1307 1 2 792 769 102 768 99 803 ICV_13 $T=245180 470560 0 0 $X=244990 $Y=470320
X1308 1 2 822 133 96 786 86 822 ICV_13 $T=258520 448800 0 0 $X=258330 $Y=448560
X1309 1 2 823 808 103 813 97 823 ICV_13 $T=258520 459680 0 0 $X=258330 $Y=459440
X1310 1 2 824 808 94 813 85 824 ICV_13 $T=258520 465120 1 0 $X=258330 $Y=462160
X1311 1 2 837 808 96 813 95 841 ICV_13 $T=272780 465120 1 0 $X=272590 $Y=462160
X1312 1 2 859 864 102 851 95 859 ICV_13 $T=286580 459680 0 0 $X=286390 $Y=459440
X1313 1 2 862 826 92 817 83 862 ICV_13 $T=287040 470560 1 0 $X=286850 $Y=467600
X1314 1 2 858 847 96 833 85 865 ICV_13 $T=288420 448800 0 0 $X=288230 $Y=448560
X1315 1 2 866 847 92 833 83 866 ICV_13 $T=288420 454240 1 0 $X=288230 $Y=451280
X1316 1 2 852 839 96 831 95 856 ICV_13 $T=288420 476000 1 0 $X=288230 $Y=473040
X1317 1 2 877 876 94 855 85 877 ICV_13 $T=297160 476000 0 0 $X=296970 $Y=475760
X1318 1 2 879 864 92 851 83 879 ICV_13 $T=300840 459680 1 0 $X=300650 $Y=456720
X1319 1 2 881 864 93 851 82 881 ICV_13 $T=300840 470560 1 0 $X=300650 $Y=467600
X1320 1 2 882 864 103 851 97 882 ICV_13 $T=302680 465120 1 0 $X=302490 $Y=462160
X1321 1 2 888 890 101 140 82 148 ICV_13 $T=308200 448800 1 0 $X=308010 $Y=445840
X1322 1 2 912 890 92 878 83 912 ICV_13 $T=317860 448800 0 0 $X=317670 $Y=448560
X1323 1 2 918 903 157 875 150 918 ICV_13 $T=321080 492320 0 0 $X=320890 $Y=492080
X1324 1 2 922 925 157 904 150 922 ICV_13 $T=321540 503200 0 0 $X=321350 $Y=502960
X1325 1 2 910 890 89 153 150 158 ICV_13 $T=322000 443360 0 0 $X=321810 $Y=443120
X1326 1 2 923 902 157 884 150 923 ICV_13 $T=322460 486880 0 0 $X=322270 $Y=486640
X1327 1 2 927 915 155 898 149 927 ICV_13 $T=324300 481440 0 0 $X=324110 $Y=481200
X1328 1 2 966 902 167 884 159 966 ICV_13 $T=342700 486880 0 0 $X=342510 $Y=486640
X1329 1 2 946 945 152 926 165 973 ICV_13 $T=345920 454240 0 0 $X=345730 $Y=454000
X1330 1 2 977 958 164 943 149 979 ICV_13 $T=350060 470560 0 0 $X=349870 $Y=470320
X1331 1 2 981 958 151 943 146 981 ICV_13 $T=350980 459680 0 0 $X=350790 $Y=459440
X1332 1 2 992 994 151 978 146 992 ICV_13 $T=356960 492320 1 0 $X=356770 $Y=489360
X1333 1 2 996 184 152 182 144 996 ICV_13 $T=358800 443360 0 0 $X=358610 $Y=443120
X1334 1 2 1005 972 155 968 149 1005 ICV_13 $T=361560 497760 1 0 $X=361370 $Y=494800
X1335 1 2 985 915 152 990 165 1012 ICV_13 $T=363400 481440 1 0 $X=363210 $Y=478480
X1336 1 2 999 1000 151 988 165 998 ICV_13 $T=367540 459680 1 0 $X=367350 $Y=456720
X1337 1 2 1026 184 155 182 149 1026 ICV_13 $T=370760 443360 0 0 $X=370570 $Y=443120
X1338 1 2 1024 994 156 978 150 1028 ICV_13 $T=370760 486880 0 0 $X=370570 $Y=486640
X1339 1 2 1038 1014 151 989 146 1038 ICV_13 $T=375820 476000 0 0 $X=375630 $Y=475760
X1340 1 2 1041 1021 167 1019 159 1041 ICV_13 $T=376740 514080 1 0 $X=376550 $Y=511120
X1341 1 2 1058 994 152 978 144 1058 ICV_13 $T=385020 492320 1 0 $X=384830 $Y=489360
X1342 1 2 1071 1046 157 1025 150 1071 ICV_13 $T=391460 448800 1 0 $X=391270 $Y=445840
X1343 1 2 1089 1046 164 1025 165 1089 ICV_13 $T=398820 454240 1 0 $X=398630 $Y=451280
X1344 1 2 1084 1080 156 1067 149 1090 ICV_13 $T=398820 476000 0 0 $X=398630 $Y=475760
X1345 1 2 1128 1105 167 1086 144 1123 ICV_13 $T=413080 497760 1 0 $X=412890 $Y=494800
X1346 1 2 1155 210 155 208 149 1155 ICV_13 $T=428720 443360 0 0 $X=428530 $Y=443120
X1347 1 2 1156 210 167 208 159 1156 ICV_13 $T=428720 454240 1 0 $X=428530 $Y=451280
X1348 1 2 1150 1143 156 1118 144 1141 ICV_13 $T=429180 492320 1 0 $X=428990 $Y=489360
X1349 1 2 1163 1142 152 1130 144 1163 ICV_13 $T=431020 465120 0 0 $X=430830 $Y=464880
X1350 1 2 1162 1142 156 1130 146 1168 ICV_13 $T=431940 476000 0 0 $X=431750 $Y=475760
X1351 1 2 1169 1143 155 1118 149 1169 ICV_13 $T=431940 481440 0 0 $X=431750 $Y=481200
X1352 1 2 1167 1138 170 1152 159 1144 ICV_13 $T=433780 514080 1 0 $X=433590 $Y=511120
X1353 1 2 1175 1176 156 1153 154 1175 ICV_13 $T=434240 459680 0 0 $X=434050 $Y=459440
X1354 1 2 1186 210 164 1153 149 1196 ICV_13 $T=447120 454240 1 0 $X=446930 $Y=451280
X1355 1 2 1194 1205 170 1184 159 1201 ICV_13 $T=448040 514080 1 0 $X=447850 $Y=511120
X1356 1 2 1224 1216 156 1180 159 1128 ICV_13 $T=455860 492320 0 0 $X=455670 $Y=492080
X1357 1 2 1207 1199 164 1214 149 1233 ICV_13 $T=462300 465120 0 0 $X=462110 $Y=464880
X1358 1 2 1248 1231 164 1232 161 1244 ICV_13 $T=467360 492320 0 0 $X=467170 $Y=492080
X1359 1 2 1250 1230 164 1232 165 1250 ICV_13 $T=469200 481440 1 0 $X=469010 $Y=478480
X1360 1 2 1251 1231 152 1225 146 1252 ICV_13 $T=469200 503200 1 0 $X=469010 $Y=500240
X1361 1 2 1238 1231 157 1225 161 1229 ICV_13 $T=469200 508640 1 0 $X=469010 $Y=505680
X1362 1 2 1234 1239 152 1213 146 1249 ICV_13 $T=470580 448800 0 0 $X=470390 $Y=448560
X1363 1 2 1253 1239 167 1213 159 1253 ICV_13 $T=470580 454240 0 0 $X=470390 $Y=454000
X1364 1 2 1274 1276 151 1261 146 1274 ICV_13 $T=484380 497760 1 0 $X=484190 $Y=494800
X1365 1 2 1286 1282 155 1265 149 1286 ICV_13 $T=488520 459680 0 0 $X=488330 $Y=459440
X1366 1 2 1287 1282 156 1265 154 1287 ICV_13 $T=488520 465120 0 0 $X=488330 $Y=464880
X1367 1 2 1320 1324 170 1290 165 1319 ICV_13 $T=501400 459680 1 0 $X=501210 $Y=456720
X1368 1 2 1326 1322 157 1297 150 1326 ICV_13 $T=511060 508640 1 0 $X=510870 $Y=505680
X1369 1 2 1330 1322 155 1297 149 1330 ICV_13 $T=511520 503200 1 0 $X=511330 $Y=500240
X1370 1 2 1332 1325 157 1296 154 1333 ICV_13 $T=511980 497760 1 0 $X=511790 $Y=494800
X1371 1 2 1334 1304 157 1290 150 1334 ICV_13 $T=512440 448800 0 0 $X=512250 $Y=448560
X1372 1 2 1333 1325 156 1296 144 1336 ICV_13 $T=512440 492320 1 0 $X=512250 $Y=489360
X1373 1 2 1340 1304 156 1290 144 1323 ICV_13 $T=512900 454240 1 0 $X=512710 $Y=451280
X1374 1 2 1338 1293 155 1298 149 1338 ICV_13 $T=512900 476000 1 0 $X=512710 $Y=473040
X1375 1 2 1390 1365 262 1355 256 1390 ICV_13 $T=539120 459680 0 0 $X=538930 $Y=459440
X1376 1 2 1381 1378 264 1375 263 1377 ICV_13 $T=539120 503200 0 0 $X=538930 $Y=502960
X1377 1 2 1420 1378 262 1375 256 1420 ICV_13 $T=553380 503200 1 0 $X=553190 $Y=500240
X1378 1 2 1421 1378 255 1375 258 1421 ICV_13 $T=553380 508640 1 0 $X=553190 $Y=505680
X1379 1 2 1428 1409 269 1386 263 1428 ICV_13 $T=558440 459680 1 0 $X=558250 $Y=456720
X1380 1 2 1431 1409 262 1386 257 1429 ICV_13 $T=558440 465120 1 0 $X=558250 $Y=462160
X1381 1 2 1433 1412 262 1397 256 1433 ICV_13 $T=560280 470560 1 0 $X=560090 $Y=467600
X1382 1 2 1445 279 266 277 259 1445 ICV_13 $T=566720 454240 1 0 $X=566530 $Y=451280
X1383 1 2 1426 1418 269 1411 267 1447 ICV_13 $T=567180 486880 1 0 $X=566990 $Y=483920
X1384 1 2 1451 1418 270 1411 265 1451 ICV_13 $T=568100 486880 0 0 $X=567910 $Y=486640
X1385 1 2 1458 1438 266 1424 267 1455 ICV_13 $T=574540 497760 0 0 $X=574350 $Y=497520
X1386 1 2 1492 1456 264 1446 257 1492 ICV_13 $T=587880 476000 1 0 $X=587690 $Y=473040
X1387 1 2 1499 1495 264 1472 257 1499 ICV_13 $T=593400 503200 1 0 $X=593210 $Y=500240
X1388 1 2 1482 283 266 1474 265 1500 ICV_13 $T=593860 454240 1 0 $X=593670 $Y=451280
X1389 1 2 1501 1495 268 1472 261 1501 ICV_13 $T=593860 508640 1 0 $X=593670 $Y=505680
X1390 1 2 1504 283 269 1474 267 1502 ICV_13 $T=595240 448800 0 0 $X=595050 $Y=448560
X1391 1 2 1503 1495 275 1472 267 1503 ICV_13 $T=595240 497760 0 0 $X=595050 $Y=497520
X1392 1 2 1500 283 270 1474 263 1504 ICV_13 $T=596160 454240 0 0 $X=595970 $Y=454000
X1393 1 2 1507 1476 266 1463 259 1507 ICV_13 $T=597540 492320 1 0 $X=597350 $Y=489360
X1394 1 2 1513 1516 275 1523 267 1532 ICV_13 $T=609500 459680 1 0 $X=609310 $Y=456720
X1395 1 2 1533 1524 262 1520 256 1533 ICV_13 $T=609500 503200 1 0 $X=609310 $Y=500240
X1396 1 2 1539 1524 266 1520 259 1539 ICV_13 $T=610880 492320 0 0 $X=610690 $Y=492080
X1397 1 2 1552 1553 275 1527 263 1559 ICV_13 $T=623300 465120 0 0 $X=623110 $Y=464880
X1398 1 2 1566 1544 269 1525 263 1566 ICV_13 $T=623300 476000 0 0 $X=623110 $Y=475760
X1399 1 2 1560 1556 268 1550 258 1555 ICV_13 $T=623300 503200 0 0 $X=623110 $Y=502960
X1400 1 2 1567 1544 270 1525 265 1567 ICV_13 $T=623760 486880 1 0 $X=623570 $Y=483920
X1401 1 2 1582 1556 264 1550 257 1582 ICV_13 $T=630660 492320 0 0 $X=630470 $Y=492080
X1402 1 2 1586 1592 264 1578 257 1586 ICV_13 $T=635260 486880 0 0 $X=635070 $Y=486640
X1403 1 2 1608 1613 255 1588 258 1608 ICV_13 $T=643540 503200 1 0 $X=643350 $Y=500240
X1404 1 2 1605 1563 262 1576 265 1611 ICV_13 $T=644920 470560 1 0 $X=644730 $Y=467600
X1405 1 2 1624 1613 275 1588 267 1624 ICV_13 $T=652280 492320 1 0 $X=652090 $Y=489360
X1406 1 2 1634 1622 268 1620 267 1641 ICV_13 $T=659180 486880 0 0 $X=658990 $Y=486640
X1407 1 2 1639 1631 264 1620 263 1629 ICV_13 $T=665620 497760 1 0 $X=665430 $Y=494800
X1408 1 2 1659 1658 268 1649 261 1659 ICV_13 $T=670680 503200 1 0 $X=670490 $Y=500240
X1409 1 2 1690 1658 275 1649 267 1690 ICV_13 $T=686780 492320 0 0 $X=686590 $Y=492080
X1410 1 2 1700 1679 268 1668 267 1699 ICV_13 $T=691840 459680 0 0 $X=691650 $Y=459440
X1411 1 2 1701 308 262 1672 256 1701 ICV_13 $T=693680 443360 0 0 $X=693490 $Y=443120
X1412 1 2 1694 1679 264 1668 258 1696 ICV_13 $T=693680 470560 1 0 $X=693490 $Y=467600
X1413 1 2 1712 308 266 1672 259 1712 ICV_13 $T=696900 454240 1 0 $X=696710 $Y=451280
X1414 1 2 1724 1705 264 1691 257 1724 ICV_13 $T=703800 497760 1 0 $X=703610 $Y=494800
X1415 1 2 1725 1733 270 1719 265 1725 ICV_13 $T=707480 465120 0 0 $X=707290 $Y=464880
X1416 1 2 1727 1705 275 1691 267 1727 ICV_13 $T=707480 497760 0 0 $X=707290 $Y=497520
X1417 1 2 1728 1705 268 1691 261 1728 ICV_13 $T=707480 503200 0 0 $X=707290 $Y=502960
X1418 1 2 1731 1738 262 1720 256 1731 ICV_13 $T=708400 492320 1 0 $X=708210 $Y=489360
X1419 1 2 1745 1744 264 313 265 316 ICV_13 $T=709780 443360 0 0 $X=709590 $Y=443120
X1420 1 2 1739 1744 270 1721 265 1739 ICV_13 $T=709780 454240 0 0 $X=709590 $Y=454000
X1421 1 2 1748 1744 275 1721 267 1748 ICV_13 $T=721740 454240 1 0 $X=721550 $Y=451280
X1422 1 2 1749 1733 275 1719 267 1749 ICV_13 $T=721740 470560 1 0 $X=721550 $Y=467600
X1423 1 2 1752 1742 275 1722 267 1752 ICV_13 $T=721740 481440 1 0 $X=721550 $Y=478480
X1424 1 2 1755 1733 266 1719 259 1755 ICV_13 $T=722200 465120 0 0 $X=722010 $Y=464880
X1425 1 2 1762 317 255 313 267 1757 ICV_13 $T=722660 448800 1 0 $X=722470 $Y=445840
X1426 1 2 325 19 353 353 339 28 ICV_14 $T=17480 465120 0 0 $X=17290 $Y=464880
X1427 1 2 370 9 384 389 385 27 ICV_14 $T=32200 470560 1 0 $X=32010 $Y=467600
X1428 1 2 371 19 400 402 382 27 ICV_14 $T=41400 497760 0 0 $X=41210 $Y=497520
X1429 1 2 404 9 415 415 420 22 ICV_14 $T=50600 486880 1 0 $X=50410 $Y=483920
X1430 1 2 404 19 417 417 420 28 ICV_14 $T=51060 470560 1 0 $X=50870 $Y=467600
X1431 1 2 407 19 432 432 428 28 ICV_14 $T=57500 503200 1 0 $X=57310 $Y=500240
X1432 1 2 445 13 458 458 459 25 ICV_14 $T=71300 486880 0 0 $X=71110 $Y=486640
X1433 1 2 536 15 545 545 533 27 ICV_14 $T=116380 497760 1 0 $X=116190 $Y=494800
X1434 1 2 536 19 546 546 533 28 ICV_14 $T=116380 503200 1 0 $X=116190 $Y=500240
X1435 1 2 511 15 553 553 513 27 ICV_14 $T=117760 459680 1 0 $X=117570 $Y=456720
X1436 1 2 682 99 699 699 705 101 ICV_14 $T=189520 486880 0 0 $X=189330 $Y=486640
X1437 1 2 719 19 742 742 735 28 ICV_14 $T=206540 476000 0 0 $X=206350 $Y=475760
X1438 1 2 718 86 753 748 734 93 ICV_14 $T=217120 459680 0 0 $X=216930 $Y=459440
X1439 1 2 786 98 132 799 133 103 ICV_14 $T=243340 443360 0 0 $X=243150 $Y=443120
X1440 1 2 895 149 908 908 897 155 ICV_14 $T=316020 470560 1 0 $X=315830 $Y=467600
X1441 1 2 943 150 982 982 958 157 ICV_14 $T=350060 465120 0 0 $X=349870 $Y=464880
X1442 1 2 1073 159 1094 1094 1095 167 ICV_14 $T=398820 486880 1 0 $X=398630 $Y=483920
X1443 1 2 1067 150 1115 1117 1095 170 ICV_14 $T=410320 476000 0 0 $X=410130 $Y=475760
X1444 1 2 1184 144 1202 1193 1205 156 ICV_14 $T=447580 503200 1 0 $X=447390 $Y=500240
X1445 1 2 1299 150 1345 1345 1324 157 ICV_14 $T=513360 459680 0 0 $X=513170 $Y=459440
X1446 1 2 1355 259 1361 1361 1365 266 ICV_14 $T=525780 459680 0 0 $X=525590 $Y=459440
X1447 1 2 1375 267 1415 1415 1378 275 ICV_14 $T=550620 503200 0 0 $X=550430 $Y=502960
X1448 1 2 271 257 1423 1423 273 264 ICV_14 $T=553380 448800 1 0 $X=553190 $Y=445840
X1449 1 2 277 265 1444 1444 279 270 ICV_14 $T=565800 448800 1 0 $X=565610 $Y=445840
X1450 1 2 1411 258 1450 1450 1418 255 ICV_14 $T=566720 492320 1 0 $X=566530 $Y=489360
X1451 1 2 1520 263 1529 1529 1524 269 ICV_14 $T=606740 497760 0 0 $X=606550 $Y=497520
X1452 1 2 1520 257 1531 1531 1524 264 ICV_14 $T=608120 503200 0 0 $X=607930 $Y=502960
X1453 1 2 1722 256 1730 1734 1742 270 ICV_14 $T=707480 476000 0 0 $X=707290 $Y=475760
X1454 1 2 1720 267 1761 1761 1738 275 ICV_14 $T=721740 492320 1 0 $X=721550 $Y=489360
X1455 1 2 29 18 32 3 19 347 347 18 28 ICV_15 $T=15640 443360 0 0 $X=15450 $Y=443120
X1456 1 2 451 448 22 433 9 451 450 448 25 ICV_15 $T=66240 459680 0 0 $X=66050 $Y=459440
X1457 1 2 496 470 20 457 15 493 493 470 27 ICV_15 $T=90160 465120 0 0 $X=89970 $Y=464880
X1458 1 2 508 485 28 464 13 505 505 485 25 ICV_15 $T=94300 454240 0 0 $X=94110 $Y=454000
X1459 1 2 506 504 20 487 8 506 503 504 21 ICV_15 $T=94300 497760 0 0 $X=94110 $Y=497520
X1460 1 2 514 484 30 474 26 514 516 484 25 ICV_15 $T=101660 486880 0 0 $X=101470 $Y=486640
X1461 1 2 73 72 21 58 19 539 540 64 32 ICV_15 $T=118220 448800 0 0 $X=118030 $Y=448560
X1462 1 2 623 624 20 588 7 605 604 597 30 ICV_15 $T=146280 486880 0 0 $X=146090 $Y=486640
X1463 1 2 729 704 22 690 9 729 723 704 21 ICV_15 $T=205620 443360 0 0 $X=205430 $Y=443120
X1464 1 2 842 839 89 831 82 838 838 839 93 ICV_15 $T=270020 476000 0 0 $X=269830 $Y=475760
X1465 1 2 854 839 94 831 85 854 856 839 102 ICV_15 $T=281980 481440 1 0 $X=281790 $Y=478480
X1466 1 2 907 890 93 878 86 906 906 890 96 ICV_15 $T=315560 454240 0 0 $X=315370 $Y=454000
X1467 1 2 1009 1000 170 988 150 1018 1018 1000 157 ICV_15 $T=366160 465120 1 0 $X=365970 $Y=462160
X1468 1 2 1266 1239 164 1213 154 1270 1270 1239 156 ICV_15 $T=483000 454240 0 0 $X=482810 $Y=454000
X1469 1 2 1323 1304 152 1290 161 1301 1303 1304 167 ICV_15 $T=497260 454240 1 0 $X=497070 $Y=451280
X1470 1 2 1373 1354 262 1358 256 1373 1366 1371 262 ICV_15 $T=529460 492320 1 0 $X=529270 $Y=489360
X1471 1 2 1401 1409 268 1397 258 1414 1414 1412 255 ICV_15 $T=550620 465120 0 0 $X=550430 $Y=464880
X1472 1 2 1448 1438 269 1424 256 1440 1440 1438 262 ICV_15 $T=564880 503200 1 0 $X=564690 $Y=500240
X1473 1 2 1573 1575 275 1523 261 1558 1561 1563 275 ICV_15 $T=621460 454240 1 0 $X=621270 $Y=451280
X1474 1 2 1598 1592 275 1578 267 1598 1587 1592 262 ICV_15 $T=640320 486880 1 0 $X=640130 $Y=483920
X1475 1 2 1651 1622 275 1615 259 1643 1643 1622 266 ICV_15 $T=659640 476000 0 0 $X=659450 $Y=475760
X1476 1 2 1702 1692 270 1681 261 1695 1693 1692 266 ICV_15 $T=689080 481440 0 0 $X=688890 $Y=481200
X1477 1 2 1706 1705 269 1691 256 1703 1703 1705 262 ICV_15 $T=693680 503200 1 0 $X=693490 $Y=500240
X1478 1 2 1765 1738 269 1720 259 1753 1753 1738 266 ICV_15 $T=721740 486880 1 0 $X=721550 $Y=483920
X1479 1 2 3 15 350 350 18 27 ICV_16 $T=17020 448800 0 0 $X=16830 $Y=448560
X1480 1 2 325 24 361 361 339 32 ICV_16 $T=20240 470560 1 0 $X=20050 $Y=467600
X1481 1 2 445 7 465 465 459 21 ICV_16 $T=75440 492320 0 0 $X=75250 $Y=492080
X1482 1 2 58 9 515 515 64 22 ICV_16 $T=101660 443360 0 0 $X=101470 $Y=443120
X1483 1 2 487 26 525 524 504 25 ICV_16 $T=104420 497760 1 0 $X=104230 $Y=494800
X1484 1 2 487 19 526 526 504 28 ICV_16 $T=104420 503200 1 0 $X=104230 $Y=500240
X1485 1 2 511 24 522 523 529 20 ICV_16 $T=105800 465120 0 0 $X=105610 $Y=464880
X1486 1 2 588 8 600 598 597 22 ICV_16 $T=143980 503200 1 0 $X=143790 $Y=500240
X1487 1 2 588 26 604 605 597 21 ICV_16 $T=145360 486880 1 0 $X=145170 $Y=483920
X1488 1 2 682 95 698 703 705 89 ICV_16 $T=189980 476000 0 0 $X=189790 $Y=475760
X1489 1 2 719 13 738 738 735 25 ICV_16 $T=206540 481440 0 0 $X=206350 $Y=481200
X1490 1 2 722 9 794 791 732 21 ICV_16 $T=239200 492320 0 0 $X=239010 $Y=492080
X1491 1 2 768 97 804 802 781 94 ICV_16 $T=244720 470560 1 0 $X=244530 $Y=467600
X1492 1 2 798 83 830 827 812 103 ICV_16 $T=259900 486880 1 0 $X=259710 $Y=483920
X1493 1 2 831 83 840 840 839 92 ICV_16 $T=270940 481440 0 0 $X=270750 $Y=481200
X1494 1 2 817 86 863 863 826 96 ICV_16 $T=286580 470560 0 0 $X=286390 $Y=470320
X1495 1 2 878 99 888 887 890 102 ICV_16 $T=304980 454240 1 0 $X=304790 $Y=451280
X1496 1 2 895 159 934 936 897 170 ICV_16 $T=327520 470560 0 0 $X=327330 $Y=470320
X1497 1 2 926 150 967 967 945 157 ICV_16 $T=344080 454240 1 0 $X=343890 $Y=451280
X1498 1 2 1034 150 1075 1069 1051 156 ICV_16 $T=392380 465120 1 0 $X=392190 $Y=462160
X1499 1 2 1067 144 1096 1074 1051 152 ICV_16 $T=399740 470560 1 0 $X=399550 $Y=467600
X1500 1 2 1086 149 1125 1125 1129 155 ICV_16 $T=413080 497760 0 0 $X=412890 $Y=497520
X1501 1 2 1153 161 1187 1190 1199 155 ICV_16 $T=445280 465120 1 0 $X=445090 $Y=462160
X1502 1 2 1184 146 1204 1204 1205 151 ICV_16 $T=448960 497760 1 0 $X=448770 $Y=494800
X1503 1 2 219 154 1220 1220 225 156 ICV_16 $T=454940 443360 0 0 $X=454750 $Y=443120
X1504 1 2 1232 144 1255 1255 1230 152 ICV_16 $T=470580 470560 0 0 $X=470390 $Y=470320
X1505 1 2 1290 159 1303 1301 1304 170 ICV_16 $T=498640 454240 0 0 $X=498450 $Y=454000
X1506 1 2 1297 144 1331 1331 1322 152 ICV_16 $T=511060 503200 0 0 $X=510870 $Y=502960
X1507 1 2 245 154 252 1337 250 157 ICV_16 $T=512440 448800 1 0 $X=512250 $Y=445840
X1508 1 2 1355 265 1380 1380 1365 270 ICV_16 $T=535900 470560 1 0 $X=535710 $Y=467600
X1509 1 2 1463 258 1477 1477 1476 255 ICV_16 $T=581440 492320 1 0 $X=581250 $Y=489360
X1510 1 2 1497 259 1514 1502 283 275 ICV_16 $T=599380 459680 0 0 $X=599190 $Y=459440
X1511 1 2 1463 261 1512 1519 1476 264 ICV_16 $T=599380 486880 0 0 $X=599190 $Y=486640
X1512 1 2 1497 263 1522 1522 1516 269 ICV_16 $T=601680 470560 0 0 $X=601490 $Y=470320
X1513 1 2 1525 258 1568 1568 1544 255 ICV_16 $T=623300 486880 0 0 $X=623110 $Y=486640
X1514 1 2 1588 261 1609 1609 1613 268 ICV_16 $T=643080 508640 1 0 $X=642890 $Y=505680
X1515 1 2 1649 257 1667 1667 1658 264 ICV_16 $T=672520 492320 1 0 $X=672330 $Y=489360
X1516 1 2 1652 265 1673 1673 1661 270 ICV_16 $T=676200 486880 1 0 $X=676010 $Y=483920
X1517 1 2 1672 263 311 1687 1679 266 ICV_16 $T=683560 454240 0 0 $X=683370 $Y=454000
X1518 1 2 1722 265 1734 1730 1742 262 ICV_16 $T=708400 481440 1 0 $X=708210 $Y=478480
X1519 1 2 1722 261 1736 1736 1742 268 ICV_16 $T=708860 476000 1 0 $X=708670 $Y=473040
X1520 1 2 1722 258 1750 1750 1742 255 ICV_16 $T=721280 470560 0 0 $X=721090 $Y=470320
X1521 1 2 1722 263 1756 1756 1742 269 ICV_16 $T=721740 476000 1 0 $X=721550 $Y=473040
X1522 1 2 323 9 332 332 334 22 ICV_17 $T=5520 481440 1 0 $X=5330 $Y=478480
X1523 1 2 407 26 437 437 428 30 ICV_17 $T=60720 492320 1 0 $X=60530 $Y=489360
X1524 1 2 429 26 444 444 436 30 ICV_17 $T=63020 476000 1 0 $X=62830 $Y=473040
X1525 1 2 563 24 572 572 579 32 ICV_17 $T=129720 497760 0 0 $X=129530 $Y=497520
X1526 1 2 563 9 573 573 579 22 ICV_17 $T=129720 503200 0 0 $X=129530 $Y=502960
X1527 1 2 559 24 581 584 568 22 ICV_17 $T=132480 465120 1 0 $X=132290 $Y=462160
X1528 1 2 81 99 628 645 616 101 ICV_17 $T=160540 454240 0 0 $X=160350 $Y=454000
X1529 1 2 718 85 754 753 734 96 ICV_17 $T=216660 465120 1 0 $X=216470 $Y=462160
X1530 1 2 817 95 821 821 826 102 ICV_17 $T=256680 470560 1 0 $X=256490 $Y=467600
X1531 1 2 135 98 835 835 137 89 ICV_17 $T=266800 443360 0 0 $X=266610 $Y=443120
X1532 1 2 943 161 957 957 958 170 ICV_17 $T=339020 465120 1 0 $X=338830 $Y=462160
X1533 1 2 978 159 1059 1059 994 167 ICV_17 $T=383640 492320 0 0 $X=383450 $Y=492080
X1534 1 2 198 154 1109 1109 204 156 ICV_17 $T=407100 443360 0 0 $X=406910 $Y=443120
X1535 1 2 1067 165 1111 1114 1080 151 ICV_17 $T=408480 470560 0 0 $X=408290 $Y=470320
X1536 1 2 1130 165 1145 1135 1143 167 ICV_17 $T=420440 481440 1 0 $X=420250 $Y=478480
X1537 1 2 208 150 1154 1154 210 157 ICV_17 $T=426880 448800 0 0 $X=426690 $Y=448560
X1538 1 2 1153 144 1178 1172 1176 164 ICV_17 $T=434240 454240 0 0 $X=434050 $Y=454000
X1539 1 2 1180 146 1209 1212 1216 152 ICV_17 $T=451720 486880 1 0 $X=451530 $Y=483920
X1540 1 2 219 161 1245 1245 225 170 ICV_17 $T=466900 443360 0 0 $X=466710 $Y=443120
X1541 1 2 1296 149 1335 1335 1325 155 ICV_17 $T=511060 486880 0 0 $X=510870 $Y=486640
X1542 1 2 1353 261 1382 1362 1351 264 ICV_17 $T=535440 454240 1 0 $X=535250 $Y=451280
X1543 1 2 1397 265 1434 1434 1412 270 ICV_17 $T=560740 476000 1 0 $X=560550 $Y=473040
X1544 1 2 1443 258 1486 1488 1459 268 ICV_17 $T=585580 465120 1 0 $X=585390 $Y=462160
X1545 1 2 1443 261 1488 1487 1459 266 ICV_17 $T=585580 470560 1 0 $X=585390 $Y=467600
X1546 1 2 1474 256 1505 1505 283 262 ICV_17 $T=595240 443360 0 0 $X=595050 $Y=443120
X1547 1 2 1474 258 1506 1506 283 255 ICV_17 $T=596160 448800 1 0 $X=595970 $Y=445840
X1548 1 2 1523 259 1536 1536 287 266 ICV_17 $T=609040 448800 0 0 $X=608850 $Y=448560
X1549 1 2 1615 258 1625 1626 1622 264 ICV_17 $T=652280 481440 1 0 $X=652090 $Y=478480
X1550 1 2 1691 258 1723 1723 1705 255 ICV_17 $T=701040 508640 1 0 $X=700850 $Y=505680
X1551 1 2 1721 256 1732 1732 1744 262 ICV_17 $T=707480 448800 0 0 $X=707290 $Y=448560
X1552 1 2 1720 265 1735 1735 1738 270 ICV_17 $T=707480 486880 0 0 $X=707290 $Y=486640
X1553 1 2 1719 261 1740 1729 1733 262 ICV_17 $T=708400 465120 1 0 $X=708210 $Y=462160
X1554 1 2 1721 258 1759 1759 1744 255 ICV_17 $T=721280 454240 0 0 $X=721090 $Y=454000
X1555 1 2 1719 258 1760 1760 1733 255 ICV_17 $T=721280 459680 0 0 $X=721090 $Y=459440
X1556 1 2 1721 263 1763 1763 1744 269 ICV_17 $T=721740 459680 1 0 $X=721550 $Y=456720
X1557 1 2 1719 263 1764 1740 1733 268 ICV_17 $T=721740 465120 1 0 $X=721550 $Y=462160
X1574 1 2 41 24 409 398 35 22 ICV_19 $T=48300 448800 1 0 $X=48110 $Y=445840
X1575 1 2 563 26 574 574 579 30 ICV_19 $T=129720 492320 0 0 $X=129530 $Y=492080
X1576 1 2 635 99 664 669 663 103 ICV_19 $T=172040 486880 1 0 $X=171850 $Y=483920
X1577 1 2 109 99 111 112 113 96 ICV_19 $T=187680 443360 0 0 $X=187490 $Y=443120
X1578 1 2 675 99 717 715 685 103 ICV_19 $T=195960 459680 1 0 $X=195770 $Y=456720
X1579 1 2 722 15 728 743 732 25 ICV_19 $T=206540 492320 0 0 $X=206350 $Y=492080
X1580 1 2 719 9 756 756 735 22 ICV_19 $T=216660 486880 1 0 $X=216470 $Y=483920
X1581 1 2 746 83 774 774 752 92 ICV_19 $T=227240 454240 1 0 $X=227050 $Y=451280
X1582 1 2 813 82 828 819 133 94 ICV_19 $T=258520 454240 0 0 $X=258330 $Y=454000
X1583 1 2 884 161 962 962 902 170 ICV_19 $T=339940 486880 1 0 $X=339750 $Y=483920
X1584 1 2 978 149 991 991 994 155 ICV_19 $T=354200 486880 0 0 $X=354010 $Y=486640
X1585 1 2 1056 146 1078 1081 1065 156 ICV_19 $T=393300 503200 1 0 $X=393110 $Y=500240
X1586 1 2 1073 149 1087 1087 1095 155 ICV_19 $T=396520 492320 1 0 $X=396330 $Y=489360
X1587 1 2 1082 161 1120 1120 1107 170 ICV_19 $T=411240 454240 0 0 $X=411050 $Y=454000
X1588 1 2 1082 146 1121 1121 1107 151 ICV_19 $T=411240 459680 0 0 $X=411050 $Y=459440
X1589 1 2 198 159 1134 1134 204 167 ICV_19 $T=417220 448800 1 0 $X=417030 $Y=445840
X1590 1 2 219 159 1210 1210 225 167 ICV_19 $T=452180 448800 1 0 $X=451990 $Y=445840
X1591 1 2 1232 149 1256 1256 1230 155 ICV_19 $T=469200 476000 1 0 $X=469010 $Y=473040
X1592 1 2 1296 159 1310 1311 1322 164 ICV_19 $T=498640 497760 1 0 $X=498450 $Y=494800
X1593 1 2 1446 256 1469 1469 1456 262 ICV_19 $T=575460 476000 0 0 $X=575270 $Y=475760
X1594 1 2 1681 267 1698 1709 1692 264 ICV_19 $T=693680 486880 1 0 $X=693490 $Y=483920
X1595 1 2 1681 263 1714 1710 1692 262 ICV_19 $T=695060 481440 1 0 $X=694870 $Y=478480
X1596 1 2 1722 259 1751 1751 1742 266 ICV_19 $T=719900 476000 0 0 $X=719710 $Y=475760
X1597 1 2 313 258 1762 1743 317 264 ICV_19 $T=721280 443360 0 0 $X=721090 $Y=443120
X1598 1 2 370 8 378 ICV_20 $T=31740 459680 1 0 $X=31550 $Y=456720
X1599 1 2 371 13 380 ICV_20 $T=31740 492320 1 0 $X=31550 $Y=489360
X1600 1 2 371 9 381 ICV_20 $T=31740 497760 1 0 $X=31550 $Y=494800
X1601 1 2 355 19 394 ICV_20 $T=40020 481440 0 0 $X=39830 $Y=481200
X1602 1 2 407 15 421 ICV_20 $T=52900 492320 1 0 $X=52710 $Y=489360
X1603 1 2 392 13 427 ICV_20 $T=55660 465120 1 0 $X=55470 $Y=462160
X1604 1 2 433 13 450 ICV_20 $T=65780 459680 1 0 $X=65590 $Y=456720
X1605 1 2 464 24 477 ICV_20 $T=81880 448800 0 0 $X=81690 $Y=448560
X1606 1 2 464 9 478 ICV_20 $T=81880 459680 0 0 $X=81690 $Y=459440
X1607 1 2 457 19 491 ICV_20 $T=87400 476000 1 0 $X=87210 $Y=473040
X1608 1 2 457 8 496 ICV_20 $T=90620 470560 1 0 $X=90430 $Y=467600
X1609 1 2 464 15 501 ICV_20 $T=93840 459680 1 0 $X=93650 $Y=456720
X1610 1 2 464 8 502 ICV_20 $T=95680 465120 1 0 $X=95490 $Y=462160
X1611 1 2 69 19 583 ICV_20 $T=134320 448800 1 0 $X=134130 $Y=445840
X1612 1 2 69 13 77 ICV_20 $T=135700 443360 0 0 $X=135510 $Y=443120
X1613 1 2 593 83 615 ICV_20 $T=148580 459680 1 0 $X=148390 $Y=456720
X1614 1 2 593 86 621 ICV_20 $T=149040 465120 1 0 $X=148850 $Y=462160
X1615 1 2 81 83 642 ICV_20 $T=160540 448800 1 0 $X=160350 $Y=445840
X1616 1 2 81 98 602 ICV_20 $T=160540 459680 1 0 $X=160350 $Y=456720
X1617 1 2 593 97 647 ICV_20 $T=162380 465120 0 0 $X=162190 $Y=464880
X1618 1 2 649 97 659 ICV_20 $T=172040 454240 1 0 $X=171850 $Y=451280
X1619 1 2 682 86 695 ICV_20 $T=188600 476000 1 0 $X=188410 $Y=473040
X1620 1 2 690 8 708 ICV_20 $T=192740 454240 0 0 $X=192550 $Y=454000
X1621 1 2 675 83 714 ICV_20 $T=195960 470560 1 0 $X=195770 $Y=467600
X1622 1 2 675 97 715 ICV_20 $T=196880 465120 1 0 $X=196690 $Y=462160
X1623 1 2 719 26 758 ICV_20 $T=218960 476000 0 0 $X=218770 $Y=475760
X1624 1 2 746 85 776 ICV_20 $T=230460 454240 0 0 $X=230270 $Y=454000
X1625 1 2 768 95 801 ICV_20 $T=244260 459680 0 0 $X=244070 $Y=459440
X1626 1 2 798 95 810 ICV_20 $T=247940 476000 0 0 $X=247750 $Y=475760
X1627 1 2 817 99 825 ICV_20 $T=258520 470560 0 0 $X=258330 $Y=470320
X1628 1 2 798 86 829 ICV_20 $T=260360 476000 0 0 $X=260170 $Y=475760
X1629 1 2 831 86 852 ICV_20 $T=280600 476000 1 0 $X=280410 $Y=473040
X1630 1 2 817 82 861 ICV_20 $T=286580 465120 0 0 $X=286390 $Y=464880
X1631 1 2 140 99 142 ICV_20 $T=287960 443360 0 0 $X=287770 $Y=443120
X1632 1 2 140 97 870 ICV_20 $T=291180 448800 1 0 $X=290990 $Y=445840
X1633 1 2 875 144 885 ICV_20 $T=302680 497760 1 0 $X=302490 $Y=494800
X1634 1 2 884 149 905 ICV_20 $T=314640 486880 0 0 $X=314450 $Y=486640
X1635 1 2 878 98 910 ICV_20 $T=316940 454240 1 0 $X=316750 $Y=451280
X1636 1 2 875 149 919 ICV_20 $T=320620 497760 1 0 $X=320430 $Y=494800
X1637 1 2 926 159 939 ICV_20 $T=330740 448800 1 0 $X=330550 $Y=445840
X1638 1 2 926 146 942 ICV_20 $T=331200 454240 0 0 $X=331010 $Y=454000
X1639 1 2 875 154 948 ICV_20 $T=332580 492320 0 0 $X=332390 $Y=492080
X1640 1 2 153 159 975 ICV_20 $T=346840 448800 0 0 $X=346650 $Y=448560
X1641 1 2 968 165 969 ICV_20 $T=350980 503200 0 0 $X=350790 $Y=502960
X1642 1 2 989 161 1003 ICV_20 $T=361100 470560 1 0 $X=360910 $Y=467600
X1643 1 2 989 154 1004 ICV_20 $T=361100 476000 0 0 $X=360910 $Y=475760
X1644 1 2 988 161 1009 ICV_20 $T=362480 459680 0 0 $X=362290 $Y=459440
X1645 1 2 990 161 1013 ICV_20 $T=362940 486880 1 0 $X=362750 $Y=483920
X1646 1 2 989 159 1023 ICV_20 $T=368920 470560 1 0 $X=368730 $Y=467600
X1647 1 2 1019 149 1030 ICV_20 $T=373060 497760 1 0 $X=372870 $Y=494800
X1648 1 2 1019 146 1031 ICV_20 $T=373060 497760 0 0 $X=372870 $Y=497520
X1649 1 2 1025 159 1043 ICV_20 $T=376740 454240 1 0 $X=376550 $Y=451280
X1650 1 2 1034 146 1052 ICV_20 $T=381800 465120 0 0 $X=381610 $Y=464880
X1651 1 2 990 154 1054 ICV_20 $T=382260 486880 0 0 $X=382070 $Y=486640
X1652 1 2 1025 146 1072 ICV_20 $T=391000 454240 1 0 $X=390810 $Y=451280
X1653 1 2 1073 144 1092 ICV_20 $T=398820 492320 0 0 $X=398630 $Y=492080
X1654 1 2 1082 159 1100 ICV_20 $T=403420 459680 0 0 $X=403230 $Y=459440
X1655 1 2 1082 165 1102 ICV_20 $T=404340 465120 1 0 $X=404150 $Y=462160
X1656 1 2 1086 146 1126 ICV_20 $T=413080 503200 1 0 $X=412890 $Y=500240
X1657 1 2 198 149 1132 ICV_20 $T=416300 448800 0 0 $X=416110 $Y=448560
X1658 1 2 1152 154 1158 ICV_20 $T=429180 508640 1 0 $X=428990 $Y=505680
X1659 1 2 1152 149 1166 ICV_20 $T=431020 497760 1 0 $X=430830 $Y=494800
X1660 1 2 208 161 1185 ICV_20 $T=442980 448800 1 0 $X=442790 $Y=445840
X1661 1 2 1213 144 1234 ICV_20 $T=460920 454240 1 0 $X=460730 $Y=451280
X1662 1 2 1214 159 230 ICV_20 $T=462760 470560 0 0 $X=462570 $Y=470320
X1663 1 2 1214 150 1254 ICV_20 $T=473800 465120 0 0 $X=473610 $Y=464880
X1664 1 2 1261 150 1271 ICV_20 $T=483000 503200 0 0 $X=482810 $Y=502960
X1665 1 2 1297 161 1306 ICV_20 $T=499560 508640 0 0 $X=499370 $Y=508400
X1666 1 2 1298 159 1315 ICV_20 $T=500480 481440 0 0 $X=500290 $Y=481200
X1667 1 2 1298 154 1329 ICV_20 $T=511060 481440 0 0 $X=510870 $Y=481200
X1668 1 2 1358 263 1403 ICV_20 $T=545100 492320 1 0 $X=544910 $Y=489360
X1669 1 2 1443 257 1454 ICV_20 $T=571780 470560 1 0 $X=571590 $Y=467600
X1670 1 2 277 263 1461 ICV_20 $T=574540 448800 0 0 $X=574350 $Y=448560
X1671 1 2 1472 256 1481 ICV_20 $T=585580 503200 1 0 $X=585390 $Y=500240
X1672 1 2 1446 258 1489 ICV_20 $T=586500 470560 0 0 $X=586310 $Y=470320
X1673 1 2 1497 261 1509 ICV_20 $T=598460 470560 1 0 $X=598270 $Y=467600
X1674 1 2 1497 267 1513 ICV_20 $T=599380 459680 1 0 $X=599190 $Y=456720
X1675 1 2 1497 256 1517 ICV_20 $T=599840 481440 1 0 $X=599650 $Y=478480
X1676 1 2 1525 257 1540 ICV_20 $T=611340 486880 0 0 $X=611150 $Y=486640
X1677 1 2 1525 261 1542 ICV_20 $T=611800 481440 0 0 $X=611610 $Y=481200
X1678 1 2 1527 257 1548 ICV_20 $T=613640 470560 1 0 $X=613450 $Y=467600
X1679 1 2 1527 256 1554 ICV_20 $T=617780 465120 1 0 $X=617590 $Y=462160
X1680 1 2 1550 261 1560 ICV_20 $T=621000 503200 1 0 $X=620810 $Y=500240
X1681 1 2 1550 256 1579 ICV_20 $T=628820 503200 1 0 $X=628630 $Y=500240
X1682 1 2 1578 256 1587 ICV_20 $T=635260 481440 0 0 $X=635070 $Y=481200
X1683 1 2 1578 259 1596 ICV_20 $T=637560 476000 1 0 $X=637370 $Y=473040
X1684 1 2 1588 263 1601 ICV_20 $T=642160 492320 0 0 $X=641970 $Y=492080
X1685 1 2 1618 267 1632 ICV_20 $T=655040 465120 1 0 $X=654850 $Y=462160
X1686 1 2 1615 261 1634 ICV_20 $T=655960 486880 1 0 $X=655770 $Y=483920
X1687 1 2 1620 256 1636 ICV_20 $T=656880 497760 1 0 $X=656690 $Y=494800
X1688 1 2 1620 265 1644 ICV_20 $T=659180 503200 0 0 $X=658990 $Y=502960
X1689 1 2 300 265 1640 ICV_20 $T=659640 454240 0 0 $X=659450 $Y=454000
X1690 1 2 1615 265 1646 ICV_20 $T=661020 481440 0 0 $X=660830 $Y=481200
X1691 1 2 1691 259 1711 ICV_20 $T=695980 497760 1 0 $X=695790 $Y=494800
X1692 1 2 1719 256 1729 ICV_20 $T=707480 459680 0 0 $X=707290 $Y=459440
X1693 1 2 1720 261 1747 ICV_20 $T=711620 492320 0 0 $X=711430 $Y=492080
X1694 1 2 325 8 342 ICV_21 $T=6900 459680 1 0 $X=6710 $Y=456720
X1695 1 2 325 13 343 ICV_21 $T=6900 465120 0 0 $X=6710 $Y=464880
X1696 1 2 328 13 337 ICV_21 $T=6900 486880 0 0 $X=6710 $Y=486640
X1697 1 2 323 24 351 ICV_21 $T=14260 481440 0 0 $X=14070 $Y=481200
X1698 1 2 355 7 396 ICV_21 $T=36340 481440 1 0 $X=36150 $Y=478480
X1699 1 2 404 15 419 ICV_21 $T=49680 470560 0 0 $X=49490 $Y=470320
X1700 1 2 433 26 447 ICV_21 $T=62560 454240 1 0 $X=62370 $Y=451280
X1701 1 2 474 8 489 ICV_21 $T=83720 492320 1 0 $X=83530 $Y=489360
X1702 1 2 487 7 503 ICV_21 $T=90160 492320 0 0 $X=89970 $Y=492080
X1703 1 2 511 19 530 ICV_21 $T=103500 459680 0 0 $X=103310 $Y=459440
X1704 1 2 58 24 540 ICV_21 $T=111320 454240 1 0 $X=111130 $Y=451280
X1705 1 2 509 26 541 ICV_21 $T=111780 476000 1 0 $X=111590 $Y=473040
X1706 1 2 511 9 544 ICV_21 $T=113620 470560 1 0 $X=113430 $Y=467600
X1707 1 2 682 85 702 ICV_21 $T=188140 470560 0 0 $X=187950 $Y=470320
X1708 1 2 746 82 760 ICV_21 $T=216660 448800 1 0 $X=216470 $Y=445840
X1709 1 2 786 99 797 ICV_21 $T=238280 454240 0 0 $X=238090 $Y=454000
X1710 1 2 831 99 853 ICV_21 $T=278300 486880 1 0 $X=278110 $Y=483920
X1711 1 2 855 98 869 ICV_21 $T=286580 476000 0 0 $X=286390 $Y=475760
X1712 1 2 898 150 911 ICV_21 $T=314180 481440 1 0 $X=313990 $Y=478480
X1713 1 2 878 97 913 ICV_21 $T=314640 459680 0 0 $X=314450 $Y=459440
X1714 1 2 988 146 999 ICV_21 $T=356960 459680 1 0 $X=356770 $Y=456720
X1715 1 2 988 154 1002 ICV_21 $T=357420 454240 0 0 $X=357230 $Y=454000
X1716 1 2 1019 150 1033 ICV_21 $T=370760 503200 0 0 $X=370570 $Y=502960
X1717 1 2 1034 165 1050 ICV_21 $T=378120 459680 0 0 $X=377930 $Y=459440
X1718 1 2 1073 146 1112 ICV_21 $T=407100 481440 0 0 $X=406910 $Y=481200
X1719 1 2 1152 150 1160 ICV_21 $T=426880 503200 0 0 $X=426690 $Y=502960
X1720 1 2 1118 146 1159 ICV_21 $T=429180 486880 1 0 $X=428990 $Y=483920
X1721 1 2 1179 154 1195 ICV_21 $T=443440 476000 0 0 $X=443250 $Y=475760
X1722 1 2 1265 165 1279 ICV_21 $T=483000 470560 0 0 $X=482810 $Y=470320
X1723 1 2 1265 161 1281 ICV_21 $T=483000 476000 0 0 $X=482810 $Y=475760
X1724 1 2 1296 161 1305 ICV_21 $T=496800 492320 0 0 $X=496610 $Y=492080
X1725 1 2 1297 159 1312 ICV_21 $T=497260 508640 1 0 $X=497070 $Y=505680
X1726 1 2 1668 263 1683 ICV_21 $T=678960 465120 1 0 $X=678770 $Y=462160
X1727 1 2 1681 256 1710 ICV_21 $T=693220 476000 0 0 $X=693030 $Y=475760
X1728 1 2 1720 263 1765 ICV_21 $T=720360 486880 0 0 $X=720170 $Y=486640
X1729 1 2 323 19 349 349 334 28 ICV_22 $T=14260 470560 0 0 $X=14070 $Y=470320
X1730 1 2 429 7 443 443 436 21 ICV_22 $T=62100 470560 0 0 $X=61910 $Y=470320
X1731 1 2 433 24 453 453 448 32 ICV_22 $T=66240 454240 0 0 $X=66050 $Y=454000
X1732 1 2 635 95 661 661 663 102 ICV_22 $T=170200 476000 1 0 $X=170010 $Y=473040
X1733 1 2 665 13 700 700 689 25 ICV_22 $T=188600 497760 1 0 $X=188410 $Y=494800
X1734 1 2 665 15 711 711 689 27 ICV_22 $T=192740 503200 1 0 $X=192550 $Y=500240
X1735 1 2 718 99 750 749 734 103 ICV_22 $T=214360 470560 0 0 $X=214170 $Y=470320
X1736 1 2 817 97 836 836 826 103 ICV_22 $T=266340 470560 0 0 $X=266150 $Y=470320
X1737 1 2 817 98 843 841 808 102 ICV_22 $T=270940 465120 0 0 $X=270750 $Y=464880
X1738 1 2 833 98 845 846 847 101 ICV_22 $T=271860 454240 0 0 $X=271670 $Y=454000
X1739 1 2 851 85 860 860 864 94 ICV_22 $T=284280 465120 1 0 $X=284090 $Y=462160
X1740 1 2 884 144 899 891 876 103 ICV_22 $T=307740 486880 1 0 $X=307550 $Y=483920
X1741 1 2 926 154 940 940 945 156 ICV_22 $T=328900 459680 1 0 $X=328710 $Y=456720
X1742 1 2 926 161 970 970 945 170 ICV_22 $T=342700 459680 1 0 $X=342510 $Y=456720
X1743 1 2 990 150 1061 1061 1016 157 ICV_22 $T=385020 486880 1 0 $X=384830 $Y=483920
X1744 1 2 1056 159 1076 1076 1065 167 ICV_22 $T=391000 514080 1 0 $X=390810 $Y=511120
X1745 1 2 1290 154 1340 1344 1324 155 ICV_22 $T=511060 454240 0 0 $X=510870 $Y=454000
X1746 1 2 1353 257 1362 1360 1351 266 ICV_22 $T=524860 454240 0 0 $X=524670 $Y=454000
X1747 1 2 1356 263 1384 1384 1371 269 ICV_22 $T=535440 486880 1 0 $X=535250 $Y=483920
X1748 1 2 1618 256 1637 1637 1619 262 ICV_22 $T=655500 465120 0 0 $X=655310 $Y=464880
X1749 1 2 1618 263 1654 1654 1619 269 ICV_22 $T=665620 459680 1 0 $X=665430 $Y=456720
X1750 1 2 1719 257 1726 1726 1733 264 ICV_22 $T=705180 470560 1 0 $X=704990 $Y=467600
X1751 1 2 1720 257 1737 1737 1738 264 ICV_22 $T=707020 486880 1 0 $X=706830 $Y=483920
X1752 1 2 1722 257 1741 1741 1742 264 ICV_22 $T=707480 470560 0 0 $X=707290 $Y=470320
X1753 1 2 1720 258 1754 1754 1738 255 ICV_22 $T=719440 492320 0 0 $X=719250 $Y=492080
X1754 1 2 1721 259 1758 1758 1744 266 ICV_22 $T=720360 448800 0 0 $X=720170 $Y=448560
X1755 1 2 ICV_23 $T=18400 448800 1 0 $X=18210 $Y=445840
X1756 1 2 ICV_23 $T=88320 443360 0 0 $X=88130 $Y=443120
X1757 1 2 ICV_23 $T=88320 503200 0 0 $X=88130 $Y=502960
X1758 1 2 ICV_23 $T=102580 448800 1 0 $X=102390 $Y=445840
X1759 1 2 ICV_23 $T=116380 508640 0 0 $X=116190 $Y=508400
X1760 1 2 ICV_23 $T=158700 459680 1 0 $X=158510 $Y=456720
X1761 1 2 ICV_23 $T=158700 508640 1 0 $X=158510 $Y=505680
X1762 1 2 ICV_23 $T=200560 454240 0 0 $X=200370 $Y=454000
X1763 1 2 ICV_23 $T=214820 465120 1 0 $X=214630 $Y=462160
X1764 1 2 ICV_23 $T=242880 454240 1 0 $X=242690 $Y=451280
X1765 1 2 ICV_23 $T=256680 470560 0 0 $X=256490 $Y=470320
X1766 1 2 ICV_23 $T=256680 486880 0 0 $X=256490 $Y=486640
X1767 1 2 ICV_23 $T=256680 503200 0 0 $X=256490 $Y=502960
X1768 1 2 ICV_23 $T=270940 497760 1 0 $X=270750 $Y=494800
X1769 1 2 ICV_23 $T=270940 503200 1 0 $X=270750 $Y=500240
X1770 1 2 ICV_23 $T=284740 465120 0 0 $X=284550 $Y=464880
X1771 1 2 ICV_23 $T=312800 486880 0 0 $X=312610 $Y=486640
X1772 1 2 ICV_23 $T=340860 486880 0 0 $X=340670 $Y=486640
X1773 1 2 ICV_23 $T=368920 476000 0 0 $X=368730 $Y=475760
X1774 1 2 ICV_23 $T=368920 497760 0 0 $X=368730 $Y=497520
X1775 1 2 ICV_23 $T=368920 503200 0 0 $X=368730 $Y=502960
X1776 1 2 ICV_23 $T=383180 486880 1 0 $X=382990 $Y=483920
X1777 1 2 ICV_23 $T=411240 459680 1 0 $X=411050 $Y=456720
X1778 1 2 ICV_23 $T=495420 470560 1 0 $X=495230 $Y=467600
X1779 1 2 ICV_23 $T=509220 476000 0 0 $X=509030 $Y=475760
X1780 1 2 ICV_23 $T=523480 497760 1 0 $X=523290 $Y=494800
X1781 1 2 ICV_23 $T=551540 508640 1 0 $X=551350 $Y=505680
X1782 1 2 ICV_23 $T=607660 481440 1 0 $X=607470 $Y=478480
X1783 1 2 ICV_23 $T=607660 497760 1 0 $X=607470 $Y=494800
X1784 1 2 ICV_23 $T=621460 497760 0 0 $X=621270 $Y=497520
X1785 1 2 ICV_23 $T=621460 508640 0 0 $X=621270 $Y=508400
X1786 1 2 ICV_23 $T=649520 508640 0 0 $X=649330 $Y=508400
X1787 1 2 ICV_23 $T=663780 459680 1 0 $X=663590 $Y=456720
X1788 1 2 ICV_23 $T=663780 470560 1 0 $X=663590 $Y=467600
X1789 1 2 ICV_23 $T=663780 486880 1 0 $X=663590 $Y=483920
X1790 1 2 ICV_23 $T=691840 486880 1 0 $X=691650 $Y=483920
X1791 1 2 ICV_23 $T=705640 448800 0 0 $X=705450 $Y=448560
X1792 1 2 ICV_23 $T=705640 459680 0 0 $X=705450 $Y=459440
X1793 1 2 ICV_23 $T=705640 486880 0 0 $X=705450 $Y=486640
X1794 1 2 ICV_23 $T=719900 492320 1 0 $X=719710 $Y=489360
X1795 1 2 ICV_24 $T=17940 497760 1 0 $X=17750 $Y=494800
X1796 1 2 ICV_24 $T=17940 508640 1 0 $X=17750 $Y=505680
X1797 1 2 ICV_24 $T=17940 514080 1 0 $X=17750 $Y=511120
X1798 1 2 ICV_24 $T=46000 476000 1 0 $X=45810 $Y=473040
X1799 1 2 ICV_24 $T=87860 465120 0 0 $X=87670 $Y=464880
X1800 1 2 ICV_24 $T=102120 497760 1 0 $X=101930 $Y=494800
X1801 1 2 ICV_24 $T=130180 459680 1 0 $X=129990 $Y=456720
X1802 1 2 ICV_24 $T=143980 459680 0 0 $X=143790 $Y=459440
X1803 1 2 ICV_24 $T=143980 476000 0 0 $X=143790 $Y=475760
X1804 1 2 ICV_24 $T=172040 470560 0 0 $X=171850 $Y=470320
X1805 1 2 ICV_24 $T=186300 508640 1 0 $X=186110 $Y=505680
X1806 1 2 ICV_24 $T=214360 486880 1 0 $X=214170 $Y=483920
X1807 1 2 ICV_24 $T=228160 476000 0 0 $X=227970 $Y=475760
X1808 1 2 ICV_24 $T=242420 470560 1 0 $X=242230 $Y=467600
X1809 1 2 ICV_24 $T=242420 486880 1 0 $X=242230 $Y=483920
X1810 1 2 ICV_24 $T=256220 497760 0 0 $X=256030 $Y=497520
X1811 1 2 ICV_24 $T=298540 470560 1 0 $X=298350 $Y=467600
X1812 1 2 ICV_24 $T=312340 459680 0 0 $X=312150 $Y=459440
X1813 1 2 ICV_24 $T=354660 476000 1 0 $X=354470 $Y=473040
X1814 1 2 ICV_24 $T=360180 514080 1 0 $X=359990 $Y=511120
X1815 1 2 ICV_24 $T=396520 443360 0 0 $X=396330 $Y=443120
X1816 1 2 ICV_24 $T=396520 476000 0 0 $X=396330 $Y=475760
X1817 1 2 ICV_24 $T=396520 492320 0 0 $X=396330 $Y=492080
X1818 1 2 ICV_24 $T=431480 514080 1 0 $X=431290 $Y=511120
X1819 1 2 ICV_24 $T=438840 497760 1 0 $X=438650 $Y=494800
X1820 1 2 ICV_24 $T=494960 492320 1 0 $X=494770 $Y=489360
X1821 1 2 ICV_24 $T=508760 443360 0 0 $X=508570 $Y=443120
X1822 1 2 ICV_24 $T=508760 459680 0 0 $X=508570 $Y=459440
X1823 1 2 ICV_24 $T=508760 470560 0 0 $X=508570 $Y=470320
X1824 1 2 ICV_24 $T=523020 481440 1 0 $X=522830 $Y=478480
X1825 1 2 ICV_24 $T=523020 503200 1 0 $X=522830 $Y=500240
X1826 1 2 ICV_24 $T=564880 476000 0 0 $X=564690 $Y=475760
X1827 1 2 ICV_24 $T=564880 508640 0 0 $X=564690 $Y=508400
X1828 1 2 ICV_24 $T=579140 492320 1 0 $X=578950 $Y=489360
X1829 1 2 ICV_24 $T=592940 448800 0 0 $X=592750 $Y=448560
X1830 1 2 ICV_24 $T=592940 492320 0 0 $X=592750 $Y=492080
X1831 1 2 ICV_24 $T=607200 459680 1 0 $X=607010 $Y=456720
X1832 1 2 ICV_24 $T=621000 465120 0 0 $X=620810 $Y=464880
X1833 1 2 ICV_24 $T=621000 470560 0 0 $X=620810 $Y=470320
X1834 1 2 ICV_24 $T=635260 476000 1 0 $X=635070 $Y=473040
X1835 1 2 ICV_24 $T=635260 486880 1 0 $X=635070 $Y=483920
X1836 1 2 ICV_24 $T=705180 443360 0 0 $X=704990 $Y=443120
X1837 1 2 ICV_24 $T=719440 459680 1 0 $X=719250 $Y=456720
X1838 1 2 ICV_24 $T=719440 508640 1 0 $X=719250 $Y=505680
X1839 1 2 10 2 334 1 sky130_fd_sc_hd__inv_1 $T=18400 470560 1 0 $X=18210 $Y=467600
X1840 1 2 4 2 339 1 sky130_fd_sc_hd__inv_1 $T=24840 454240 0 0 $X=24650 $Y=454000
X1841 1 2 11 2 340 1 sky130_fd_sc_hd__inv_1 $T=27600 486880 1 0 $X=27410 $Y=483920
X1842 1 2 34 2 385 1 sky130_fd_sc_hd__inv_1 $T=41400 454240 0 0 $X=41210 $Y=454000
X1843 1 2 31 2 369 1 sky130_fd_sc_hd__inv_1 $T=44620 476000 1 0 $X=44430 $Y=473040
X1844 1 2 38 2 382 1 sky130_fd_sc_hd__inv_1 $T=50600 492320 0 0 $X=50410 $Y=492080
X1845 1 2 40 2 364 1 sky130_fd_sc_hd__inv_1 $T=59340 465120 0 0 $X=59150 $Y=464880
X1846 1 2 39 2 420 1 sky130_fd_sc_hd__inv_1 $T=60260 470560 0 0 $X=60070 $Y=470320
X1847 1 2 45 2 428 1 sky130_fd_sc_hd__inv_1 $T=70380 492320 0 0 $X=70190 $Y=492080
X1848 1 2 51 2 436 1 sky130_fd_sc_hd__inv_1 $T=80500 465120 1 0 $X=80310 $Y=462160
X1849 1 2 55 2 459 1 sky130_fd_sc_hd__inv_1 $T=88320 486880 1 0 $X=88130 $Y=483920
X1850 1 2 46 2 448 1 sky130_fd_sc_hd__inv_1 $T=89240 448800 1 0 $X=89050 $Y=445840
X1851 1 2 61 2 485 1 sky130_fd_sc_hd__inv_1 $T=98440 454240 1 0 $X=98250 $Y=451280
X1852 1 2 49 2 470 1 sky130_fd_sc_hd__inv_1 $T=98440 470560 1 0 $X=98250 $Y=467600
X1853 1 2 53 2 484 1 sky130_fd_sc_hd__inv_1 $T=104420 481440 1 0 $X=104230 $Y=478480
X1854 1 2 56 2 529 1 sky130_fd_sc_hd__inv_1 $T=122360 470560 0 0 $X=122170 $Y=470320
X1855 1 2 68 2 513 1 sky130_fd_sc_hd__inv_1 $T=124660 454240 0 0 $X=124470 $Y=454000
X1856 1 2 66 2 533 1 sky130_fd_sc_hd__inv_1 $T=129720 486880 0 0 $X=129530 $Y=486640
X1857 1 2 71 2 579 1 sky130_fd_sc_hd__inv_1 $T=143980 486880 1 0 $X=143790 $Y=483920
X1858 1 2 78 2 597 1 sky130_fd_sc_hd__inv_1 $T=154560 481440 0 0 $X=154370 $Y=481200
X1859 1 2 14 2 603 1 sky130_fd_sc_hd__inv_1 $T=160540 443360 0 0 $X=160350 $Y=443120
X1860 1 2 4 2 616 1 sky130_fd_sc_hd__inv_1 $T=168820 459680 1 0 $X=168630 $Y=456720
X1861 1 2 10 2 618 1 sky130_fd_sc_hd__inv_1 $T=168820 476000 1 0 $X=168630 $Y=473040
X1862 1 2 11 2 663 1 sky130_fd_sc_hd__inv_1 $T=181700 476000 0 0 $X=181510 $Y=475760
X1863 1 2 34 2 655 1 sky130_fd_sc_hd__inv_1 $T=186300 454240 1 0 $X=186110 $Y=451280
X1864 1 2 100 2 624 1 sky130_fd_sc_hd__inv_1 $T=186300 492320 1 0 $X=186110 $Y=489360
X1865 1 2 31 2 705 1 sky130_fd_sc_hd__inv_1 $T=200100 470560 0 0 $X=199910 $Y=470320
X1866 1 2 39 2 685 1 sky130_fd_sc_hd__inv_1 $T=204700 465120 1 0 $X=204510 $Y=462160
X1867 1 2 108 2 704 1 sky130_fd_sc_hd__inv_1 $T=213900 448800 1 0 $X=213710 $Y=445840
X1868 1 2 53 2 752 1 sky130_fd_sc_hd__inv_1 $T=225860 454240 1 0 $X=225670 $Y=451280
X1869 1 2 118 2 735 1 sky130_fd_sc_hd__inv_1 $T=226780 476000 0 0 $X=226590 $Y=475760
X1870 1 2 51 2 734 1 sky130_fd_sc_hd__inv_1 $T=229540 465120 1 0 $X=229350 $Y=462160
X1871 1 2 38 2 769 1 sky130_fd_sc_hd__inv_1 $T=232760 476000 0 0 $X=232570 $Y=475760
X1872 1 2 40 2 781 1 sky130_fd_sc_hd__inv_1 $T=240580 465120 1 0 $X=240390 $Y=462160
X1873 1 2 119 2 736 1 sky130_fd_sc_hd__inv_1 $T=242420 497760 1 0 $X=242230 $Y=494800
X1874 1 2 116 2 732 1 sky130_fd_sc_hd__inv_1 $T=248860 486880 0 0 $X=248670 $Y=486640
X1875 1 2 45 2 812 1 sky130_fd_sc_hd__inv_1 $T=255300 486880 0 0 $X=255110 $Y=486640
X1876 1 2 49 2 826 1 sky130_fd_sc_hd__inv_1 $T=269560 465120 0 0 $X=269370 $Y=464880
X1877 1 2 68 2 808 1 sky130_fd_sc_hd__inv_1 $T=270020 448800 0 0 $X=269830 $Y=448560
X1878 1 2 56 2 839 1 sky130_fd_sc_hd__inv_1 $T=279220 476000 1 0 $X=279030 $Y=473040
X1879 1 2 139 2 847 1 sky130_fd_sc_hd__inv_1 $T=286580 443360 0 0 $X=286390 $Y=443120
X1880 1 2 70 2 876 1 sky130_fd_sc_hd__inv_1 $T=309120 470560 0 0 $X=308930 $Y=470320
X1881 1 2 166 2 902 1 sky130_fd_sc_hd__inv_1 $T=338560 486880 1 0 $X=338370 $Y=483920
X1882 1 2 160 2 903 1 sky130_fd_sc_hd__inv_1 $T=340860 492320 0 0 $X=340670 $Y=492080
X1883 1 2 177 2 174 1 sky130_fd_sc_hd__inv_1 $T=353280 443360 0 0 $X=353090 $Y=443120
X1884 1 2 169 2 945 1 sky130_fd_sc_hd__inv_1 $T=354660 448800 0 0 $X=354470 $Y=448560
X1885 1 2 176 2 915 1 sky130_fd_sc_hd__inv_1 $T=355120 481440 1 0 $X=354930 $Y=478480
X1886 1 2 171 2 958 1 sky130_fd_sc_hd__inv_1 $T=356960 465120 1 0 $X=356770 $Y=462160
X1887 1 2 178 2 972 1 sky130_fd_sc_hd__inv_1 $T=367540 497760 0 0 $X=367350 $Y=497520
X1888 1 2 187 2 994 1 sky130_fd_sc_hd__inv_1 $T=376740 492320 1 0 $X=376550 $Y=489360
X1889 1 2 183 2 1014 1 sky130_fd_sc_hd__inv_1 $T=379500 470560 0 0 $X=379310 $Y=470320
X1890 1 2 186 2 1021 1 sky130_fd_sc_hd__inv_1 $T=382720 497760 1 0 $X=382530 $Y=494800
X1891 1 2 193 2 1016 1 sky130_fd_sc_hd__inv_1 $T=391000 476000 1 0 $X=390810 $Y=473040
X1892 1 2 188 2 1051 1 sky130_fd_sc_hd__inv_1 $T=397440 459680 1 0 $X=397250 $Y=456720
X1893 1 2 190 2 1065 1 sky130_fd_sc_hd__inv_1 $T=402040 497760 1 0 $X=401850 $Y=494800
X1894 1 2 185 2 1046 1 sky130_fd_sc_hd__inv_1 $T=402960 448800 1 0 $X=402770 $Y=445840
X1895 1 2 200 2 1080 1 sky130_fd_sc_hd__inv_1 $T=417680 465120 0 0 $X=417490 $Y=464880
X1896 1 2 197 2 1095 1 sky130_fd_sc_hd__inv_1 $T=417680 481440 0 0 $X=417490 $Y=481200
X1897 1 2 206 2 1107 1 sky130_fd_sc_hd__inv_1 $T=425040 454240 0 0 $X=424850 $Y=454000
X1898 1 2 201 2 1129 1 sky130_fd_sc_hd__inv_1 $T=425040 497760 0 0 $X=424850 $Y=497520
X1899 1 2 205 2 1142 1 sky130_fd_sc_hd__inv_1 $T=437000 470560 1 0 $X=436810 $Y=467600
X1900 1 2 209 2 1143 1 sky130_fd_sc_hd__inv_1 $T=441140 486880 1 0 $X=440950 $Y=483920
X1901 1 2 207 2 1138 1 sky130_fd_sc_hd__inv_1 $T=441140 497760 1 0 $X=440950 $Y=494800
X1902 1 2 218 2 210 1 sky130_fd_sc_hd__inv_1 $T=450800 448800 1 0 $X=450610 $Y=445840
X1903 1 2 212 2 1176 1 sky130_fd_sc_hd__inv_1 $T=454940 454240 0 0 $X=454750 $Y=454000
X1904 1 2 213 2 1199 1 sky130_fd_sc_hd__inv_1 $T=460000 470560 1 0 $X=459810 $Y=467600
X1905 1 2 217 2 1205 1 sky130_fd_sc_hd__inv_1 $T=463220 497760 1 0 $X=463030 $Y=494800
X1906 1 2 215 2 1105 1 sky130_fd_sc_hd__inv_1 $T=465060 481440 1 0 $X=464870 $Y=478480
X1907 1 2 223 2 1231 1 sky130_fd_sc_hd__inv_1 $T=476560 497760 1 0 $X=476370 $Y=494800
X1908 1 2 222 2 228 1 sky130_fd_sc_hd__inv_1 $T=479320 459680 1 0 $X=479130 $Y=456720
X1909 1 2 226 2 1230 1 sky130_fd_sc_hd__inv_1 $T=482540 476000 1 0 $X=482350 $Y=473040
X1910 1 2 221 2 1239 1 sky130_fd_sc_hd__inv_1 $T=494500 454240 1 0 $X=494310 $Y=451280
X1911 1 2 236 2 1282 1 sky130_fd_sc_hd__inv_1 $T=495420 465120 1 0 $X=495230 $Y=462160
X1912 1 2 227 2 1216 1 sky130_fd_sc_hd__inv_1 $T=497260 481440 1 0 $X=497070 $Y=478480
X1913 1 2 234 2 1276 1 sky130_fd_sc_hd__inv_1 $T=497260 497760 1 0 $X=497070 $Y=494800
X1914 1 2 247 2 1322 1 sky130_fd_sc_hd__inv_1 $T=509220 497760 0 0 $X=509030 $Y=497520
X1915 1 2 243 2 1304 1 sky130_fd_sc_hd__inv_1 $T=511060 448800 0 0 $X=510870 $Y=448560
X1916 1 2 240 2 1293 1 sky130_fd_sc_hd__inv_1 $T=520260 476000 0 0 $X=520070 $Y=475760
X1917 1 2 251 2 1324 1 sky130_fd_sc_hd__inv_1 $T=521180 459680 1 0 $X=520990 $Y=456720
X1918 1 2 244 2 1325 1 sky130_fd_sc_hd__inv_1 $T=522560 486880 1 0 $X=522370 $Y=483920
X1919 1 2 162 2 1351 1 sky130_fd_sc_hd__inv_1 $T=534060 454240 1 0 $X=533870 $Y=451280
X1920 1 2 193 2 1365 1 sky130_fd_sc_hd__inv_1 $T=534520 470560 1 0 $X=534330 $Y=467600
X1921 1 2 197 2 1371 1 sky130_fd_sc_hd__inv_1 $T=546480 476000 0 0 $X=546290 $Y=475760
X1922 1 2 168 2 1378 1 sky130_fd_sc_hd__inv_1 $T=551080 497760 0 0 $X=550890 $Y=497520
X1923 1 2 160 2 1354 1 sky130_fd_sc_hd__inv_1 $T=553380 492320 1 0 $X=553190 $Y=489360
X1924 1 2 176 2 1409 1 sky130_fd_sc_hd__inv_1 $T=555680 454240 0 0 $X=555490 $Y=454000
X1925 1 2 187 2 1412 1 sky130_fd_sc_hd__inv_1 $T=557060 470560 0 0 $X=556870 $Y=470320
X1926 1 2 186 2 1438 1 sky130_fd_sc_hd__inv_1 $T=571320 497760 1 0 $X=571130 $Y=494800
X1927 1 2 177 2 279 1 sky130_fd_sc_hd__inv_1 $T=574540 443360 0 0 $X=574350 $Y=443120
X1928 1 2 183 2 1456 1 sky130_fd_sc_hd__inv_1 $T=579600 470560 1 0 $X=579410 $Y=467600
X1929 1 2 209 2 1418 1 sky130_fd_sc_hd__inv_1 $T=579600 481440 1 0 $X=579410 $Y=478480
X1930 1 2 166 2 1476 1 sky130_fd_sc_hd__inv_1 $T=587420 486880 0 0 $X=587230 $Y=486640
X1931 1 2 188 2 283 1 sky130_fd_sc_hd__inv_1 $T=591560 448800 0 0 $X=591370 $Y=448560
X1932 1 2 178 2 1495 1 sky130_fd_sc_hd__inv_1 $T=601220 497760 1 0 $X=601030 $Y=494800
X1933 1 2 200 2 1516 1 sky130_fd_sc_hd__inv_1 $T=606740 470560 1 0 $X=606550 $Y=467600
X1934 1 2 201 2 1524 1 sky130_fd_sc_hd__inv_1 $T=609500 492320 0 0 $X=609310 $Y=492080
X1935 1 2 185 2 287 1 sky130_fd_sc_hd__inv_1 $T=615940 448800 1 0 $X=615750 $Y=445840
X1936 1 2 215 2 1544 1 sky130_fd_sc_hd__inv_1 $T=619160 481440 1 0 $X=618970 $Y=478480
X1937 1 2 190 2 1556 1 sky130_fd_sc_hd__inv_1 $T=625600 497760 1 0 $X=625410 $Y=494800
X1938 1 2 205 2 1553 1 sky130_fd_sc_hd__inv_1 $T=630200 465120 1 0 $X=630010 $Y=462160
X1939 1 2 181 2 1575 1 sky130_fd_sc_hd__inv_1 $T=640320 448800 0 0 $X=640130 $Y=448560
X1940 1 2 213 2 1592 1 sky130_fd_sc_hd__inv_1 $T=645380 476000 1 0 $X=645190 $Y=473040
X1941 1 2 217 2 1613 1 sky130_fd_sc_hd__inv_1 $T=655500 497760 1 0 $X=655310 $Y=494800
X1942 1 2 212 2 1619 1 sky130_fd_sc_hd__inv_1 $T=655960 459680 1 0 $X=655770 $Y=456720
X1943 1 2 234 2 1622 1 sky130_fd_sc_hd__inv_1 $T=658260 476000 0 0 $X=658070 $Y=475760
X1944 1 2 207 2 1631 1 sky130_fd_sc_hd__inv_1 $T=663780 492320 1 0 $X=663590 $Y=489360
X1945 1 2 223 2 1658 1 sky130_fd_sc_hd__inv_1 $T=676200 492320 0 0 $X=676010 $Y=492080
X1946 1 2 226 2 1661 1 sky130_fd_sc_hd__inv_1 $T=677580 470560 0 0 $X=677390 $Y=470320
X1947 1 2 227 2 1692 1 sky130_fd_sc_hd__inv_1 $T=693680 481440 1 0 $X=693490 $Y=478480
X1948 1 2 247 2 1705 1 sky130_fd_sc_hd__inv_1 $T=701960 497760 0 0 $X=701770 $Y=497520
X1949 1 2 222 2 308 1 sky130_fd_sc_hd__inv_1 $T=704260 448800 0 0 $X=704070 $Y=448560
X1950 1 2 236 2 1733 1 sky130_fd_sc_hd__inv_1 $T=715300 459680 0 0 $X=715110 $Y=459440
X1951 1 2 244 2 1738 1 sky130_fd_sc_hd__inv_1 $T=715760 481440 0 0 $X=715570 $Y=481200
X1952 1 2 251 2 1744 1 sky130_fd_sc_hd__inv_1 $T=718060 459680 1 0 $X=717870 $Y=456720
X1953 1 2 240 2 1742 1 sky130_fd_sc_hd__inv_1 $T=718980 470560 1 0 $X=718790 $Y=467600
X1954 1 2 ICV_25 $T=30360 508640 0 0 $X=30170 $Y=508400
X1955 1 2 ICV_25 $T=44620 470560 1 0 $X=44430 $Y=467600
X1956 1 2 ICV_25 $T=100740 481440 1 0 $X=100550 $Y=478480
X1957 1 2 ICV_25 $T=114540 497760 0 0 $X=114350 $Y=497520
X1958 1 2 ICV_25 $T=128800 492320 1 0 $X=128610 $Y=489360
X1959 1 2 ICV_25 $T=128800 503200 1 0 $X=128610 $Y=500240
X1960 1 2 ICV_25 $T=156860 465120 1 0 $X=156670 $Y=462160
X1961 1 2 ICV_25 $T=170660 459680 0 0 $X=170470 $Y=459440
X1962 1 2 ICV_25 $T=226780 508640 0 0 $X=226590 $Y=508400
X1963 1 2 ICV_25 $T=297160 503200 1 0 $X=296970 $Y=500240
X1964 1 2 ICV_25 $T=339020 448800 0 0 $X=338830 $Y=448560
X1965 1 2 ICV_25 $T=339020 454240 0 0 $X=338830 $Y=454000
X1966 1 2 ICV_25 $T=353280 486880 1 0 $X=353090 $Y=483920
X1967 1 2 ICV_25 $T=465520 465120 1 0 $X=465330 $Y=462160
X1968 1 2 ICV_25 $T=507380 492320 0 0 $X=507190 $Y=492080
X1969 1 2 ICV_25 $T=521640 465120 1 0 $X=521450 $Y=462160
X1970 1 2 ICV_25 $T=619620 443360 0 0 $X=619430 $Y=443120
X1971 1 2 ICV_25 $T=619620 481440 0 0 $X=619430 $Y=481200
X1972 1 2 ICV_25 $T=703800 476000 0 0 $X=703610 $Y=475760
X1973 1 2 ICV_25 $T=718060 454240 1 0 $X=717870 $Y=451280
X1974 1 2 362 364 21 ICV_26 $T=27600 454240 1 0 $X=27410 $Y=451280
X1975 1 2 368 369 32 ICV_26 $T=28980 486880 0 0 $X=28790 $Y=486640
X1976 1 2 376 382 32 ICV_26 $T=37720 503200 0 0 $X=37530 $Y=502960
X1977 1 2 397 35 27 ICV_26 $T=45540 443360 0 0 $X=45350 $Y=443120
X1978 1 2 401 382 30 ICV_26 $T=48300 492320 1 0 $X=48110 $Y=489360
X1979 1 2 412 364 28 ICV_26 $T=57040 459680 0 0 $X=56850 $Y=459440
X1980 1 2 491 470 28 ICV_26 $T=94300 476000 0 0 $X=94110 $Y=475760
X1981 1 2 520 504 27 ICV_26 $T=109940 497760 0 0 $X=109750 $Y=497520
X1982 1 2 525 504 30 ICV_26 $T=110860 492320 1 0 $X=110670 $Y=489360
X1983 1 2 530 513 28 ICV_26 $T=112700 454240 0 0 $X=112510 $Y=454000
X1984 1 2 527 529 32 ICV_26 $T=112700 476000 0 0 $X=112510 $Y=475760
X1985 1 2 532 533 20 ICV_26 $T=113160 492320 0 0 $X=112970 $Y=492080
X1986 1 2 549 533 21 ICV_26 $T=124200 492320 1 0 $X=124010 $Y=489360
X1987 1 2 566 568 21 ICV_26 $T=132480 459680 1 0 $X=132290 $Y=456720
X1988 1 2 567 561 25 ICV_26 $T=132480 481440 1 0 $X=132290 $Y=478480
X1989 1 2 607 616 93 ICV_26 $T=154560 459680 0 0 $X=154370 $Y=459440
X1990 1 2 610 616 94 ICV_26 $T=155020 470560 1 0 $X=154830 $Y=467600
X1991 1 2 647 616 103 ICV_26 $T=169280 470560 1 0 $X=169090 $Y=467600
X1992 1 2 674 624 25 ICV_26 $T=184460 492320 0 0 $X=184270 $Y=492080
X1993 1 2 692 685 96 ICV_26 $T=194580 459680 0 0 $X=194390 $Y=459440
X1994 1 2 694 705 103 ICV_26 $T=197340 481440 0 0 $X=197150 $Y=481200
X1995 1 2 714 685 92 ICV_26 $T=202400 470560 0 0 $X=202210 $Y=470320
X1996 1 2 733 736 25 ICV_26 $T=211600 497760 1 0 $X=211410 $Y=494800
X1997 1 2 759 735 21 ICV_26 $T=225400 481440 0 0 $X=225210 $Y=481200
X1998 1 2 770 769 94 ICV_26 $T=233220 465120 0 0 $X=233030 $Y=464880
X1999 1 2 793 732 32 ICV_26 $T=244260 486880 0 0 $X=244070 $Y=486640
X2000 1 2 800 133 93 ICV_26 $T=252080 448800 1 0 $X=251890 $Y=445840
X2001 1 2 825 826 101 ICV_26 $T=264960 465120 0 0 $X=264770 $Y=464880
X2002 1 2 830 812 92 ICV_26 $T=266340 481440 0 0 $X=266150 $Y=481200
X2003 1 2 834 808 92 ICV_26 $T=271400 448800 0 0 $X=271210 $Y=448560
X2004 1 2 896 897 151 ICV_26 $T=314640 465120 0 0 $X=314450 $Y=464880
X2005 1 2 944 915 170 ICV_26 $T=337640 476000 0 0 $X=337450 $Y=475760
X2006 1 2 984 972 151 ICV_26 $T=356960 497760 1 0 $X=356770 $Y=494800
X2007 1 2 1030 1021 155 ICV_26 $T=380880 497760 0 0 $X=380690 $Y=497520
X2008 1 2 1036 1021 170 ICV_26 $T=381800 508640 0 0 $X=381610 $Y=508400
X2009 1 2 1042 1046 152 ICV_26 $T=386400 448800 0 0 $X=386210 $Y=448560
X2010 1 2 1075 1051 157 ICV_26 $T=398820 459680 0 0 $X=398630 $Y=459440
X2011 1 2 1127 1129 170 ICV_26 $T=420900 508640 0 0 $X=420710 $Y=508400
X2012 1 2 1144 1138 167 ICV_26 $T=426880 508640 0 0 $X=426690 $Y=508400
X2013 1 2 1147 1107 155 ICV_26 $T=427800 465120 1 0 $X=427610 $Y=462160
X2014 1 2 1195 1199 156 ICV_26 $T=454940 476000 0 0 $X=454750 $Y=475760
X2015 1 2 1200 1205 155 ICV_26 $T=454940 497760 0 0 $X=454750 $Y=497520
X2016 1 2 1203 1205 157 ICV_26 $T=456320 508640 1 0 $X=456130 $Y=505680
X2017 1 2 1281 1282 170 ICV_26 $T=492200 486880 1 0 $X=492010 $Y=483920
X2018 1 2 1294 1293 151 ICV_26 $T=497260 476000 1 0 $X=497070 $Y=473040
X2019 1 2 1302 1304 151 ICV_26 $T=505080 448800 0 0 $X=504890 $Y=448560
X2020 1 2 1318 250 151 ICV_26 $T=507840 448800 1 0 $X=507650 $Y=445840
X2021 1 2 1349 1351 255 ICV_26 $T=523940 448800 0 0 $X=523750 $Y=448560
X2022 1 2 1413 1412 266 ICV_26 $T=556140 476000 1 0 $X=555950 $Y=473040
X2023 1 2 1441 279 275 ICV_26 $T=571320 454240 0 0 $X=571130 $Y=454000
X2024 1 2 1455 1438 275 ICV_26 $T=578680 492320 0 0 $X=578490 $Y=492080
X2025 1 2 1453 1459 270 ICV_26 $T=579600 465120 0 0 $X=579410 $Y=464880
X2026 1 2 1494 1495 266 ICV_26 $T=596620 497760 1 0 $X=596430 $Y=494800
X2027 1 2 1511 1516 255 ICV_26 $T=606280 465120 0 0 $X=606090 $Y=464880
X2028 1 2 1530 1524 255 ICV_26 $T=614100 514080 1 0 $X=613910 $Y=511120
X2029 1 2 1534 1524 270 ICV_26 $T=616860 508640 0 0 $X=616670 $Y=508400
X2030 1 2 1551 287 255 ICV_26 $T=621460 448800 1 0 $X=621270 $Y=445840
X2031 1 2 1546 1553 268 ICV_26 $T=621460 470560 1 0 $X=621270 $Y=467600
X2032 1 2 1554 1553 262 ICV_26 $T=625600 465120 1 0 $X=625410 $Y=462160
X2033 1 2 1585 1563 264 ICV_26 $T=640320 465120 1 0 $X=640130 $Y=462160
X2034 1 2 1595 1592 255 ICV_26 $T=645380 470560 0 0 $X=645190 $Y=470320
X2035 1 2 1610 1563 266 ICV_26 $T=650440 459680 1 0 $X=650250 $Y=456720
X2036 1 2 1606 1613 264 ICV_26 $T=650900 497760 1 0 $X=650710 $Y=494800
X2037 1 2 1603 1575 269 ICV_26 $T=651360 443360 0 0 $X=651170 $Y=443120
X2038 1 2 1612 1613 266 ICV_26 $T=651360 492320 0 0 $X=651170 $Y=492080
X2039 1 2 1642 1631 266 ICV_26 $T=665620 492320 1 0 $X=665430 $Y=489360
X2040 1 2 1697 1679 270 ICV_26 $T=698740 465120 0 0 $X=698550 $Y=464880
X2041 1 2 1704 1705 270 ICV_26 $T=699660 508640 0 0 $X=699470 $Y=508400
X2042 1 2 1746 1744 268 ICV_26 $T=716680 459680 0 0 $X=716490 $Y=459440
X2043 1 2 487 13 524 62 504 ICV_27 $T=104420 492320 0 0 $X=104230 $Y=492080
X2044 1 2 559 15 586 74 568 ICV_27 $T=136160 448800 0 0 $X=135970 $Y=448560
X2045 1 2 547 19 585 70 561 ICV_27 $T=136620 470560 1 0 $X=136430 $Y=467600
X2046 1 2 636 26 654 88 630 ICV_27 $T=167900 492320 1 0 $X=167710 $Y=489360
X2047 1 2 665 26 706 110 689 ICV_27 $T=191820 492320 1 0 $X=191630 $Y=489360
X2048 1 2 786 83 818 130 133 ICV_27 $T=256680 448800 1 0 $X=256490 $Y=445840
X2049 1 2 851 98 868 138 864 ICV_27 $T=289340 459680 1 0 $X=289150 $Y=456720
X2050 1 2 878 95 887 61 890 ICV_27 $T=304980 448800 0 0 $X=304790 $Y=448560
X2051 1 2 895 161 936 162 897 ICV_27 $T=329360 465120 0 0 $X=329170 $Y=464880
X2052 1 2 904 165 959 168 925 ICV_27 $T=341320 503200 1 0 $X=341130 $Y=500240
X2053 1 2 988 149 1022 181 1000 ICV_27 $T=368000 454240 1 0 $X=367810 $Y=451280
X2054 1 2 1443 267 1468 171 1459 ICV_27 $T=576840 459680 0 0 $X=576650 $Y=459440
X2055 1 2 1576 267 1561 206 1563 ICV_27 $T=633880 454240 0 0 $X=633690 $Y=454000
X2056 1 2 300 256 1666 218 301 ICV_27 $T=672520 448800 1 0 $X=672330 $Y=445840
X2057 1 2 1668 259 1687 221 1679 ICV_27 $T=684480 459680 1 0 $X=684290 $Y=456720
X2058 1 2 313 257 1743 243 317 ICV_27 $T=710240 448800 1 0 $X=710050 $Y=445840
X2059 1 2 325 9 335 ICV_28 $T=6900 470560 1 0 $X=6710 $Y=467600
X2060 1 2 33 26 374 ICV_28 $T=28520 448800 1 0 $X=28330 $Y=445840
X2061 1 2 33 15 397 ICV_28 $T=37720 448800 1 0 $X=37530 $Y=445840
X2062 1 2 371 15 402 ICV_28 $T=41400 492320 0 0 $X=41210 $Y=492080
X2063 1 2 407 7 423 ICV_28 $T=51980 492320 0 0 $X=51790 $Y=492080
X2064 1 2 445 15 476 ICV_28 $T=78660 497760 0 0 $X=78470 $Y=497520
X2065 1 2 58 15 507 ICV_28 $T=94300 448800 0 0 $X=94110 $Y=448560
X2066 1 2 464 19 508 ICV_28 $T=94300 459680 0 0 $X=94110 $Y=459440
X2067 1 2 511 8 512 ICV_28 $T=104420 470560 1 0 $X=104230 $Y=467600
X2068 1 2 593 85 610 ICV_28 $T=146280 465120 0 0 $X=146090 $Y=464880
X2069 1 2 649 98 653 ICV_28 $T=170200 459680 1 0 $X=170010 $Y=456720
X2070 1 2 675 82 684 ICV_28 $T=185380 459680 0 0 $X=185190 $Y=459440
X2071 1 2 720 13 733 ICV_28 $T=206540 497760 0 0 $X=206350 $Y=497520
X2072 1 2 746 95 755 ICV_28 $T=216660 454240 1 0 $X=216470 $Y=451280
X2073 1 2 813 99 807 ICV_28 $T=256220 459680 1 0 $X=256030 $Y=456720
X2074 1 2 833 99 846 ICV_28 $T=272780 454240 1 0 $X=272590 $Y=451280
X2075 1 2 833 97 867 ICV_28 $T=286580 454240 0 0 $X=286390 $Y=454000
X2076 1 2 898 154 983 ICV_28 $T=350060 481440 0 0 $X=349870 $Y=481200
X2077 1 2 1179 149 1190 ICV_28 $T=442520 465120 0 0 $X=442330 $Y=464880
X2078 1 2 1180 144 1131 ICV_28 $T=442520 486880 1 0 $X=442330 $Y=483920
X2079 1 2 1298 161 1308 ICV_28 $T=498640 481440 1 0 $X=498450 $Y=478480
X2080 1 2 245 150 1337 ICV_28 $T=511060 443360 0 0 $X=510870 $Y=443120
X2081 1 2 1298 144 1339 ICV_28 $T=511060 476000 0 0 $X=510870 $Y=475760
X2082 1 2 1355 257 1364 ICV_28 $T=525320 470560 1 0 $X=525130 $Y=467600
X2083 1 2 1375 257 1381 ICV_28 $T=534520 503200 1 0 $X=534330 $Y=500240
X2084 1 2 1358 261 1399 ICV_28 $T=543260 492320 0 0 $X=543070 $Y=492080
X2085 1 2 1386 259 1406 ICV_28 $T=546480 454240 0 0 $X=546290 $Y=454000
X2086 1 2 1525 267 1562 ICV_28 $T=620540 481440 1 0 $X=620350 $Y=478480
X2087 1 2 1527 259 1570 ICV_28 $T=623300 459680 0 0 $X=623110 $Y=459440
X2088 1 2 293 267 1573 ICV_28 $T=630660 448800 0 0 $X=630470 $Y=448560
X2089 1 2 1588 257 1606 ICV_28 $T=641700 497760 1 0 $X=641510 $Y=494800
X2090 1 2 1618 258 1650 ICV_28 $T=665620 470560 1 0 $X=665430 $Y=467600
X2091 1 2 1618 265 1655 ICV_28 $T=666540 459680 0 0 $X=666350 $Y=459440
X2092 1 2 300 267 306 ICV_28 $T=669760 443360 0 0 $X=669570 $Y=443120
X2093 1 2 1649 256 1665 ICV_28 $T=669760 497760 0 0 $X=669570 $Y=497520
X2094 1 2 1672 267 312 ICV_28 $T=693680 448800 1 0 $X=693490 $Y=445840
X2095 1 2 1721 261 1746 ICV_28 $T=708860 459680 1 0 $X=708670 $Y=456720
X2096 1 2 325 7 336 ICV_29 $T=6900 459680 0 0 $X=6710 $Y=459440
X2097 1 2 404 13 410 ICV_29 $T=48300 476000 0 0 $X=48110 $Y=475760
X2098 1 2 429 8 441 ICV_29 $T=62100 465120 0 0 $X=61910 $Y=464880
X2099 1 2 547 9 564 ICV_29 $T=122360 476000 1 0 $X=122170 $Y=473040
X2100 1 2 619 9 626 ICV_29 $T=153640 503200 0 0 $X=153450 $Y=502960
X2101 1 2 635 83 656 ICV_29 $T=167900 481440 1 0 $X=167710 $Y=478480
X2102 1 2 636 15 657 ICV_29 $T=168820 503200 1 0 $X=168630 $Y=500240
X2103 1 2 636 7 677 ICV_29 $T=176640 492320 1 0 $X=176450 $Y=489360
X2104 1 2 649 83 678 ICV_29 $T=177560 448800 1 0 $X=177370 $Y=445840
X2105 1 2 665 8 681 ICV_29 $T=178480 503200 1 0 $X=178290 $Y=500240
X2106 1 2 720 19 744 ICV_29 $T=206540 503200 1 0 $X=206350 $Y=500240
X2107 1 2 746 86 773 ICV_29 $T=227240 448800 1 0 $X=227050 $Y=445840
X2108 1 2 768 86 779 ICV_29 $T=230920 465120 1 0 $X=230730 $Y=462160
X2109 1 2 786 95 806 ICV_29 $T=244720 454240 1 0 $X=244530 $Y=451280
X2110 1 2 833 86 858 ICV_29 $T=281520 448800 1 0 $X=281330 $Y=445840
X2111 1 2 855 83 874 ICV_29 $T=293940 481440 0 0 $X=293750 $Y=481200
X2112 1 2 898 146 909 ICV_29 $T=314640 481440 0 0 $X=314450 $Y=481200
X2113 1 2 926 149 941 ICV_29 $T=329360 448800 0 0 $X=329170 $Y=448560
X2114 1 2 943 154 954 ICV_29 $T=337180 470560 1 0 $X=336990 $Y=467600
X2115 1 2 943 165 977 ICV_29 $T=346840 470560 1 0 $X=346650 $Y=467600
X2116 1 2 1034 154 1069 ICV_29 $T=388700 459680 0 0 $X=388510 $Y=459440
X2117 1 2 1056 165 1063 ICV_29 $T=388700 503200 0 0 $X=388510 $Y=502960
X2118 1 2 1086 159 1116 ICV_29 $T=409400 514080 1 0 $X=409210 $Y=511120
X2119 1 2 1179 159 1188 ICV_29 $T=441140 476000 1 0 $X=440950 $Y=473040
X2120 1 2 1184 161 1194 ICV_29 $T=443900 508640 0 0 $X=443710 $Y=508400
X2121 1 2 1225 150 1238 ICV_29 $T=462300 503200 0 0 $X=462110 $Y=502960
X2122 1 2 1232 150 1240 ICV_29 $T=463680 481440 0 0 $X=463490 $Y=481200
X2123 1 2 1265 150 1280 ICV_29 $T=483920 476000 1 0 $X=483730 $Y=473040
X2124 1 2 1297 165 1311 ICV_29 $T=498180 503200 0 0 $X=497990 $Y=502960
X2125 1 2 1299 149 1344 ICV_29 $T=511980 465120 1 0 $X=511790 $Y=462160
X2126 1 2 1375 265 1383 ICV_29 $T=534520 508640 1 0 $X=534330 $Y=505680
X2127 1 2 1375 259 1395 ICV_29 $T=539120 497760 0 0 $X=538930 $Y=497520
X2128 1 2 1397 259 1413 ICV_29 $T=547860 476000 0 0 $X=547670 $Y=475760
X2129 1 2 1411 261 1417 ICV_29 $T=554760 492320 1 0 $X=554570 $Y=489360
X2130 1 2 1443 263 1452 ICV_29 $T=569940 465120 1 0 $X=569750 $Y=462160
X2131 1 2 1463 265 1480 ICV_29 $T=583740 486880 1 0 $X=583550 $Y=483920
X2132 1 2 1523 263 288 ICV_29 $T=607660 454240 0 0 $X=607470 $Y=454000
X2133 1 2 1615 257 1626 ICV_29 $T=651360 481440 0 0 $X=651170 $Y=481200
X2134 1 2 1672 257 1686 ICV_29 $T=681260 448800 1 0 $X=681070 $Y=445840
X2135 1 2 1668 257 1694 ICV_29 $T=686780 470560 0 0 $X=686590 $Y=470320
X2136 1 2 1721 257 1745 ICV_29 $T=708400 454240 1 0 $X=708210 $Y=451280
X2137 1 2 341 340 22 346 340 27 ICV_30 $T=16100 492320 0 0 $X=15910 $Y=492080
X2138 1 2 345 334 27 348 334 25 ICV_30 $T=18400 476000 0 0 $X=18210 $Y=475760
X2139 1 2 338 18 25 352 18 30 ICV_30 $T=20240 448800 1 0 $X=20050 $Y=445840
X2140 1 2 343 339 25 335 339 22 ICV_30 $T=20240 465120 1 0 $X=20050 $Y=462160
X2141 1 2 372 369 22 380 382 25 ICV_30 $T=34960 486880 0 0 $X=34770 $Y=486640
X2142 1 2 375 369 27 390 369 20 ICV_30 $T=37260 470560 0 0 $X=37070 $Y=470320
X2143 1 2 421 428 27 423 428 21 ICV_30 $T=62100 492320 0 0 $X=61910 $Y=492080
X2144 1 2 416 420 32 414 420 20 ICV_30 $T=63020 486880 1 0 $X=62830 $Y=483920
X2145 1 2 462 448 28 426 364 30 ICV_30 $T=80960 454240 0 0 $X=80770 $Y=454000
X2146 1 2 469 470 32 475 470 21 ICV_30 $T=83260 465120 1 0 $X=83070 $Y=462160
X2147 1 2 480 484 32 490 484 21 ICV_30 $T=89700 486880 1 0 $X=89510 $Y=483920
X2148 1 2 512 513 20 522 513 32 ICV_30 $T=106720 465120 1 0 $X=106530 $Y=462160
X2149 1 2 538 529 27 541 529 30 ICV_30 $T=118220 476000 0 0 $X=118030 $Y=475760
X2150 1 2 528 529 28 542 529 21 ICV_30 $T=118220 481440 0 0 $X=118030 $Y=481200
X2151 1 2 543 513 30 554 513 21 ICV_30 $T=122820 465120 1 0 $X=122630 $Y=462160
X2152 1 2 556 72 20 562 72 32 ICV_30 $T=126040 454240 0 0 $X=125850 $Y=454000
X2153 1 2 560 561 20 564 561 22 ICV_30 $T=128800 481440 0 0 $X=128610 $Y=481200
X2154 1 2 587 561 27 590 561 32 ICV_30 $T=146280 481440 0 0 $X=146090 $Y=481200
X2155 1 2 602 603 89 614 603 94 ICV_30 $T=151340 454240 1 0 $X=151150 $Y=451280
X2156 1 2 617 618 94 608 618 93 ICV_30 $T=155940 476000 0 0 $X=155750 $Y=475760
X2157 1 2 622 618 96 631 618 102 ICV_30 $T=160540 476000 1 0 $X=160350 $Y=473040
X2158 1 2 628 603 101 642 603 92 ICV_30 $T=163300 448800 0 0 $X=163110 $Y=448560
X2159 1 2 651 630 28 658 624 28 ICV_30 $T=174340 503200 0 0 $X=174150 $Y=502960
X2160 1 2 660 663 93 662 655 101 ICV_30 $T=178940 470560 1 0 $X=178750 $Y=467600
X2161 1 2 670 663 89 677 624 21 ICV_30 $T=181240 486880 0 0 $X=181050 $Y=486640
X2162 1 2 684 685 93 691 685 102 ICV_30 $T=188600 465120 1 0 $X=188410 $Y=462160
X2163 1 2 688 689 32 681 689 20 ICV_30 $T=190900 508640 0 0 $X=190710 $Y=508400
X2164 1 2 695 705 96 698 705 102 ICV_30 $T=197800 476000 1 0 $X=197610 $Y=473040
X2165 1 2 693 685 94 717 685 101 ICV_30 $T=202400 465120 0 0 $X=202210 $Y=464880
X2166 1 2 710 685 89 741 734 92 ICV_30 $T=210680 465120 0 0 $X=210490 $Y=464880
X2167 1 2 796 781 93 801 781 102 ICV_30 $T=247480 465120 0 0 $X=247290 $Y=464880
X2168 1 2 810 812 102 815 812 94 ICV_30 $T=254840 476000 1 0 $X=254650 $Y=473040
X2169 1 2 778 781 89 818 133 92 ICV_30 $T=258520 443360 0 0 $X=258330 $Y=443120
X2170 1 2 820 812 93 804 781 103 ICV_30 $T=264040 476000 1 0 $X=263850 $Y=473040
X2171 1 2 861 826 93 869 876 89 ICV_30 $T=298540 470560 0 0 $X=298350 $Y=470320
X2172 1 2 916 897 157 928 897 152 ICV_30 $T=328900 470560 1 0 $X=328710 $Y=467600
X2173 1 2 924 915 164 934 897 167 ICV_30 $T=329360 476000 0 0 $X=329170 $Y=475760
X2174 1 2 932 902 156 919 903 155 ICV_30 $T=332580 492320 1 0 $X=332390 $Y=489360
X2175 1 2 933 925 156 921 925 152 ICV_30 $T=333040 503200 0 0 $X=332850 $Y=502960
X2176 1 2 952 174 151 917 174 152 ICV_30 $T=342700 443360 0 0 $X=342510 $Y=443120
X2177 1 2 942 945 151 956 958 167 ICV_30 $T=342700 459680 0 0 $X=342510 $Y=459440
X2178 1 2 950 925 151 959 925 164 ICV_30 $T=342700 503200 0 0 $X=342510 $Y=502960
X2179 1 2 955 903 167 960 903 164 ICV_30 $T=345920 492320 1 0 $X=345730 $Y=489360
X2180 1 2 954 958 156 964 958 152 ICV_30 $T=346380 476000 1 0 $X=346190 $Y=473040
X2181 1 2 995 972 170 1007 972 156 ICV_30 $T=363860 514080 1 0 $X=363670 $Y=511120
X2182 1 2 1002 1000 156 1022 1000 155 ICV_30 $T=370760 454240 0 0 $X=370570 $Y=454000
X2183 1 2 1004 1014 156 1010 1014 152 ICV_30 $T=370760 470560 0 0 $X=370570 $Y=470320
X2184 1 2 1013 1016 170 1011 1016 167 ICV_30 $T=371680 481440 0 0 $X=371490 $Y=481200
X2185 1 2 1031 1021 151 1037 1021 152 ICV_30 $T=385020 503200 1 0 $X=384830 $Y=500240
X2186 1 2 1033 1021 157 1044 1021 156 ICV_30 $T=385020 508640 1 0 $X=384830 $Y=505680
X2187 1 2 1050 1051 164 1043 1046 167 ICV_30 $T=388240 454240 0 0 $X=388050 $Y=454000
X2188 1 2 1054 1016 156 1060 994 164 ICV_30 $T=389620 481440 0 0 $X=389430 $Y=481200
X2189 1 2 1068 1046 156 199 196 170 ICV_30 $T=398820 443360 0 0 $X=398630 $Y=443120
X2190 1 2 1079 1080 170 1093 1095 164 ICV_30 $T=402040 481440 1 0 $X=401850 $Y=478480
X2191 1 2 1070 1051 167 1096 1080 152 ICV_30 $T=409400 465120 0 0 $X=409210 $Y=464880
X2192 1 2 1104 1105 170 1110 1095 156 ICV_30 $T=411700 486880 0 0 $X=411510 $Y=486640
X2193 1 2 1099 1107 156 1106 204 152 ICV_30 $T=413080 454240 1 0 $X=412890 $Y=451280
X2194 1 2 1098 1107 157 1102 1107 164 ICV_30 $T=413080 459680 1 0 $X=412890 $Y=456720
X2195 1 2 1185 210 170 1197 1176 151 ICV_30 $T=454940 448800 0 0 $X=454750 $Y=448560
X2196 1 2 1191 1199 151 1218 1199 152 ICV_30 $T=457240 465120 1 0 $X=457050 $Y=462160
X2197 1 2 1202 1205 152 1219 1205 164 ICV_30 $T=460000 503200 1 0 $X=459810 $Y=500240
X2198 1 2 1237 1239 155 1249 1239 151 ICV_30 $T=471040 454240 1 0 $X=470850 $Y=451280
X2199 1 2 1240 1230 157 1244 1230 170 ICV_30 $T=472880 486880 1 0 $X=472690 $Y=483920
X2200 1 2 1275 1276 170 1289 1276 167 ICV_30 $T=492200 514080 1 0 $X=492010 $Y=511120
X2201 1 2 1283 1282 151 1284 1282 167 ICV_30 $T=497260 465120 1 0 $X=497070 $Y=462160
X2202 1 2 1308 1293 170 1315 1293 167 ICV_30 $T=507380 486880 1 0 $X=507190 $Y=483920
X2203 1 2 1306 1322 170 1312 1322 167 ICV_30 $T=510140 514080 1 0 $X=509950 $Y=511120
X2204 1 2 1314 1324 167 1321 1324 164 ICV_30 $T=511060 470560 0 0 $X=510870 $Y=470320
X2205 1 2 1317 1322 151 1305 1325 170 ICV_30 $T=511060 497760 0 0 $X=510870 $Y=497520
X2206 1 2 1341 1304 155 1319 1304 164 ICV_30 $T=525320 459680 1 0 $X=525130 $Y=456720
X2207 1 2 1342 1324 152 1235 228 170 ICV_30 $T=525320 465120 0 0 $X=525130 $Y=464880
X2208 1 2 1339 1293 152 1316 1325 164 ICV_30 $T=525320 476000 1 0 $X=525130 $Y=473040
X2209 1 2 1369 1371 264 1370 1371 255 ICV_30 $T=534980 476000 1 0 $X=534790 $Y=473040
X2210 1 2 1377 1378 269 1383 1378 270 ICV_30 $T=540500 508640 0 0 $X=540310 $Y=508400
X2211 1 2 1379 1351 270 272 273 269 ICV_30 $T=542800 443360 0 0 $X=542610 $Y=443120
X2212 1 2 1398 273 262 1408 273 266 ICV_30 $T=551080 443360 0 0 $X=550890 $Y=443120
X2213 1 2 1388 1351 269 1389 1351 275 ICV_30 $T=553380 454240 1 0 $X=553190 $Y=451280
X2214 1 2 1405 1354 270 1399 1354 268 ICV_30 $T=553380 492320 0 0 $X=553190 $Y=492080
X2215 1 2 1417 1418 268 1425 1418 264 ICV_30 $T=558900 486880 1 0 $X=558710 $Y=483920
X2216 1 2 1419 1412 269 1435 1412 275 ICV_30 $T=567180 476000 0 0 $X=566990 $Y=475760
X2217 1 2 1430 1418 266 1439 1418 262 ICV_30 $T=567180 481440 0 0 $X=566990 $Y=481200
X2218 1 2 1436 1438 264 1447 1418 275 ICV_30 $T=570400 492320 0 0 $X=570210 $Y=492080
X2219 1 2 1467 279 262 1475 279 264 ICV_30 $T=583280 448800 0 0 $X=583090 $Y=448560
X2220 1 2 1484 1456 268 1498 1476 262 ICV_30 $T=595240 481440 0 0 $X=595050 $Y=481200
X2221 1 2 1481 1495 262 1491 1495 269 ICV_30 $T=596160 503200 0 0 $X=595970 $Y=502960
X2222 1 2 1538 1524 275 1540 1544 264 ICV_30 $T=617320 492320 1 0 $X=617130 $Y=489360
X2223 1 2 1548 1553 264 1559 1553 269 ICV_30 $T=623300 470560 0 0 $X=623110 $Y=470320
X2224 1 2 1549 1544 266 1542 1544 268 ICV_30 $T=623300 481440 0 0 $X=623110 $Y=481200
X2225 1 2 1589 1575 262 1593 1575 264 ICV_30 $T=642620 448800 0 0 $X=642430 $Y=448560
X2226 1 2 1591 1592 270 1599 1592 269 ICV_30 $T=644000 481440 1 0 $X=643810 $Y=478480
X2227 1 2 1627 1622 262 1625 1622 255 ICV_30 $T=665620 481440 1 0 $X=665430 $Y=478480
X2228 1 2 1644 1631 270 1638 1631 255 ICV_30 $T=667000 508640 1 0 $X=666810 $Y=505680
X2229 1 2 1646 1622 270 1641 1631 275 ICV_30 $T=667920 486880 1 0 $X=667730 $Y=483920
X2230 1 2 1647 301 266 305 301 269 ICV_30 $T=669300 448800 0 0 $X=669110 $Y=448560
X2231 1 2 1650 1619 255 1655 1619 270 ICV_30 $T=670680 465120 1 0 $X=670490 $Y=462160
X2232 1 2 1657 1619 264 1670 1661 269 ICV_30 $T=676200 470560 1 0 $X=676010 $Y=467600
X2233 1 2 1665 1658 262 1674 1658 269 ICV_30 $T=678960 497760 1 0 $X=678770 $Y=494800
X2234 1 2 1675 1661 266 1684 1661 275 ICV_30 $T=684480 470560 1 0 $X=684290 $Y=467600
X2235 1 2 1676 308 268 1686 308 264 ICV_30 $T=685860 448800 0 0 $X=685670 $Y=448560
X2236 1 2 1683 1679 269 1696 1679 255 ICV_30 $T=693680 465120 1 0 $X=693490 $Y=462160
X2237 1 2 1688 1658 266 1698 1692 275 ICV_30 $T=693680 492320 1 0 $X=693490 $Y=489360
X2238 1 2 1699 1679 275 1708 308 255 ICV_30 $T=698740 454240 0 0 $X=698550 $Y=454000
X2239 1 2 1695 1692 268 1714 1692 269 ICV_30 $T=707480 481440 0 0 $X=707290 $Y=481200
X2240 1 2 4 6 2 324 1 sky130_fd_sc_hd__and2_1 $T=6900 454240 0 0 $X=6710 $Y=454000
X2241 1 2 10 6 2 326 1 sky130_fd_sc_hd__and2_1 $T=8740 476000 1 0 $X=8550 $Y=473040
X2242 1 2 11 6 2 327 1 sky130_fd_sc_hd__and2_1 $T=8740 486880 1 0 $X=8550 $Y=483920
X2243 1 2 14 6 2 16 1 sky130_fd_sc_hd__and2_1 $T=11500 443360 0 0 $X=11310 $Y=443120
X2244 1 2 31 6 2 367 1 sky130_fd_sc_hd__and2_1 $T=27600 476000 1 0 $X=27410 $Y=473040
X2245 1 2 34 6 2 365 1 sky130_fd_sc_hd__and2_1 $T=30360 448800 0 0 $X=30170 $Y=448560
X2246 1 2 38 6 2 391 1 sky130_fd_sc_hd__and2_1 $T=48300 486880 1 0 $X=48110 $Y=483920
X2247 1 2 39 6 2 403 1 sky130_fd_sc_hd__and2_1 $T=48760 470560 1 0 $X=48570 $Y=467600
X2248 1 2 40 6 2 405 1 sky130_fd_sc_hd__and2_1 $T=49680 454240 1 0 $X=49490 $Y=451280
X2249 1 2 45 6 2 430 1 sky130_fd_sc_hd__and2_1 $T=62560 486880 0 0 $X=62370 $Y=486640
X2250 1 2 46 6 2 431 1 sky130_fd_sc_hd__and2_1 $T=63480 448800 0 0 $X=63290 $Y=448560
X2251 1 2 49 6 2 452 1 sky130_fd_sc_hd__and2_1 $T=71760 465120 0 0 $X=71570 $Y=464880
X2252 1 2 51 6 2 442 1 sky130_fd_sc_hd__and2_1 $T=75900 470560 0 0 $X=75710 $Y=470320
X2253 1 2 53 6 2 471 1 sky130_fd_sc_hd__and2_1 $T=83720 481440 1 0 $X=83530 $Y=478480
X2254 1 2 55 6 2 463 1 sky130_fd_sc_hd__and2_1 $T=86020 486880 1 0 $X=85830 $Y=483920
X2255 1 2 56 6 2 479 1 sky130_fd_sc_hd__and2_1 $T=87400 470560 0 0 $X=87210 $Y=470320
X2256 1 2 61 6 2 488 1 sky130_fd_sc_hd__and2_1 $T=100280 448800 1 0 $X=100090 $Y=445840
X2257 1 2 62 6 2 510 1 sky130_fd_sc_hd__and2_1 $T=102120 492320 0 0 $X=101930 $Y=492080
X2258 1 2 66 6 2 531 1 sky130_fd_sc_hd__and2_1 $T=113620 481440 1 0 $X=113430 $Y=478480
X2259 1 2 68 6 2 537 1 sky130_fd_sc_hd__and2_1 $T=115460 459680 1 0 $X=115270 $Y=456720
X2260 1 2 70 6 2 555 1 sky130_fd_sc_hd__and2_1 $T=125580 465120 0 0 $X=125390 $Y=464880
X2261 1 2 71 6 2 558 1 sky130_fd_sc_hd__and2_1 $T=126500 481440 0 0 $X=126310 $Y=481200
X2262 1 2 74 6 2 557 1 sky130_fd_sc_hd__and2_1 $T=133860 448800 0 0 $X=133670 $Y=448560
X2263 1 2 78 6 2 582 1 sky130_fd_sc_hd__and2_1 $T=143060 481440 0 0 $X=142870 $Y=481200
X2264 1 2 10 79 2 591 1 sky130_fd_sc_hd__and2_1 $T=145360 470560 1 0 $X=145170 $Y=467600
X2265 1 2 14 79 2 80 1 sky130_fd_sc_hd__and2_1 $T=146740 443360 0 0 $X=146550 $Y=443120
X2266 1 2 88 6 2 612 1 sky130_fd_sc_hd__and2_1 $T=153640 492320 0 0 $X=153450 $Y=492080
X2267 1 2 4 79 2 595 1 sky130_fd_sc_hd__and2_1 $T=156400 459680 1 0 $X=156210 $Y=456720
X2268 1 2 100 6 2 629 1 sky130_fd_sc_hd__and2_1 $T=163300 492320 0 0 $X=163110 $Y=492080
X2269 1 2 11 79 2 634 1 sky130_fd_sc_hd__and2_1 $T=164220 476000 0 0 $X=164030 $Y=475760
X2270 1 2 34 79 2 650 1 sky130_fd_sc_hd__and2_1 $T=171580 448800 0 0 $X=171390 $Y=448560
X2271 1 2 39 79 2 667 1 sky130_fd_sc_hd__and2_1 $T=180320 465120 1 0 $X=180130 $Y=462160
X2272 1 2 108 6 2 679 1 sky130_fd_sc_hd__and2_1 $T=185380 443360 0 0 $X=185190 $Y=443120
X2273 1 2 31 79 2 676 1 sky130_fd_sc_hd__and2_1 $T=185840 470560 0 0 $X=185650 $Y=470320
X2274 1 2 110 6 2 687 1 sky130_fd_sc_hd__and2_1 $T=189520 492320 1 0 $X=189330 $Y=489360
X2275 1 2 116 6 2 716 1 sky130_fd_sc_hd__and2_1 $T=203320 486880 1 0 $X=203130 $Y=483920
X2276 1 2 118 6 2 721 1 sky130_fd_sc_hd__and2_1 $T=206080 476000 1 0 $X=205890 $Y=473040
X2277 1 2 119 6 2 713 1 sky130_fd_sc_hd__and2_1 $T=208840 486880 0 0 $X=208650 $Y=486640
X2278 1 2 51 79 2 724 1 sky130_fd_sc_hd__and2_1 $T=214820 459680 0 0 $X=214630 $Y=459440
X2279 1 2 53 79 2 737 1 sky130_fd_sc_hd__and2_1 $T=216660 448800 0 0 $X=216470 $Y=448560
X2280 1 2 40 79 2 765 1 sky130_fd_sc_hd__and2_1 $T=230460 459680 0 0 $X=230270 $Y=459440
X2281 1 2 38 79 2 766 1 sky130_fd_sc_hd__and2_1 $T=230460 476000 0 0 $X=230270 $Y=475760
X2282 1 2 130 79 2 777 1 sky130_fd_sc_hd__and2_1 $T=240580 454240 1 0 $X=240390 $Y=451280
X2283 1 2 45 79 2 795 1 sky130_fd_sc_hd__and2_1 $T=245640 476000 0 0 $X=245450 $Y=475760
X2284 1 2 68 79 2 805 1 sky130_fd_sc_hd__and2_1 $T=254380 454240 1 0 $X=254190 $Y=451280
X2285 1 2 49 79 2 814 1 sky130_fd_sc_hd__and2_1 $T=255760 465120 0 0 $X=255570 $Y=464880
X2286 1 2 56 79 2 832 1 sky130_fd_sc_hd__and2_1 $T=269560 470560 1 0 $X=269370 $Y=467600
X2287 1 2 138 79 2 848 1 sky130_fd_sc_hd__and2_1 $T=280600 459680 1 0 $X=280410 $Y=456720
X2288 1 2 61 79 2 871 1 sky130_fd_sc_hd__and2_1 $T=297160 454240 0 0 $X=296970 $Y=454000
X2289 1 2 70 79 2 872 1 sky130_fd_sc_hd__and2_1 $T=306820 470560 0 0 $X=306630 $Y=470320
X2290 1 2 162 163 2 929 1 sky130_fd_sc_hd__and2_1 $T=330280 465120 1 0 $X=330090 $Y=462160
X2291 1 2 160 163 2 930 1 sky130_fd_sc_hd__and2_1 $T=330280 492320 1 0 $X=330090 $Y=489360
X2292 1 2 166 163 2 937 1 sky130_fd_sc_hd__and2_1 $T=336260 486880 1 0 $X=336070 $Y=483920
X2293 1 2 168 163 2 931 1 sky130_fd_sc_hd__and2_1 $T=337180 497760 0 0 $X=336990 $Y=497520
X2294 1 2 169 163 2 949 1 sky130_fd_sc_hd__and2_1 $T=338560 448800 1 0 $X=338370 $Y=445840
X2295 1 2 171 163 2 935 1 sky130_fd_sc_hd__and2_1 $T=339020 459680 0 0 $X=338830 $Y=459440
X2296 1 2 176 163 2 961 1 sky130_fd_sc_hd__and2_1 $T=346380 481440 1 0 $X=346190 $Y=478480
X2297 1 2 177 163 2 179 1 sky130_fd_sc_hd__and2_1 $T=350980 443360 0 0 $X=350790 $Y=443120
X2298 1 2 178 163 2 971 1 sky130_fd_sc_hd__and2_1 $T=351440 497760 0 0 $X=351250 $Y=497520
X2299 1 2 181 163 2 980 1 sky130_fd_sc_hd__and2_1 $T=356960 454240 1 0 $X=356770 $Y=451280
X2300 1 2 183 163 2 987 1 sky130_fd_sc_hd__and2_1 $T=358800 476000 0 0 $X=358610 $Y=475760
X2301 1 2 185 163 2 1008 1 sky130_fd_sc_hd__and2_1 $T=368000 448800 0 0 $X=367810 $Y=448560
X2302 1 2 186 163 2 1017 1 sky130_fd_sc_hd__and2_1 $T=370760 497760 0 0 $X=370570 $Y=497520
X2303 1 2 187 163 2 1029 1 sky130_fd_sc_hd__and2_1 $T=381340 492320 0 0 $X=381150 $Y=492080
X2304 1 2 188 163 2 1040 1 sky130_fd_sc_hd__and2_1 $T=381800 465120 1 0 $X=381610 $Y=462160
X2305 1 2 190 163 2 1049 1 sky130_fd_sc_hd__and2_1 $T=385480 497760 0 0 $X=385290 $Y=497520
X2306 1 2 193 163 2 1053 1 sky130_fd_sc_hd__and2_1 $T=390540 481440 1 0 $X=390350 $Y=478480
X2307 1 2 197 163 2 1064 1 sky130_fd_sc_hd__and2_1 $T=394220 476000 0 0 $X=394030 $Y=475760
X2308 1 2 200 163 2 1085 1 sky130_fd_sc_hd__and2_1 $T=406180 470560 0 0 $X=405990 $Y=470320
X2309 1 2 201 163 2 1097 1 sky130_fd_sc_hd__and2_1 $T=407560 497760 1 0 $X=407370 $Y=494800
X2310 1 2 205 163 2 1122 1 sky130_fd_sc_hd__and2_1 $T=418140 465120 1 0 $X=417950 $Y=462160
X2311 1 2 206 163 2 1133 1 sky130_fd_sc_hd__and2_1 $T=424120 448800 0 0 $X=423930 $Y=448560
X2312 1 2 207 163 2 1136 1 sky130_fd_sc_hd__and2_1 $T=424120 486880 0 0 $X=423930 $Y=486640
X2313 1 2 209 163 2 1149 1 sky130_fd_sc_hd__and2_1 $T=433320 481440 1 0 $X=433130 $Y=478480
X2314 1 2 212 163 2 1151 1 sky130_fd_sc_hd__and2_1 $T=439760 448800 0 0 $X=439570 $Y=448560
X2315 1 2 213 163 2 1177 1 sky130_fd_sc_hd__and2_1 $T=441140 470560 1 0 $X=440950 $Y=467600
X2316 1 2 215 163 2 1182 1 sky130_fd_sc_hd__and2_1 $T=443900 481440 0 0 $X=443710 $Y=481200
X2317 1 2 217 163 2 1181 1 sky130_fd_sc_hd__and2_1 $T=445280 503200 1 0 $X=445090 $Y=500240
X2318 1 2 221 163 2 1208 1 sky130_fd_sc_hd__and2_1 $T=458620 454240 1 0 $X=458430 $Y=451280
X2319 1 2 222 163 2 1211 1 sky130_fd_sc_hd__and2_1 $T=459080 459680 1 0 $X=458890 $Y=456720
X2320 1 2 223 163 2 1217 1 sky130_fd_sc_hd__and2_1 $T=460920 497760 1 0 $X=460730 $Y=494800
X2321 1 2 226 163 2 1223 1 sky130_fd_sc_hd__and2_1 $T=465520 476000 1 0 $X=465330 $Y=473040
X2322 1 2 227 163 2 1236 1 sky130_fd_sc_hd__and2_1 $T=466440 481440 1 0 $X=466250 $Y=478480
X2323 1 2 234 163 2 1257 1 sky130_fd_sc_hd__and2_1 $T=478860 492320 0 0 $X=478670 $Y=492080
X2324 1 2 236 163 2 1260 1 sky130_fd_sc_hd__and2_1 $T=480240 459680 0 0 $X=480050 $Y=459440
X2325 1 2 240 163 2 1288 1 sky130_fd_sc_hd__and2_1 $T=494500 476000 1 0 $X=494310 $Y=473040
X2326 1 2 243 163 2 1278 1 sky130_fd_sc_hd__and2_1 $T=497260 448800 1 0 $X=497070 $Y=445840
X2327 1 2 244 163 2 1295 1 sky130_fd_sc_hd__and2_1 $T=498180 486880 0 0 $X=497990 $Y=486640
X2328 1 2 247 163 2 1300 1 sky130_fd_sc_hd__and2_1 $T=506920 497760 0 0 $X=506730 $Y=497520
X2329 1 2 251 163 2 1307 1 sky130_fd_sc_hd__and2_1 $T=511060 459680 0 0 $X=510870 $Y=459440
X2330 1 2 193 253 2 1346 1 sky130_fd_sc_hd__and2_1 $T=519340 470560 0 0 $X=519150 $Y=470320
X2331 1 2 162 253 2 1347 1 sky130_fd_sc_hd__and2_1 $T=521640 443360 0 0 $X=521450 $Y=443120
X2332 1 2 160 253 2 1350 1 sky130_fd_sc_hd__and2_1 $T=523940 486880 0 0 $X=523750 $Y=486640
X2333 1 2 197 253 2 1348 1 sky130_fd_sc_hd__and2_1 $T=525320 481440 1 0 $X=525130 $Y=478480
X2334 1 2 168 253 2 1357 1 sky130_fd_sc_hd__and2_1 $T=526700 497760 1 0 $X=526510 $Y=494800
X2335 1 2 176 253 2 1385 1 sky130_fd_sc_hd__and2_1 $T=543260 465120 1 0 $X=543070 $Y=462160
X2336 1 2 187 253 2 1392 1 sky130_fd_sc_hd__and2_1 $T=546480 470560 0 0 $X=546290 $Y=470320
X2337 1 2 209 253 2 1402 1 sky130_fd_sc_hd__and2_1 $T=550620 486880 1 0 $X=550430 $Y=483920
X2338 1 2 186 253 2 1416 1 sky130_fd_sc_hd__and2_1 $T=564420 492320 1 0 $X=564230 $Y=489360
X2339 1 2 171 253 2 1442 1 sky130_fd_sc_hd__and2_1 $T=570860 459680 1 0 $X=570670 $Y=456720
X2340 1 2 183 253 2 1449 1 sky130_fd_sc_hd__and2_1 $T=577300 481440 1 0 $X=577110 $Y=478480
X2341 1 2 166 253 2 1466 1 sky130_fd_sc_hd__and2_1 $T=581440 486880 1 0 $X=581250 $Y=483920
X2342 1 2 188 253 2 1471 1 sky130_fd_sc_hd__and2_1 $T=587420 459680 1 0 $X=587230 $Y=456720
X2343 1 2 178 253 2 1470 1 sky130_fd_sc_hd__and2_1 $T=590640 492320 0 0 $X=590450 $Y=492080
X2344 1 2 200 253 2 1496 1 sky130_fd_sc_hd__and2_1 $T=599380 470560 0 0 $X=599190 $Y=470320
X2345 1 2 201 253 2 1518 1 sky130_fd_sc_hd__and2_1 $T=605360 497760 1 0 $X=605170 $Y=494800
X2346 1 2 185 253 2 1521 1 sky130_fd_sc_hd__and2_1 $T=606740 448800 0 0 $X=606550 $Y=448560
X2347 1 2 205 253 2 1526 1 sky130_fd_sc_hd__and2_1 $T=611340 465120 0 0 $X=611150 $Y=464880
X2348 1 2 215 253 2 1528 1 sky130_fd_sc_hd__and2_1 $T=613640 476000 1 0 $X=613450 $Y=473040
X2349 1 2 190 253 2 1547 1 sky130_fd_sc_hd__and2_1 $T=619160 497760 0 0 $X=618970 $Y=497520
X2350 1 2 181 253 2 1557 1 sky130_fd_sc_hd__and2_1 $T=624680 443360 0 0 $X=624490 $Y=443120
X2351 1 2 206 253 2 1571 1 sky130_fd_sc_hd__and2_1 $T=631580 454240 0 0 $X=631390 $Y=454000
X2352 1 2 213 253 2 1569 1 sky130_fd_sc_hd__and2_1 $T=632960 476000 1 0 $X=632770 $Y=473040
X2353 1 2 217 253 2 1581 1 sky130_fd_sc_hd__and2_1 $T=634800 497760 1 0 $X=634610 $Y=494800
X2354 1 2 234 253 2 1600 1 sky130_fd_sc_hd__and2_1 $T=651360 470560 0 0 $X=651170 $Y=470320
X2355 1 2 207 253 2 1617 1 sky130_fd_sc_hd__and2_1 $T=655960 492320 0 0 $X=655770 $Y=492080
X2356 1 2 212 253 2 1623 1 sky130_fd_sc_hd__and2_1 $T=657340 454240 0 0 $X=657150 $Y=454000
X2357 1 2 218 253 2 1621 1 sky130_fd_sc_hd__and2_1 $T=661940 448800 1 0 $X=661750 $Y=445840
X2358 1 2 223 253 2 1653 1 sky130_fd_sc_hd__and2_1 $T=670220 492320 1 0 $X=670030 $Y=489360
X2359 1 2 226 253 2 1648 1 sky130_fd_sc_hd__and2_1 $T=675280 470560 0 0 $X=675090 $Y=470320
X2360 1 2 221 253 2 1662 1 sky130_fd_sc_hd__and2_1 $T=676660 459680 0 0 $X=676470 $Y=459440
X2361 1 2 222 253 2 1669 1 sky130_fd_sc_hd__and2_1 $T=683560 448800 0 0 $X=683370 $Y=448560
X2362 1 2 227 253 2 1680 1 sky130_fd_sc_hd__and2_1 $T=690000 481440 1 0 $X=689810 $Y=478480
X2363 1 2 247 253 2 1689 1 sky130_fd_sc_hd__and2_1 $T=693680 497760 1 0 $X=693490 $Y=494800
X2364 1 2 236 253 2 1713 1 sky130_fd_sc_hd__and2_1 $T=703340 459680 0 0 $X=703150 $Y=459440
X2365 1 2 244 253 2 1715 1 sky130_fd_sc_hd__and2_1 $T=703340 486880 0 0 $X=703150 $Y=486640
X2366 1 2 240 253 2 1717 1 sky130_fd_sc_hd__and2_1 $T=703800 470560 0 0 $X=703610 $Y=470320
X2367 1 2 243 253 2 1718 1 sky130_fd_sc_hd__and2_1 $T=707480 443360 0 0 $X=707290 $Y=443120
X2368 1 2 251 253 2 1716 1 sky130_fd_sc_hd__and2_1 $T=707480 454240 0 0 $X=707290 $Y=454000
X2369 1 2 ICV_31 $T=17480 459680 1 0 $X=17290 $Y=456720
X2370 1 2 ICV_31 $T=31280 443360 0 0 $X=31090 $Y=443120
X2371 1 2 ICV_31 $T=87400 492320 0 0 $X=87210 $Y=492080
X2372 1 2 ICV_31 $T=101660 459680 1 0 $X=101470 $Y=456720
X2373 1 2 ICV_31 $T=143520 443360 0 0 $X=143330 $Y=443120
X2374 1 2 ICV_31 $T=255760 443360 0 0 $X=255570 $Y=443120
X2375 1 2 ICV_31 $T=270020 465120 1 0 $X=269830 $Y=462160
X2376 1 2 ICV_31 $T=298080 459680 1 0 $X=297890 $Y=456720
X2377 1 2 ICV_31 $T=354200 492320 1 0 $X=354010 $Y=489360
X2378 1 2 ICV_31 $T=368000 454240 0 0 $X=367810 $Y=454000
X2379 1 2 ICV_31 $T=382260 503200 1 0 $X=382070 $Y=500240
X2380 1 2 ICV_31 $T=388240 514080 1 0 $X=388050 $Y=511120
X2381 1 2 ICV_31 $T=410320 454240 1 0 $X=410130 $Y=451280
X2382 1 2 ICV_31 $T=438380 470560 1 0 $X=438190 $Y=467600
X2383 1 2 ICV_31 $T=445280 514080 1 0 $X=445090 $Y=511120
X2384 1 2 ICV_31 $T=473800 514080 1 0 $X=473610 $Y=511120
X2385 1 2 ICV_31 $T=508300 465120 0 0 $X=508110 $Y=464880
X2386 1 2 ICV_31 $T=508300 481440 0 0 $X=508110 $Y=481200
X2387 1 2 ICV_31 $T=522560 459680 1 0 $X=522370 $Y=456720
X2388 1 2 ICV_31 $T=522560 508640 1 0 $X=522370 $Y=505680
X2389 1 2 ICV_31 $T=530840 514080 1 0 $X=530650 $Y=511120
X2390 1 2 ICV_31 $T=536360 443360 0 0 $X=536170 $Y=443120
X2391 1 2 ICV_31 $T=550620 476000 1 0 $X=550430 $Y=473040
X2392 1 2 ICV_31 $T=578680 486880 1 0 $X=578490 $Y=483920
X2393 1 2 ICV_31 $T=620540 503200 0 0 $X=620350 $Y=502960
X2394 1 2 ICV_31 $T=690920 448800 1 0 $X=690730 $Y=445840
X2395 1 2 ICV_31 $T=704720 481440 0 0 $X=704530 $Y=481200
X2396 1 2 320 326 2 323 1 sky130_fd_sc_hd__dlclkp_1 $T=7820 470560 0 0 $X=7630 $Y=470320
X2397 1 2 320 327 2 328 1 sky130_fd_sc_hd__dlclkp_1 $T=7820 492320 1 0 $X=7630 $Y=489360
X2398 1 2 320 324 2 325 1 sky130_fd_sc_hd__dlclkp_1 $T=9200 454240 0 0 $X=9010 $Y=454000
X2399 1 2 320 365 2 370 1 sky130_fd_sc_hd__dlclkp_1 $T=27140 454240 0 0 $X=26950 $Y=454000
X2400 1 2 320 367 2 355 1 sky130_fd_sc_hd__dlclkp_1 $T=27140 476000 0 0 $X=26950 $Y=475760
X2401 1 2 320 391 2 371 1 sky130_fd_sc_hd__dlclkp_1 $T=41400 492320 1 0 $X=41210 $Y=489360
X2402 1 2 320 403 2 404 1 sky130_fd_sc_hd__dlclkp_1 $T=48760 465120 0 0 $X=48570 $Y=464880
X2403 1 2 320 405 2 392 1 sky130_fd_sc_hd__dlclkp_1 $T=51980 454240 1 0 $X=51790 $Y=451280
X2404 1 2 320 431 2 433 1 sky130_fd_sc_hd__dlclkp_1 $T=63480 448800 1 0 $X=63290 $Y=445840
X2405 1 2 320 430 2 407 1 sky130_fd_sc_hd__dlclkp_1 $T=64860 486880 0 0 $X=64670 $Y=486640
X2406 1 2 320 442 2 429 1 sky130_fd_sc_hd__dlclkp_1 $T=69460 470560 1 0 $X=69270 $Y=467600
X2407 1 2 320 463 2 445 1 sky130_fd_sc_hd__dlclkp_1 $T=79580 486880 1 0 $X=79390 $Y=483920
X2408 1 2 320 471 2 474 1 sky130_fd_sc_hd__dlclkp_1 $T=83260 481440 0 0 $X=83070 $Y=481200
X2409 1 2 320 488 2 464 1 sky130_fd_sc_hd__dlclkp_1 $T=92000 454240 1 0 $X=91810 $Y=451280
X2410 1 2 320 479 2 509 1 sky130_fd_sc_hd__dlclkp_1 $T=97060 476000 1 0 $X=96870 $Y=473040
X2411 1 2 320 510 2 487 1 sky130_fd_sc_hd__dlclkp_1 $T=104420 492320 1 0 $X=104230 $Y=489360
X2412 1 2 320 537 2 511 1 sky130_fd_sc_hd__dlclkp_1 $T=118220 454240 0 0 $X=118030 $Y=454000
X2413 1 2 320 555 2 547 1 sky130_fd_sc_hd__dlclkp_1 $T=124200 470560 1 0 $X=124010 $Y=467600
X2414 1 2 320 557 2 559 1 sky130_fd_sc_hd__dlclkp_1 $T=125580 454240 1 0 $X=125390 $Y=451280
X2415 1 2 320 558 2 563 1 sky130_fd_sc_hd__dlclkp_1 $T=125580 486880 1 0 $X=125390 $Y=483920
X2416 1 2 320 582 2 588 1 sky130_fd_sc_hd__dlclkp_1 $T=139380 486880 0 0 $X=139190 $Y=486640
X2417 1 2 320 591 2 594 1 sky130_fd_sc_hd__dlclkp_1 $T=142600 476000 1 0 $X=142410 $Y=473040
X2418 1 2 320 595 2 593 1 sky130_fd_sc_hd__dlclkp_1 $T=148120 459680 0 0 $X=147930 $Y=459440
X2419 1 2 320 612 2 619 1 sky130_fd_sc_hd__dlclkp_1 $T=153640 492320 1 0 $X=153450 $Y=489360
X2420 1 2 320 629 2 636 1 sky130_fd_sc_hd__dlclkp_1 $T=161920 486880 0 0 $X=161730 $Y=486640
X2421 1 2 320 634 2 635 1 sky130_fd_sc_hd__dlclkp_1 $T=165600 470560 0 0 $X=165410 $Y=470320
X2422 1 2 320 650 2 649 1 sky130_fd_sc_hd__dlclkp_1 $T=171120 448800 1 0 $X=170930 $Y=445840
X2423 1 2 320 676 2 682 1 sky130_fd_sc_hd__dlclkp_1 $T=183540 476000 0 0 $X=183350 $Y=475760
X2424 1 2 320 679 2 690 1 sky130_fd_sc_hd__dlclkp_1 $T=189060 448800 0 0 $X=188870 $Y=448560
X2425 1 2 320 687 2 665 1 sky130_fd_sc_hd__dlclkp_1 $T=189520 492320 0 0 $X=189330 $Y=492080
X2426 1 2 320 716 2 722 1 sky130_fd_sc_hd__dlclkp_1 $T=202400 486880 0 0 $X=202210 $Y=486640
X2427 1 2 320 721 2 719 1 sky130_fd_sc_hd__dlclkp_1 $T=205620 481440 1 0 $X=205430 $Y=478480
X2428 1 2 320 724 2 718 1 sky130_fd_sc_hd__dlclkp_1 $T=208380 465120 1 0 $X=208190 $Y=462160
X2429 1 2 320 737 2 746 1 sky130_fd_sc_hd__dlclkp_1 $T=212060 454240 0 0 $X=211870 $Y=454000
X2430 1 2 320 765 2 768 1 sky130_fd_sc_hd__dlclkp_1 $T=228160 459680 1 0 $X=227970 $Y=456720
X2431 1 2 320 766 2 762 1 sky130_fd_sc_hd__dlclkp_1 $T=228160 481440 1 0 $X=227970 $Y=478480
X2432 1 2 320 777 2 786 1 sky130_fd_sc_hd__dlclkp_1 $T=237820 448800 1 0 $X=237630 $Y=445840
X2433 1 2 320 795 2 798 1 sky130_fd_sc_hd__dlclkp_1 $T=245640 476000 1 0 $X=245450 $Y=473040
X2434 1 2 320 805 2 813 1 sky130_fd_sc_hd__dlclkp_1 $T=250700 454240 0 0 $X=250510 $Y=454000
X2435 1 2 320 814 2 817 1 sky130_fd_sc_hd__dlclkp_1 $T=258520 465120 0 0 $X=258330 $Y=464880
X2436 1 2 320 134 2 833 1 sky130_fd_sc_hd__dlclkp_1 $T=265880 448800 1 0 $X=265690 $Y=445840
X2437 1 2 320 832 2 831 1 sky130_fd_sc_hd__dlclkp_1 $T=272780 476000 1 0 $X=272590 $Y=473040
X2438 1 2 320 848 2 851 1 sky130_fd_sc_hd__dlclkp_1 $T=282900 459680 1 0 $X=282710 $Y=456720
X2439 1 2 320 872 2 855 1 sky130_fd_sc_hd__dlclkp_1 $T=300840 476000 1 0 $X=300650 $Y=473040
X2440 1 2 241 931 2 904 1 sky130_fd_sc_hd__dlclkp_1 $T=330740 497760 0 0 $X=330550 $Y=497520
X2441 1 2 241 930 2 875 1 sky130_fd_sc_hd__dlclkp_1 $T=331660 497760 1 0 $X=331470 $Y=494800
X2442 1 2 241 929 2 895 1 sky130_fd_sc_hd__dlclkp_1 $T=332580 459680 0 0 $X=332390 $Y=459440
X2443 1 2 241 935 2 943 1 sky130_fd_sc_hd__dlclkp_1 $T=332580 465120 1 0 $X=332390 $Y=462160
X2444 1 2 241 937 2 884 1 sky130_fd_sc_hd__dlclkp_1 $T=334420 486880 0 0 $X=334230 $Y=486640
X2445 1 2 241 949 2 926 1 sky130_fd_sc_hd__dlclkp_1 $T=340860 448800 1 0 $X=340670 $Y=445840
X2446 1 2 241 961 2 898 1 sky130_fd_sc_hd__dlclkp_1 $T=348680 481440 1 0 $X=348490 $Y=478480
X2447 1 2 241 971 2 968 1 sky130_fd_sc_hd__dlclkp_1 $T=350060 503200 1 0 $X=349870 $Y=500240
X2448 1 2 241 980 2 988 1 sky130_fd_sc_hd__dlclkp_1 $T=356040 448800 0 0 $X=355850 $Y=448560
X2449 1 2 241 987 2 989 1 sky130_fd_sc_hd__dlclkp_1 $T=356960 476000 1 0 $X=356770 $Y=473040
X2450 1 2 241 1017 2 1019 1 sky130_fd_sc_hd__dlclkp_1 $T=370760 492320 0 0 $X=370570 $Y=492080
X2451 1 2 241 1008 2 1025 1 sky130_fd_sc_hd__dlclkp_1 $T=371220 448800 0 0 $X=371030 $Y=448560
X2452 1 2 241 1029 2 978 1 sky130_fd_sc_hd__dlclkp_1 $T=378120 492320 1 0 $X=377930 $Y=489360
X2453 1 2 241 1040 2 1034 1 sky130_fd_sc_hd__dlclkp_1 $T=385020 459680 1 0 $X=384830 $Y=456720
X2454 1 2 241 1053 2 990 1 sky130_fd_sc_hd__dlclkp_1 $T=387780 476000 0 0 $X=387590 $Y=475760
X2455 1 2 241 1049 2 1056 1 sky130_fd_sc_hd__dlclkp_1 $T=387780 497760 0 0 $X=387590 $Y=497520
X2456 1 2 241 1064 2 1073 1 sky130_fd_sc_hd__dlclkp_1 $T=393300 481440 1 0 $X=393110 $Y=478480
X2457 1 2 241 1085 2 1067 1 sky130_fd_sc_hd__dlclkp_1 $T=402960 465120 0 0 $X=402770 $Y=464880
X2458 1 2 241 1097 2 1086 1 sky130_fd_sc_hd__dlclkp_1 $T=406640 497760 0 0 $X=406450 $Y=497520
X2459 1 2 241 1122 2 1130 1 sky130_fd_sc_hd__dlclkp_1 $T=419980 465120 0 0 $X=419790 $Y=464880
X2460 1 2 241 1133 2 1082 1 sky130_fd_sc_hd__dlclkp_1 $T=421360 459680 1 0 $X=421170 $Y=456720
X2461 1 2 241 1136 2 1152 1 sky130_fd_sc_hd__dlclkp_1 $T=424580 497760 1 0 $X=424390 $Y=494800
X2462 1 2 241 1149 2 1118 1 sky130_fd_sc_hd__dlclkp_1 $T=426880 486880 0 0 $X=426690 $Y=486640
X2463 1 2 241 1151 2 1153 1 sky130_fd_sc_hd__dlclkp_1 $T=427800 454240 0 0 $X=427610 $Y=454000
X2464 1 2 241 1177 2 1179 1 sky130_fd_sc_hd__dlclkp_1 $T=440220 470560 0 0 $X=440030 $Y=470320
X2465 1 2 241 1181 2 1184 1 sky130_fd_sc_hd__dlclkp_1 $T=442520 497760 1 0 $X=442330 $Y=494800
X2466 1 2 241 216 2 208 1 sky130_fd_sc_hd__dlclkp_1 $T=442980 443360 0 0 $X=442790 $Y=443120
X2467 1 2 241 1182 2 1180 1 sky130_fd_sc_hd__dlclkp_1 $T=445280 481440 1 0 $X=445090 $Y=478480
X2468 1 2 241 1208 2 1213 1 sky130_fd_sc_hd__dlclkp_1 $T=457700 454240 0 0 $X=457510 $Y=454000
X2469 1 2 241 1211 2 1214 1 sky130_fd_sc_hd__dlclkp_1 $T=461840 459680 0 0 $X=461650 $Y=459440
X2470 1 2 241 1223 2 1232 1 sky130_fd_sc_hd__dlclkp_1 $T=461840 476000 0 0 $X=461650 $Y=475760
X2471 1 2 241 1236 2 1258 1 sky130_fd_sc_hd__dlclkp_1 $T=474260 481440 0 0 $X=474070 $Y=481200
X2472 1 2 241 1257 2 1261 1 sky130_fd_sc_hd__dlclkp_1 $T=477940 497760 1 0 $X=477750 $Y=494800
X2473 1 2 241 1295 2 1296 1 sky130_fd_sc_hd__dlclkp_1 $T=499560 486880 1 0 $X=499370 $Y=483920
X2474 1 2 241 1300 2 1297 1 sky130_fd_sc_hd__dlclkp_1 $T=500480 497760 0 0 $X=500290 $Y=497520
X2475 1 2 241 1307 2 1299 1 sky130_fd_sc_hd__dlclkp_1 $T=505540 465120 1 0 $X=505350 $Y=462160
X2476 1 2 241 1348 2 1356 1 sky130_fd_sc_hd__dlclkp_1 $T=522100 476000 0 0 $X=521910 $Y=475760
X2477 1 2 241 1347 2 1353 1 sky130_fd_sc_hd__dlclkp_1 $T=523940 443360 0 0 $X=523750 $Y=443120
X2478 1 2 241 1357 2 1375 1 sky130_fd_sc_hd__dlclkp_1 $T=536360 497760 1 0 $X=536170 $Y=494800
X2479 1 2 241 1385 2 1386 1 sky130_fd_sc_hd__dlclkp_1 $T=544180 465120 0 0 $X=543990 $Y=464880
X2480 1 2 241 1392 2 1397 1 sky130_fd_sc_hd__dlclkp_1 $T=544180 476000 1 0 $X=543990 $Y=473040
X2481 1 2 241 1402 2 1411 1 sky130_fd_sc_hd__dlclkp_1 $T=551080 481440 0 0 $X=550890 $Y=481200
X2482 1 2 241 1442 2 1443 1 sky130_fd_sc_hd__dlclkp_1 $T=570400 459680 0 0 $X=570210 $Y=459440
X2483 1 2 241 1466 2 1463 1 sky130_fd_sc_hd__dlclkp_1 $T=580980 486880 0 0 $X=580790 $Y=486640
X2484 1 2 241 1471 2 1474 1 sky130_fd_sc_hd__dlclkp_1 $T=583280 454240 0 0 $X=583090 $Y=454000
X2485 1 2 241 1496 2 1497 1 sky130_fd_sc_hd__dlclkp_1 $T=597080 465120 0 0 $X=596890 $Y=464880
X2486 1 2 241 1521 2 1523 1 sky130_fd_sc_hd__dlclkp_1 $T=609500 448800 1 0 $X=609310 $Y=445840
X2487 1 2 241 1518 2 1520 1 sky130_fd_sc_hd__dlclkp_1 $T=609500 492320 1 0 $X=609310 $Y=489360
X2488 1 2 241 1526 2 1527 1 sky130_fd_sc_hd__dlclkp_1 $T=611340 465120 1 0 $X=611150 $Y=462160
X2489 1 2 241 1528 2 1525 1 sky130_fd_sc_hd__dlclkp_1 $T=612720 481440 1 0 $X=612530 $Y=478480
X2490 1 2 241 1547 2 1550 1 sky130_fd_sc_hd__dlclkp_1 $T=618700 497760 1 0 $X=618510 $Y=494800
X2491 1 2 241 1557 2 293 1 sky130_fd_sc_hd__dlclkp_1 $T=626060 448800 1 0 $X=625870 $Y=445840
X2492 1 2 241 1569 2 1578 1 sky130_fd_sc_hd__dlclkp_1 $T=629740 481440 1 0 $X=629550 $Y=478480
X2493 1 2 241 1571 2 1576 1 sky130_fd_sc_hd__dlclkp_1 $T=630660 459680 1 0 $X=630470 $Y=456720
X2494 1 2 241 1600 2 1615 1 sky130_fd_sc_hd__dlclkp_1 $T=647680 476000 1 0 $X=647490 $Y=473040
X2495 1 2 241 1617 2 1620 1 sky130_fd_sc_hd__dlclkp_1 $T=652740 486880 0 0 $X=652550 $Y=486640
X2496 1 2 241 1623 2 1618 1 sky130_fd_sc_hd__dlclkp_1 $T=657340 459680 1 0 $X=657150 $Y=456720
X2497 1 2 241 1648 2 1652 1 sky130_fd_sc_hd__dlclkp_1 $T=668840 470560 0 0 $X=668650 $Y=470320
X2498 1 2 241 1653 2 1649 1 sky130_fd_sc_hd__dlclkp_1 $T=669760 492320 0 0 $X=669570 $Y=492080
X2499 1 2 241 1662 2 1668 1 sky130_fd_sc_hd__dlclkp_1 $T=679420 459680 0 0 $X=679230 $Y=459440
X2500 1 2 241 1680 2 1681 1 sky130_fd_sc_hd__dlclkp_1 $T=686780 476000 0 0 $X=686590 $Y=475760
X2501 1 2 241 1689 2 1691 1 sky130_fd_sc_hd__dlclkp_1 $T=691380 497760 0 0 $X=691190 $Y=497520
X2502 1 2 241 1713 2 1719 1 sky130_fd_sc_hd__dlclkp_1 $T=701960 465120 1 0 $X=701770 $Y=462160
X2503 1 2 241 1715 2 1720 1 sky130_fd_sc_hd__dlclkp_1 $T=701960 492320 1 0 $X=701770 $Y=489360
X2504 1 2 241 1716 2 1721 1 sky130_fd_sc_hd__dlclkp_1 $T=702420 459680 1 0 $X=702230 $Y=456720
X2505 1 2 241 1717 2 1722 1 sky130_fd_sc_hd__dlclkp_1 $T=702420 476000 1 0 $X=702230 $Y=473040
X2506 1 2 241 1718 2 313 1 sky130_fd_sc_hd__dlclkp_1 $T=703800 448800 1 0 $X=703610 $Y=445840
X2507 1 2 ICV_32 $T=100280 503200 1 0 $X=100090 $Y=500240
X2508 1 2 ICV_32 $T=114080 459680 0 0 $X=113890 $Y=459440
X2509 1 2 ICV_32 $T=170200 481440 0 0 $X=170010 $Y=481200
X2510 1 2 ICV_32 $T=240580 459680 1 0 $X=240390 $Y=456720
X2511 1 2 ICV_32 $T=268640 492320 1 0 $X=268450 $Y=489360
X2512 1 2 ICV_32 $T=324760 454240 1 0 $X=324570 $Y=451280
X2513 1 2 ICV_32 $T=324760 481440 1 0 $X=324570 $Y=478480
X2514 1 2 ICV_32 $T=352820 508640 1 0 $X=352630 $Y=505680
X2515 1 2 ICV_32 $T=422740 476000 0 0 $X=422550 $Y=475760
X2516 1 2 ICV_32 $T=450800 448800 0 0 $X=450610 $Y=448560
X2517 1 2 ICV_32 $T=450800 470560 0 0 $X=450610 $Y=470320
X2518 1 2 ICV_32 $T=478860 486880 0 0 $X=478670 $Y=486640
X2519 1 2 ICV_32 $T=521180 470560 1 0 $X=520990 $Y=467600
X2520 1 2 ICV_32 $T=605360 454240 1 0 $X=605170 $Y=451280
X2521 1 2 ICV_32 $T=619160 486880 0 0 $X=618970 $Y=486640
X2522 1 2 ICV_32 $T=689540 465120 1 0 $X=689350 $Y=462160
X2523 1 2 ICV_32 $T=703340 465120 0 0 $X=703150 $Y=464880
X2524 1 2 ICV_32 $T=703340 497760 0 0 $X=703150 $Y=497520
X2525 1 2 ICV_33 $T=86940 508640 0 0 $X=86750 $Y=508400
X2526 1 2 ICV_33 $T=255300 492320 0 0 $X=255110 $Y=492080
X2527 1 2 ICV_33 $T=287960 514080 1 0 $X=287770 $Y=511120
X2528 1 2 ICV_33 $T=573160 514080 1 0 $X=572970 $Y=511120
X2529 1 2 ICV_34 $T=31280 514080 1 0 $X=31090 $Y=511120
X2530 1 2 ICV_34 $T=59800 514080 1 0 $X=59610 $Y=511120
X2531 1 2 ICV_34 $T=88320 514080 1 0 $X=88130 $Y=511120
X2532 1 2 ICV_34 $T=116840 514080 1 0 $X=116650 $Y=511120
X2533 1 2 ICV_34 $T=145360 514080 1 0 $X=145170 $Y=511120
X2534 1 2 ICV_34 $T=173880 514080 1 0 $X=173690 $Y=511120
X2535 1 2 ICV_34 $T=202400 514080 1 0 $X=202210 $Y=511120
X2536 1 2 ICV_34 $T=230920 514080 1 0 $X=230730 $Y=511120
X2537 1 2 ICV_34 $T=259440 514080 1 0 $X=259250 $Y=511120
X2538 1 2 ICV_34 $T=644460 514080 1 0 $X=644270 $Y=511120
X2539 1 2 ICV_34 $T=672980 514080 1 0 $X=672790 $Y=511120
X2540 1 2 ICV_34 $T=701500 514080 1 0 $X=701310 $Y=511120
X2541 1 2 323 15 345 ICV_35 $T=11040 476000 1 0 $X=10850 $Y=473040
X2542 1 2 404 24 416 ICV_35 $T=50600 486880 0 0 $X=50410 $Y=486640
X2543 1 2 457 26 472 ICV_35 $T=78200 470560 0 0 $X=78010 $Y=470320
X2544 1 2 511 7 554 ICV_35 $T=118220 459680 0 0 $X=118030 $Y=459440
X2545 1 2 563 15 575 ICV_35 $T=131100 486880 0 0 $X=130910 $Y=486640
X2546 1 2 594 95 631 ICV_35 $T=157320 470560 0 0 $X=157130 $Y=470320
X2547 1 2 619 8 643 ICV_35 $T=160540 503200 1 0 $X=160350 $Y=500240
X2548 1 2 636 8 623 ICV_35 $T=165600 492320 0 0 $X=165410 $Y=492080
X2549 1 2 665 9 686 ICV_35 $T=182620 503200 0 0 $X=182430 $Y=502960
X2550 1 2 682 82 696 ICV_35 $T=188600 481440 1 0 $X=188410 $Y=478480
X2551 1 2 690 7 723 ICV_35 $T=202400 448800 0 0 $X=202210 $Y=448560
X2552 1 2 718 95 740 ICV_35 $T=206540 459680 0 0 $X=206350 $Y=459440
X2553 1 2 746 99 757 ICV_35 $T=218960 448800 0 0 $X=218770 $Y=448560
X2554 1 2 762 99 790 ICV_35 $T=235980 486880 0 0 $X=235790 $Y=486640
X2555 1 2 813 83 834 ICV_35 $T=264040 454240 1 0 $X=263850 $Y=451280
X2556 1 2 140 83 892 ICV_35 $T=305900 443360 0 0 $X=305710 $Y=443120
X2557 1 2 904 146 950 ICV_35 $T=333040 503200 1 0 $X=332850 $Y=500240
X2558 1 2 153 161 976 ICV_35 $T=347300 448800 1 0 $X=347110 $Y=445840
X2559 1 2 978 154 1024 ICV_35 $T=368460 492320 1 0 $X=368270 $Y=489360
X2560 1 2 1025 161 1047 ICV_35 $T=379040 454240 0 0 $X=378850 $Y=454000
X2561 1 2 1056 150 1077 ICV_35 $T=393300 508640 1 0 $X=393110 $Y=505680
X2562 1 2 1073 165 1093 ICV_35 $T=398820 481440 0 0 $X=398630 $Y=481200
X2563 1 2 1082 150 1098 ICV_35 $T=402960 454240 0 0 $X=402770 $Y=454000
X2564 1 2 1153 159 1173 ICV_35 $T=432400 465120 1 0 $X=432210 $Y=462160
X2565 1 2 1179 146 1191 ICV_35 $T=443440 470560 1 0 $X=443250 $Y=467600
X2566 1 2 1214 154 1259 ICV_35 $T=473340 470560 1 0 $X=473150 $Y=467600
X2567 1 2 1258 149 1262 ICV_35 $T=480700 481440 1 0 $X=480510 $Y=478480
X2568 1 2 1258 144 1212 ICV_35 $T=481160 486880 1 0 $X=480970 $Y=483920
X2569 1 2 1261 149 1273 ICV_35 $T=483000 497760 0 0 $X=482810 $Y=497520
X2570 1 2 245 161 248 ICV_35 $T=499560 448800 1 0 $X=499370 $Y=445840
X2571 1 2 1299 146 1313 ICV_35 $T=500020 465120 0 0 $X=499830 $Y=464880
X2572 1 2 1296 150 1332 ICV_35 $T=511060 492320 0 0 $X=510870 $Y=492080
X2573 1 2 1290 149 1341 ICV_35 $T=512900 459680 1 0 $X=512710 $Y=456720
X2574 1 2 1353 256 1359 ICV_35 $T=525320 448800 1 0 $X=525130 $Y=445840
X2575 1 2 1356 258 1370 ICV_35 $T=527620 481440 1 0 $X=527430 $Y=478480
X2576 1 2 1358 258 1352 ICV_35 $T=529460 497760 0 0 $X=529270 $Y=497520
X2577 1 2 1397 257 1410 ICV_35 $T=548780 470560 0 0 $X=548590 $Y=470320
X2578 1 2 1386 265 1407 ICV_35 $T=550620 459680 0 0 $X=550430 $Y=459440
X2579 1 2 1411 259 1430 ICV_35 $T=557520 481440 0 0 $X=557330 $Y=481200
X2580 1 2 1397 261 1432 ICV_35 $T=558440 470560 0 0 $X=558250 $Y=470320
X2581 1 2 1424 259 1458 ICV_35 $T=572700 497760 1 0 $X=572510 $Y=494800
X2582 1 2 1443 256 1483 ICV_35 $T=585580 459680 0 0 $X=585390 $Y=459440
X2583 1 2 1472 265 1485 ICV_35 $T=585580 508640 1 0 $X=585390 $Y=505680
X2584 1 2 1497 258 1511 ICV_35 $T=598460 465120 1 0 $X=598270 $Y=462160
X2585 1 2 1497 257 1515 ICV_35 $T=599380 476000 1 0 $X=599190 $Y=473040
X2586 1 2 1520 261 1535 ICV_35 $T=608580 508640 0 0 $X=608390 $Y=508400
X2587 1 2 1523 258 1551 ICV_35 $T=621000 459680 1 0 $X=620810 $Y=456720
X2588 1 2 293 258 1604 ICV_35 $T=642620 454240 0 0 $X=642430 $Y=454000
X2589 1 2 293 259 1614 ICV_35 $T=644920 448800 1 0 $X=644730 $Y=445840
X2590 1 2 1620 259 1642 ICV_35 $T=658260 492320 0 0 $X=658070 $Y=492080
X2591 1 2 1652 256 1664 ICV_35 $T=670680 486880 0 0 $X=670490 $Y=486640
X2592 1 2 1668 256 1677 ICV_35 $T=679420 465120 0 0 $X=679230 $Y=464880
X2593 1 2 1649 259 1688 ICV_35 $T=684480 492320 1 0 $X=684290 $Y=489360
X2594 1 2 1691 263 1706 ICV_35 $T=694140 503200 0 0 $X=693950 $Y=502960
X2595 1 2 3 13 338 ICV_36 $T=6900 448800 0 0 $X=6710 $Y=448560
X2596 1 2 392 26 426 ICV_36 $T=51520 454240 0 0 $X=51330 $Y=454000
X2597 1 2 619 19 651 ICV_36 $T=163300 503200 0 0 $X=163110 $Y=502960
X2598 1 2 636 9 671 ICV_36 $T=174340 492320 0 0 $X=174150 $Y=492080
X2599 1 2 722 8 764 ICV_36 $T=219880 492320 0 0 $X=219690 $Y=492080
X2600 1 2 140 95 145 ICV_36 $T=295780 443360 0 0 $X=295590 $Y=443120
X2601 1 2 855 97 891 ICV_36 $T=303600 481440 0 0 $X=303410 $Y=481200
X2602 1 2 968 150 1006 ICV_36 $T=358800 503200 0 0 $X=358610 $Y=502960
X2603 1 2 1019 144 1037 ICV_36 $T=372140 503200 1 0 $X=371950 $Y=500240
X2604 1 2 1214 144 232 ICV_36 $T=469200 459680 1 0 $X=469010 $Y=456720
X2605 1 2 1356 259 1368 ICV_36 $T=525320 486880 1 0 $X=525130 $Y=483920
X2606 1 2 1353 265 1379 ICV_36 $T=533600 448800 1 0 $X=533410 $Y=445840
X2607 1 2 1358 267 1404 ICV_36 $T=542800 497760 1 0 $X=542610 $Y=494800
X2608 1 2 1443 259 1487 ICV_36 $T=584200 465120 0 0 $X=584010 $Y=464880
X2609 1 2 1474 261 1490 ICV_36 $T=584660 443360 0 0 $X=584470 $Y=443120
X2610 1 2 1620 258 1638 ICV_36 $T=655040 508640 1 0 $X=654850 $Y=505680
X2611 1 2 300 261 1628 ICV_36 $T=657800 448800 0 0 $X=657610 $Y=448560
X2612 1 2 1652 257 1663 ICV_36 $T=668840 481440 0 0 $X=668650 $Y=481200
X2613 1 2 1672 258 1708 ICV_36 $T=694140 448800 0 0 $X=693950 $Y=448560
X2614 1 2 3 26 352 ICV_37 $T=19780 454240 1 0 $X=19590 $Y=451280
X2615 1 2 323 26 358 ICV_37 $T=19780 476000 1 0 $X=19590 $Y=473040
X2616 1 2 323 13 348 ICV_37 $T=19780 481440 1 0 $X=19590 $Y=478480
X2617 1 2 328 7 356 ICV_37 $T=19780 486880 1 0 $X=19590 $Y=483920
X2618 1 2 370 7 387 ICV_37 $T=33580 454240 0 0 $X=33390 $Y=454000
X2619 1 2 370 15 389 ICV_37 $T=33580 465120 0 0 $X=33390 $Y=464880
X2620 1 2 371 7 379 ICV_37 $T=33580 492320 0 0 $X=33390 $Y=492080
X2621 1 2 371 24 376 ICV_37 $T=33580 497760 0 0 $X=33390 $Y=497520
X2622 1 2 392 15 366 ICV_37 $T=47840 459680 1 0 $X=47650 $Y=456720
X2623 1 2 392 9 408 ICV_37 $T=47840 465120 1 0 $X=47650 $Y=462160
X2624 1 2 433 8 466 ICV_37 $T=75900 454240 1 0 $X=75710 $Y=451280
X2625 1 2 433 19 462 ICV_37 $T=75900 459680 1 0 $X=75710 $Y=456720
X2626 1 2 429 19 460 ICV_37 $T=75900 481440 1 0 $X=75710 $Y=478480
X2627 1 2 445 26 467 ICV_37 $T=75900 492320 1 0 $X=75710 $Y=489360
X2628 1 2 509 8 523 ICV_37 $T=103960 476000 1 0 $X=103770 $Y=473040
X2629 1 2 474 13 516 ICV_37 $T=103960 486880 1 0 $X=103770 $Y=483920
X2630 1 2 58 26 535 ICV_37 $T=117760 443360 0 0 $X=117570 $Y=443120
X2631 1 2 511 26 543 ICV_37 $T=117760 465120 0 0 $X=117570 $Y=464880
X2632 1 2 559 19 570 ICV_37 $T=132020 454240 1 0 $X=131830 $Y=451280
X2633 1 2 547 7 565 ICV_37 $T=132020 476000 1 0 $X=131830 $Y=473040
X2634 1 2 563 7 578 ICV_37 $T=132020 497760 1 0 $X=131830 $Y=494800
X2635 1 2 588 13 599 ICV_37 $T=145820 492320 0 0 $X=145630 $Y=492080
X2636 1 2 588 24 606 ICV_37 $T=145820 497760 0 0 $X=145630 $Y=497520
X2637 1 2 588 19 601 ICV_37 $T=145820 503200 0 0 $X=145630 $Y=502960
X2638 1 2 594 98 638 ICV_37 $T=160080 481440 1 0 $X=159890 $Y=478480
X2639 1 2 619 7 640 ICV_37 $T=160080 492320 1 0 $X=159890 $Y=489360
X2640 1 2 104 95 107 ICV_37 $T=173880 443360 0 0 $X=173690 $Y=443120
X2641 1 2 649 95 666 ICV_37 $T=173880 448800 0 0 $X=173690 $Y=448560
X2642 1 2 635 82 660 ICV_37 $T=173880 476000 0 0 $X=173690 $Y=475760
X2643 1 2 636 19 658 ICV_37 $T=173880 497760 0 0 $X=173690 $Y=497520
X2644 1 2 675 86 692 ICV_37 $T=188140 459680 1 0 $X=187950 $Y=456720
X2645 1 2 675 85 693 ICV_37 $T=188140 470560 1 0 $X=187950 $Y=467600
X2646 1 2 682 97 694 ICV_37 $T=188140 486880 1 0 $X=187950 $Y=483920
X2647 1 2 718 97 749 ICV_37 $T=216200 470560 1 0 $X=216010 $Y=467600
X2648 1 2 722 19 745 ICV_37 $T=216200 492320 1 0 $X=216010 $Y=489360
X2649 1 2 762 85 770 ICV_37 $T=230000 470560 0 0 $X=229810 $Y=470320
X2650 1 2 786 82 800 ICV_37 $T=244260 448800 1 0 $X=244070 $Y=445840
X2651 1 2 768 85 802 ICV_37 $T=244260 465120 1 0 $X=244070 $Y=462160
X2652 1 2 722 24 793 ICV_37 $T=244260 492320 1 0 $X=244070 $Y=489360
X2653 1 2 813 98 809 ICV_37 $T=272320 459680 1 0 $X=272130 $Y=456720
X2654 1 2 831 98 842 ICV_37 $T=272320 481440 1 0 $X=272130 $Y=478480
X2655 1 2 831 97 857 ICV_37 $T=286120 481440 0 0 $X=285930 $Y=481200
X2656 1 2 884 154 932 ICV_37 $T=328440 486880 1 0 $X=328250 $Y=483920
X2657 1 2 904 154 933 ICV_37 $T=328440 508640 1 0 $X=328250 $Y=505680
X2658 1 2 943 159 956 ICV_37 $T=342240 465120 0 0 $X=342050 $Y=464880
X2659 1 2 943 144 964 ICV_37 $T=342240 470560 0 0 $X=342050 $Y=470320
X2660 1 2 898 161 944 ICV_37 $T=342240 476000 0 0 $X=342050 $Y=475760
X2661 1 2 884 165 965 ICV_37 $T=342240 481440 0 0 $X=342050 $Y=481200
X2662 1 2 875 159 955 ICV_37 $T=342240 492320 0 0 $X=342050 $Y=492080
X2663 1 2 875 161 963 ICV_37 $T=342240 497760 0 0 $X=342050 $Y=497520
X2664 1 2 968 144 974 ICV_37 $T=356500 503200 1 0 $X=356310 $Y=500240
X2665 1 2 988 159 1027 ICV_37 $T=370300 459680 0 0 $X=370110 $Y=459440
X2666 1 2 1034 161 1057 ICV_37 $T=384560 465120 1 0 $X=384370 $Y=462160
X2667 1 2 1034 149 1055 ICV_37 $T=384560 470560 1 0 $X=384370 $Y=467600
X2668 1 2 978 165 1060 ICV_37 $T=384560 497760 1 0 $X=384370 $Y=494800
X2669 1 2 198 165 1088 ICV_37 $T=398360 448800 0 0 $X=398170 $Y=448560
X2670 1 2 1067 161 1079 ICV_37 $T=398360 470560 0 0 $X=398170 $Y=470320
X2671 1 2 1056 149 1083 ICV_37 $T=398360 497760 0 0 $X=398170 $Y=497520
X2672 1 2 1056 161 1091 ICV_37 $T=398360 508640 0 0 $X=398170 $Y=508400
X2673 1 2 1067 146 1114 ICV_37 $T=412620 470560 1 0 $X=412430 $Y=467600
X2674 1 2 1067 159 1108 ICV_37 $T=412620 481440 1 0 $X=412430 $Y=478480
X2675 1 2 1073 161 1117 ICV_37 $T=412620 486880 1 0 $X=412430 $Y=483920
X2676 1 2 1073 150 1113 ICV_37 $T=412620 492320 1 0 $X=412430 $Y=489360
X2677 1 2 1086 154 1124 ICV_37 $T=412620 508640 1 0 $X=412430 $Y=505680
X2678 1 2 1082 149 1147 ICV_37 $T=426420 459680 0 0 $X=426230 $Y=459440
X2679 1 2 1179 144 1218 ICV_37 $T=454480 465120 0 0 $X=454290 $Y=464880
X2680 1 2 1184 165 1219 ICV_37 $T=454480 503200 0 0 $X=454290 $Y=502960
X2681 1 2 219 165 231 ICV_37 $T=468740 448800 1 0 $X=468550 $Y=445840
X2682 1 2 1232 154 1247 ICV_37 $T=468740 492320 1 0 $X=468550 $Y=489360
X2683 1 2 1225 144 1251 ICV_37 $T=468740 497760 1 0 $X=468550 $Y=494800
X2684 1 2 237 161 1267 ICV_37 $T=482540 443360 0 0 $X=482350 $Y=443120
X2685 1 2 1213 150 1268 ICV_37 $T=482540 448800 0 0 $X=482350 $Y=448560
X2686 1 2 1258 146 1264 ICV_37 $T=482540 481440 0 0 $X=482350 $Y=481200
X2687 1 2 1258 159 1228 ICV_37 $T=482540 492320 0 0 $X=482350 $Y=492080
X2688 1 2 1297 154 1327 ICV_37 $T=510600 508640 0 0 $X=510410 $Y=508400
X2689 1 2 1353 263 1388 ICV_37 $T=538660 448800 0 0 $X=538470 $Y=448560
X2690 1 2 1353 267 1389 ICV_37 $T=538660 454240 0 0 $X=538470 $Y=454000
X2691 1 2 1355 267 1391 ICV_37 $T=538660 470560 0 0 $X=538470 $Y=470320
X2692 1 2 1356 265 1393 ICV_37 $T=538660 476000 0 0 $X=538470 $Y=475760
X2693 1 2 1356 267 1394 ICV_37 $T=538660 486880 0 0 $X=538470 $Y=486640
X2694 1 2 1397 263 1419 ICV_37 $T=552920 481440 1 0 $X=552730 $Y=478480
X2695 1 2 277 261 280 ICV_37 $T=566720 443360 0 0 $X=566530 $Y=443120
X2696 1 2 277 267 1441 ICV_37 $T=566720 448800 0 0 $X=566530 $Y=448560
X2697 1 2 1424 263 1448 ICV_37 $T=566720 497760 0 0 $X=566530 $Y=497520
X2698 1 2 1424 258 1437 ICV_37 $T=566720 503200 0 0 $X=566530 $Y=502960
X2699 1 2 277 257 1475 ICV_37 $T=580980 448800 1 0 $X=580790 $Y=445840
X2700 1 2 1520 265 1534 ICV_37 $T=609040 508640 1 0 $X=608850 $Y=505680
X2701 1 2 1523 256 1565 ICV_37 $T=622840 448800 0 0 $X=622650 $Y=448560
X2702 1 2 1523 257 1541 ICV_37 $T=622840 454240 0 0 $X=622650 $Y=454000
X2703 1 2 1550 259 1564 ICV_37 $T=622840 492320 0 0 $X=622650 $Y=492080
X2704 1 2 293 257 1593 ICV_37 $T=637100 448800 1 0 $X=636910 $Y=445840
X2705 1 2 293 256 1589 ICV_37 $T=637100 454240 1 0 $X=636910 $Y=451280
X2706 1 2 1576 258 1590 ICV_37 $T=637100 470560 1 0 $X=636910 $Y=467600
X2707 1 2 1578 261 1594 ICV_37 $T=637100 492320 1 0 $X=636910 $Y=489360
X2708 1 2 1615 267 1651 ICV_37 $T=665160 476000 1 0 $X=664970 $Y=473040
X2709 1 2 1652 259 1675 ICV_37 $T=678960 470560 0 0 $X=678770 $Y=470320
X2710 1 2 1652 258 1678 ICV_37 $T=678960 476000 0 0 $X=678770 $Y=475760
X2711 1 2 1649 263 1674 ICV_37 $T=678960 492320 0 0 $X=678770 $Y=492080
X2712 1 2 1668 261 1700 ICV_37 $T=693220 459680 1 0 $X=693030 $Y=456720
X2713 1 2 1681 265 1702 ICV_37 $T=693220 476000 1 0 $X=693030 $Y=473040
X2714 1 2 1691 265 1704 ICV_37 $T=693220 508640 1 0 $X=693030 $Y=505680
X2715 1 2 355 15 375 355 26 393 ICV_38 $T=29900 476000 1 0 $X=29710 $Y=473040
X2716 1 2 474 15 486 474 19 498 ICV_38 $T=86020 481440 1 0 $X=85830 $Y=478480
X2717 1 2 559 7 566 559 9 584 ICV_38 $T=129260 459680 0 0 $X=129070 $Y=459440
X2718 1 2 762 86 771 768 83 782 ICV_38 $T=227700 470560 1 0 $X=227510 $Y=467600
X2719 1 2 720 26 772 720 7 788 ICV_38 $T=227700 497760 1 0 $X=227510 $Y=494800
X2720 1 2 798 85 815 798 82 820 ICV_38 $T=250700 481440 1 0 $X=250510 $Y=478480
X2721 1 2 855 86 893 855 95 894 ICV_38 $T=307280 476000 1 0 $X=307090 $Y=473040
X2722 1 2 1130 149 1140 1130 161 1157 ICV_38 $T=422280 470560 1 0 $X=422090 $Y=467600
X2723 1 2 1118 150 1174 1118 165 1170 ICV_38 $T=433320 486880 0 0 $X=433130 $Y=486640
X2724 1 2 1179 150 1206 1179 161 1215 ICV_38 $T=450800 476000 1 0 $X=450610 $Y=473040
X2725 1 2 1258 154 1224 1258 161 1221 ICV_38 $T=480240 492320 1 0 $X=480050 $Y=489360
X2726 1 2 1261 161 1275 1261 159 1289 ICV_38 $T=484840 508640 0 0 $X=484650 $Y=508400
X2727 1 2 1355 258 1363 1355 263 1376 ICV_38 $T=527160 465120 1 0 $X=526970 $Y=462160
X2728 1 2 271 259 1408 271 261 1422 ICV_38 $T=548320 448800 0 0 $X=548130 $Y=448560
X2729 1 2 1397 267 1435 1411 256 1439 ICV_38 $T=562580 481440 1 0 $X=562390 $Y=478480
X2730 1 2 1424 265 1460 1424 261 1464 ICV_38 $T=574540 503200 0 0 $X=574350 $Y=502960
X2731 1 2 1463 256 1498 1463 257 1519 ICV_38 $T=593400 486880 1 0 $X=593210 $Y=483920
X2732 1 2 1652 263 1670 1652 267 1684 ICV_38 $T=676660 476000 1 0 $X=676470 $Y=473040
X2733 1 2 1681 259 1693 1681 258 1707 ICV_38 $T=688620 486880 0 0 $X=688430 $Y=486640
X2734 1 2 379 382 21 ICV_39 $T=38640 486880 1 0 $X=38450 $Y=483920
X2735 1 2 424 428 25 ICV_39 $T=62100 497760 0 0 $X=61910 $Y=497520
X2736 1 2 456 459 32 ICV_39 $T=78200 497760 1 0 $X=78010 $Y=494800
X2737 1 2 581 568 32 ICV_39 $T=140760 465120 0 0 $X=140570 $Y=464880
X2738 1 2 600 597 20 ICV_39 $T=155020 497760 1 0 $X=154830 $Y=494800
X2739 1 2 643 630 20 ICV_39 $T=168820 508640 0 0 $X=168630 $Y=508400
X2740 1 2 678 655 92 ICV_39 $T=188600 454240 1 0 $X=188410 $Y=451280
X2741 1 2 761 735 20 ICV_39 $T=230000 486880 1 0 $X=229810 $Y=483920
X2742 1 2 787 769 103 ICV_39 $T=245640 481440 0 0 $X=245450 $Y=481200
X2743 1 2 844 847 102 ICV_39 $T=281060 443360 0 0 $X=280870 $Y=443120
X2744 1 2 845 847 89 ICV_39 $T=281060 459680 0 0 $X=280870 $Y=459440
X2745 1 2 865 847 94 ICV_39 $T=299920 448800 0 0 $X=299730 $Y=448560
X2746 1 2 911 915 157 ICV_39 $T=324300 476000 0 0 $X=324110 $Y=475760
X2747 1 2 948 903 156 ICV_39 $T=340860 492320 1 0 $X=340670 $Y=489360
X2748 1 2 1100 1107 167 ICV_39 $T=413080 465120 1 0 $X=412890 $Y=462160
X2749 1 2 1111 1080 164 ICV_39 $T=421360 470560 0 0 $X=421170 $Y=470320
X2750 1 2 1178 1176 152 ICV_39 $T=442060 454240 1 0 $X=441870 $Y=451280
X2751 1 2 1161 210 151 ICV_39 $T=449420 443360 0 0 $X=449230 $Y=443120
X2752 1 2 1196 1176 155 ICV_39 $T=454020 459680 1 0 $X=453830 $Y=456720
X2753 1 2 1243 1231 167 ICV_39 $T=480700 503200 1 0 $X=480510 $Y=500240
X2754 1 2 1269 1239 170 ICV_39 $T=491740 448800 1 0 $X=491550 $Y=445840
X2755 1 2 1271 1276 157 ICV_39 $T=491740 508640 1 0 $X=491550 $Y=505680
X2756 1 2 1364 1365 264 ICV_39 $T=533600 465120 0 0 $X=533410 $Y=464880
X2757 1 2 1391 1365 275 ICV_39 $T=547860 470560 1 0 $X=547670 $Y=467600
X2758 1 2 1400 1409 275 ICV_39 $T=561660 454240 1 0 $X=561470 $Y=451280
X2759 1 2 1403 1354 269 ICV_39 $T=561660 492320 0 0 $X=561470 $Y=492080
X2760 1 2 1404 1354 275 ICV_39 $T=561660 497760 0 0 $X=561470 $Y=497520
X2761 1 2 1429 1409 264 ICV_39 $T=567180 465120 0 0 $X=566990 $Y=464880
X2762 1 2 1461 279 269 ICV_39 $T=589720 454240 0 0 $X=589530 $Y=454000
X2763 1 2 1596 1592 266 ICV_39 $T=645840 476000 0 0 $X=645650 $Y=475760
X2764 1 2 1604 1575 255 ICV_39 $T=652280 454240 0 0 $X=652090 $Y=454000
X2765 1 2 304 299 255 ICV_39 $T=667460 448800 1 0 $X=667270 $Y=445840
X2766 1 2 1632 1619 275 ICV_39 $T=679420 459680 1 0 $X=679230 $Y=456720
X2767 1 2 1682 1658 255 ICV_39 $T=688160 497760 1 0 $X=687970 $Y=494800
X2768 1 2 419 420 27 ICV_40 $T=63480 470560 1 0 $X=63290 $Y=467600
X2769 1 2 425 428 20 ICV_40 $T=69920 503200 1 0 $X=69730 $Y=500240
X2770 1 2 467 459 30 ICV_40 $T=83720 486880 0 0 $X=83530 $Y=486640
X2771 1 2 489 484 20 ICV_40 $T=97980 486880 1 0 $X=97790 $Y=483920
X2772 1 2 498 484 28 ICV_40 $T=99360 476000 0 0 $X=99170 $Y=475760
X2773 1 2 518 529 22 ICV_40 $T=111780 481440 0 0 $X=111590 $Y=481200
X2774 1 2 586 568 27 ICV_40 $T=142600 448800 1 0 $X=142410 $Y=445840
X2775 1 2 621 616 96 ICV_40 $T=156400 465120 0 0 $X=156210 $Y=464880
X2776 1 2 626 630 22 ICV_40 $T=162840 508640 0 0 $X=162650 $Y=508400
X2777 1 2 640 630 21 ICV_40 $T=167900 497760 0 0 $X=167710 $Y=497520
X2778 1 2 625 630 30 ICV_40 $T=172040 497760 1 0 $X=171850 $Y=494800
X2779 1 2 654 624 30 ICV_40 $T=175260 486880 0 0 $X=175070 $Y=486640
X2780 1 2 680 655 94 ICV_40 $T=186760 454240 0 0 $X=186570 $Y=454000
X2781 1 2 671 624 22 ICV_40 $T=195960 492320 0 0 $X=195770 $Y=492080
X2782 1 2 758 735 30 ICV_40 $T=228160 476000 1 0 $X=227970 $Y=473040
X2783 1 2 771 769 96 ICV_40 $T=234140 476000 1 0 $X=233950 $Y=473040
X2784 1 2 843 826 89 ICV_40 $T=280140 470560 0 0 $X=279950 $Y=470320
X2785 1 2 905 902 155 ICV_40 $T=322460 492320 1 0 $X=322270 $Y=489360
X2786 1 2 965 902 164 ICV_40 $T=356960 486880 1 0 $X=356770 $Y=483920
X2787 1 2 983 915 156 ICV_40 $T=357420 481440 1 0 $X=357230 $Y=478480
X2788 1 2 1001 1000 152 ICV_40 $T=371220 448800 1 0 $X=371030 $Y=445840
X2789 1 2 1023 1014 167 ICV_40 $T=375820 465120 0 0 $X=375630 $Y=464880
X2790 1 2 1057 1051 170 ICV_40 $T=391460 459680 1 0 $X=391270 $Y=456720
X2791 1 2 1092 1095 152 ICV_40 $T=405720 486880 0 0 $X=405530 $Y=486640
X2792 1 2 1078 1065 151 ICV_40 $T=406640 503200 1 0 $X=406450 $Y=500240
X2793 1 2 1119 1129 157 ICV_40 $T=420440 503200 0 0 $X=420250 $Y=502960
X2794 1 2 1132 204 155 ICV_40 $T=422740 454240 1 0 $X=422550 $Y=451280
X2795 1 2 1170 1143 164 ICV_40 $T=438840 492320 0 0 $X=438650 $Y=492080
X2796 1 2 1246 1230 151 ICV_40 $T=476560 476000 0 0 $X=476370 $Y=475760
X2797 1 2 1387 1371 268 ICV_40 $T=545100 481440 0 0 $X=544910 $Y=481200
X2798 1 2 1422 273 268 ICV_40 $T=560740 443360 0 0 $X=560550 $Y=443120
X2799 1 2 1457 1456 269 ICV_40 $T=581900 476000 1 0 $X=581710 $Y=473040
X2800 1 2 1473 1456 275 ICV_40 $T=588800 476000 0 0 $X=588610 $Y=475760
X2801 1 2 1486 1459 255 ICV_40 $T=593400 459680 1 0 $X=593210 $Y=456720
X2802 1 2 1512 1476 268 ICV_40 $T=605820 481440 0 0 $X=605630 $Y=481200
X2803 1 2 1572 1553 270 ICV_40 $T=632040 470560 0 0 $X=631850 $Y=470320
X2804 1 2 1579 1556 262 ICV_40 $T=637560 503200 1 0 $X=637370 $Y=500240
X2805 1 2 1601 1613 269 ICV_40 $T=655040 503200 1 0 $X=654850 $Y=500240
X2806 1 2 1677 1679 262 ICV_40 $T=685860 459680 0 0 $X=685670 $Y=459440
X2807 1 2 41 8 411 ICV_41 $T=51060 448800 0 0 $X=50870 $Y=448560
X2808 1 2 404 8 414 ICV_41 $T=51520 481440 0 0 $X=51330 $Y=481200
X2809 1 2 392 19 412 ICV_41 $T=55660 459680 1 0 $X=55470 $Y=456720
X2810 1 2 457 24 469 ICV_41 $T=80500 470560 1 0 $X=80310 $Y=467600
X2811 1 2 464 7 483 ICV_41 $T=83720 459680 1 0 $X=83530 $Y=456720
X2812 1 2 69 24 562 ICV_41 $T=125580 443360 0 0 $X=125390 $Y=443120
X2813 1 2 635 98 670 ICV_41 $T=177560 481440 1 0 $X=177370 $Y=478480
X2814 1 2 636 13 674 ICV_41 $T=178020 497760 1 0 $X=177830 $Y=494800
X2815 1 2 719 8 761 ICV_41 $T=219880 486880 0 0 $X=219690 $Y=486640
X2816 1 2 833 82 850 ICV_41 $T=276000 448800 0 0 $X=275810 $Y=448560
X2817 1 2 875 146 901 ICV_41 $T=310500 497760 1 0 $X=310310 $Y=494800
X2818 1 2 895 150 916 ICV_41 $T=319240 465120 0 0 $X=319050 $Y=464880
X2819 1 2 978 161 993 ICV_41 $T=359720 492320 0 0 $X=359530 $Y=492080
X2820 1 2 989 150 1015 ICV_41 $T=366160 476000 1 0 $X=365970 $Y=473040
X2821 1 2 198 144 1106 ICV_41 $T=406180 448800 0 0 $X=405990 $Y=448560
X2822 1 2 208 146 1161 ICV_41 $T=430560 448800 1 0 $X=430370 $Y=445840
X2823 1 2 1225 165 1248 ICV_41 $T=471960 503200 0 0 $X=471770 $Y=502960
X2824 1 2 1258 165 1263 ICV_41 $T=490360 481440 0 0 $X=490170 $Y=481200
X2825 1 2 1296 146 1309 ICV_41 $T=500480 486880 0 0 $X=500290 $Y=486640
X2826 1 2 1353 258 1349 ICV_41 $T=528540 448800 0 0 $X=528350 $Y=448560
X2827 1 2 1356 257 1369 ICV_41 $T=528540 476000 0 0 $X=528350 $Y=475760
X2828 1 2 1358 265 1405 ICV_41 $T=546480 486880 0 0 $X=546290 $Y=486640
X2829 1 2 1411 257 1425 ICV_41 $T=556600 486880 0 0 $X=556410 $Y=486640
X2830 1 2 1520 258 1530 ICV_41 $T=616860 508640 1 0 $X=616670 $Y=505680
X2831 1 2 1550 265 1574 ICV_41 $T=626980 508640 1 0 $X=626790 $Y=505680
X2832 1 2 1576 259 1610 ICV_41 $T=644920 465120 1 0 $X=644730 $Y=462160
X2833 1 2 1672 265 310 ICV_41 $T=683560 443360 0 0 $X=683370 $Y=443120
X2834 1 2 371 8 395 ICV_42 $T=39560 497760 1 0 $X=39370 $Y=494800
X2835 1 2 407 9 422 ICV_42 $T=53360 503200 0 0 $X=53170 $Y=502960
X2836 1 2 429 24 435 ICV_42 $T=70840 481440 0 0 $X=70650 $Y=481200
X2837 1 2 464 26 482 ICV_42 $T=83720 454240 1 0 $X=83530 $Y=451280
X2838 1 2 989 149 1039 ICV_42 $T=376280 476000 1 0 $X=376090 $Y=473040
X2839 1 2 990 144 1066 ICV_42 $T=390080 486880 0 0 $X=389890 $Y=486640
X2840 1 2 198 150 1101 ICV_42 $T=404340 448800 1 0 $X=404150 $Y=445840
X2841 1 2 1086 150 1119 ICV_42 $T=412160 503200 0 0 $X=411970 $Y=502960
X2842 1 2 1184 154 1193 ICV_42 $T=446200 503200 0 0 $X=446010 $Y=502960
X2843 1 2 1179 165 1207 ICV_42 $T=451720 470560 1 0 $X=451530 $Y=467600
X2844 1 2 1180 154 1189 ICV_42 $T=456320 492320 1 0 $X=456130 $Y=489360
X2845 1 2 1225 154 1242 ICV_42 $T=466440 508640 0 0 $X=466250 $Y=508400
X2846 1 2 1232 146 1246 ICV_42 $T=468280 476000 0 0 $X=468090 $Y=475760
X2847 1 2 1214 165 233 ICV_42 $T=471960 459680 0 0 $X=471770 $Y=459440
X2848 1 2 1261 154 1272 ICV_42 $T=483460 508640 1 0 $X=483270 $Y=505680
X2849 1 2 1265 144 1285 ICV_42 $T=488520 459680 1 0 $X=488330 $Y=456720
X2850 1 2 1588 265 1602 ICV_42 $T=642620 503200 0 0 $X=642430 $Y=502960
X2851 1 2 1649 265 1685 ICV_42 $T=683100 497760 0 0 $X=682910 $Y=497520
X2852 1 2 328 8 344 ICV_43 $T=10580 497760 0 0 $X=10390 $Y=497520
X2853 1 2 407 24 434 ICV_43 $T=63940 497760 1 0 $X=63750 $Y=494800
X2854 1 2 594 85 617 ICV_43 $T=149040 476000 1 0 $X=148850 $Y=473040
X2855 1 2 665 24 688 ICV_43 $T=190900 503200 0 0 $X=190710 $Y=502960
X2856 1 2 813 86 837 ICV_43 $T=270020 459680 0 0 $X=269830 $Y=459440
X2857 1 2 1056 154 1081 ICV_43 $T=401580 508640 1 0 $X=401390 $Y=505680
X2858 1 2 1152 165 1137 ICV_43 $T=429640 503200 1 0 $X=429450 $Y=500240
X2859 1 2 1180 150 1192 ICV_43 $T=445280 492320 1 0 $X=445090 $Y=489360
X2860 1 2 1261 144 1277 ICV_43 $T=485760 503200 1 0 $X=485570 $Y=500240
X2861 1 2 237 159 242 ICV_43 $T=490360 443360 0 0 $X=490170 $Y=443120
X2862 1 2 1298 146 1294 ICV_43 $T=501860 476000 1 0 $X=501670 $Y=473040
X2863 1 2 1446 265 1462 ICV_43 $T=575460 481440 0 0 $X=575270 $Y=481200
X2864 1 2 1527 265 1572 ICV_43 $T=626060 470560 1 0 $X=625870 $Y=467600
X2865 1 2 1615 256 1627 ICV_43 $T=654120 476000 1 0 $X=653930 $Y=473040
X2866 1 2 1620 261 1645 ICV_43 $T=667000 503200 0 0 $X=666810 $Y=502960
X2867 1 2 1649 258 1682 ICV_43 $T=682180 503200 1 0 $X=681990 $Y=500240
X2868 1 2 381 382 22 395 382 20 ICV_44 $T=39100 503200 1 0 $X=38910 $Y=500240
X2869 1 2 461 448 21 466 448 20 ICV_44 $T=80500 448800 1 0 $X=80310 $Y=445840
X2870 1 2 535 64 30 539 64 28 ICV_44 $T=115920 448800 1 0 $X=115730 $Y=445840
X2871 1 2 659 655 103 672 655 93 ICV_44 $T=179400 459680 1 0 $X=179210 $Y=456720
X2872 1 2 728 732 27 745 732 28 ICV_44 $T=211140 486880 0 0 $X=210950 $Y=486640
X2873 1 2 124 125 103 757 752 101 ICV_44 $T=221260 443360 0 0 $X=221070 $Y=443120
X2874 1 2 764 732 20 772 736 30 ICV_44 $T=230460 492320 0 0 $X=230270 $Y=492080
X2875 1 2 773 752 96 129 125 94 ICV_44 $T=234600 443360 0 0 $X=234410 $Y=443120
X2876 1 2 1108 1080 167 1115 1080 157 ICV_44 $T=413080 476000 1 0 $X=412890 $Y=473040
X2877 1 2 1124 1129 156 1103 1129 164 ICV_44 $T=420440 508640 1 0 $X=420250 $Y=505680
X2878 1 2 1126 1129 151 1137 1138 164 ICV_44 $T=420900 503200 1 0 $X=420710 $Y=500240
X2879 1 2 1166 1138 155 1165 1138 151 ICV_44 $T=438380 497760 0 0 $X=438190 $Y=497520
X2880 1 2 1183 1105 164 1187 1176 170 ICV_44 $T=445280 459680 1 0 $X=445090 $Y=456720
X2881 1 2 1241 1231 155 1252 1231 151 ICV_44 $T=473340 497760 0 0 $X=473150 $Y=497520
X2882 1 2 1272 1276 156 1273 1276 155 ICV_44 $T=491280 497760 0 0 $X=491090 $Y=497520
X2883 1 2 1614 1575 266 298 299 275 ICV_44 $T=653200 448800 1 0 $X=653010 $Y=445840
X2884 1 2 1671 1661 268 1678 1661 255 ICV_44 $T=681260 481440 1 0 $X=681070 $Y=478480
X2885 1 2 333 334 20 ICV_45 $T=11040 486880 1 0 $X=10850 $Y=483920
X2886 1 2 473 470 22 ICV_45 $T=83260 476000 0 0 $X=83070 $Y=475760
X2887 1 2 686 689 22 ICV_45 $T=188600 508640 1 0 $X=188410 $Y=505680
X2888 1 2 754 734 94 ICV_45 $T=223100 465120 0 0 $X=222910 $Y=464880
X2889 1 2 809 808 89 ICV_45 $T=252080 465120 1 0 $X=251890 $Y=462160
X2890 1 2 899 902 152 ICV_45 $T=314640 492320 0 0 $X=314450 $Y=492080
X2891 1 2 909 915 151 ICV_45 $T=321540 486880 1 0 $X=321350 $Y=483920
X2892 1 2 993 994 170 ICV_45 $T=361100 497760 0 0 $X=360910 $Y=497520
X2893 1 2 1116 1129 167 ICV_45 $T=419520 514080 1 0 $X=419330 $Y=511120
X2894 1 2 1189 1105 156 ICV_45 $T=448040 486880 0 0 $X=447850 $Y=486640
X2895 1 2 1233 228 155 ICV_45 $T=464140 454240 0 0 $X=463950 $Y=454000
X2896 1 2 1277 1276 152 ICV_45 $T=490360 492320 0 0 $X=490170 $Y=492080
X2897 1 2 1376 1365 269 ICV_45 $T=537740 459680 1 0 $X=537550 $Y=456720
X2898 1 2 1545 1553 255 ICV_45 $T=620080 476000 1 0 $X=619890 $Y=473040
X2899 1 2 1562 1544 275 ICV_45 $T=626520 476000 1 0 $X=626330 $Y=473040
X2900 1 2 297 1575 270 ICV_45 $T=651360 448800 0 0 $X=651170 $Y=448560
X2901 1 2 1663 1661 264 ICV_45 $T=679420 481440 0 0 $X=679230 $Y=481200
X2902 1 2 1664 1661 262 ICV_45 $T=679420 486880 0 0 $X=679230 $Y=486640
X2903 1 2 457 7 475 452 457 320 ICV_46 $T=74060 465120 0 0 $X=73870 $Y=464880
X2904 1 2 536 26 548 531 536 320 ICV_46 $T=111780 486880 1 0 $X=111590 $Y=483920
X2905 1 2 675 95 691 667 675 320 ICV_46 $T=179400 465120 0 0 $X=179210 $Y=464880
X2906 1 2 722 13 743 713 720 320 ICV_46 $T=201020 492320 1 0 $X=200830 $Y=489360
X2907 1 2 878 85 889 871 878 320 ICV_46 $T=299460 454240 0 0 $X=299270 $Y=454000
X2908 1 2 1225 149 1241 1217 1225 241 ICV_46 $T=459540 497760 0 0 $X=459350 $Y=497520
X2909 1 2 1265 146 1283 1260 1265 241 ICV_46 $T=481160 465120 1 0 $X=480970 $Y=462160
X2910 1 2 1290 146 1302 1278 1290 241 ICV_46 $T=491280 448800 0 0 $X=491090 $Y=448560
X2911 1 2 1298 165 1291 1288 1298 241 ICV_46 $T=495420 476000 0 0 $X=495230 $Y=475760
X2912 1 2 1355 261 1367 1346 1355 241 ICV_46 $T=521640 470560 0 0 $X=521450 $Y=470320
X2913 1 2 1358 259 1374 1350 1358 241 ICV_46 $T=523020 492320 0 0 $X=522830 $Y=492080
X2914 1 2 1424 257 1436 1416 1424 241 ICV_46 $T=557060 497760 1 0 $X=556870 $Y=494800
X2915 1 2 1446 267 1473 1449 1446 241 ICV_46 $T=572700 470560 0 0 $X=572510 $Y=470320
X2916 1 2 1472 259 1494 1470 1472 241 ICV_46 $T=582820 497760 1 0 $X=582630 $Y=494800
X2917 1 2 1588 256 1607 1581 1588 241 ICV_46 $T=637100 497760 0 0 $X=636910 $Y=497520
X2918 1 2 300 259 1647 1621 300 241 ICV_46 $T=655960 443360 0 0 $X=655770 $Y=443120
X2919 1 2 1672 261 1676 1669 1672 241 ICV_46 $T=678960 454240 1 0 $X=678770 $Y=451280
X2920 1 2 323 8 333 ICV_47 $T=5520 481440 0 0 $X=5330 $Y=481200
X2921 1 2 355 24 368 ICV_47 $T=24840 481440 0 0 $X=24650 $Y=481200
X2922 1 2 355 9 372 ICV_47 $T=27600 481440 1 0 $X=27410 $Y=478480
X2923 1 2 392 7 362 ICV_47 $T=42780 454240 0 0 $X=42590 $Y=454000
X2924 1 2 41 19 42 ICV_47 $T=50140 443360 0 0 $X=49950 $Y=443120
X2925 1 2 407 13 424 ICV_47 $T=52440 497760 1 0 $X=52250 $Y=494800
X2926 1 2 429 9 440 ICV_47 $T=62100 481440 0 0 $X=61910 $Y=481200
X2927 1 2 433 7 461 ICV_47 $T=73140 448800 0 0 $X=72950 $Y=448560
X2928 1 2 487 9 499 ICV_47 $T=91540 503200 1 0 $X=91350 $Y=500240
X2929 1 2 474 9 497 ICV_47 $T=94300 492320 1 0 $X=94110 $Y=489360
X2930 1 2 509 13 517 ICV_47 $T=101660 470560 0 0 $X=101470 $Y=470320
X2931 1 2 509 9 518 ICV_47 $T=101660 481440 0 0 $X=101470 $Y=481200
X2932 1 2 536 8 532 ICV_47 $T=115460 492320 1 0 $X=115270 $Y=489360
X2933 1 2 547 8 560 ICV_47 $T=123280 481440 1 0 $X=123090 $Y=478480
X2934 1 2 547 13 567 ICV_47 $T=126500 476000 0 0 $X=126310 $Y=475760
X2935 1 2 547 15 587 ICV_47 $T=135240 476000 0 0 $X=135050 $Y=475760
X2936 1 2 594 82 608 ICV_47 $T=146280 476000 0 0 $X=146090 $Y=475760
X2937 1 2 593 99 645 ICV_47 $T=160540 465120 1 0 $X=160350 $Y=462160
X2938 1 2 593 98 646 ICV_47 $T=160540 470560 1 0 $X=160350 $Y=467600
X2939 1 2 675 98 710 ICV_47 $T=193200 465120 0 0 $X=193010 $Y=464880
X2940 1 2 690 15 725 ICV_47 $T=202400 454240 0 0 $X=202210 $Y=454000
X2941 1 2 690 13 727 ICV_47 $T=203780 448800 1 0 $X=203590 $Y=445840
X2942 1 2 719 15 739 ICV_47 $T=205620 486880 1 0 $X=205430 $Y=483920
X2943 1 2 720 9 789 ICV_47 $T=233680 503200 1 0 $X=233490 $Y=500240
X2944 1 2 762 98 780 ICV_47 $T=234600 481440 1 0 $X=234410 $Y=478480
X2945 1 2 722 7 791 ICV_47 $T=235520 492320 1 0 $X=235330 $Y=489360
X2946 1 2 786 97 799 ICV_47 $T=241960 448800 0 0 $X=241770 $Y=448560
X2947 1 2 798 97 827 ICV_47 $T=258520 486880 0 0 $X=258330 $Y=486640
X2948 1 2 833 95 844 ICV_47 $T=272780 448800 1 0 $X=272590 $Y=445840
X2949 1 2 895 146 896 ICV_47 $T=314180 465120 1 0 $X=313990 $Y=462160
X2950 1 2 895 154 914 ICV_47 $T=318780 470560 0 0 $X=318590 $Y=470320
X2951 1 2 153 144 917 ICV_47 $T=319700 448800 1 0 $X=319510 $Y=445840
X2952 1 2 898 159 938 ICV_47 $T=328900 481440 1 0 $X=328710 $Y=478480
X2953 1 2 153 146 952 ICV_47 $T=333500 443360 0 0 $X=333310 $Y=443120
X2954 1 2 898 144 985 ICV_47 $T=350060 476000 0 0 $X=349870 $Y=475760
X2955 1 2 968 159 986 ICV_47 $T=351900 508640 0 0 $X=351710 $Y=508400
X2956 1 2 988 144 1001 ICV_47 $T=359260 454240 1 0 $X=359070 $Y=451280
X2957 1 2 968 161 995 ICV_47 $T=360640 508640 0 0 $X=360450 $Y=508400
X2958 1 2 989 144 1010 ICV_47 $T=361560 470560 0 0 $X=361370 $Y=470320
X2959 1 2 1025 149 1045 ICV_47 $T=377660 448800 0 0 $X=377470 $Y=448560
X2960 1 2 1034 159 1070 ICV_47 $T=389620 465120 0 0 $X=389430 $Y=464880
X2961 1 2 1056 144 1062 ICV_47 $T=392380 497760 1 0 $X=392190 $Y=494800
X2962 1 2 1067 154 1084 ICV_47 $T=396060 476000 1 0 $X=395870 $Y=473040
X2963 1 2 1082 154 1099 ICV_47 $T=402500 459680 1 0 $X=402310 $Y=456720
X2964 1 2 1118 161 1146 ICV_47 $T=420440 486880 1 0 $X=420250 $Y=483920
X2965 1 2 1118 154 1150 ICV_47 $T=420440 492320 1 0 $X=420250 $Y=489360
X2966 1 2 1130 154 1162 ICV_47 $T=429180 476000 1 0 $X=428990 $Y=473040
X2967 1 2 1153 165 1172 ICV_47 $T=431940 459680 1 0 $X=431750 $Y=456720
X2968 1 2 208 165 1186 ICV_47 $T=442060 448800 0 0 $X=441870 $Y=448560
X2969 1 2 1153 150 1198 ICV_47 $T=445740 459680 0 0 $X=445550 $Y=459440
X2970 1 2 1180 149 1222 ICV_47 $T=454940 481440 0 0 $X=454750 $Y=481200
X2971 1 2 1258 150 1226 ICV_47 $T=483000 486880 0 0 $X=482810 $Y=486640
X2972 1 2 1299 161 1320 ICV_47 $T=500020 459680 0 0 $X=499830 $Y=459440
X2973 1 2 1299 154 1343 ICV_47 $T=512440 470560 1 0 $X=512250 $Y=467600
X2974 1 2 1353 259 1360 ICV_47 $T=525320 454240 1 0 $X=525130 $Y=451280
X2975 1 2 1356 256 1366 ICV_47 $T=526240 486880 0 0 $X=526050 $Y=486640
X2976 1 2 271 256 1398 ICV_47 $T=543720 448800 1 0 $X=543530 $Y=445840
X2977 1 2 1386 267 1400 ICV_47 $T=544180 459680 1 0 $X=543990 $Y=456720
X2978 1 2 1386 258 1427 ICV_47 $T=557060 454240 0 0 $X=556870 $Y=454000
X2979 1 2 277 256 1467 ICV_47 $T=575920 443360 0 0 $X=575730 $Y=443120
X2980 1 2 1472 258 1479 ICV_47 $T=584200 508640 0 0 $X=584010 $Y=508400
X2981 1 2 1472 263 1491 ICV_47 $T=586040 497760 0 0 $X=585850 $Y=497520
X2982 1 2 1523 265 1537 ICV_47 $T=609500 454240 1 0 $X=609310 $Y=451280
X2983 1 2 1520 267 1538 ICV_47 $T=609500 497760 1 0 $X=609310 $Y=494800
X2984 1 2 1576 257 1585 ICV_47 $T=634800 465120 0 0 $X=634610 $Y=464880
X2985 1 2 1578 265 1591 ICV_47 $T=634800 476000 0 0 $X=634610 $Y=475760
X2986 1 2 1618 257 1657 ICV_47 $T=669300 465120 0 0 $X=669110 $Y=464880
X2987 1 2 336 339 21 ICV_48 $T=15640 465120 1 0 $X=15450 $Y=462160
X2988 1 2 337 340 25 ICV_48 $T=15640 492320 1 0 $X=15450 $Y=489360
X2989 1 2 387 385 21 ICV_48 $T=43700 454240 1 0 $X=43510 $Y=451280
X2990 1 2 394 369 28 ICV_48 $T=43700 486880 1 0 $X=43510 $Y=483920
X2991 1 2 501 485 27 ICV_48 $T=99820 454240 1 0 $X=99630 $Y=451280
X2992 1 2 502 485 20 ICV_48 $T=99820 470560 1 0 $X=99630 $Y=467600
X2993 1 2 500 504 32 ICV_48 $T=99820 508640 1 0 $X=99630 $Y=505680
X2994 1 2 585 561 28 ICV_48 $T=141680 470560 0 0 $X=141490 $Y=470320
X2995 1 2 606 597 32 ICV_48 $T=155940 503200 1 0 $X=155750 $Y=500240
X2996 1 2 673 655 96 ICV_48 $T=184000 465120 1 0 $X=183810 $Y=462160
X2997 1 2 652 663 94 ICV_48 $T=184000 476000 1 0 $X=183810 $Y=473040
X2998 1 2 701 704 32 ICV_48 $T=197800 448800 0 0 $X=197610 $Y=448560
X2999 1 2 730 734 89 ICV_48 $T=212060 476000 1 0 $X=211870 $Y=473040
X3000 1 2 731 735 32 ICV_48 $T=212060 481440 1 0 $X=211870 $Y=478480
X3001 1 2 780 769 89 ICV_48 $T=240120 476000 1 0 $X=239930 $Y=473040
X3002 1 2 807 808 101 ICV_48 $T=253920 459680 0 0 $X=253730 $Y=459440
X3003 1 2 913 890 103 ICV_48 $T=324300 465120 1 0 $X=324110 $Y=462160
X3004 1 2 914 897 156 ICV_48 $T=324300 476000 1 0 $X=324110 $Y=473040
X3005 1 2 974 972 152 ICV_48 $T=352360 497760 1 0 $X=352170 $Y=494800
X3006 1 2 1032 1016 151 ICV_48 $T=380420 481440 1 0 $X=380230 $Y=478480
X3007 1 2 1226 1216 157 ICV_48 $T=464600 486880 1 0 $X=464410 $Y=483920
X3008 1 2 1229 1231 170 ICV_48 $T=464600 508640 1 0 $X=464410 $Y=505680
X3009 1 2 1280 1282 157 ICV_48 $T=492660 481440 1 0 $X=492470 $Y=478480
X3010 1 2 1292 1276 164 ICV_48 $T=500480 514080 1 0 $X=500290 $Y=511120
X3011 1 2 1597 1563 268 ICV_48 $T=646760 459680 0 0 $X=646570 $Y=459440
X3012 1 2 1594 1592 268 ICV_48 $T=646760 486880 0 0 $X=646570 $Y=486640
X3013 1 2 1629 1631 269 ICV_48 $T=661020 503200 1 0 $X=660830 $Y=500240
X3014 1 2 325 26 354 354 339 30 ICV_49 $T=16560 459680 0 0 $X=16370 $Y=459440
X3015 1 2 355 8 390 393 369 30 ICV_49 $T=34040 476000 0 0 $X=33850 $Y=475760
X3016 1 2 487 24 500 499 504 22 ICV_49 $T=90160 503200 0 0 $X=89970 $Y=502960
X3017 1 2 81 85 614 615 616 92 ICV_49 $T=146280 454240 0 0 $X=146090 $Y=454000
X3018 1 2 619 15 627 627 630 27 ICV_49 $T=153640 497760 0 0 $X=153450 $Y=497520
X3019 1 2 594 97 632 632 618 103 ICV_49 $T=155940 481440 0 0 $X=155750 $Y=481200
X3020 1 2 817 85 849 849 826 94 ICV_49 $T=272780 470560 1 0 $X=272590 $Y=467600
X3021 1 2 851 99 880 880 864 101 ICV_49 $T=298080 459680 0 0 $X=297890 $Y=459440
X3022 1 2 851 86 883 883 864 96 ICV_49 $T=299920 465120 0 0 $X=299730 $Y=464880
X3023 1 2 875 165 960 963 903 170 ICV_49 $T=338100 497760 1 0 $X=337910 $Y=494800
X3024 1 2 182 165 997 997 184 164 ICV_49 $T=356960 448800 1 0 $X=356770 $Y=445840
X3025 1 2 189 146 194 195 196 155 ICV_49 $T=382260 443360 0 0 $X=382070 $Y=443120
X3026 1 2 1073 154 1110 1113 1095 157 ICV_49 $T=406640 492320 0 0 $X=406450 $Y=492080
X3027 1 2 1299 144 1342 1343 1324 156 ICV_49 $T=511060 465120 0 0 $X=510870 $Y=464880
X3028 1 2 1356 261 1387 1393 1371 270 ICV_49 $T=535900 481440 1 0 $X=535710 $Y=478480
X3029 1 2 1446 259 1493 1493 1456 266 ICV_49 $T=585580 481440 1 0 $X=585390 $Y=478480
X3030 1 2 1463 263 1508 1508 1476 269 ICV_49 $T=595240 492320 0 0 $X=595050 $Y=492080
X3031 1 2 1525 256 1543 1543 1544 262 ICV_49 $T=609500 486880 1 0 $X=609310 $Y=483920
X3032 1 2 1576 263 1584 1590 1563 255 ICV_49 $T=632500 459680 0 0 $X=632310 $Y=459440
X3033 1 2 293 261 1616 1616 1575 268 ICV_49 $T=644920 454240 1 0 $X=644730 $Y=451280
X3034 1 2 1620 257 1639 1636 1631 262 ICV_49 $T=655500 497760 0 0 $X=655310 $Y=497520
X3035 1 2 404 26 418 418 420 30 ICV_50 $T=48300 481440 1 0 $X=48110 $Y=478480
X3036 1 2 588 15 596 599 597 25 ICV_50 $T=139840 497760 1 0 $X=139650 $Y=494800
X3037 1 2 690 26 707 707 704 30 ICV_50 $T=188600 448800 1 0 $X=188410 $Y=445840
X3038 1 2 762 83 784 784 769 92 ICV_50 $T=230460 481440 0 0 $X=230270 $Y=481200
X3039 1 2 720 24 785 785 736 32 ICV_50 $T=230460 503200 0 0 $X=230270 $Y=502960
X3040 1 2 798 99 811 811 812 101 ICV_50 $T=244720 486880 1 0 $X=244530 $Y=483920
X3041 1 2 884 146 900 900 902 151 ICV_50 $T=306360 492320 1 0 $X=306170 $Y=489360
X3042 1 2 878 82 907 889 890 94 ICV_50 $T=312340 459680 1 0 $X=312150 $Y=456720
X3043 1 2 926 144 946 941 945 155 ICV_50 $T=328900 454240 1 0 $X=328710 $Y=451280
X3044 1 2 895 165 947 947 897 164 ICV_50 $T=328900 476000 1 0 $X=328710 $Y=473040
X3045 1 2 1213 165 1266 1267 239 170 ICV_50 $T=476560 448800 1 0 $X=476370 $Y=445840
X3046 1 2 1213 161 1269 1268 1239 157 ICV_50 $T=479320 454240 1 0 $X=479130 $Y=451280
X3047 1 2 1299 159 1314 1313 1324 151 ICV_50 $T=497260 470560 1 0 $X=497070 $Y=467600
X3048 1 2 1296 165 1316 1309 1325 151 ICV_50 $T=497260 492320 1 0 $X=497070 $Y=489360
X3049 1 2 1298 150 1328 1328 1293 157 ICV_50 $T=507840 481440 1 0 $X=507650 $Y=478480
X3050 1 2 1497 265 1510 1510 1516 270 ICV_50 $T=595240 476000 0 0 $X=595050 $Y=475760
X3051 1 2 1618 259 1630 1630 1619 266 ICV_50 $T=651360 459680 0 0 $X=651170 $Y=459440
X3052 1 2 1615 263 1635 1635 1622 269 ICV_50 $T=653660 470560 0 0 $X=653470 $Y=470320
X3053 1 2 374 35 30 33 9 398 ICV_51 $T=35880 448800 0 0 $X=35690 $Y=448560
X3054 1 2 434 428 32 445 9 454 ICV_51 $T=67160 497760 0 0 $X=66970 $Y=497520
X3055 1 2 653 655 89 649 82 672 ICV_51 $T=174340 454240 0 0 $X=174150 $Y=454000
X3056 1 2 664 663 101 682 83 697 ICV_51 $T=185840 481440 0 0 $X=185650 $Y=481200
X3057 1 2 873 876 101 855 82 886 ICV_51 $T=302680 481440 1 0 $X=302490 $Y=478480
X3058 1 2 901 903 151 904 144 921 ICV_51 $T=317400 497760 0 0 $X=317210 $Y=497520
X3059 1 2 986 972 167 968 154 1007 ICV_51 $T=357880 508640 1 0 $X=357690 $Y=505680
X3060 1 2 1012 1016 164 990 146 1032 ICV_51 $T=371680 486880 1 0 $X=371490 $Y=483920
X3061 1 2 1020 1021 164 1019 154 1044 ICV_51 $T=373060 508640 1 0 $X=372870 $Y=505680
X3062 1 2 1077 1065 157 1086 165 1103 ICV_51 $T=400660 503200 0 0 $X=400470 $Y=502960
X3063 1 2 1148 1142 157 1130 159 1171 ICV_51 $T=428720 470560 0 0 $X=428530 $Y=470320
X3064 1 2 1221 1216 170 1232 159 1227 ICV_51 $T=461840 486880 0 0 $X=461650 $Y=486640
X3065 1 2 1262 1216 155 1265 159 1284 ICV_51 $T=483920 470560 1 0 $X=483730 $Y=467600
X3066 1 2 1291 1293 164 1299 165 1321 ICV_51 $T=497260 470560 0 0 $X=497070 $Y=470320
X3067 1 2 1465 279 255 1474 259 1482 ICV_51 $T=582360 454240 1 0 $X=582170 $Y=451280
X3068 1 2 1490 283 268 286 263 289 ICV_51 $T=608120 443360 0 0 $X=607930 $Y=443120
X3069 1 2 1517 1516 262 1525 259 1549 ICV_51 $T=610420 476000 0 0 $X=610230 $Y=475760
X3070 1 2 1514 1516 266 1527 267 1552 ICV_51 $T=611340 459680 0 0 $X=611150 $Y=459440
X3071 1 2 1555 1556 255 1550 267 1580 ICV_51 $T=625600 497760 0 0 $X=625410 $Y=497520
X3072 1 2 1558 287 268 292 265 1583 ICV_51 $T=626980 443360 0 0 $X=626790 $Y=443120
X3073 1 2 1584 1563 269 1576 261 1597 ICV_51 $T=638940 459680 1 0 $X=638750 $Y=456720
X3074 1 2 1583 294 270 293 263 1603 ICV_51 $T=639400 443360 0 0 $X=639210 $Y=443120
X3075 1 2 358 334 30 ICV_52 $T=28060 470560 0 0 $X=27870 $Y=470320
X3076 1 2 477 485 32 ICV_52 $T=90620 448800 1 0 $X=90430 $Y=445840
X3077 1 2 544 513 22 ICV_52 $T=123740 470560 0 0 $X=123550 $Y=470320
X3078 1 2 570 568 28 ICV_52 $T=135700 454240 0 0 $X=135510 $Y=454000
X3079 1 2 577 579 20 ICV_52 $T=143980 492320 1 0 $X=143790 $Y=489360
X3080 1 2 638 618 89 ICV_52 $T=168360 486880 0 0 $X=168170 $Y=486640
X3081 1 2 666 655 102 ICV_52 $T=180780 454240 1 0 $X=180590 $Y=451280
X3082 1 2 725 704 27 ICV_52 $T=210680 459680 1 0 $X=210490 $Y=456720
X3083 1 2 828 808 93 ICV_52 $T=266800 459680 1 0 $X=266610 $Y=456720
X3084 1 2 829 812 96 ICV_52 $T=266800 481440 1 0 $X=266610 $Y=478480
X3085 1 2 850 847 93 ICV_52 $T=282900 454240 1 0 $X=282710 $Y=451280
X3086 1 2 938 915 167 ICV_52 $T=336720 481440 0 0 $X=336530 $Y=481200
X3087 1 2 975 174 167 ICV_52 $T=362480 448800 0 0 $X=362290 $Y=448560
X3088 1 2 1027 1000 167 ICV_52 $T=379040 459680 1 0 $X=378850 $Y=456720
X3089 1 2 1045 1046 155 ICV_52 $T=385940 448800 1 0 $X=385750 $Y=445840
X3090 1 2 1310 1325 167 ICV_52 $T=523020 503200 0 0 $X=522830 $Y=502960
X3091 1 2 1336 1325 152 ICV_52 $T=529000 481440 0 0 $X=528810 $Y=481200
X3092 1 2 1395 1378 266 ICV_52 $T=547400 503200 1 0 $X=547210 $Y=500240
X3093 1 2 1570 1553 266 ICV_52 $T=631580 465120 1 0 $X=631390 $Y=462160
X3094 1 2 342 339 20 ICV_53 $T=15640 454240 0 0 $X=15450 $Y=454000
X3095 1 2 384 385 22 ICV_53 $T=39560 459680 1 0 $X=39370 $Y=456720
X3096 1 2 435 436 32 ICV_53 $T=66240 476000 0 0 $X=66050 $Y=475760
X3097 1 2 476 459 27 ICV_53 $T=86020 503200 1 0 $X=85830 $Y=500240
X3098 1 2 696 705 93 ICV_53 $T=196880 481440 1 0 $X=196690 $Y=478480
X3099 1 2 744 736 28 ICV_53 $T=216660 503200 1 0 $X=216470 $Y=500240
X3100 1 2 868 864 89 ICV_53 $T=294400 465120 0 0 $X=294210 $Y=464880
X3101 1 2 886 876 93 ICV_53 $T=308660 476000 0 0 $X=308470 $Y=475760
X3102 1 2 951 925 170 ICV_53 $T=339480 514080 1 0 $X=339290 $Y=511120
X3103 1 2 1048 1016 155 ICV_53 $T=385020 481440 1 0 $X=384830 $Y=478480
X3104 1 2 1131 1105 152 ICV_53 $T=420900 492320 0 0 $X=420710 $Y=492080
X3105 1 2 1188 1199 167 ICV_53 $T=451720 481440 1 0 $X=451530 $Y=478480
X3106 1 2 1247 1230 156 ICV_53 $T=473340 486880 0 0 $X=473150 $Y=486640
X3107 1 2 1263 1216 164 ICV_53 $T=483000 459680 0 0 $X=482810 $Y=459440
X3108 1 2 1264 1216 151 ICV_53 $T=483000 465120 0 0 $X=482810 $Y=464880
X3109 1 2 1541 287 264 ICV_53 $T=617320 454240 0 0 $X=617130 $Y=454000
X3110 1 2 ICV_54 $T=33580 481440 0 0 $X=33390 $Y=481200
X3111 1 2 ICV_54 $T=75900 503200 1 0 $X=75710 $Y=500240
X3112 1 2 ICV_54 $T=132020 448800 1 0 $X=131830 $Y=445840
X3113 1 2 ICV_54 $T=216200 497760 1 0 $X=216010 $Y=494800
X3114 1 2 ICV_54 $T=258060 476000 0 0 $X=257870 $Y=475760
X3115 1 2 ICV_54 $T=286120 448800 0 0 $X=285930 $Y=448560
X3116 1 2 ICV_54 $T=286120 486880 0 0 $X=285930 $Y=486640
X3117 1 2 ICV_54 $T=300380 465120 1 0 $X=300190 $Y=462160
X3118 1 2 ICV_54 $T=300380 497760 1 0 $X=300190 $Y=494800
X3119 1 2 ICV_54 $T=328440 448800 1 0 $X=328250 $Y=445840
X3120 1 2 ICV_54 $T=384560 454240 1 0 $X=384370 $Y=451280
X3121 1 2 ICV_54 $T=398360 503200 0 0 $X=398170 $Y=502960
X3122 1 2 ICV_54 $T=426420 443360 0 0 $X=426230 $Y=443120
X3123 1 2 ICV_54 $T=426420 470560 0 0 $X=426230 $Y=470320
X3124 1 2 ICV_54 $T=440680 448800 1 0 $X=440490 $Y=445840
X3125 1 2 ICV_54 $T=468740 454240 1 0 $X=468550 $Y=451280
X3126 1 2 ICV_54 $T=482540 508640 0 0 $X=482350 $Y=508400
X3127 1 2 ICV_54 $T=580980 459680 1 0 $X=580790 $Y=456720
X3128 1 2 ICV_54 $T=609040 465120 1 0 $X=608850 $Y=462160
X3129 1 2 114 2 13 1 sky130_fd_sc_hd__clkbuf_16 $T=202400 497760 1 0 $X=202210 $Y=494800
X3130 1 2 117 2 15 1 sky130_fd_sc_hd__clkbuf_16 $T=205160 503200 0 0 $X=204970 $Y=502960
X3131 1 2 120 2 19 1 sky130_fd_sc_hd__clkbuf_16 $T=210220 508640 0 0 $X=210030 $Y=508400
X3132 1 2 121 2 26 1 sky130_fd_sc_hd__clkbuf_16 $T=218500 497760 1 0 $X=218310 $Y=494800
X3133 1 2 122 2 8 1 sky130_fd_sc_hd__clkbuf_16 $T=220340 503200 0 0 $X=220150 $Y=502960
X3134 1 2 126 2 24 1 sky130_fd_sc_hd__clkbuf_16 $T=225860 508640 1 0 $X=225670 $Y=505680
X3135 1 2 127 2 7 1 sky130_fd_sc_hd__clkbuf_16 $T=230460 497760 0 0 $X=230270 $Y=497520
X3136 1 2 128 2 9 1 sky130_fd_sc_hd__clkbuf_16 $T=235060 508640 1 0 $X=234870 $Y=505680
X3137 1 2 121 2 146 1 sky130_fd_sc_hd__clkbuf_16 $T=304060 492320 0 0 $X=303870 $Y=492080
X3138 1 2 127 2 144 1 sky130_fd_sc_hd__clkbuf_16 $T=304520 497760 0 0 $X=304330 $Y=497520
X3139 1 2 117 2 149 1 sky130_fd_sc_hd__clkbuf_16 $T=311880 503200 1 0 $X=311690 $Y=500240
X3140 1 2 114 2 150 1 sky130_fd_sc_hd__clkbuf_16 $T=312340 508640 1 0 $X=312150 $Y=505680
X3141 1 2 120 2 154 1 sky130_fd_sc_hd__clkbuf_16 $T=315560 508640 0 0 $X=315370 $Y=508400
X3142 1 2 128 2 161 1 sky130_fd_sc_hd__clkbuf_16 $T=325680 508640 0 0 $X=325490 $Y=508400
X3143 1 2 126 2 159 1 sky130_fd_sc_hd__clkbuf_16 $T=343620 508640 1 0 $X=343430 $Y=505680
X3144 1 2 122 2 165 1 sky130_fd_sc_hd__clkbuf_16 $T=350520 492320 0 0 $X=350330 $Y=492080
X3145 1 2 249 2 258 1 sky130_fd_sc_hd__clkbuf_16 $T=518880 508640 0 0 $X=518690 $Y=508400
X3146 1 2 192 2 259 1 sky130_fd_sc_hd__clkbuf_16 $T=519800 481440 0 0 $X=519610 $Y=481200
X3147 1 2 224 2 257 1 sky130_fd_sc_hd__clkbuf_16 $T=520260 497760 0 0 $X=520070 $Y=497520
X3148 1 2 214 2 256 1 sky130_fd_sc_hd__clkbuf_16 $T=525320 503200 1 0 $X=525130 $Y=500240
X3149 1 2 238 2 261 1 sky130_fd_sc_hd__clkbuf_16 $T=525320 508640 1 0 $X=525130 $Y=505680
X3150 1 2 260 2 263 1 sky130_fd_sc_hd__clkbuf_16 $T=528540 503200 0 0 $X=528350 $Y=502960
X3151 1 2 203 2 265 1 sky130_fd_sc_hd__clkbuf_16 $T=528540 508640 0 0 $X=528350 $Y=508400
X3152 1 2 276 2 267 1 sky130_fd_sc_hd__clkbuf_16 $T=552460 497760 0 0 $X=552270 $Y=497520
.ENDS
***************************************
.SUBCKT ICV_56 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=14
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=4140 0 0 0 $X=3950 $Y=-240
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__ebufn_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_57 1 2 3 4 5 6 7 8 9 10 11 12 13 14
** N=14 EP=14 IP=16 FDC=72
*.SEEDPROM
X0 1 2 6 7 8 3 4 5 ICV_13 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 12 13 14 9 10 11 ICV_13 $T=0 5440 1 0 $X=-190 $Y=2480
.ENDS
***************************************
.SUBCKT ICV_58 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=10 FDC=38
*.SEEDPROM
X0 1 2 ICV_4 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 6 7 8 3 4 5 ICV_13 $T=3220 0 0 0 $X=3030 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_59 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=10 FDC=36
*.SEEDPROM
X1 1 2 6 7 8 3 4 5 ICV_13 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_60 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=38
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=11500 0 0 0 $X=11310 $Y=-240
X1 1 2 6 7 8 3 4 5 ICV_13 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_61 1 2 3 4
** N=4 EP=4 IP=10 FDC=4
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=1380 0 0 0 $X=1190 $Y=-240
X1 1 2 3 2 4 1 sky130_fd_sc_hd__inv_1 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_62 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=12
*.SEEDPROM
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__ebufn_2 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_63 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=12
*.SEEDPROM
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__ebufn_2 $T=920 0 0 0 $X=730 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_64 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=48
*.SEEDPROM
X0 1 2 3 4 2 5 1 sky130_fd_sc_hd__dfxtp_1 $T=7820 0 0 0 $X=7630 $Y=-240
X1 1 2 6 7 8 ICV_37 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_65 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=6
*.SEEDPROM
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__and2_1 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_66 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=24
*.SEEDPROM
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__dfxtp_1 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__and4b_2 VNB VPB A_N B C D VPWR X VGND
** N=81 EP=9 IP=0 FDC=14
*.SEEDPROM
M0 10 A_N VGND VNB nshort L=0.15 W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75000.2 a=0.063 p=1.14 mult=1 $X=395 $Y=235 $D=9
M1 12 10 11 VNB nshort L=0.15 W=0.42 AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 m=1 r=2.8 sa=75000.2 sb=75002.4 a=0.063 p=1.14 mult=1 $X=1335 $Y=235 $D=9
M2 13 B 12 VNB nshort L=0.15 W=0.42 AD=0.0735 AS=0.0441 PD=0.77 PS=0.63 NRD=34.284 NRS=14.28 m=1 r=2.8 sa=75000.5 sb=75002.1 a=0.063 p=1.14 mult=1 $X=1695 $Y=235 $D=8
M3 14 C 13 VNB nshort L=0.15 W=0.42 AD=0.06195 AS=0.0735 PD=0.715 PS=0.77 NRD=26.424 NRS=34.284 m=1 r=2.8 sa=75001 sb=75001.6 a=0.063 p=1.14 mult=1 $X=2195 $Y=235 $D=8
M4 VGND D 14 VNB nshort L=0.15 W=0.42 AD=0.0816252 AS=0.06195 PD=0.785047 PS=0.715 NRD=0 NRS=26.424 m=1 r=2.8 sa=75001.5 sb=75001.1 a=0.063 p=1.14 mult=1 $X=2640 $Y=235 $D=9
M5 X 11 VGND VNB nshort L=0.15 W=0.65 AD=0.099125 AS=0.126325 PD=0.955 PS=1.21495 NRD=5.532 NRS=13.836 m=1 r=4.33333 sa=75001.4 sb=75000.6 a=0.0975 p=1.6 mult=1 $X=3140 $Y=235 $D=9
M6 VGND 11 X VNB nshort L=0.15 W=0.65 AD=0.169 AS=0.099125 PD=1.82 PS=0.955 NRD=0 NRS=0 m=1 r=4.33333 sa=75001.8 sb=75000.2 a=0.0975 p=1.6 mult=1 $X=3595 $Y=235 $D=9
M7 VPWR A_N 10 VPB phighvt L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75003.4 a=0.063 p=1.14 mult=1 $X=395 $Y=2065 $D=89
M8 11 10 VPWR VPB phighvt L=0.15 W=0.42 AD=0.0987 AS=0.0567 PD=0.89 PS=0.69 NRD=0 NRS=0 m=1 r=2.8 sa=75000.6 sb=75003 a=0.063 p=1.14 mult=1 $X=815 $Y=2065 $D=89
M9 VPWR B 11 VPB phighvt L=0.15 W=0.42 AD=0.1281 AS=0.0987 PD=1.03 PS=0.89 NRD=0 NRS=91.4474 m=1 r=2.8 sa=75001.2 sb=75002.3 a=0.063 p=1.14 mult=1 $X=1435 $Y=2065 $D=89
M10 11 C VPWR VPB phighvt L=0.15 W=0.42 AD=0.06615 AS=0.1281 PD=0.735 PS=1.03 NRD=18.7544 NRS=0 m=1 r=2.8 sa=75002 sb=75001.6 a=0.063 p=1.14 mult=1 $X=2195 $Y=2065 $D=89
M11 VPWR D 11 VPB phighvt L=0.15 W=0.42 AD=0.0847394 AS=0.06615 PD=0.786761 PS=0.735 NRD=25.7873 NRS=0 m=1 r=2.8 sa=75002.4 sb=75001.1 a=0.063 p=1.14 mult=1 $X=2660 $Y=2065 $D=89
M12 X 11 VPWR VPB phighvt L=0.15 W=1 AD=0.1525 AS=0.201761 PD=1.305 PS=1.87324 NRD=5.8903 NRS=0 m=1 r=6.66667 sa=75001.3 sb=75000.6 a=0.15 p=2.3 mult=1 $X=3140 $Y=1485 $D=89
M13 VPWR 11 X VPB phighvt L=0.15 W=1 AD=0.26 AS=0.1525 PD=2.52 PS=1.305 NRD=0 NRS=0 m=1 r=6.66667 sa=75001.8 sb=75000.2 a=0.15 p=2.3 mult=1 $X=3595 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__and4_2 VNB VPB A B C D VPWR X VGND
** N=74 EP=9 IP=0 FDC=12
*.SEEDPROM
M0 13 A 12 VNB nshort L=0.15 W=0.42 AD=0.06195 AS=0.1092 PD=0.715 PS=1.36 NRD=26.424 NRS=0 m=1 r=2.8 sa=75000.2 sb=75002.9 a=0.063 p=1.14 mult=1 $X=395 $Y=235 $D=9
M1 14 B 13 VNB nshort L=0.15 W=0.42 AD=0.0798 AS=0.06195 PD=0.8 PS=0.715 NRD=38.568 NRS=26.424 m=1 r=2.8 sa=75000.6 sb=75002.5 a=0.063 p=1.14 mult=1 $X=840 $Y=235 $D=8
M2 15 C 14 VNB nshort L=0.15 W=0.42 AD=0.0693 AS=0.0798 PD=0.75 PS=0.8 NRD=31.428 NRS=38.568 m=1 r=2.8 sa=75001.2 sb=75001.9 a=0.063 p=1.14 mult=1 $X=1370 $Y=235 $D=8
M3 VGND D 15 VNB nshort L=0.15 W=0.42 AD=0.137501 AS=0.0693 PD=0.993084 PS=0.75 NRD=94.992 NRS=31.428 m=1 r=2.8 sa=75001.6 sb=75001.5 a=0.063 p=1.14 mult=1 $X=1850 $Y=235 $D=9
M4 X 12 VGND VNB nshort L=0.15 W=0.65 AD=0.10725 AS=0.212799 PD=0.98 PS=1.53692 NRD=0 NRS=0.912 m=1 r=4.33333 sa=75001.7 sb=75000.7 a=0.0975 p=1.6 mult=1 $X=2615 $Y=235 $D=9
M5 VGND 12 X VNB nshort L=0.15 W=0.65 AD=0.195 AS=0.10725 PD=1.9 PS=0.98 NRD=6.456 NRS=10.152 m=1 r=4.33333 sa=75002.1 sb=75000.2 a=0.0975 p=1.6 mult=1 $X=3095 $Y=235 $D=9
M6 12 A VPWR VPB phighvt L=0.15 W=0.42 AD=0.07455 AS=0.1092 PD=0.775 PS=1.36 NRD=18.7544 NRS=0 m=1 r=2.8 sa=75000.2 sb=75002.9 a=0.063 p=1.14 mult=1 $X=395 $Y=2065 $D=89
M7 VPWR B 12 VPB phighvt L=0.15 W=0.42 AD=0.0777 AS=0.07455 PD=0.79 PS=0.775 NRD=21.0987 NRS=16.4101 m=1 r=2.8 sa=75000.7 sb=75002.4 a=0.063 p=1.14 mult=1 $X=900 $Y=2065 $D=89
M8 12 C VPWR VPB phighvt L=0.15 W=0.42 AD=0.0588 AS=0.0777 PD=0.7 PS=0.79 NRD=0 NRS=21.0987 m=1 r=2.8 sa=75001.2 sb=75001.9 a=0.063 p=1.14 mult=1 $X=1420 $Y=2065 $D=89
M9 VPWR D 12 VPB phighvt L=0.15 W=0.42 AD=0.165604 AS=0.0588 PD=0.955352 PS=0.7 NRD=123.105 NRS=0 m=1 r=2.8 sa=75001.6 sb=75001.5 a=0.063 p=1.14 mult=1 $X=1850 $Y=2065 $D=89
M10 X 12 VPWR VPB phighvt L=0.15 W=1 AD=0.165 AS=0.394296 PD=1.33 PS=2.27465 NRD=0 NRS=14.7553 m=1 r=6.66667 sa=75001.3 sb=75000.7 a=0.15 p=2.3 mult=1 $X=2615 $Y=1485 $D=89
M11 VPWR 12 X VPB phighvt L=0.15 W=1 AD=0.3 AS=0.165 PD=2.6 PS=1.33 NRD=4.9053 NRS=10.8153 m=1 r=6.66667 sa=75001.7 sb=75000.2 a=0.15 p=2.3 mult=1 $X=3095 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__ebufn_4 VNB VPB A TE_B VPWR Z VGND
** N=111 EP=7 IP=0 FDC=20
*.SEEDPROM
M0 VGND A 9 VNB nshort L=0.15 W=0.65 AD=0.121875 AS=0.169 PD=1.025 PS=1.82 NRD=0 NRS=0 m=1 r=4.33333 sa=75000.2 sb=75000.7 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 8 TE_B VGND VNB nshort L=0.15 W=0.65 AD=0.169 AS=0.121875 PD=1.82 PS=1.025 NRD=0 NRS=18.456 m=1 r=4.33333 sa=75000.7 sb=75000.2 a=0.0975 p=1.6 mult=1 $X=920 $Y=235 $D=9
M2 VGND 8 11 VNB nshort L=0.15 W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 m=1 r=4.33333 sa=75000.2 sb=75003.3 a=0.0975 p=1.6 mult=1 $X=2225 $Y=235 $D=9
M3 11 8 VGND VNB nshort L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75000.6 sb=75002.8 a=0.0975 p=1.6 mult=1 $X=2645 $Y=235 $D=9
M4 VGND 8 11 VNB nshort L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75001 sb=75002.4 a=0.0975 p=1.6 mult=1 $X=3065 $Y=235 $D=9
M5 11 8 VGND VNB nshort L=0.15 W=0.65 AD=0.12675 AS=0.08775 PD=1.04 PS=0.92 NRD=10.152 NRS=0 m=1 r=4.33333 sa=75001.4 sb=75002 a=0.0975 p=1.6 mult=1 $X=3485 $Y=235 $D=9
M6 Z 9 11 VNB nshort L=0.15 W=0.65 AD=0.08775 AS=0.12675 PD=0.92 PS=1.04 NRD=0 NRS=10.152 m=1 r=4.33333 sa=75002 sb=75001.5 a=0.0975 p=1.6 mult=1 $X=4025 $Y=235 $D=9
M7 11 9 Z VNB nshort L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75002.4 sb=75001 a=0.0975 p=1.6 mult=1 $X=4445 $Y=235 $D=9
M8 Z 9 11 VNB nshort L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75002.8 sb=75000.6 a=0.0975 p=1.6 mult=1 $X=4865 $Y=235 $D=9
M9 11 9 Z VNB nshort L=0.15 W=0.65 AD=0.182 AS=0.08775 PD=1.86 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75003.2 sb=75000.2 a=0.0975 p=1.6 mult=1 $X=5285 $Y=235 $D=9
M10 VPWR A 9 VPB phighvt L=0.15 W=1 AD=0.1875 AS=0.26 PD=1.375 PS=2.52 NRD=6.8753 NRS=0 m=1 r=6.66667 sa=75000.2 sb=75000.7 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M11 8 TE_B VPWR VPB phighvt L=0.15 W=1 AD=0.26 AS=0.1875 PD=2.52 PS=1.375 NRD=0 NRS=11.8003 m=1 r=6.66667 sa=75000.7 sb=75000.2 a=0.15 p=2.3 mult=1 $X=920 $Y=1485 $D=89
M12 VPWR TE_B 10 VPB phighvt L=0.15 W=0.94 AD=0.1269 AS=0.2444 PD=1.21 PS=2.4 NRD=0 NRS=0 m=1 r=6.26667 sa=75000.2 sb=75003.6 a=0.141 p=2.18 mult=1 $X=1860 $Y=1545 $D=89
M13 10 TE_B VPWR VPB phighvt L=0.15 W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 m=1 r=6.26667 sa=75000.6 sb=75003.2 a=0.141 p=2.18 mult=1 $X=2280 $Y=1545 $D=89
M14 VPWR TE_B 10 VPB phighvt L=0.15 W=0.94 AD=0.1269 AS=0.1269 PD=1.21 PS=1.21 NRD=0 NRS=0 m=1 r=6.26667 sa=75001 sb=75002.8 a=0.141 p=2.18 mult=1 $X=2700 $Y=1545 $D=89
M15 10 TE_B VPWR VPB phighvt L=0.15 W=0.94 AD=0.363644 AS=0.1269 PD=1.70072 PS=1.21 NRD=17.8088 NRS=0 m=1 r=6.26667 sa=75001.4 sb=75002.4 a=0.141 p=2.18 mult=1 $X=3120 $Y=1545 $D=89
M16 Z 9 10 VPB phighvt L=0.15 W=1 AD=0.135 AS=0.386856 PD=1.27 PS=1.80928 NRD=0 NRS=9.8303 m=1 r=6.66667 sa=75002.2 sb=75001.5 a=0.15 p=2.3 mult=1 $X=4025 $Y=1485 $D=89
M17 10 9 Z VPB phighvt L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75002.7 sb=75001 a=0.15 p=2.3 mult=1 $X=4445 $Y=1485 $D=89
M18 Z 9 10 VPB phighvt L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75003.1 sb=75000.6 a=0.15 p=2.3 mult=1 $X=4865 $Y=1485 $D=89
M19 10 9 Z VPB phighvt L=0.15 W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75003.5 sb=75000.2 a=0.15 p=2.3 mult=1 $X=5285 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__nor4b_2 VNB VPB A B C D_N VPWR Y VGND
** N=132 EP=9 IP=0 FDC=18
*.SEEDPROM
M0 Y A VGND VNB nshort L=0.15 W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 m=1 r=4.33333 sa=75000.2 sb=75001.4 a=0.0975 p=1.6 mult=1 $X=395 $Y=235 $D=9
M1 VGND A Y VNB nshort L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75000.6 sb=75001 a=0.0975 p=1.6 mult=1 $X=815 $Y=235 $D=9
M2 Y B VGND VNB nshort L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75001 sb=75000.6 a=0.0975 p=1.6 mult=1 $X=1235 $Y=235 $D=9
M3 VGND B Y VNB nshort L=0.15 W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75001.4 sb=75000.2 a=0.0975 p=1.6 mult=1 $X=1655 $Y=235 $D=9
M4 Y C VGND VNB nshort L=0.15 W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 m=1 r=4.33333 sa=75000.2 sb=75001.4 a=0.0975 p=1.6 mult=1 $X=2630 $Y=235 $D=9
M5 VGND C Y VNB nshort L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75000.6 sb=75001 a=0.0975 p=1.6 mult=1 $X=3050 $Y=235 $D=9
M6 Y 10 VGND VNB nshort L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75001 sb=75000.6 a=0.0975 p=1.6 mult=1 $X=3470 $Y=235 $D=9
M7 VGND 10 Y VNB nshort L=0.15 W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75001.4 sb=75000.2 a=0.0975 p=1.6 mult=1 $X=3890 $Y=235 $D=9
M8 VGND D_N 10 VNB nshort L=0.15 W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75000.2 a=0.063 p=1.14 mult=1 $X=4830 $Y=465 $D=9
M9 VPWR A 11 VPB phighvt L=0.15 W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 m=1 r=6.66667 sa=75000.2 sb=75001.4 a=0.15 p=2.3 mult=1 $X=395 $Y=1485 $D=89
M10 11 A VPWR VPB phighvt L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75000.6 sb=75001 a=0.15 p=2.3 mult=1 $X=815 $Y=1485 $D=89
M11 12 B 11 VPB phighvt L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75001 sb=75000.6 a=0.15 p=2.3 mult=1 $X=1235 $Y=1485 $D=89
M12 11 B 12 VPB phighvt L=0.15 W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75001.4 sb=75000.2 a=0.15 p=2.3 mult=1 $X=1655 $Y=1485 $D=89
M13 12 C 13 VPB phighvt L=0.15 W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 m=1 r=6.66667 sa=75000.2 sb=75001.4 a=0.15 p=2.3 mult=1 $X=2630 $Y=1485 $D=89
M14 13 C 12 VPB phighvt L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75000.6 sb=75001 a=0.15 p=2.3 mult=1 $X=3050 $Y=1485 $D=89
M15 Y 10 13 VPB phighvt L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75001 sb=75000.6 a=0.15 p=2.3 mult=1 $X=3470 $Y=1485 $D=89
M16 13 10 Y VPB phighvt L=0.15 W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75001.4 sb=75000.2 a=0.15 p=2.3 mult=1 $X=3890 $Y=1485 $D=89
M17 VPWR D_N 10 VPB phighvt L=0.15 W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75000.2 a=0.063 p=1.14 mult=1 $X=4830 $Y=2065 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__and4bb_2 VNB VPB A_N C D B_N VPWR X VGND
** N=85 EP=9 IP=0 FDC=16
*.SEEDPROM
M0 VGND A_N 11 VNB nshort L=0.15 W=0.42 AD=0.0761495 AS=0.1092 PD=0.765421 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75001.1 a=0.063 p=1.14 mult=1 $X=395 $Y=235 $D=9
M1 X 10 VGND VNB nshort L=0.15 W=0.65 AD=0.08775 AS=0.11785 PD=0.92 PS=1.18458 NRD=0 NRS=9.228 m=1 r=4.33333 sa=75000.5 sb=75000.6 a=0.0975 p=1.6 mult=1 $X=870 $Y=235 $D=9
M2 VGND 10 X VNB nshort L=0.15 W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75000.9 sb=75000.2 a=0.0975 p=1.6 mult=1 $X=1290 $Y=235 $D=9
M3 13 11 10 VNB nshort L=0.15 W=0.42 AD=0.0441 AS=0.1092 PD=0.63 PS=1.36 NRD=14.28 NRS=0 m=1 r=2.8 sa=75000.2 sb=75002 a=0.063 p=1.14 mult=1 $X=2230 $Y=235 $D=9
M4 14 12 13 VNB nshort L=0.15 W=0.42 AD=0.06405 AS=0.0441 PD=0.725 PS=0.63 NRD=27.852 NRS=14.28 m=1 r=2.8 sa=75000.5 sb=75001.6 a=0.063 p=1.14 mult=1 $X=2590 $Y=235 $D=8
M5 15 C 14 VNB nshort L=0.15 W=0.42 AD=0.0567 AS=0.06405 PD=0.69 PS=0.725 NRD=22.848 NRS=27.852 m=1 r=2.8 sa=75001 sb=75001.2 a=0.063 p=1.14 mult=1 $X=3045 $Y=235 $D=8
M6 VGND D 15 VNB nshort L=0.15 W=0.42 AD=0.0924 AS=0.0567 PD=0.86 PS=0.69 NRD=47.136 NRS=22.848 m=1 r=2.8 sa=75001.4 sb=75000.8 a=0.063 p=1.14 mult=1 $X=3465 $Y=235 $D=9
M7 12 B_N VGND VNB nshort L=0.15 W=0.42 AD=0.1092 AS=0.0924 PD=1.36 PS=0.86 NRD=0 NRS=0 m=1 r=2.8 sa=75002 sb=75000.2 a=0.063 p=1.14 mult=1 $X=4055 $Y=235 $D=9
M8 VPWR A_N 11 VPB phighvt L=0.15 W=0.42 AD=0.0832606 AS=0.1092 PD=0.783803 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75003.8 a=0.063 p=1.14 mult=1 $X=395 $Y=2065 $D=89
M9 X 10 VPWR VPB phighvt L=0.15 W=1 AD=0.135 AS=0.198239 PD=1.27 PS=1.8662 NRD=0 NRS=9.8303 m=1 r=6.66667 sa=75000.4 sb=75002 a=0.15 p=2.3 mult=1 $X=870 $Y=1485 $D=89
M10 VPWR 10 X VPB phighvt L=0.15 W=1 AD=0.465845 AS=0.135 PD=2.40141 PS=1.27 NRD=14.7553 NRS=0 m=1 r=6.66667 sa=75000.8 sb=75001.6 a=0.15 p=2.3 mult=1 $X=1290 $Y=1485 $D=89
M11 10 11 VPWR VPB phighvt L=0.15 W=0.42 AD=0.0672 AS=0.195655 PD=0.74 PS=1.00859 NRD=21.0987 NRS=4.6886 m=1 r=2.8 sa=75001.9 sb=75002.1 a=0.063 p=1.14 mult=1 $X=2145 $Y=2065 $D=89
M12 VPWR 12 10 VPB phighvt L=0.15 W=0.42 AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=0 m=1 r=2.8 sa=75002.4 sb=75001.6 a=0.063 p=1.14 mult=1 $X=2615 $Y=2065 $D=89
M13 10 C VPWR VPB phighvt L=0.15 W=0.42 AD=0.0567 AS=0.0588 PD=0.69 PS=0.7 NRD=0 NRS=2.3443 m=1 r=2.8 sa=75002.8 sb=75001.2 a=0.063 p=1.14 mult=1 $X=3045 $Y=2065 $D=89
M14 VPWR D 10 VPB phighvt L=0.15 W=0.42 AD=0.0924 AS=0.0567 PD=0.86 PS=0.69 NRD=77.3816 NRS=0 m=1 r=2.8 sa=75003.3 sb=75000.8 a=0.063 p=1.14 mult=1 $X=3465 $Y=2065 $D=89
M15 12 B_N VPWR VPB phighvt L=0.15 W=0.42 AD=0.1092 AS=0.0924 PD=1.36 PS=0.86 NRD=0 NRS=0 m=1 r=2.8 sa=75003.8 sb=75000.2 a=0.063 p=1.14 mult=1 $X=4055 $Y=2065 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__clkbuf_4 VNB VPB A VPWR X VGND
** N=74 EP=6 IP=0 FDC=10
*.SEEDPROM
M0 VGND A 8 VNB nshort L=0.15 W=0.42 AD=0.07035 AS=0.1113 PD=0.755 PS=1.37 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75002 a=0.063 p=1.14 mult=1 $X=400 $Y=235 $D=9
M1 X 8 VGND VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.07035 PD=0.7 PS=0.755 NRD=0 NRS=15.708 m=1 r=2.8 sa=75000.7 sb=75001.5 a=0.063 p=1.14 mult=1 $X=885 $Y=235 $D=9
M2 VGND 8 X VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75001.1 sb=75001.1 a=0.063 p=1.14 mult=1 $X=1315 $Y=235 $D=9
M3 X 8 VGND VNB nshort L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75001.5 sb=75000.6 a=0.063 p=1.14 mult=1 $X=1745 $Y=235 $D=9
M4 VGND 8 X VNB nshort L=0.15 W=0.42 AD=0.1218 AS=0.0588 PD=1.42 PS=0.7 NRD=0 NRS=0 m=1 r=2.8 sa=75002 sb=75000.2 a=0.063 p=1.14 mult=1 $X=2175 $Y=235 $D=9
M5 VPWR A 8 VPB phighvt L=0.15 W=1 AD=0.165 AS=0.265 PD=1.33 PS=2.53 NRD=0 NRS=0 m=1 r=6.66667 sa=75000.2 sb=75002 a=0.15 p=2.3 mult=1 $X=400 $Y=1485 $D=89
M6 X 8 VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.165 PD=1.28 PS=1.33 NRD=0 NRS=9.8303 m=1 r=6.66667 sa=75000.7 sb=75001.5 a=0.15 p=2.3 mult=1 $X=880 $Y=1485 $D=89
M7 VPWR 8 X VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75001.1 sb=75001.1 a=0.15 p=2.3 mult=1 $X=1310 $Y=1485 $D=89
M8 X 8 VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75001.5 sb=75000.7 a=0.15 p=2.3 mult=1 $X=1740 $Y=1485 $D=89
M9 VPWR 8 X VPB phighvt L=0.15 W=1 AD=0.3 AS=0.14 PD=2.6 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75002 sb=75000.2 a=0.15 p=2.3 mult=1 $X=2170 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__conb_1 VPWR VGND LO
** N=16 EP=3 IP=0 FDC=2
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VNB VPB
R0 HI VPWR 0.01 m=1 $[short] $X=105 $Y=1160 $D=280
R1 VGND LO 0.01 m=1 $[short] $X=795 $Y=1160 $D=280
.ENDS
***************************************
.SUBCKT ICV_67 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380
+ 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400
+ 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420
+ 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440
+ 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460
+ 461 462 463 464 465 466 472
** N=1934 EP=467 IP=16805 FDC=47624
X0 1 2 Dpar a=2090.71 p=1485.24 m=1 $[nwdiode] $X=5330 $Y=379385 $D=191
X1 1 2 Dpar a=2090.79 p=1485.14 m=1 $[nwdiode] $X=5330 $Y=384825 $D=191
X2 1 2 Dpar a=2091.36 p=1484.44 m=1 $[nwdiode] $X=5330 $Y=390265 $D=191
X3 1 2 Dpar a=2090.87 p=1485.04 m=1 $[nwdiode] $X=5330 $Y=395705 $D=191
X4 1 2 Dpar a=2090.3 p=1485.74 m=1 $[nwdiode] $X=5330 $Y=401145 $D=191
X5 1 2 Dpar a=2090.3 p=1485.74 m=1 $[nwdiode] $X=5330 $Y=406585 $D=191
X6 1 2 Dpar a=2090.95 p=1484.94 m=1 $[nwdiode] $X=5330 $Y=412025 $D=191
X7 1 2 Dpar a=2091.03 p=1484.84 m=1 $[nwdiode] $X=5330 $Y=417465 $D=191
X8 1 2 Dpar a=2090.63 p=1485.34 m=1 $[nwdiode] $X=5330 $Y=422905 $D=191
X9 1 2 Dpar a=2090.87 p=1485.04 m=1 $[nwdiode] $X=5330 $Y=428345 $D=191
X10 1 2 Dpar a=2090.79 p=1485.14 m=1 $[nwdiode] $X=5330 $Y=433785 $D=191
X11 1 2 Dpar a=2090.63 p=1485.34 m=1 $[nwdiode] $X=5330 $Y=439225 $D=191
X12 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 405280 0 0 $X=5330 $Y=405040
X13 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 421600 1 0 $X=5330 $Y=418640
X14 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 421600 0 0 $X=5330 $Y=421360
X15 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 427040 1 0 $X=5330 $Y=424080
X16 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 427040 0 0 $X=5330 $Y=426800
X17 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=6900 394400 0 0 $X=6710 $Y=394160
X18 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=14260 378080 0 0 $X=14070 $Y=377840
X19 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=14260 405280 1 0 $X=14070 $Y=402320
X20 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=18400 410720 1 0 $X=18210 $Y=407760
X21 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=18400 421600 1 0 $X=18210 $Y=418640
X22 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=25760 437920 0 0 $X=25570 $Y=437680
X23 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=29900 383520 0 0 $X=29710 $Y=383280
X24 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=49680 405280 1 0 $X=49490 $Y=402320
X25 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=65780 416160 1 0 $X=65590 $Y=413200
X26 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=76360 388960 1 0 $X=76170 $Y=386000
X27 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=88320 399840 0 0 $X=88130 $Y=399600
X28 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=94760 405280 1 0 $X=94570 $Y=402320
X29 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=101660 378080 0 0 $X=101470 $Y=377840
X30 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=118220 383520 1 0 $X=118030 $Y=380560
X31 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=118220 388960 0 0 $X=118030 $Y=388720
X32 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=139840 410720 1 0 $X=139650 $Y=407760
X33 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=144440 399840 0 0 $X=144250 $Y=399600
X34 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=154560 416160 0 0 $X=154370 $Y=415920
X35 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=157320 427040 0 0 $X=157130 $Y=426800
X36 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=164680 394400 1 0 $X=164490 $Y=391440
X37 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=166060 399840 0 0 $X=165870 $Y=399600
X38 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=182620 405280 0 0 $X=182430 $Y=405040
X39 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=185840 432480 0 0 $X=185650 $Y=432240
X40 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=195040 427040 1 0 $X=194850 $Y=424080
X41 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=202400 432480 0 0 $X=202210 $Y=432240
X42 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=208840 443360 1 0 $X=208650 $Y=440400
X43 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=220340 437920 0 0 $X=220150 $Y=437680
X44 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=221260 405280 1 0 $X=221070 $Y=402320
X45 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=224480 410720 0 0 $X=224290 $Y=410480
X46 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=228160 437920 1 0 $X=227970 $Y=434960
X47 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=237820 388960 0 0 $X=237630 $Y=388720
X48 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=238740 443360 1 0 $X=238550 $Y=440400
X49 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=240580 410720 1 0 $X=240390 $Y=407760
X50 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=256680 383520 0 0 $X=256490 $Y=383280
X51 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=269560 383520 1 0 $X=269370 $Y=380560
X52 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=270020 378080 0 0 $X=269830 $Y=377840
X53 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=276920 399840 1 0 $X=276730 $Y=396880
X54 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=280140 443360 1 0 $X=279950 $Y=440400
X55 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=296700 399840 0 0 $X=296510 $Y=399600
X56 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=310960 443360 1 0 $X=310770 $Y=440400
X57 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=333960 427040 0 0 $X=333770 $Y=426800
X58 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=336260 399840 1 0 $X=336070 $Y=396880
X59 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=339940 388960 1 0 $X=339750 $Y=386000
X60 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=340400 383520 1 0 $X=340210 $Y=380560
X61 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=342700 421600 0 0 $X=342510 $Y=421360
X62 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=368920 437920 0 0 $X=368730 $Y=437680
X63 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=370760 405280 0 0 $X=370570 $Y=405040
X64 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=378120 437920 0 0 $X=377930 $Y=437680
X65 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=390080 405280 0 0 $X=389890 $Y=405040
X66 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=396980 378080 0 0 $X=396790 $Y=377840
X67 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=396980 416160 0 0 $X=396790 $Y=415920
X68 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=413080 427040 1 0 $X=412890 $Y=424080
X69 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=414920 399840 0 0 $X=414730 $Y=399600
X70 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=420900 416160 0 0 $X=420710 $Y=415920
X71 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=428260 437920 0 0 $X=428070 $Y=437680
X72 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=453100 383520 0 0 $X=452910 $Y=383280
X73 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=455860 405280 1 0 $X=455670 $Y=402320
X74 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=467360 405280 0 0 $X=467170 $Y=405040
X75 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=467360 432480 1 0 $X=467170 $Y=429520
X76 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=476560 432480 1 0 $X=476370 $Y=429520
X77 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=488060 399840 0 0 $X=487870 $Y=399600
X78 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=497260 388960 1 0 $X=497070 $Y=386000
X79 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=497260 410720 1 0 $X=497070 $Y=407760
X80 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=497260 421600 1 0 $X=497070 $Y=418640
X81 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=497720 383520 0 0 $X=497530 $Y=383280
X82 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=505080 410720 1 0 $X=504890 $Y=407760
X83 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=507840 427040 0 0 $X=507650 $Y=426800
X84 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=509220 378080 0 0 $X=509030 $Y=377840
X85 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=515200 383520 1 0 $X=515010 $Y=380560
X86 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=515200 421600 0 0 $X=515010 $Y=421360
X87 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=517960 394400 1 0 $X=517770 $Y=391440
X88 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=522560 427040 0 0 $X=522370 $Y=426800
X89 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=532680 388960 1 0 $X=532490 $Y=386000
X90 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=537740 405280 1 0 $X=537550 $Y=402320
X91 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=539120 410720 0 0 $X=538930 $Y=410480
X92 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=579600 410720 1 0 $X=579410 $Y=407760
X93 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=595240 427040 0 0 $X=595050 $Y=426800
X94 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=603520 437920 1 0 $X=603330 $Y=434960
X95 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=607660 421600 1 0 $X=607470 $Y=418640
X96 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=621460 427040 0 0 $X=621270 $Y=426800
X97 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=622840 416160 1 0 $X=622650 $Y=413200
X98 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=623300 383520 0 0 $X=623110 $Y=383280
X99 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=635720 421600 1 0 $X=635530 $Y=418640
X100 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=652740 405280 1 0 $X=652550 $Y=402320
X101 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=657340 388960 1 0 $X=657150 $Y=386000
X102 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=662860 405280 0 0 $X=662670 $Y=405040
X103 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=677580 378080 0 0 $X=677390 $Y=377840
X104 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=677580 427040 0 0 $X=677390 $Y=426800
X105 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=683100 405280 1 0 $X=682910 $Y=402320
X106 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=687700 388960 1 0 $X=687510 $Y=386000
X107 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=691840 410720 1 0 $X=691650 $Y=407760
X108 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=698740 416160 0 0 $X=698550 $Y=415920
X109 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=720360 421600 0 0 $X=720170 $Y=421360
X110 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 378080 1 180 $X=742710 $Y=377840
X111 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 443360 0 180 $X=742710 $Y=440400
X112 1 2 ICV_1 $T=5520 383520 1 0 $X=5330 $Y=380560
X113 1 2 ICV_1 $T=5520 388960 1 0 $X=5330 $Y=386000
X114 1 2 ICV_1 $T=5520 394400 1 0 $X=5330 $Y=391440
X115 1 2 ICV_1 $T=5520 399840 1 0 $X=5330 $Y=396880
X116 1 2 ICV_1 $T=5520 410720 1 0 $X=5330 $Y=407760
X117 1 2 ICV_1 $T=5520 416160 1 0 $X=5330 $Y=413200
X118 1 2 ICV_1 $T=5520 432480 1 0 $X=5330 $Y=429520
X119 1 2 ICV_1 $T=5520 437920 1 0 $X=5330 $Y=434960
X120 1 2 ICV_1 $T=551540 388960 1 0 $X=551350 $Y=386000
X121 1 2 ICV_1 $T=744280 383520 0 180 $X=742710 $Y=380560
X122 1 2 ICV_1 $T=744280 388960 0 180 $X=742710 $Y=386000
X123 1 2 ICV_1 $T=744280 394400 0 180 $X=742710 $Y=391440
X124 1 2 ICV_1 $T=744280 399840 0 180 $X=742710 $Y=396880
X125 1 2 ICV_1 $T=744280 405280 0 180 $X=742710 $Y=402320
X126 1 2 ICV_1 $T=744280 410720 0 180 $X=742710 $Y=407760
X127 1 2 ICV_1 $T=744280 416160 0 180 $X=742710 $Y=413200
X128 1 2 ICV_1 $T=744280 421600 0 180 $X=742710 $Y=418640
X129 1 2 ICV_1 $T=744280 427040 0 180 $X=742710 $Y=424080
X130 1 2 ICV_1 $T=744280 432480 0 180 $X=742710 $Y=429520
X131 1 2 ICV_1 $T=744280 437920 0 180 $X=742710 $Y=434960
X302 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=6900 405280 0 0 $X=6710 $Y=405040
X303 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=16560 383520 0 0 $X=16370 $Y=383280
X304 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=31740 399840 1 0 $X=31550 $Y=396880
X305 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=34040 416160 0 0 $X=33850 $Y=415920
X306 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=41400 378080 0 0 $X=41210 $Y=377840
X307 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=86480 388960 0 0 $X=86290 $Y=388720
X308 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=98440 388960 0 0 $X=98250 $Y=388720
X309 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=102120 394400 1 0 $X=101930 $Y=391440
X310 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=103960 383520 0 0 $X=103770 $Y=383280
X311 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=111320 378080 0 0 $X=111130 $Y=377840
X312 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=115920 437920 1 0 $X=115730 $Y=434960
X313 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=125580 432480 0 0 $X=125390 $Y=432240
X314 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=126500 378080 0 0 $X=126310 $Y=377840
X315 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=136620 383520 1 0 $X=136430 $Y=380560
X316 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=153640 437920 0 0 $X=153450 $Y=437680
X317 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=166520 388960 0 0 $X=166330 $Y=388720
X318 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=172040 383520 1 0 $X=171850 $Y=380560
X319 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=172040 394400 0 0 $X=171850 $Y=394160
X320 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=172960 405280 1 0 $X=172770 $Y=402320
X321 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=173420 421600 1 0 $X=173230 $Y=418640
X322 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=182160 394400 1 0 $X=181970 $Y=391440
X323 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=186300 405280 1 0 $X=186110 $Y=402320
X324 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=207920 394400 1 0 $X=207730 $Y=391440
X325 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=244720 437920 1 0 $X=244530 $Y=434960
X326 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=256220 383520 1 0 $X=256030 $Y=380560
X327 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=270480 443360 1 0 $X=270290 $Y=440400
X328 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=277840 416160 0 0 $X=277650 $Y=415920
X329 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=298080 378080 0 0 $X=297890 $Y=377840
X330 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=326600 394400 1 0 $X=326410 $Y=391440
X331 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=326600 437920 1 0 $X=326410 $Y=434960
X332 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=327060 437920 0 0 $X=326870 $Y=437680
X333 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=328900 421600 1 0 $X=328710 $Y=418640
X334 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=340400 388960 0 0 $X=340210 $Y=388720
X335 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=340400 437920 0 0 $X=340210 $Y=437680
X336 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=351900 405280 0 0 $X=351710 $Y=405040
X337 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=354200 416160 0 0 $X=354010 $Y=415920
X338 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=378120 421600 0 0 $X=377930 $Y=421360
X339 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=396520 432480 0 0 $X=396330 $Y=432240
X340 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=396520 437920 1 0 $X=396330 $Y=434960
X341 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=410780 399840 1 0 $X=410590 $Y=396880
X342 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=424580 410720 1 0 $X=424390 $Y=407760
X343 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=426880 378080 0 0 $X=426690 $Y=377840
X344 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=435620 399840 0 0 $X=435430 $Y=399600
X345 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=452640 378080 0 0 $X=452450 $Y=377840
X346 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=480700 432480 0 0 $X=480510 $Y=432240
X347 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=496800 416160 0 0 $X=496610 $Y=415920
X348 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=504620 432480 1 0 $X=504430 $Y=429520
X349 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=510140 421600 1 0 $X=509950 $Y=418640
X350 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=511060 388960 0 0 $X=510870 $Y=388720
X351 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=522100 378080 0 0 $X=521910 $Y=377840
X352 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=523020 427040 1 0 $X=522830 $Y=424080
X353 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=536820 421600 0 0 $X=536630 $Y=421360
X354 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=537740 416160 1 0 $X=537550 $Y=413200
X355 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=538660 399840 1 0 $X=538470 $Y=396880
X356 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=549240 394400 0 0 $X=549050 $Y=394160
X357 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=553380 416160 1 0 $X=553190 $Y=413200
X358 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=569020 399840 1 0 $X=568830 $Y=396880
X359 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=579140 432480 1 0 $X=578950 $Y=429520
X360 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=581440 399840 1 0 $X=581250 $Y=396880
X361 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=603520 410720 0 0 $X=603330 $Y=410480
X362 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=607200 416160 1 0 $X=607010 $Y=413200
X363 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=607200 427040 1 0 $X=607010 $Y=424080
X364 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=616860 410720 0 0 $X=616670 $Y=410480
X365 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=623300 437920 0 0 $X=623110 $Y=437680
X366 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=630660 427040 0 0 $X=630470 $Y=426800
X367 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=635720 432480 0 0 $X=635530 $Y=432240
X368 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=651360 405280 0 0 $X=651170 $Y=405040
X369 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=667920 388960 0 0 $X=667730 $Y=388720
X370 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=668380 437920 0 0 $X=668190 $Y=437680
X371 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=677120 394400 1 0 $X=676930 $Y=391440
X372 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=682180 421600 1 0 $X=681990 $Y=418640
X373 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=693220 405280 0 0 $X=693030 $Y=405040
X374 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=707480 383520 0 0 $X=707290 $Y=383280
X375 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=716680 388960 0 0 $X=716490 $Y=388720
X376 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 405280 0 0 $X=740870 $Y=405040
X377 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 410720 0 0 $X=740870 $Y=410480
X378 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 416160 1 0 $X=740870 $Y=413200
X379 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 416160 0 0 $X=740870 $Y=415920
X380 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 421600 0 0 $X=740870 $Y=421360
X381 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 427040 0 0 $X=740870 $Y=426800
X382 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 437920 0 0 $X=740870 $Y=437680
X383 1 2 ICV_3 $T=20240 416160 0 0 $X=20050 $Y=415920
X384 1 2 ICV_3 $T=55200 405280 0 0 $X=55010 $Y=405040
X385 1 2 ICV_3 $T=59340 416160 0 0 $X=59150 $Y=415920
X386 1 2 ICV_3 $T=59340 421600 0 0 $X=59150 $Y=421360
X387 1 2 ICV_3 $T=59340 427040 0 0 $X=59150 $Y=426800
X388 1 2 ICV_3 $T=74060 383520 0 0 $X=73870 $Y=383280
X389 1 2 ICV_3 $T=76360 421600 1 0 $X=76170 $Y=418640
X390 1 2 ICV_3 $T=87400 421600 0 0 $X=87210 $Y=421360
X391 1 2 ICV_3 $T=90160 383520 0 0 $X=89970 $Y=383280
X392 1 2 ICV_3 $T=90160 394400 0 0 $X=89970 $Y=394160
X393 1 2 ICV_3 $T=93380 394400 1 0 $X=93190 $Y=391440
X394 1 2 ICV_3 $T=94300 416160 1 0 $X=94110 $Y=413200
X395 1 2 ICV_3 $T=101660 388960 1 0 $X=101470 $Y=386000
X396 1 2 ICV_3 $T=124660 416160 0 0 $X=124470 $Y=415920
X397 1 2 ICV_3 $T=129720 383520 1 0 $X=129530 $Y=380560
X398 1 2 ICV_3 $T=132480 427040 1 0 $X=132290 $Y=424080
X399 1 2 ICV_3 $T=136160 421600 0 0 $X=135970 $Y=421360
X400 1 2 ICV_3 $T=168820 416160 1 0 $X=168630 $Y=413200
X401 1 2 ICV_3 $T=179400 388960 1 0 $X=179210 $Y=386000
X402 1 2 ICV_3 $T=188140 405280 0 0 $X=187950 $Y=405040
X403 1 2 ICV_3 $T=202400 405280 1 0 $X=202210 $Y=402320
X404 1 2 ICV_3 $T=209760 394400 0 0 $X=209570 $Y=394160
X405 1 2 ICV_3 $T=213900 421600 1 0 $X=213710 $Y=418640
X406 1 2 ICV_3 $T=213900 427040 1 0 $X=213710 $Y=424080
X407 1 2 ICV_3 $T=216660 421600 1 0 $X=216470 $Y=418640
X408 1 2 ICV_3 $T=226320 388960 0 0 $X=226130 $Y=388720
X409 1 2 ICV_3 $T=230460 399840 0 0 $X=230270 $Y=399600
X410 1 2 ICV_3 $T=235520 394400 0 0 $X=235330 $Y=394160
X411 1 2 ICV_3 $T=236900 427040 1 0 $X=236710 $Y=424080
X412 1 2 ICV_3 $T=249780 427040 0 0 $X=249590 $Y=426800
X413 1 2 ICV_3 $T=263580 405280 1 0 $X=263390 $Y=402320
X414 1 2 ICV_3 $T=294860 427040 0 0 $X=294670 $Y=426800
X415 1 2 ICV_3 $T=298080 432480 1 0 $X=297890 $Y=429520
X416 1 2 ICV_3 $T=311880 383520 0 0 $X=311690 $Y=383280
X417 1 2 ICV_3 $T=326140 416160 1 0 $X=325950 $Y=413200
X418 1 2 ICV_3 $T=327060 432480 0 0 $X=326870 $Y=432240
X419 1 2 ICV_3 $T=364780 443360 1 0 $X=364590 $Y=440400
X420 1 2 ICV_3 $T=370760 394400 0 0 $X=370570 $Y=394160
X421 1 2 ICV_3 $T=396060 399840 0 0 $X=395870 $Y=399600
X422 1 2 ICV_3 $T=396060 437920 0 0 $X=395870 $Y=437680
X423 1 2 ICV_3 $T=403420 383520 1 0 $X=403230 $Y=380560
X424 1 2 ICV_3 $T=419060 383520 0 0 $X=418870 $Y=383280
X425 1 2 ICV_3 $T=424120 394400 0 0 $X=423930 $Y=394160
X426 1 2 ICV_3 $T=449420 388960 1 0 $X=449230 $Y=386000
X427 1 2 ICV_3 $T=452180 388960 0 0 $X=451990 $Y=388720
X428 1 2 ICV_3 $T=452180 432480 0 0 $X=451990 $Y=432240
X429 1 2 ICV_3 $T=480240 437920 0 0 $X=480050 $Y=437680
X430 1 2 ICV_3 $T=494500 388960 1 0 $X=494310 $Y=386000
X431 1 2 ICV_3 $T=508300 399840 0 0 $X=508110 $Y=399600
X432 1 2 ICV_3 $T=508300 437920 0 0 $X=508110 $Y=437680
X433 1 2 ICV_3 $T=509220 405280 1 0 $X=509030 $Y=402320
X434 1 2 ICV_3 $T=515200 378080 0 0 $X=515010 $Y=377840
X435 1 2 ICV_3 $T=522560 388960 1 0 $X=522370 $Y=386000
X436 1 2 ICV_3 $T=536360 383520 1 0 $X=536170 $Y=380560
X437 1 2 ICV_3 $T=536360 383520 0 0 $X=536170 $Y=383280
X438 1 2 ICV_3 $T=536360 437920 0 0 $X=536170 $Y=437680
X439 1 2 ICV_3 $T=539120 388960 0 0 $X=538930 $Y=388720
X440 1 2 ICV_3 $T=564420 388960 0 0 $X=564230 $Y=388720
X441 1 2 ICV_3 $T=576380 405280 1 0 $X=576190 $Y=402320
X442 1 2 ICV_3 $T=578680 416160 1 0 $X=578490 $Y=413200
X443 1 2 ICV_3 $T=578680 437920 1 0 $X=578490 $Y=434960
X444 1 2 ICV_3 $T=592480 388960 0 0 $X=592290 $Y=388720
X445 1 2 ICV_3 $T=595240 399840 0 0 $X=595050 $Y=399600
X446 1 2 ICV_3 $T=597540 405280 1 0 $X=597350 $Y=402320
X447 1 2 ICV_3 $T=604440 388960 1 0 $X=604250 $Y=386000
X448 1 2 ICV_3 $T=606740 443360 1 0 $X=606550 $Y=440400
X449 1 2 ICV_3 $T=609500 432480 1 0 $X=609310 $Y=429520
X450 1 2 ICV_3 $T=620540 421600 0 0 $X=620350 $Y=421360
X451 1 2 ICV_3 $T=623300 378080 0 0 $X=623110 $Y=377840
X452 1 2 ICV_3 $T=627440 421600 0 0 $X=627250 $Y=421360
X453 1 2 ICV_3 $T=637560 416160 1 0 $X=637370 $Y=413200
X454 1 2 ICV_3 $T=662860 388960 1 0 $X=662670 $Y=386000
X455 1 2 ICV_3 $T=662860 416160 1 0 $X=662670 $Y=413200
X456 1 2 ICV_3 $T=676660 410720 0 0 $X=676470 $Y=410480
X457 1 2 ICV_3 $T=676660 421600 0 0 $X=676470 $Y=421360
X458 1 2 ICV_3 $T=676660 437920 0 0 $X=676470 $Y=437680
X459 1 2 ICV_3 $T=683560 378080 0 0 $X=683370 $Y=377840
X460 1 2 ICV_3 $T=718980 394400 1 0 $X=718790 $Y=391440
X461 1 2 ICV_3 $T=732780 394400 0 0 $X=732590 $Y=394160
X462 1 2 ICV_3 $T=740600 388960 1 0 $X=740410 $Y=386000
X463 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=6900 394400 1 0 $X=6710 $Y=391440
X464 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=16560 388960 1 0 $X=16370 $Y=386000
X465 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=45080 394400 1 0 $X=44890 $Y=391440
X466 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=45080 432480 1 0 $X=44890 $Y=429520
X467 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=48300 443360 1 0 $X=48110 $Y=440400
X468 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=73140 410720 1 0 $X=72950 $Y=407760
X469 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=101200 410720 1 0 $X=101010 $Y=407760
X470 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=128800 427040 1 0 $X=128610 $Y=424080
X471 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=128800 443360 1 0 $X=128610 $Y=440400
X472 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=129260 405280 1 0 $X=129070 $Y=402320
X473 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=132480 443360 1 0 $X=132290 $Y=440400
X474 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=139840 399840 1 0 $X=139650 $Y=396880
X475 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=142600 378080 0 0 $X=142410 $Y=377840
X476 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=185380 432480 1 0 $X=185190 $Y=429520
X477 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=212980 399840 0 0 $X=212790 $Y=399600
X478 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=216660 388960 1 0 $X=216470 $Y=386000
X479 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=227240 378080 0 0 $X=227050 $Y=377840
X480 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=230460 416160 0 0 $X=230270 $Y=415920
X481 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=244720 399840 1 0 $X=244530 $Y=396880
X482 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=244720 405280 1 0 $X=244530 $Y=402320
X483 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=297160 443360 1 0 $X=296970 $Y=440400
X484 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=297620 405280 1 0 $X=297430 $Y=402320
X485 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=363860 405280 1 0 $X=363670 $Y=402320
X486 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=367540 427040 0 0 $X=367350 $Y=426800
X487 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=395140 427040 0 0 $X=394950 $Y=426800
X488 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=401580 432480 1 0 $X=401390 $Y=429520
X489 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=409860 405280 1 0 $X=409670 $Y=402320
X490 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=420440 437920 1 0 $X=420250 $Y=434960
X491 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=444360 421600 0 0 $X=444170 $Y=421360
X492 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=448500 410720 1 0 $X=448310 $Y=407760
X493 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=451260 410720 0 0 $X=451070 $Y=410480
X494 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=465520 443360 1 0 $X=465330 $Y=440400
X495 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=469200 383520 1 0 $X=469010 $Y=380560
X496 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=507380 410720 0 0 $X=507190 $Y=410480
X497 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=529460 383520 1 0 $X=529270 $Y=380560
X498 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=535900 388960 0 0 $X=535710 $Y=388720
X499 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=539120 399840 0 0 $X=538930 $Y=399600
X500 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=539120 405280 0 0 $X=538930 $Y=405040
X501 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=581440 437920 1 0 $X=581250 $Y=434960
X502 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=609500 383520 1 0 $X=609310 $Y=380560
X503 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=651820 416160 1 0 $X=651630 $Y=413200
X504 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=658720 410720 0 0 $X=658530 $Y=410480
X505 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=690000 416160 1 0 $X=689810 $Y=413200
X506 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=690000 437920 1 0 $X=689810 $Y=434960
X507 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=704260 437920 0 0 $X=704070 $Y=437680
X508 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=731860 399840 0 0 $X=731670 $Y=399600
X509 1 2 ICV_4 $T=6900 437920 0 0 $X=6710 $Y=437680
X510 1 2 ICV_4 $T=17020 394400 0 0 $X=16830 $Y=394160
X511 1 2 ICV_4 $T=20240 405280 0 0 $X=20050 $Y=405040
X512 1 2 ICV_4 $T=34040 437920 1 0 $X=33850 $Y=434960
X513 1 2 ICV_4 $T=36800 383520 1 0 $X=36610 $Y=380560
X514 1 2 ICV_4 $T=40020 388960 1 0 $X=39830 $Y=386000
X515 1 2 ICV_4 $T=97520 416160 0 0 $X=97330 $Y=415920
X516 1 2 ICV_4 $T=100740 443360 1 0 $X=100550 $Y=440400
X517 1 2 ICV_4 $T=104420 399840 1 0 $X=104230 $Y=396880
X518 1 2 ICV_4 $T=139840 405280 1 0 $X=139650 $Y=402320
X519 1 2 ICV_4 $T=188600 383520 1 0 $X=188410 $Y=380560
X520 1 2 ICV_4 $T=202400 394400 0 0 $X=202210 $Y=394160
X521 1 2 ICV_4 $T=212980 399840 1 0 $X=212790 $Y=396880
X522 1 2 ICV_4 $T=236900 405280 1 0 $X=236710 $Y=402320
X523 1 2 ICV_4 $T=262200 437920 1 0 $X=262010 $Y=434960
X524 1 2 ICV_4 $T=272780 388960 1 0 $X=272590 $Y=386000
X525 1 2 ICV_4 $T=272780 437920 1 0 $X=272590 $Y=434960
X526 1 2 ICV_4 $T=290720 421600 0 0 $X=290530 $Y=421360
X527 1 2 ICV_4 $T=302220 421600 0 0 $X=302030 $Y=421360
X528 1 2 ICV_4 $T=306820 421600 0 0 $X=306630 $Y=421360
X529 1 2 ICV_4 $T=310960 427040 0 0 $X=310770 $Y=426800
X530 1 2 ICV_4 $T=334880 399840 0 0 $X=334690 $Y=399600
X531 1 2 ICV_4 $T=382260 410720 0 0 $X=382070 $Y=410480
X532 1 2 ICV_4 $T=395140 394400 0 0 $X=394950 $Y=394160
X533 1 2 ICV_4 $T=410320 437920 0 0 $X=410130 $Y=437680
X534 1 2 ICV_4 $T=434700 421600 0 0 $X=434510 $Y=421360
X535 1 2 ICV_4 $T=441140 427040 1 0 $X=440950 $Y=424080
X536 1 2 ICV_4 $T=467820 427040 0 0 $X=467630 $Y=426800
X537 1 2 ICV_4 $T=539120 427040 0 0 $X=538930 $Y=426800
X538 1 2 ICV_4 $T=567180 388960 0 0 $X=566990 $Y=388720
X539 1 2 ICV_4 $T=581440 421600 1 0 $X=581250 $Y=418640
X540 1 2 ICV_4 $T=600760 427040 0 0 $X=600570 $Y=426800
X541 1 2 ICV_4 $T=633880 427040 1 0 $X=633690 $Y=424080
X542 1 2 ICV_4 $T=635720 437920 0 0 $X=635530 $Y=437680
X543 1 2 ICV_4 $T=657800 427040 0 0 $X=657610 $Y=426800
X544 1 2 ICV_4 $T=661940 443360 1 0 $X=661750 $Y=440400
X545 1 2 ICV_4 $T=721740 388960 1 0 $X=721550 $Y=386000
X546 1 2 ICV_4 $T=739680 378080 0 0 $X=739490 $Y=377840
X547 1 2 ICV_4 $T=739680 383520 0 0 $X=739490 $Y=383280
X548 1 2 ICV_4 $T=739680 388960 0 0 $X=739490 $Y=388720
X549 1 2 ICV_4 $T=739680 394400 0 0 $X=739490 $Y=394160
X550 1 2 ICV_4 $T=739680 399840 0 0 $X=739490 $Y=399600
X551 1 2 ICV_4 $T=739680 410720 1 0 $X=739490 $Y=407760
X552 1 2 ICV_4 $T=739680 432480 0 0 $X=739490 $Y=432240
X553 1 2 ICV_4 $T=739680 437920 1 0 $X=739490 $Y=434960
X554 1 2 ICV_4 $T=739680 443360 1 0 $X=739490 $Y=440400
X555 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 432480 0 0 $X=6710 $Y=432240
X556 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=15180 410720 0 0 $X=14990 $Y=410480
X557 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=22080 437920 0 0 $X=21890 $Y=437680
X558 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=26680 410720 1 0 $X=26490 $Y=407760
X559 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=29900 388960 0 0 $X=29710 $Y=388720
X560 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=29900 405280 0 0 $X=29710 $Y=405040
X561 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=44160 383520 1 0 $X=43970 $Y=380560
X562 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=66240 416160 0 0 $X=66050 $Y=415920
X563 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=71760 427040 0 0 $X=71570 $Y=426800
X564 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=84640 437920 0 0 $X=84450 $Y=437680
X565 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=101660 427040 0 0 $X=101470 $Y=426800
X566 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=106720 399840 0 0 $X=106530 $Y=399600
X567 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=108560 410720 1 0 $X=108370 $Y=407760
X568 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=118220 383520 0 0 $X=118030 $Y=383280
X569 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=139840 421600 1 0 $X=139650 $Y=418640
X570 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=146280 427040 1 0 $X=146090 $Y=424080
X571 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=146280 427040 0 0 $X=146090 $Y=426800
X572 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=156400 437920 1 0 $X=156210 $Y=434960
X573 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=172040 443360 1 0 $X=171850 $Y=440400
X574 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=186760 437920 0 0 $X=186570 $Y=437680
X575 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=193660 432480 0 0 $X=193470 $Y=432240
X576 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=194120 399840 0 0 $X=193930 $Y=399600
X577 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=196880 394400 1 0 $X=196690 $Y=391440
X578 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=216660 437920 0 0 $X=216470 $Y=437680
X579 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=224020 394400 1 0 $X=223830 $Y=391440
X580 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=272780 383520 1 0 $X=272590 $Y=380560
X581 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=272780 410720 1 0 $X=272590 $Y=407760
X582 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=275080 388960 0 0 $X=274890 $Y=388720
X583 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=277380 437920 1 0 $X=277190 $Y=434960
X584 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=284280 427040 1 0 $X=284090 $Y=424080
X585 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=310500 405280 1 0 $X=310310 $Y=402320
X586 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=314640 383520 0 0 $X=314450 $Y=383280
X587 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=315560 388960 1 0 $X=315370 $Y=386000
X588 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=316020 410720 1 0 $X=315830 $Y=407760
X589 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=322000 427040 0 0 $X=321810 $Y=426800
X590 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=324760 399840 1 0 $X=324570 $Y=396880
X591 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=326600 405280 0 0 $X=326410 $Y=405040
X592 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=336260 437920 1 0 $X=336070 $Y=434960
X593 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=348680 416160 1 0 $X=348490 $Y=413200
X594 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=355120 410720 0 0 $X=354930 $Y=410480
X595 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=364780 432480 1 0 $X=364590 $Y=429520
X596 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=379040 383520 0 0 $X=378850 $Y=383280
X597 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=387780 437920 0 0 $X=387590 $Y=437680
X598 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=393300 443360 1 0 $X=393110 $Y=440400
X599 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=397900 421600 1 0 $X=397710 $Y=418640
X600 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=408480 432480 1 0 $X=408290 $Y=429520
X601 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=437000 383520 1 0 $X=436810 $Y=380560
X602 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=457700 383520 1 0 $X=457510 $Y=380560
X603 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=460000 427040 1 0 $X=459810 $Y=424080
X604 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=463680 405280 0 0 $X=463490 $Y=405040
X605 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=467360 394400 0 0 $X=467170 $Y=394160
X606 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=473340 388960 1 0 $X=473150 $Y=386000
X607 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=484380 399840 0 0 $X=484190 $Y=399600
X608 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=515660 443360 1 0 $X=515470 $Y=440400
X609 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=525320 399840 0 0 $X=525130 $Y=399600
X610 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=525320 405280 1 0 $X=525130 $Y=402320
X611 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=533600 405280 0 0 $X=533410 $Y=405040
X612 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=533600 427040 0 0 $X=533410 $Y=426800
X613 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=534980 416160 0 0 $X=534790 $Y=415920
X614 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=547860 410720 1 0 $X=547670 $Y=407760
X615 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=548780 394400 1 0 $X=548590 $Y=391440
X616 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=553380 421600 1 0 $X=553190 $Y=418640
X617 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=558900 427040 0 0 $X=558710 $Y=426800
X618 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=569020 421600 1 0 $X=568830 $Y=418640
X619 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=581900 410720 0 0 $X=581710 $Y=410480
X620 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=586500 383520 1 0 $X=586310 $Y=380560
X621 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=588340 437920 1 0 $X=588150 $Y=434960
X622 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=596160 427040 1 0 $X=595970 $Y=424080
X623 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=619160 432480 0 0 $X=618970 $Y=432240
X624 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=623300 388960 0 0 $X=623110 $Y=388720
X625 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=635720 416160 0 0 $X=635530 $Y=415920
X626 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=647220 437920 0 0 $X=647030 $Y=437680
X627 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=658720 378080 0 0 $X=658530 $Y=377840
X628 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=697820 443360 1 0 $X=697630 $Y=440400
X629 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=707480 416160 1 0 $X=707290 $Y=413200
X630 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=718980 432480 0 0 $X=718790 $Y=432240
X631 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=720820 383520 0 0 $X=720630 $Y=383280
X632 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=721740 383520 1 0 $X=721550 $Y=380560
X633 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=731400 378080 0 0 $X=731210 $Y=377840
X634 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=738760 405280 1 0 $X=738570 $Y=402320
X635 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=738760 427040 1 0 $X=738570 $Y=424080
X636 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=739220 421600 1 0 $X=739030 $Y=418640
X637 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=16560 437920 0 0 $X=16370 $Y=437680
X638 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=76360 416160 1 0 $X=76170 $Y=413200
X639 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=125580 399840 0 0 $X=125390 $Y=399600
X640 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=146280 405280 0 0 $X=146090 $Y=405040
X641 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=228160 421600 1 0 $X=227970 $Y=418640
X642 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=291180 399840 0 0 $X=290990 $Y=399600
X643 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=378580 399840 1 0 $X=378390 $Y=396880
X644 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=435160 432480 1 0 $X=434970 $Y=429520
X645 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=559820 405280 1 0 $X=559630 $Y=402320
X646 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=560280 416160 0 0 $X=560090 $Y=415920
X647 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=561200 410720 0 0 $X=561010 $Y=410480
X648 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=665160 427040 0 0 $X=664970 $Y=426800
X649 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=730020 416160 1 0 $X=729830 $Y=413200
X650 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=733240 405280 1 0 $X=733050 $Y=402320
X651 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=733240 427040 1 0 $X=733050 $Y=424080
X652 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=733700 421600 1 0 $X=733510 $Y=418640
X653 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=734160 410720 1 0 $X=733970 $Y=407760
X654 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=734160 437920 1 0 $X=733970 $Y=434960
X655 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=734160 443360 1 0 $X=733970 $Y=440400
X656 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 405280 0 0 $X=735350 $Y=405040
X657 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 410720 0 0 $X=735350 $Y=410480
X658 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 416160 1 0 $X=735350 $Y=413200
X659 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 416160 0 0 $X=735350 $Y=415920
X660 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 421600 0 0 $X=735350 $Y=421360
X661 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 427040 0 0 $X=735350 $Y=426800
X662 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 437920 0 0 $X=735350 $Y=437680
X663 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=736460 399840 1 0 $X=736270 $Y=396880
X664 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=737380 432480 1 0 $X=737190 $Y=429520
X665 1 2 4 2 14 1 sky130_fd_sc_hd__clkbuf_8 $T=6900 399840 1 0 $X=6710 $Y=396880
X666 1 2 19 2 27 1 sky130_fd_sc_hd__clkbuf_8 $T=14720 427040 1 0 $X=14530 $Y=424080
X667 1 2 535 534 2 23 1 sky130_fd_sc_hd__ebufn_2 $T=16100 416160 0 0 $X=15910 $Y=415920
X668 1 2 573 580 2 36 1 sky130_fd_sc_hd__ebufn_2 $T=40020 383520 1 0 $X=39830 $Y=380560
X669 1 2 586 554 2 34 1 sky130_fd_sc_hd__ebufn_2 $T=41400 427040 0 0 $X=41210 $Y=426800
X670 1 2 584 576 2 16 1 sky130_fd_sc_hd__ebufn_2 $T=42320 421600 1 0 $X=42130 $Y=418640
X671 1 2 44 45 2 34 1 sky130_fd_sc_hd__ebufn_2 $T=43240 378080 0 0 $X=43050 $Y=377840
X672 1 2 589 580 2 23 1 sky130_fd_sc_hd__ebufn_2 $T=43240 388960 1 0 $X=43050 $Y=386000
X673 1 2 572 576 2 24 1 sky130_fd_sc_hd__ebufn_2 $T=43240 410720 1 0 $X=43050 $Y=407760
X674 1 2 603 605 2 31 1 sky130_fd_sc_hd__ebufn_2 $T=51060 405280 1 0 $X=50870 $Y=402320
X675 1 2 607 51 2 36 1 sky130_fd_sc_hd__ebufn_2 $T=62100 378080 0 0 $X=61910 $Y=377840
X676 1 2 671 644 2 24 1 sky130_fd_sc_hd__ebufn_2 $T=83260 421600 0 0 $X=83070 $Y=421360
X677 1 2 688 634 2 23 1 sky130_fd_sc_hd__ebufn_2 $T=92460 394400 0 0 $X=92270 $Y=394160
X678 1 2 715 716 2 23 1 sky130_fd_sc_hd__ebufn_2 $T=107640 399840 1 0 $X=107450 $Y=396880
X679 1 2 777 768 2 16 1 sky130_fd_sc_hd__ebufn_2 $T=138460 437920 1 0 $X=138270 $Y=434960
X680 1 2 812 120 2 118 1 sky130_fd_sc_hd__ebufn_2 $T=155480 437920 0 0 $X=155290 $Y=437680
X681 1 2 871 854 2 118 1 sky130_fd_sc_hd__ebufn_2 $T=184000 405280 0 0 $X=183810 $Y=405040
X682 1 2 862 844 2 129 1 sky130_fd_sc_hd__ebufn_2 $T=185840 427040 0 0 $X=185650 $Y=426800
X683 1 2 883 888 2 131 1 sky130_fd_sc_hd__ebufn_2 $T=196880 383520 1 0 $X=196690 $Y=380560
X684 1 2 894 140 2 131 1 sky130_fd_sc_hd__ebufn_2 $T=197340 432480 0 0 $X=197150 $Y=432240
X685 1 2 896 873 2 118 1 sky130_fd_sc_hd__ebufn_2 $T=198260 405280 1 0 $X=198070 $Y=402320
X686 1 2 892 845 2 119 1 sky130_fd_sc_hd__ebufn_2 $T=201940 410720 1 0 $X=201750 $Y=407760
X687 1 2 903 873 2 128 1 sky130_fd_sc_hd__ebufn_2 $T=205620 394400 0 0 $X=205430 $Y=394160
X688 1 2 893 845 2 118 1 sky130_fd_sc_hd__ebufn_2 $T=213900 410720 0 0 $X=213710 $Y=410480
X689 1 2 947 918 2 122 1 sky130_fd_sc_hd__ebufn_2 $T=224020 405280 1 0 $X=223830 $Y=402320
X690 1 2 948 949 2 130 1 sky130_fd_sc_hd__ebufn_2 $T=224020 421600 1 0 $X=223830 $Y=418640
X691 1 2 998 976 2 122 1 sky130_fd_sc_hd__ebufn_2 $T=252080 427040 0 0 $X=251890 $Y=426800
X692 1 2 1002 1008 2 129 1 sky130_fd_sc_hd__ebufn_2 $T=252540 399840 1 0 $X=252350 $Y=396880
X693 1 2 993 1008 2 118 1 sky130_fd_sc_hd__ebufn_2 $T=256680 394400 1 0 $X=256490 $Y=391440
X694 1 2 1030 162 2 129 1 sky130_fd_sc_hd__ebufn_2 $T=265420 437920 1 0 $X=265230 $Y=434960
X695 1 2 1044 1019 2 129 1 sky130_fd_sc_hd__ebufn_2 $T=271860 427040 0 0 $X=271670 $Y=426800
X696 1 2 1064 1067 2 130 1 sky130_fd_sc_hd__ebufn_2 $T=283360 437920 1 0 $X=283170 $Y=434960
X697 1 2 1071 1053 2 118 1 sky130_fd_sc_hd__ebufn_2 $T=286580 399840 1 0 $X=286390 $Y=396880
X698 1 2 1069 1067 2 129 1 sky130_fd_sc_hd__ebufn_2 $T=286580 421600 0 0 $X=286390 $Y=421360
X699 1 2 1075 1053 2 129 1 sky130_fd_sc_hd__ebufn_2 $T=287960 394400 0 0 $X=287770 $Y=394160
X700 1 2 1085 1067 2 131 1 sky130_fd_sc_hd__ebufn_2 $T=293940 432480 1 0 $X=293750 $Y=429520
X701 1 2 1094 1097 2 130 1 sky130_fd_sc_hd__ebufn_2 $T=296240 410720 1 0 $X=296050 $Y=407760
X702 1 2 1099 1097 2 128 1 sky130_fd_sc_hd__ebufn_2 $T=298080 399840 0 0 $X=297890 $Y=399600
X703 1 2 1122 1107 2 130 1 sky130_fd_sc_hd__ebufn_2 $T=310040 421600 0 0 $X=309850 $Y=421360
X704 1 2 1114 1097 2 129 1 sky130_fd_sc_hd__ebufn_2 $T=314640 405280 0 0 $X=314450 $Y=405040
X705 1 2 1139 1102 2 130 1 sky130_fd_sc_hd__ebufn_2 $T=324300 432480 1 0 $X=324110 $Y=429520
X706 1 2 1157 1144 2 230 1 sky130_fd_sc_hd__ebufn_2 $T=333500 388960 1 0 $X=333310 $Y=386000
X707 1 2 1166 1168 2 221 1 sky130_fd_sc_hd__ebufn_2 $T=337640 399840 1 0 $X=337450 $Y=396880
X708 1 2 1224 1225 2 205 1 sky130_fd_sc_hd__ebufn_2 $T=366620 405280 1 0 $X=366430 $Y=402320
X709 1 2 1227 1223 2 180 1 sky130_fd_sc_hd__ebufn_2 $T=368460 432480 1 0 $X=368270 $Y=429520
X710 1 2 1253 1225 2 222 1 sky130_fd_sc_hd__ebufn_2 $T=379960 388960 0 0 $X=379770 $Y=388720
X711 1 2 1293 264 2 220 1 sky130_fd_sc_hd__ebufn_2 $T=404340 432480 1 0 $X=404150 $Y=429520
X712 1 2 1295 1290 2 222 1 sky130_fd_sc_hd__ebufn_2 $T=408480 394400 1 0 $X=408290 $Y=391440
X713 1 2 1303 1305 2 192 1 sky130_fd_sc_hd__ebufn_2 $T=408480 421600 1 0 $X=408290 $Y=418640
X714 1 2 1309 276 2 192 1 sky130_fd_sc_hd__ebufn_2 $T=413540 437920 0 0 $X=413350 $Y=437680
X715 1 2 1315 1317 2 230 1 sky130_fd_sc_hd__ebufn_2 $T=414920 383520 0 0 $X=414730 $Y=383280
X716 1 2 1324 1317 2 221 1 sky130_fd_sc_hd__ebufn_2 $T=419060 405280 0 0 $X=418870 $Y=405040
X717 1 2 1310 1305 2 239 1 sky130_fd_sc_hd__ebufn_2 $T=423200 427040 1 0 $X=423010 $Y=424080
X718 1 2 1382 295 2 222 1 sky130_fd_sc_hd__ebufn_2 $T=448040 388960 0 0 $X=447850 $Y=388720
X719 1 2 1392 1380 2 180 1 sky130_fd_sc_hd__ebufn_2 $T=454940 410720 0 0 $X=454750 $Y=410480
X720 1 2 1419 1403 2 187 1 sky130_fd_sc_hd__ebufn_2 $T=469200 410720 1 0 $X=469010 $Y=407760
X721 1 2 1437 1443 2 222 1 sky130_fd_sc_hd__ebufn_2 $T=477940 388960 0 0 $X=477750 $Y=388720
X722 1 2 1446 1447 2 220 1 sky130_fd_sc_hd__ebufn_2 $T=481160 410720 1 0 $X=480970 $Y=407760
X723 1 2 1468 326 2 206 1 sky130_fd_sc_hd__ebufn_2 $T=497260 383520 1 0 $X=497070 $Y=380560
X724 1 2 1485 1487 2 192 1 sky130_fd_sc_hd__ebufn_2 $T=500020 421600 0 0 $X=499830 $Y=421360
X725 1 2 1497 336 2 239 1 sky130_fd_sc_hd__ebufn_2 $T=506460 432480 1 0 $X=506270 $Y=429520
X726 1 2 1499 336 2 220 1 sky130_fd_sc_hd__ebufn_2 $T=511520 443360 1 0 $X=511330 $Y=440400
X727 1 2 1509 1480 2 187 1 sky130_fd_sc_hd__ebufn_2 $T=525320 410720 0 0 $X=525130 $Y=410480
X728 1 2 1555 1545 2 343 1 sky130_fd_sc_hd__ebufn_2 $T=555220 416160 1 0 $X=555030 $Y=413200
X729 1 2 1593 1589 2 355 1 sky130_fd_sc_hd__ebufn_2 $T=573160 427040 0 0 $X=572970 $Y=426800
X730 1 2 1613 1586 2 388 1 sky130_fd_sc_hd__ebufn_2 $T=583280 399840 1 0 $X=583090 $Y=396880
X731 1 2 1615 1589 2 368 1 sky130_fd_sc_hd__ebufn_2 $T=584200 437920 1 0 $X=584010 $Y=434960
X732 1 2 1639 1637 2 363 1 sky130_fd_sc_hd__ebufn_2 $T=596620 405280 0 0 $X=596430 $Y=405040
X733 1 2 1640 1638 2 368 1 sky130_fd_sc_hd__ebufn_2 $T=596620 427040 0 0 $X=596430 $Y=426800
X734 1 2 1684 1643 2 371 1 sky130_fd_sc_hd__ebufn_2 $T=631580 437920 0 0 $X=631390 $Y=437680
X735 1 2 1714 1690 2 363 1 sky130_fd_sc_hd__ebufn_2 $T=632500 427040 0 0 $X=632310 $Y=426800
X736 1 2 1724 1689 2 363 1 sky130_fd_sc_hd__ebufn_2 $T=639860 416160 1 0 $X=639670 $Y=413200
X737 1 2 1746 1754 2 371 1 sky130_fd_sc_hd__ebufn_2 $T=653200 416160 0 0 $X=653010 $Y=415920
X738 1 2 1745 1754 2 366 1 sky130_fd_sc_hd__ebufn_2 $T=657800 410720 1 0 $X=657610 $Y=407760
X739 1 2 1762 440 2 355 1 sky130_fd_sc_hd__ebufn_2 $T=657800 443360 1 0 $X=657610 $Y=440400
X740 1 2 1763 439 2 397 1 sky130_fd_sc_hd__ebufn_2 $T=658720 388960 1 0 $X=658530 $Y=386000
X741 1 2 1768 440 2 363 1 sky130_fd_sc_hd__ebufn_2 $T=661020 427040 0 0 $X=660830 $Y=426800
X742 1 2 1796 447 2 391 1 sky130_fd_sc_hd__ebufn_2 $T=674820 388960 0 0 $X=674630 $Y=388720
X743 1 2 1807 447 2 352 1 sky130_fd_sc_hd__ebufn_2 $T=684020 394400 0 0 $X=683830 $Y=394160
X744 1 2 1817 447 2 397 1 sky130_fd_sc_hd__ebufn_2 $T=688620 399840 1 0 $X=688430 $Y=396880
X745 1 2 1845 1851 2 392 1 sky130_fd_sc_hd__ebufn_2 $T=706100 388960 1 0 $X=705910 $Y=386000
X746 1 2 1835 1842 2 345 1 sky130_fd_sc_hd__ebufn_2 $T=707480 399840 0 0 $X=707290 $Y=399600
X747 1 2 1908 1885 2 386 1 sky130_fd_sc_hd__ebufn_2 $T=735540 383520 0 0 $X=735350 $Y=383280
X748 1 2 1909 1885 2 387 1 sky130_fd_sc_hd__ebufn_2 $T=735540 388960 0 0 $X=735350 $Y=388720
X749 1 2 1911 1865 2 388 1 sky130_fd_sc_hd__ebufn_2 $T=735540 399840 0 0 $X=735350 $Y=399600
X875 1 2 529 534 24 ICV_6 $T=19780 410720 1 0 $X=19590 $Y=407760
X876 1 2 568 554 36 ICV_6 $T=33580 421600 0 0 $X=33390 $Y=421360
X877 1 2 559 533 36 ICV_6 $T=33580 432480 0 0 $X=33390 $Y=432240
X878 1 2 629 51 34 ICV_6 $T=61640 383520 0 0 $X=61450 $Y=383280
X879 1 2 627 615 31 ICV_6 $T=61640 410720 0 0 $X=61450 $Y=410480
X880 1 2 620 615 23 ICV_6 $T=61640 416160 0 0 $X=61450 $Y=415920
X881 1 2 618 52 25 ICV_6 $T=61640 432480 0 0 $X=61450 $Y=432240
X882 1 2 619 52 23 ICV_6 $T=61640 437920 0 0 $X=61450 $Y=437680
X883 1 2 682 683 16 ICV_6 $T=89700 410720 0 0 $X=89510 $Y=410480
X884 1 2 704 683 31 ICV_6 $T=103960 410720 1 0 $X=103770 $Y=407760
X885 1 2 778 758 37 ICV_6 $T=145820 399840 0 0 $X=145630 $Y=399600
X886 1 2 804 802 118 ICV_6 $T=160080 394400 1 0 $X=159890 $Y=391440
X887 1 2 828 798 131 ICV_6 $T=173880 394400 0 0 $X=173690 $Y=394160
X888 1 2 1031 1008 130 ICV_6 $T=272320 399840 1 0 $X=272130 $Y=396880
X889 1 2 1034 1019 130 ICV_6 $T=272320 432480 1 0 $X=272130 $Y=429520
X890 1 2 1170 1152 180 ICV_6 $T=342240 416160 0 0 $X=342050 $Y=415920
X891 1 2 1187 1168 222 ICV_6 $T=356500 399840 1 0 $X=356310 $Y=396880
X892 1 2 1228 1207 236 ICV_6 $T=370300 378080 0 0 $X=370110 $Y=377840
X893 1 2 1280 1223 220 ICV_6 $T=398360 421600 0 0 $X=398170 $Y=421360
X894 1 2 1297 1290 221 ICV_6 $T=412620 394400 1 0 $X=412430 $Y=391440
X895 1 2 1312 1305 195 ICV_6 $T=412620 416160 1 0 $X=412430 $Y=413200
X896 1 2 1345 282 221 ICV_6 $T=440680 399840 1 0 $X=440490 $Y=396880
X897 1 2 1397 1380 187 ICV_6 $T=454480 416160 0 0 $X=454290 $Y=415920
X898 1 2 1417 1399 222 ICV_6 $T=468740 388960 1 0 $X=468550 $Y=386000
X899 1 2 321 307 180 ICV_6 $T=482540 432480 0 0 $X=482350 $Y=432240
X900 1 2 1481 323 206 ICV_6 $T=496800 399840 1 0 $X=496610 $Y=396880
X901 1 2 1477 322 239 ICV_6 $T=496800 437920 1 0 $X=496610 $Y=434960
X902 1 2 1500 326 236 ICV_6 $T=510600 378080 0 0 $X=510410 $Y=377840
X903 1 2 1498 1487 220 ICV_6 $T=510600 421600 0 0 $X=510410 $Y=421360
X904 1 2 1582 1553 388 ICV_6 $T=566720 399840 0 0 $X=566530 $Y=399600
X905 1 2 1576 1545 368 ICV_6 $T=566720 416160 0 0 $X=566530 $Y=415920
X906 1 2 1578 1550 368 ICV_6 $T=566720 421600 0 0 $X=566530 $Y=421360
X907 1 2 1606 1597 363 ICV_6 $T=580980 410720 1 0 $X=580790 $Y=407760
X908 1 2 1604 1597 343 ICV_6 $T=580980 427040 1 0 $X=580790 $Y=424080
X909 1 2 1661 1638 367 ICV_6 $T=609040 427040 1 0 $X=608850 $Y=424080
X910 1 2 1681 1655 386 ICV_6 $T=622840 399840 0 0 $X=622650 $Y=399600
X911 1 2 1692 1690 345 ICV_6 $T=622840 421600 0 0 $X=622650 $Y=421360
X912 1 2 1758 440 368 ICV_6 $T=665160 437920 1 0 $X=664970 $Y=434960
X913 1 2 1798 448 397 ICV_6 $T=678960 378080 0 0 $X=678770 $Y=377840
X914 1 2 458 455 371 ICV_6 $T=693220 443360 1 0 $X=693030 $Y=440400
X915 1 2 1889 464 389 ICV_6 $T=735080 378080 0 0 $X=734890 $Y=377840
X916 1 2 1910 1865 387 ICV_6 $T=735080 394400 0 0 $X=734890 $Y=394160
X917 1 2 1903 1874 366 ICV_6 $T=735080 432480 0 0 $X=734890 $Y=432240
X1047 1 2 517 9 2 536 1 sky130_fd_sc_hd__dfxtp_1 $T=9200 383520 0 0 $X=9010 $Y=383280
X1048 1 2 514 28 2 553 1 sky130_fd_sc_hd__dfxtp_1 $T=18860 432480 0 0 $X=18670 $Y=432240
X1049 1 2 555 9 2 552 1 sky130_fd_sc_hd__dfxtp_1 $T=26220 432480 0 0 $X=26030 $Y=432240
X1050 1 2 564 28 2 596 1 sky130_fd_sc_hd__dfxtp_1 $T=40020 416160 1 0 $X=39830 $Y=413200
X1051 1 2 604 29 2 622 1 sky130_fd_sc_hd__dfxtp_1 $T=51980 427040 0 0 $X=51790 $Y=426800
X1052 1 2 597 28 2 629 1 sky130_fd_sc_hd__dfxtp_1 $T=55660 388960 1 0 $X=55470 $Y=386000
X1053 1 2 637 17 2 654 1 sky130_fd_sc_hd__dfxtp_1 $T=68080 394400 1 0 $X=67890 $Y=391440
X1054 1 2 635 30 2 655 1 sky130_fd_sc_hd__dfxtp_1 $T=68080 399840 0 0 $X=67890 $Y=399600
X1055 1 2 637 9 2 633 1 sky130_fd_sc_hd__dfxtp_1 $T=68540 394400 0 0 $X=68350 $Y=394160
X1056 1 2 664 28 2 684 1 sky130_fd_sc_hd__dfxtp_1 $T=84640 388960 1 0 $X=84450 $Y=386000
X1057 1 2 64 29 2 693 1 sky130_fd_sc_hd__dfxtp_1 $T=87400 437920 1 0 $X=87210 $Y=434960
X1058 1 2 664 30 2 733 1 sky130_fd_sc_hd__dfxtp_1 $T=107180 388960 0 0 $X=106990 $Y=388720
X1059 1 2 712 10 2 718 1 sky130_fd_sc_hd__dfxtp_1 $T=108560 416160 0 0 $X=108370 $Y=415920
X1060 1 2 711 11 2 755 1 sky130_fd_sc_hd__dfxtp_1 $T=120060 421600 0 0 $X=119870 $Y=421360
X1061 1 2 794 109 2 808 1 sky130_fd_sc_hd__dfxtp_1 $T=149040 399840 1 0 $X=148850 $Y=396880
X1062 1 2 108 109 2 812 1 sky130_fd_sc_hd__dfxtp_1 $T=149040 437920 1 0 $X=148850 $Y=434960
X1063 1 2 795 113 2 815 1 sky130_fd_sc_hd__dfxtp_1 $T=149960 421600 1 0 $X=149770 $Y=418640
X1064 1 2 795 112 2 817 1 sky130_fd_sc_hd__dfxtp_1 $T=149960 427040 0 0 $X=149770 $Y=426800
X1065 1 2 794 113 2 818 1 sky130_fd_sc_hd__dfxtp_1 $T=150420 399840 0 0 $X=150230 $Y=399600
X1066 1 2 794 112 2 797 1 sky130_fd_sc_hd__dfxtp_1 $T=152260 405280 1 0 $X=152070 $Y=402320
X1067 1 2 121 111 2 821 1 sky130_fd_sc_hd__dfxtp_1 $T=158240 383520 0 0 $X=158050 $Y=383280
X1068 1 2 793 127 2 851 1 sky130_fd_sc_hd__dfxtp_1 $T=172040 388960 1 0 $X=171850 $Y=386000
X1069 1 2 846 124 2 847 1 sky130_fd_sc_hd__dfxtp_1 $T=176180 410720 1 0 $X=175990 $Y=407760
X1070 1 2 855 127 2 869 1 sky130_fd_sc_hd__dfxtp_1 $T=180780 394400 0 0 $X=180590 $Y=394160
X1071 1 2 846 127 2 877 1 sky130_fd_sc_hd__dfxtp_1 $T=182620 410720 0 0 $X=182430 $Y=410480
X1072 1 2 135 109 2 142 1 sky130_fd_sc_hd__dfxtp_1 $T=192280 378080 0 0 $X=192090 $Y=377840
X1073 1 2 855 124 2 903 1 sky130_fd_sc_hd__dfxtp_1 $T=198260 399840 1 0 $X=198070 $Y=396880
X1074 1 2 874 113 2 905 1 sky130_fd_sc_hd__dfxtp_1 $T=200560 394400 1 0 $X=200370 $Y=391440
X1075 1 2 855 111 2 924 1 sky130_fd_sc_hd__dfxtp_1 $T=205620 399840 1 0 $X=205430 $Y=396880
X1076 1 2 931 112 2 154 1 sky130_fd_sc_hd__dfxtp_1 $T=231380 443360 1 0 $X=231190 $Y=440400
X1077 1 2 965 111 2 975 1 sky130_fd_sc_hd__dfxtp_1 $T=233220 410720 1 0 $X=233030 $Y=407760
X1078 1 2 926 113 2 960 1 sky130_fd_sc_hd__dfxtp_1 $T=233680 399840 1 0 $X=233490 $Y=396880
X1079 1 2 1014 124 2 1027 1 sky130_fd_sc_hd__dfxtp_1 $T=258520 421600 1 0 $X=258330 $Y=418640
X1080 1 2 169 127 2 170 1 sky130_fd_sc_hd__dfxtp_1 $T=276460 383520 1 0 $X=276270 $Y=380560
X1081 1 2 160 112 2 1047 1 sky130_fd_sc_hd__dfxtp_1 $T=276460 383520 0 0 $X=276270 $Y=383280
X1082 1 2 1050 124 2 1070 1 sky130_fd_sc_hd__dfxtp_1 $T=278300 432480 0 0 $X=278110 $Y=432240
X1083 1 2 1066 109 2 1100 1 sky130_fd_sc_hd__dfxtp_1 $T=291640 421600 1 0 $X=291450 $Y=418640
X1084 1 2 1072 109 2 1116 1 sky130_fd_sc_hd__dfxtp_1 $T=303140 388960 0 0 $X=302950 $Y=388720
X1085 1 2 1104 125 2 1123 1 sky130_fd_sc_hd__dfxtp_1 $T=303600 427040 0 0 $X=303410 $Y=426800
X1086 1 2 1129 191 2 1145 1 sky130_fd_sc_hd__dfxtp_1 $T=319240 388960 1 0 $X=319050 $Y=386000
X1087 1 2 1128 191 2 1149 1 sky130_fd_sc_hd__dfxtp_1 $T=322460 394400 0 0 $X=322270 $Y=394160
X1088 1 2 1129 219 2 1175 1 sky130_fd_sc_hd__dfxtp_1 $T=334880 378080 0 0 $X=334690 $Y=377840
X1089 1 2 1167 190 2 1178 1 sky130_fd_sc_hd__dfxtp_1 $T=338100 405280 1 0 $X=337910 $Y=402320
X1090 1 2 1173 224 2 1186 1 sky130_fd_sc_hd__dfxtp_1 $T=341320 416160 1 0 $X=341130 $Y=413200
X1091 1 2 1173 199 2 1193 1 sky130_fd_sc_hd__dfxtp_1 $T=346840 416160 0 0 $X=346650 $Y=415920
X1092 1 2 1173 227 2 1190 1 sky130_fd_sc_hd__dfxtp_1 $T=349140 410720 1 0 $X=348950 $Y=407760
X1093 1 2 1185 196 2 1205 1 sky130_fd_sc_hd__dfxtp_1 $T=350520 421600 0 0 $X=350330 $Y=421360
X1094 1 2 241 212 2 1238 1 sky130_fd_sc_hd__dfxtp_1 $T=366160 388960 1 0 $X=365970 $Y=386000
X1095 1 2 1210 184 2 1253 1 sky130_fd_sc_hd__dfxtp_1 $T=373520 388960 1 0 $X=373330 $Y=386000
X1096 1 2 248 228 2 1251 1 sky130_fd_sc_hd__dfxtp_1 $T=373520 437920 1 0 $X=373330 $Y=434960
X1097 1 2 248 204 2 1252 1 sky130_fd_sc_hd__dfxtp_1 $T=373520 443360 1 0 $X=373330 $Y=440400
X1098 1 2 1211 227 2 1237 1 sky130_fd_sc_hd__dfxtp_1 $T=374900 410720 1 0 $X=374710 $Y=407760
X1099 1 2 268 189 2 269 1 sky130_fd_sc_hd__dfxtp_1 $T=396060 383520 1 0 $X=395870 $Y=380560
X1100 1 2 258 228 2 271 1 sky130_fd_sc_hd__dfxtp_1 $T=396980 443360 1 0 $X=396790 $Y=440400
X1101 1 2 1259 228 2 1284 1 sky130_fd_sc_hd__dfxtp_1 $T=400660 410720 1 0 $X=400470 $Y=407760
X1102 1 2 1282 189 2 1307 1 sky130_fd_sc_hd__dfxtp_1 $T=404800 388960 1 0 $X=404610 $Y=386000
X1103 1 2 1286 228 2 1303 1 sky130_fd_sc_hd__dfxtp_1 $T=413540 416160 0 0 $X=413350 $Y=415920
X1104 1 2 277 219 2 1332 1 sky130_fd_sc_hd__dfxtp_1 $T=415380 388960 0 0 $X=415190 $Y=388720
X1105 1 2 1321 227 2 1333 1 sky130_fd_sc_hd__dfxtp_1 $T=417220 416160 1 0 $X=417030 $Y=413200
X1106 1 2 1300 185 2 1339 1 sky130_fd_sc_hd__dfxtp_1 $T=418600 399840 0 0 $X=418410 $Y=399600
X1107 1 2 1340 185 2 1356 1 sky130_fd_sc_hd__dfxtp_1 $T=428260 399840 0 0 $X=428070 $Y=399600
X1108 1 2 277 185 2 1360 1 sky130_fd_sc_hd__dfxtp_1 $T=429640 383520 1 0 $X=429450 $Y=380560
X1109 1 2 277 189 2 1363 1 sky130_fd_sc_hd__dfxtp_1 $T=431480 388960 1 0 $X=431290 $Y=386000
X1110 1 2 1364 204 2 1375 1 sky130_fd_sc_hd__dfxtp_1 $T=438380 416160 0 0 $X=438190 $Y=415920
X1111 1 2 298 196 2 1409 1 sky130_fd_sc_hd__dfxtp_1 $T=455400 437920 1 0 $X=455210 $Y=434960
X1112 1 2 1377 219 2 1415 1 sky130_fd_sc_hd__dfxtp_1 $T=460920 399840 0 0 $X=460730 $Y=399600
X1113 1 2 1408 190 2 1445 1 sky130_fd_sc_hd__dfxtp_1 $T=474260 378080 0 0 $X=474070 $Y=377840
X1114 1 2 319 196 2 1454 1 sky130_fd_sc_hd__dfxtp_1 $T=477940 437920 1 0 $X=477750 $Y=434960
X1115 1 2 1456 191 2 1452 1 sky130_fd_sc_hd__dfxtp_1 $T=487140 388960 1 0 $X=486950 $Y=386000
X1116 1 2 1470 213 2 1498 1 sky130_fd_sc_hd__dfxtp_1 $T=500480 427040 0 0 $X=500290 $Y=426800
X1117 1 2 1519 359 2 1528 1 sky130_fd_sc_hd__dfxtp_1 $T=526240 427040 0 0 $X=526050 $Y=426800
X1118 1 2 179 371 2 382 1 sky130_fd_sc_hd__dfxtp_1 $T=534060 410720 1 0 $X=533870 $Y=407760
X1119 1 2 1539 357 2 1551 1 sky130_fd_sc_hd__dfxtp_1 $T=547860 405280 0 0 $X=547670 $Y=405040
X1120 1 2 1587 403 2 1599 1 sky130_fd_sc_hd__dfxtp_1 $T=571780 394400 1 0 $X=571590 $Y=391440
X1121 1 2 1587 402 2 1601 1 sky130_fd_sc_hd__dfxtp_1 $T=572240 399840 1 0 $X=572050 $Y=396880
X1122 1 2 1585 381 2 1602 1 sky130_fd_sc_hd__dfxtp_1 $T=572240 410720 1 0 $X=572050 $Y=407760
X1123 1 2 1585 358 2 1603 1 sky130_fd_sc_hd__dfxtp_1 $T=572700 421600 1 0 $X=572510 $Y=418640
X1124 1 2 1585 365 2 1606 1 sky130_fd_sc_hd__dfxtp_1 $T=573160 405280 0 0 $X=572970 $Y=405040
X1125 1 2 1618 358 2 1627 1 sky130_fd_sc_hd__dfxtp_1 $T=585580 410720 1 0 $X=585390 $Y=407760
X1126 1 2 1618 378 2 1628 1 sky130_fd_sc_hd__dfxtp_1 $T=585580 410720 0 0 $X=585390 $Y=410480
X1127 1 2 1587 395 2 1629 1 sky130_fd_sc_hd__dfxtp_1 $T=586040 399840 0 0 $X=585850 $Y=399600
X1128 1 2 1592 406 2 1631 1 sky130_fd_sc_hd__dfxtp_1 $T=586960 383520 0 0 $X=586770 $Y=383280
X1129 1 2 1621 357 2 1661 1 sky130_fd_sc_hd__dfxtp_1 $T=599840 427040 1 0 $X=599650 $Y=424080
X1130 1 2 1641 402 2 1665 1 sky130_fd_sc_hd__dfxtp_1 $T=601680 399840 1 0 $X=601490 $Y=396880
X1131 1 2 421 402 2 1674 1 sky130_fd_sc_hd__dfxtp_1 $T=605820 383520 0 0 $X=605630 $Y=383280
X1132 1 2 1671 360 2 1682 1 sky130_fd_sc_hd__dfxtp_1 $T=611800 432480 0 0 $X=611610 $Y=432240
X1133 1 2 418 381 2 1701 1 sky130_fd_sc_hd__dfxtp_1 $T=619160 443360 1 0 $X=618970 $Y=440400
X1134 1 2 1685 395 2 1709 1 sky130_fd_sc_hd__dfxtp_1 $T=623760 399840 1 0 $X=623570 $Y=396880
X1135 1 2 1685 393 2 1712 1 sky130_fd_sc_hd__dfxtp_1 $T=624680 405280 1 0 $X=624490 $Y=402320
X1136 1 2 1671 365 2 1714 1 sky130_fd_sc_hd__dfxtp_1 $T=626520 427040 1 0 $X=626330 $Y=424080
X1137 1 2 1685 406 2 1718 1 sky130_fd_sc_hd__dfxtp_1 $T=628360 388960 1 0 $X=628170 $Y=386000
X1138 1 2 1721 407 2 1727 1 sky130_fd_sc_hd__dfxtp_1 $T=641240 383520 0 0 $X=641050 $Y=383280
X1139 1 2 1751 358 2 1766 1 sky130_fd_sc_hd__dfxtp_1 $T=653660 421600 0 0 $X=653470 $Y=421360
X1140 1 2 1747 381 2 441 1 sky130_fd_sc_hd__dfxtp_1 $T=657800 437920 1 0 $X=657610 $Y=434960
X1141 1 2 1751 372 2 1792 1 sky130_fd_sc_hd__dfxtp_1 $T=667920 421600 0 0 $X=667730 $Y=421360
X1142 1 2 445 395 2 1798 1 sky130_fd_sc_hd__dfxtp_1 $T=668840 378080 0 0 $X=668650 $Y=377840
X1143 1 2 1765 402 2 1800 1 sky130_fd_sc_hd__dfxtp_1 $T=669300 394400 0 0 $X=669110 $Y=394160
X1144 1 2 1786 372 2 1803 1 sky130_fd_sc_hd__dfxtp_1 $T=672060 437920 1 0 $X=671870 $Y=434960
X1145 1 2 1802 372 2 1830 1 sky130_fd_sc_hd__dfxtp_1 $T=688160 427040 0 0 $X=687970 $Y=426800
X1146 1 2 1828 395 2 1846 1 sky130_fd_sc_hd__dfxtp_1 $T=694600 394400 0 0 $X=694410 $Y=394160
X1147 1 2 1826 378 2 1860 1 sky130_fd_sc_hd__dfxtp_1 $T=698740 410720 0 0 $X=698550 $Y=410480
X1148 1 2 524 521 25 513 9 524 ICV_13 $T=6900 399840 0 0 $X=6710 $Y=399600
X1149 1 2 525 521 24 513 10 518 ICV_13 $T=6900 410720 1 0 $X=6710 $Y=407760
X1150 1 2 526 533 24 514 11 526 ICV_13 $T=6900 432480 1 0 $X=6710 $Y=429520
X1151 1 2 527 533 25 514 9 527 ICV_13 $T=6900 437920 1 0 $X=6710 $Y=434960
X1152 1 2 544 533 23 514 13 544 ICV_13 $T=13800 427040 0 0 $X=13610 $Y=426800
X1153 1 2 546 543 34 517 28 546 ICV_13 $T=18400 383520 0 0 $X=18210 $Y=383280
X1154 1 2 561 543 37 517 30 549 ICV_13 $T=20240 388960 1 0 $X=20050 $Y=386000
X1155 1 2 558 534 36 515 30 558 ICV_13 $T=20240 416160 1 0 $X=20050 $Y=413200
X1156 1 2 553 533 34 514 30 559 ICV_13 $T=20240 437920 1 0 $X=20050 $Y=434960
X1157 1 2 547 543 31 517 29 561 ICV_13 $T=21160 394400 1 0 $X=20970 $Y=391440
X1158 1 2 577 580 25 567 10 582 ICV_13 $T=34040 394400 0 0 $X=33850 $Y=394160
X1159 1 2 583 580 37 567 29 583 ICV_13 $T=34040 399840 0 0 $X=33850 $Y=399600
X1160 1 2 593 43 37 555 17 590 ICV_13 $T=38180 432480 0 0 $X=37990 $Y=432240
X1161 1 2 599 580 24 567 11 599 ICV_13 $T=41400 388960 0 0 $X=41210 $Y=388720
X1162 1 2 579 45 16 597 9 49 ICV_13 $T=47380 378080 0 0 $X=47190 $Y=377840
X1163 1 2 611 52 31 48 17 611 ICV_13 $T=50600 432480 1 0 $X=50410 $Y=429520
X1164 1 2 625 615 24 604 11 625 ICV_13 $T=53820 410720 1 0 $X=53630 $Y=407760
X1165 1 2 616 615 34 604 17 627 ICV_13 $T=54280 416160 1 0 $X=54090 $Y=413200
X1166 1 2 628 605 37 594 29 628 ICV_13 $T=55200 405280 1 0 $X=55010 $Y=402320
X1167 1 2 650 51 37 597 29 650 ICV_13 $T=66240 378080 0 0 $X=66050 $Y=377840
X1168 1 2 643 58 31 56 13 651 ICV_13 $T=66240 432480 0 0 $X=66050 $Y=432240
X1169 1 2 653 58 25 56 11 647 ICV_13 $T=66240 437920 0 0 $X=66050 $Y=437680
X1170 1 2 663 648 31 635 9 662 ICV_13 $T=73140 405280 0 0 $X=72950 $Y=405040
X1171 1 2 669 648 34 635 11 660 ICV_13 $T=75440 399840 0 0 $X=75250 $Y=399600
X1172 1 2 672 58 34 56 28 672 ICV_13 $T=76360 443360 1 0 $X=76170 $Y=440400
X1173 1 2 674 63 37 61 29 674 ICV_13 $T=77740 378080 0 0 $X=77550 $Y=377840
X1174 1 2 675 58 36 56 30 675 ICV_13 $T=77740 432480 0 0 $X=77550 $Y=432240
X1175 1 2 699 71 31 64 17 699 ICV_13 $T=90160 432480 0 0 $X=89970 $Y=432240
X1176 1 2 693 71 37 64 10 70 ICV_13 $T=90160 437920 0 0 $X=89970 $Y=437680
X1177 1 2 686 673 23 665 30 691 ICV_13 $T=92460 421600 1 0 $X=92270 $Y=418640
X1178 1 2 722 71 36 64 30 722 ICV_13 $T=104420 437920 1 0 $X=104230 $Y=434960
X1179 1 2 725 732 23 711 17 726 ICV_13 $T=105340 427040 0 0 $X=105150 $Y=426800
X1180 1 2 721 66 31 664 11 727 ICV_13 $T=105800 383520 0 0 $X=105610 $Y=383280
X1181 1 2 729 720 34 712 28 729 ICV_13 $T=106260 405280 0 0 $X=106070 $Y=405040
X1182 1 2 742 716 31 695 17 742 ICV_13 $T=111780 394400 1 0 $X=111590 $Y=391440
X1183 1 2 713 716 34 695 9 743 ICV_13 $T=111780 399840 1 0 $X=111590 $Y=396880
X1184 1 2 744 720 36 712 30 744 ICV_13 $T=112240 410720 1 0 $X=112050 $Y=407760
X1185 1 2 751 720 31 712 17 751 ICV_13 $T=119140 416160 1 0 $X=118950 $Y=413200
X1186 1 2 753 732 25 711 9 753 ICV_13 $T=119600 421600 1 0 $X=119410 $Y=418640
X1187 1 2 754 720 25 712 9 754 ICV_13 $T=120060 410720 0 0 $X=119870 $Y=410480
X1188 1 2 760 758 34 746 28 760 ICV_13 $T=124200 394400 0 0 $X=124010 $Y=394160
X1189 1 2 761 758 31 746 9 764 ICV_13 $T=126040 388960 0 0 $X=125850 $Y=388720
X1190 1 2 767 768 34 749 28 767 ICV_13 $T=127420 432480 0 0 $X=127230 $Y=432240
X1191 1 2 775 773 23 759 13 775 ICV_13 $T=132020 416160 0 0 $X=131830 $Y=415920
X1192 1 2 790 768 25 749 11 791 ICV_13 $T=139840 432480 1 0 $X=139650 $Y=429520
X1193 1 2 801 809 123 792 111 801 ICV_13 $T=147660 410720 1 0 $X=147470 $Y=407760
X1194 1 2 803 802 123 793 111 803 ICV_13 $T=148120 388960 1 0 $X=147930 $Y=386000
X1195 1 2 805 809 119 792 112 805 ICV_13 $T=148120 410720 0 0 $X=147930 $Y=410480
X1196 1 2 806 120 123 108 111 806 ICV_13 $T=148120 443360 1 0 $X=147930 $Y=440400
X1197 1 2 807 798 123 794 111 807 ICV_13 $T=148580 394400 0 0 $X=148390 $Y=394160
X1198 1 2 832 120 129 108 125 832 ICV_13 $T=160540 443360 1 0 $X=160350 $Y=440400
X1199 1 2 835 819 130 795 126 835 ICV_13 $T=161000 427040 0 0 $X=160810 $Y=426800
X1200 1 2 859 116 128 121 125 133 ICV_13 $T=173880 383520 1 0 $X=173690 $Y=380560
X1201 1 2 863 844 123 132 111 863 ICV_13 $T=174340 432480 0 0 $X=174150 $Y=432240
X1202 1 2 838 819 131 848 111 866 ICV_13 $T=175260 421600 1 0 $X=175070 $Y=418640
X1203 1 2 134 844 128 132 113 867 ICV_13 $T=175720 443360 1 0 $X=175530 $Y=440400
X1204 1 2 884 888 129 874 127 883 ICV_13 $T=189520 388960 1 0 $X=189330 $Y=386000
X1205 1 2 887 888 128 874 124 887 ICV_13 $T=189980 383520 0 0 $X=189790 $Y=383280
X1206 1 2 141 140 129 137 127 894 ICV_13 $T=190440 437920 0 0 $X=190250 $Y=437680
X1207 1 2 908 888 119 874 112 908 ICV_13 $T=202400 383520 0 0 $X=202210 $Y=383280
X1208 1 2 909 888 123 874 111 909 ICV_13 $T=202400 388960 0 0 $X=202210 $Y=388720
X1209 1 2 913 890 119 879 112 913 ICV_13 $T=202400 427040 1 0 $X=202210 $Y=424080
X1210 1 2 939 147 118 931 127 937 ICV_13 $T=216660 437920 1 0 $X=216470 $Y=434960
X1211 1 2 968 936 119 926 109 967 ICV_13 $T=227700 394400 1 0 $X=227510 $Y=391440
X1212 1 2 971 949 131 932 127 971 ICV_13 $T=230460 421600 0 0 $X=230270 $Y=421360
X1213 1 2 974 976 123 957 124 973 ICV_13 $T=232760 432480 1 0 $X=232570 $Y=429520
X1214 1 2 985 951 123 927 124 987 ICV_13 $T=237820 383520 0 0 $X=237630 $Y=383280
X1215 1 2 1001 976 129 957 125 1001 ICV_13 $T=245640 432480 1 0 $X=245450 $Y=429520
X1216 1 2 1012 1008 131 969 127 991 ICV_13 $T=246560 399840 0 0 $X=246370 $Y=399600
X1217 1 2 1024 165 118 160 109 1024 ICV_13 $T=258060 383520 1 0 $X=257870 $Y=380560
X1218 1 2 1028 1019 119 1014 112 1028 ICV_13 $T=258520 427040 0 0 $X=258330 $Y=426800
X1219 1 2 1039 1038 118 1023 126 1040 ICV_13 $T=264040 410720 0 0 $X=263850 $Y=410480
X1220 1 2 1043 1019 123 1014 111 1043 ICV_13 $T=265420 421600 0 0 $X=265230 $Y=421360
X1221 1 2 1045 1038 123 1023 127 1037 ICV_13 $T=273240 405280 0 0 $X=273050 $Y=405040
X1222 1 2 1062 1038 122 1023 113 1062 ICV_13 $T=276460 410720 1 0 $X=276270 $Y=407760
X1223 1 2 1065 1067 122 1050 113 1065 ICV_13 $T=276920 432480 1 0 $X=276730 $Y=429520
X1224 1 2 1080 171 128 169 124 1080 ICV_13 $T=286580 378080 0 0 $X=286390 $Y=377840
X1225 1 2 1086 1067 123 1050 127 1085 ICV_13 $T=287500 437920 1 0 $X=287310 $Y=434960
X1226 1 2 1087 1092 128 1072 124 1087 ICV_13 $T=287960 388960 1 0 $X=287770 $Y=386000
X1227 1 2 1088 1067 119 1050 112 1088 ICV_13 $T=287960 427040 1 0 $X=287770 $Y=424080
X1228 1 2 173 174 129 1072 127 1089 ICV_13 $T=288420 383520 1 0 $X=288230 $Y=380560
X1229 1 2 1093 1092 122 1041 127 1073 ICV_13 $T=288880 394400 1 0 $X=288690 $Y=391440
X1230 1 2 1105 1079 119 1066 112 1105 ICV_13 $T=297160 416160 0 0 $X=296970 $Y=415920
X1231 1 2 1109 171 130 169 126 1109 ICV_13 $T=300840 383520 1 0 $X=300650 $Y=380560
X1232 1 2 1119 1097 122 1076 111 1113 ICV_13 $T=302220 399840 0 0 $X=302030 $Y=399600
X1233 1 2 1115 1102 122 1103 113 1115 ICV_13 $T=302220 432480 0 0 $X=302030 $Y=432240
X1234 1 2 1120 1102 119 1103 112 1120 ICV_13 $T=303140 437920 1 0 $X=302950 $Y=434960
X1235 1 2 1125 1092 123 1072 112 1124 ICV_13 $T=304060 388960 1 0 $X=303870 $Y=386000
X1236 1 2 1127 1107 122 1104 109 1134 ICV_13 $T=314640 416160 1 0 $X=314450 $Y=413200
X1237 1 2 1116 1092 118 1128 184 1136 ICV_13 $T=315100 394400 1 0 $X=314910 $Y=391440
X1238 1 2 210 214 221 1129 189 1148 ICV_13 $T=322000 378080 0 0 $X=321810 $Y=377840
X1239 1 2 1162 1144 236 1128 211 1162 ICV_13 $T=328900 388960 0 0 $X=328710 $Y=388720
X1240 1 2 1147 218 195 1146 213 229 ICV_13 $T=328900 437920 0 0 $X=328710 $Y=437680
X1241 1 2 1164 1144 237 1128 219 1164 ICV_13 $T=329820 394400 0 0 $X=329630 $Y=394160
X1242 1 2 1174 218 183 193 199 1174 ICV_13 $T=334420 443360 1 0 $X=334230 $Y=440400
X1243 1 2 1184 215 195 1146 196 1184 ICV_13 $T=339940 437920 1 0 $X=339750 $Y=434960
X1244 1 2 1178 1168 206 1167 191 1166 ICV_13 $T=341780 399840 1 0 $X=341590 $Y=396880
X1245 1 2 1190 1183 239 1167 185 1169 ICV_13 $T=342700 399840 0 0 $X=342510 $Y=399600
X1246 1 2 1201 1207 221 241 191 1201 ICV_13 $T=349600 388960 0 0 $X=349410 $Y=388720
X1247 1 2 1212 1183 188 1173 204 1212 ICV_13 $T=356040 416160 0 0 $X=355850 $Y=415920
X1248 1 2 1215 1183 195 1173 196 1215 ICV_13 $T=356960 416160 1 0 $X=356770 $Y=413200
X1249 1 2 1226 1207 209 241 189 1226 ICV_13 $T=362020 383520 1 0 $X=361830 $Y=380560
X1250 1 2 1232 1239 220 1233 228 1222 ICV_13 $T=369840 427040 1 0 $X=369650 $Y=424080
X1251 1 2 1245 1239 195 1211 204 1244 ICV_13 $T=370760 416160 0 0 $X=370570 $Y=415920
X1252 1 2 1250 1223 195 1233 196 1250 ICV_13 $T=372600 432480 1 0 $X=372410 $Y=429520
X1253 1 2 1262 1264 205 1256 185 1262 ICV_13 $T=383640 394400 0 0 $X=383450 $Y=394160
X1254 1 2 1266 1264 236 1256 211 1266 ICV_13 $T=385020 388960 1 0 $X=384830 $Y=386000
X1255 1 2 1267 1264 209 1256 189 1267 ICV_13 $T=385020 394400 1 0 $X=384830 $Y=391440
X1256 1 2 1269 1264 237 1256 191 1268 ICV_13 $T=385020 399840 1 0 $X=384830 $Y=396880
X1257 1 2 1292 1290 236 1282 184 1295 ICV_13 $T=398820 383520 0 0 $X=398630 $Y=383280
X1258 1 2 1311 281 236 268 191 280 ICV_13 $T=413540 378080 0 0 $X=413350 $Y=377840
X1259 1 2 1332 282 237 1300 184 1337 ICV_13 $T=417220 394400 1 0 $X=417030 $Y=391440
X1260 1 2 1348 1334 195 1321 224 1346 ICV_13 $T=424580 416160 1 0 $X=424390 $Y=413200
X1261 1 2 1352 1334 187 1321 202 1352 ICV_13 $T=426420 410720 1 0 $X=426230 $Y=407760
X1262 1 2 1354 1334 192 1321 228 1354 ICV_13 $T=426880 410720 0 0 $X=426690 $Y=410480
X1263 1 2 1341 1334 183 1321 213 1351 ICV_13 $T=426880 416160 0 0 $X=426690 $Y=415920
X1264 1 2 1367 1371 220 1353 227 1368 ICV_13 $T=434700 437920 0 0 $X=434510 $Y=437680
X1265 1 2 1373 1350 206 1340 190 1373 ICV_13 $T=437460 399840 0 0 $X=437270 $Y=399600
X1266 1 2 1378 295 206 293 190 1378 ICV_13 $T=441140 378080 0 0 $X=440950 $Y=377840
X1267 1 2 1394 1380 183 1364 199 1394 ICV_13 $T=448040 421600 1 0 $X=447850 $Y=418640
X1268 1 2 1395 1399 205 1377 185 1395 ICV_13 $T=448500 399840 1 0 $X=448310 $Y=396880
X1269 1 2 1411 1414 187 1400 202 1411 ICV_13 $T=455860 432480 1 0 $X=455670 $Y=429520
X1270 1 2 1433 305 188 298 204 1433 ICV_13 $T=468740 437920 0 0 $X=468550 $Y=437680
X1271 1 2 1439 1443 209 1427 184 1437 ICV_13 $T=471040 394400 0 0 $X=470850 $Y=394160
X1272 1 2 1453 1447 195 1431 224 1450 ICV_13 $T=476560 416160 1 0 $X=476370 $Y=413200
X1273 1 2 1448 1447 239 1427 219 1463 ICV_13 $T=483920 405280 0 0 $X=483730 $Y=405040
X1274 1 2 1464 1447 192 1431 228 1464 ICV_13 $T=485300 410720 1 0 $X=485110 $Y=407760
X1275 1 2 1454 322 195 319 204 1451 ICV_13 $T=485300 437920 1 0 $X=485110 $Y=434960
X1276 1 2 1472 326 237 324 219 1472 ICV_13 $T=487600 378080 0 0 $X=487410 $Y=377840
X1277 1 2 1476 322 180 319 224 1476 ICV_13 $T=488520 432480 0 0 $X=488330 $Y=432240
X1278 1 2 1502 326 205 324 185 1502 ICV_13 $T=503700 383520 1 0 $X=503510 $Y=380560
X1279 1 2 1503 323 205 1456 185 1503 ICV_13 $T=503700 399840 1 0 $X=503510 $Y=396880
X1280 1 2 1508 1487 180 1470 224 1508 ICV_13 $T=511060 432480 0 0 $X=510870 $Y=432240
X1281 1 2 1514 336 180 332 224 1514 ICV_13 $T=512900 437920 0 0 $X=512710 $Y=437680
X1282 1 2 1529 1516 368 1519 358 1529 ICV_13 $T=526240 427040 1 0 $X=526050 $Y=424080
X1283 1 2 1536 1516 371 1519 372 1536 ICV_13 $T=537740 427040 1 0 $X=537550 $Y=424080
X1284 1 2 1562 1553 392 1543 400 1562 ICV_13 $T=552920 388960 0 0 $X=552730 $Y=388720
X1285 1 2 1549 401 371 385 357 1564 ICV_13 $T=555220 437920 0 0 $X=555030 $Y=437680
X1286 1 2 1570 1545 345 1539 381 1570 ICV_13 $T=558440 410720 1 0 $X=558250 $Y=407760
X1287 1 2 1577 1553 389 1543 406 1577 ICV_13 $T=560280 394400 1 0 $X=560090 $Y=391440
X1288 1 2 1581 1553 391 1543 407 1581 ICV_13 $T=560740 388960 1 0 $X=560550 $Y=386000
X1289 1 2 1594 1545 371 1539 372 1594 ICV_13 $T=567180 416160 1 0 $X=566990 $Y=413200
X1290 1 2 1566 401 345 1580 360 1595 ICV_13 $T=567180 437920 1 0 $X=566990 $Y=434960
X1291 1 2 1595 1589 343 1580 359 1593 ICV_13 $T=567640 432480 1 0 $X=567450 $Y=429520
X1292 1 2 1601 1586 352 1587 407 1600 ICV_13 $T=572240 394400 0 0 $X=572050 $Y=394160
X1293 1 2 1616 1589 363 1580 381 1614 ICV_13 $T=577300 427040 0 0 $X=577110 $Y=426800
X1294 1 2 1622 1590 386 1592 393 1622 ICV_13 $T=581440 388960 1 0 $X=581250 $Y=386000
X1295 1 2 1624 1589 371 1580 372 1624 ICV_13 $T=581440 443360 1 0 $X=581250 $Y=440400
X1296 1 2 1630 1586 389 1587 406 1630 ICV_13 $T=586500 394400 1 0 $X=586310 $Y=391440
X1297 1 2 1626 1586 392 1587 405 1613 ICV_13 $T=587420 399840 1 0 $X=587230 $Y=396880
X1298 1 2 1596 1589 366 418 359 1644 ICV_13 $T=592020 437920 1 0 $X=591830 $Y=434960
X1299 1 2 1645 1590 388 1592 405 1645 ICV_13 $T=592940 388960 1 0 $X=592750 $Y=386000
X1300 1 2 1663 1638 355 1621 359 1663 ICV_13 $T=600300 432480 0 0 $X=600110 $Y=432240
X1301 1 2 1672 1667 368 1658 358 1672 ICV_13 $T=605360 410720 0 0 $X=605170 $Y=410480
X1302 1 2 1676 1655 397 1658 381 1668 ICV_13 $T=607200 405280 0 0 $X=607010 $Y=405040
X1303 1 2 1691 1690 367 1671 357 1691 ICV_13 $T=613640 427040 1 0 $X=613450 $Y=424080
X1304 1 2 427 422 389 421 395 1695 ICV_13 $T=616860 383520 1 0 $X=616670 $Y=380560
X1305 1 2 1713 1689 368 1698 358 1713 ICV_13 $T=625600 416160 1 0 $X=625410 $Y=413200
X1306 1 2 1718 1707 389 1685 403 1704 ICV_13 $T=626980 388960 0 0 $X=626790 $Y=388720
X1307 1 2 1701 1643 345 1698 359 1726 ICV_13 $T=634340 421600 0 0 $X=634150 $Y=421360
X1308 1 2 1731 434 368 429 358 1731 ICV_13 $T=636640 427040 0 0 $X=636450 $Y=426800
X1309 1 2 1733 434 355 429 357 1732 ICV_13 $T=637560 432480 1 0 $X=637370 $Y=429520
X1310 1 2 1738 1728 352 1721 402 1738 ICV_13 $T=639400 399840 1 0 $X=639210 $Y=396880
X1311 1 2 1781 440 371 1747 378 1778 ICV_13 $T=661480 432480 0 0 $X=661290 $Y=432240
X1312 1 2 1787 1770 389 1765 406 1787 ICV_13 $T=665620 394400 1 0 $X=665430 $Y=391440
X1313 1 2 1789 1772 345 1751 378 1783 ICV_13 $T=666080 416160 0 0 $X=665890 $Y=415920
X1314 1 2 1800 1770 352 1784 395 1817 ICV_13 $T=679420 399840 0 0 $X=679230 $Y=399600
X1315 1 2 1818 1799 355 1777 360 1819 ICV_13 $T=679420 416160 0 0 $X=679230 $Y=415920
X1316 1 2 1816 447 388 1784 402 1807 ICV_13 $T=680340 394400 1 0 $X=680150 $Y=391440
X1317 1 2 1836 1842 367 1826 381 1835 ICV_13 $T=693680 405280 1 0 $X=693490 $Y=402320
X1318 1 2 1847 1810 355 1786 381 1838 ICV_13 $T=693680 432480 1 0 $X=693490 $Y=429520
X1319 1 2 1839 1804 363 1786 365 1839 ICV_13 $T=693680 437920 1 0 $X=693490 $Y=434960
X1320 1 2 1850 1842 363 1826 365 1850 ICV_13 $T=695060 405280 0 0 $X=694870 $Y=405040
X1321 1 2 1855 1842 355 1802 359 1847 ICV_13 $T=695520 427040 0 0 $X=695330 $Y=426800
X1322 1 2 1870 1878 343 1857 360 1870 ICV_13 $T=707480 421600 0 0 $X=707290 $Y=421360
X1323 1 2 1873 1878 355 1857 359 1873 ICV_13 $T=707940 427040 1 0 $X=707750 $Y=424080
X1324 1 2 1880 1885 392 1862 395 1879 ICV_13 $T=709320 383520 0 0 $X=709130 $Y=383280
X1325 1 2 1881 1869 371 1864 372 1881 ICV_13 $T=709780 410720 1 0 $X=709590 $Y=407760
X1326 1 2 1883 462 363 1859 359 1882 ICV_13 $T=709780 437920 1 0 $X=709590 $Y=434960
X1327 1 2 1886 1865 392 1866 395 1887 ICV_13 $T=711620 399840 0 0 $X=711430 $Y=399600
X1328 1 2 1900 1869 368 1864 358 1900 ICV_13 $T=722660 410720 1 0 $X=722470 $Y=407760
X1329 1 2 1914 1885 391 1862 407 1914 ICV_13 $T=725420 383520 1 0 $X=725230 $Y=380560
X1330 1 2 515 29 556 530 534 16 ICV_14 $T=18860 421600 0 0 $X=18670 $Y=421360
X1331 1 2 567 9 577 581 580 34 ICV_14 $T=32660 394400 1 0 $X=32470 $Y=391440
X1332 1 2 594 28 630 633 634 25 ICV_14 $T=55660 394400 1 0 $X=55470 $Y=391440
X1333 1 2 637 11 685 685 634 24 ICV_14 $T=83720 399840 1 0 $X=83530 $Y=396880
X1334 1 2 712 29 735 735 720 37 ICV_14 $T=106720 416160 1 0 $X=106530 $Y=413200
X1335 1 2 749 29 766 762 768 31 ICV_14 $T=125580 427040 0 0 $X=125390 $Y=426800
X1336 1 2 794 125 836 823 798 128 ICV_14 $T=160540 405280 1 0 $X=160350 $Y=402320
X1337 1 2 795 127 838 840 819 129 ICV_14 $T=160540 421600 0 0 $X=160350 $Y=421360
X1338 1 2 132 126 857 853 844 118 ICV_14 $T=172960 432480 1 0 $X=172770 $Y=429520
X1339 1 2 848 109 871 866 854 123 ICV_14 $T=176640 416160 0 0 $X=176450 $Y=415920
X1340 1 2 848 113 885 885 854 122 ICV_14 $T=188600 416160 1 0 $X=188410 $Y=413200
X1341 1 2 137 126 902 902 140 130 ICV_14 $T=196420 443360 1 0 $X=196230 $Y=440400
X1342 1 2 926 126 934 934 936 130 ICV_14 $T=213900 388960 0 0 $X=213710 $Y=388720
X1343 1 2 901 111 940 940 918 123 ICV_14 $T=215280 405280 0 0 $X=215090 $Y=405040
X1344 1 2 957 109 977 977 976 118 ICV_14 $T=232760 432480 0 0 $X=232570 $Y=432240
X1345 1 2 957 112 1005 1005 976 119 ICV_14 $T=245180 432480 0 0 $X=244990 $Y=432240
X1346 1 2 1104 112 1112 1112 1107 119 ICV_14 $T=300840 421600 1 0 $X=300650 $Y=418640
X1347 1 2 1076 125 1114 1113 1097 123 ICV_14 $T=301300 405280 0 0 $X=301110 $Y=405040
X1348 1 2 1103 126 1139 1135 1102 129 ICV_14 $T=314640 432480 0 0 $X=314450 $Y=432240
X1349 1 2 1103 127 1140 1140 1102 131 ICV_14 $T=314640 437920 0 0 $X=314450 $Y=437680
X1350 1 2 1173 213 1191 1186 1183 180 ICV_14 $T=342700 410720 0 0 $X=342510 $Y=410480
X1351 1 2 241 219 1206 1206 1207 237 ICV_14 $T=350060 378080 0 0 $X=349870 $Y=377840
X1352 1 2 248 202 1219 1219 251 187 ICV_14 $T=356500 437920 0 0 $X=356310 $Y=437680
X1353 1 2 1185 227 1220 1200 1199 180 ICV_14 $T=357420 432480 0 0 $X=357230 $Y=432240
X1354 1 2 1185 202 1221 1221 1199 187 ICV_14 $T=357880 421600 0 0 $X=357690 $Y=421360
X1355 1 2 1210 190 1234 1234 1225 206 ICV_14 $T=362480 399840 1 0 $X=362290 $Y=396880
X1356 1 2 1256 190 1265 1265 1264 206 ICV_14 $T=383640 399840 0 0 $X=383450 $Y=399600
X1357 1 2 1259 224 1285 1285 1274 180 ICV_14 $T=392840 416160 1 0 $X=392650 $Y=413200
X1358 1 2 286 199 1357 1357 290 183 ICV_14 $T=427800 443360 1 0 $X=427610 $Y=440400
X1359 1 2 1340 184 1362 1363 282 209 ICV_14 $T=429640 388960 0 0 $X=429450 $Y=388720
X1360 1 2 1427 190 1460 1463 1443 237 ICV_14 $T=483000 405280 1 0 $X=482810 $Y=402320
X1361 1 2 324 191 1469 1469 326 221 ICV_14 $T=485300 383520 0 0 $X=485110 $Y=383280
X1362 1 2 1483 213 1492 1492 1480 220 ICV_14 $T=497260 416160 1 0 $X=497070 $Y=413200
X1363 1 2 1592 400 1610 1607 1590 387 ICV_14 $T=574540 383520 0 0 $X=574350 $Y=383280
X1364 1 2 418 358 1680 425 426 366 ICV_14 $T=609960 437920 0 0 $X=609770 $Y=437680
X1365 1 2 421 393 1696 1695 422 397 ICV_14 $T=615940 388960 1 0 $X=615750 $Y=386000
X1366 1 2 437 395 1763 1759 439 386 ICV_14 $T=651360 383520 1 0 $X=651170 $Y=380560
X1367 1 2 1751 360 1767 1767 1772 343 ICV_14 $T=652740 427040 1 0 $X=652550 $Y=424080
X1368 1 2 1828 400 1845 1840 1851 389 ICV_14 $T=693680 388960 1 0 $X=693490 $Y=386000
X1369 1 2 1857 372 1877 1877 1878 371 ICV_14 $T=707940 421600 1 0 $X=707750 $Y=418640
X1370 1 2 1866 400 1886 1884 1885 352 ICV_14 $T=709780 394400 0 0 $X=709590 $Y=394160
X1371 1 2 587 576 37 564 10 584 575 576 36 ICV_15 $T=34040 410720 0 0 $X=33850 $Y=410480
X1372 1 2 595 554 37 564 17 588 588 576 31 ICV_15 $T=35880 416160 0 0 $X=35690 $Y=415920
X1373 1 2 54 52 34 48 11 614 592 43 16 ICV_15 $T=51060 443360 1 0 $X=50870 $Y=440400
X1374 1 2 697 683 37 676 30 707 707 683 36 ICV_15 $T=94300 410720 0 0 $X=94110 $Y=410480
X1375 1 2 774 773 16 759 17 780 780 773 31 ICV_15 $T=132480 416160 1 0 $X=132290 $Y=413200
X1376 1 2 860 116 130 121 126 860 851 802 131 ICV_15 $T=174340 383520 0 0 $X=174150 $Y=383280
X1377 1 2 944 951 129 927 112 952 952 951 119 ICV_15 $T=219420 388960 1 0 $X=219230 $Y=386000
X1378 1 2 1009 162 119 157 112 1009 1006 162 122 ICV_15 $T=246560 437920 1 0 $X=246370 $Y=434960
X1379 1 2 1022 1008 123 984 111 1022 1017 990 118 ICV_15 $T=256680 399840 1 0 $X=256490 $Y=396880
X1380 1 2 1148 217 209 1129 185 201 1142 1144 209 ICV_15 $T=318320 383520 0 0 $X=318130 $Y=383280
X1381 1 2 1381 1380 220 1353 202 1386 1386 1371 187 ICV_15 $T=444360 427040 1 0 $X=444170 $Y=424080
X1382 1 2 1612 1590 352 1592 402 1612 1600 1586 391 ICV_15 $T=576840 388960 0 0 $X=576650 $Y=388720
X1383 1 2 1633 1637 367 1618 381 1642 1647 1637 355 ICV_15 $T=592940 410720 1 0 $X=592750 $Y=407760
X1384 1 2 1675 422 391 421 407 1675 423 422 392 ICV_15 $T=606740 378080 0 0 $X=606550 $Y=377840
X1385 1 2 1897 1874 345 1859 381 1897 1867 1874 363 ICV_15 $T=721740 432480 1 0 $X=721550 $Y=429520
X1386 1 2 465 464 387 1862 405 1912 1912 1885 388 ICV_15 $T=724960 388960 1 0 $X=724770 $Y=386000
X1387 1 2 515 11 529 532 534 25 ICV_16 $T=6900 416160 1 0 $X=6710 $Y=413200
X1388 1 2 515 10 530 531 533 16 ICV_16 $T=6900 421600 0 0 $X=6710 $Y=421360
X1389 1 2 631 28 640 640 644 34 ICV_16 $T=63020 421600 1 0 $X=62830 $Y=418640
X1390 1 2 664 13 723 723 66 23 ICV_16 $T=104420 388960 1 0 $X=104230 $Y=386000
X1391 1 2 711 30 745 726 732 31 ICV_16 $T=112240 432480 1 0 $X=112050 $Y=429520
X1392 1 2 759 30 772 772 773 36 ICV_16 $T=131100 399840 0 0 $X=130910 $Y=399600
X1393 1 2 759 10 774 779 773 25 ICV_16 $T=131560 410720 0 0 $X=131370 $Y=410480
X1394 1 2 848 127 886 878 854 129 ICV_16 $T=189060 416160 0 0 $X=188870 $Y=415920
X1395 1 2 846 109 893 886 854 131 ICV_16 $T=189980 410720 0 0 $X=189790 $Y=410480
X1396 1 2 137 111 900 900 140 123 ICV_16 $T=190900 437920 1 0 $X=190710 $Y=434960
X1397 1 2 879 124 916 916 890 128 ICV_16 $T=202400 421600 0 0 $X=202210 $Y=421360
X1398 1 2 932 125 962 962 949 129 ICV_16 $T=224940 427040 1 0 $X=224750 $Y=424080
X1399 1 2 984 124 996 996 1008 128 ICV_16 $T=244720 394400 1 0 $X=244530 $Y=391440
X1400 1 2 965 112 997 997 980 119 ICV_16 $T=244720 416160 0 0 $X=244530 $Y=415920
X1401 1 2 957 113 998 992 976 131 ICV_16 $T=244720 427040 1 0 $X=244530 $Y=424080
X1402 1 2 1066 124 1078 1083 1079 123 ICV_16 $T=287040 416160 1 0 $X=286850 $Y=413200
X1403 1 2 1103 111 1132 1132 1102 123 ICV_16 $T=312340 432480 1 0 $X=312150 $Y=429520
X1404 1 2 1103 109 1138 1138 1102 118 ICV_16 $T=314640 437920 1 0 $X=314450 $Y=434960
X1405 1 2 241 185 1203 1203 1207 205 ICV_16 $T=350060 383520 0 0 $X=349870 $Y=383280
X1406 1 2 1167 211 1204 1179 1168 230 ICV_16 $T=350060 394400 0 0 $X=349870 $Y=394160
X1407 1 2 1256 184 1261 1261 1264 222 ICV_16 $T=382720 383520 0 0 $X=382530 $Y=383280
X1408 1 2 1233 227 1278 1278 1223 239 ICV_16 $T=386400 421600 0 0 $X=386210 $Y=421360
X1409 1 2 1282 190 1291 1291 1290 206 ICV_16 $T=396520 394400 1 0 $X=396330 $Y=391440
X1410 1 2 1306 202 1320 1320 1323 187 ICV_16 $T=409400 427040 0 0 $X=409210 $Y=426800
X1411 1 2 1340 211 1358 1362 1350 222 ICV_16 $T=428720 394400 1 0 $X=428530 $Y=391440
X1412 1 2 293 211 1383 1383 295 236 ICV_16 $T=441140 383520 0 0 $X=440950 $Y=383280
X1413 1 2 298 224 1410 1409 305 195 ICV_16 $T=454940 437920 0 0 $X=454750 $Y=437680
X1414 1 2 1408 191 310 1426 312 236 ICV_16 $T=462300 383520 0 0 $X=462110 $Y=383280
X1415 1 2 1400 204 1455 1455 1414 188 ICV_16 $T=478860 427040 1 0 $X=478670 $Y=424080
X1416 1 2 1470 196 1510 1510 1487 195 ICV_16 $T=511060 427040 1 0 $X=510870 $Y=424080
X1417 1 2 1517 358 1524 1524 1527 368 ICV_16 $T=524400 437920 0 0 $X=524210 $Y=437680
X1418 1 2 1540 365 1568 1568 1550 363 ICV_16 $T=557060 421600 1 0 $X=556870 $Y=418640
X1419 1 2 1540 358 1578 1571 1550 355 ICV_16 $T=559820 427040 1 0 $X=559630 $Y=424080
X1420 1 2 390 407 1583 1557 398 397 ICV_16 $T=560740 383520 1 0 $X=560550 $Y=380560
X1421 1 2 1641 407 1679 1678 1655 392 ICV_16 $T=609500 394400 0 0 $X=609310 $Y=394160
X1422 1 2 1698 381 1687 1717 1689 367 ICV_16 $T=625140 410720 1 0 $X=624950 $Y=407760
X1423 1 2 1721 393 1761 1760 1728 388 ICV_16 $T=650900 399840 1 0 $X=650710 $Y=396880
X1424 1 2 445 393 1795 1795 448 386 ICV_16 $T=667920 383520 1 0 $X=667730 $Y=380560
X1425 1 2 1786 358 1805 1805 1804 368 ICV_16 $T=672980 443360 1 0 $X=672790 $Y=440400
X1426 1 2 1802 378 1829 1829 1810 366 ICV_16 $T=686780 421600 0 0 $X=686590 $Y=421360
X1427 1 2 1786 378 1834 1834 1804 366 ICV_16 $T=692760 432480 0 0 $X=692570 $Y=432240
X1428 1 2 5 11 528 528 20 24 ICV_17 $T=5520 443360 1 0 $X=5330 $Y=440400
X1429 1 2 517 17 547 539 543 23 ICV_17 $T=17020 388960 0 0 $X=16830 $Y=388720
X1430 1 2 513 29 562 562 521 37 ICV_17 $T=20240 405280 1 0 $X=20050 $Y=402320
X1431 1 2 564 11 572 574 576 23 ICV_17 $T=30360 410720 1 0 $X=30170 $Y=407760
X1432 1 2 555 29 595 590 554 31 ICV_17 $T=38180 421600 0 0 $X=37990 $Y=421360
X1433 1 2 56 17 643 647 58 24 ICV_17 $T=63020 437920 1 0 $X=62830 $Y=434960
X1434 1 2 631 13 661 659 644 36 ICV_17 $T=70380 421600 0 0 $X=70190 $Y=421360
X1435 1 2 64 13 694 694 71 23 ICV_17 $T=87860 443360 1 0 $X=87670 $Y=440400
X1436 1 2 712 11 728 709 716 16 ICV_17 $T=104420 405280 1 0 $X=104230 $Y=402320
X1437 1 2 711 29 730 730 732 37 ICV_17 $T=104880 421600 0 0 $X=104690 $Y=421360
X1438 1 2 89 30 756 756 87 36 ICV_17 $T=119600 437920 0 0 $X=119410 $Y=437680
X1439 1 2 108 124 822 822 120 128 ICV_17 $T=156860 432480 0 0 $X=156670 $Y=432240
X1440 1 2 795 125 840 811 819 118 ICV_17 $T=160540 421600 1 0 $X=160350 $Y=418640
X1441 1 2 848 124 889 889 854 128 ICV_17 $T=188600 421600 1 0 $X=188410 $Y=418640
X1442 1 2 901 112 917 917 918 119 ICV_17 $T=202400 405280 0 0 $X=202210 $Y=405040
X1443 1 2 137 124 921 919 140 118 ICV_17 $T=202400 437920 0 0 $X=202210 $Y=437680
X1444 1 2 984 112 999 999 1008 119 ICV_17 $T=244260 394400 0 0 $X=244070 $Y=394160
X1445 1 2 969 126 1003 1003 990 130 ICV_17 $T=244720 410720 1 0 $X=244530 $Y=407760
X1446 1 2 157 113 1006 159 161 131 ICV_17 $T=244720 443360 1 0 $X=244530 $Y=440400
X1447 1 2 157 111 1010 1010 162 123 ICV_17 $T=245180 437920 0 0 $X=244990 $Y=437680
X1448 1 2 157 125 1030 1032 162 130 ICV_17 $T=257600 443360 1 0 $X=257410 $Y=440400
X1449 1 2 1023 112 1046 1046 1038 119 ICV_17 $T=264960 416160 0 0 $X=264770 $Y=415920
X1450 1 2 157 124 1048 1048 162 128 ICV_17 $T=267260 437920 0 0 $X=267070 $Y=437680
X1451 1 2 1104 127 1131 1133 1107 128 ICV_17 $T=310960 427040 1 0 $X=310770 $Y=424080
X1452 1 2 1210 191 1249 1249 1225 221 ICV_17 $T=370760 399840 0 0 $X=370570 $Y=399600
X1453 1 2 1259 196 1277 1277 1274 195 ICV_17 $T=385020 421600 1 0 $X=384830 $Y=418640
X1454 1 2 1300 219 1314 1314 1317 237 ICV_17 $T=406180 405280 0 0 $X=405990 $Y=405040
X1455 1 2 1340 191 1349 1356 1350 205 ICV_17 $T=426880 405280 1 0 $X=426690 $Y=402320
X1456 1 2 1364 228 1376 1375 1380 188 ICV_17 $T=438380 410720 0 0 $X=438190 $Y=410480
X1457 1 2 1400 224 1412 1412 1414 180 ICV_17 $T=454940 427040 0 0 $X=454750 $Y=426800
X1458 1 2 1400 213 1413 1388 1371 192 ICV_17 $T=454940 432480 0 0 $X=454750 $Y=432240
X1459 1 2 1407 228 1424 1420 1403 180 ICV_17 $T=460460 410720 0 0 $X=460270 $Y=410480
X1460 1 2 1400 196 1436 1436 1414 195 ICV_17 $T=467820 432480 0 0 $X=467630 $Y=432240
X1461 1 2 1427 211 1457 1457 1443 236 ICV_17 $T=478860 394400 1 0 $X=478670 $Y=391440
X1462 1 2 1517 372 1531 1531 1527 371 ICV_17 $T=532680 443360 1 0 $X=532490 $Y=440400
X1463 1 2 1585 360 1604 1603 1597 368 ICV_17 $T=571320 421600 0 0 $X=571130 $Y=421360
X1464 1 2 1580 357 1611 1611 1589 367 ICV_17 $T=574080 432480 0 0 $X=573890 $Y=432240
X1465 1 2 415 407 1625 416 417 387 ICV_17 $T=581900 378080 0 0 $X=581710 $Y=377840
X1466 1 2 1730 365 1752 1748 1754 355 ICV_17 $T=644920 410720 1 0 $X=644730 $Y=407760
X1467 1 2 436 372 438 1736 434 345 ICV_17 $T=644920 443360 1 0 $X=644730 $Y=440400
X1468 1 2 1777 372 1813 1813 1799 371 ICV_17 $T=677120 416160 1 0 $X=676930 $Y=413200
X1469 1 2 456 402 1848 1848 457 352 ICV_17 $T=693680 378080 0 0 $X=693490 $Y=377840
X1470 1 2 1864 360 1876 1860 1842 366 ICV_17 $T=707480 410720 0 0 $X=707290 $Y=410480
X1471 1 2 461 406 1889 1879 1885 397 ICV_17 $T=709780 378080 0 0 $X=709590 $Y=377840
X1492 1 2 514 10 531 ICV_20 $T=6900 427040 1 0 $X=6710 $Y=424080
X1493 1 2 513 17 542 ICV_20 $T=11960 399840 1 0 $X=11770 $Y=396880
X1494 1 2 33 13 41 ICV_20 $T=25760 378080 0 0 $X=25570 $Y=377840
X1495 1 2 604 13 620 ICV_20 $T=51520 416160 0 0 $X=51330 $Y=415920
X1496 1 2 594 10 626 ICV_20 $T=53820 399840 0 0 $X=53630 $Y=399600
X1497 1 2 631 10 641 ICV_20 $T=63480 427040 1 0 $X=63290 $Y=424080
X1498 1 2 631 9 642 ICV_20 $T=63940 427040 0 0 $X=63750 $Y=426800
X1499 1 2 635 13 649 ICV_20 $T=65320 405280 0 0 $X=65130 $Y=405040
X1500 1 2 635 10 646 ICV_20 $T=65320 410720 1 0 $X=65130 $Y=407760
X1501 1 2 597 13 652 ICV_20 $T=66240 383520 0 0 $X=66050 $Y=383280
X1502 1 2 56 9 653 ICV_20 $T=66700 443360 1 0 $X=66510 $Y=440400
X1503 1 2 665 9 670 ICV_20 $T=81880 416160 0 0 $X=81690 $Y=415920
X1504 1 2 664 10 67 ICV_20 $T=84640 383520 1 0 $X=84450 $Y=380560
X1505 1 2 665 13 686 ICV_20 $T=84640 421600 1 0 $X=84450 $Y=418640
X1506 1 2 695 10 709 ICV_20 $T=96140 399840 1 0 $X=95950 $Y=396880
X1507 1 2 64 9 717 ICV_20 $T=101660 437920 0 0 $X=101470 $Y=437680
X1508 1 2 711 13 725 ICV_20 $T=104420 432480 1 0 $X=104230 $Y=429520
X1509 1 2 746 10 757 ICV_20 $T=123280 399840 1 0 $X=123090 $Y=396880
X1510 1 2 749 17 762 ICV_20 $T=124200 432480 1 0 $X=124010 $Y=429520
X1511 1 2 749 10 777 ICV_20 $T=138000 427040 0 0 $X=137810 $Y=426800
X1512 1 2 793 109 804 ICV_20 $T=147660 394400 1 0 $X=147470 $Y=391440
X1513 1 2 793 125 824 ICV_20 $T=158700 388960 0 0 $X=158510 $Y=388720
X1514 1 2 855 126 881 ICV_20 $T=186300 399840 0 0 $X=186110 $Y=399600
X1515 1 2 137 113 139 ICV_20 $T=188600 443360 1 0 $X=188410 $Y=440400
X1516 1 2 879 113 899 ICV_20 $T=191360 421600 0 0 $X=191170 $Y=421360
X1517 1 2 874 109 906 ICV_20 $T=201020 383520 1 0 $X=200830 $Y=380560
X1518 1 2 901 109 928 ICV_20 $T=208380 410720 1 0 $X=208190 $Y=407760
X1519 1 2 931 109 939 ICV_20 $T=215280 432480 0 0 $X=215090 $Y=432240
X1520 1 2 146 126 149 ICV_20 $T=219420 378080 0 0 $X=219230 $Y=377840
X1521 1 2 927 111 985 ICV_20 $T=236440 383520 1 0 $X=236250 $Y=380560
X1522 1 2 969 111 989 ICV_20 $T=238740 399840 0 0 $X=238550 $Y=399600
X1523 1 2 969 125 1015 ICV_20 $T=250240 405280 0 0 $X=250050 $Y=405040
X1524 1 2 969 109 1017 ICV_20 $T=254380 405280 1 0 $X=254190 $Y=402320
X1525 1 2 1014 127 1018 ICV_20 $T=256680 427040 1 0 $X=256490 $Y=424080
X1526 1 2 984 113 1035 ICV_20 $T=260820 394400 1 0 $X=260630 $Y=391440
X1527 1 2 1014 113 1042 ICV_20 $T=264500 427040 1 0 $X=264310 $Y=424080
X1528 1 2 1041 113 1052 ICV_20 $T=271860 394400 0 0 $X=271670 $Y=394160
X1529 1 2 1050 126 1064 ICV_20 $T=276000 427040 0 0 $X=275810 $Y=426800
X1530 1 2 1041 112 1074 ICV_20 $T=280140 405280 1 0 $X=279950 $Y=402320
X1531 1 2 1041 125 1075 ICV_20 $T=281060 394400 1 0 $X=280870 $Y=391440
X1532 1 2 1076 113 1119 ICV_20 $T=302680 405280 1 0 $X=302490 $Y=402320
X1533 1 2 1104 126 1122 ICV_20 $T=303140 427040 1 0 $X=302950 $Y=424080
X1534 1 2 1104 113 1127 ICV_20 $T=306820 416160 1 0 $X=306630 $Y=413200
X1535 1 2 179 180 182 ICV_20 $T=308200 410720 1 0 $X=308010 $Y=407760
X1536 1 2 1128 185 1137 ICV_20 $T=314640 394400 0 0 $X=314450 $Y=394160
X1537 1 2 179 192 203 ICV_20 $T=318780 405280 0 0 $X=318590 $Y=405040
X1538 1 2 193 196 1147 ICV_20 $T=320620 443360 1 0 $X=320430 $Y=440400
X1539 1 2 1141 202 1151 ICV_20 $T=323840 410720 0 0 $X=323650 $Y=410480
X1540 1 2 1185 199 1194 ICV_20 $T=346840 427040 1 0 $X=346650 $Y=424080
X1541 1 2 241 184 1197 ICV_20 $T=348680 383520 1 0 $X=348490 $Y=380560
X1542 1 2 1167 219 1209 ICV_20 $T=354200 399840 0 0 $X=354010 $Y=399600
X1543 1 2 1185 213 1217 ICV_20 $T=356960 427040 1 0 $X=356770 $Y=424080
X1544 1 2 1185 228 1216 ICV_20 $T=356960 432480 1 0 $X=356770 $Y=429520
X1545 1 2 248 199 1218 ICV_20 $T=356960 443360 1 0 $X=356770 $Y=440400
X1546 1 2 1210 185 1224 ICV_20 $T=362020 399840 0 0 $X=361830 $Y=399600
X1547 1 2 241 211 1228 ICV_20 $T=362480 378080 0 0 $X=362290 $Y=377840
X1548 1 2 1210 211 1235 ICV_20 $T=365240 394400 1 0 $X=365050 $Y=391440
X1549 1 2 1211 224 1241 ICV_20 $T=368460 416160 1 0 $X=368270 $Y=413200
X1550 1 2 1210 219 1248 ICV_20 $T=373060 394400 1 0 $X=372870 $Y=391440
X1551 1 2 1259 213 1275 ICV_20 $T=385020 416160 1 0 $X=384830 $Y=413200
X1552 1 2 1282 185 1289 ICV_20 $T=395600 405280 1 0 $X=395410 $Y=402320
X1553 1 2 1300 211 1316 ICV_20 $T=407560 394400 0 0 $X=407370 $Y=394160
X1554 1 2 1321 204 1355 ICV_20 $T=426880 421600 0 0 $X=426690 $Y=421360
X1555 1 2 1340 212 1359 ICV_20 $T=428720 394400 0 0 $X=428530 $Y=394160
X1556 1 2 1377 189 1398 ICV_20 $T=448500 394400 1 0 $X=448310 $Y=391440
X1557 1 2 1377 184 1417 ICV_20 $T=459540 394400 0 0 $X=459350 $Y=394160
X1558 1 2 1377 190 1418 ICV_20 $T=460000 399840 1 0 $X=459810 $Y=396880
X1559 1 2 1431 196 1453 ICV_20 $T=476560 421600 1 0 $X=476370 $Y=418640
X1560 1 2 319 199 1458 ICV_20 $T=479780 443360 1 0 $X=479590 $Y=440400
X1561 1 2 324 211 1500 ICV_20 $T=501400 378080 0 0 $X=501210 $Y=377840
X1562 1 2 1456 211 1495 ICV_20 $T=501860 388960 0 0 $X=501670 $Y=388720
X1563 1 2 1483 202 1509 ICV_20 $T=511060 410720 0 0 $X=510870 $Y=410480
X1564 1 2 1517 360 1526 ICV_20 $T=525320 432480 1 0 $X=525130 $Y=429520
X1565 1 2 179 366 374 ICV_20 $T=529460 410720 0 0 $X=529270 $Y=410480
X1566 1 2 1540 357 1567 ICV_20 $T=556600 432480 1 0 $X=556410 $Y=429520
X1567 1 2 1539 365 1569 ICV_20 $T=557520 405280 0 0 $X=557330 $Y=405040
X1568 1 2 390 405 1573 ICV_20 $T=558900 378080 0 0 $X=558710 $Y=377840
X1569 1 2 1539 358 1576 ICV_20 $T=559360 416160 1 0 $X=559170 $Y=413200
X1570 1 2 1621 360 1635 ICV_20 $T=586960 432480 0 0 $X=586770 $Y=432240
X1571 1 2 1618 365 1639 ICV_20 $T=589720 405280 1 0 $X=589530 $Y=402320
X1572 1 2 1621 372 1657 ICV_20 $T=597540 432480 1 0 $X=597350 $Y=429520
X1573 1 2 418 357 1660 ICV_20 $T=598920 443360 1 0 $X=598730 $Y=440400
X1574 1 2 1641 400 1678 ICV_20 $T=609500 394400 1 0 $X=609310 $Y=391440
X1575 1 2 418 372 1684 ICV_20 $T=611340 443360 1 0 $X=611150 $Y=440400
X1576 1 2 1685 402 1708 ICV_20 $T=623300 394400 0 0 $X=623110 $Y=394160
X1577 1 2 1730 359 1748 ICV_20 $T=644000 416160 1 0 $X=643810 $Y=413200
X1578 1 2 1730 381 1750 ICV_20 $T=644920 405280 1 0 $X=644730 $Y=402320
X1579 1 2 1765 407 1780 ICV_20 $T=661940 383520 0 0 $X=661750 $Y=383280
X1580 1 2 1802 381 1827 ICV_20 $T=685400 427040 1 0 $X=685210 $Y=424080
X1581 1 2 1826 360 1831 ICV_20 $T=690920 410720 0 0 $X=690730 $Y=410480
X1582 1 2 1826 372 1832 ICV_20 $T=690920 416160 0 0 $X=690730 $Y=415920
X1583 1 2 1859 365 1867 ICV_20 $T=705180 432480 1 0 $X=704990 $Y=429520
X1584 1 2 1866 406 1892 ICV_20 $T=711160 394400 1 0 $X=710970 $Y=391440
X1585 1 2 604 9 617 ICV_21 $T=48300 427040 1 0 $X=48110 $Y=424080
X1586 1 2 597 11 656 ICV_21 $T=65320 388960 1 0 $X=65130 $Y=386000
X1587 1 2 665 28 690 ICV_21 $T=83720 427040 1 0 $X=83530 $Y=424080
X1588 1 2 695 29 738 ICV_21 $T=107180 394400 0 0 $X=106990 $Y=394160
X1589 1 2 135 112 880 ICV_21 $T=181700 378080 0 0 $X=181510 $Y=377840
X1590 1 2 855 113 925 ICV_21 $T=202400 399840 0 0 $X=202210 $Y=399600
X1591 1 2 1141 204 1155 ICV_21 $T=322000 416160 0 0 $X=321810 $Y=415920
X1592 1 2 1167 189 1198 ICV_21 $T=345920 394400 1 0 $X=345730 $Y=391440
X1593 1 2 1286 204 1304 ICV_21 $T=398820 427040 0 0 $X=398630 $Y=426800
X1594 1 2 1407 196 1425 ICV_21 $T=459080 416160 0 0 $X=458890 $Y=415920
X1595 1 2 1431 202 1466 ICV_21 $T=483000 410720 0 0 $X=482810 $Y=410480
X1596 1 2 1621 365 1636 ICV_21 $T=585580 427040 1 0 $X=585390 $Y=424080
X1597 1 2 1721 406 1740 ICV_21 $T=637560 388960 1 0 $X=637370 $Y=386000
X1598 1 2 1765 405 1779 ICV_21 $T=658720 394400 0 0 $X=658530 $Y=394160
X1599 1 2 1802 357 1811 ICV_21 $T=674820 427040 1 0 $X=674630 $Y=424080
X1600 1 2 1866 407 1915 ICV_21 $T=722200 394400 0 0 $X=722010 $Y=394160
X1601 1 2 513 30 560 557 521 34 ICV_22 $T=18400 399840 0 0 $X=18210 $Y=399600
X1602 1 2 879 127 898 897 890 123 ICV_22 $T=188600 432480 1 0 $X=188410 $Y=429520
X1603 1 2 932 124 942 942 949 128 ICV_22 $T=214360 421600 0 0 $X=214170 $Y=421360
X1604 1 2 146 112 155 963 951 131 ICV_22 $T=230460 378080 0 0 $X=230270 $Y=377840
X1605 1 2 146 109 1007 1007 158 118 ICV_22 $T=244260 378080 0 0 $X=244070 $Y=377840
X1606 1 2 965 113 1011 1011 980 122 ICV_22 $T=244720 421600 1 0 $X=244530 $Y=418640
X1607 1 2 1072 126 1091 1091 1092 130 ICV_22 $T=286580 383520 0 0 $X=286390 $Y=383280
X1608 1 2 1076 127 1118 1117 1097 119 ICV_22 $T=300840 399840 1 0 $X=300650 $Y=396880
X1609 1 2 254 185 1273 1273 259 205 ICV_22 $T=383180 378080 0 0 $X=382990 $Y=377840
X1610 1 2 1427 191 1441 1440 1443 205 ICV_22 $T=469200 405280 1 0 $X=469010 $Y=402320
X1611 1 2 1431 199 1465 1465 1447 183 ICV_22 $T=483000 416160 0 0 $X=482810 $Y=415920
X1612 1 2 1519 378 1534 1537 1516 343 ICV_22 $T=534980 421600 1 0 $X=534790 $Y=418640
X1613 1 2 1585 372 1609 1609 1597 371 ICV_22 $T=571320 416160 0 0 $X=571130 $Y=415920
X1614 1 2 1621 381 1656 1656 1638 345 ICV_22 $T=595240 421600 0 0 $X=595050 $Y=421360
X1615 1 2 1671 359 1683 1682 1690 343 ICV_22 $T=609500 437920 1 0 $X=609310 $Y=434960
X1616 1 2 1784 403 453 1822 447 389 ICV_22 $T=679420 383520 0 0 $X=679230 $Y=383280
X1617 1 2 1826 358 1854 1854 1842 368 ICV_22 $T=693680 416160 1 0 $X=693490 $Y=413200
X1618 1 2 1864 357 1894 1894 1869 367 ICV_22 $T=719440 405280 0 0 $X=719250 $Y=405040
X1619 1 2 1859 358 1901 1901 1874 368 ICV_22 $T=720360 427040 0 0 $X=720170 $Y=426800
X1620 1 2 ICV_23 $T=18400 432480 1 0 $X=18210 $Y=429520
X1621 1 2 ICV_23 $T=18400 437920 1 0 $X=18210 $Y=434960
X1622 1 2 ICV_23 $T=32200 399840 0 0 $X=32010 $Y=399600
X1623 1 2 ICV_23 $T=32200 416160 0 0 $X=32010 $Y=415920
X1624 1 2 ICV_23 $T=74520 443360 1 0 $X=74330 $Y=440400
X1625 1 2 ICV_23 $T=88320 437920 0 0 $X=88130 $Y=437680
X1626 1 2 ICV_23 $T=130640 416160 1 0 $X=130450 $Y=413200
X1627 1 2 ICV_23 $T=172500 405280 0 0 $X=172310 $Y=405040
X1628 1 2 ICV_23 $T=172500 410720 0 0 $X=172310 $Y=410480
X1629 1 2 ICV_23 $T=172500 416160 0 0 $X=172310 $Y=415920
X1630 1 2 ICV_23 $T=186760 421600 1 0 $X=186570 $Y=418640
X1631 1 2 ICV_23 $T=200560 421600 0 0 $X=200370 $Y=421360
X1632 1 2 ICV_23 $T=228620 416160 0 0 $X=228430 $Y=415920
X1633 1 2 ICV_23 $T=242880 421600 1 0 $X=242690 $Y=418640
X1634 1 2 ICV_23 $T=256680 416160 0 0 $X=256490 $Y=415920
X1635 1 2 ICV_23 $T=270940 416160 1 0 $X=270750 $Y=413200
X1636 1 2 ICV_23 $T=284740 405280 0 0 $X=284550 $Y=405040
X1637 1 2 ICV_23 $T=299000 416160 1 0 $X=298810 $Y=413200
X1638 1 2 ICV_23 $T=299000 421600 1 0 $X=298810 $Y=418640
X1639 1 2 ICV_23 $T=327060 421600 1 0 $X=326870 $Y=418640
X1640 1 2 ICV_23 $T=368920 416160 0 0 $X=368730 $Y=415920
X1641 1 2 ICV_23 $T=425040 378080 0 0 $X=424850 $Y=377840
X1642 1 2 ICV_23 $T=453100 405280 0 0 $X=452910 $Y=405040
X1643 1 2 ICV_23 $T=453100 427040 0 0 $X=452910 $Y=426800
X1644 1 2 ICV_23 $T=467360 394400 1 0 $X=467170 $Y=391440
X1645 1 2 ICV_23 $T=481160 399840 0 0 $X=480970 $Y=399600
X1646 1 2 ICV_23 $T=495420 405280 1 0 $X=495230 $Y=402320
X1647 1 2 ICV_23 $T=509220 432480 0 0 $X=509030 $Y=432240
X1648 1 2 ICV_23 $T=523480 399840 1 0 $X=523290 $Y=396880
X1649 1 2 ICV_23 $T=523480 421600 1 0 $X=523290 $Y=418640
X1650 1 2 ICV_23 $T=537280 405280 0 0 $X=537090 $Y=405040
X1651 1 2 ICV_23 $T=537280 410720 0 0 $X=537090 $Y=410480
X1652 1 2 ICV_23 $T=537280 427040 0 0 $X=537090 $Y=426800
X1653 1 2 ICV_23 $T=551540 437920 1 0 $X=551350 $Y=434960
X1654 1 2 ICV_23 $T=565340 405280 0 0 $X=565150 $Y=405040
X1655 1 2 ICV_23 $T=579600 399840 1 0 $X=579410 $Y=396880
X1656 1 2 ICV_23 $T=593400 399840 0 0 $X=593210 $Y=399600
X1657 1 2 ICV_23 $T=607660 394400 1 0 $X=607470 $Y=391440
X1658 1 2 ICV_23 $T=621460 394400 0 0 $X=621270 $Y=394160
X1659 1 2 ICV_23 $T=635720 388960 1 0 $X=635530 $Y=386000
X1660 1 2 ICV_23 $T=635720 432480 1 0 $X=635530 $Y=429520
X1661 1 2 ICV_23 $T=635720 437920 1 0 $X=635530 $Y=434960
X1662 1 2 ICV_23 $T=663780 383520 1 0 $X=663590 $Y=380560
X1663 1 2 ICV_23 $T=663780 394400 1 0 $X=663590 $Y=391440
X1664 1 2 ICV_23 $T=677580 416160 0 0 $X=677390 $Y=415920
X1665 1 2 ICV_23 $T=691840 394400 1 0 $X=691650 $Y=391440
X1666 1 2 ICV_23 $T=733700 416160 0 0 $X=733510 $Y=415920
X1667 1 2 ICV_24 $T=46000 427040 1 0 $X=45810 $Y=424080
X1668 1 2 ICV_24 $T=46000 443360 1 0 $X=45810 $Y=440400
X1669 1 2 ICV_24 $T=74060 383520 1 0 $X=73870 $Y=380560
X1670 1 2 ICV_24 $T=102120 405280 1 0 $X=101930 $Y=402320
X1671 1 2 ICV_24 $T=102120 437920 1 0 $X=101930 $Y=434960
X1672 1 2 ICV_24 $T=115920 416160 0 0 $X=115730 $Y=415920
X1673 1 2 ICV_24 $T=200100 388960 0 0 $X=199910 $Y=388720
X1674 1 2 ICV_24 $T=228160 421600 0 0 $X=227970 $Y=421360
X1675 1 2 ICV_24 $T=326600 388960 1 0 $X=326410 $Y=386000
X1676 1 2 ICV_24 $T=340400 405280 0 0 $X=340210 $Y=405040
X1677 1 2 ICV_24 $T=354660 427040 1 0 $X=354470 $Y=424080
X1678 1 2 ICV_24 $T=368460 405280 0 0 $X=368270 $Y=405040
X1679 1 2 ICV_24 $T=480700 383520 0 0 $X=480510 $Y=383280
X1680 1 2 ICV_24 $T=551080 405280 1 0 $X=550890 $Y=402320
X1681 1 2 ICV_24 $T=564880 432480 0 0 $X=564690 $Y=432240
X1682 1 2 ICV_24 $T=579140 394400 1 0 $X=578950 $Y=391440
X1683 1 2 ICV_24 $T=592940 394400 0 0 $X=592750 $Y=394160
X1684 1 2 ICV_24 $T=592940 410720 0 0 $X=592750 $Y=410480
X1685 1 2 ICV_24 $T=607200 432480 1 0 $X=607010 $Y=429520
X1686 1 2 ICV_24 $T=649060 432480 0 0 $X=648870 $Y=432240
X1687 1 2 ICV_24 $T=705180 421600 0 0 $X=704990 $Y=421360
X1688 1 2 ICV_24 $T=719440 427040 1 0 $X=719250 $Y=424080
X1689 1 2 ICV_24 $T=733240 405280 0 0 $X=733050 $Y=405040
X1690 1 2 ICV_24 $T=733240 421600 0 0 $X=733050 $Y=421360
X1691 1 2 26 2 20 1 sky130_fd_sc_hd__inv_1 $T=18400 443360 1 0 $X=18210 $Y=440400
X1692 1 2 7 2 534 1 sky130_fd_sc_hd__inv_1 $T=22540 416160 0 0 $X=22350 $Y=415920
X1693 1 2 6 2 543 1 sky130_fd_sc_hd__inv_1 $T=24380 378080 0 0 $X=24190 $Y=377840
X1694 1 2 12 2 521 1 sky130_fd_sc_hd__inv_1 $T=28520 394400 0 0 $X=28330 $Y=394160
X1695 1 2 22 2 533 1 sky130_fd_sc_hd__inv_1 $T=31280 421600 0 0 $X=31090 $Y=421360
X1696 1 2 40 2 43 1 sky130_fd_sc_hd__inv_1 $T=45540 437920 1 0 $X=45350 $Y=434960
X1697 1 2 42 2 554 1 sky130_fd_sc_hd__inv_1 $T=46460 421600 1 0 $X=46270 $Y=418640
X1698 1 2 32 2 576 1 sky130_fd_sc_hd__inv_1 $T=48300 405280 1 0 $X=48110 $Y=402320
X1699 1 2 50 2 605 1 sky130_fd_sc_hd__inv_1 $T=60260 394400 0 0 $X=60070 $Y=394160
X1700 1 2 53 2 51 1 sky130_fd_sc_hd__inv_1 $T=64400 383520 1 0 $X=64210 $Y=380560
X1701 1 2 62 2 58 1 sky130_fd_sc_hd__inv_1 $T=83260 437920 0 0 $X=83070 $Y=437680
X1702 1 2 60 2 648 1 sky130_fd_sc_hd__inv_1 $T=86940 399840 0 0 $X=86750 $Y=399600
X1703 1 2 55 2 634 1 sky130_fd_sc_hd__inv_1 $T=88320 388960 0 0 $X=88130 $Y=388720
X1704 1 2 65 2 683 1 sky130_fd_sc_hd__inv_1 $T=100740 405280 1 0 $X=100550 $Y=402320
X1705 1 2 76 2 673 1 sky130_fd_sc_hd__inv_1 $T=107180 416160 0 0 $X=106990 $Y=415920
X1706 1 2 73 2 66 1 sky130_fd_sc_hd__inv_1 $T=111780 383520 1 0 $X=111590 $Y=380560
X1707 1 2 72 2 71 1 sky130_fd_sc_hd__inv_1 $T=118220 437920 0 0 $X=118030 $Y=437680
X1708 1 2 86 2 732 1 sky130_fd_sc_hd__inv_1 $T=118680 421600 0 0 $X=118490 $Y=421360
X1709 1 2 80 2 88 1 sky130_fd_sc_hd__inv_1 $T=118680 443360 1 0 $X=118490 $Y=440400
X1710 1 2 69 2 716 1 sky130_fd_sc_hd__inv_1 $T=122820 394400 0 0 $X=122630 $Y=394160
X1711 1 2 77 2 720 1 sky130_fd_sc_hd__inv_1 $T=124660 410720 1 0 $X=124470 $Y=407760
X1712 1 2 82 2 758 1 sky130_fd_sc_hd__inv_1 $T=138460 388960 0 0 $X=138270 $Y=388720
X1713 1 2 93 2 773 1 sky130_fd_sc_hd__inv_1 $T=143060 399840 0 0 $X=142870 $Y=399600
X1714 1 2 97 2 87 1 sky130_fd_sc_hd__inv_1 $T=143980 437920 0 0 $X=143790 $Y=437680
X1715 1 2 81 2 768 1 sky130_fd_sc_hd__inv_1 $T=146280 432480 0 0 $X=146090 $Y=432240
X1716 1 2 7 2 819 1 sky130_fd_sc_hd__inv_1 $T=157780 421600 1 0 $X=157590 $Y=418640
X1717 1 2 50 2 802 1 sky130_fd_sc_hd__inv_1 $T=160540 388960 1 0 $X=160350 $Y=386000
X1718 1 2 60 2 798 1 sky130_fd_sc_hd__inv_1 $T=166060 394400 1 0 $X=165870 $Y=391440
X1719 1 2 40 2 120 1 sky130_fd_sc_hd__inv_1 $T=167900 437920 1 0 $X=167710 $Y=434960
X1720 1 2 6 2 116 1 sky130_fd_sc_hd__inv_1 $T=172040 378080 0 0 $X=171850 $Y=377840
X1721 1 2 22 2 844 1 sky130_fd_sc_hd__inv_1 $T=172500 427040 0 0 $X=172310 $Y=426800
X1722 1 2 32 2 809 1 sky130_fd_sc_hd__inv_1 $T=174800 410720 1 0 $X=174610 $Y=407760
X1723 1 2 12 2 873 1 sky130_fd_sc_hd__inv_1 $T=188140 394400 0 0 $X=187950 $Y=394160
X1724 1 2 46 2 890 1 sky130_fd_sc_hd__inv_1 $T=196420 427040 1 0 $X=196230 $Y=424080
X1725 1 2 57 2 845 1 sky130_fd_sc_hd__inv_1 $T=196880 405280 1 0 $X=196690 $Y=402320
X1726 1 2 42 2 854 1 sky130_fd_sc_hd__inv_1 $T=199180 421600 0 0 $X=198990 $Y=421360
X1727 1 2 39 2 888 1 sky130_fd_sc_hd__inv_1 $T=199640 378080 0 0 $X=199450 $Y=377840
X1728 1 2 136 2 140 1 sky130_fd_sc_hd__inv_1 $T=215280 437920 0 0 $X=215090 $Y=437680
X1729 1 2 47 2 918 1 sky130_fd_sc_hd__inv_1 $T=222640 405280 1 0 $X=222450 $Y=402320
X1730 1 2 55 2 936 1 sky130_fd_sc_hd__inv_1 $T=228620 388960 0 0 $X=228430 $Y=388720
X1731 1 2 77 2 949 1 sky130_fd_sc_hd__inv_1 $T=230460 410720 0 0 $X=230270 $Y=410480
X1732 1 2 65 2 147 1 sky130_fd_sc_hd__inv_1 $T=230460 427040 0 0 $X=230270 $Y=426800
X1733 1 2 151 2 980 1 sky130_fd_sc_hd__inv_1 $T=241960 410720 1 0 $X=241770 $Y=407760
X1734 1 2 153 2 976 1 sky130_fd_sc_hd__inv_1 $T=256220 427040 0 0 $X=256030 $Y=426800
X1735 1 2 150 2 990 1 sky130_fd_sc_hd__inv_1 $T=262200 405280 1 0 $X=262010 $Y=402320
X1736 1 2 101 2 1019 1 sky130_fd_sc_hd__inv_1 $T=270480 427040 0 0 $X=270290 $Y=426800
X1737 1 2 166 2 165 1 sky130_fd_sc_hd__inv_1 $T=270940 383520 1 0 $X=270750 $Y=380560
X1738 1 2 97 2 1008 1 sky130_fd_sc_hd__inv_1 $T=270940 394400 1 0 $X=270750 $Y=391440
X1739 1 2 156 2 162 1 sky130_fd_sc_hd__inv_1 $T=276000 437920 1 0 $X=275810 $Y=434960
X1740 1 2 163 2 1038 1 sky130_fd_sc_hd__inv_1 $T=283820 410720 0 0 $X=283630 $Y=410480
X1741 1 2 62 2 1067 1 sky130_fd_sc_hd__inv_1 $T=283820 427040 0 0 $X=283630 $Y=426800
X1742 1 2 80 2 1053 1 sky130_fd_sc_hd__inv_1 $T=286580 394400 0 0 $X=286390 $Y=394160
X1743 1 2 177 2 1102 1 sky130_fd_sc_hd__inv_1 $T=299000 437920 1 0 $X=298810 $Y=434960
X1744 1 2 82 2 1097 1 sky130_fd_sc_hd__inv_1 $T=300840 394400 0 0 $X=300650 $Y=394160
X1745 1 2 100 2 1107 1 sky130_fd_sc_hd__inv_1 $T=305440 421600 0 0 $X=305250 $Y=421360
X1746 1 2 81 2 176 1 sky130_fd_sc_hd__inv_1 $T=309580 443360 1 0 $X=309390 $Y=440400
X1747 1 2 226 2 214 1 sky130_fd_sc_hd__inv_1 $T=333500 378080 0 0 $X=333310 $Y=377840
X1748 1 2 223 2 1144 1 sky130_fd_sc_hd__inv_1 $T=336260 394400 1 0 $X=336070 $Y=391440
X1749 1 2 233 2 217 1 sky130_fd_sc_hd__inv_1 $T=340400 383520 0 0 $X=340210 $Y=383280
X1750 1 2 247 2 1183 1 sky130_fd_sc_hd__inv_1 $T=360180 405280 0 0 $X=359990 $Y=405040
X1751 1 2 245 2 1168 1 sky130_fd_sc_hd__inv_1 $T=361100 399840 1 0 $X=360910 $Y=396880
X1752 1 2 240 2 1199 1 sky130_fd_sc_hd__inv_1 $T=367540 416160 0 0 $X=367350 $Y=415920
X1753 1 2 249 2 251 1 sky130_fd_sc_hd__inv_1 $T=372140 437920 1 0 $X=371950 $Y=434960
X1754 1 2 252 2 1207 1 sky130_fd_sc_hd__inv_1 $T=373520 383520 1 0 $X=373330 $Y=380560
X1755 1 2 253 2 1225 1 sky130_fd_sc_hd__inv_1 $T=377200 399840 1 0 $X=377010 $Y=396880
X1756 1 2 250 2 1239 1 sky130_fd_sc_hd__inv_1 $T=382260 410720 1 0 $X=382070 $Y=407760
X1757 1 2 255 2 1223 1 sky130_fd_sc_hd__inv_1 $T=382260 427040 0 0 $X=382070 $Y=426800
X1758 1 2 260 2 1274 1 sky130_fd_sc_hd__inv_1 $T=396980 410720 0 0 $X=396790 $Y=410480
X1759 1 2 270 2 1290 1 sky130_fd_sc_hd__inv_1 $T=406180 394400 0 0 $X=405990 $Y=394160
X1760 1 2 263 2 264 1 sky130_fd_sc_hd__inv_1 $T=406180 432480 0 0 $X=405990 $Y=432240
X1761 1 2 274 2 1305 1 sky130_fd_sc_hd__inv_1 $T=411240 410720 1 0 $X=411050 $Y=407760
X1762 1 2 278 2 1317 1 sky130_fd_sc_hd__inv_1 $T=426880 399840 0 0 $X=426690 $Y=399600
X1763 1 2 279 2 276 1 sky130_fd_sc_hd__inv_1 $T=426880 437920 0 0 $X=426690 $Y=437680
X1764 1 2 275 2 1323 1 sky130_fd_sc_hd__inv_1 $T=427340 427040 1 0 $X=427150 $Y=424080
X1765 1 2 284 2 1334 1 sky130_fd_sc_hd__inv_1 $T=431480 405280 0 0 $X=431290 $Y=405040
X1766 1 2 285 2 282 1 sky130_fd_sc_hd__inv_1 $T=438840 388960 1 0 $X=438650 $Y=386000
X1767 1 2 291 2 1371 1 sky130_fd_sc_hd__inv_1 $T=451720 427040 0 0 $X=451530 $Y=426800
X1768 1 2 300 2 295 1 sky130_fd_sc_hd__inv_1 $T=457240 394400 1 0 $X=457050 $Y=391440
X1769 1 2 301 2 1380 1 sky130_fd_sc_hd__inv_1 $T=459080 410720 0 0 $X=458890 $Y=410480
X1770 1 2 302 2 1399 1 sky130_fd_sc_hd__inv_1 $T=459540 399840 0 0 $X=459350 $Y=399600
X1771 1 2 308 2 305 1 sky130_fd_sc_hd__inv_1 $T=467360 437920 0 0 $X=467170 $Y=437680
X1772 1 2 314 2 312 1 sky130_fd_sc_hd__inv_1 $T=472880 378080 0 0 $X=472690 $Y=377840
X1773 1 2 304 2 1403 1 sky130_fd_sc_hd__inv_1 $T=473340 410720 1 0 $X=473150 $Y=407760
X1774 1 2 320 2 1443 1 sky130_fd_sc_hd__inv_1 $T=483000 399840 0 0 $X=482810 $Y=399600
X1775 1 2 318 2 322 1 sky130_fd_sc_hd__inv_1 $T=487140 432480 0 0 $X=486950 $Y=432240
X1776 1 2 315 2 1447 1 sky130_fd_sc_hd__inv_1 $T=493580 410720 0 0 $X=493390 $Y=410480
X1777 1 2 334 2 323 1 sky130_fd_sc_hd__inv_1 $T=506920 399840 0 0 $X=506730 $Y=399600
X1778 1 2 338 2 1487 1 sky130_fd_sc_hd__inv_1 $T=509220 427040 0 0 $X=509030 $Y=426800
X1779 1 2 333 2 326 1 sky130_fd_sc_hd__inv_1 $T=511060 383520 0 0 $X=510870 $Y=383280
X1780 1 2 335 2 336 1 sky130_fd_sc_hd__inv_1 $T=522560 432480 0 0 $X=522370 $Y=432240
X1781 1 2 328 2 1480 1 sky130_fd_sc_hd__inv_1 $T=523480 410720 1 0 $X=523290 $Y=407760
X1782 1 2 235 2 1527 1 sky130_fd_sc_hd__inv_1 $T=533140 432480 1 0 $X=532950 $Y=429520
X1783 1 2 240 2 1516 1 sky130_fd_sc_hd__inv_1 $T=533600 421600 1 0 $X=533410 $Y=418640
X1784 1 2 233 2 398 1 sky130_fd_sc_hd__inv_1 $T=551540 383520 1 0 $X=551350 $Y=380560
X1785 1 2 247 2 1545 1 sky130_fd_sc_hd__inv_1 $T=551540 410720 1 0 $X=551350 $Y=407760
X1786 1 2 384 2 401 1 sky130_fd_sc_hd__inv_1 $T=553840 437920 0 0 $X=553650 $Y=437680
X1787 1 2 223 2 1553 1 sky130_fd_sc_hd__inv_1 $T=554300 394400 1 0 $X=554110 $Y=391440
X1788 1 2 253 2 1586 1 sky130_fd_sc_hd__inv_1 $T=570860 399840 1 0 $X=570670 $Y=396880
X1789 1 2 255 2 1589 1 sky130_fd_sc_hd__inv_1 $T=571780 427040 0 0 $X=571590 $Y=426800
X1790 1 2 285 2 1590 1 sky130_fd_sc_hd__inv_1 $T=572240 388960 1 0 $X=572050 $Y=386000
X1791 1 2 260 2 1597 1 sky130_fd_sc_hd__inv_1 $T=575000 405280 1 0 $X=574810 $Y=402320
X1792 1 2 250 2 1637 1 sky130_fd_sc_hd__inv_1 $T=595240 405280 0 0 $X=595050 $Y=405040
X1793 1 2 279 2 1643 1 sky130_fd_sc_hd__inv_1 $T=597540 443360 1 0 $X=597350 $Y=440400
X1794 1 2 249 2 1638 1 sky130_fd_sc_hd__inv_1 $T=605820 432480 1 0 $X=605630 $Y=429520
X1795 1 2 245 2 1655 1 sky130_fd_sc_hd__inv_1 $T=609040 399840 0 0 $X=608850 $Y=399600
X1796 1 2 284 2 1667 1 sky130_fd_sc_hd__inv_1 $T=609500 410720 1 0 $X=609310 $Y=407760
X1797 1 2 270 2 422 1 sky130_fd_sc_hd__inv_1 $T=613180 383520 0 0 $X=612990 $Y=383280
X1798 1 2 274 2 1689 1 sky130_fd_sc_hd__inv_1 $T=624220 416160 1 0 $X=624030 $Y=413200
X1799 1 2 275 2 1690 1 sky130_fd_sc_hd__inv_1 $T=625140 427040 1 0 $X=624950 $Y=424080
X1800 1 2 256 2 1707 1 sky130_fd_sc_hd__inv_1 $T=631120 394400 0 0 $X=630930 $Y=394160
X1801 1 2 351 2 435 1 sky130_fd_sc_hd__inv_1 $T=640780 378080 0 0 $X=640590 $Y=377840
X1802 1 2 263 2 434 1 sky130_fd_sc_hd__inv_1 $T=644920 427040 1 0 $X=644730 $Y=424080
X1803 1 2 292 2 1728 1 sky130_fd_sc_hd__inv_1 $T=648600 399840 0 0 $X=648410 $Y=399600
X1804 1 2 304 2 1754 1 sky130_fd_sc_hd__inv_1 $T=653200 405280 0 0 $X=653010 $Y=405040
X1805 1 2 278 2 1770 1 sky130_fd_sc_hd__inv_1 $T=663780 399840 1 0 $X=663590 $Y=396880
X1806 1 2 318 2 440 1 sky130_fd_sc_hd__inv_1 $T=663780 432480 1 0 $X=663590 $Y=429520
X1807 1 2 291 2 1772 1 sky130_fd_sc_hd__inv_1 $T=675280 421600 0 0 $X=675090 $Y=421360
X1808 1 2 302 2 448 1 sky130_fd_sc_hd__inv_1 $T=676200 378080 0 0 $X=676010 $Y=377840
X1809 1 2 300 2 447 1 sky130_fd_sc_hd__inv_1 $T=678960 394400 1 0 $X=678770 $Y=391440
X1810 1 2 308 2 1804 1 sky130_fd_sc_hd__inv_1 $T=679420 437920 1 0 $X=679230 $Y=434960
X1811 1 2 335 2 1810 1 sky130_fd_sc_hd__inv_1 $T=686780 427040 0 0 $X=686590 $Y=426800
X1812 1 2 314 2 457 1 sky130_fd_sc_hd__inv_1 $T=692300 378080 0 0 $X=692110 $Y=377840
X1813 1 2 315 2 1842 1 sky130_fd_sc_hd__inv_1 $T=701960 410720 1 0 $X=701770 $Y=407760
X1814 1 2 301 2 1869 1 sky130_fd_sc_hd__inv_1 $T=718060 405280 0 0 $X=717870 $Y=405040
X1815 1 2 330 2 1885 1 sky130_fd_sc_hd__inv_1 $T=718980 388960 1 0 $X=718790 $Y=386000
X1816 1 2 311 2 1878 1 sky130_fd_sc_hd__inv_1 $T=718980 421600 0 0 $X=718790 $Y=421360
X1817 1 2 338 2 1874 1 sky130_fd_sc_hd__inv_1 $T=718980 427040 0 0 $X=718790 $Y=426800
X1818 1 2 334 2 1865 1 sky130_fd_sc_hd__inv_1 $T=719900 399840 1 0 $X=719710 $Y=396880
X1819 1 2 617 615 25 ICV_26 $T=58880 427040 1 0 $X=58690 $Y=424080
X1820 1 2 645 634 16 ICV_26 $T=71300 399840 1 0 $X=71110 $Y=396880
X1821 1 2 642 644 25 ICV_26 $T=71300 427040 1 0 $X=71110 $Y=424080
X1822 1 2 657 648 37 ICV_26 $T=76360 410720 0 0 $X=76170 $Y=410480
X1823 1 2 743 716 25 ICV_26 $T=118220 394400 0 0 $X=118030 $Y=394160
X1824 1 2 800 802 122 ICV_26 $T=153640 383520 0 0 $X=153450 $Y=383280
X1825 1 2 808 798 118 ICV_26 $T=155480 394400 1 0 $X=155290 $Y=391440
X1826 1 2 824 802 129 ICV_26 $T=165600 383520 0 0 $X=165410 $Y=383280
X1827 1 2 829 809 130 ICV_26 $T=167900 410720 0 0 $X=167710 $Y=410480
X1828 1 2 842 845 129 ICV_26 $T=172040 399840 1 0 $X=171850 $Y=396880
X1829 1 2 856 844 131 ICV_26 $T=181240 427040 1 0 $X=181050 $Y=424080
X1830 1 2 872 854 119 ICV_26 $T=183540 410720 1 0 $X=183350 $Y=407760
X1831 1 2 907 918 130 ICV_26 $T=209300 416160 1 0 $X=209110 $Y=413200
X1832 1 2 928 918 118 ICV_26 $T=216660 405280 1 0 $X=216470 $Y=402320
X1833 1 2 955 147 128 ICV_26 $T=228160 432480 1 0 $X=227970 $Y=429520
X1834 1 2 988 990 128 ICV_26 $T=245640 405280 0 0 $X=245450 $Y=405040
X1835 1 2 1018 1019 131 ICV_26 $T=260820 421600 0 0 $X=260630 $Y=421360
X1836 1 2 1068 171 122 ICV_26 $T=283820 383520 1 0 $X=283630 $Y=380560
X1837 1 2 1074 1053 119 ICV_26 $T=286580 399840 0 0 $X=286390 $Y=399600
X1838 1 2 1181 1183 192 ICV_26 $T=345460 405280 1 0 $X=345270 $Y=402320
X1839 1 2 1209 1168 237 ICV_26 $T=359260 405280 1 0 $X=359070 $Y=402320
X1840 1 2 262 264 188 ICV_26 $T=391460 437920 0 0 $X=391270 $Y=437680
X1841 1 2 1398 1399 209 ICV_26 $T=454940 394400 0 0 $X=454750 $Y=394160
X1842 1 2 1393 1380 195 ICV_26 $T=454940 421600 0 0 $X=454750 $Y=421360
X1843 1 2 1406 305 187 ICV_26 $T=460920 443360 1 0 $X=460730 $Y=440400
X1844 1 2 1425 1403 195 ICV_26 $T=469660 416160 0 0 $X=469470 $Y=415920
X1845 1 2 1452 323 221 ICV_26 $T=483000 388960 0 0 $X=482810 $Y=388720
X1846 1 2 1558 1553 387 ICV_26 $T=555680 394400 1 0 $X=555490 $Y=391440
X1847 1 2 1559 1545 355 ICV_26 $T=555680 416160 0 0 $X=555490 $Y=415920
X1848 1 2 419 420 355 ICV_26 $T=592940 443360 1 0 $X=592750 $Y=440400
X1849 1 2 1833 1804 367 ICV_26 $T=699660 437920 0 0 $X=699470 $Y=437680
X1850 1 2 1849 1851 387 ICV_26 $T=702420 388960 0 0 $X=702230 $Y=388720
X1851 1 2 1852 1851 352 ICV_26 $T=703340 394400 1 0 $X=703150 $Y=391440
X1852 1 2 515 13 535 ICV_28 $T=6900 421600 1 0 $X=6710 $Y=418640
X1853 1 2 637 28 658 ICV_28 $T=68540 388960 0 0 $X=68350 $Y=388720
X1854 1 2 676 11 687 ICV_28 $T=83720 410720 1 0 $X=83530 $Y=407760
X1855 1 2 68 10 706 ICV_28 $T=92460 383520 1 0 $X=92270 $Y=380560
X1856 1 2 665 10 677 ICV_28 $T=94300 427040 1 0 $X=94110 $Y=424080
X1857 1 2 695 28 713 ICV_28 $T=97520 399840 0 0 $X=97330 $Y=399600
X1858 1 2 711 10 731 ICV_28 $T=104420 427040 1 0 $X=104230 $Y=424080
X1859 1 2 746 11 782 ICV_28 $T=132480 388960 1 0 $X=132290 $Y=386000
X1860 1 2 108 112 814 ICV_28 $T=147660 432480 0 0 $X=147470 $Y=432240
X1861 1 2 132 127 856 ICV_28 $T=172040 427040 1 0 $X=171850 $Y=424080
X1862 1 2 931 124 955 ICV_28 $T=220800 427040 0 0 $X=220610 $Y=426800
X1863 1 2 965 109 981 ICV_28 $T=233680 421600 1 0 $X=233490 $Y=418640
X1864 1 2 1014 109 1029 ICV_28 $T=257140 432480 1 0 $X=256950 $Y=429520
X1865 1 2 172 127 1090 ICV_28 $T=286580 437920 0 0 $X=286390 $Y=437680
X1866 1 2 172 113 1095 ICV_28 $T=287960 443360 1 0 $X=287770 $Y=440400
X1867 1 2 179 188 198 ICV_28 $T=314640 410720 0 0 $X=314450 $Y=410480
X1868 1 2 1141 199 1153 ICV_28 $T=322000 421600 0 0 $X=321810 $Y=421360
X1869 1 2 179 220 234 ICV_28 $T=328900 410720 1 0 $X=328710 $Y=407760
X1870 1 2 179 239 243 ICV_28 $T=342700 405280 0 0 $X=342510 $Y=405040
X1871 1 2 1210 189 1230 ICV_28 $T=361100 388960 0 0 $X=360910 $Y=388720
X1872 1 2 1300 212 1315 ICV_28 $T=406180 388960 0 0 $X=405990 $Y=388720
X1873 1 2 1306 199 1319 ICV_28 $T=407560 432480 0 0 $X=407370 $Y=432240
X1874 1 2 277 190 1331 ICV_28 $T=413080 388960 1 0 $X=412890 $Y=386000
X1875 1 2 277 191 1345 ICV_28 $T=422280 388960 1 0 $X=422090 $Y=386000
X1876 1 2 1353 199 1369 ICV_28 $T=434240 427040 0 0 $X=434050 $Y=426800
X1877 1 2 1353 196 1370 ICV_28 $T=434240 432480 0 0 $X=434050 $Y=432240
X1878 1 2 286 224 1384 ICV_28 $T=441140 443360 1 0 $X=440950 $Y=440400
X1879 1 2 293 189 299 ICV_28 $T=448500 383520 1 0 $X=448310 $Y=380560
X1880 1 2 1431 227 1448 ICV_28 $T=473340 410720 0 0 $X=473150 $Y=410480
X1881 1 2 1456 219 1474 ICV_28 $T=486680 399840 1 0 $X=486490 $Y=396880
X1882 1 2 319 202 1479 ICV_28 $T=487600 443360 1 0 $X=487410 $Y=440400
X1883 1 2 1539 360 1555 ICV_28 $T=546480 416160 0 0 $X=546290 $Y=415920
X1884 1 2 1587 400 1626 ICV_28 $T=583740 394400 0 0 $X=583550 $Y=394160
X1885 1 2 1618 360 1632 ICV_28 $T=585120 416160 0 0 $X=584930 $Y=415920
X1886 1 2 1671 381 1692 ICV_28 $T=612260 427040 0 0 $X=612070 $Y=426800
X1887 1 2 1685 407 1700 ICV_28 $T=617320 394400 1 0 $X=617130 $Y=391440
X1888 1 2 1721 400 1756 ICV_28 $T=648140 388960 1 0 $X=647950 $Y=386000
X1889 1 2 1777 358 1791 ICV_28 $T=665620 410720 1 0 $X=665430 $Y=407760
X1890 1 2 1751 359 1793 ICV_28 $T=665620 427040 1 0 $X=665430 $Y=424080
X1891 1 2 1784 407 1796 ICV_28 $T=669760 383520 0 0 $X=669570 $Y=383280
X1892 1 2 1786 360 1823 ICV_28 $T=680800 437920 1 0 $X=680610 $Y=434960
X1893 1 2 1862 400 1880 ICV_28 $T=707480 388960 0 0 $X=707290 $Y=388720
X1894 1 2 517 11 537 ICV_29 $T=6900 388960 1 0 $X=6710 $Y=386000
X1895 1 2 38 9 571 ICV_29 $T=27600 443360 1 0 $X=27410 $Y=440400
X1896 1 2 604 10 613 ICV_29 $T=51980 410720 0 0 $X=51790 $Y=410480
X1897 1 2 637 13 688 ICV_29 $T=83720 394400 1 0 $X=83530 $Y=391440
X1898 1 2 664 29 703 ICV_29 $T=92000 388960 1 0 $X=91810 $Y=386000
X1899 1 2 759 29 770 ICV_29 $T=126960 405280 0 0 $X=126770 $Y=405040
X1900 1 2 855 109 896 ICV_29 $T=188600 399840 1 0 $X=188410 $Y=396880
X1901 1 2 926 111 964 ICV_29 $T=224020 399840 1 0 $X=223830 $Y=396880
X1902 1 2 957 127 992 ICV_29 $T=240120 427040 0 0 $X=239930 $Y=426800
X1903 1 2 1014 126 1034 ICV_29 $T=258520 432480 0 0 $X=258330 $Y=432240
X1904 1 2 1023 109 1039 ICV_29 $T=261280 416160 1 0 $X=261090 $Y=413200
X1905 1 2 1076 109 1096 ICV_29 $T=287960 405280 1 0 $X=287770 $Y=402320
X1906 1 2 193 227 1195 ICV_29 $T=345920 443360 1 0 $X=345730 $Y=440400
X1907 1 2 1185 224 1200 ICV_29 $T=346840 432480 1 0 $X=346650 $Y=429520
X1908 1 2 1286 199 1302 ICV_29 $T=399280 427040 1 0 $X=399090 $Y=424080
X1909 1 2 1321 199 1341 ICV_29 $T=420440 421600 1 0 $X=420250 $Y=418640
X1910 1 2 1408 185 313 ICV_29 $T=462300 378080 0 0 $X=462110 $Y=377840
X1911 1 2 1427 189 1439 ICV_29 $T=469200 394400 1 0 $X=469010 $Y=391440
X1912 1 2 319 227 1477 ICV_29 $T=486680 432480 1 0 $X=486490 $Y=429520
X1913 1 2 1540 372 1556 ICV_29 $T=546480 421600 0 0 $X=546290 $Y=421360
X1914 1 2 1540 378 1565 ICV_29 $T=555220 432480 0 0 $X=555030 $Y=432240
X1915 1 2 1540 359 1571 ICV_29 $T=556140 421600 0 0 $X=555950 $Y=421360
X1916 1 2 1641 406 1662 ICV_29 $T=598000 394400 1 0 $X=597810 $Y=391440
X1917 1 2 1730 378 1745 ICV_29 $T=641240 410720 0 0 $X=641050 $Y=410480
X1918 1 2 1747 357 444 ICV_29 $T=658720 437920 0 0 $X=658530 $Y=437680
X1919 1 2 1784 406 1822 ICV_29 $T=679880 383520 1 0 $X=679690 $Y=380560
X1920 1 2 1828 402 1852 ICV_29 $T=693680 394400 1 0 $X=693490 $Y=391440
X1921 1 2 1828 405 1853 ICV_29 $T=693680 399840 1 0 $X=693490 $Y=396880
X1922 1 2 21 18 23 537 543 24 ICV_30 $T=15640 378080 0 0 $X=15450 $Y=377840
X1923 1 2 542 521 31 540 543 16 ICV_30 $T=20240 394400 0 0 $X=20050 $Y=394160
X1924 1 2 545 534 34 556 534 37 ICV_30 $T=23920 416160 0 0 $X=23730 $Y=415920
X1925 1 2 551 533 37 565 554 24 ICV_30 $T=25300 427040 0 0 $X=25110 $Y=426800
X1926 1 2 571 43 25 585 43 23 ICV_30 $T=37260 437920 1 0 $X=37070 $Y=434960
X1927 1 2 621 615 36 622 615 37 ICV_30 $T=62100 421600 0 0 $X=61910 $Y=421360
X1928 1 2 652 51 23 656 51 24 ICV_30 $T=76360 383520 1 0 $X=76170 $Y=380560
X1929 1 2 649 648 23 655 648 36 ICV_30 $T=76360 405280 1 0 $X=76170 $Y=402320
X1930 1 2 677 673 16 681 673 37 ICV_30 $T=85100 432480 1 0 $X=84910 $Y=429520
X1931 1 2 678 634 36 680 634 37 ICV_30 $T=90160 388960 0 0 $X=89970 $Y=388720
X1932 1 2 691 673 36 698 673 24 ICV_30 $T=93380 432480 1 0 $X=93190 $Y=429520
X1933 1 2 705 74 37 706 74 16 ICV_30 $T=103040 378080 0 0 $X=102850 $Y=377840
X1934 1 2 718 720 16 731 732 16 ICV_30 $T=109020 421600 1 0 $X=108830 $Y=418640
X1935 1 2 733 66 36 727 66 24 ICV_30 $T=116380 388960 1 0 $X=116190 $Y=386000
X1936 1 2 745 732 36 750 732 34 ICV_30 $T=120520 427040 1 0 $X=120330 $Y=424080
X1937 1 2 771 773 34 770 773 37 ICV_30 $T=137540 405280 0 0 $X=137350 $Y=405040
X1938 1 2 115 116 118 813 116 119 ICV_30 $T=151800 383520 1 0 $X=151610 $Y=380560
X1939 1 2 797 798 119 818 798 122 ICV_30 $T=152720 405280 0 0 $X=152530 $Y=405040
X1940 1 2 810 809 122 799 809 118 ICV_30 $T=155940 416160 0 0 $X=155750 $Y=415920
X1941 1 2 815 819 122 837 809 129 ICV_30 $T=164220 416160 0 0 $X=164030 $Y=415920
X1942 1 2 847 845 128 852 854 130 ICV_30 $T=174340 410720 0 0 $X=174150 $Y=410480
X1943 1 2 905 888 122 906 888 118 ICV_30 $T=207000 388960 1 0 $X=206810 $Y=386000
X1944 1 2 924 873 123 925 873 122 ICV_30 $T=212060 394400 0 0 $X=211870 $Y=394160
X1945 1 2 935 936 129 938 936 131 ICV_30 $T=221260 394400 0 0 $X=221070 $Y=394160
X1946 1 2 937 147 131 954 147 129 ICV_30 $T=221720 437920 0 0 $X=221530 $Y=437680
X1947 1 2 981 980 118 986 980 130 ICV_30 $T=241960 421600 0 0 $X=241770 $Y=421360
X1948 1 2 983 951 122 987 951 128 ICV_30 $T=244720 388960 1 0 $X=244530 $Y=386000
X1949 1 2 1051 1053 128 1054 1053 130 ICV_30 $T=278300 399840 1 0 $X=278110 $Y=396880
X1950 1 2 1063 1038 128 1078 1079 128 ICV_30 $T=287960 410720 1 0 $X=287770 $Y=407760
X1951 1 2 1084 1067 118 1081 1079 130 ICV_30 $T=293940 421600 0 0 $X=293750 $Y=421360
X1952 1 2 175 176 129 1090 176 131 ICV_30 $T=296700 437920 0 0 $X=296510 $Y=437680
X1953 1 2 1095 176 122 178 176 128 ICV_30 $T=300840 443360 1 0 $X=300650 $Y=440400
X1954 1 2 1126 176 119 186 176 118 ICV_30 $T=312340 443360 1 0 $X=312150 $Y=440400
X1955 1 2 1130 1107 123 1134 1107 118 ICV_30 $T=318780 421600 1 0 $X=318590 $Y=418640
X1956 1 2 1143 1144 206 1149 1144 221 ICV_30 $T=324300 399840 0 0 $X=324110 $Y=399600
X1957 1 2 1150 215 188 1156 215 187 ICV_30 $T=329360 432480 0 0 $X=329170 $Y=432240
X1958 1 2 1153 1152 183 1159 1152 195 ICV_30 $T=330740 421600 1 0 $X=330550 $Y=418640
X1959 1 2 1155 1152 188 1172 1152 192 ICV_30 $T=339020 421600 1 0 $X=338830 $Y=418640
X1960 1 2 1176 1152 220 1182 215 192 ICV_30 $T=342700 427040 0 0 $X=342510 $Y=426800
X1961 1 2 1188 215 239 1194 1199 183 ICV_30 $T=350980 427040 0 0 $X=350790 $Y=426800
X1962 1 2 1204 1168 236 1198 1168 209 ICV_30 $T=356960 394400 1 0 $X=356770 $Y=391440
X1963 1 2 1171 1152 239 1205 1199 195 ICV_30 $T=356960 421600 1 0 $X=356770 $Y=418640
X1964 1 2 1202 1199 188 1216 1199 192 ICV_30 $T=359260 427040 0 0 $X=359070 $Y=426800
X1965 1 2 1218 251 183 1220 1199 239 ICV_30 $T=363860 437920 1 0 $X=363670 $Y=434960
X1966 1 2 1229 1207 206 1238 1207 230 ICV_30 $T=370760 383520 0 0 $X=370570 $Y=383280
X1967 1 2 1230 1225 209 1231 1225 230 ICV_30 $T=371680 388960 0 0 $X=371490 $Y=388720
X1968 1 2 1237 1239 239 1240 1239 187 ICV_30 $T=372140 405280 0 0 $X=371950 $Y=405040
X1969 1 2 1252 251 188 1247 251 220 ICV_30 $T=379500 437920 0 0 $X=379310 $Y=437680
X1970 1 2 1255 259 236 261 259 230 ICV_30 $T=385020 383520 1 0 $X=384830 $Y=380560
X1971 1 2 1288 1290 237 1289 1290 205 ICV_30 $T=402500 399840 1 0 $X=402310 $Y=396880
X1972 1 2 1313 1317 206 1316 1317 236 ICV_30 $T=414920 399840 1 0 $X=414730 $Y=396880
X1973 1 2 1304 1305 188 1327 1305 220 ICV_30 $T=417220 421600 0 0 $X=417030 $Y=421360
X1974 1 2 1319 1323 183 1328 1323 180 ICV_30 $T=417220 432480 0 0 $X=417030 $Y=432240
X1975 1 2 1336 1317 209 1339 1317 205 ICV_30 $T=423200 399840 1 0 $X=423010 $Y=396880
X1976 1 2 1342 1323 220 1344 1323 239 ICV_30 $T=429640 427040 1 0 $X=429450 $Y=424080
X1977 1 2 1349 1350 221 1359 1350 230 ICV_30 $T=432400 399840 1 0 $X=432210 $Y=396880
X1978 1 2 1369 1371 183 1370 1371 195 ICV_30 $T=442980 432480 1 0 $X=442790 $Y=429520
X1979 1 2 1374 1350 237 1376 1380 192 ICV_30 $T=444820 405280 0 0 $X=444630 $Y=405040
X1980 1 2 1368 1371 239 1384 290 180 ICV_30 $T=446200 437920 0 0 $X=446010 $Y=437680
X1981 1 2 1391 1399 230 1405 295 237 ICV_30 $T=455400 388960 0 0 $X=455210 $Y=388720
X1982 1 2 1418 1399 206 1423 312 209 ICV_30 $T=469200 399840 1 0 $X=469010 $Y=396880
X1983 1 2 1421 1403 183 1422 1403 188 ICV_30 $T=469200 421600 0 0 $X=469010 $Y=421360
X1984 1 2 1429 1414 183 317 307 188 ICV_30 $T=471040 427040 0 0 $X=470850 $Y=426800
X1985 1 2 1441 1443 221 1449 312 222 ICV_30 $T=478400 399840 1 0 $X=478210 $Y=396880
X1986 1 2 1451 322 188 1458 322 183 ICV_30 $T=483000 437920 0 0 $X=482810 $Y=437680
X1987 1 2 1450 1447 180 1466 1447 187 ICV_30 $T=488060 416160 1 0 $X=487870 $Y=413200
X1988 1 2 325 307 220 329 322 220 ICV_30 $T=491280 437920 0 0 $X=491090 $Y=437680
X1989 1 2 1490 1487 239 337 336 192 ICV_30 $T=503240 443360 1 0 $X=503050 $Y=440400
X1990 1 2 1495 323 236 1501 326 222 ICV_30 $T=505540 388960 1 0 $X=505350 $Y=386000
X1991 1 2 1521 1516 367 1528 1516 355 ICV_30 $T=528540 421600 0 0 $X=528350 $Y=421360
X1992 1 2 1525 1527 355 1523 1527 367 ICV_30 $T=531760 437920 1 0 $X=531570 $Y=434960
X1993 1 2 1533 1527 363 1542 1527 366 ICV_30 $T=542340 427040 0 0 $X=542150 $Y=426800
X1994 1 2 1541 1516 345 1556 1550 371 ICV_30 $T=550620 427040 0 0 $X=550430 $Y=426800
X1995 1 2 1552 1550 343 1548 1550 345 ICV_30 $T=554300 437920 1 0 $X=554110 $Y=434960
X1996 1 2 1561 1553 386 1560 1553 397 ICV_30 $T=557520 394400 0 0 $X=557330 $Y=394160
X1997 1 2 1563 398 352 1583 398 391 ICV_30 $T=572700 383520 1 0 $X=572510 $Y=380560
X1998 1 2 410 412 387 414 398 387 ICV_30 $T=573620 378080 0 0 $X=573430 $Y=377840
X1999 1 2 1602 1597 345 1617 1586 386 ICV_30 $T=581440 405280 1 0 $X=581250 $Y=402320
X2000 1 2 1605 1597 355 1636 1638 363 ICV_30 $T=591100 421600 1 0 $X=590910 $Y=418640
X2001 1 2 1627 1637 368 1632 1637 343 ICV_30 $T=595240 410720 0 0 $X=595050 $Y=410480
X2002 1 2 1634 1638 366 1628 1637 366 ICV_30 $T=599380 421600 1 0 $X=599190 $Y=418640
X2003 1 2 1654 1655 387 1662 1655 389 ICV_30 $T=603060 388960 0 0 $X=602870 $Y=388720
X2004 1 2 1657 1638 371 1644 1643 355 ICV_30 $T=603980 427040 0 0 $X=603790 $Y=426800
X2005 1 2 1673 1667 371 1677 1667 343 ICV_30 $T=612260 421600 0 0 $X=612070 $Y=421360
X2006 1 2 1683 1690 355 1680 1643 368 ICV_30 $T=619160 432480 1 0 $X=618970 $Y=429520
X2007 1 2 1693 1667 363 1703 1689 366 ICV_30 $T=623300 405280 0 0 $X=623110 $Y=405040
X2008 1 2 1651 1643 363 1660 1643 367 ICV_30 $T=627440 432480 1 0 $X=627250 $Y=429520
X2009 1 2 1694 422 388 1700 1707 391 ICV_30 $T=628360 383520 1 0 $X=628170 $Y=380560
X2010 1 2 1715 1707 392 1708 1707 352 ICV_30 $T=633420 394400 0 0 $X=633230 $Y=394160
X2011 1 2 1719 434 366 1732 434 367 ICV_30 $T=638940 437920 0 0 $X=638750 $Y=437680
X2012 1 2 1727 1728 391 1737 1728 387 ICV_30 $T=641240 394400 1 0 $X=641050 $Y=391440
X2013 1 2 1729 435 388 1725 435 397 ICV_30 $T=642160 378080 0 0 $X=641970 $Y=377840
X2014 1 2 1752 1754 363 1750 1754 345 ICV_30 $T=654580 405280 0 0 $X=654390 $Y=405040
X2015 1 2 1755 1754 368 1749 1754 343 ICV_30 $T=654580 416160 1 0 $X=654390 $Y=413200
X2016 1 2 1756 1728 392 1761 1728 386 ICV_30 $T=655500 394400 1 0 $X=655310 $Y=391440
X2017 1 2 1771 1772 367 1783 1772 366 ICV_30 $T=665620 421600 1 0 $X=665430 $Y=418640
X2018 1 2 1792 1772 371 1793 1772 355 ICV_30 $T=673900 421600 1 0 $X=673710 $Y=418640
X2019 1 2 1791 1799 368 1801 1799 366 ICV_30 $T=674820 405280 1 0 $X=674630 $Y=402320
X2020 1 2 1808 1810 363 1811 1810 367 ICV_30 $T=684020 421600 1 0 $X=683830 $Y=418640
X2021 1 2 1809 1799 367 1780 1770 391 ICV_30 $T=684480 405280 1 0 $X=684290 $Y=402320
X2022 1 2 1812 1810 343 1823 1804 343 ICV_30 $T=684480 432480 0 0 $X=684290 $Y=432240
X2023 1 2 450 451 345 454 455 366 ICV_30 $T=684940 443360 1 0 $X=684750 $Y=440400
X2024 1 2 1868 1869 363 1887 1865 397 ICV_30 $T=713000 405280 1 0 $X=712810 $Y=402320
X2025 1 2 1876 1869 343 1890 1869 355 ICV_30 $T=721740 416160 1 0 $X=721550 $Y=413200
X2026 1 2 6 8 2 516 1 sky130_fd_sc_hd__and2_1 $T=6900 383520 0 0 $X=6710 $Y=383280
X2027 1 2 12 8 2 522 1 sky130_fd_sc_hd__and2_1 $T=8280 394400 0 0 $X=8090 $Y=394160
X2028 1 2 22 8 2 520 1 sky130_fd_sc_hd__and2_1 $T=16100 421600 1 0 $X=15910 $Y=418640
X2029 1 2 32 8 2 548 1 sky130_fd_sc_hd__and2_1 $T=24380 410720 1 0 $X=24190 $Y=407760
X2030 1 2 39 8 2 566 1 sky130_fd_sc_hd__and2_1 $T=31280 383520 0 0 $X=31090 $Y=383280
X2031 1 2 40 8 2 563 1 sky130_fd_sc_hd__and2_1 $T=31740 437920 1 0 $X=31550 $Y=434960
X2032 1 2 42 8 2 570 1 sky130_fd_sc_hd__and2_1 $T=34960 427040 1 0 $X=34770 $Y=424080
X2033 1 2 46 8 2 598 1 sky130_fd_sc_hd__and2_1 $T=48300 432480 1 0 $X=48110 $Y=429520
X2034 1 2 47 8 2 601 1 sky130_fd_sc_hd__and2_1 $T=49680 410720 0 0 $X=49490 $Y=410480
X2035 1 2 50 8 2 602 1 sky130_fd_sc_hd__and2_1 $T=55660 383520 1 0 $X=55470 $Y=380560
X2036 1 2 53 8 2 623 1 sky130_fd_sc_hd__and2_1 $T=58880 378080 0 0 $X=58690 $Y=377840
X2037 1 2 55 8 2 632 1 sky130_fd_sc_hd__and2_1 $T=63020 388960 1 0 $X=62830 $Y=386000
X2038 1 2 57 8 2 638 1 sky130_fd_sc_hd__and2_1 $T=67160 416160 1 0 $X=66970 $Y=413200
X2039 1 2 60 8 2 636 1 sky130_fd_sc_hd__and2_1 $T=75900 394400 0 0 $X=75710 $Y=394160
X2040 1 2 62 8 2 668 1 sky130_fd_sc_hd__and2_1 $T=82340 432480 1 0 $X=82150 $Y=429520
X2041 1 2 65 8 2 667 1 sky130_fd_sc_hd__and2_1 $T=87400 410720 0 0 $X=87210 $Y=410480
X2042 1 2 69 8 2 700 1 sky130_fd_sc_hd__and2_1 $T=96600 394400 0 0 $X=96410 $Y=394160
X2043 1 2 73 8 2 702 1 sky130_fd_sc_hd__and2_1 $T=101660 383520 1 0 $X=101470 $Y=380560
X2044 1 2 72 8 2 701 1 sky130_fd_sc_hd__and2_1 $T=101660 432480 1 0 $X=101470 $Y=429520
X2045 1 2 76 8 2 708 1 sky130_fd_sc_hd__and2_1 $T=104420 416160 1 0 $X=104230 $Y=413200
X2046 1 2 77 8 2 724 1 sky130_fd_sc_hd__and2_1 $T=109940 410720 0 0 $X=109750 $Y=410480
X2047 1 2 80 8 2 734 1 sky130_fd_sc_hd__and2_1 $T=114540 437920 0 0 $X=114350 $Y=437680
X2048 1 2 82 8 2 737 1 sky130_fd_sc_hd__and2_1 $T=115460 388960 0 0 $X=115270 $Y=388720
X2049 1 2 81 8 2 740 1 sky130_fd_sc_hd__and2_1 $T=115460 432480 0 0 $X=115270 $Y=432240
X2050 1 2 86 8 2 736 1 sky130_fd_sc_hd__and2_1 $T=117300 421600 1 0 $X=117110 $Y=418640
X2051 1 2 93 8 2 748 1 sky130_fd_sc_hd__and2_1 $T=123280 399840 0 0 $X=123090 $Y=399600
X2052 1 2 32 107 2 785 1 sky130_fd_sc_hd__and2_1 $T=143520 410720 0 0 $X=143330 $Y=410480
X2053 1 2 7 107 2 789 1 sky130_fd_sc_hd__and2_1 $T=143520 416160 0 0 $X=143330 $Y=415920
X2054 1 2 40 107 2 788 1 sky130_fd_sc_hd__and2_1 $T=143520 432480 0 0 $X=143330 $Y=432240
X2055 1 2 50 107 2 786 1 sky130_fd_sc_hd__and2_1 $T=146280 388960 0 0 $X=146090 $Y=388720
X2056 1 2 60 107 2 787 1 sky130_fd_sc_hd__and2_1 $T=146280 394400 0 0 $X=146090 $Y=394160
X2057 1 2 6 107 2 796 1 sky130_fd_sc_hd__and2_1 $T=157780 378080 0 0 $X=157590 $Y=377840
X2058 1 2 22 107 2 820 1 sky130_fd_sc_hd__and2_1 $T=158700 427040 0 0 $X=158510 $Y=426800
X2059 1 2 57 107 2 841 1 sky130_fd_sc_hd__and2_1 $T=172500 410720 1 0 $X=172310 $Y=407760
X2060 1 2 42 107 2 843 1 sky130_fd_sc_hd__and2_1 $T=174340 416160 0 0 $X=174150 $Y=415920
X2061 1 2 12 107 2 850 1 sky130_fd_sc_hd__and2_1 $T=178480 394400 0 0 $X=178290 $Y=394160
X2062 1 2 39 107 2 868 1 sky130_fd_sc_hd__and2_1 $T=185380 383520 1 0 $X=185190 $Y=380560
X2063 1 2 46 107 2 875 1 sky130_fd_sc_hd__and2_1 $T=185840 427040 1 0 $X=185650 $Y=424080
X2064 1 2 136 107 2 876 1 sky130_fd_sc_hd__and2_1 $T=188600 437920 1 0 $X=188410 $Y=434960
X2065 1 2 47 107 2 904 1 sky130_fd_sc_hd__and2_1 $T=206080 410720 1 0 $X=205890 $Y=407760
X2066 1 2 73 107 2 922 1 sky130_fd_sc_hd__and2_1 $T=210680 378080 0 0 $X=210490 $Y=377840
X2067 1 2 55 107 2 923 1 sky130_fd_sc_hd__and2_1 $T=213900 383520 0 0 $X=213710 $Y=383280
X2068 1 2 77 107 2 929 1 sky130_fd_sc_hd__and2_1 $T=213900 416160 1 0 $X=213710 $Y=413200
X2069 1 2 65 107 2 930 1 sky130_fd_sc_hd__and2_1 $T=213900 432480 1 0 $X=213710 $Y=429520
X2070 1 2 151 107 2 956 1 sky130_fd_sc_hd__and2_1 $T=227700 405280 0 0 $X=227510 $Y=405040
X2071 1 2 150 107 2 958 1 sky130_fd_sc_hd__and2_1 $T=228160 405280 1 0 $X=227970 $Y=402320
X2072 1 2 153 107 2 950 1 sky130_fd_sc_hd__and2_1 $T=230460 432480 0 0 $X=230270 $Y=432240
X2073 1 2 97 107 2 972 1 sky130_fd_sc_hd__and2_1 $T=241040 399840 1 0 $X=240850 $Y=396880
X2074 1 2 156 107 2 979 1 sky130_fd_sc_hd__and2_1 $T=241040 437920 1 0 $X=240850 $Y=434960
X2075 1 2 101 107 2 1000 1 sky130_fd_sc_hd__and2_1 $T=258520 421600 0 0 $X=258330 $Y=421360
X2076 1 2 163 107 2 1016 1 sky130_fd_sc_hd__and2_1 $T=258980 416160 1 0 $X=258790 $Y=413200
X2077 1 2 166 107 2 995 1 sky130_fd_sc_hd__and2_1 $T=265880 383520 0 0 $X=265690 $Y=383280
X2078 1 2 80 107 2 1033 1 sky130_fd_sc_hd__and2_1 $T=268640 394400 1 0 $X=268450 $Y=391440
X2079 1 2 86 107 2 167 1 sky130_fd_sc_hd__and2_1 $T=269560 437920 1 0 $X=269370 $Y=434960
X2080 1 2 93 107 2 168 1 sky130_fd_sc_hd__and2_1 $T=271400 378080 0 0 $X=271210 $Y=377840
X2081 1 2 62 107 2 1055 1 sky130_fd_sc_hd__and2_1 $T=277840 421600 1 0 $X=277650 $Y=418640
X2082 1 2 81 107 2 1060 1 sky130_fd_sc_hd__and2_1 $T=281060 437920 1 0 $X=280870 $Y=434960
X2083 1 2 152 107 2 1061 1 sky130_fd_sc_hd__and2_1 $T=283820 383520 0 0 $X=283630 $Y=383280
X2084 1 2 82 107 2 1082 1 sky130_fd_sc_hd__and2_1 $T=292100 394400 0 0 $X=291910 $Y=394160
X2085 1 2 100 107 2 1101 1 sky130_fd_sc_hd__and2_1 $T=300840 427040 1 0 $X=300650 $Y=424080
X2086 1 2 177 107 2 1098 1 sky130_fd_sc_hd__and2_1 $T=300840 437920 1 0 $X=300650 $Y=434960
X2087 1 2 223 225 2 1154 1 sky130_fd_sc_hd__and2_1 $T=332580 399840 0 0 $X=332390 $Y=399600
X2088 1 2 231 232 2 1165 1 sky130_fd_sc_hd__and2_1 $T=336260 432480 1 0 $X=336070 $Y=429520
X2089 1 2 233 225 2 1161 1 sky130_fd_sc_hd__and2_1 $T=337640 388960 1 0 $X=337450 $Y=386000
X2090 1 2 235 232 2 1158 1 sky130_fd_sc_hd__and2_1 $T=338100 410720 1 0 $X=337910 $Y=407760
X2091 1 2 245 225 2 1192 1 sky130_fd_sc_hd__and2_1 $T=353280 399840 1 0 $X=353090 $Y=396880
X2092 1 2 247 232 2 1196 1 sky130_fd_sc_hd__and2_1 $T=356960 405280 1 0 $X=356770 $Y=402320
X2093 1 2 249 232 2 1213 1 sky130_fd_sc_hd__and2_1 $T=361560 437920 1 0 $X=361370 $Y=434960
X2094 1 2 250 232 2 1214 1 sky130_fd_sc_hd__and2_1 $T=364320 410720 1 0 $X=364130 $Y=407760
X2095 1 2 253 225 2 1236 1 sky130_fd_sc_hd__and2_1 $T=374900 399840 1 0 $X=374710 $Y=396880
X2096 1 2 255 232 2 1254 1 sky130_fd_sc_hd__and2_1 $T=381340 427040 1 0 $X=381150 $Y=424080
X2097 1 2 256 225 2 1257 1 sky130_fd_sc_hd__and2_1 $T=382260 405280 1 0 $X=382070 $Y=402320
X2098 1 2 260 232 2 1260 1 sky130_fd_sc_hd__and2_1 $T=387780 405280 0 0 $X=387590 $Y=405040
X2099 1 2 270 225 2 1294 1 sky130_fd_sc_hd__and2_1 $T=403880 405280 0 0 $X=403690 $Y=405040
X2100 1 2 274 232 2 1301 1 sky130_fd_sc_hd__and2_1 $T=408020 410720 1 0 $X=407830 $Y=407760
X2101 1 2 275 232 2 1318 1 sky130_fd_sc_hd__and2_1 $T=414460 427040 1 0 $X=414270 $Y=424080
X2102 1 2 278 225 2 1322 1 sky130_fd_sc_hd__and2_1 $T=416300 399840 0 0 $X=416110 $Y=399600
X2103 1 2 279 232 2 1325 1 sky130_fd_sc_hd__and2_1 $T=417680 437920 0 0 $X=417490 $Y=437680
X2104 1 2 284 232 2 1330 1 sky130_fd_sc_hd__and2_1 $T=423200 405280 0 0 $X=423010 $Y=405040
X2105 1 2 296 232 2 297 1 sky130_fd_sc_hd__and2_1 $T=450340 443360 1 0 $X=450150 $Y=440400
X2106 1 2 301 232 2 1389 1 sky130_fd_sc_hd__and2_1 $T=457700 410720 1 0 $X=457510 $Y=407760
X2107 1 2 300 225 2 1390 1 sky130_fd_sc_hd__and2_1 $T=458160 388960 1 0 $X=457970 $Y=386000
X2108 1 2 304 232 2 1401 1 sky130_fd_sc_hd__and2_1 $T=461380 405280 0 0 $X=461190 $Y=405040
X2109 1 2 302 225 2 1404 1 sky130_fd_sc_hd__and2_1 $T=468280 399840 0 0 $X=468090 $Y=399600
X2110 1 2 311 232 2 1430 1 sky130_fd_sc_hd__and2_1 $T=470120 427040 1 0 $X=469930 $Y=424080
X2111 1 2 315 232 2 1432 1 sky130_fd_sc_hd__and2_1 $T=473800 405280 0 0 $X=473610 $Y=405040
X2112 1 2 308 232 2 1428 1 sky130_fd_sc_hd__and2_1 $T=475640 437920 1 0 $X=475450 $Y=434960
X2113 1 2 318 232 2 1444 1 sky130_fd_sc_hd__and2_1 $T=477940 432480 1 0 $X=477750 $Y=429520
X2114 1 2 320 225 2 1438 1 sky130_fd_sc_hd__and2_1 $T=478860 399840 0 0 $X=478670 $Y=399600
X2115 1 2 314 225 2 1434 1 sky130_fd_sc_hd__and2_1 $T=483000 383520 0 0 $X=482810 $Y=383280
X2116 1 2 330 225 2 331 1 sky130_fd_sc_hd__and2_1 $T=499100 378080 0 0 $X=498910 $Y=377840
X2117 1 2 333 225 2 1486 1 sky130_fd_sc_hd__and2_1 $T=501400 383520 1 0 $X=501210 $Y=380560
X2118 1 2 334 225 2 1488 1 sky130_fd_sc_hd__and2_1 $T=501400 399840 1 0 $X=501210 $Y=396880
X2119 1 2 335 232 2 1489 1 sky130_fd_sc_hd__and2_1 $T=506920 432480 0 0 $X=506730 $Y=432240
X2120 1 2 338 232 2 1496 1 sky130_fd_sc_hd__and2_1 $T=508760 427040 1 0 $X=508570 $Y=424080
X2121 1 2 235 353 2 1518 1 sky130_fd_sc_hd__and2_1 $T=523940 427040 0 0 $X=523750 $Y=426800
X2122 1 2 240 353 2 1520 1 sky130_fd_sc_hd__and2_1 $T=525780 421600 0 0 $X=525590 $Y=421360
X2123 1 2 384 353 2 1538 1 sky130_fd_sc_hd__and2_1 $T=543260 432480 1 0 $X=543070 $Y=429520
X2124 1 2 233 394 2 1535 1 sky130_fd_sc_hd__and2_1 $T=549240 388960 1 0 $X=549050 $Y=386000
X2125 1 2 231 353 2 1544 1 sky130_fd_sc_hd__and2_1 $T=550160 427040 1 0 $X=549970 $Y=424080
X2126 1 2 247 353 2 1554 1 sky130_fd_sc_hd__and2_1 $T=555220 405280 0 0 $X=555030 $Y=405040
X2127 1 2 255 353 2 1579 1 sky130_fd_sc_hd__and2_1 $T=565340 432480 1 0 $X=565150 $Y=429520
X2128 1 2 260 353 2 1584 1 sky130_fd_sc_hd__and2_1 $T=569940 410720 1 0 $X=569750 $Y=407760
X2129 1 2 285 394 2 1588 1 sky130_fd_sc_hd__and2_1 $T=572240 383520 0 0 $X=572050 $Y=383280
X2130 1 2 253 394 2 1591 1 sky130_fd_sc_hd__and2_1 $T=572700 405280 1 0 $X=572510 $Y=402320
X2131 1 2 250 353 2 1608 1 sky130_fd_sc_hd__and2_1 $T=578680 405280 1 0 $X=578490 $Y=402320
X2132 1 2 249 353 2 1619 1 sky130_fd_sc_hd__and2_1 $T=585120 421600 0 0 $X=584930 $Y=421360
X2133 1 2 284 353 2 1652 1 sky130_fd_sc_hd__and2_1 $T=606280 405280 1 0 $X=606090 $Y=402320
X2134 1 2 270 394 2 1664 1 sky130_fd_sc_hd__and2_1 $T=606740 388960 1 0 $X=606550 $Y=386000
X2135 1 2 275 353 2 1670 1 sky130_fd_sc_hd__and2_1 $T=609960 421600 0 0 $X=609770 $Y=421360
X2136 1 2 263 353 2 1702 1 sky130_fd_sc_hd__and2_1 $T=626520 443360 1 0 $X=626330 $Y=440400
X2137 1 2 304 353 2 1720 1 sky130_fd_sc_hd__and2_1 $T=637100 399840 0 0 $X=636910 $Y=399600
X2138 1 2 292 394 2 1723 1 sky130_fd_sc_hd__and2_1 $T=638480 394400 1 0 $X=638290 $Y=391440
X2139 1 2 318 353 2 1743 1 sky130_fd_sc_hd__and2_1 $T=648140 427040 0 0 $X=647950 $Y=426800
X2140 1 2 320 394 2 1739 1 sky130_fd_sc_hd__and2_1 $T=648600 383520 0 0 $X=648410 $Y=383280
X2141 1 2 291 353 2 1741 1 sky130_fd_sc_hd__and2_1 $T=651360 421600 0 0 $X=651170 $Y=421360
X2142 1 2 328 353 2 1773 1 sky130_fd_sc_hd__and2_1 $T=661940 410720 1 0 $X=661750 $Y=407760
X2143 1 2 302 394 2 1774 1 sky130_fd_sc_hd__and2_1 $T=665620 383520 1 0 $X=665430 $Y=380560
X2144 1 2 308 353 2 1785 1 sky130_fd_sc_hd__and2_1 $T=669760 437920 1 0 $X=669570 $Y=434960
X2145 1 2 335 353 2 1790 1 sky130_fd_sc_hd__and2_1 $T=672980 432480 1 0 $X=672790 $Y=429520
X2146 1 2 300 394 2 1794 1 sky130_fd_sc_hd__and2_1 $T=676660 394400 0 0 $X=676470 $Y=394160
X2147 1 2 315 353 2 1821 1 sky130_fd_sc_hd__and2_1 $T=689540 410720 1 0 $X=689350 $Y=407760
X2148 1 2 333 394 2 1825 1 sky130_fd_sc_hd__and2_1 $T=690920 399840 0 0 $X=690730 $Y=399600
X2149 1 2 338 353 2 1843 1 sky130_fd_sc_hd__and2_1 $T=704720 432480 0 0 $X=704530 $Y=432240
X2150 1 2 311 353 2 1837 1 sky130_fd_sc_hd__and2_1 $T=705640 427040 1 0 $X=705450 $Y=424080
X2151 1 2 330 394 2 1856 1 sky130_fd_sc_hd__and2_1 $T=707480 378080 0 0 $X=707290 $Y=377840
X2152 1 2 334 394 2 1861 1 sky130_fd_sc_hd__and2_1 $T=707480 394400 0 0 $X=707290 $Y=394160
X2153 1 2 301 353 2 1858 1 sky130_fd_sc_hd__and2_1 $T=707480 405280 0 0 $X=707290 $Y=405040
X2154 1 2 466 516 2 517 1 sky130_fd_sc_hd__dlclkp_1 $T=6900 383520 1 0 $X=6710 $Y=380560
X2155 1 2 466 520 2 514 1 sky130_fd_sc_hd__dlclkp_1 $T=7360 427040 0 0 $X=7170 $Y=426800
X2156 1 2 466 519 2 515 1 sky130_fd_sc_hd__dlclkp_1 $T=9660 416160 0 0 $X=9470 $Y=415920
X2157 1 2 466 15 2 5 1 sky130_fd_sc_hd__dlclkp_1 $T=10120 437920 0 0 $X=9930 $Y=437680
X2158 1 2 466 522 2 513 1 sky130_fd_sc_hd__dlclkp_1 $T=10580 394400 0 0 $X=10390 $Y=394160
X2159 1 2 466 548 2 564 1 sky130_fd_sc_hd__dlclkp_1 $T=23460 405280 0 0 $X=23270 $Y=405040
X2160 1 2 466 563 2 38 1 sky130_fd_sc_hd__dlclkp_1 $T=27140 437920 0 0 $X=26950 $Y=437680
X2161 1 2 466 566 2 567 1 sky130_fd_sc_hd__dlclkp_1 $T=30360 383520 1 0 $X=30170 $Y=380560
X2162 1 2 466 570 2 555 1 sky130_fd_sc_hd__dlclkp_1 $T=35880 421600 1 0 $X=35690 $Y=418640
X2163 1 2 466 598 2 48 1 sky130_fd_sc_hd__dlclkp_1 $T=45540 427040 0 0 $X=45350 $Y=426800
X2164 1 2 466 601 2 604 1 sky130_fd_sc_hd__dlclkp_1 $T=48760 405280 0 0 $X=48570 $Y=405040
X2165 1 2 466 602 2 594 1 sky130_fd_sc_hd__dlclkp_1 $T=49220 388960 1 0 $X=49030 $Y=386000
X2166 1 2 466 623 2 597 1 sky130_fd_sc_hd__dlclkp_1 $T=57960 383520 1 0 $X=57770 $Y=380560
X2167 1 2 466 632 2 637 1 sky130_fd_sc_hd__dlclkp_1 $T=62100 388960 0 0 $X=61910 $Y=388720
X2168 1 2 466 636 2 635 1 sky130_fd_sc_hd__dlclkp_1 $T=64860 399840 1 0 $X=64670 $Y=396880
X2169 1 2 466 638 2 631 1 sky130_fd_sc_hd__dlclkp_1 $T=69460 416160 1 0 $X=69270 $Y=413200
X2170 1 2 466 667 2 676 1 sky130_fd_sc_hd__dlclkp_1 $T=80960 410720 0 0 $X=80770 $Y=410480
X2171 1 2 466 668 2 56 1 sky130_fd_sc_hd__dlclkp_1 $T=80960 437920 1 0 $X=80770 $Y=434960
X2172 1 2 466 700 2 695 1 sky130_fd_sc_hd__dlclkp_1 $T=95680 394400 1 0 $X=95490 $Y=391440
X2173 1 2 466 701 2 64 1 sky130_fd_sc_hd__dlclkp_1 $T=95680 437920 1 0 $X=95490 $Y=434960
X2174 1 2 466 702 2 664 1 sky130_fd_sc_hd__dlclkp_1 $T=97520 383520 0 0 $X=97330 $Y=383280
X2175 1 2 466 708 2 665 1 sky130_fd_sc_hd__dlclkp_1 $T=100740 416160 0 0 $X=100550 $Y=415920
X2176 1 2 466 734 2 75 1 sky130_fd_sc_hd__dlclkp_1 $T=112240 443360 1 0 $X=112050 $Y=440400
X2177 1 2 466 736 2 711 1 sky130_fd_sc_hd__dlclkp_1 $T=114080 427040 1 0 $X=113890 $Y=424080
X2178 1 2 466 724 2 712 1 sky130_fd_sc_hd__dlclkp_1 $T=118220 416160 0 0 $X=118030 $Y=415920
X2179 1 2 466 740 2 749 1 sky130_fd_sc_hd__dlclkp_1 $T=119140 432480 0 0 $X=118950 $Y=432240
X2180 1 2 466 737 2 746 1 sky130_fd_sc_hd__dlclkp_1 $T=119600 388960 0 0 $X=119410 $Y=388720
X2181 1 2 466 748 2 759 1 sky130_fd_sc_hd__dlclkp_1 $T=122820 405280 1 0 $X=122630 $Y=402320
X2182 1 2 466 763 2 89 1 sky130_fd_sc_hd__dlclkp_1 $T=135240 443360 1 0 $X=135050 $Y=440400
X2183 1 2 466 785 2 792 1 sky130_fd_sc_hd__dlclkp_1 $T=141220 410720 1 0 $X=141030 $Y=407760
X2184 1 2 466 786 2 793 1 sky130_fd_sc_hd__dlclkp_1 $T=141680 388960 1 0 $X=141490 $Y=386000
X2185 1 2 466 787 2 794 1 sky130_fd_sc_hd__dlclkp_1 $T=142600 399840 1 0 $X=142410 $Y=396880
X2186 1 2 466 788 2 108 1 sky130_fd_sc_hd__dlclkp_1 $T=142600 437920 1 0 $X=142410 $Y=434960
X2187 1 2 466 789 2 795 1 sky130_fd_sc_hd__dlclkp_1 $T=143520 421600 1 0 $X=143330 $Y=418640
X2188 1 2 466 110 2 117 1 sky130_fd_sc_hd__dlclkp_1 $T=147200 437920 0 0 $X=147010 $Y=437680
X2189 1 2 466 796 2 121 1 sky130_fd_sc_hd__dlclkp_1 $T=151340 378080 0 0 $X=151150 $Y=377840
X2190 1 2 466 820 2 132 1 sky130_fd_sc_hd__dlclkp_1 $T=166520 432480 1 0 $X=166330 $Y=429520
X2191 1 2 466 841 2 846 1 sky130_fd_sc_hd__dlclkp_1 $T=167440 399840 0 0 $X=167250 $Y=399600
X2192 1 2 466 843 2 848 1 sky130_fd_sc_hd__dlclkp_1 $T=171120 416160 1 0 $X=170930 $Y=413200
X2193 1 2 466 850 2 855 1 sky130_fd_sc_hd__dlclkp_1 $T=176640 399840 1 0 $X=176450 $Y=396880
X2194 1 2 466 868 2 874 1 sky130_fd_sc_hd__dlclkp_1 $T=181700 388960 1 0 $X=181510 $Y=386000
X2195 1 2 466 876 2 137 1 sky130_fd_sc_hd__dlclkp_1 $T=187220 432480 0 0 $X=187030 $Y=432240
X2196 1 2 466 875 2 879 1 sky130_fd_sc_hd__dlclkp_1 $T=188600 427040 1 0 $X=188410 $Y=424080
X2197 1 2 466 904 2 901 1 sky130_fd_sc_hd__dlclkp_1 $T=204700 405280 1 0 $X=204510 $Y=402320
X2198 1 2 466 922 2 927 1 sky130_fd_sc_hd__dlclkp_1 $T=209760 383520 1 0 $X=209570 $Y=380560
X2199 1 2 466 923 2 926 1 sky130_fd_sc_hd__dlclkp_1 $T=209760 394400 1 0 $X=209570 $Y=391440
X2200 1 2 466 145 2 146 1 sky130_fd_sc_hd__dlclkp_1 $T=212980 378080 0 0 $X=212790 $Y=377840
X2201 1 2 466 930 2 931 1 sky130_fd_sc_hd__dlclkp_1 $T=214360 427040 0 0 $X=214170 $Y=426800
X2202 1 2 466 929 2 932 1 sky130_fd_sc_hd__dlclkp_1 $T=218040 410720 0 0 $X=217850 $Y=410480
X2203 1 2 466 950 2 957 1 sky130_fd_sc_hd__dlclkp_1 $T=223560 432480 0 0 $X=223370 $Y=432240
X2204 1 2 466 958 2 969 1 sky130_fd_sc_hd__dlclkp_1 $T=230460 405280 1 0 $X=230270 $Y=402320
X2205 1 2 466 956 2 965 1 sky130_fd_sc_hd__dlclkp_1 $T=230460 405280 0 0 $X=230270 $Y=405040
X2206 1 2 466 972 2 984 1 sky130_fd_sc_hd__dlclkp_1 $T=237820 394400 0 0 $X=237630 $Y=394160
X2207 1 2 466 979 2 157 1 sky130_fd_sc_hd__dlclkp_1 $T=238740 437920 0 0 $X=238550 $Y=437680
X2208 1 2 466 995 2 160 1 sky130_fd_sc_hd__dlclkp_1 $T=250240 383520 0 0 $X=250050 $Y=383280
X2209 1 2 466 1000 2 1014 1 sky130_fd_sc_hd__dlclkp_1 $T=250700 421600 0 0 $X=250510 $Y=421360
X2210 1 2 466 1016 2 1023 1 sky130_fd_sc_hd__dlclkp_1 $T=258520 416160 0 0 $X=258330 $Y=415920
X2211 1 2 466 1033 2 1041 1 sky130_fd_sc_hd__dlclkp_1 $T=265880 405280 1 0 $X=265690 $Y=402320
X2212 1 2 466 1055 2 1050 1 sky130_fd_sc_hd__dlclkp_1 $T=277840 427040 1 0 $X=277650 $Y=424080
X2213 1 2 466 1058 2 1066 1 sky130_fd_sc_hd__dlclkp_1 $T=279680 416160 0 0 $X=279490 $Y=415920
X2214 1 2 466 1061 2 1072 1 sky130_fd_sc_hd__dlclkp_1 $T=281520 388960 1 0 $X=281330 $Y=386000
X2215 1 2 466 1060 2 172 1 sky130_fd_sc_hd__dlclkp_1 $T=281520 443360 1 0 $X=281330 $Y=440400
X2216 1 2 466 1082 2 1076 1 sky130_fd_sc_hd__dlclkp_1 $T=294400 394400 0 0 $X=294210 $Y=394160
X2217 1 2 466 1098 2 1103 1 sky130_fd_sc_hd__dlclkp_1 $T=295780 432480 0 0 $X=295590 $Y=432240
X2218 1 2 466 1101 2 1104 1 sky130_fd_sc_hd__dlclkp_1 $T=297160 427040 0 0 $X=296970 $Y=426800
X2219 1 2 472 1154 2 1128 1 sky130_fd_sc_hd__dlclkp_1 $T=329820 399840 1 0 $X=329630 $Y=396880
X2220 1 2 472 1158 2 1141 1 sky130_fd_sc_hd__dlclkp_1 $T=332580 416160 0 0 $X=332390 $Y=415920
X2221 1 2 472 1161 2 1129 1 sky130_fd_sc_hd__dlclkp_1 $T=333960 383520 0 0 $X=333770 $Y=383280
X2222 1 2 472 1165 2 1146 1 sky130_fd_sc_hd__dlclkp_1 $T=335340 427040 0 0 $X=335150 $Y=426800
X2223 1 2 472 1180 2 1185 1 sky130_fd_sc_hd__dlclkp_1 $T=344080 421600 0 0 $X=343890 $Y=421360
X2224 1 2 472 1192 2 1167 1 sky130_fd_sc_hd__dlclkp_1 $T=350060 405280 1 0 $X=349870 $Y=402320
X2225 1 2 472 244 2 193 1 sky130_fd_sc_hd__dlclkp_1 $T=350060 437920 0 0 $X=349870 $Y=437680
X2226 1 2 472 1196 2 1173 1 sky130_fd_sc_hd__dlclkp_1 $T=353740 405280 0 0 $X=353550 $Y=405040
X2227 1 2 472 1214 2 1211 1 sky130_fd_sc_hd__dlclkp_1 $T=362020 405280 0 0 $X=361830 $Y=405040
X2228 1 2 472 1213 2 248 1 sky130_fd_sc_hd__dlclkp_1 $T=367080 443360 1 0 $X=366890 $Y=440400
X2229 1 2 472 1236 2 1210 1 sky130_fd_sc_hd__dlclkp_1 $T=370760 405280 1 0 $X=370570 $Y=402320
X2230 1 2 472 1254 2 1233 1 sky130_fd_sc_hd__dlclkp_1 $T=379960 421600 0 0 $X=379770 $Y=421360
X2231 1 2 472 1257 2 1256 1 sky130_fd_sc_hd__dlclkp_1 $T=381340 405280 0 0 $X=381150 $Y=405040
X2232 1 2 472 1260 2 1259 1 sky130_fd_sc_hd__dlclkp_1 $T=385480 410720 0 0 $X=385290 $Y=410480
X2233 1 2 472 1281 2 258 1 sky130_fd_sc_hd__dlclkp_1 $T=395140 432480 1 0 $X=394950 $Y=429520
X2234 1 2 472 1294 2 1282 1 sky130_fd_sc_hd__dlclkp_1 $T=403420 405280 1 0 $X=403230 $Y=402320
X2235 1 2 472 1301 2 1286 1 sky130_fd_sc_hd__dlclkp_1 $T=406180 416160 1 0 $X=405990 $Y=413200
X2236 1 2 472 1318 2 1306 1 sky130_fd_sc_hd__dlclkp_1 $T=416760 427040 1 0 $X=416570 $Y=424080
X2237 1 2 472 1330 2 1321 1 sky130_fd_sc_hd__dlclkp_1 $T=419520 410720 0 0 $X=419330 $Y=410480
X2238 1 2 472 1325 2 272 1 sky130_fd_sc_hd__dlclkp_1 $T=419980 437920 0 0 $X=419790 $Y=437680
X2239 1 2 472 1322 2 1300 1 sky130_fd_sc_hd__dlclkp_1 $T=420440 405280 1 0 $X=420250 $Y=402320
X2240 1 2 472 1338 2 277 1 sky130_fd_sc_hd__dlclkp_1 $T=423200 383520 1 0 $X=423010 $Y=380560
X2241 1 2 472 287 2 288 1 sky130_fd_sc_hd__dlclkp_1 $T=428720 378080 0 0 $X=428530 $Y=377840
X2242 1 2 472 1365 2 1353 1 sky130_fd_sc_hd__dlclkp_1 $T=437920 421600 0 0 $X=437730 $Y=421360
X2243 1 2 472 1366 2 1340 1 sky130_fd_sc_hd__dlclkp_1 $T=438380 405280 0 0 $X=438190 $Y=405040
X2244 1 2 472 1389 2 1364 1 sky130_fd_sc_hd__dlclkp_1 $T=451260 410720 1 0 $X=451070 $Y=407760
X2245 1 2 472 1390 2 293 1 sky130_fd_sc_hd__dlclkp_1 $T=451720 388960 1 0 $X=451530 $Y=386000
X2246 1 2 472 1401 2 1407 1 sky130_fd_sc_hd__dlclkp_1 $T=454940 405280 0 0 $X=454750 $Y=405040
X2247 1 2 472 1404 2 1377 1 sky130_fd_sc_hd__dlclkp_1 $T=457240 405280 1 0 $X=457050 $Y=402320
X2248 1 2 472 1428 2 298 1 sky130_fd_sc_hd__dlclkp_1 $T=469200 437920 1 0 $X=469010 $Y=434960
X2249 1 2 472 1430 2 1400 1 sky130_fd_sc_hd__dlclkp_1 $T=472420 427040 1 0 $X=472230 $Y=424080
X2250 1 2 472 1434 2 1408 1 sky130_fd_sc_hd__dlclkp_1 $T=474260 383520 0 0 $X=474070 $Y=383280
X2251 1 2 472 1432 2 1431 1 sky130_fd_sc_hd__dlclkp_1 $T=474720 410720 1 0 $X=474530 $Y=407760
X2252 1 2 472 1438 2 1427 1 sky130_fd_sc_hd__dlclkp_1 $T=476100 405280 0 0 $X=475910 $Y=405040
X2253 1 2 472 1444 2 319 1 sky130_fd_sc_hd__dlclkp_1 $T=480240 432480 1 0 $X=480050 $Y=429520
X2254 1 2 472 1486 2 324 1 sky130_fd_sc_hd__dlclkp_1 $T=498640 388960 1 0 $X=498450 $Y=386000
X2255 1 2 472 1482 2 1483 1 sky130_fd_sc_hd__dlclkp_1 $T=498640 410720 1 0 $X=498450 $Y=407760
X2256 1 2 472 1488 2 1456 1 sky130_fd_sc_hd__dlclkp_1 $T=500480 399840 0 0 $X=500290 $Y=399600
X2257 1 2 472 1489 2 332 1 sky130_fd_sc_hd__dlclkp_1 $T=500480 432480 0 0 $X=500290 $Y=432240
X2258 1 2 472 1496 2 1470 1 sky130_fd_sc_hd__dlclkp_1 $T=504160 421600 0 0 $X=503970 $Y=421360
X2259 1 2 472 1520 2 1519 1 sky130_fd_sc_hd__dlclkp_1 $T=525320 416160 1 0 $X=525130 $Y=413200
X2260 1 2 472 1518 2 1517 1 sky130_fd_sc_hd__dlclkp_1 $T=525320 437920 1 0 $X=525130 $Y=434960
X2261 1 2 472 1535 2 390 1 sky130_fd_sc_hd__dlclkp_1 $T=542800 383520 0 0 $X=542610 $Y=383280
X2262 1 2 472 1538 2 385 1 sky130_fd_sc_hd__dlclkp_1 $T=545100 437920 1 0 $X=544910 $Y=434960
X2263 1 2 472 1546 2 1543 1 sky130_fd_sc_hd__dlclkp_1 $T=551080 394400 0 0 $X=550890 $Y=394160
X2264 1 2 472 1554 2 1539 1 sky130_fd_sc_hd__dlclkp_1 $T=553380 405280 1 0 $X=553190 $Y=402320
X2265 1 2 472 1544 2 1540 1 sky130_fd_sc_hd__dlclkp_1 $T=553380 427040 1 0 $X=553190 $Y=424080
X2266 1 2 472 1584 2 1585 1 sky130_fd_sc_hd__dlclkp_1 $T=566260 405280 1 0 $X=566070 $Y=402320
X2267 1 2 472 1572 2 409 1 sky130_fd_sc_hd__dlclkp_1 $T=566260 443360 1 0 $X=566070 $Y=440400
X2268 1 2 472 1579 2 1580 1 sky130_fd_sc_hd__dlclkp_1 $T=567640 432480 0 0 $X=567450 $Y=432240
X2269 1 2 472 1588 2 1592 1 sky130_fd_sc_hd__dlclkp_1 $T=570400 388960 0 0 $X=570210 $Y=388720
X2270 1 2 472 1591 2 1587 1 sky130_fd_sc_hd__dlclkp_1 $T=571320 399840 0 0 $X=571130 $Y=399600
X2271 1 2 472 1608 2 1618 1 sky130_fd_sc_hd__dlclkp_1 $T=580980 405280 0 0 $X=580790 $Y=405040
X2272 1 2 472 1619 2 1621 1 sky130_fd_sc_hd__dlclkp_1 $T=584660 421600 1 0 $X=584470 $Y=418640
X2273 1 2 472 1620 2 418 1 sky130_fd_sc_hd__dlclkp_1 $T=587420 437920 0 0 $X=587230 $Y=437680
X2274 1 2 472 1648 2 1641 1 sky130_fd_sc_hd__dlclkp_1 $T=599840 405280 1 0 $X=599650 $Y=402320
X2275 1 2 472 1652 2 1658 1 sky130_fd_sc_hd__dlclkp_1 $T=600760 405280 0 0 $X=600570 $Y=405040
X2276 1 2 472 1664 2 421 1 sky130_fd_sc_hd__dlclkp_1 $T=609500 388960 1 0 $X=609310 $Y=386000
X2277 1 2 472 1670 2 1671 1 sky130_fd_sc_hd__dlclkp_1 $T=611800 432480 1 0 $X=611610 $Y=429520
X2278 1 2 472 1686 2 1685 1 sky130_fd_sc_hd__dlclkp_1 $T=617320 399840 1 0 $X=617130 $Y=396880
X2279 1 2 472 1699 2 1698 1 sky130_fd_sc_hd__dlclkp_1 $T=623300 410720 0 0 $X=623110 $Y=410480
X2280 1 2 472 1702 2 429 1 sky130_fd_sc_hd__dlclkp_1 $T=625140 437920 0 0 $X=624950 $Y=437680
X2281 1 2 472 428 2 430 1 sky130_fd_sc_hd__dlclkp_1 $T=625600 378080 0 0 $X=625410 $Y=377840
X2282 1 2 472 1720 2 1730 1 sky130_fd_sc_hd__dlclkp_1 $T=637100 405280 0 0 $X=636910 $Y=405040
X2283 1 2 472 1723 2 1721 1 sky130_fd_sc_hd__dlclkp_1 $T=638480 405280 1 0 $X=638290 $Y=402320
X2284 1 2 472 1739 2 437 1 sky130_fd_sc_hd__dlclkp_1 $T=644920 383520 1 0 $X=644730 $Y=380560
X2285 1 2 472 1741 2 1751 1 sky130_fd_sc_hd__dlclkp_1 $T=646300 427040 1 0 $X=646110 $Y=424080
X2286 1 2 472 1743 2 1747 1 sky130_fd_sc_hd__dlclkp_1 $T=651360 427040 0 0 $X=651170 $Y=426800
X2287 1 2 472 1753 2 1765 1 sky130_fd_sc_hd__dlclkp_1 $T=654120 399840 0 0 $X=653930 $Y=399600
X2288 1 2 472 1773 2 1777 1 sky130_fd_sc_hd__dlclkp_1 $T=661480 410720 0 0 $X=661290 $Y=410480
X2289 1 2 472 1774 2 445 1 sky130_fd_sc_hd__dlclkp_1 $T=662400 378080 0 0 $X=662210 $Y=377840
X2290 1 2 472 1785 2 1786 1 sky130_fd_sc_hd__dlclkp_1 $T=670220 437920 0 0 $X=670030 $Y=437680
X2291 1 2 472 1790 2 1802 1 sky130_fd_sc_hd__dlclkp_1 $T=671140 427040 0 0 $X=670950 $Y=426800
X2292 1 2 472 1794 2 1784 1 sky130_fd_sc_hd__dlclkp_1 $T=672980 399840 1 0 $X=672790 $Y=396880
X2293 1 2 472 452 2 456 1 sky130_fd_sc_hd__dlclkp_1 $T=685860 378080 0 0 $X=685670 $Y=377840
X2294 1 2 472 1821 2 1826 1 sky130_fd_sc_hd__dlclkp_1 $T=686780 405280 0 0 $X=686590 $Y=405040
X2295 1 2 472 1825 2 1828 1 sky130_fd_sc_hd__dlclkp_1 $T=688160 394400 0 0 $X=687970 $Y=394160
X2296 1 2 472 1837 2 1857 1 sky130_fd_sc_hd__dlclkp_1 $T=698740 421600 0 0 $X=698550 $Y=421360
X2297 1 2 472 1843 2 1859 1 sky130_fd_sc_hd__dlclkp_1 $T=699200 427040 1 0 $X=699010 $Y=424080
X2298 1 2 472 1856 2 1862 1 sky130_fd_sc_hd__dlclkp_1 $T=702880 383520 1 0 $X=702690 $Y=380560
X2299 1 2 472 1858 2 1864 1 sky130_fd_sc_hd__dlclkp_1 $T=703340 410720 1 0 $X=703150 $Y=407760
X2300 1 2 472 1861 2 1866 1 sky130_fd_sc_hd__dlclkp_1 $T=705640 405280 1 0 $X=705450 $Y=402320
X2301 1 2 ICV_32 $T=29900 394400 0 0 $X=29710 $Y=394160
X2302 1 2 ICV_32 $T=156400 399840 1 0 $X=156210 $Y=396880
X2303 1 2 ICV_32 $T=156400 416160 1 0 $X=156210 $Y=413200
X2304 1 2 ICV_32 $T=170200 383520 0 0 $X=170010 $Y=383280
X2305 1 2 ICV_32 $T=184460 437920 1 0 $X=184270 $Y=434960
X2306 1 2 ICV_32 $T=198260 394400 0 0 $X=198070 $Y=394160
X2307 1 2 ICV_32 $T=198260 427040 0 0 $X=198070 $Y=426800
X2308 1 2 ICV_32 $T=310500 388960 0 0 $X=310310 $Y=388720
X2309 1 2 ICV_32 $T=310500 394400 0 0 $X=310310 $Y=394160
X2310 1 2 ICV_32 $T=380880 388960 1 0 $X=380690 $Y=386000
X2311 1 2 ICV_32 $T=380880 394400 1 0 $X=380690 $Y=391440
X2312 1 2 ICV_32 $T=380880 437920 1 0 $X=380690 $Y=434960
X2313 1 2 ICV_32 $T=380880 443360 1 0 $X=380690 $Y=440400
X2314 1 2 ICV_32 $T=394680 383520 0 0 $X=394490 $Y=383280
X2315 1 2 ICV_32 $T=408940 427040 1 0 $X=408750 $Y=424080
X2316 1 2 ICV_32 $T=422740 388960 0 0 $X=422550 $Y=388720
X2317 1 2 ICV_32 $T=493120 421600 1 0 $X=492930 $Y=418640
X2318 1 2 ICV_32 $T=647220 388960 0 0 $X=647030 $Y=388720
X2319 1 2 ICV_32 $T=689540 383520 1 0 $X=689350 $Y=380560
X2320 1 2 ICV_32 $T=689540 432480 1 0 $X=689350 $Y=429520
X2321 1 2 ICV_32 $T=717600 383520 1 0 $X=717410 $Y=380560
X2322 1 2 515 9 532 ICV_35 $T=6900 410720 0 0 $X=6710 $Y=410480
X2323 1 2 514 17 541 ICV_35 $T=10580 432480 0 0 $X=10390 $Y=432240
X2324 1 2 555 11 565 ICV_35 $T=27600 421600 1 0 $X=27410 $Y=418640
X2325 1 2 567 30 573 ICV_35 $T=31740 388960 1 0 $X=31550 $Y=386000
X2326 1 2 564 30 575 ICV_35 $T=31740 416160 1 0 $X=31550 $Y=413200
X2327 1 2 555 28 586 ICV_35 $T=36800 432480 1 0 $X=36610 $Y=429520
X2328 1 2 594 17 603 ICV_35 $T=45540 399840 0 0 $X=45350 $Y=399600
X2329 1 2 48 30 612 ICV_35 $T=49680 432480 0 0 $X=49490 $Y=432240
X2330 1 2 604 30 621 ICV_35 $T=51060 421600 0 0 $X=50870 $Y=421360
X2331 1 2 594 9 624 ICV_35 $T=52900 388960 0 0 $X=52710 $Y=388720
X2332 1 2 631 17 639 ICV_35 $T=62100 432480 1 0 $X=61910 $Y=429520
X2333 1 2 597 10 59 ICV_35 $T=65780 383520 1 0 $X=65590 $Y=380560
X2334 1 2 676 17 704 ICV_35 $T=92920 410720 1 0 $X=92730 $Y=407760
X2335 1 2 695 11 714 ICV_35 $T=98900 394400 0 0 $X=98710 $Y=394160
X2336 1 2 64 11 719 ICV_35 $T=101660 432480 0 0 $X=101470 $Y=432240
X2337 1 2 792 109 799 ICV_35 $T=146280 416160 0 0 $X=146090 $Y=415920
X2338 1 2 792 113 810 ICV_35 $T=148120 416160 1 0 $X=147930 $Y=413200
X2339 1 2 794 124 823 ICV_35 $T=157780 399840 0 0 $X=157590 $Y=399600
X2340 1 2 792 126 829 ICV_35 $T=159620 410720 0 0 $X=159430 $Y=410480
X2341 1 2 792 125 837 ICV_35 $T=160540 416160 1 0 $X=160350 $Y=413200
X2342 1 2 846 113 865 ICV_35 $T=174340 405280 0 0 $X=174150 $Y=405040
X2343 1 2 848 125 878 ICV_35 $T=183080 421600 0 0 $X=182890 $Y=421360
X2344 1 2 874 125 884 ICV_35 $T=188600 394400 1 0 $X=188410 $Y=391440
X2345 1 2 879 111 897 ICV_35 $T=189980 427040 0 0 $X=189790 $Y=426800
X2346 1 2 901 126 907 ICV_35 $T=201020 416160 1 0 $X=200830 $Y=413200
X2347 1 2 927 125 944 ICV_35 $T=216200 383520 0 0 $X=216010 $Y=383280
X2348 1 2 927 126 946 ICV_35 $T=216660 383520 1 0 $X=216470 $Y=380560
X2349 1 2 901 113 947 ICV_35 $T=216660 410720 1 0 $X=216470 $Y=407760
X2350 1 2 932 126 948 ICV_35 $T=216660 427040 1 0 $X=216470 $Y=424080
X2351 1 2 927 127 963 ICV_35 $T=224940 383520 1 0 $X=224750 $Y=380560
X2352 1 2 932 109 953 ICV_35 $T=224940 410720 1 0 $X=224750 $Y=407760
X2353 1 2 957 111 974 ICV_35 $T=231840 427040 0 0 $X=231650 $Y=426800
X2354 1 2 984 125 1002 ICV_35 $T=258520 388960 0 0 $X=258330 $Y=388720
X2355 1 2 984 126 1031 ICV_35 $T=258520 394400 0 0 $X=258330 $Y=394160
X2356 1 2 160 126 1036 ICV_35 $T=266800 388960 0 0 $X=266610 $Y=388720
X2357 1 2 160 113 1049 ICV_35 $T=268180 383520 0 0 $X=267990 $Y=383280
X2358 1 2 1041 111 1057 ICV_35 $T=272780 394400 1 0 $X=272590 $Y=391440
X2359 1 2 1023 124 1063 ICV_35 $T=275540 410720 0 0 $X=275350 $Y=410480
X2360 1 2 1066 111 1083 ICV_35 $T=286580 410720 0 0 $X=286390 $Y=410480
X2361 1 2 1050 109 1084 ICV_35 $T=286580 427040 0 0 $X=286390 $Y=426800
X2362 1 2 1050 111 1086 ICV_35 $T=286580 432480 0 0 $X=286390 $Y=432240
X2363 1 2 1076 112 1117 ICV_35 $T=302220 394400 0 0 $X=302030 $Y=394160
X2364 1 2 172 112 1126 ICV_35 $T=304980 437920 0 0 $X=304790 $Y=437680
X2365 1 2 1146 202 1156 ICV_35 $T=325680 427040 0 0 $X=325490 $Y=426800
X2366 1 2 1167 212 1179 ICV_35 $T=337640 394400 1 0 $X=337450 $Y=391440
X2367 1 2 1146 228 1182 ICV_35 $T=338560 432480 1 0 $X=338370 $Y=429520
X2368 1 2 241 190 1229 ICV_35 $T=362020 383520 0 0 $X=361830 $Y=383280
X2369 1 2 1210 212 1231 ICV_35 $T=362020 394400 0 0 $X=361830 $Y=394160
X2370 1 2 1211 202 1240 ICV_35 $T=366620 410720 1 0 $X=366430 $Y=407760
X2371 1 2 254 211 1255 ICV_35 $T=374900 378080 0 0 $X=374710 $Y=377840
X2372 1 2 258 196 265 ICV_35 $T=385020 443360 1 0 $X=384830 $Y=440400
X2373 1 2 1259 202 1283 ICV_35 $T=392380 410720 1 0 $X=392190 $Y=407760
X2374 1 2 1282 211 1292 ICV_35 $T=396520 388960 1 0 $X=396330 $Y=386000
X2375 1 2 272 228 1309 ICV_35 $T=404340 443360 1 0 $X=404150 $Y=440400
X2376 1 2 293 184 1382 ICV_35 $T=441140 388960 1 0 $X=440950 $Y=386000
X2377 1 2 1353 224 1387 ICV_35 $T=443440 427040 0 0 $X=443250 $Y=426800
X2378 1 2 298 202 1406 ICV_35 $T=452640 443360 1 0 $X=452450 $Y=440400
X2379 1 2 1407 202 1419 ICV_35 $T=460000 410720 1 0 $X=459810 $Y=407760
X2380 1 2 1408 189 1423 ICV_35 $T=460460 388960 1 0 $X=460270 $Y=386000
X2381 1 2 1427 185 1440 ICV_35 $T=470580 399840 0 0 $X=470390 $Y=399600
X2382 1 2 1431 213 1446 ICV_35 $T=474260 416160 0 0 $X=474070 $Y=415920
X2383 1 2 332 227 1497 ICV_35 $T=501400 437920 1 0 $X=501210 $Y=434960
X2384 1 2 179 343 356 ICV_35 $T=517040 399840 0 0 $X=516850 $Y=399600
X2385 1 2 1517 357 1523 ICV_35 $T=523940 432480 0 0 $X=523750 $Y=432240
X2386 1 2 1519 357 1521 ICV_35 $T=525320 421600 1 0 $X=525130 $Y=418640
X2387 1 2 1543 405 1582 ICV_35 $T=560740 399840 1 0 $X=560550 $Y=396880
X2388 1 2 1585 359 1605 ICV_35 $T=571780 427040 1 0 $X=571590 $Y=424080
X2389 1 2 1587 393 1617 ICV_35 $T=577760 399840 0 0 $X=577570 $Y=399600
X2390 1 2 421 405 1694 ICV_35 $T=614560 383520 0 0 $X=614370 $Y=383280
X2391 1 2 429 378 1719 ICV_35 $T=628820 443360 1 0 $X=628630 $Y=440400
X2392 1 2 430 393 433 ICV_35 $T=632040 378080 0 0 $X=631850 $Y=377840
X2393 1 2 1721 395 1742 ICV_35 $T=641700 394400 0 0 $X=641510 $Y=394160
X2394 1 2 1765 393 1769 ICV_35 $T=660560 399840 0 0 $X=660370 $Y=399600
X2395 1 2 1828 406 1840 ICV_35 $T=693220 383520 0 0 $X=693030 $Y=383280
X2396 1 2 1828 393 1841 ICV_35 $T=693220 399840 0 0 $X=693030 $Y=399600
X2397 1 2 1828 407 1844 ICV_35 $T=693680 383520 1 0 $X=693490 $Y=380560
X2398 1 2 1828 403 1849 ICV_35 $T=694140 388960 0 0 $X=693950 $Y=388720
X2399 1 2 1862 402 1884 ICV_35 $T=709320 383520 1 0 $X=709130 $Y=380560
X2400 1 2 1864 365 1868 ICV_35 $T=709780 405280 0 0 $X=709590 $Y=405040
X2401 1 2 517 13 539 ICV_36 $T=6900 388960 0 0 $X=6710 $Y=388720
X2402 1 2 567 13 589 ICV_36 $T=34040 383520 0 0 $X=33850 $Y=383280
X2403 1 2 635 29 657 ICV_36 $T=66240 410720 0 0 $X=66050 $Y=410480
X2404 1 2 676 28 692 ICV_36 $T=84640 405280 1 0 $X=84450 $Y=402320
X2405 1 2 132 109 853 ICV_36 $T=169280 437920 1 0 $X=169090 $Y=434960
X2406 1 2 932 111 966 ICV_36 $T=224020 416160 1 0 $X=223830 $Y=413200
X2407 1 2 1128 190 1143 ICV_36 $T=314640 399840 1 0 $X=314450 $Y=396880
X2408 1 2 1141 228 1172 ICV_36 $T=331200 421600 0 0 $X=331010 $Y=421360
X2409 1 2 277 211 283 ICV_36 $T=413080 383520 1 0 $X=412890 $Y=380560
X2410 1 2 1470 228 1485 ICV_36 $T=490360 427040 0 0 $X=490170 $Y=426800
X2411 1 2 179 363 369 ICV_36 $T=523480 405280 0 0 $X=523290 $Y=405040
X2412 1 2 1543 395 1560 ICV_36 $T=547860 399840 0 0 $X=547670 $Y=399600
X2413 1 2 385 381 1566 ICV_36 $T=553380 443360 1 0 $X=553190 $Y=440400
X2414 1 2 1580 358 1615 ICV_36 $T=574540 437920 0 0 $X=574350 $Y=437680
X2415 1 2 1658 372 1673 ICV_36 $T=602600 416160 0 0 $X=602410 $Y=415920
X2416 1 2 1747 365 1768 ICV_36 $T=651360 432480 0 0 $X=651170 $Y=432240
X2417 1 2 515 28 545 ICV_37 $T=19780 421600 1 0 $X=19590 $Y=418640
X2418 1 2 5 29 35 ICV_37 $T=19780 443360 1 0 $X=19590 $Y=440400
X2419 1 2 33 10 579 ICV_37 $T=33580 378080 0 0 $X=33390 $Y=377840
X2420 1 2 567 28 581 ICV_37 $T=33580 388960 0 0 $X=33390 $Y=388720
X2421 1 2 38 13 585 ICV_37 $T=33580 437920 0 0 $X=33390 $Y=437680
X2422 1 2 597 30 607 ICV_37 $T=47840 383520 1 0 $X=47650 $Y=380560
X2423 1 2 594 11 608 ICV_37 $T=47840 394400 1 0 $X=47650 $Y=391440
X2424 1 2 637 10 645 ICV_37 $T=75900 394400 1 0 $X=75710 $Y=391440
X2425 1 2 635 28 669 ICV_37 $T=75900 399840 1 0 $X=75710 $Y=396880
X2426 1 2 635 17 663 ICV_37 $T=75900 410720 1 0 $X=75710 $Y=407760
X2427 1 2 631 11 671 ICV_37 $T=75900 427040 1 0 $X=75710 $Y=424080
X2428 1 2 676 13 696 ICV_37 $T=89700 399840 0 0 $X=89510 $Y=399600
X2429 1 2 676 10 682 ICV_37 $T=89700 416160 0 0 $X=89510 $Y=415920
X2430 1 2 664 17 721 ICV_37 $T=103960 383520 1 0 $X=103770 $Y=380560
X2431 1 2 695 13 715 ICV_37 $T=103960 394400 1 0 $X=103770 $Y=391440
X2432 1 2 75 10 78 ICV_37 $T=103960 443360 1 0 $X=103770 $Y=440400
X2433 1 2 711 28 750 ICV_37 $T=117760 427040 0 0 $X=117570 $Y=426800
X2434 1 2 746 29 778 ICV_37 $T=132020 399840 1 0 $X=131830 $Y=396880
X2435 1 2 759 28 771 ICV_37 $T=132020 405280 1 0 $X=131830 $Y=402320
X2436 1 2 759 9 779 ICV_37 $T=132020 410720 1 0 $X=131830 $Y=407760
X2437 1 2 759 11 776 ICV_37 $T=132020 421600 1 0 $X=131830 $Y=418640
X2438 1 2 749 13 781 ICV_37 $T=132020 432480 1 0 $X=131830 $Y=429520
X2439 1 2 108 127 831 ICV_37 $T=160080 437920 1 0 $X=159890 $Y=434960
X2440 1 2 121 124 859 ICV_37 $T=173880 378080 0 0 $X=173690 $Y=377840
X2441 1 2 132 112 858 ICV_37 $T=173880 437920 0 0 $X=173690 $Y=437680
X2442 1 2 855 125 870 ICV_37 $T=188140 405280 1 0 $X=187950 $Y=402320
X2443 1 2 135 124 144 ICV_37 $T=201940 378080 0 0 $X=201750 $Y=377840
X2444 1 2 926 125 935 ICV_37 $T=216200 394400 1 0 $X=216010 $Y=391440
X2445 1 2 926 124 941 ICV_37 $T=216200 399840 1 0 $X=216010 $Y=396880
X2446 1 2 901 124 933 ICV_37 $T=216200 416160 1 0 $X=216010 $Y=413200
X2447 1 2 927 109 970 ICV_37 $T=230000 383520 0 0 $X=229810 $Y=383280
X2448 1 2 926 112 968 ICV_37 $T=230000 388960 0 0 $X=229810 $Y=388720
X2449 1 2 931 125 954 ICV_37 $T=230000 437920 0 0 $X=229810 $Y=437680
X2450 1 2 160 111 1020 ICV_37 $T=258060 383520 0 0 $X=257870 $Y=383280
X2451 1 2 1041 126 1054 ICV_37 $T=272320 405280 1 0 $X=272130 $Y=402320
X2452 1 2 157 109 1056 ICV_37 $T=272320 443360 1 0 $X=272130 $Y=440400
X2453 1 2 1066 126 1081 ICV_37 $T=286120 416160 0 0 $X=285930 $Y=415920
X2454 1 2 1066 127 1110 ICV_37 $T=300380 410720 1 0 $X=300190 $Y=407760
X2455 1 2 179 183 194 ICV_37 $T=314180 378080 0 0 $X=313990 $Y=377840
X2456 1 2 1104 111 1130 ICV_37 $T=314180 416160 0 0 $X=313990 $Y=415920
X2457 1 2 1104 124 1133 ICV_37 $T=314180 421600 0 0 $X=313990 $Y=421360
X2458 1 2 1103 125 1135 ICV_37 $T=314180 427040 0 0 $X=313990 $Y=426800
X2459 1 2 1128 212 1157 ICV_37 $T=328440 394400 1 0 $X=328250 $Y=391440
X2460 1 2 1146 204 1150 ICV_37 $T=328440 432480 1 0 $X=328250 $Y=429520
X2461 1 2 1146 199 1163 ICV_37 $T=328440 437920 1 0 $X=328250 $Y=434960
X2462 1 2 1129 212 242 ICV_37 $T=342240 378080 0 0 $X=342050 $Y=377840
X2463 1 2 1129 211 1177 ICV_37 $T=342240 383520 0 0 $X=342050 $Y=383280
X2464 1 2 1167 184 1187 ICV_37 $T=342240 394400 0 0 $X=342050 $Y=394160
X2465 1 2 1146 224 1189 ICV_37 $T=342240 437920 0 0 $X=342050 $Y=437680
X2466 1 2 1173 202 1208 ICV_37 $T=356500 410720 1 0 $X=356310 $Y=407760
X2467 1 2 1211 196 1245 ICV_37 $T=370300 421600 0 0 $X=370110 $Y=421360
X2468 1 2 1233 224 1227 ICV_37 $T=370300 432480 0 0 $X=370110 $Y=432240
X2469 1 2 248 213 1247 ICV_37 $T=370300 437920 0 0 $X=370110 $Y=437680
X2470 1 2 1256 219 1269 ICV_37 $T=384560 405280 1 0 $X=384370 $Y=402320
X2471 1 2 1259 227 1270 ICV_37 $T=384560 410720 1 0 $X=384370 $Y=407760
X2472 1 2 1233 204 1258 ICV_37 $T=384560 432480 1 0 $X=384370 $Y=429520
X2473 1 2 1282 212 1296 ICV_37 $T=398360 388960 0 0 $X=398170 $Y=388720
X2474 1 2 1282 191 1297 ICV_37 $T=398360 394400 0 0 $X=398170 $Y=394160
X2475 1 2 1282 219 1288 ICV_37 $T=398360 399840 0 0 $X=398170 $Y=399600
X2476 1 2 258 199 1298 ICV_37 $T=398360 432480 0 0 $X=398170 $Y=432240
X2477 1 2 1300 191 1324 ICV_37 $T=412620 405280 1 0 $X=412430 $Y=402320
X2478 1 2 1286 213 1327 ICV_37 $T=412620 421600 1 0 $X=412430 $Y=418640
X2479 1 2 1306 224 1328 ICV_37 $T=412620 432480 1 0 $X=412430 $Y=429520
X2480 1 2 1306 228 1329 ICV_37 $T=412620 437920 1 0 $X=412430 $Y=434960
X2481 1 2 1306 213 1342 ICV_37 $T=426420 427040 0 0 $X=426230 $Y=426800
X2482 1 2 1306 196 1347 ICV_37 $T=426420 432480 0 0 $X=426230 $Y=432240
X2483 1 2 293 212 294 ICV_37 $T=440680 383520 1 0 $X=440490 $Y=380560
X2484 1 2 1340 189 1372 ICV_37 $T=440680 394400 1 0 $X=440490 $Y=391440
X2485 1 2 1364 227 1379 ICV_37 $T=440680 410720 1 0 $X=440490 $Y=407760
X2486 1 2 293 191 303 ICV_37 $T=454480 378080 0 0 $X=454290 $Y=377840
X2487 1 2 293 219 1405 ICV_37 $T=454480 383520 0 0 $X=454290 $Y=383280
X2488 1 2 1407 227 1402 ICV_37 $T=468740 416160 1 0 $X=468550 $Y=413200
X2489 1 2 1407 213 1435 ICV_37 $T=468740 421600 1 0 $X=468550 $Y=418640
X2490 1 2 1400 199 1429 ICV_37 $T=468740 432480 1 0 $X=468550 $Y=429520
X2491 1 2 1400 228 1462 ICV_37 $T=482540 427040 0 0 $X=482350 $Y=426800
X2492 1 2 1470 227 1490 ICV_37 $T=496800 432480 1 0 $X=496610 $Y=429520
X2493 1 2 1517 359 1525 ICV_37 $T=524860 443360 1 0 $X=524670 $Y=440400
X2494 1 2 1519 360 1537 ICV_37 $T=538660 416160 0 0 $X=538470 $Y=415920
X2495 1 2 1519 381 1541 ICV_37 $T=538660 421600 0 0 $X=538470 $Y=421360
X2496 1 2 1517 378 1542 ICV_37 $T=538660 432480 0 0 $X=538470 $Y=432240
X2497 1 2 390 402 1563 ICV_37 $T=552920 383520 1 0 $X=552730 $Y=380560
X2498 1 2 1543 403 1558 ICV_37 $T=552920 388960 1 0 $X=552730 $Y=386000
X2499 1 2 1543 393 1561 ICV_37 $T=552920 399840 1 0 $X=552730 $Y=396880
X2500 1 2 1580 378 1596 ICV_37 $T=566720 437920 0 0 $X=566530 $Y=437680
X2501 1 2 1580 365 1616 ICV_37 $T=580980 432480 1 0 $X=580790 $Y=429520
X2502 1 2 1592 395 1646 ICV_37 $T=594780 388960 0 0 $X=594590 $Y=388720
X2503 1 2 1618 359 1647 ICV_37 $T=594780 416160 0 0 $X=594590 $Y=415920
X2504 1 2 1641 395 1676 ICV_37 $T=609040 399840 1 0 $X=608850 $Y=396880
X2505 1 2 1671 378 1706 ICV_37 $T=622840 427040 0 0 $X=622650 $Y=426800
X2506 1 2 430 405 1729 ICV_37 $T=637100 383520 1 0 $X=636910 $Y=380560
X2507 1 2 1698 357 1717 ICV_37 $T=637100 410720 1 0 $X=636910 $Y=407760
X2508 1 2 1698 372 1722 ICV_37 $T=637100 421600 1 0 $X=636910 $Y=418640
X2509 1 2 429 359 1733 ICV_37 $T=637100 427040 1 0 $X=636910 $Y=424080
X2510 1 2 429 381 1736 ICV_37 $T=637100 443360 1 0 $X=636910 $Y=440400
X2511 1 2 437 393 1759 ICV_37 $T=650900 378080 0 0 $X=650710 $Y=377840
X2512 1 2 437 402 1757 ICV_37 $T=650900 383520 0 0 $X=650710 $Y=383280
X2513 1 2 1721 405 1760 ICV_37 $T=650900 394400 0 0 $X=650710 $Y=394160
X2514 1 2 1730 358 1755 ICV_37 $T=650900 410720 0 0 $X=650710 $Y=410480
X2515 1 2 1747 359 1762 ICV_37 $T=650900 437920 0 0 $X=650710 $Y=437680
X2516 1 2 1765 400 1782 ICV_37 $T=665160 388960 1 0 $X=664970 $Y=386000
X2517 1 2 1765 395 1788 ICV_37 $T=665160 399840 1 0 $X=664970 $Y=396880
X2518 1 2 1747 372 1781 ICV_37 $T=665160 432480 1 0 $X=664970 $Y=429520
X2519 1 2 443 378 446 ICV_37 $T=665160 443360 1 0 $X=664970 $Y=440400
X2520 1 2 1777 365 1814 ICV_37 $T=678960 405280 0 0 $X=678770 $Y=405040
X2521 1 2 1802 365 1808 ICV_37 $T=678960 421600 0 0 $X=678770 $Y=421360
X2522 1 2 1802 358 1815 ICV_37 $T=678960 427040 0 0 $X=678770 $Y=426800
X2523 1 2 1826 357 1836 ICV_37 $T=693220 410720 1 0 $X=693030 $Y=407760
X2524 1 2 536 543 25 ICV_39 $T=20240 383520 1 0 $X=20050 $Y=380560
X2525 1 2 549 543 36 ICV_39 $T=25300 383520 1 0 $X=25110 $Y=380560
X2526 1 2 626 605 16 ICV_39 $T=66700 405280 1 0 $X=66510 $Y=402320
X2527 1 2 639 644 31 ICV_39 $T=70840 432480 1 0 $X=70650 $Y=429520
X2528 1 2 662 648 25 ICV_39 $T=84640 405280 0 0 $X=84450 $Y=405040
X2529 1 2 684 66 34 ICV_39 $T=92460 383520 0 0 $X=92270 $Y=383280
X2530 1 2 738 716 37 ICV_39 $T=117760 405280 1 0 $X=117570 $Y=402320
X2531 1 2 755 732 24 ICV_39 $T=126960 416160 0 0 $X=126770 $Y=415920
X2532 1 2 766 768 37 ICV_39 $T=133400 437920 1 0 $X=133210 $Y=434960
X2533 1 2 783 758 36 ICV_39 $T=140760 388960 0 0 $X=140570 $Y=388720
X2534 1 2 880 138 119 ICV_39 $T=191820 383520 1 0 $X=191630 $Y=380560
X2535 1 2 877 845 131 ICV_39 $T=211140 405280 1 0 $X=210950 $Y=402320
X2536 1 2 933 918 128 ICV_39 $T=218960 421600 1 0 $X=218770 $Y=418640
X2537 1 2 946 951 130 ICV_39 $T=224940 383520 0 0 $X=224750 $Y=383280
X2538 1 2 967 936 118 ICV_39 $T=239200 394400 1 0 $X=239010 $Y=391440
X2539 1 2 973 976 128 ICV_39 $T=239200 427040 1 0 $X=239010 $Y=424080
X2540 1 2 991 990 131 ICV_39 $T=247480 399840 1 0 $X=247290 $Y=396880
X2541 1 2 1029 1019 118 ICV_39 $T=267260 432480 1 0 $X=267070 $Y=429520
X2542 1 2 1040 1038 130 ICV_39 $T=272780 421600 1 0 $X=272590 $Y=418640
X2543 1 2 1042 1019 122 ICV_39 $T=272780 427040 1 0 $X=272590 $Y=424080
X2544 1 2 1110 1079 131 ICV_39 $T=309120 410720 0 0 $X=308930 $Y=410480
X2545 1 2 1137 1144 205 ICV_39 $T=323380 405280 1 0 $X=323190 $Y=402320
X2546 1 2 1177 217 236 ICV_39 $T=344540 388960 0 0 $X=344350 $Y=388720
X2547 1 2 1189 215 180 ICV_39 $T=351440 437920 1 0 $X=351250 $Y=434960
X2548 1 2 1217 1199 220 ICV_39 $T=365240 421600 1 0 $X=365050 $Y=418640
X2549 1 2 1248 1225 237 ICV_39 $T=378580 394400 0 0 $X=378390 $Y=394160
X2550 1 2 1331 282 206 ICV_39 $T=421360 383520 0 0 $X=421170 $Y=383280
X2551 1 2 1329 1323 192 ICV_39 $T=421360 427040 0 0 $X=421170 $Y=426800
X2552 1 2 1343 1323 188 ICV_39 $T=429640 437920 0 0 $X=429450 $Y=437680
X2553 1 2 1413 1414 220 ICV_39 $T=463680 437920 1 0 $X=463490 $Y=434960
X2554 1 2 1424 1403 192 ICV_39 $T=468740 405280 0 0 $X=468550 $Y=405040
X2555 1 2 1435 1403 220 ICV_39 $T=477480 421600 0 0 $X=477290 $Y=421360
X2556 1 2 1460 1443 206 ICV_39 $T=489440 399840 0 0 $X=489250 $Y=399600
X2557 1 2 1459 1443 230 ICV_39 $T=491740 394400 1 0 $X=491550 $Y=391440
X2558 1 2 1575 1553 352 ICV_39 $T=567180 394400 0 0 $X=566990 $Y=394160
X2559 1 2 1599 1586 387 ICV_39 $T=581440 394400 1 0 $X=581250 $Y=391440
X2560 1 2 1635 1638 343 ICV_39 $T=595240 432480 0 0 $X=595050 $Y=432240
X2561 1 2 1696 422 386 ICV_39 $T=624680 383520 0 0 $X=624490 $Y=383280
X2562 1 2 1712 1707 386 ICV_39 $T=632040 399840 1 0 $X=631850 $Y=396880
X2563 1 2 1726 1689 355 ICV_39 $T=645840 421600 0 0 $X=645650 $Y=421360
X2564 1 2 1740 1728 389 ICV_39 $T=651360 388960 0 0 $X=651170 $Y=388720
X2565 1 2 1782 1770 392 ICV_39 $T=669760 388960 0 0 $X=669570 $Y=388720
X2566 1 2 1779 1770 388 ICV_39 $T=669760 399840 0 0 $X=669570 $Y=399600
X2567 1 2 1803 1804 371 ICV_39 $T=679420 432480 0 0 $X=679230 $Y=432240
X2568 1 2 523 18 16 ICV_40 $T=13800 383520 1 0 $X=13610 $Y=380560
X2569 1 2 596 576 34 ICV_40 $T=48300 416160 1 0 $X=48110 $Y=413200
X2570 1 2 608 605 24 ICV_40 $T=62100 399840 0 0 $X=61910 $Y=399600
X2571 1 2 630 605 34 ICV_40 $T=62560 394400 0 0 $X=62370 $Y=394160
X2572 1 2 654 634 31 ICV_40 $T=76360 383520 0 0 $X=76170 $Y=383280
X2573 1 2 641 644 16 ICV_40 $T=76360 432480 1 0 $X=76170 $Y=429520
X2574 1 2 661 644 23 ICV_40 $T=78660 421600 1 0 $X=78470 $Y=418640
X2575 1 2 752 720 23 ICV_40 $T=126040 410720 1 0 $X=125850 $Y=407760
X2576 1 2 784 758 23 ICV_40 $T=141680 394400 1 0 $X=141490 $Y=391440
X2577 1 2 106 87 23 ICV_40 $T=142140 443360 1 0 $X=141950 $Y=440400
X2578 1 2 817 819 119 ICV_40 $T=160540 432480 1 0 $X=160350 $Y=429520
X2579 1 2 143 116 131 ICV_40 $T=201020 388960 1 0 $X=200830 $Y=386000
X2580 1 2 921 140 128 ICV_40 $T=210220 443360 1 0 $X=210030 $Y=440400
X2581 1 2 964 936 123 ICV_40 $T=232760 399840 0 0 $X=232570 $Y=399600
X2582 1 2 1020 165 123 ICV_40 $T=262200 388960 1 0 $X=262010 $Y=386000
X2583 1 2 1021 990 119 ICV_40 $T=262200 410720 1 0 $X=262010 $Y=407760
X2584 1 2 1027 1019 128 ICV_40 $T=266340 421600 1 0 $X=266150 $Y=418640
X2585 1 2 1057 1053 123 ICV_40 $T=280140 394400 0 0 $X=279950 $Y=394160
X2586 1 2 1056 162 118 ICV_40 $T=280140 437920 0 0 $X=279950 $Y=437680
X2587 1 2 1073 1053 131 ICV_40 $T=287040 388960 0 0 $X=286850 $Y=388720
X2588 1 2 1100 1079 118 ICV_40 $T=300840 416160 1 0 $X=300650 $Y=413200
X2589 1 2 1124 1092 119 ICV_40 $T=312340 383520 1 0 $X=312150 $Y=380560
X2590 1 2 1145 217 221 ICV_40 $T=350520 388960 1 0 $X=350330 $Y=386000
X2591 1 2 1191 1183 220 ICV_40 $T=350520 421600 1 0 $X=350330 $Y=418640
X2592 1 2 1251 251 192 ICV_40 $T=379040 432480 0 0 $X=378850 $Y=432240
X2593 1 2 1268 1264 221 ICV_40 $T=396520 399840 1 0 $X=396330 $Y=396880
X2594 1 2 289 282 230 ICV_40 $T=435160 378080 0 0 $X=434970 $Y=377840
X2595 1 2 1358 1350 236 ICV_40 $T=437000 394400 0 0 $X=436810 $Y=394160
X2596 1 2 1361 282 222 ICV_40 $T=442060 388960 0 0 $X=441870 $Y=388720
X2597 1 2 316 305 239 ICV_40 $T=473800 443360 1 0 $X=473610 $Y=440400
X2598 1 2 1462 1414 192 ICV_40 $T=490820 427040 1 0 $X=490630 $Y=424080
X2599 1 2 1479 322 187 ICV_40 $T=497260 443360 1 0 $X=497070 $Y=440400
X2600 1 2 1526 1527 343 ICV_40 $T=532680 432480 0 0 $X=532490 $Y=432240
X2601 1 2 1569 1545 363 ICV_40 $T=567180 405280 0 0 $X=566990 $Y=405040
X2602 1 2 1614 1589 345 ICV_40 $T=588800 427040 0 0 $X=588610 $Y=426800
X2603 1 2 1646 1590 397 ICV_40 $T=599840 383520 0 0 $X=599650 $Y=383280
X2604 1 2 1666 1655 388 ICV_40 $T=609500 405280 1 0 $X=609310 $Y=402320
X2605 1 2 1679 1655 391 ICV_40 $T=616860 388960 0 0 $X=616670 $Y=388720
X2606 1 2 1742 1728 397 ICV_40 $T=649520 394400 1 0 $X=649330 $Y=391440
X2607 1 2 1766 1772 368 ICV_40 $T=661940 421600 0 0 $X=661750 $Y=421360
X2608 1 2 1778 440 366 ICV_40 $T=672980 432480 0 0 $X=672790 $Y=432240
X2609 1 2 1891 1885 389 ICV_40 $T=718520 388960 0 0 $X=718330 $Y=388720
X2610 1 2 1907 464 386 ICV_40 $T=736920 383520 1 0 $X=736730 $Y=380560
X2611 1 2 517 10 540 ICV_41 $T=9660 394400 1 0 $X=9470 $Y=391440
X2612 1 2 38 29 593 ICV_41 $T=41400 437920 0 0 $X=41210 $Y=437680
X2613 1 2 48 13 619 ICV_41 $T=51520 437920 0 0 $X=51330 $Y=437680
X2614 1 2 746 13 784 ICV_41 $T=135700 394400 0 0 $X=135510 $Y=394160
X2615 1 2 793 113 800 ICV_41 $T=148580 388960 0 0 $X=148390 $Y=388720
X2616 1 2 795 111 816 ICV_41 $T=149960 427040 1 0 $X=149770 $Y=424080
X2617 1 2 793 124 839 ICV_41 $T=161920 388960 1 0 $X=161730 $Y=386000
X2618 1 2 848 112 872 ICV_41 $T=177560 416160 1 0 $X=177370 $Y=413200
X2619 1 2 932 112 961 ICV_41 $T=234140 416160 1 0 $X=233950 $Y=413200
X2620 1 2 1014 125 1044 ICV_41 $T=268180 432480 0 0 $X=267990 $Y=432240
X2621 1 2 1072 113 1093 ICV_41 $T=293020 388960 0 0 $X=292830 $Y=388720
X2622 1 2 1129 184 200 ICV_41 $T=318320 383520 1 0 $X=318130 $Y=380560
X2623 1 2 1141 224 1170 ICV_41 $T=331660 410720 0 0 $X=331470 $Y=410480
X2624 1 2 1306 204 1343 ICV_41 $T=423200 437920 1 0 $X=423010 $Y=434960
X2625 1 2 1321 196 1348 ICV_41 $T=430100 421600 1 0 $X=429910 $Y=418640
X2626 1 2 1408 184 1449 ICV_41 $T=477020 388960 1 0 $X=476830 $Y=386000
X2627 1 2 324 190 1468 ICV_41 $T=486220 383520 1 0 $X=486030 $Y=380560
X2628 1 2 390 393 404 ICV_41 $T=548780 378080 0 0 $X=548590 $Y=377840
X2629 1 2 390 395 1557 ICV_41 $T=549240 383520 0 0 $X=549050 $Y=383280
X2630 1 2 1658 359 1669 ICV_41 $T=612720 416160 0 0 $X=612530 $Y=415920
X2631 1 2 1685 400 1715 ICV_41 $T=626520 394400 1 0 $X=626330 $Y=391440
X2632 1 2 1730 360 1749 ICV_41 $T=644920 421600 1 0 $X=644730 $Y=418640
X2633 1 2 1751 357 1771 ICV_41 $T=655040 421600 1 0 $X=654850 $Y=418640
X2634 1 2 1864 359 1890 ICV_41 $T=711160 416160 1 0 $X=710970 $Y=413200
X2635 1 2 1862 393 1908 ICV_41 $T=724500 383520 0 0 $X=724310 $Y=383280
X2636 1 2 1862 403 1909 ICV_41 $T=724500 388960 0 0 $X=724310 $Y=388720
X2637 1 2 3 10 523 ICV_47 $T=5520 378080 0 0 $X=5330 $Y=377840
X2638 1 2 513 11 525 ICV_47 $T=5520 405280 1 0 $X=5330 $Y=402320
X2639 1 2 555 10 591 ICV_47 $T=37260 427040 1 0 $X=37070 $Y=424080
X2640 1 2 38 10 592 ICV_47 $T=37260 443360 1 0 $X=37070 $Y=440400
X2641 1 2 631 30 659 ICV_47 $T=69920 416160 0 0 $X=69730 $Y=415920
X2642 1 2 637 30 678 ICV_47 $T=77740 388960 0 0 $X=77550 $Y=388720
X2643 1 2 712 13 752 ICV_47 $T=118220 405280 0 0 $X=118030 $Y=405040
X2644 1 2 89 9 95 ICV_47 $T=120060 443360 1 0 $X=119870 $Y=440400
X2645 1 2 749 30 769 ICV_47 $T=127420 421600 0 0 $X=127230 $Y=421360
X2646 1 2 746 30 783 ICV_47 $T=132480 394400 1 0 $X=132290 $Y=391440
X2647 1 2 848 126 852 ICV_47 $T=174340 421600 0 0 $X=174150 $Y=421360
X2648 1 2 855 112 895 ICV_47 $T=189520 394400 0 0 $X=189330 $Y=394160
X2649 1 2 927 113 983 ICV_47 $T=235060 388960 1 0 $X=234870 $Y=386000
X2650 1 2 969 124 988 ICV_47 $T=236900 405280 0 0 $X=236710 $Y=405040
X2651 1 2 160 125 164 ICV_47 $T=253000 388960 1 0 $X=252810 $Y=386000
X2652 1 2 157 126 1032 ICV_47 $T=258520 437920 0 0 $X=258330 $Y=437680
X2653 1 2 1041 124 1051 ICV_47 $T=270020 399840 0 0 $X=269830 $Y=399600
X2654 1 2 1050 125 1069 ICV_47 $T=276920 421600 0 0 $X=276730 $Y=421360
X2655 1 2 1066 125 1077 ICV_47 $T=282900 421600 1 0 $X=282710 $Y=418640
X2656 1 2 1076 124 1099 ICV_47 $T=290720 399840 1 0 $X=290530 $Y=396880
X2657 1 2 179 187 197 ICV_47 $T=314640 399840 0 0 $X=314450 $Y=399600
X2658 1 2 179 195 207 ICV_47 $T=319700 410720 1 0 $X=319510 $Y=407760
X2659 1 2 1173 228 1181 ICV_47 $T=340400 410720 1 0 $X=340210 $Y=407760
X2660 1 2 254 189 257 ICV_47 $T=374900 383520 1 0 $X=374710 $Y=380560
X2661 1 2 1300 190 1313 ICV_47 $T=406180 399840 0 0 $X=405990 $Y=399600
X2662 1 2 1300 189 1336 ICV_47 $T=415380 394400 0 0 $X=415190 $Y=394160
X2663 1 2 1353 228 1388 ICV_47 $T=443440 432480 0 0 $X=443250 $Y=432240
X2664 1 2 1364 224 1392 ICV_47 $T=445740 416160 0 0 $X=445550 $Y=415920
X2665 1 2 1377 211 1416 ICV_47 $T=458620 394400 1 0 $X=458430 $Y=391440
X2666 1 2 1407 199 1421 ICV_47 $T=459540 421600 1 0 $X=459350 $Y=418640
X2667 1 2 1407 204 1422 ICV_47 $T=459540 421600 0 0 $X=459350 $Y=421360
X2668 1 2 1431 204 1467 ICV_47 $T=484380 421600 1 0 $X=484190 $Y=418640
X2669 1 2 332 213 1499 ICV_47 $T=499560 437920 0 0 $X=499370 $Y=437680
X2670 1 2 1483 224 1504 ICV_47 $T=509680 416160 1 0 $X=509490 $Y=413200
X2671 1 2 179 355 327 ICV_47 $T=525320 410720 1 0 $X=525130 $Y=407760
X2672 1 2 179 367 376 ICV_47 $T=529000 399840 0 0 $X=528810 $Y=399600
X2673 1 2 179 368 377 ICV_47 $T=529000 405280 1 0 $X=528810 $Y=402320
X2674 1 2 1517 365 1533 ICV_47 $T=534520 432480 1 0 $X=534330 $Y=429520
X2675 1 2 1540 360 1552 ICV_47 $T=546480 432480 0 0 $X=546290 $Y=432240
X2676 1 2 1543 402 1575 ICV_47 $T=557980 399840 0 0 $X=557790 $Y=399600
X2677 1 2 1621 358 1640 ICV_47 $T=588800 432480 1 0 $X=588610 $Y=429520
X2678 1 2 1641 393 1681 ICV_47 $T=610420 399840 0 0 $X=610230 $Y=399600
X2679 1 2 1685 405 1716 ICV_47 $T=627440 399840 0 0 $X=627250 $Y=399600
X2680 1 2 1721 403 1737 ICV_47 $T=638480 388960 0 0 $X=638290 $Y=388720
X2681 1 2 1747 358 1758 ICV_47 $T=649060 437920 1 0 $X=648870 $Y=434960
X2682 1 2 1751 365 1776 ICV_47 $T=657340 416160 0 0 $X=657150 $Y=415920
X2683 1 2 1777 378 1801 ICV_47 $T=667920 410720 0 0 $X=667730 $Y=410480
X2684 1 2 1786 357 1833 ICV_47 $T=690920 437920 0 0 $X=690730 $Y=437680
X2685 1 2 1862 406 1891 ICV_47 $T=710240 388960 1 0 $X=710050 $Y=386000
X2686 1 2 461 393 1907 ICV_47 $T=722660 378080 0 0 $X=722470 $Y=377840
X2687 1 2 1866 405 1911 ICV_47 $T=723120 399840 0 0 $X=722930 $Y=399600
X2688 1 2 538 521 23 ICV_48 $T=15640 405280 1 0 $X=15450 $Y=402320
X2689 1 2 613 615 16 ICV_48 $T=57500 405280 0 0 $X=57310 $Y=405040
X2690 1 2 646 648 16 ICV_48 $T=71760 405280 1 0 $X=71570 $Y=402320
X2691 1 2 757 758 16 ICV_48 $T=127880 394400 1 0 $X=127690 $Y=391440
X2692 1 2 814 120 119 ICV_48 $T=155940 432480 1 0 $X=155750 $Y=429520
X2693 1 2 831 120 131 ICV_48 $T=169740 432480 0 0 $X=169550 $Y=432240
X2694 1 2 869 873 131 ICV_48 $T=184000 394400 1 0 $X=183810 $Y=391440
X2695 1 2 870 873 129 ICV_48 $T=184000 399840 1 0 $X=183810 $Y=396880
X2696 1 2 895 873 119 ICV_48 $T=197800 399840 0 0 $X=197610 $Y=399600
X2697 1 2 953 949 118 ICV_48 $T=225860 410720 0 0 $X=225670 $Y=410480
X2698 1 2 975 980 123 ICV_48 $T=240120 405280 1 0 $X=239930 $Y=402320
X2699 1 2 978 976 130 ICV_48 $T=240120 443360 1 0 $X=239930 $Y=440400
X2700 1 2 1036 165 130 ICV_48 $T=268180 388960 1 0 $X=267990 $Y=386000
X2701 1 2 1037 1038 131 ICV_48 $T=268180 410720 1 0 $X=267990 $Y=407760
X2702 1 2 1169 1168 205 ICV_48 $T=338100 399840 0 0 $X=337910 $Y=399600
X2703 1 2 1193 1183 183 ICV_48 $T=352360 416160 1 0 $X=352170 $Y=413200
X2704 1 2 1333 1334 239 ICV_48 $T=422280 416160 0 0 $X=422090 $Y=415920
X2705 1 2 1415 1399 237 ICV_48 $T=464600 405280 1 0 $X=464410 $Y=402320
X2706 1 2 306 307 239 ICV_48 $T=464600 427040 1 0 $X=464410 $Y=424080
X2707 1 2 1534 1516 366 ICV_48 $T=548780 421600 1 0 $X=548590 $Y=418640
X2708 1 2 1565 1550 366 ICV_48 $T=562580 427040 0 0 $X=562390 $Y=426800
X2709 1 2 1659 1643 343 ICV_48 $T=604900 437920 1 0 $X=604710 $Y=434960
X2710 1 2 1687 1689 345 ICV_48 $T=618700 405280 0 0 $X=618510 $Y=405040
X2711 1 2 1688 1667 367 ICV_48 $T=618700 410720 0 0 $X=618510 $Y=410480
X2712 1 2 1716 1707 388 ICV_48 $T=632960 405280 1 0 $X=632770 $Y=402320
X2713 1 2 1769 1770 386 ICV_48 $T=661020 405280 1 0 $X=660830 $Y=402320
X2714 1 2 1797 1799 345 ICV_48 $T=674820 399840 0 0 $X=674630 $Y=399600
X2715 1 2 1824 447 386 ICV_48 $T=689080 388960 1 0 $X=688890 $Y=386000
X2716 1 2 1846 1851 397 ICV_48 $T=702880 394400 0 0 $X=702690 $Y=394160
X2717 1 2 564 29 587 582 580 16 ICV_49 $T=33120 405280 1 0 $X=32930 $Y=402320
X2718 1 2 795 109 811 816 819 123 ICV_49 $T=146280 421600 0 0 $X=146090 $Y=421360
X2719 1 2 874 126 882 882 888 130 ICV_49 $T=185840 388960 0 0 $X=185650 $Y=388720
X2720 1 2 965 127 1004 982 980 129 ICV_49 $T=243340 410720 0 0 $X=243150 $Y=410480
X2721 1 2 965 124 1013 1013 980 128 ICV_49 $T=244720 416160 1 0 $X=244530 $Y=413200
X2722 1 2 1023 125 1059 1059 1038 129 ICV_49 $T=272780 416160 1 0 $X=272590 $Y=413200
X2723 1 2 1066 113 1106 1106 1079 122 ICV_49 $T=294860 410720 0 0 $X=294670 $Y=410480
X2724 1 2 1072 125 1121 1118 1097 131 ICV_49 $T=300840 394400 1 0 $X=300650 $Y=391440
X2725 1 2 1128 189 1142 1121 1092 129 ICV_49 $T=314640 388960 0 0 $X=314450 $Y=388720
X2726 1 2 1233 199 1279 1279 1223 183 ICV_49 $T=385020 427040 1 0 $X=384830 $Y=424080
X2727 1 2 1286 227 1310 1302 1305 183 ICV_49 $T=402960 421600 0 0 $X=402770 $Y=421360
X2728 1 2 277 184 1361 1360 282 205 ICV_49 $T=426880 383520 0 0 $X=426690 $Y=383280
X2729 1 2 1353 204 1385 1385 1371 188 ICV_49 $T=441140 437920 1 0 $X=440950 $Y=434960
X2730 1 2 1618 372 1653 1653 1637 371 ICV_49 $T=592940 416160 1 0 $X=592750 $Y=413200
X2731 1 2 1641 403 1654 1629 1586 397 ICV_49 $T=595240 394400 0 0 $X=595050 $Y=394160
X2732 1 2 1802 360 1812 1815 1810 368 ICV_49 $T=675280 432480 1 0 $X=675090 $Y=429520
X2733 1 2 1826 359 1855 1831 1842 343 ICV_49 $T=693680 421600 1 0 $X=693490 $Y=418640
X2734 1 2 1864 378 1906 1906 1869 366 ICV_49 $T=720360 410720 0 0 $X=720170 $Y=410480
X2735 1 2 1866 403 1910 1892 1865 389 ICV_49 $T=721740 394400 1 0 $X=721550 $Y=391440
X2736 1 2 518 521 16 513 13 538 ICV_51 $T=8740 405280 0 0 $X=8550 $Y=405040
X2737 1 2 552 554 25 555 13 569 ICV_51 $T=25300 432480 1 0 $X=25110 $Y=429520
X2738 1 2 660 648 24 637 29 680 ICV_51 $T=78200 394400 0 0 $X=78010 $Y=394160
X2739 1 2 670 673 25 676 9 689 ICV_51 $T=82800 416160 1 0 $X=82610 $Y=413200
X2740 1 2 679 66 25 68 29 705 ICV_51 $T=90160 378080 0 0 $X=89970 $Y=377840
X2741 1 2 741 87 24 89 11 741 ICV_51 $T=117760 437920 1 0 $X=117570 $Y=434960
X2742 1 2 765 87 31 89 17 765 ICV_51 $T=132480 437920 0 0 $X=132290 $Y=437680
X2743 1 2 769 768 36 749 9 790 ICV_51 $T=134780 427040 1 0 $X=134590 $Y=424080
X2744 1 2 959 147 123 957 126 978 ICV_51 $T=229540 437920 1 0 $X=229350 $Y=434960
X2745 1 2 961 949 119 965 125 982 ICV_51 $T=231840 410720 0 0 $X=231650 $Y=410480
X2746 1 2 966 949 123 965 126 986 ICV_51 $T=233220 416160 0 0 $X=233030 $Y=415920
X2747 1 2 970 951 118 984 109 993 ICV_51 $T=239200 388960 0 0 $X=239010 $Y=388720
X2748 1 2 1047 165 119 169 113 1068 ICV_51 $T=273700 378080 0 0 $X=273510 $Y=377840
X2749 1 2 1089 1092 131 1072 111 1125 ICV_51 $T=300380 383520 0 0 $X=300190 $Y=383280
X2750 1 2 1151 1152 187 1141 227 1171 ICV_51 $T=329820 416160 1 0 $X=329630 $Y=413200
X2751 1 2 1208 1183 187 1211 213 1232 ICV_51 $T=358800 410720 0 0 $X=358610 $Y=410480
X2752 1 2 1258 1223 188 1233 213 1280 ICV_51 $T=383640 427040 0 0 $X=383450 $Y=426800
X2753 1 2 1372 1350 209 1377 212 1391 ICV_51 $T=442980 394400 0 0 $X=442790 $Y=394160
X2754 1 2 1402 1403 239 1407 224 1420 ICV_51 $T=456780 416160 1 0 $X=456590 $Y=413200
X2755 1 2 1478 1480 239 1483 227 1478 ICV_51 $T=495880 410720 0 0 $X=495690 $Y=410480
X2756 1 2 1484 323 230 324 184 1501 ICV_51 $T=499100 383520 0 0 $X=498910 $Y=383280
X2757 1 2 1515 1516 363 1519 365 1515 ICV_51 $T=523480 416160 0 0 $X=523290 $Y=415920
X2758 1 2 1642 1637 345 1641 405 1666 ICV_51 $T=597540 399840 0 0 $X=597350 $Y=399600
X2759 1 2 1668 1667 345 1658 365 1693 ICV_51 $T=610880 410720 1 0 $X=610690 $Y=407760
X2760 1 2 1669 1667 355 1658 357 1688 ICV_51 $T=611340 416160 1 0 $X=611150 $Y=413200
X2761 1 2 1704 1707 387 430 395 1725 ICV_51 $T=629740 383520 0 0 $X=629550 $Y=383280
X2762 1 2 1705 1689 343 1698 365 1724 ICV_51 $T=629740 410720 0 0 $X=629550 $Y=410480
X2763 1 2 1722 1689 371 1730 372 1746 ICV_51 $T=639400 416160 0 0 $X=639210 $Y=415920
X2764 1 2 1757 439 352 1765 403 1775 ICV_51 $T=656420 388960 0 0 $X=656230 $Y=388720
X2765 1 2 1775 1770 387 1777 381 1797 ICV_51 $T=664240 405280 0 0 $X=664050 $Y=405040
X2766 1 2 1863 1865 352 1866 402 1863 ICV_51 $T=708400 399840 1 0 $X=708210 $Y=396880
X2767 1 2 569 554 23 ICV_52 $T=35880 427040 0 0 $X=35690 $Y=426800
X2768 1 2 600 576 25 ICV_52 $T=48300 410720 1 0 $X=48110 $Y=407760
X2769 1 2 614 52 24 ICV_52 $T=77740 437920 0 0 $X=77550 $Y=437680
X2770 1 2 728 720 24 ICV_52 $T=112240 410720 0 0 $X=112050 $Y=410480
X2771 1 2 764 758 25 ICV_52 $T=134780 383520 0 0 $X=134590 $Y=383280
X2772 1 2 782 758 24 ICV_52 $T=140300 383520 0 0 $X=140110 $Y=383280
X2773 1 2 839 802 128 ICV_52 $T=168360 388960 0 0 $X=168170 $Y=388720
X2774 1 2 1004 980 131 ICV_52 $T=258520 410720 0 0 $X=258330 $Y=410480
X2775 1 2 1049 165 122 ICV_52 $T=276000 388960 1 0 $X=275810 $Y=386000
X2776 1 2 1070 1067 128 ICV_52 $T=288420 432480 1 0 $X=288230 $Y=429520
X2777 1 2 1077 1079 129 ICV_52 $T=308660 416160 0 0 $X=308470 $Y=415920
X2778 1 2 1123 1107 129 ICV_52 $T=313260 421600 1 0 $X=313070 $Y=418640
X2779 1 2 1235 1225 236 ICV_52 $T=373060 394400 0 0 $X=372870 $Y=394160
X2780 1 2 1283 1274 187 ICV_52 $T=399740 410720 0 0 $X=399550 $Y=410480
X2781 1 2 1351 1334 220 ICV_52 $T=432860 405280 0 0 $X=432670 $Y=405040
X2782 1 2 1379 1380 239 ICV_52 $T=448960 399840 0 0 $X=448770 $Y=399600
X2783 1 2 1467 1447 188 ICV_52 $T=494500 421600 0 0 $X=494310 $Y=421360
X2784 1 2 349 336 183 ICV_52 $T=519340 443360 1 0 $X=519150 $Y=440400
X2785 1 2 1573 398 388 ICV_52 $T=568100 378080 0 0 $X=567910 $Y=377840
X2786 1 2 1665 1655 352 ICV_52 $T=611340 388960 0 0 $X=611150 $Y=388720
X2787 1 2 1709 1707 397 ICV_52 $T=631580 405280 0 0 $X=631390 $Y=405040
X2788 1 2 ICV_54 $T=33580 427040 0 0 $X=33390 $Y=426800
X2789 1 2 ICV_54 $T=61640 427040 0 0 $X=61450 $Y=426800
X2790 1 2 ICV_54 $T=117760 410720 0 0 $X=117570 $Y=410480
X2791 1 2 ICV_54 $T=145820 410720 0 0 $X=145630 $Y=410480
X2792 1 2 ICV_54 $T=188140 410720 1 0 $X=187950 $Y=407760
X2793 1 2 ICV_54 $T=300380 405280 1 0 $X=300190 $Y=402320
X2794 1 2 ICV_54 $T=342240 388960 0 0 $X=342050 $Y=388720
X2795 1 2 ICV_54 $T=412620 399840 1 0 $X=412430 $Y=396880
X2796 1 2 ICV_54 $T=426420 394400 0 0 $X=426230 $Y=394160
X2797 1 2 ICV_54 $T=440680 432480 1 0 $X=440490 $Y=429520
X2798 1 2 ICV_54 $T=510600 437920 0 0 $X=510410 $Y=437680
X2799 1 2 ICV_54 $T=524860 388960 1 0 $X=524670 $Y=386000
X2800 1 2 ICV_54 $T=609040 416160 1 0 $X=608850 $Y=413200
X2801 1 2 ICV_54 $T=609040 443360 1 0 $X=608850 $Y=440400
X2802 1 2 ICV_54 $T=637100 399840 1 0 $X=636910 $Y=396880
X2803 1 2 ICV_54 $T=650900 416160 0 0 $X=650710 $Y=415920
X2804 1 2 27 2 107 1 sky130_fd_sc_hd__clkbuf_16 $T=143060 405280 1 0 $X=142870 $Y=402320
X2805 1 2 181 2 190 1 sky130_fd_sc_hd__clkbuf_16 $T=314180 405280 1 0 $X=313990 $Y=402320
X2806 1 2 208 2 219 1 sky130_fd_sc_hd__clkbuf_16 $T=328900 405280 1 0 $X=328710 $Y=402320
X2807 1 2 14 2 232 1 sky130_fd_sc_hd__clkbuf_16 $T=331200 405280 0 0 $X=331010 $Y=405040
X2808 1 2 238 2 111 1 sky130_fd_sc_hd__clkbuf_16 $T=341320 388960 1 0 $X=341130 $Y=386000
X2809 1 2 246 2 126 1 sky130_fd_sc_hd__clkbuf_16 $T=356960 388960 1 0 $X=356770 $Y=386000
X2810 1 2 27 2 353 1 sky130_fd_sc_hd__clkbuf_16 $T=516580 421600 0 0 $X=516390 $Y=421360
X2811 1 2 424 2 405 1 sky130_fd_sc_hd__clkbuf_16 $T=615480 405280 1 0 $X=615290 $Y=402320
X2812 1 2 432 2 393 1 sky130_fd_sc_hd__clkbuf_16 $T=639400 399840 0 0 $X=639210 $Y=399600
X2813 1 2 442 2 395 1 sky130_fd_sc_hd__clkbuf_16 $T=665620 405280 1 0 $X=665430 $Y=402320
X2814 1 2 449 2 402 1 sky130_fd_sc_hd__clkbuf_16 $T=679420 399840 1 0 $X=679230 $Y=396880
X2815 1 2 658 634 34 ICV_56 $T=77740 388960 1 0 $X=77550 $Y=386000
X2816 1 2 689 683 25 ICV_56 $T=96600 416160 1 0 $X=96410 $Y=413200
X2817 1 2 703 66 37 ICV_56 $T=100280 388960 0 0 $X=100090 $Y=388720
X2818 1 2 776 773 24 ICV_56 $T=138460 421600 0 0 $X=138270 $Y=421360
X2819 1 2 989 990 123 ICV_56 $T=247480 405280 1 0 $X=247290 $Y=402320
X2820 1 2 1052 1053 122 ICV_56 $T=278760 388960 0 0 $X=278570 $Y=388720
X2821 1 2 1175 217 237 ICV_56 $T=341780 383520 1 0 $X=341590 $Y=380560
X2822 1 2 1244 1239 188 ICV_56 $T=377200 416160 1 0 $X=377010 $Y=413200
X2823 1 2 1270 1274 239 ICV_56 $T=391460 405280 0 0 $X=391270 $Y=405040
X2824 1 2 1287 1274 183 ICV_56 $T=401580 421600 1 0 $X=401390 $Y=418640
X2825 1 2 1296 1290 230 ICV_56 $T=405720 383520 1 0 $X=405530 $Y=380560
X2826 1 2 1355 1334 188 ICV_56 $T=441140 421600 1 0 $X=440950 $Y=418640
X2827 1 2 1474 323 237 ICV_56 $T=503700 394400 0 0 $X=503510 $Y=394160
X2828 1 2 411 413 363 ICV_56 $T=573620 443360 1 0 $X=573430 $Y=440400
X2829 1 2 1744 1754 367 ICV_56 $T=654120 405280 1 0 $X=653930 $Y=402320
X2830 1 2 1832 1842 371 ICV_56 $T=700120 416160 0 0 $X=699930 $Y=415920
X2831 1 2 1871 1874 371 ICV_56 $T=713920 432480 1 0 $X=713730 $Y=429520
X2832 1 2 1915 1865 391 ICV_56 $T=736000 394400 1 0 $X=735810 $Y=391440
X2833 1 2 121 113 826 826 116 122 121 112 813 821 116 123 ICV_57 $T=160540 378080 0 0 $X=160350 $Y=377840
X2834 1 2 794 126 827 827 798 130 794 127 828 836 798 129 ICV_57 $T=160540 394400 0 0 $X=160350 $Y=394160
X2835 1 2 792 127 833 833 809 131 792 124 834 834 809 128 ICV_57 $T=161000 405280 0 0 $X=160810 $Y=405040
X2836 1 2 846 126 864 864 845 130 846 125 842 865 845 122 ICV_57 $T=174800 399840 0 0 $X=174610 $Y=399600
X2837 1 2 846 111 891 881 873 130 846 112 892 891 845 123 ICV_57 $T=190440 405280 0 0 $X=190250 $Y=405040
X2838 1 2 901 125 911 911 918 129 879 109 912 912 890 118 ICV_57 $T=202400 416160 0 0 $X=202210 $Y=415920
X2839 1 2 879 126 914 914 890 130 879 125 915 915 890 129 ICV_57 $T=202400 427040 0 0 $X=202210 $Y=426800
X2840 1 2 137 109 919 898 890 131 137 112 920 920 140 119 ICV_57 $T=203780 432480 0 0 $X=203590 $Y=432240
X2841 1 2 258 227 1271 1271 264 239 258 224 1272 1272 264 180 ICV_57 $T=385020 432480 0 0 $X=384830 $Y=432240
X2842 1 2 1483 204 1493 1493 1480 188 1483 228 1494 1494 1480 192 ICV_57 $T=498640 416160 0 0 $X=498450 $Y=415920
X2843 1 2 1483 199 1511 1511 1480 183 1483 196 1512 1512 1480 195 ICV_57 $T=511980 416160 0 0 $X=511790 $Y=415920
X2844 1 2 1698 378 1703 1697 1667 366 1698 360 1705 431 1643 366 ICV_57 $T=624220 416160 0 0 $X=624030 $Y=415920
X2845 1 2 1671 358 1710 1710 1690 368 1671 372 1711 1711 1690 371 ICV_57 $T=624220 432480 0 0 $X=624030 $Y=432240
X2846 1 2 429 365 1734 1734 434 363 429 360 1735 1735 434 343 ICV_57 $T=637560 432480 0 0 $X=637370 $Y=432240
X2847 1 2 1857 358 1895 1895 1878 368 1857 381 1896 1896 1878 345 ICV_57 $T=721740 421600 0 0 $X=721550 $Y=421360
X2848 1 2 1857 357 1898 1898 1878 367 1857 378 1899 1899 1878 366 ICV_57 $T=722200 416160 0 0 $X=722010 $Y=415920
X2849 1 2 1859 357 1902 1882 1874 355 1859 378 1903 1902 1874 367 ICV_57 $T=722660 432480 0 0 $X=722470 $Y=432240
X2850 1 2 460 358 1904 1904 462 368 460 378 1905 1905 462 366 ICV_57 $T=722660 437920 0 0 $X=722470 $Y=437680
X2851 1 2 594 30 610 610 605 36 ICV_58 $T=45540 394400 0 0 $X=45350 $Y=394160
X2852 1 2 604 28 616 591 554 16 ICV_58 $T=48300 421600 1 0 $X=48110 $Y=418640
X2853 1 2 48 9 618 612 52 36 ICV_58 $T=48300 437920 1 0 $X=48110 $Y=434960
X2854 1 2 793 112 849 849 802 119 ICV_58 $T=167440 394400 1 0 $X=167250 $Y=391440
X2855 1 2 932 113 945 945 949 122 ICV_58 $T=213900 416160 0 0 $X=213710 $Y=415920
X2856 1 2 1076 126 1094 1096 1097 118 ICV_58 $T=286580 405280 0 0 $X=286390 $Y=405040
X2857 1 2 1259 204 1276 1276 1274 188 ICV_58 $T=382260 416160 0 0 $X=382070 $Y=415920
X2858 1 2 272 204 1335 1335 276 188 ICV_58 $T=413080 443360 1 0 $X=412890 $Y=440400
X2859 1 2 1306 227 1344 1347 1323 195 ICV_58 $T=420440 432480 1 0 $X=420250 $Y=429520
X2860 1 2 332 196 1513 1513 336 195 ICV_58 $T=509680 437920 1 0 $X=509490 $Y=434960
X2861 1 2 1539 359 1559 1547 1545 366 ICV_58 $T=546480 410720 0 0 $X=546290 $Y=410480
X2862 1 2 1585 357 1598 1598 1597 367 ICV_58 $T=567180 410720 0 0 $X=566990 $Y=410480
X2863 1 2 1747 360 1764 1764 440 343 ICV_58 $T=649060 432480 1 0 $X=648870 $Y=429520
X2864 1 2 1784 400 1806 1806 447 392 ICV_58 $T=672980 388960 1 0 $X=672790 $Y=386000
X2865 1 2 1777 357 1809 1814 1799 363 ICV_58 $T=674820 410720 1 0 $X=674630 $Y=407760
X2866 1 2 460 365 1883 463 462 371 ICV_58 $T=706560 443360 1 0 $X=706370 $Y=440400
X2867 1 2 1857 365 1888 1888 1878 363 ICV_58 $T=707480 416160 0 0 $X=707290 $Y=415920
X2868 1 2 1866 393 1913 1913 1865 386 ICV_58 $T=721740 399840 1 0 $X=721550 $Y=396880
X2869 1 2 513 28 557 560 521 36 ICV_59 $T=19780 399840 1 0 $X=19590 $Y=396880
X2870 1 2 594 13 609 609 605 23 ICV_59 $T=47840 399840 1 0 $X=47650 $Y=396880
X2871 1 2 676 29 697 692 683 34 ICV_59 $T=89700 405280 0 0 $X=89510 $Y=405040
X2872 1 2 665 11 698 690 673 34 ICV_59 $T=89700 427040 0 0 $X=89510 $Y=426800
X2873 1 2 795 124 830 830 819 128 ICV_59 $T=160080 427040 1 0 $X=159890 $Y=424080
X2874 1 2 793 126 861 861 802 130 ICV_59 $T=173880 388960 0 0 $X=173690 $Y=388720
X2875 1 2 132 125 862 857 844 130 ICV_59 $T=173880 427040 0 0 $X=173690 $Y=426800
X2876 1 2 901 127 910 910 918 131 ICV_59 $T=201940 410720 0 0 $X=201750 $Y=410480
X2877 1 2 931 113 943 943 147 122 ICV_59 $T=216200 432480 1 0 $X=216010 $Y=429520
X2878 1 2 146 127 994 994 158 131 ICV_59 $T=244260 383520 1 0 $X=244070 $Y=380560
X2879 1 2 160 124 1025 1025 165 128 ICV_59 $T=258060 378080 0 0 $X=257870 $Y=377840
X2880 1 2 969 113 1026 1026 990 122 ICV_59 $T=258060 399840 0 0 $X=257870 $Y=399600
X2881 1 2 1103 124 1111 1111 1102 128 ICV_59 $T=300380 432480 1 0 $X=300190 $Y=429520
X2882 1 2 1129 190 1160 1160 217 206 ICV_59 $T=328440 383520 1 0 $X=328250 $Y=380560
X2883 1 2 1211 228 1243 1241 1239 180 ICV_59 $T=370300 410720 0 0 $X=370110 $Y=410480
X2884 1 2 1233 202 1246 1246 1223 187 ICV_59 $T=370300 427040 0 0 $X=370110 $Y=426800
X2885 1 2 258 202 1299 1299 264 187 ICV_59 $T=398360 437920 0 0 $X=398170 $Y=437680
X2886 1 2 1286 202 1326 1326 1305 187 ICV_59 $T=412620 410720 1 0 $X=412430 $Y=407760
X2887 1 2 1400 227 1461 1461 1414 239 ICV_59 $T=482540 421600 0 0 $X=482350 $Y=421360
X2888 1 2 1470 204 1491 1491 1487 188 ICV_59 $T=496800 427040 1 0 $X=496610 $Y=424080
X2889 1 2 1470 199 1507 1507 1487 183 ICV_59 $T=510600 427040 0 0 $X=510410 $Y=426800
X2890 1 2 1585 378 1623 1623 1597 366 ICV_59 $T=580980 416160 1 0 $X=580790 $Y=413200
X2891 1 2 415 402 1650 1650 417 352 ICV_59 $T=594780 378080 0 0 $X=594590 $Y=377840
X2892 1 2 1751 381 1789 1776 1772 363 ICV_59 $T=665160 416160 1 0 $X=664970 $Y=413200
X2893 1 2 1777 359 1818 1819 1799 343 ICV_59 $T=678960 410720 0 0 $X=678770 $Y=410480
X2894 1 2 1786 359 1820 1820 1804 355 ICV_59 $T=678960 437920 0 0 $X=678770 $Y=437680
X2895 1 2 1859 372 1871 1827 1810 345 ICV_59 $T=707020 427040 0 0 $X=706830 $Y=426800
X2896 1 2 1859 360 1872 1872 1874 343 ICV_59 $T=707020 432480 0 0 $X=706830 $Y=432240
X2897 1 2 1864 381 1893 1893 1869 345 ICV_59 $T=721280 405280 1 0 $X=721090 $Y=402320
X2898 1 2 515 17 550 550 534 31 ICV_60 $T=18860 410720 0 0 $X=18670 $Y=410480
X2899 1 2 567 17 578 578 580 31 ICV_60 $T=33580 399840 1 0 $X=33390 $Y=396880
X2900 1 2 597 17 606 606 51 31 ICV_60 $T=47380 383520 0 0 $X=47190 $Y=383280
X2901 1 2 631 29 666 666 644 37 ICV_60 $T=75440 427040 0 0 $X=75250 $Y=426800
X2902 1 2 108 126 825 825 120 130 ICV_60 $T=159620 437920 0 0 $X=159430 $Y=437680
X2903 1 2 926 127 938 941 936 128 ICV_60 $T=215740 399840 0 0 $X=215550 $Y=399600
X2904 1 2 169 112 1108 1108 171 119 ICV_60 $T=299920 378080 0 0 $X=299730 $Y=377840
X2905 1 2 1211 199 1242 1242 1239 183 ICV_60 $T=370300 421600 1 0 $X=370110 $Y=418640
X2906 1 2 1256 212 1263 1263 1264 230 ICV_60 $T=384100 388960 0 0 $X=383910 $Y=388720
X2907 1 2 258 213 1293 1298 264 183 ICV_60 $T=398360 437920 1 0 $X=398170 $Y=434960
X2908 1 2 1286 224 1308 1308 1305 180 ICV_60 $T=405260 410720 0 0 $X=405070 $Y=410480
X2909 1 2 1408 211 1426 1416 1399 236 ICV_60 $T=463680 388960 0 0 $X=463490 $Y=388720
X2910 1 2 1408 219 1442 1442 312 237 ICV_60 $T=471960 383520 1 0 $X=471770 $Y=380560
X2911 1 2 1456 189 1473 1473 323 209 ICV_60 $T=487600 388960 0 0 $X=487410 $Y=388720
X2912 1 2 1470 202 1506 1506 1487 187 ICV_60 $T=510600 432480 1 0 $X=510410 $Y=429520
X2913 1 2 1592 407 1649 1649 1590 391 ICV_60 $T=594780 383520 1 0 $X=594590 $Y=380560
X2914 1 2 460 360 1875 1875 462 343 ICV_60 $T=708400 437920 0 0 $X=708210 $Y=437680
X2915 1 2 39 580 ICV_61 $T=44160 383520 0 0 $X=43970 $Y=383280
X2916 1 2 46 52 ICV_61 $T=58420 432480 0 0 $X=58230 $Y=432240
X2917 1 2 47 615 ICV_61 $T=62100 405280 0 0 $X=61910 $Y=405040
X2918 1 2 57 644 ICV_61 $T=78660 416160 0 0 $X=78470 $Y=415920
X2919 1 2 73 951 ICV_61 $T=233220 383520 1 0 $X=233030 $Y=380560
X2920 1 2 76 1079 ICV_61 $T=293940 416160 0 0 $X=293750 $Y=415920
X2921 1 2 152 1092 ICV_61 $T=300840 388960 1 0 $X=300650 $Y=386000
X2922 1 2 235 1152 ICV_61 $T=339020 416160 0 0 $X=338830 $Y=415920
X2923 1 2 231 215 ICV_61 $T=343620 427040 1 0 $X=343430 $Y=424080
X2924 1 2 256 1264 ICV_61 $T=392380 405280 1 0 $X=392190 $Y=402320
X2925 1 2 292 1350 ICV_61 $T=445280 399840 1 0 $X=445090 $Y=396880
X2926 1 2 311 1414 ICV_61 $T=479320 427040 0 0 $X=479130 $Y=426800
X2927 1 2 231 1550 ICV_61 $T=553380 432480 1 0 $X=553190 $Y=429520
X2928 1 2 320 439 ICV_61 $T=658720 383520 0 0 $X=658530 $Y=383280
X2929 1 2 328 1799 ICV_61 $T=675740 405280 0 0 $X=675550 $Y=405040
X2930 1 2 333 1851 ICV_61 $T=707940 394400 1 0 $X=707750 $Y=391440
X2931 1 2 541 533 31 ICV_62 $T=20700 432480 1 0 $X=20510 $Y=429520
X2932 1 2 651 58 23 ICV_62 $T=76360 437920 1 0 $X=76170 $Y=434960
X2933 1 2 696 683 23 ICV_62 $T=96140 405280 1 0 $X=95950 $Y=402320
X2934 1 2 687 683 24 ICV_62 $T=101660 405280 0 0 $X=101470 $Y=405040
X2935 1 2 710 673 31 ICV_62 $T=104420 421600 1 0 $X=104230 $Y=418640
X2936 1 2 719 71 24 ICV_62 $T=110860 432480 0 0 $X=110670 $Y=432240
X2937 1 2 714 716 24 ICV_62 $T=123280 394400 1 0 $X=123090 $Y=391440
X2938 1 2 781 768 23 ICV_62 $T=138920 432480 0 0 $X=138730 $Y=432240
X2939 1 2 791 768 24 ICV_62 $T=151340 432480 1 0 $X=151150 $Y=429520
X2940 1 2 899 890 122 ICV_62 $T=197800 427040 1 0 $X=197610 $Y=424080
X2941 1 2 1015 990 129 ICV_62 $T=257600 410720 1 0 $X=257410 $Y=407760
X2942 1 2 1131 1107 131 ICV_62 $T=323840 427040 1 0 $X=323650 $Y=424080
X2943 1 2 1136 1144 222 ICV_62 $T=328900 388960 1 0 $X=328710 $Y=386000
X2944 1 2 216 218 187 ICV_62 $T=329820 443360 1 0 $X=329630 $Y=440400
X2945 1 2 1163 215 183 ICV_62 $T=337640 432480 0 0 $X=337450 $Y=432240
X2946 1 2 1195 218 239 ICV_62 $T=356960 437920 1 0 $X=356770 $Y=434960
X2947 1 2 1243 1239 192 ICV_62 $T=377660 405280 1 0 $X=377470 $Y=402320
X2948 1 2 1275 1274 220 ICV_62 $T=392380 410720 0 0 $X=392190 $Y=410480
X2949 1 2 1307 1290 209 ICV_62 $T=410320 383520 0 0 $X=410130 $Y=383280
X2950 1 2 1337 1317 222 ICV_62 $T=426880 405280 0 0 $X=426690 $Y=405040
X2951 1 2 1346 1334 180 ICV_62 $T=436080 416160 1 0 $X=435890 $Y=413200
X2952 1 2 1387 1371 180 ICV_62 $T=451260 432480 1 0 $X=451070 $Y=429520
X2953 1 2 1396 1399 221 ICV_62 $T=454940 399840 0 0 $X=454750 $Y=399600
X2954 1 2 1410 305 180 ICV_62 $T=469200 443360 1 0 $X=469010 $Y=440400
X2955 1 2 1445 312 206 ICV_62 $T=483000 378080 0 0 $X=482810 $Y=377840
X2956 1 2 1551 1545 367 ICV_62 $T=553840 410720 1 0 $X=553650 $Y=407760
X2957 1 2 1564 401 367 ICV_62 $T=562580 437920 1 0 $X=562390 $Y=434960
X2958 1 2 1567 1550 367 ICV_62 $T=567180 427040 0 0 $X=566990 $Y=426800
X2959 1 2 1625 417 391 ICV_62 $T=590180 383520 1 0 $X=589990 $Y=380560
X2960 1 2 1631 1590 389 ICV_62 $T=595240 383520 0 0 $X=595050 $Y=383280
X2961 1 2 1674 422 352 ICV_62 $T=612260 383520 1 0 $X=612070 $Y=380560
X2962 1 2 1706 1690 366 ICV_62 $T=629740 421600 0 0 $X=629550 $Y=421360
X2963 1 2 1788 1770 397 ICV_62 $T=679420 394400 0 0 $X=679230 $Y=394160
X2964 1 2 1830 1810 371 ICV_62 $T=694600 427040 1 0 $X=694410 $Y=424080
X2965 1 2 1853 1851 388 ICV_62 $T=703800 399840 1 0 $X=703610 $Y=396880
X2966 1 2 1838 1804 345 ICV_62 $T=705180 437920 1 0 $X=704990 $Y=434960
X2967 1 2 624 605 25 ICV_63 $T=59800 399840 1 0 $X=59610 $Y=396880
X2968 1 2 717 71 25 ICV_63 $T=109480 437920 0 0 $X=109290 $Y=437680
X2969 1 2 739 716 36 ICV_63 $T=118220 399840 0 0 $X=118030 $Y=399600
X2970 1 2 858 844 119 ICV_63 $T=179400 437920 1 0 $X=179210 $Y=434960
X2971 1 2 867 844 122 ICV_63 $T=181700 437920 0 0 $X=181510 $Y=437680
X2972 1 2 960 936 122 ICV_63 $T=230460 394400 0 0 $X=230270 $Y=394160
X2973 1 2 1035 1008 122 ICV_63 $T=266800 394400 0 0 $X=266610 $Y=394160
X2974 1 2 1197 1207 222 ICV_63 $T=356960 383520 1 0 $X=356770 $Y=380560
X2975 1 2 1222 1223 192 ICV_63 $T=364780 427040 1 0 $X=364590 $Y=424080
X2976 1 2 1284 1274 192 ICV_63 $T=398820 405280 0 0 $X=398630 $Y=405040
X2977 1 2 1504 1480 180 ICV_63 $T=512440 410720 1 0 $X=512250 $Y=407760
X2978 1 2 1532 1527 345 ICV_63 $T=540040 437920 1 0 $X=539850 $Y=434960
X2979 1 2 1574 398 389 ICV_63 $T=567180 383520 0 0 $X=566990 $Y=383280
X2980 1 2 1610 1590 392 ICV_63 $T=581440 383520 1 0 $X=581250 $Y=380560
X2981 1 2 1844 1851 391 ICV_63 $T=701500 383520 0 0 $X=701310 $Y=383280
X2982 1 2 1841 1851 386 ICV_63 $T=701500 399840 0 0 $X=701310 $Y=399600
X2983 1 2 459 455 345 ICV_63 $T=701500 443360 1 0 $X=701310 $Y=440400
X2984 1 2 555 30 568 514 29 551 ICV_64 $T=19780 427040 1 0 $X=19590 $Y=424080
X2985 1 2 564 9 600 564 13 574 ICV_64 $T=33580 405280 0 0 $X=33390 $Y=405040
X2986 1 2 665 17 710 665 29 681 ICV_64 $T=89700 421600 0 0 $X=89510 $Y=421360
X2987 1 2 931 111 959 931 126 148 ICV_64 $T=216200 443360 1 0 $X=216010 $Y=440400
X2988 1 2 1023 111 1045 969 112 1021 ICV_64 $T=258060 405280 0 0 $X=257870 $Y=405040
X2989 1 2 1141 213 1176 1141 196 1159 ICV_64 $T=328440 427040 1 0 $X=328250 $Y=424080
X2990 1 2 1185 204 1202 1146 227 1188 ICV_64 $T=342240 432480 0 0 $X=342050 $Y=432240
X2991 1 2 268 211 1311 268 219 273 ICV_64 $T=398360 378080 0 0 $X=398170 $Y=377840
X2992 1 2 1286 196 1312 1259 199 1287 ICV_64 $T=398360 416160 0 0 $X=398170 $Y=415920
X2993 1 2 1377 191 1396 1340 219 1374 ICV_64 $T=440680 405280 1 0 $X=440490 $Y=402320
X2994 1 2 1364 202 1397 1364 213 1381 ICV_64 $T=440680 416160 1 0 $X=440490 $Y=413200
X2995 1 2 1456 190 1481 1427 212 1459 ICV_64 $T=482540 394400 0 0 $X=482350 $Y=394160
X2996 1 2 1456 184 339 1456 212 1484 ICV_64 $T=496800 394400 1 0 $X=496610 $Y=391440
X2997 1 2 385 372 1549 1517 381 1532 ICV_64 $T=538660 437920 0 0 $X=538470 $Y=437680
X2998 1 2 418 360 1659 418 365 1651 ICV_64 $T=594780 437920 0 0 $X=594590 $Y=437680
X2999 1 2 1658 378 1697 1658 360 1677 ICV_64 $T=609040 421600 1 0 $X=608850 $Y=418640
X3000 1 2 1784 393 1824 1784 405 1816 ICV_64 $T=678960 388960 0 0 $X=678770 $Y=388720
X3001 1 2 7 8 519 ICV_65 $T=6900 416160 0 0 $X=6710 $Y=415920
X3002 1 2 97 8 763 ICV_65 $T=129260 437920 1 0 $X=129070 $Y=434960
X3003 1 2 76 107 1058 ICV_65 $T=280140 421600 1 0 $X=279950 $Y=418640
X3004 1 2 240 232 1180 ICV_65 $T=347300 421600 1 0 $X=347110 $Y=418640
X3005 1 2 263 232 1281 ICV_65 $T=392380 432480 1 0 $X=392190 $Y=429520
X3006 1 2 266 225 267 ICV_65 $T=393300 383520 1 0 $X=393110 $Y=380560
X3007 1 2 285 225 1338 ICV_65 $T=426880 388960 0 0 $X=426690 $Y=388720
X3008 1 2 292 225 1366 ICV_65 $T=437920 410720 1 0 $X=437730 $Y=407760
X3009 1 2 291 232 1365 ICV_65 $T=437920 427040 1 0 $X=437730 $Y=424080
X3010 1 2 328 232 1482 ICV_65 $T=495420 405280 0 0 $X=495230 $Y=405040
X3011 1 2 223 394 1546 ICV_65 $T=550160 399840 1 0 $X=549970 $Y=396880
X3012 1 2 408 353 1572 ICV_65 $T=563500 443360 1 0 $X=563310 $Y=440400
X3013 1 2 279 353 1620 ICV_65 $T=584660 437920 0 0 $X=584470 $Y=437680
X3014 1 2 245 394 1648 ICV_65 $T=598920 399840 1 0 $X=598730 $Y=396880
X3015 1 2 256 394 1686 ICV_65 $T=619160 399840 0 0 $X=618970 $Y=399600
X3016 1 2 274 353 1699 ICV_65 $T=622380 410720 1 0 $X=622190 $Y=407760
X3017 1 2 278 394 1753 ICV_65 $T=651360 399840 0 0 $X=651170 $Y=399600
X3018 1 2 664 9 679 ICV_66 $T=82340 383520 0 0 $X=82150 $Y=383280
X3019 1 2 695 30 739 ICV_66 $T=110400 399840 0 0 $X=110210 $Y=399600
X3020 1 2 746 17 761 ICV_66 $T=124660 388960 1 0 $X=124470 $Y=386000
X3021 1 2 984 127 1012 ICV_66 $T=250700 388960 0 0 $X=250510 $Y=388720
X3022 1 2 1041 109 1071 ICV_66 $T=278760 399840 0 0 $X=278570 $Y=399600
X3023 1 2 1353 213 1367 ICV_66 $T=433320 437920 1 0 $X=433130 $Y=434960
X3024 1 2 1364 196 1393 ICV_66 $T=447120 421600 0 0 $X=446930 $Y=421360
X3025 1 2 1408 212 309 ICV_66 $T=461380 383520 1 0 $X=461190 $Y=380560
X3026 1 2 179 345 354 ICV_66 $T=517500 405280 1 0 $X=517310 $Y=402320
X3027 1 2 1539 378 1547 ICV_66 $T=545560 416160 1 0 $X=545370 $Y=413200
X3028 1 2 1540 381 1548 ICV_66 $T=545560 432480 1 0 $X=545370 $Y=429520
X3029 1 2 385 378 399 ICV_66 $T=545560 443360 1 0 $X=545370 $Y=440400
X3030 1 2 390 406 1574 ICV_66 $T=559360 383520 0 0 $X=559170 $Y=383280
X3031 1 2 1592 403 1607 ICV_66 $T=573620 388960 1 0 $X=573430 $Y=386000
X3032 1 2 1618 357 1633 ICV_66 $T=587420 405280 0 0 $X=587230 $Y=405040
X3033 1 2 1621 378 1634 ICV_66 $T=587420 421600 0 0 $X=587230 $Y=421360
X3034 1 2 1730 357 1744 ICV_66 $T=643540 405280 0 0 $X=643350 $Y=405040
X3035 1 2 94 96 98 99 2 747 1 sky130_fd_sc_hd__and4b_2 $T=128340 378080 0 0 $X=128150 $Y=377840
X3036 1 2 85 83 79 747 2 100 1 sky130_fd_sc_hd__and4b_2 $T=130640 383520 0 0 $X=130450 $Y=383280
X3037 1 2 83 85 79 747 2 101 1 sky130_fd_sc_hd__and4b_2 $T=132480 378080 0 0 $X=132290 $Y=377840
X3038 1 2 79 85 83 747 2 102 1 sky130_fd_sc_hd__and4b_2 $T=132480 383520 1 0 $X=132290 $Y=380560
X3039 1 2 79 85 83 105 2 114 1 sky130_fd_sc_hd__and4b_2 $T=147660 383520 1 0 $X=147470 $Y=380560
X3040 1 2 340 342 341 1505 2 330 1 sky130_fd_sc_hd__and4b_2 $T=513360 383520 0 0 $X=513170 $Y=383280
X3041 1 2 341 340 342 1505 2 344 1 sky130_fd_sc_hd__and4b_2 $T=513820 388960 1 0 $X=513630 $Y=386000
X3042 1 2 342 340 341 346 2 315 1 sky130_fd_sc_hd__and4b_2 $T=516580 383520 1 0 $X=516390 $Y=380560
X3043 1 2 341 340 342 346 2 250 1 sky130_fd_sc_hd__and4b_2 $T=520720 383520 1 0 $X=520530 $Y=380560
X3044 1 2 340 342 341 346 2 318 1 sky130_fd_sc_hd__and4b_2 $T=523020 383520 0 0 $X=522830 $Y=383280
X3045 1 2 96 98 94 361 2 1505 1 sky130_fd_sc_hd__and4b_2 $T=525320 383520 1 0 $X=525130 $Y=380560
X3046 1 2 342 340 341 1505 2 320 1 sky130_fd_sc_hd__and4b_2 $T=525320 399840 1 0 $X=525130 $Y=396880
X3047 1 2 341 340 342 1522 2 300 1 sky130_fd_sc_hd__and4b_2 $T=527620 394400 0 0 $X=527430 $Y=394160
X3048 1 2 342 340 341 1522 2 370 1 sky130_fd_sc_hd__and4b_2 $T=531760 388960 0 0 $X=531570 $Y=388720
X3049 1 2 98 96 94 361 2 1530 1 sky130_fd_sc_hd__and4b_2 $T=532220 383520 1 0 $X=532030 $Y=380560
X3050 1 2 340 342 341 1522 2 373 1 sky130_fd_sc_hd__and4b_2 $T=532220 383520 0 0 $X=532030 $Y=383280
X3051 1 2 94 96 98 361 2 375 1 sky130_fd_sc_hd__and4b_2 $T=534060 378080 0 0 $X=533870 $Y=377840
X3052 1 2 341 340 342 1530 2 383 1 sky130_fd_sc_hd__and4b_2 $T=538200 394400 1 0 $X=538010 $Y=391440
X3053 1 2 340 342 341 1530 2 334 1 sky130_fd_sc_hd__and4b_2 $T=539120 394400 0 0 $X=538930 $Y=394160
X3054 1 2 341 340 342 375 2 333 1 sky130_fd_sc_hd__and4b_2 $T=543260 383520 1 0 $X=543070 $Y=380560
X3055 1 2 340 342 341 375 2 308 1 sky130_fd_sc_hd__and4b_2 $T=544640 378080 0 0 $X=544450 $Y=377840
X3056 1 2 342 340 341 375 2 396 1 sky130_fd_sc_hd__and4b_2 $T=547400 383520 1 0 $X=547210 $Y=380560
X3057 1 2 342 340 341 1530 2 314 1 sky130_fd_sc_hd__and4b_2 $T=547400 388960 0 0 $X=547210 $Y=388720
X3058 1 2 83 85 79 84 2 76 1 sky130_fd_sc_hd__and4_2 $T=118220 378080 0 0 $X=118030 $Y=377840
X3059 1 2 83 85 79 747 2 80 1 sky130_fd_sc_hd__and4_2 $T=126960 383520 0 0 $X=126770 $Y=383280
X3060 1 2 98 96 94 99 2 105 1 sky130_fd_sc_hd__and4_2 $T=146280 383520 0 0 $X=146090 $Y=383280
X3061 1 2 83 85 79 105 2 97 1 sky130_fd_sc_hd__and4_2 $T=149960 383520 0 0 $X=149770 $Y=383280
X3062 1 2 342 340 341 346 2 233 1 sky130_fd_sc_hd__and4_2 $T=523480 388960 0 0 $X=523290 $Y=388720
X3063 1 2 342 340 341 1505 2 292 1 sky130_fd_sc_hd__and4_2 $T=523940 394400 0 0 $X=523750 $Y=394160
X3064 1 2 342 340 341 1522 2 245 1 sky130_fd_sc_hd__and4_2 $T=529460 399840 1 0 $X=529270 $Y=396880
X3065 1 2 342 340 341 375 2 302 1 sky130_fd_sc_hd__and4_2 $T=539120 383520 0 0 $X=538930 $Y=383280
X3066 1 2 342 340 341 1530 2 278 1 sky130_fd_sc_hd__and4_2 $T=546480 399840 1 0 $X=546290 $Y=396880
X3067 1 2 1471 1475 2 221 1 sky130_fd_sc_hd__ebufn_4 $T=494500 399840 0 0 $X=494310 $Y=399600
X3068 1 2 1471 1475 2 206 1 sky130_fd_sc_hd__ebufn_4 $T=497260 405280 1 0 $X=497070 $Y=402320
X3069 1 2 1471 1475 2 209 1 sky130_fd_sc_hd__ebufn_4 $T=497720 394400 0 0 $X=497530 $Y=394160
X3070 1 2 1471 1475 2 188 1 sky130_fd_sc_hd__ebufn_4 $T=498180 405280 0 0 $X=497990 $Y=405040
X3071 1 2 1471 1475 2 237 1 sky130_fd_sc_hd__ebufn_4 $T=503240 405280 1 0 $X=503050 $Y=402320
X3072 1 2 1471 1475 2 220 1 sky130_fd_sc_hd__ebufn_4 $T=504620 405280 0 0 $X=504430 $Y=405040
X3073 1 2 1471 1475 2 192 1 sky130_fd_sc_hd__ebufn_4 $T=506460 410720 1 0 $X=506270 $Y=407760
X3074 1 2 1471 1475 2 230 1 sky130_fd_sc_hd__ebufn_4 $T=511060 394400 0 0 $X=510870 $Y=394160
X3075 1 2 1471 1475 2 205 1 sky130_fd_sc_hd__ebufn_4 $T=511060 399840 0 0 $X=510870 $Y=399600
X3076 1 2 1471 1475 2 239 1 sky130_fd_sc_hd__ebufn_4 $T=511060 405280 0 0 $X=510870 $Y=405040
X3077 1 2 1471 1475 2 343 1 sky130_fd_sc_hd__ebufn_4 $T=511520 405280 1 0 $X=511330 $Y=402320
X3078 1 2 1471 1475 2 236 1 sky130_fd_sc_hd__ebufn_4 $T=511980 394400 1 0 $X=511790 $Y=391440
X3079 1 2 1471 1475 2 222 1 sky130_fd_sc_hd__ebufn_4 $T=512900 388960 0 0 $X=512710 $Y=388720
X3080 1 2 1471 1475 2 352 1 sky130_fd_sc_hd__ebufn_4 $T=516120 399840 1 0 $X=515930 $Y=396880
X3081 1 2 1471 1475 2 195 1 sky130_fd_sc_hd__ebufn_4 $T=517500 405280 0 0 $X=517310 $Y=405040
X3082 1 2 1471 1475 2 187 1 sky130_fd_sc_hd__ebufn_4 $T=517500 410720 1 0 $X=517310 $Y=407760
X3083 1 2 1471 1475 2 183 1 sky130_fd_sc_hd__ebufn_4 $T=517960 394400 0 0 $X=517770 $Y=394160
X3084 1 2 1471 1475 2 355 1 sky130_fd_sc_hd__ebufn_4 $T=518880 416160 1 0 $X=518690 $Y=413200
X3085 1 2 1471 1475 2 180 1 sky130_fd_sc_hd__ebufn_4 $T=519340 410720 0 0 $X=519150 $Y=410480
X3086 1 2 1471 1475 2 368 1 sky130_fd_sc_hd__ebufn_4 $T=531760 416160 1 0 $X=531570 $Y=413200
X3087 1 2 1471 1475 2 367 1 sky130_fd_sc_hd__ebufn_4 $T=539120 405280 1 0 $X=538930 $Y=402320
X3088 1 2 1471 1475 2 366 1 sky130_fd_sc_hd__ebufn_4 $T=539580 416160 1 0 $X=539390 $Y=413200
X3089 1 2 1471 1475 2 386 1 sky130_fd_sc_hd__ebufn_4 $T=540500 399840 1 0 $X=540310 $Y=396880
X3090 1 2 1471 1475 2 371 1 sky130_fd_sc_hd__ebufn_4 $T=540500 410720 0 0 $X=540310 $Y=410480
X3091 1 2 1471 1475 2 387 1 sky130_fd_sc_hd__ebufn_4 $T=541420 388960 0 0 $X=541230 $Y=388720
X3092 1 2 1471 1475 2 388 1 sky130_fd_sc_hd__ebufn_4 $T=541880 399840 0 0 $X=541690 $Y=399600
X3093 1 2 1471 1475 2 345 1 sky130_fd_sc_hd__ebufn_4 $T=541880 405280 0 0 $X=541690 $Y=405040
X3094 1 2 1471 1475 2 363 1 sky130_fd_sc_hd__ebufn_4 $T=541880 410720 1 0 $X=541690 $Y=407760
X3095 1 2 1471 1475 2 389 1 sky130_fd_sc_hd__ebufn_4 $T=542800 394400 1 0 $X=542610 $Y=391440
X3096 1 2 1471 1475 2 391 1 sky130_fd_sc_hd__ebufn_4 $T=543260 388960 1 0 $X=543070 $Y=386000
X3097 1 2 1471 1475 2 392 1 sky130_fd_sc_hd__ebufn_4 $T=543260 394400 0 0 $X=543070 $Y=394160
X3098 1 2 1471 1475 2 397 1 sky130_fd_sc_hd__ebufn_4 $T=545100 405280 1 0 $X=544910 $Y=402320
X3099 1 2 83 85 79 747 2 92 1 sky130_fd_sc_hd__nor4b_2 $T=119600 383520 1 0 $X=119410 $Y=380560
X3100 1 2 83 85 79 105 2 104 1 sky130_fd_sc_hd__nor4b_2 $T=137080 378080 0 0 $X=136890 $Y=377840
X3101 1 2 342 340 341 1505 2 351 1 sky130_fd_sc_hd__nor4b_2 $T=517500 383520 0 0 $X=517310 $Y=383280
X3102 1 2 342 340 341 1522 2 270 1 sky130_fd_sc_hd__nor4b_2 $T=527160 388960 1 0 $X=526970 $Y=386000
X3103 1 2 98 96 94 361 2 1522 1 sky130_fd_sc_hd__nor4b_2 $T=528540 378080 0 0 $X=528350 $Y=377840
X3104 1 2 342 340 341 1530 2 256 1 sky130_fd_sc_hd__nor4b_2 $T=532220 394400 0 0 $X=532030 $Y=394160
X3105 1 2 342 340 341 375 2 379 1 sky130_fd_sc_hd__nor4b_2 $T=539120 378080 0 0 $X=538930 $Y=377840
X3106 1 2 79 83 84 85 2 32 1 sky130_fd_sc_hd__and4bb_2 $T=113160 378080 0 0 $X=112970 $Y=377840
X3107 1 2 79 85 84 83 2 12 1 sky130_fd_sc_hd__and4bb_2 $T=113620 383520 1 0 $X=113430 $Y=380560
X3108 1 2 83 79 747 85 2 90 1 sky130_fd_sc_hd__and4bb_2 $T=121900 378080 0 0 $X=121710 $Y=377840
X3109 1 2 79 85 747 83 2 91 1 sky130_fd_sc_hd__and4bb_2 $T=121900 383520 0 0 $X=121710 $Y=383280
X3110 1 2 79 83 747 85 2 47 1 sky130_fd_sc_hd__and4bb_2 $T=125120 383520 1 0 $X=124930 $Y=380560
X3111 1 2 79 83 105 85 2 103 1 sky130_fd_sc_hd__and4bb_2 $T=138460 383520 1 0 $X=138270 $Y=380560
X3112 1 2 79 85 105 83 2 81 1 sky130_fd_sc_hd__and4bb_2 $T=143060 383520 1 0 $X=142870 $Y=380560
X3113 1 2 83 79 105 85 2 77 1 sky130_fd_sc_hd__and4bb_2 $T=146280 378080 0 0 $X=146090 $Y=377840
X3114 1 2 341 340 346 342 2 252 1 sky130_fd_sc_hd__and4bb_2 $T=517500 378080 0 0 $X=517310 $Y=377840
X3115 1 2 341 340 1505 342 2 347 1 sky130_fd_sc_hd__and4bb_2 $T=517960 388960 1 0 $X=517770 $Y=386000
X3116 1 2 342 341 1505 340 2 348 1 sky130_fd_sc_hd__and4bb_2 $T=518880 388960 0 0 $X=518690 $Y=388720
X3117 1 2 341 342 1505 340 2 350 1 sky130_fd_sc_hd__and4bb_2 $T=519340 394400 1 0 $X=519150 $Y=391440
X3118 1 2 98 94 361 96 2 346 1 sky130_fd_sc_hd__and4bb_2 $T=523940 378080 0 0 $X=523750 $Y=377840
X3119 1 2 341 342 1522 340 2 362 1 sky130_fd_sc_hd__and4bb_2 $T=526240 394400 1 0 $X=526050 $Y=391440
X3120 1 2 342 341 1522 340 2 364 1 sky130_fd_sc_hd__and4bb_2 $T=527160 388960 0 0 $X=526970 $Y=388720
X3121 1 2 341 340 1522 342 2 226 1 sky130_fd_sc_hd__and4bb_2 $T=527620 383520 0 0 $X=527430 $Y=383280
X3122 1 2 342 341 1530 340 2 285 1 sky130_fd_sc_hd__and4bb_2 $T=533600 394400 1 0 $X=533410 $Y=391440
X3123 1 2 341 342 1530 340 2 296 1 sky130_fd_sc_hd__and4bb_2 $T=534060 388960 1 0 $X=533870 $Y=386000
X3124 1 2 341 340 1530 342 2 253 1 sky130_fd_sc_hd__and4bb_2 $T=534060 399840 1 0 $X=533870 $Y=396880
X3125 1 2 341 340 375 342 2 380 1 sky130_fd_sc_hd__and4bb_2 $T=538660 383520 1 0 $X=538470 $Y=380560
X3126 1 2 341 342 375 340 2 223 1 sky130_fd_sc_hd__and4bb_2 $T=538660 388960 1 0 $X=538470 $Y=386000
X3127 1 2 361 2 1475 1 sky130_fd_sc_hd__clkbuf_4 $T=530840 394400 1 0 $X=530650 $Y=391440
X3128 2 1 1471 sky130_fd_sc_hd__conb_1 $T=522100 399840 1 0 $X=521910 $Y=396880
.ENDS
***************************************
.SUBCKT ICV_68 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=38
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=11500 0 0 0 $X=11310 $Y=-240
X1 1 2 6 7 8 3 4 5 ICV_13 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_69 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=26
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=7360 0 0 0 $X=7170 $Y=-240
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__dfxtp_1 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_70 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=10 FDC=36
*.SEEDPROM
X1 1 2 6 7 8 3 4 5 ICV_13 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_71 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=12 FDC=36
*.SEEDPROM
X1 1 2 6 7 8 3 4 5 ICV_13 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_72 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=24
*.SEEDPROM
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__dfxtp_1 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_73 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=10 FDC=24
*.SEEDPROM
X1 1 2 3 4 5 6 7 8 ICV_30 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_74 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=14 FDC=26
*.SEEDPROM
X0 1 2 3 4 2 5 1 sky130_fd_sc_hd__and2_1 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 8 6 2 7 1 sky130_fd_sc_hd__dlclkp_1 $T=2300 0 0 0 $X=2110 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_75 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380
+ 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400
+ 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420
+ 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440
+ 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460
+ 461 462 463 464 465 466 467 468 469 470
** N=2170 EP=470 IP=17032 FDC=47888
M0 1 3 518 1 nshort L=0.15 W=0.65 AD=0.08775 AS=0.182 PD=0.92 PS=1.86 NRD=0 NRS=0 m=1 r=4.33333 sa=75000.2 sb=75005.7 a=0.0975 p=1.6 mult=1 $X=121855 $Y=356555 $D=9
M1 6 4 1 1 nshort L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75000.6 sb=75005.3 a=0.0975 p=1.6 mult=1 $X=122275 $Y=356555 $D=9
M2 1 4 6 1 nshort L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75001 sb=75004.9 a=0.0975 p=1.6 mult=1 $X=122695 $Y=356555 $D=9
M3 6 4 1 1 nshort L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75001.5 sb=75004.5 a=0.0975 p=1.6 mult=1 $X=123115 $Y=356555 $D=9
M4 1 4 6 1 nshort L=0.15 W=0.65 AD=0.25675 AS=0.08775 PD=1.44 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75001.9 sb=75004.1 a=0.0975 p=1.6 mult=1 $X=123535 $Y=356555 $D=9
M5 6 5 1 1 nshort L=0.15 W=0.65 AD=0.08775 AS=0.25675 PD=0.92 PS=1.44 NRD=0 NRS=0 m=1 r=4.33333 sa=75002.8 sb=75003.1 a=0.0975 p=1.6 mult=1 $X=124475 $Y=356555 $D=9
M6 1 5 6 1 nshort L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75003.2 sb=75002.7 a=0.0975 p=1.6 mult=1 $X=124895 $Y=356555 $D=9
M7 6 5 1 1 nshort L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75003.7 sb=75002.3 a=0.0975 p=1.6 mult=1 $X=125315 $Y=356555 $D=9
M8 1 5 6 1 nshort L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75004.1 sb=75001.9 a=0.0975 p=1.6 mult=1 $X=125735 $Y=356555 $D=9
M9 6 518 1 1 nshort L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75004.5 sb=75001.4 a=0.0975 p=1.6 mult=1 $X=126155 $Y=356555 $D=9
M10 1 518 6 1 nshort L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75004.9 sb=75001 a=0.0975 p=1.6 mult=1 $X=126575 $Y=356555 $D=9
M11 6 518 1 1 nshort L=0.15 W=0.65 AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75005.3 sb=75000.6 a=0.0975 p=1.6 mult=1 $X=126995 $Y=356555 $D=9
M12 1 518 6 1 nshort L=0.15 W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 m=1 r=4.33333 sa=75005.8 sb=75000.2 a=0.0975 p=1.6 mult=1 $X=127415 $Y=356555 $D=9
M13 522 5 519 1 nshort L=0.15 W=0.65 AD=0.128375 AS=0.19825 PD=1.045 PS=1.91 NRD=26.304 NRS=0 m=1 r=4.33333 sa=75000.2 sb=75003 a=0.0975 p=1.6 mult=1 $X=527015 $Y=356555 $D=9
M14 523 4 522 1 nshort L=0.15 W=0.65 AD=0.06825 AS=0.128375 PD=0.86 PS=1.045 NRD=9.228 NRS=26.304 m=1 r=4.33333 sa=75000.8 sb=75002.4 a=0.0975 p=1.6 mult=1 $X=527560 $Y=356555 $D=8
M15 1 3 523 1 nshort L=0.15 W=0.65 AD=0.138125 AS=0.06825 PD=1.075 PS=0.86 NRD=18.456 NRS=9.228 m=1 r=4.33333 sa=75001.1 sb=75002.1 a=0.0975 p=1.6 mult=1 $X=527920 $Y=356555 $D=9
M16 7 519 1 1 nshort L=0.15 W=0.65 AD=0.091 AS=0.138125 PD=0.93 PS=1.075 NRD=0 NRS=8.304 m=1 r=4.33333 sa=75001.7 sb=75001.5 a=0.0975 p=1.6 mult=1 $X=528495 $Y=356555 $D=9
M17 1 519 7 1 nshort L=0.15 W=0.65 AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 m=1 r=4.33333 sa=75002.1 sb=75001.1 a=0.0975 p=1.6 mult=1 $X=528925 $Y=356555 $D=9
M18 7 519 1 1 nshort L=0.15 W=0.65 AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 m=1 r=4.33333 sa=75002.6 sb=75000.6 a=0.0975 p=1.6 mult=1 $X=529355 $Y=356555 $D=9
M19 1 519 7 1 nshort L=0.15 W=0.65 AD=0.18525 AS=0.091 PD=1.87 PS=0.93 NRD=0 NRS=0 m=1 r=4.33333 sa=75003 sb=75000.2 a=0.0975 p=1.6 mult=1 $X=529785 $Y=356555 $D=9
M20 2 3 518 2 phighvt L=0.15 W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 m=1 r=6.66667 sa=75000.2 sb=75001.9 a=0.15 p=2.3 mult=1 $X=121855 $Y=357805 $D=89
M21 520 4 2 2 phighvt L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75000.6 sb=75001.4 a=0.15 p=2.3 mult=1 $X=122275 $Y=357805 $D=89
M22 2 4 520 2 phighvt L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75001 sb=75001 a=0.15 p=2.3 mult=1 $X=122695 $Y=357805 $D=89
M23 520 4 2 2 phighvt L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75001.5 sb=75000.6 a=0.15 p=2.3 mult=1 $X=123115 $Y=357805 $D=89
M24 2 4 520 2 phighvt L=0.15 W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75001.9 sb=75000.2 a=0.15 p=2.3 mult=1 $X=123535 $Y=357805 $D=89
M25 520 5 521 2 phighvt L=0.15 W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 m=1 r=6.66667 sa=75000.2 sb=75003.1 a=0.15 p=2.3 mult=1 $X=124475 $Y=357805 $D=89
M26 521 5 520 2 phighvt L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75000.6 sb=75002.7 a=0.15 p=2.3 mult=1 $X=124895 $Y=357805 $D=89
M27 520 5 521 2 phighvt L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75001 sb=75002.3 a=0.15 p=2.3 mult=1 $X=125315 $Y=357805 $D=89
M28 521 5 520 2 phighvt L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75001.4 sb=75001.9 a=0.15 p=2.3 mult=1 $X=125735 $Y=357805 $D=89
M29 6 518 521 2 phighvt L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75001.9 sb=75001.4 a=0.15 p=2.3 mult=1 $X=126155 $Y=357805 $D=89
M30 521 518 6 2 phighvt L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75002.3 sb=75001 a=0.15 p=2.3 mult=1 $X=126575 $Y=357805 $D=89
M31 6 518 521 2 phighvt L=0.15 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75002.7 sb=75000.6 a=0.15 p=2.3 mult=1 $X=126995 $Y=357805 $D=89
M32 521 518 6 2 phighvt L=0.15 W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75003.1 sb=75000.2 a=0.15 p=2.3 mult=1 $X=127415 $Y=357805 $D=89
M33 2 5 519 2 phighvt L=0.15 W=1 AD=0.1975 AS=0.305 PD=1.395 PS=2.61 NRD=12.7853 NRS=0 m=1 r=6.66667 sa=75000.2 sb=75003 a=0.15 p=2.3 mult=1 $X=527015 $Y=357805 $D=89
M34 519 4 2 2 phighvt L=0.15 W=1 AD=0.14 AS=0.1975 PD=1.28 PS=1.395 NRD=0 NRS=9.8303 m=1 r=6.66667 sa=75000.8 sb=75002.4 a=0.15 p=2.3 mult=1 $X=527560 $Y=357805 $D=89
M35 2 3 519 2 phighvt L=0.15 W=1 AD=0.1775 AS=0.14 PD=1.355 PS=1.28 NRD=6.8753 NRS=0 m=1 r=6.66667 sa=75001.2 sb=75002 a=0.15 p=2.3 mult=1 $X=527990 $Y=357805 $D=89
M36 7 519 2 2 phighvt L=0.15 W=1 AD=0.14 AS=0.1775 PD=1.28 PS=1.355 NRD=0 NRS=7.8603 m=1 r=6.66667 sa=75001.7 sb=75001.5 a=0.15 p=2.3 mult=1 $X=528495 $Y=357805 $D=89
M37 2 519 7 2 phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75002.1 sb=75001.1 a=0.15 p=2.3 mult=1 $X=528925 $Y=357805 $D=89
M38 7 519 2 2 phighvt L=0.15 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75002.6 sb=75000.6 a=0.15 p=2.3 mult=1 $X=529355 $Y=357805 $D=89
M39 2 519 7 2 phighvt L=0.15 W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75003 sb=75000.2 a=0.15 p=2.3 mult=1 $X=529785 $Y=357805 $D=89
X40 1 2 Dpar a=2090.3 p=1485.74 m=1 $[nwdiode] $X=5330 $Y=314105 $D=191
X41 1 2 Dpar a=2091.12 p=1484.74 m=1 $[nwdiode] $X=5330 $Y=319545 $D=191
X42 1 2 Dpar a=2091.03 p=1484.84 m=1 $[nwdiode] $X=5330 $Y=324985 $D=191
X43 1 2 Dpar a=2090.3 p=1485.74 m=1 $[nwdiode] $X=5330 $Y=330425 $D=191
X44 1 2 Dpar a=2090.95 p=1484.94 m=1 $[nwdiode] $X=5330 $Y=335865 $D=191
X45 1 2 Dpar a=2090.95 p=1484.94 m=1 $[nwdiode] $X=5330 $Y=341305 $D=191
X46 1 2 Dpar a=2091.03 p=1484.84 m=1 $[nwdiode] $X=5330 $Y=346745 $D=191
X47 1 2 Dpar a=2090.79 p=1485.14 m=1 $[nwdiode] $X=5330 $Y=352185 $D=191
X48 1 2 Dpar a=2090.79 p=1485.14 m=1 $[nwdiode] $X=5330 $Y=357625 $D=191
X49 1 2 Dpar a=2090.14 p=1485.94 m=1 $[nwdiode] $X=5330 $Y=363065 $D=191
X50 1 2 Dpar a=2091.28 p=1484.54 m=1 $[nwdiode] $X=5330 $Y=368505 $D=191
X51 1 2 Dpar a=2090.95 p=1484.94 m=1 $[nwdiode] $X=5330 $Y=373945 $D=191
X52 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 312800 0 0 $X=5330 $Y=312560
X53 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 367200 1 0 $X=5330 $Y=364240
X54 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 378080 1 0 $X=5330 $Y=375120
X55 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=6900 312800 0 0 $X=6710 $Y=312560
X56 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=6900 329120 0 0 $X=6710 $Y=328880
X57 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=6900 361760 1 0 $X=6710 $Y=358800
X58 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=18400 334560 1 0 $X=18210 $Y=331600
X59 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=27600 361760 1 0 $X=27410 $Y=358800
X60 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=57960 350880 1 0 $X=57770 $Y=347920
X61 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=101660 367200 0 0 $X=101470 $Y=366960
X62 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=102580 372640 1 0 $X=102390 $Y=369680
X63 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=104420 350880 1 0 $X=104230 $Y=347920
X64 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=106260 329120 0 0 $X=106070 $Y=328880
X65 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=109940 345440 0 0 $X=109750 $Y=345200
X66 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=118220 361760 0 0 $X=118030 $Y=361520
X67 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=118220 378080 1 0 $X=118030 $Y=375120
X68 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=122360 372640 0 0 $X=122170 $Y=372400
X69 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=126500 372640 1 0 $X=126310 $Y=369680
X70 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=128800 361760 0 0 $X=128610 $Y=361520
X71 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=136620 372640 0 0 $X=136430 $Y=372400
X72 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=150420 356320 1 0 $X=150230 $Y=353360
X73 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=154560 378080 1 0 $X=154370 $Y=375120
X74 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=158700 329120 1 0 $X=158510 $Y=326160
X75 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=170660 345440 1 0 $X=170470 $Y=342480
X76 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=174340 356320 1 0 $X=174150 $Y=353360
X77 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=186760 372640 1 0 $X=186570 $Y=369680
X78 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=189060 334560 0 0 $X=188870 $Y=334320
X79 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=220800 340000 1 0 $X=220610 $Y=337040
X80 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=228620 329120 0 0 $X=228430 $Y=328880
X81 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=232300 356320 1 0 $X=232110 $Y=353360
X82 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=242880 361760 1 0 $X=242690 $Y=358800
X83 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=247020 318240 1 0 $X=246830 $Y=315280
X84 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=258520 340000 0 0 $X=258330 $Y=339760
X85 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=260820 323680 1 0 $X=260630 $Y=320720
X86 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=268640 372640 1 0 $X=268450 $Y=369680
X87 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=270940 323680 1 0 $X=270750 $Y=320720
X88 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=277380 312800 0 0 $X=277190 $Y=312560
X89 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=277840 350880 0 0 $X=277650 $Y=350640
X90 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=278300 318240 0 0 $X=278110 $Y=318000
X91 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=284280 372640 1 0 $X=284090 $Y=369680
X92 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=286580 334560 0 0 $X=286390 $Y=334320
X93 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=290720 372640 0 0 $X=290530 $Y=372400
X94 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=299000 318240 1 0 $X=298810 $Y=315280
X95 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=306360 356320 1 0 $X=306170 $Y=353360
X96 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=308660 334560 0 0 $X=308470 $Y=334320
X97 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=314640 356320 0 0 $X=314450 $Y=356080
X98 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=325680 334560 0 0 $X=325490 $Y=334320
X99 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=328900 378080 1 0 $X=328710 $Y=375120
X100 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=340860 372640 0 0 $X=340670 $Y=372400
X101 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=352820 350880 1 0 $X=352630 $Y=347920
X102 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=355120 329120 1 0 $X=354930 $Y=326160
X103 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=368920 312800 0 0 $X=368730 $Y=312560
X104 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=383180 356320 1 0 $X=382990 $Y=353360
X105 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=383180 367200 1 0 $X=382990 $Y=364240
X106 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=396980 367200 0 0 $X=396790 $Y=366960
X107 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=411240 345440 1 0 $X=411050 $Y=342480
X108 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=413540 367200 0 0 $X=413350 $Y=366960
X109 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=414920 312800 0 0 $X=414730 $Y=312560
X110 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=422280 334560 1 0 $X=422090 $Y=331600
X111 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=426880 345440 0 0 $X=426690 $Y=345200
X112 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=426880 361760 0 0 $X=426690 $Y=361520
X113 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=435160 329120 1 0 $X=434970 $Y=326160
X114 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=460920 372640 1 0 $X=460730 $Y=369680
X115 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=465060 350880 0 0 $X=464870 $Y=350640
X116 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=467360 318240 1 0 $X=467170 $Y=315280
X117 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=481160 350880 0 0 $X=480970 $Y=350640
X118 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=483000 367200 0 0 $X=482810 $Y=366960
X119 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=495420 345440 0 0 $X=495230 $Y=345200
X120 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=512440 312800 0 0 $X=512250 $Y=312560
X121 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=515660 334560 0 0 $X=515470 $Y=334320
X122 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=519340 361760 1 0 $X=519150 $Y=358800
X123 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=529000 372640 1 0 $X=528810 $Y=369680
X124 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=547860 367200 0 0 $X=547670 $Y=366960
X125 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=559360 372640 0 0 $X=559170 $Y=372400
X126 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=571320 350880 0 0 $X=571130 $Y=350640
X127 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=572240 356320 1 0 $X=572050 $Y=353360
X128 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=601220 361760 1 0 $X=601030 $Y=358800
X129 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=607660 372640 1 0 $X=607470 $Y=369680
X130 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=621460 334560 0 0 $X=621270 $Y=334320
X131 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=628820 323680 1 0 $X=628630 $Y=320720
X132 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=658720 329120 0 0 $X=658530 $Y=328880
X133 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=673440 334560 0 0 $X=673250 $Y=334320
X134 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=680340 345440 1 0 $X=680150 $Y=342480
X135 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=687700 367200 1 0 $X=687510 $Y=364240
X136 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=733700 323680 0 0 $X=733510 $Y=323440
X137 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=733700 329120 0 0 $X=733510 $Y=328880
X138 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=741520 323680 1 0 $X=741330 $Y=320720
X139 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 312800 1 180 $X=742710 $Y=312560
X140 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 378080 0 180 $X=742710 $Y=375120
X141 1 2 ICV_1 $T=5520 361760 1 0 $X=5330 $Y=358800
X142 1 2 ICV_1 $T=5520 372640 1 0 $X=5330 $Y=369680
X143 1 2 ICV_1 $T=744280 372640 0 180 $X=742710 $Y=369680
X144 1 2 ICV_2 $T=5520 318240 1 0 $X=5330 $Y=315280
X145 1 2 ICV_2 $T=5520 329120 1 0 $X=5330 $Y=326160
X146 1 2 ICV_2 $T=5520 340000 1 0 $X=5330 $Y=337040
X147 1 2 ICV_2 $T=5520 350880 1 0 $X=5330 $Y=347920
X148 1 2 ICV_2 $T=744280 318240 0 180 $X=742710 $Y=315280
X149 1 2 ICV_2 $T=744280 329120 0 180 $X=742710 $Y=326160
X150 1 2 ICV_2 $T=744280 340000 0 180 $X=742710 $Y=337040
X151 1 2 ICV_2 $T=744280 350880 0 180 $X=742710 $Y=347920
X152 1 2 ICV_2 $T=744280 361760 0 180 $X=742710 $Y=358800
X354 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=6900 350880 0 0 $X=6710 $Y=350640
X355 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=46000 367200 1 0 $X=45810 $Y=364240
X356 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=62100 323680 1 0 $X=61910 $Y=320720
X357 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=65780 334560 1 0 $X=65590 $Y=331600
X358 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=66240 350880 0 0 $X=66050 $Y=350640
X359 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=76360 361760 1 0 $X=76170 $Y=358800
X360 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=88320 356320 1 0 $X=88130 $Y=353360
X361 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=124660 350880 0 0 $X=124470 $Y=350640
X362 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=125120 378080 1 0 $X=124930 $Y=375120
X363 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=143520 323680 0 0 $X=143330 $Y=323440
X364 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=143520 367200 0 0 $X=143330 $Y=366960
X365 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=143520 372640 0 0 $X=143330 $Y=372400
X366 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=158240 323680 0 0 $X=158050 $Y=323440
X367 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=162380 312800 0 0 $X=162190 $Y=312560
X368 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=164680 323680 1 0 $X=164490 $Y=320720
X369 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=171580 367200 0 0 $X=171390 $Y=366960
X370 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=174340 345440 0 0 $X=174150 $Y=345200
X371 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=183540 361760 0 0 $X=183350 $Y=361520
X372 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=185840 323680 1 0 $X=185650 $Y=320720
X373 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=220340 329120 0 0 $X=220150 $Y=328880
X374 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=226780 318240 1 0 $X=226590 $Y=315280
X375 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=236900 318240 1 0 $X=236710 $Y=315280
X376 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=266340 350880 1 0 $X=266150 $Y=347920
X377 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=266800 345440 0 0 $X=266610 $Y=345200
X378 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=274160 350880 1 0 $X=273970 $Y=347920
X379 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=280600 329120 1 0 $X=280410 $Y=326160
X380 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=304980 372640 1 0 $X=304790 $Y=369680
X381 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=326140 356320 1 0 $X=325950 $Y=353360
X382 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=326600 372640 1 0 $X=326410 $Y=369680
X383 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=333040 318240 1 0 $X=332850 $Y=315280
X384 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=337180 329120 1 0 $X=336990 $Y=326160
X385 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=346840 356320 0 0 $X=346650 $Y=356080
X386 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=353740 340000 0 0 $X=353550 $Y=339760
X387 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=354200 323680 1 0 $X=354010 $Y=320720
X388 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=354200 372640 1 0 $X=354010 $Y=369680
X389 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=356960 323680 1 0 $X=356770 $Y=320720
X390 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=356960 372640 1 0 $X=356770 $Y=369680
X391 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=373520 323680 1 0 $X=373330 $Y=320720
X392 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=396520 312800 0 0 $X=396330 $Y=312560
X393 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=410320 350880 1 0 $X=410130 $Y=347920
X394 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=413080 323680 1 0 $X=412890 $Y=320720
X395 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=414920 378080 1 0 $X=414730 $Y=375120
X396 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=438840 323680 1 0 $X=438650 $Y=320720
X397 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=445280 378080 1 0 $X=445090 $Y=375120
X398 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=494960 378080 1 0 $X=494770 $Y=375120
X399 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=497260 367200 1 0 $X=497070 $Y=364240
X400 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=513820 367200 1 0 $X=513630 $Y=364240
X401 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=515200 367200 0 0 $X=515010 $Y=366960
X402 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=516580 350880 1 0 $X=516390 $Y=347920
X403 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=527160 350880 0 0 $X=526970 $Y=350640
X404 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=528540 340000 1 0 $X=528350 $Y=337040
X405 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=532220 318240 1 0 $X=532030 $Y=315280
X406 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=532680 356320 0 0 $X=532490 $Y=356080
X407 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=536360 312800 0 0 $X=536170 $Y=312560
X408 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=539120 312800 0 0 $X=538930 $Y=312560
X409 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=564420 350880 1 0 $X=564230 $Y=347920
X410 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=578680 323680 1 0 $X=578490 $Y=320720
X411 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=581440 329120 0 0 $X=581250 $Y=328880
X412 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=584200 334560 0 0 $X=584010 $Y=334320
X413 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=588800 329120 1 0 $X=588610 $Y=326160
X414 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=588800 367200 1 0 $X=588610 $Y=364240
X415 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=592480 334560 0 0 $X=592290 $Y=334320
X416 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=593400 318240 1 0 $X=593210 $Y=315280
X417 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=607200 378080 1 0 $X=607010 $Y=375120
X418 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=620540 361760 0 0 $X=620350 $Y=361520
X419 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=623300 361760 1 0 $X=623110 $Y=358800
X420 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=627900 350880 1 0 $X=627710 $Y=347920
X421 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=637560 345440 1 0 $X=637370 $Y=342480
X422 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=651360 318240 0 0 $X=651170 $Y=318000
X423 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=665620 334560 1 0 $X=665430 $Y=331600
X424 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=690920 361760 1 0 $X=690730 $Y=358800
X425 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=691380 372640 1 0 $X=691190 $Y=369680
X426 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=696440 312800 0 0 $X=696250 $Y=312560
X427 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=701040 329120 1 0 $X=700850 $Y=326160
X428 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=707480 345440 0 0 $X=707290 $Y=345200
X429 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=707940 361760 1 0 $X=707750 $Y=358800
X430 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=711620 361760 0 0 $X=711430 $Y=361520
X431 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=716220 318240 0 0 $X=716030 $Y=318000
X432 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=720360 356320 0 0 $X=720170 $Y=356080
X433 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=732780 318240 0 0 $X=732590 $Y=318000
X434 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=733240 367200 0 0 $X=733050 $Y=366960
X435 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 318240 0 0 $X=740870 $Y=318000
X436 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 350880 0 0 $X=740870 $Y=350640
X437 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 356320 0 0 $X=740870 $Y=356080
X438 1 2 ICV_3 $T=40020 372640 1 0 $X=39830 $Y=369680
X439 1 2 ICV_3 $T=69460 378080 1 0 $X=69270 $Y=375120
X440 1 2 ICV_3 $T=70840 340000 0 0 $X=70650 $Y=339760
X441 1 2 ICV_3 $T=101660 323680 0 0 $X=101470 $Y=323440
X442 1 2 ICV_3 $T=101660 378080 1 0 $X=101470 $Y=375120
X443 1 2 ICV_3 $T=102580 340000 0 0 $X=102390 $Y=339760
X444 1 2 ICV_3 $T=118220 318240 0 0 $X=118030 $Y=318000
X445 1 2 ICV_3 $T=143980 378080 1 0 $X=143790 $Y=375120
X446 1 2 ICV_3 $T=160540 334560 1 0 $X=160350 $Y=331600
X447 1 2 ICV_3 $T=160540 345440 1 0 $X=160350 $Y=342480
X448 1 2 ICV_3 $T=174340 372640 0 0 $X=174150 $Y=372400
X449 1 2 ICV_3 $T=192740 378080 1 0 $X=192550 $Y=375120
X450 1 2 ICV_3 $T=199640 345440 0 0 $X=199450 $Y=345200
X451 1 2 ICV_3 $T=213900 340000 1 0 $X=213710 $Y=337040
X452 1 2 ICV_3 $T=231380 361760 1 0 $X=231190 $Y=358800
X453 1 2 ICV_3 $T=239660 312800 0 0 $X=239470 $Y=312560
X454 1 2 ICV_3 $T=243800 361760 0 0 $X=243610 $Y=361520
X455 1 2 ICV_3 $T=266800 312800 0 0 $X=266610 $Y=312560
X456 1 2 ICV_3 $T=270020 323680 0 0 $X=269830 $Y=323440
X457 1 2 ICV_3 $T=276920 323680 1 0 $X=276730 $Y=320720
X458 1 2 ICV_3 $T=297620 312800 0 0 $X=297430 $Y=312560
X459 1 2 ICV_3 $T=298080 356320 0 0 $X=297890 $Y=356080
X460 1 2 ICV_3 $T=322000 378080 1 0 $X=321810 $Y=375120
X461 1 2 ICV_3 $T=326140 318240 1 0 $X=325950 $Y=315280
X462 1 2 ICV_3 $T=345460 323680 1 0 $X=345270 $Y=320720
X463 1 2 ICV_3 $T=354200 361760 0 0 $X=354010 $Y=361520
X464 1 2 ICV_3 $T=382260 378080 1 0 $X=382070 $Y=375120
X465 1 2 ICV_3 $T=383180 323680 0 0 $X=382990 $Y=323440
X466 1 2 ICV_3 $T=391460 378080 1 0 $X=391270 $Y=375120
X467 1 2 ICV_3 $T=411700 334560 0 0 $X=411510 $Y=334320
X468 1 2 ICV_3 $T=438380 356320 1 0 $X=438190 $Y=353360
X469 1 2 ICV_3 $T=442520 372640 0 0 $X=442330 $Y=372400
X470 1 2 ICV_3 $T=469200 334560 1 0 $X=469010 $Y=331600
X471 1 2 ICV_3 $T=480240 340000 0 0 $X=480050 $Y=339760
X472 1 2 ICV_3 $T=517500 372640 1 0 $X=517310 $Y=369680
X473 1 2 ICV_3 $T=547400 312800 0 0 $X=547210 $Y=312560
X474 1 2 ICV_3 $T=564420 318240 0 0 $X=564230 $Y=318000
X475 1 2 ICV_3 $T=564420 329120 0 0 $X=564230 $Y=328880
X476 1 2 ICV_3 $T=568100 378080 1 0 $X=567910 $Y=375120
X477 1 2 ICV_3 $T=571780 340000 1 0 $X=571590 $Y=337040
X478 1 2 ICV_3 $T=574540 329120 1 0 $X=574350 $Y=326160
X479 1 2 ICV_3 $T=595240 356320 0 0 $X=595050 $Y=356080
X480 1 2 ICV_3 $T=615940 329120 1 0 $X=615750 $Y=326160
X481 1 2 ICV_3 $T=637560 367200 1 0 $X=637370 $Y=364240
X482 1 2 ICV_3 $T=649060 350880 1 0 $X=648870 $Y=347920
X483 1 2 ICV_3 $T=652280 361760 1 0 $X=652090 $Y=358800
X484 1 2 ICV_3 $T=659180 345440 0 0 $X=658990 $Y=345200
X485 1 2 ICV_3 $T=665620 372640 1 0 $X=665430 $Y=369680
X486 1 2 ICV_3 $T=679420 334560 0 0 $X=679230 $Y=334320
X487 1 2 ICV_3 $T=683100 329120 1 0 $X=682910 $Y=326160
X488 1 2 ICV_3 $T=697360 323680 0 0 $X=697170 $Y=323440
X489 1 2 ICV_3 $T=698280 329120 0 0 $X=698090 $Y=328880
X490 1 2 ICV_3 $T=740600 318240 1 0 $X=740410 $Y=315280
X491 1 2 ICV_3 $T=740600 340000 1 0 $X=740410 $Y=337040
X492 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=14260 367200 0 0 $X=14070 $Y=366960
X493 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=20240 372640 1 0 $X=20050 $Y=369680
X494 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=28520 345440 1 0 $X=28330 $Y=342480
X495 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=41400 312800 0 0 $X=41210 $Y=312560
X496 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=45080 378080 1 0 $X=44890 $Y=375120
X497 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=57040 345440 1 0 $X=56850 $Y=342480
X498 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=76360 356320 1 0 $X=76170 $Y=353360
X499 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=89240 345440 1 0 $X=89050 $Y=342480
X500 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=90160 334560 0 0 $X=89970 $Y=334320
X501 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=90160 345440 0 0 $X=89970 $Y=345200
X502 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=120980 334560 1 0 $X=120790 $Y=331600
X503 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=120980 367200 1 0 $X=120790 $Y=364240
X504 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=130180 312800 0 0 $X=129990 $Y=312560
X505 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=132480 334560 1 0 $X=132290 $Y=331600
X506 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=132480 334560 0 0 $X=132290 $Y=334320
X507 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=136160 367200 0 0 $X=135970 $Y=366960
X508 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=136620 378080 1 0 $X=136430 $Y=375120
X509 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=138920 329120 0 0 $X=138730 $Y=328880
X510 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=139840 350880 1 0 $X=139650 $Y=347920
X511 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=143060 345440 0 0 $X=142870 $Y=345200
X512 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=150420 345440 0 0 $X=150230 $Y=345200
X513 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=157320 340000 1 0 $X=157130 $Y=337040
X514 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=161000 345440 0 0 $X=160810 $Y=345200
X515 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=174340 356320 0 0 $X=174150 $Y=356080
X516 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=188600 323680 1 0 $X=188410 $Y=320720
X517 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=189520 318240 0 0 $X=189330 $Y=318000
X518 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=189980 350880 0 0 $X=189790 $Y=350640
X519 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=199180 323680 0 0 $X=198990 $Y=323440
X520 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=199180 340000 0 0 $X=198990 $Y=339760
X521 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=213440 334560 1 0 $X=213250 $Y=331600
X522 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=213440 345440 1 0 $X=213250 $Y=342480
X523 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=216660 329120 1 0 $X=216470 $Y=326160
X524 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=218500 345440 0 0 $X=218310 $Y=345200
X525 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=220800 345440 1 0 $X=220610 $Y=342480
X526 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=234600 340000 0 0 $X=234410 $Y=339760
X527 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=237820 329120 0 0 $X=237630 $Y=328880
X528 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=237820 367200 0 0 $X=237630 $Y=366960
X529 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=242420 356320 0 0 $X=242230 $Y=356080
X530 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=248860 350880 1 0 $X=248670 $Y=347920
X531 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=255300 356320 0 0 $X=255110 $Y=356080
X532 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=259900 329120 1 0 $X=259710 $Y=326160
X533 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=281060 361760 1 0 $X=280870 $Y=358800
X534 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=286580 340000 0 0 $X=286390 $Y=339760
X535 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=290720 312800 0 0 $X=290530 $Y=312560
X536 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=300840 345440 1 0 $X=300650 $Y=342480
X537 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=314640 329120 0 0 $X=314450 $Y=328880
X538 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=314640 367200 0 0 $X=314450 $Y=366960
X539 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=314640 372640 0 0 $X=314450 $Y=372400
X540 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=322920 323680 0 0 $X=322730 $Y=323440
X541 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=342700 318240 0 0 $X=342510 $Y=318000
X542 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=353740 356320 1 0 $X=353550 $Y=353360
X543 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=370760 372640 0 0 $X=370570 $Y=372400
X544 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=396520 340000 1 0 $X=396330 $Y=337040
X545 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=409860 367200 1 0 $X=409670 $Y=364240
X546 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=413080 350880 1 0 $X=412890 $Y=347920
X547 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=415840 318240 0 0 $X=415650 $Y=318000
X548 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=419520 323680 0 0 $X=419330 $Y=323440
X549 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=426880 318240 0 0 $X=426690 $Y=318000
X550 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=426880 323680 0 0 $X=426690 $Y=323440
X551 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=434240 334560 0 0 $X=434050 $Y=334320
X552 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=445280 356320 1 0 $X=445090 $Y=353360
X553 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=454940 350880 0 0 $X=454750 $Y=350640
X554 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=467360 318240 0 0 $X=467170 $Y=318000
X555 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=469200 345440 1 0 $X=469010 $Y=342480
X556 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=485300 372640 1 0 $X=485110 $Y=369680
X557 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=489440 361760 0 0 $X=489250 $Y=361520
X558 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=500480 329120 0 0 $X=500290 $Y=328880
X559 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=514280 323680 1 0 $X=514090 $Y=320720
X560 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=551080 334560 0 0 $X=550890 $Y=334320
X561 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=563960 340000 0 0 $X=563770 $Y=339760
X562 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=574540 323680 0 0 $X=574350 $Y=323440
X563 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=581440 345440 1 0 $X=581250 $Y=342480
X564 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=592020 367200 0 0 $X=591830 $Y=366960
X565 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=602140 329120 1 0 $X=601950 $Y=326160
X566 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=609500 323680 1 0 $X=609310 $Y=320720
X567 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=609500 367200 1 0 $X=609310 $Y=364240
X568 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=640780 361760 0 0 $X=640590 $Y=361520
X569 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=642160 361760 1 0 $X=641970 $Y=358800
X570 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=662400 345440 1 0 $X=662210 $Y=342480
X571 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=690460 323680 1 0 $X=690270 $Y=320720
X572 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=690920 318240 0 0 $X=690730 $Y=318000
X573 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=695520 345440 0 0 $X=695330 $Y=345200
X574 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=721740 340000 0 0 $X=721550 $Y=339760
X575 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=722200 334560 0 0 $X=722010 $Y=334320
X576 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=732320 312800 0 0 $X=732130 $Y=312560
X577 1 2 ICV_4 $T=19780 361760 0 0 $X=19590 $Y=361520
X578 1 2 ICV_4 $T=80040 361760 0 0 $X=79850 $Y=361520
X579 1 2 ICV_4 $T=86480 372640 0 0 $X=86290 $Y=372400
X580 1 2 ICV_4 $T=100740 323680 1 0 $X=100550 $Y=320720
X581 1 2 ICV_4 $T=118220 367200 0 0 $X=118030 $Y=366960
X582 1 2 ICV_4 $T=136160 372640 1 0 $X=135970 $Y=369680
X583 1 2 ICV_4 $T=143980 372640 1 0 $X=143790 $Y=369680
X584 1 2 ICV_4 $T=161460 356320 0 0 $X=161270 $Y=356080
X585 1 2 ICV_4 $T=174340 361760 0 0 $X=174150 $Y=361520
X586 1 2 ICV_4 $T=180780 318240 1 0 $X=180590 $Y=315280
X587 1 2 ICV_4 $T=180780 350880 0 0 $X=180590 $Y=350640
X588 1 2 ICV_4 $T=182620 329120 0 0 $X=182430 $Y=328880
X589 1 2 ICV_4 $T=183080 356320 0 0 $X=182890 $Y=356080
X590 1 2 ICV_4 $T=210680 356320 0 0 $X=210490 $Y=356080
X591 1 2 ICV_4 $T=211140 312800 0 0 $X=210950 $Y=312560
X592 1 2 ICV_4 $T=226780 372640 0 0 $X=226590 $Y=372400
X593 1 2 ICV_4 $T=227700 329120 1 0 $X=227510 $Y=326160
X594 1 2 ICV_4 $T=234600 372640 0 0 $X=234410 $Y=372400
X595 1 2 ICV_4 $T=264960 345440 1 0 $X=264770 $Y=342480
X596 1 2 ICV_4 $T=304980 350880 0 0 $X=304790 $Y=350640
X597 1 2 ICV_4 $T=325220 340000 1 0 $X=325030 $Y=337040
X598 1 2 ICV_4 $T=405260 323680 1 0 $X=405070 $Y=320720
X599 1 2 ICV_4 $T=429180 340000 0 0 $X=428990 $Y=339760
X600 1 2 ICV_4 $T=473800 361760 0 0 $X=473610 $Y=361520
X601 1 2 ICV_4 $T=493580 350880 1 0 $X=493390 $Y=347920
X602 1 2 ICV_4 $T=523020 372640 0 0 $X=522830 $Y=372400
X603 1 2 ICV_4 $T=535440 367200 1 0 $X=535250 $Y=364240
X604 1 2 ICV_4 $T=539120 334560 1 0 $X=538930 $Y=331600
X605 1 2 ICV_4 $T=563040 323680 1 0 $X=562850 $Y=320720
X606 1 2 ICV_4 $T=602600 340000 0 0 $X=602410 $Y=339760
X607 1 2 ICV_4 $T=608120 372640 0 0 $X=607930 $Y=372400
X608 1 2 ICV_4 $T=611340 318240 0 0 $X=611150 $Y=318000
X609 1 2 ICV_4 $T=629740 312800 0 0 $X=629550 $Y=312560
X610 1 2 ICV_4 $T=637560 378080 1 0 $X=637370 $Y=375120
X611 1 2 ICV_4 $T=699660 340000 0 0 $X=699470 $Y=339760
X612 1 2 ICV_4 $T=731860 340000 0 0 $X=731670 $Y=339760
X613 1 2 ICV_4 $T=731860 345440 0 0 $X=731670 $Y=345200
X614 1 2 ICV_4 $T=731860 372640 0 0 $X=731670 $Y=372400
X615 1 2 ICV_4 $T=739680 312800 0 0 $X=739490 $Y=312560
X616 1 2 ICV_4 $T=739680 323680 0 0 $X=739490 $Y=323440
X617 1 2 ICV_4 $T=739680 329120 0 0 $X=739490 $Y=328880
X618 1 2 ICV_4 $T=739680 334560 0 0 $X=739490 $Y=334320
X619 1 2 ICV_4 $T=739680 340000 0 0 $X=739490 $Y=339760
X620 1 2 ICV_4 $T=739680 345440 0 0 $X=739490 $Y=345200
X621 1 2 ICV_4 $T=739680 361760 0 0 $X=739490 $Y=361520
X622 1 2 ICV_4 $T=739680 367200 0 0 $X=739490 $Y=366960
X623 1 2 ICV_4 $T=739680 372640 0 0 $X=739490 $Y=372400
X624 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 334560 1 0 $X=6710 $Y=331600
X625 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 356320 1 0 $X=6710 $Y=353360
X626 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=16100 345440 1 0 $X=15910 $Y=342480
X627 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=16100 378080 1 0 $X=15910 $Y=375120
X628 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=23920 340000 0 0 $X=23730 $Y=339760
X629 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=27600 367200 1 0 $X=27410 $Y=364240
X630 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=29900 329120 0 0 $X=29710 $Y=328880
X631 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=35880 334560 1 0 $X=35690 $Y=331600
X632 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=45540 329120 0 0 $X=45350 $Y=328880
X633 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=55660 334560 1 0 $X=55470 $Y=331600
X634 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=79120 312800 0 0 $X=78930 $Y=312560
X635 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=90160 361760 0 0 $X=89970 $Y=361520
X636 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=100280 350880 1 0 $X=100090 $Y=347920
X637 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=113160 318240 0 0 $X=112970 $Y=318000
X638 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=114080 329120 0 0 $X=113890 $Y=328880
X639 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=114080 334560 0 0 $X=113890 $Y=334320
X640 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=120980 340000 1 0 $X=120790 $Y=337040
X641 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=130640 350880 0 0 $X=130450 $Y=350640
X642 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=146280 334560 0 0 $X=146090 $Y=334320
X643 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=156400 318240 1 0 $X=156210 $Y=315280
X644 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=174340 329120 1 0 $X=174150 $Y=326160
X645 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=174340 334560 1 0 $X=174150 $Y=331600
X646 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=175260 340000 1 0 $X=175070 $Y=337040
X647 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=188600 350880 1 0 $X=188410 $Y=347920
X648 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=202400 367200 1 0 $X=202210 $Y=364240
X649 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=218960 340000 0 0 $X=218770 $Y=339760
X650 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=225400 356320 0 0 $X=225210 $Y=356080
X651 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=226320 367200 0 0 $X=226130 $Y=366960
X652 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=240120 356320 1 0 $X=239930 $Y=353360
X653 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=248860 340000 1 0 $X=248670 $Y=337040
X654 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=257600 361760 1 0 $X=257410 $Y=358800
X655 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=258520 367200 0 0 $X=258330 $Y=366960
X656 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=272780 318240 1 0 $X=272590 $Y=315280
X657 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=280140 367200 1 0 $X=279950 $Y=364240
X658 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=282440 356320 0 0 $X=282250 $Y=356080
X659 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=286580 367200 0 0 $X=286390 $Y=366960
X660 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=310500 323680 0 0 $X=310310 $Y=323440
X661 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=313720 329120 1 0 $X=313530 $Y=326160
X662 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=314640 334560 0 0 $X=314450 $Y=334320
X663 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=324760 329120 1 0 $X=324570 $Y=326160
X664 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=337640 334560 1 0 $X=337450 $Y=331600
X665 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=356960 378080 1 0 $X=356770 $Y=375120
X666 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=359720 350880 0 0 $X=359530 $Y=350640
X667 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=369840 378080 1 0 $X=369650 $Y=375120
X668 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=371680 367200 1 0 $X=371490 $Y=364240
X669 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=373520 345440 1 0 $X=373330 $Y=342480
X670 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=393300 367200 0 0 $X=393110 $Y=366960
X671 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=422280 361760 0 0 $X=422090 $Y=361520
X672 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=441140 350880 1 0 $X=440950 $Y=347920
X673 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=450340 340000 0 0 $X=450150 $Y=339760
X674 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=451260 367200 1 0 $X=451070 $Y=364240
X675 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=462760 361760 0 0 $X=462570 $Y=361520
X676 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=474260 345440 0 0 $X=474070 $Y=345200
X677 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=496340 318240 0 0 $X=496150 $Y=318000
X678 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=525320 361760 1 0 $X=525130 $Y=358800
X679 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=525320 378080 1 0 $X=525130 $Y=375120
X680 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=530380 345440 0 0 $X=530190 $Y=345200
X681 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=530840 323680 0 0 $X=530650 $Y=323440
X682 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=535900 372640 1 0 $X=535710 $Y=369680
X683 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=536820 356320 1 0 $X=536630 $Y=353360
X684 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=539120 340000 0 0 $X=538930 $Y=339760
X685 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=562120 312800 0 0 $X=561930 $Y=312560
X686 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=562120 372640 1 0 $X=561930 $Y=369680
X687 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=589720 356320 0 0 $X=589530 $Y=356080
X688 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=591100 345440 0 0 $X=590910 $Y=345200
X689 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=605360 367200 1 0 $X=605170 $Y=364240
X690 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=606740 345440 0 0 $X=606550 $Y=345200
X691 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=609500 350880 1 0 $X=609310 $Y=347920
X692 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=623300 318240 0 0 $X=623110 $Y=318000
X693 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=632500 345440 0 0 $X=632310 $Y=345200
X694 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=639860 356320 0 0 $X=639670 $Y=356080
X695 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=644920 345440 1 0 $X=644730 $Y=342480
X696 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=647220 350880 0 0 $X=647030 $Y=350640
X697 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=649980 356320 1 0 $X=649790 $Y=353360
X698 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=660560 323680 1 0 $X=660370 $Y=320720
X699 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=661480 329120 1 0 $X=661290 $Y=326160
X700 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=669760 345440 1 0 $X=669570 $Y=342480
X701 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=675280 345440 0 0 $X=675090 $Y=345200
X702 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=675280 361760 0 0 $X=675090 $Y=361520
X703 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=679880 378080 1 0 $X=679690 $Y=375120
X704 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=683560 356320 0 0 $X=683370 $Y=356080
X705 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=689540 329120 1 0 $X=689350 $Y=326160
X706 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=695980 356320 0 0 $X=695790 $Y=356080
X707 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=707020 372640 1 0 $X=706830 $Y=369680
X708 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=707480 318240 1 0 $X=707290 $Y=315280
X709 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=717600 378080 1 0 $X=717410 $Y=375120
X710 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=720820 345440 0 0 $X=720630 $Y=345200
X711 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=737840 323680 1 0 $X=737650 $Y=320720
X712 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=738300 356320 1 0 $X=738110 $Y=353360
X713 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=738760 361760 1 0 $X=738570 $Y=358800
X714 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 323680 0 0 $X=6710 $Y=323440
X715 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 372640 0 0 $X=6710 $Y=372400
X716 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=48760 356320 0 0 $X=48570 $Y=356080
X717 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=107180 361760 0 0 $X=106990 $Y=361520
X718 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=107640 372640 0 0 $X=107450 $Y=372400
X719 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=236900 356320 0 0 $X=236710 $Y=356080
X720 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=247020 367200 0 0 $X=246830 $Y=366960
X721 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=266800 367200 1 0 $X=266610 $Y=364240
X722 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=280140 312800 0 0 $X=279950 $Y=312560
X723 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=300840 356320 1 0 $X=300650 $Y=353360
X724 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=322000 361760 1 0 $X=321810 $Y=358800
X725 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=416760 361760 0 0 $X=416570 $Y=361520
X726 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=430560 318240 1 0 $X=430370 $Y=315280
X727 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=445280 323680 1 0 $X=445090 $Y=320720
X728 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=463220 323680 1 0 $X=463030 $Y=320720
X729 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=516580 334560 1 0 $X=516390 $Y=331600
X730 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=590180 372640 1 0 $X=589990 $Y=369680
X731 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=631580 378080 1 0 $X=631390 $Y=375120
X732 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=633880 350880 0 0 $X=633690 $Y=350640
X733 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=647220 323680 1 0 $X=647030 $Y=320720
X734 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=679420 312800 0 0 $X=679230 $Y=312560
X735 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=733240 361760 1 0 $X=733050 $Y=358800
X736 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 318240 0 0 $X=735350 $Y=318000
X737 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 350880 0 0 $X=735350 $Y=350640
X738 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 356320 0 0 $X=735350 $Y=356080
X739 1 2 8 2 24 1 sky130_fd_sc_hd__clkbuf_8 $T=6900 345440 0 0 $X=6710 $Y=345200
X740 1 2 159 2 165 1 sky130_fd_sc_hd__clkbuf_8 $T=160540 318240 1 0 $X=160350 $Y=315280
X741 1 2 543 533 2 39 1 sky130_fd_sc_hd__ebufn_2 $T=14720 361760 1 0 $X=14530 $Y=358800
X742 1 2 567 548 2 52 1 sky130_fd_sc_hd__ebufn_2 $T=27600 340000 0 0 $X=27410 $Y=339760
X743 1 2 572 51 2 37 1 sky130_fd_sc_hd__ebufn_2 $T=29440 312800 0 0 $X=29250 $Y=312560
X744 1 2 606 72 2 36 1 sky130_fd_sc_hd__ebufn_2 $T=50140 323680 1 0 $X=49950 $Y=320720
X745 1 2 618 72 2 34 1 sky130_fd_sc_hd__ebufn_2 $T=56580 323680 0 0 $X=56390 $Y=323440
X746 1 2 613 609 2 33 1 sky130_fd_sc_hd__ebufn_2 $T=57500 367200 0 0 $X=57310 $Y=366960
X747 1 2 636 609 2 59 1 sky130_fd_sc_hd__ebufn_2 $T=63020 367200 1 0 $X=62830 $Y=364240
X748 1 2 655 645 2 37 1 sky130_fd_sc_hd__ebufn_2 $T=73140 340000 0 0 $X=72950 $Y=339760
X749 1 2 662 664 2 54 1 sky130_fd_sc_hd__ebufn_2 $T=75900 361760 0 0 $X=75710 $Y=361520
X750 1 2 667 653 2 54 1 sky130_fd_sc_hd__ebufn_2 $T=77280 329120 1 0 $X=77090 $Y=326160
X751 1 2 666 90 2 33 1 sky130_fd_sc_hd__ebufn_2 $T=83260 361760 0 0 $X=83070 $Y=361520
X752 1 2 709 690 2 28 1 sky130_fd_sc_hd__ebufn_2 $T=98440 340000 0 0 $X=98250 $Y=339760
X753 1 2 712 713 2 28 1 sky130_fd_sc_hd__ebufn_2 $T=99820 334560 1 0 $X=99630 $Y=331600
X754 1 2 714 100 2 55 1 sky130_fd_sc_hd__ebufn_2 $T=103040 361760 0 0 $X=102850 $Y=361520
X755 1 2 721 699 2 36 1 sky130_fd_sc_hd__ebufn_2 $T=103960 323680 0 0 $X=103770 $Y=323440
X756 1 2 733 713 2 36 1 sky130_fd_sc_hd__ebufn_2 $T=113160 340000 0 0 $X=112970 $Y=339760
X757 1 2 754 759 2 28 1 sky130_fd_sc_hd__ebufn_2 $T=126500 350880 0 0 $X=126310 $Y=350640
X758 1 2 740 747 2 39 1 sky130_fd_sc_hd__ebufn_2 $T=126960 318240 0 0 $X=126770 $Y=318000
X759 1 2 139 126 2 34 1 sky130_fd_sc_hd__ebufn_2 $T=141220 312800 0 0 $X=141030 $Y=312560
X760 1 2 792 791 2 54 1 sky130_fd_sc_hd__ebufn_2 $T=148120 318240 0 0 $X=147930 $Y=318000
X761 1 2 796 783 2 37 1 sky130_fd_sc_hd__ebufn_2 $T=149960 334560 0 0 $X=149770 $Y=334320
X762 1 2 794 791 2 28 1 sky130_fd_sc_hd__ebufn_2 $T=154100 323680 1 0 $X=153910 $Y=320720
X763 1 2 803 741 2 52 1 sky130_fd_sc_hd__ebufn_2 $T=168360 350880 0 0 $X=168170 $Y=350640
X764 1 2 823 821 2 180 1 sky130_fd_sc_hd__ebufn_2 $T=169280 361760 0 0 $X=169090 $Y=361520
X765 1 2 802 741 2 34 1 sky130_fd_sc_hd__ebufn_2 $T=178020 350880 1 0 $X=177830 $Y=347920
X766 1 2 206 205 2 176 1 sky130_fd_sc_hd__ebufn_2 $T=195040 378080 1 0 $X=194850 $Y=375120
X767 1 2 873 852 2 186 1 sky130_fd_sc_hd__ebufn_2 $T=200560 345440 1 0 $X=200370 $Y=342480
X768 1 2 861 854 2 197 1 sky130_fd_sc_hd__ebufn_2 $T=203780 318240 1 0 $X=203590 $Y=315280
X769 1 2 210 205 2 180 1 sky130_fd_sc_hd__ebufn_2 $T=210680 378080 1 0 $X=210490 $Y=375120
X770 1 2 216 217 2 179 1 sky130_fd_sc_hd__ebufn_2 $T=218960 334560 0 0 $X=218770 $Y=334320
X771 1 2 941 911 2 179 1 sky130_fd_sc_hd__ebufn_2 $T=239200 329120 1 0 $X=239010 $Y=326160
X772 1 2 983 987 2 198 1 sky130_fd_sc_hd__ebufn_2 $T=259900 350880 1 0 $X=259710 $Y=347920
X773 1 2 1019 1004 2 199 1 sky130_fd_sc_hd__ebufn_2 $T=276000 350880 1 0 $X=275810 $Y=347920
X774 1 2 1044 239 2 167 1 sky130_fd_sc_hd__ebufn_2 $T=290260 367200 0 0 $X=290070 $Y=366960
X775 1 2 1053 245 2 179 1 sky130_fd_sc_hd__ebufn_2 $T=293480 312800 0 0 $X=293290 $Y=312560
X776 1 2 1055 1039 2 179 1 sky130_fd_sc_hd__ebufn_2 $T=293940 350880 1 0 $X=293750 $Y=347920
X777 1 2 1075 1076 2 198 1 sky130_fd_sc_hd__ebufn_2 $T=303600 345440 1 0 $X=303410 $Y=342480
X778 1 2 1090 254 2 201 1 sky130_fd_sc_hd__ebufn_2 $T=313720 323680 1 0 $X=313530 $Y=320720
X779 1 2 1091 1094 2 167 1 sky130_fd_sc_hd__ebufn_2 $T=317860 361760 1 0 $X=317670 $Y=358800
X780 1 2 282 284 2 268 1 sky130_fd_sc_hd__ebufn_2 $T=339020 378080 1 0 $X=338830 $Y=375120
X781 1 2 1130 1138 2 275 1 sky130_fd_sc_hd__ebufn_2 $T=341320 323680 1 0 $X=341130 $Y=320720
X782 1 2 1149 1120 2 263 1 sky130_fd_sc_hd__ebufn_2 $T=344080 350880 0 0 $X=343890 $Y=350640
X783 1 2 1151 1138 2 268 1 sky130_fd_sc_hd__ebufn_2 $T=345460 318240 0 0 $X=345270 $Y=318000
X784 1 2 1155 1158 2 263 1 sky130_fd_sc_hd__ebufn_2 $T=348680 356320 0 0 $X=348490 $Y=356080
X785 1 2 1175 1158 2 280 1 sky130_fd_sc_hd__ebufn_2 $T=358800 372640 1 0 $X=358610 $Y=369680
X786 1 2 1194 1173 2 280 1 sky130_fd_sc_hd__ebufn_2 $T=371680 345440 0 0 $X=371490 $Y=345200
X787 1 2 318 289 2 277 1 sky130_fd_sc_hd__ebufn_2 $T=379040 323680 0 0 $X=378850 $Y=323440
X788 1 2 1207 315 2 263 1 sky130_fd_sc_hd__ebufn_2 $T=379500 318240 1 0 $X=379310 $Y=315280
X789 1 2 1211 319 2 280 1 sky130_fd_sc_hd__ebufn_2 $T=380420 367200 0 0 $X=380230 $Y=366960
X790 1 2 1212 1223 2 275 1 sky130_fd_sc_hd__ebufn_2 $T=385480 323680 0 0 $X=385290 $Y=323440
X791 1 2 1259 1261 2 268 1 sky130_fd_sc_hd__ebufn_2 $T=403880 345440 0 0 $X=403690 $Y=345200
X792 1 2 1272 328 2 296 1 sky130_fd_sc_hd__ebufn_2 $T=421360 318240 1 0 $X=421170 $Y=315280
X793 1 2 1292 1261 2 269 1 sky130_fd_sc_hd__ebufn_2 $T=421820 345440 0 0 $X=421630 $Y=345200
X794 1 2 1300 1295 2 280 1 sky130_fd_sc_hd__ebufn_2 $T=426420 318240 1 0 $X=426230 $Y=315280
X795 1 2 357 358 2 277 1 sky130_fd_sc_hd__ebufn_2 $T=447120 378080 1 0 $X=446930 $Y=375120
X796 1 2 1363 1350 2 269 1 sky130_fd_sc_hd__ebufn_2 $T=459080 323680 1 0 $X=458890 $Y=320720
X797 1 2 1380 1356 2 280 1 sky130_fd_sc_hd__ebufn_2 $T=464140 356320 1 0 $X=463950 $Y=353360
X798 1 2 1387 1356 2 277 1 sky130_fd_sc_hd__ebufn_2 $T=470120 345440 0 0 $X=469930 $Y=345200
X799 1 2 1401 1382 2 263 1 sky130_fd_sc_hd__ebufn_2 $T=474720 318240 0 0 $X=474530 $Y=318000
X800 1 2 1405 1391 2 275 1 sky130_fd_sc_hd__ebufn_2 $T=477020 361760 0 0 $X=476830 $Y=361520
X801 1 2 372 370 2 296 1 sky130_fd_sc_hd__ebufn_2 $T=477480 372640 0 0 $X=477290 $Y=372400
X802 1 2 1402 371 2 275 1 sky130_fd_sc_hd__ebufn_2 $T=477940 312800 0 0 $X=477750 $Y=312560
X803 1 2 1437 1450 2 280 1 sky130_fd_sc_hd__ebufn_2 $T=495880 334560 0 0 $X=495690 $Y=334320
X804 1 2 1481 1425 2 275 1 sky130_fd_sc_hd__ebufn_2 $T=512900 323680 0 0 $X=512710 $Y=323440
X805 1 2 1470 1450 2 263 1 sky130_fd_sc_hd__ebufn_2 $T=512900 340000 1 0 $X=512710 $Y=337040
X806 1 2 1474 1434 2 263 1 sky130_fd_sc_hd__ebufn_2 $T=513360 372640 1 0 $X=513170 $Y=369680
X807 1 2 1487 1456 2 263 1 sky130_fd_sc_hd__ebufn_2 $T=517040 356320 1 0 $X=516850 $Y=353360
X808 1 2 1502 1506 2 407 1 sky130_fd_sc_hd__ebufn_2 $T=526240 334560 1 0 $X=526050 $Y=331600
X809 1 2 1547 1543 2 422 1 sky130_fd_sc_hd__ebufn_2 $T=551080 340000 0 0 $X=550890 $Y=339760
X810 1 2 1535 1507 2 418 1 sky130_fd_sc_hd__ebufn_2 $T=557980 312800 0 0 $X=557790 $Y=312560
X811 1 2 1573 1543 2 409 1 sky130_fd_sc_hd__ebufn_2 $T=567640 340000 1 0 $X=567450 $Y=337040
X812 1 2 1579 426 2 418 1 sky130_fd_sc_hd__ebufn_2 $T=570400 378080 1 0 $X=570210 $Y=375120
X813 1 2 1597 1580 2 424 1 sky130_fd_sc_hd__ebufn_2 $T=576840 329120 1 0 $X=576650 $Y=326160
X814 1 2 1615 1604 2 424 1 sky130_fd_sc_hd__ebufn_2 $T=585580 356320 0 0 $X=585390 $Y=356080
X815 1 2 1623 437 2 424 1 sky130_fd_sc_hd__ebufn_2 $T=589720 378080 1 0 $X=589530 $Y=375120
X816 1 2 1619 1604 2 418 1 sky130_fd_sc_hd__ebufn_2 $T=590640 361760 0 0 $X=590450 $Y=361520
X817 1 2 1639 1604 2 405 1 sky130_fd_sc_hd__ebufn_2 $T=597540 356320 0 0 $X=597350 $Y=356080
X818 1 2 1670 1668 2 407 1 sky130_fd_sc_hd__ebufn_2 $T=612260 367200 1 0 $X=612070 $Y=364240
X819 1 2 1723 1694 2 424 1 sky130_fd_sc_hd__ebufn_2 $T=639860 367200 1 0 $X=639670 $Y=364240
X820 1 2 1725 1722 2 409 1 sky130_fd_sc_hd__ebufn_2 $T=640780 345440 1 0 $X=640590 $Y=342480
X821 1 2 1737 1722 2 408 1 sky130_fd_sc_hd__ebufn_2 $T=645840 356320 1 0 $X=645650 $Y=353360
X822 1 2 1738 1719 2 424 1 sky130_fd_sc_hd__ebufn_2 $T=646760 323680 0 0 $X=646570 $Y=323440
X823 1 2 1751 453 2 418 1 sky130_fd_sc_hd__ebufn_2 $T=654580 361760 1 0 $X=654390 $Y=358800
X824 1 2 1772 455 2 418 1 sky130_fd_sc_hd__ebufn_2 $T=667920 372640 1 0 $X=667730 $Y=369680
X825 1 2 1785 1749 2 405 1 sky130_fd_sc_hd__ebufn_2 $T=672520 312800 0 0 $X=672330 $Y=312560
X826 1 2 1803 1781 2 407 1 sky130_fd_sc_hd__ebufn_2 $T=678960 329120 1 0 $X=678770 $Y=326160
X827 1 2 1813 1781 2 409 1 sky130_fd_sc_hd__ebufn_2 $T=685400 329120 1 0 $X=685210 $Y=326160
X828 1 2 1838 1818 2 409 1 sky130_fd_sc_hd__ebufn_2 $T=699660 356320 0 0 $X=699470 $Y=356080
X829 1 2 1844 462 2 407 1 sky130_fd_sc_hd__ebufn_2 $T=700120 372640 0 0 $X=699930 $Y=372400
X830 1 2 1835 456 2 405 1 sky130_fd_sc_hd__ebufn_2 $T=701960 318240 0 0 $X=701770 $Y=318000
X831 1 2 1872 1881 2 407 1 sky130_fd_sc_hd__ebufn_2 $T=717140 367200 1 0 $X=716950 $Y=364240
X832 1 2 1896 1869 2 408 1 sky130_fd_sc_hd__ebufn_2 $T=733700 323680 1 0 $X=733510 $Y=320720
X833 1 2 1900 1871 2 418 1 sky130_fd_sc_hd__ebufn_2 $T=734160 356320 1 0 $X=733970 $Y=353360
X834 1 2 1912 469 2 418 1 sky130_fd_sc_hd__ebufn_2 $T=736460 318240 1 0 $X=736270 $Y=315280
X835 1 2 1910 1889 2 417 1 sky130_fd_sc_hd__ebufn_2 $T=736460 340000 1 0 $X=736270 $Y=337040
X836 1 2 1918 468 2 418 1 sky130_fd_sc_hd__ebufn_2 $T=738760 367200 1 0 $X=738570 $Y=364240
X951 1 2 544 548 39 ICV_6 $T=19780 334560 1 0 $X=19590 $Y=331600
X952 1 2 601 590 54 ICV_6 $T=47840 361760 1 0 $X=47650 $Y=358800
X953 1 2 631 80 39 ICV_6 $T=61640 312800 0 0 $X=61450 $Y=312560
X954 1 2 619 596 39 ICV_6 $T=61640 340000 0 0 $X=61450 $Y=339760
X955 1 2 621 624 34 ICV_6 $T=61640 350880 0 0 $X=61450 $Y=350640
X956 1 2 630 624 52 ICV_6 $T=61640 361760 0 0 $X=61450 $Y=361520
X957 1 2 654 653 36 ICV_6 $T=75900 334560 1 0 $X=75710 $Y=331600
X958 1 2 665 645 34 ICV_6 $T=75900 340000 1 0 $X=75710 $Y=337040
X959 1 2 660 645 54 ICV_6 $T=75900 345440 1 0 $X=75710 $Y=342480
X960 1 2 658 664 37 ICV_6 $T=75900 350880 1 0 $X=75710 $Y=347920
X961 1 2 675 90 38 ICV_6 $T=89700 367200 0 0 $X=89510 $Y=366960
X962 1 2 684 90 75 ICV_6 $T=89700 372640 0 0 $X=89510 $Y=372400
X963 1 2 723 699 34 ICV_6 $T=103960 323680 1 0 $X=103770 $Y=320720
X964 1 2 719 100 33 ICV_6 $T=103960 372640 1 0 $X=103770 $Y=369680
X965 1 2 715 100 49 ICV_6 $T=103960 378080 1 0 $X=103770 $Y=375120
X966 1 2 767 747 57 ICV_6 $T=132020 323680 1 0 $X=131830 $Y=320720
X967 1 2 762 701 52 ICV_6 $T=132020 345440 1 0 $X=131830 $Y=342480
X968 1 2 784 701 37 ICV_6 $T=145820 345440 0 0 $X=145630 $Y=345200
X969 1 2 810 791 39 ICV_6 $T=160080 323680 1 0 $X=159890 $Y=320720
X970 1 2 809 791 37 ICV_6 $T=160080 329120 1 0 $X=159890 $Y=326160
X971 1 2 799 783 36 ICV_6 $T=160080 340000 1 0 $X=159890 $Y=337040
X972 1 2 846 820 199 ICV_6 $T=188140 334560 1 0 $X=187950 $Y=331600
X973 1 2 848 820 201 ICV_6 $T=188140 340000 1 0 $X=187950 $Y=337040
X974 1 2 202 203 185 ICV_6 $T=188140 378080 1 0 $X=187950 $Y=375120
X975 1 2 865 854 201 ICV_6 $T=201940 323680 0 0 $X=201750 $Y=323440
X976 1 2 866 852 197 ICV_6 $T=201940 334560 0 0 $X=201750 $Y=334320
X977 1 2 877 852 184 ICV_6 $T=201940 340000 0 0 $X=201750 $Y=339760
X978 1 2 872 852 199 ICV_6 $T=201940 345440 0 0 $X=201750 $Y=345200
X979 1 2 876 852 179 ICV_6 $T=201940 350880 0 0 $X=201750 $Y=350640
X980 1 2 880 868 174 ICV_6 $T=201940 361760 0 0 $X=201750 $Y=361520
X981 1 2 881 868 193 ICV_6 $T=201940 367200 0 0 $X=201750 $Y=366960
X982 1 2 901 888 184 ICV_6 $T=216200 340000 1 0 $X=216010 $Y=337040
X983 1 2 894 888 199 ICV_6 $T=216200 345440 1 0 $X=216010 $Y=342480
X984 1 2 900 888 179 ICV_6 $T=216200 350880 1 0 $X=216010 $Y=347920
X985 1 2 933 922 166 ICV_6 $T=230000 334560 0 0 $X=229810 $Y=334320
X986 1 2 927 922 184 ICV_6 $T=230000 340000 0 0 $X=229810 $Y=339760
X987 1 2 934 922 179 ICV_6 $T=230000 356320 0 0 $X=229810 $Y=356080
X988 1 2 920 924 193 ICV_6 $T=230000 372640 0 0 $X=229810 $Y=372400
X989 1 2 957 961 184 ICV_6 $T=244260 340000 1 0 $X=244070 $Y=337040
X990 1 2 960 961 201 ICV_6 $T=244260 350880 1 0 $X=244070 $Y=347920
X991 1 2 985 958 186 ICV_6 $T=258060 323680 0 0 $X=257870 $Y=323440
X992 1 2 981 958 199 ICV_6 $T=258060 329120 0 0 $X=257870 $Y=328880
X993 1 2 1005 1010 184 ICV_6 $T=272320 323680 1 0 $X=272130 $Y=320720
X994 1 2 1036 238 186 ICV_6 $T=286120 312800 0 0 $X=285930 $Y=312560
X995 1 2 1037 239 180 ICV_6 $T=286120 361760 0 0 $X=285930 $Y=361520
X996 1 2 246 243 194 ICV_6 $T=286120 372640 0 0 $X=285930 $Y=372400
X997 1 2 1067 1047 199 ICV_6 $T=300380 329120 1 0 $X=300190 $Y=326160
X998 1 2 1068 1021 185 ICV_6 $T=300380 372640 1 0 $X=300190 $Y=369680
X999 1 2 1096 254 197 ICV_6 $T=314180 312800 0 0 $X=313990 $Y=312560
X1000 1 2 270 254 179 ICV_6 $T=328440 318240 1 0 $X=328250 $Y=315280
X1001 1 2 1110 1083 201 ICV_6 $T=328440 340000 1 0 $X=328250 $Y=337040
X1002 1 2 1117 1094 185 ICV_6 $T=328440 372640 1 0 $X=328250 $Y=369680
X1003 1 2 1125 1131 277 ICV_6 $T=342240 356320 0 0 $X=342050 $Y=356080
X1004 1 2 1140 1094 176 ICV_6 $T=342240 372640 0 0 $X=342050 $Y=372400
X1005 1 2 1167 1138 296 ICV_6 $T=356500 329120 1 0 $X=356310 $Y=326160
X1006 1 2 1189 1186 268 ICV_6 $T=370300 329120 0 0 $X=370110 $Y=328880
X1007 1 2 1183 1186 269 ICV_6 $T=370300 334560 0 0 $X=370110 $Y=334320
X1008 1 2 1218 315 267 ICV_6 $T=384560 318240 1 0 $X=384370 $Y=315280
X1009 1 2 1213 1223 269 ICV_6 $T=384560 334560 1 0 $X=384370 $Y=331600
X1010 1 2 1216 1188 268 ICV_6 $T=384560 350880 1 0 $X=384370 $Y=347920
X1011 1 2 1221 1188 269 ICV_6 $T=384560 361760 1 0 $X=384370 $Y=358800
X1012 1 2 1210 319 263 ICV_6 $T=384560 367200 1 0 $X=384370 $Y=364240
X1013 1 2 323 319 269 ICV_6 $T=384560 378080 1 0 $X=384370 $Y=375120
X1014 1 2 1239 328 275 ICV_6 $T=398360 312800 0 0 $X=398170 $Y=312560
X1015 1 2 1245 1225 269 ICV_6 $T=398360 345440 0 0 $X=398170 $Y=345200
X1016 1 2 1247 1227 268 ICV_6 $T=398360 361760 0 0 $X=398170 $Y=361520
X1017 1 2 1274 1227 263 ICV_6 $T=412620 361760 1 0 $X=412430 $Y=358800
X1018 1 2 1276 1227 269 ICV_6 $T=412620 367200 1 0 $X=412430 $Y=364240
X1019 1 2 1297 349 267 ICV_6 $T=426420 312800 0 0 $X=426230 $Y=312560
X1020 1 2 1304 1295 263 ICV_6 $T=426420 329120 0 0 $X=426230 $Y=328880
X1021 1 2 1296 1261 277 ICV_6 $T=426420 350880 0 0 $X=426230 $Y=350640
X1022 1 2 1299 1306 269 ICV_6 $T=426420 372640 0 0 $X=426230 $Y=372400
X1023 1 2 1327 1295 268 ICV_6 $T=440680 323680 1 0 $X=440490 $Y=320720
X1024 1 2 1326 1308 267 ICV_6 $T=440680 356320 1 0 $X=440490 $Y=353360
X1025 1 2 1332 1306 267 ICV_6 $T=440680 378080 1 0 $X=440490 $Y=375120
X1026 1 2 1344 1350 296 ICV_6 $T=454480 334560 0 0 $X=454290 $Y=334320
X1027 1 2 1414 1382 277 ICV_6 $T=482540 323680 0 0 $X=482350 $Y=323440
X1028 1 2 1412 1371 280 ICV_6 $T=482540 334560 0 0 $X=482350 $Y=334320
X1029 1 2 1415 1400 263 ICV_6 $T=482540 340000 0 0 $X=482350 $Y=339760
X1030 1 2 1383 1356 263 ICV_6 $T=482540 345440 0 0 $X=482350 $Y=345200
X1031 1 2 1406 1400 268 ICV_6 $T=482540 350880 0 0 $X=482350 $Y=350640
X1032 1 2 1395 1391 268 ICV_6 $T=482540 372640 0 0 $X=482350 $Y=372400
X1033 1 2 1449 381 269 ICV_6 $T=496800 318240 1 0 $X=496610 $Y=315280
X1034 1 2 1447 1450 267 ICV_6 $T=496800 334560 1 0 $X=496610 $Y=331600
X1035 1 2 1441 1457 267 ICV_6 $T=496800 345440 1 0 $X=496610 $Y=342480
X1036 1 2 1451 1456 296 ICV_6 $T=496800 350880 1 0 $X=496610 $Y=347920
X1037 1 2 1448 1434 267 ICV_6 $T=496800 372640 1 0 $X=496610 $Y=369680
X1038 1 2 1440 382 269 ICV_6 $T=496800 378080 1 0 $X=496610 $Y=375120
X1039 1 2 1476 1457 268 ICV_6 $T=510600 340000 0 0 $X=510410 $Y=339760
X1040 1 2 1433 1457 269 ICV_6 $T=510600 345440 0 0 $X=510410 $Y=345200
X1041 1 2 1477 1434 268 ICV_6 $T=510600 367200 0 0 $X=510410 $Y=366960
X1042 1 2 1519 1506 424 ICV_6 $T=538660 329120 0 0 $X=538470 $Y=328880
X1043 1 2 1518 1506 417 ICV_6 $T=538660 334560 0 0 $X=538470 $Y=334320
X1044 1 2 1523 1503 422 ICV_6 $T=538660 345440 0 0 $X=538470 $Y=345200
X1045 1 2 1571 430 409 ICV_6 $T=566720 312800 0 0 $X=566530 $Y=312560
X1046 1 2 1562 1542 409 ICV_6 $T=566720 318240 0 0 $X=566530 $Y=318000
X1047 1 2 1568 1542 417 ICV_6 $T=566720 329120 0 0 $X=566530 $Y=328880
X1048 1 2 1576 1557 417 ICV_6 $T=566720 350880 0 0 $X=566530 $Y=350640
X1049 1 2 1600 1599 407 ICV_6 $T=580980 318240 1 0 $X=580790 $Y=315280
X1050 1 2 1627 1599 418 ICV_6 $T=594780 312800 0 0 $X=594590 $Y=312560
X1051 1 2 1628 1599 405 ICV_6 $T=594780 318240 0 0 $X=594590 $Y=318000
X1052 1 2 1630 1599 409 ICV_6 $T=594780 323680 0 0 $X=594590 $Y=323440
X1053 1 2 1643 1616 418 ICV_6 $T=609040 361760 1 0 $X=608850 $Y=358800
X1054 1 2 1685 1678 405 ICV_6 $T=622840 334560 0 0 $X=622650 $Y=334320
X1055 1 2 1687 1668 405 ICV_6 $T=622840 367200 0 0 $X=622650 $Y=366960
X1056 1 2 452 445 417 ICV_6 $T=650900 312800 0 0 $X=650710 $Y=312560
X1057 1 2 1773 1740 417 ICV_6 $T=665160 345440 1 0 $X=664970 $Y=342480
X1058 1 2 1804 1780 422 ICV_6 $T=678960 356320 0 0 $X=678770 $Y=356080
X1059 1 2 1800 455 422 ICV_6 $T=678960 367200 0 0 $X=678770 $Y=366960
X1060 1 2 1816 1797 405 ICV_6 $T=693220 340000 1 0 $X=693030 $Y=337040
X1061 1 2 1826 462 418 ICV_6 $T=707020 361760 0 0 $X=706830 $Y=361520
X1062 1 2 1870 468 407 ICV_6 $T=721280 367200 1 0 $X=721090 $Y=364240
X1063 1 2 1908 469 408 ICV_6 $T=735080 312800 0 0 $X=734890 $Y=312560
X1064 1 2 1897 1869 417 ICV_6 $T=735080 323680 0 0 $X=734890 $Y=323440
X1065 1 2 1876 1889 409 ICV_6 $T=735080 329120 0 0 $X=734890 $Y=328880
X1066 1 2 1885 1889 407 ICV_6 $T=735080 334560 0 0 $X=734890 $Y=334320
X1067 1 2 1903 1891 418 ICV_6 $T=735080 340000 0 0 $X=734890 $Y=339760
X1068 1 2 1905 1891 424 ICV_6 $T=735080 345440 0 0 $X=734890 $Y=345200
X1069 1 2 1914 1881 417 ICV_6 $T=735080 361760 0 0 $X=734890 $Y=361520
X1070 1 2 1915 1881 424 ICV_6 $T=735080 367200 0 0 $X=734890 $Y=366960
X1071 1 2 1907 468 424 ICV_6 $T=735080 372640 0 0 $X=734890 $Y=372400
X1194 1 2 ICV_10 $T=73140 329120 1 0 $X=72950 $Y=326160
X1195 1 2 ICV_10 $T=129260 361760 1 0 $X=129070 $Y=358800
X1196 1 2 ICV_10 $T=143060 334560 0 0 $X=142870 $Y=334320
X1197 1 2 ICV_10 $T=255300 318240 0 0 $X=255110 $Y=318000
X1198 1 2 ICV_10 $T=269560 361760 1 0 $X=269370 $Y=358800
X1199 1 2 ICV_10 $T=283360 345440 0 0 $X=283170 $Y=345200
X1200 1 2 ICV_10 $T=311420 372640 0 0 $X=311230 $Y=372400
X1201 1 2 ICV_10 $T=395600 372640 0 0 $X=395410 $Y=372400
X1202 1 2 ICV_10 $T=465980 340000 1 0 $X=465790 $Y=337040
X1203 1 2 ICV_10 $T=465980 361760 1 0 $X=465790 $Y=358800
X1204 1 2 ICV_10 $T=522100 334560 1 0 $X=521910 $Y=331600
X1205 1 2 ICV_10 $T=522100 378080 1 0 $X=521910 $Y=375120
X1206 1 2 ICV_10 $T=563960 356320 0 0 $X=563770 $Y=356080
X1207 1 2 ICV_10 $T=563960 367200 0 0 $X=563770 $Y=366960
X1208 1 2 ICV_10 $T=620080 345440 0 0 $X=619890 $Y=345200
X1209 1 2 ICV_10 $T=718520 340000 1 0 $X=718330 $Y=337040
X1210 1 2 526 25 2 532 1 sky130_fd_sc_hd__dfxtp_1 $T=17940 350880 0 0 $X=17750 $Y=350640
X1211 1 2 9 45 2 554 1 sky130_fd_sc_hd__dfxtp_1 $T=20240 367200 1 0 $X=20050 $Y=364240
X1212 1 2 531 15 2 583 1 sky130_fd_sc_hd__dfxtp_1 $T=34040 323680 0 0 $X=33850 $Y=323440
X1213 1 2 580 18 2 612 1 sky130_fd_sc_hd__dfxtp_1 $T=48300 334560 1 0 $X=48110 $Y=331600
X1214 1 2 591 13 2 618 1 sky130_fd_sc_hd__dfxtp_1 $T=49680 318240 0 0 $X=49490 $Y=318000
X1215 1 2 66 15 2 631 1 sky130_fd_sc_hd__dfxtp_1 $T=54280 312800 0 0 $X=54090 $Y=312560
X1216 1 2 627 44 2 642 1 sky130_fd_sc_hd__dfxtp_1 $T=59800 345440 1 0 $X=59610 $Y=342480
X1217 1 2 627 43 2 643 1 sky130_fd_sc_hd__dfxtp_1 $T=60260 340000 1 0 $X=60070 $Y=337040
X1218 1 2 83 70 2 684 1 sky130_fd_sc_hd__dfxtp_1 $T=79120 372640 0 0 $X=78930 $Y=372400
X1219 1 2 687 44 2 697 1 sky130_fd_sc_hd__dfxtp_1 $T=87860 329120 1 0 $X=87670 $Y=326160
X1220 1 2 672 15 2 708 1 sky130_fd_sc_hd__dfxtp_1 $T=92920 334560 0 0 $X=92730 $Y=334320
X1221 1 2 98 40 2 714 1 sky130_fd_sc_hd__dfxtp_1 $T=94300 367200 0 0 $X=94110 $Y=366960
X1222 1 2 94 13 2 104 1 sky130_fd_sc_hd__dfxtp_1 $T=100280 312800 0 0 $X=100090 $Y=312560
X1223 1 2 732 15 2 740 1 sky130_fd_sc_hd__dfxtp_1 $T=110400 323680 0 0 $X=110210 $Y=323440
X1224 1 2 732 42 2 746 1 sky130_fd_sc_hd__dfxtp_1 $T=112700 329120 1 0 $X=112510 $Y=326160
X1225 1 2 750 42 2 763 1 sky130_fd_sc_hd__dfxtp_1 $T=123740 334560 1 0 $X=123550 $Y=331600
X1226 1 2 772 42 2 792 1 sky130_fd_sc_hd__dfxtp_1 $T=141220 318240 1 0 $X=141030 $Y=315280
X1227 1 2 785 14 2 795 1 sky130_fd_sc_hd__dfxtp_1 $T=142600 350880 1 0 $X=142410 $Y=347920
X1228 1 2 786 18 2 796 1 sky130_fd_sc_hd__dfxtp_1 $T=144440 334560 1 0 $X=144250 $Y=331600
X1229 1 2 786 14 2 799 1 sky130_fd_sc_hd__dfxtp_1 $T=145820 345440 1 0 $X=145630 $Y=342480
X1230 1 2 800 161 2 827 1 sky130_fd_sc_hd__dfxtp_1 $T=160540 367200 1 0 $X=160350 $Y=364240
X1231 1 2 825 172 2 834 1 sky130_fd_sc_hd__dfxtp_1 $T=166980 329120 1 0 $X=166790 $Y=326160
X1232 1 2 800 181 2 839 1 sky130_fd_sc_hd__dfxtp_1 $T=177100 372640 1 0 $X=176910 $Y=369680
X1233 1 2 826 189 2 846 1 sky130_fd_sc_hd__dfxtp_1 $T=178020 334560 1 0 $X=177830 $Y=331600
X1234 1 2 855 190 2 874 1 sky130_fd_sc_hd__dfxtp_1 $T=192280 356320 1 0 $X=192090 $Y=353360
X1235 1 2 882 187 2 890 1 sky130_fd_sc_hd__dfxtp_1 $T=205160 329120 0 0 $X=204970 $Y=328880
X1236 1 2 913 189 2 925 1 sky130_fd_sc_hd__dfxtp_1 $T=221260 345440 0 0 $X=221070 $Y=345200
X1237 1 2 913 187 2 921 1 sky130_fd_sc_hd__dfxtp_1 $T=222640 340000 0 0 $X=222450 $Y=339760
X1238 1 2 914 172 2 936 1 sky130_fd_sc_hd__dfxtp_1 $T=225400 334560 1 0 $X=225210 $Y=331600
X1239 1 2 939 170 2 954 1 sky130_fd_sc_hd__dfxtp_1 $T=236900 340000 1 0 $X=236710 $Y=337040
X1240 1 2 939 168 2 957 1 sky130_fd_sc_hd__dfxtp_1 $T=237360 340000 0 0 $X=237170 $Y=339760
X1241 1 2 950 189 2 981 1 sky130_fd_sc_hd__dfxtp_1 $T=250700 329120 0 0 $X=250510 $Y=328880
X1242 1 2 968 189 2 984 1 sky130_fd_sc_hd__dfxtp_1 $T=251620 350880 1 0 $X=251430 $Y=347920
X1243 1 2 968 168 2 986 1 sky130_fd_sc_hd__dfxtp_1 $T=252540 340000 1 0 $X=252350 $Y=337040
X1244 1 2 968 190 2 989 1 sky130_fd_sc_hd__dfxtp_1 $T=253460 356320 1 0 $X=253270 $Y=353360
X1245 1 2 992 168 2 1005 1 sky130_fd_sc_hd__dfxtp_1 $T=262660 323680 0 0 $X=262470 $Y=323440
X1246 1 2 1008 175 2 1020 1 sky130_fd_sc_hd__dfxtp_1 $T=270020 361760 0 0 $X=269830 $Y=361520
X1247 1 2 995 171 2 1003 1 sky130_fd_sc_hd__dfxtp_1 $T=270480 350880 0 0 $X=270290 $Y=350640
X1248 1 2 233 172 2 1036 1 sky130_fd_sc_hd__dfxtp_1 $T=276460 318240 1 0 $X=276270 $Y=315280
X1249 1 2 1022 177 2 1018 1 sky130_fd_sc_hd__dfxtp_1 $T=278760 372640 0 0 $X=278570 $Y=372400
X1250 1 2 1030 187 2 1059 1 sky130_fd_sc_hd__dfxtp_1 $T=289340 340000 0 0 $X=289150 $Y=339760
X1251 1 2 1073 171 2 1107 1 sky130_fd_sc_hd__dfxtp_1 $T=317400 329120 1 0 $X=317210 $Y=326160
X1252 1 2 1061 187 2 1104 1 sky130_fd_sc_hd__dfxtp_1 $T=317860 340000 1 0 $X=317670 $Y=337040
X1253 1 2 1073 168 2 1111 1 sky130_fd_sc_hd__dfxtp_1 $T=318320 334560 0 0 $X=318130 $Y=334320
X1254 1 2 1095 264 2 274 1 sky130_fd_sc_hd__dfxtp_1 $T=325220 372640 0 0 $X=325030 $Y=372400
X1255 1 2 278 253 2 1156 1 sky130_fd_sc_hd__dfxtp_1 $T=342700 312800 0 0 $X=342510 $Y=312560
X1256 1 2 1102 257 2 1154 1 sky130_fd_sc_hd__dfxtp_1 $T=342700 345440 0 0 $X=342510 $Y=345200
X1257 1 2 1171 264 2 1191 1 sky130_fd_sc_hd__dfxtp_1 $T=362940 334560 0 0 $X=362750 $Y=334320
X1258 1 2 165 188 2 311 1 sky130_fd_sc_hd__dfxtp_1 $T=364320 356320 1 0 $X=364130 $Y=353360
X1259 1 2 1169 253 2 1198 1 sky130_fd_sc_hd__dfxtp_1 $T=366160 345440 1 0 $X=365970 $Y=342480
X1260 1 2 1187 264 2 1185 1 sky130_fd_sc_hd__dfxtp_1 $T=370760 356320 0 0 $X=370570 $Y=356080
X1261 1 2 312 253 2 1210 1 sky130_fd_sc_hd__dfxtp_1 $T=373520 372640 0 0 $X=373330 $Y=372400
X1262 1 2 1203 262 2 1213 1 sky130_fd_sc_hd__dfxtp_1 $T=377200 334560 1 0 $X=377010 $Y=331600
X1263 1 2 1230 262 2 1276 1 sky130_fd_sc_hd__dfxtp_1 $T=406180 367200 0 0 $X=405990 $Y=366960
X1264 1 2 1257 264 2 1285 1 sky130_fd_sc_hd__dfxtp_1 $T=412620 356320 0 0 $X=412430 $Y=356080
X1265 1 2 1294 273 2 1323 1 sky130_fd_sc_hd__dfxtp_1 $T=430100 361760 1 0 $X=429910 $Y=358800
X1266 1 2 1294 260 2 1326 1 sky130_fd_sc_hd__dfxtp_1 $T=431020 350880 0 0 $X=430830 $Y=350640
X1267 1 2 343 264 2 1329 1 sky130_fd_sc_hd__dfxtp_1 $T=431940 372640 1 0 $X=431750 $Y=369680
X1268 1 2 343 253 2 1324 1 sky130_fd_sc_hd__dfxtp_1 $T=434240 367200 0 0 $X=434050 $Y=366960
X1269 1 2 1301 273 2 1337 1 sky130_fd_sc_hd__dfxtp_1 $T=438380 340000 0 0 $X=438190 $Y=339760
X1270 1 2 1339 260 2 1361 1 sky130_fd_sc_hd__dfxtp_1 $T=448040 356320 1 0 $X=447850 $Y=353360
X1271 1 2 1334 273 2 1362 1 sky130_fd_sc_hd__dfxtp_1 $T=454940 372640 0 0 $X=454750 $Y=372400
X1272 1 2 1339 273 2 1380 1 sky130_fd_sc_hd__dfxtp_1 $T=457700 350880 0 0 $X=457510 $Y=350640
X1273 1 2 1385 260 2 1399 1 sky130_fd_sc_hd__dfxtp_1 $T=466440 361760 0 0 $X=466250 $Y=361520
X1274 1 2 1384 273 2 1426 1 sky130_fd_sc_hd__dfxtp_1 $T=480700 356320 1 0 $X=480510 $Y=353360
X1275 1 2 365 264 2 1422 1 sky130_fd_sc_hd__dfxtp_1 $T=483000 312800 0 0 $X=482810 $Y=312560
X1276 1 2 1413 262 2 1433 1 sky130_fd_sc_hd__dfxtp_1 $T=486220 350880 1 0 $X=486030 $Y=347920
X1277 1 2 1413 273 2 1436 1 sky130_fd_sc_hd__dfxtp_1 $T=487140 340000 0 0 $X=486950 $Y=339760
X1278 1 2 378 262 2 1449 1 sky130_fd_sc_hd__dfxtp_1 $T=489440 318240 1 0 $X=489250 $Y=315280
X1279 1 2 1413 265 2 1471 1 sky130_fd_sc_hd__dfxtp_1 $T=503240 345440 0 0 $X=503050 $Y=345200
X1280 1 2 1428 266 2 1475 1 sky130_fd_sc_hd__dfxtp_1 $T=504620 340000 1 0 $X=504430 $Y=337040
X1281 1 2 1485 400 2 1502 1 sky130_fd_sc_hd__dfxtp_1 $T=519340 334560 0 0 $X=519150 $Y=334320
X1282 1 2 1496 400 2 1515 1 sky130_fd_sc_hd__dfxtp_1 $T=529000 361760 1 0 $X=528810 $Y=358800
X1283 1 2 1486 414 2 1523 1 sky130_fd_sc_hd__dfxtp_1 $T=531760 345440 1 0 $X=531570 $Y=342480
X1284 1 2 1527 400 2 1544 1 sky130_fd_sc_hd__dfxtp_1 $T=542800 340000 0 0 $X=542610 $Y=339760
X1285 1 2 1529 414 2 1549 1 sky130_fd_sc_hd__dfxtp_1 $T=545560 329120 0 0 $X=545370 $Y=328880
X1286 1 2 427 398 2 1572 1 sky130_fd_sc_hd__dfxtp_1 $T=557060 318240 0 0 $X=556870 $Y=318000
X1287 1 2 431 410 2 432 1 sky130_fd_sc_hd__dfxtp_1 $T=560740 378080 1 0 $X=560550 $Y=375120
X1288 1 2 1578 400 2 1600 1 sky130_fd_sc_hd__dfxtp_1 $T=571320 318240 0 0 $X=571130 $Y=318000
X1289 1 2 1612 400 2 1614 1 sky130_fd_sc_hd__dfxtp_1 $T=584200 345440 1 0 $X=584010 $Y=342480
X1290 1 2 1578 398 2 1628 1 sky130_fd_sc_hd__dfxtp_1 $T=586500 312800 0 0 $X=586310 $Y=312560
X1291 1 2 1618 415 2 1645 1 sky130_fd_sc_hd__dfxtp_1 $T=595240 340000 0 0 $X=595050 $Y=339760
X1292 1 2 1652 398 2 1669 1 sky130_fd_sc_hd__dfxtp_1 $T=609500 356320 1 0 $X=609310 $Y=353360
X1293 1 2 1663 410 2 1695 1 sky130_fd_sc_hd__dfxtp_1 $T=621460 323680 1 0 $X=621270 $Y=320720
X1294 1 2 1655 415 2 1702 1 sky130_fd_sc_hd__dfxtp_1 $T=623300 361760 0 0 $X=623110 $Y=361520
X1295 1 2 1699 410 2 1745 1 sky130_fd_sc_hd__dfxtp_1 $T=644920 361760 1 0 $X=644730 $Y=358800
X1296 1 2 451 415 2 1751 1 sky130_fd_sc_hd__dfxtp_1 $T=649060 372640 1 0 $X=648870 $Y=369680
X1297 1 2 1712 410 2 1757 1 sky130_fd_sc_hd__dfxtp_1 $T=651360 329120 0 0 $X=651170 $Y=328880
X1298 1 2 1756 398 2 1777 1 sky130_fd_sc_hd__dfxtp_1 $T=659640 356320 0 0 $X=659450 $Y=356080
X1299 1 2 1756 397 2 1778 1 sky130_fd_sc_hd__dfxtp_1 $T=659640 361760 0 0 $X=659450 $Y=361520
X1300 1 2 454 410 2 1783 1 sky130_fd_sc_hd__dfxtp_1 $T=662860 367200 0 0 $X=662670 $Y=366960
X1301 1 2 1779 400 2 1793 1 sky130_fd_sc_hd__dfxtp_1 $T=667920 345440 0 0 $X=667730 $Y=345200
X1302 1 2 1756 414 2 1804 1 sky130_fd_sc_hd__dfxtp_1 $T=672520 356320 1 0 $X=672330 $Y=353360
X1303 1 2 1779 399 2 1806 1 sky130_fd_sc_hd__dfxtp_1 $T=675280 340000 1 0 $X=675090 $Y=337040
X1304 1 2 1779 415 2 1809 1 sky130_fd_sc_hd__dfxtp_1 $T=677120 350880 1 0 $X=676930 $Y=347920
X1305 1 2 1779 398 2 1816 1 sky130_fd_sc_hd__dfxtp_1 $T=679420 340000 0 0 $X=679230 $Y=339760
X1306 1 2 457 410 2 1825 1 sky130_fd_sc_hd__dfxtp_1 $T=683560 378080 1 0 $X=683370 $Y=375120
X1307 1 2 1862 400 2 1872 1 sky130_fd_sc_hd__dfxtp_1 $T=708860 367200 1 0 $X=708670 $Y=364240
X1308 1 2 467 397 2 1882 1 sky130_fd_sc_hd__dfxtp_1 $T=710240 378080 1 0 $X=710050 $Y=375120
X1309 1 2 1861 415 2 1903 1 sky130_fd_sc_hd__dfxtp_1 $T=724500 340000 0 0 $X=724310 $Y=339760
X1310 1 2 1861 412 2 1905 1 sky130_fd_sc_hd__dfxtp_1 $T=724500 345440 0 0 $X=724310 $Y=345200
X1311 1 2 536 27 38 9 11 535 ICV_13 $T=6900 372640 1 0 $X=6710 $Y=369680
X1312 1 2 550 553 36 531 25 557 ICV_13 $T=18400 329120 0 0 $X=18210 $Y=328880
X1313 1 2 562 533 36 526 14 562 ICV_13 $T=20240 350880 1 0 $X=20050 $Y=347920
X1314 1 2 563 533 57 526 43 561 ICV_13 $T=20240 356320 1 0 $X=20050 $Y=353360
X1315 1 2 570 553 57 531 44 570 ICV_13 $T=22080 329120 1 0 $X=21890 $Y=326160
X1316 1 2 574 553 52 531 43 574 ICV_13 $T=24380 334560 1 0 $X=24190 $Y=331600
X1317 1 2 585 553 54 531 42 585 ICV_13 $T=34040 329120 0 0 $X=33850 $Y=328880
X1318 1 2 581 590 34 575 18 587 ICV_13 $T=34040 350880 0 0 $X=33850 $Y=350640
X1319 1 2 588 590 52 575 43 588 ICV_13 $T=34040 361760 0 0 $X=33850 $Y=361520
X1320 1 2 589 53 33 48 11 589 ICV_13 $T=34040 372640 0 0 $X=33850 $Y=372400
X1321 1 2 594 545 57 524 44 594 ICV_13 $T=36340 323680 1 0 $X=36150 $Y=320720
X1322 1 2 605 590 28 575 25 605 ICV_13 $T=41400 345440 0 0 $X=41210 $Y=345200
X1323 1 2 620 624 37 608 13 621 ICV_13 $T=50140 350880 0 0 $X=49950 $Y=350640
X1324 1 2 634 72 28 591 25 634 ICV_13 $T=54740 318240 1 0 $X=54550 $Y=315280
X1325 1 2 659 664 34 644 13 659 ICV_13 $T=68080 350880 0 0 $X=67890 $Y=350640
X1326 1 2 661 664 28 627 25 663 ICV_13 $T=69460 345440 0 0 $X=69270 $Y=345200
X1327 1 2 669 90 63 83 10 675 ICV_13 $T=76360 372640 1 0 $X=76170 $Y=369680
X1328 1 2 679 664 57 644 44 679 ICV_13 $T=77280 356320 0 0 $X=77090 $Y=356080
X1329 1 2 682 664 52 644 43 682 ICV_13 $T=78200 361760 1 0 $X=78010 $Y=358800
X1330 1 2 691 690 34 672 18 692 ICV_13 $T=82800 334560 1 0 $X=82610 $Y=331600
X1331 1 2 697 699 57 687 25 696 ICV_13 $T=90160 323680 0 0 $X=89970 $Y=323440
X1332 1 2 707 705 57 694 44 707 ICV_13 $T=90160 356320 0 0 $X=89970 $Y=356080
X1333 1 2 726 705 54 694 42 726 ICV_13 $T=101660 356320 0 0 $X=101470 $Y=356080
X1334 1 2 734 705 37 694 18 734 ICV_13 $T=104420 356320 1 0 $X=104230 $Y=353360
X1335 1 2 758 759 39 744 15 758 ICV_13 $T=120520 345440 1 0 $X=120330 $Y=342480
X1336 1 2 760 759 57 744 44 760 ICV_13 $T=120520 356320 1 0 $X=120330 $Y=353360
X1337 1 2 764 747 37 732 44 767 ICV_13 $T=125580 323680 0 0 $X=125390 $Y=323440
X1338 1 2 763 701 54 732 13 769 ICV_13 $T=127420 329120 0 0 $X=127230 $Y=328880
X1339 1 2 766 701 57 750 15 698 ICV_13 $T=132480 340000 1 0 $X=132290 $Y=337040
X1340 1 2 787 791 52 772 25 794 ICV_13 $T=142600 323680 1 0 $X=142410 $Y=320720
X1341 1 2 765 701 28 785 13 802 ICV_13 $T=146280 350880 0 0 $X=146090 $Y=350640
X1342 1 2 806 791 36 772 13 811 ICV_13 $T=152260 318240 0 0 $X=152070 $Y=318000
X1343 1 2 814 783 54 786 42 814 ICV_13 $T=154100 334560 0 0 $X=153910 $Y=334320
X1344 1 2 827 821 174 800 158 823 ICV_13 $T=158700 367200 0 0 $X=158510 $Y=366960
X1345 1 2 813 741 28 160 152 169 ICV_13 $T=160540 378080 1 0 $X=160350 $Y=375120
X1346 1 2 829 830 179 786 15 781 ICV_13 $T=162380 329120 0 0 $X=162190 $Y=328880
X1347 1 2 831 830 184 825 170 832 ICV_13 $T=166520 323680 1 0 $X=166330 $Y=320720
X1348 1 2 847 830 198 173 190 196 ICV_13 $T=178940 312800 0 0 $X=178750 $Y=312560
X1349 1 2 833 820 179 826 191 843 ICV_13 $T=178940 340000 0 0 $X=178750 $Y=339760
X1350 1 2 875 854 186 853 172 875 ICV_13 $T=192740 334560 1 0 $X=192550 $Y=331600
X1351 1 2 885 205 174 195 161 885 ICV_13 $T=199180 378080 1 0 $X=198990 $Y=375120
X1352 1 2 886 205 185 195 163 886 ICV_13 $T=202400 372640 0 0 $X=202210 $Y=372400
X1353 1 2 891 868 188 859 175 891 ICV_13 $T=204700 361760 1 0 $X=204510 $Y=358800
X1354 1 2 895 868 167 859 152 897 ICV_13 $T=206540 367200 0 0 $X=206350 $Y=366960
X1355 1 2 945 911 197 914 187 945 ICV_13 $T=231840 323680 1 0 $X=231650 $Y=320720
X1356 1 2 948 924 174 907 161 948 ICV_13 $T=232300 361760 0 0 $X=232110 $Y=361520
X1357 1 2 962 961 199 939 189 962 ICV_13 $T=238740 345440 0 0 $X=238550 $Y=345200
X1358 1 2 967 958 184 950 191 956 ICV_13 $T=244720 323680 1 0 $X=244530 $Y=320720
X1359 1 2 225 211 167 214 163 969 ICV_13 $T=244720 378080 1 0 $X=244530 $Y=375120
X1360 1 2 970 961 179 939 171 970 ICV_13 $T=245640 350880 0 0 $X=245450 $Y=350640
X1361 1 2 980 958 179 950 170 976 ICV_13 $T=251160 334560 1 0 $X=250970 $Y=331600
X1362 1 2 996 975 180 963 158 996 ICV_13 $T=258520 361760 0 0 $X=258330 $Y=361520
X1363 1 2 998 975 193 963 177 998 ICV_13 $T=258520 372640 0 0 $X=258330 $Y=372400
X1364 1 2 1001 987 179 968 171 1001 ICV_13 $T=260820 356320 1 0 $X=260630 $Y=353360
X1365 1 2 1011 1004 184 995 168 1011 ICV_13 $T=264500 340000 0 0 $X=264310 $Y=339760
X1366 1 2 1016 238 201 233 190 1016 ICV_13 $T=266800 318240 0 0 $X=266610 $Y=318000
X1367 1 2 1027 1004 186 995 172 1027 ICV_13 $T=272780 345440 1 0 $X=272590 $Y=342480
X1368 1 2 1028 1004 201 995 190 1028 ICV_13 $T=272780 356320 1 0 $X=272590 $Y=353360
X1369 1 2 1029 1021 193 1008 177 1029 ICV_13 $T=272780 372640 1 0 $X=272590 $Y=369680
X1370 1 2 1033 1010 197 992 187 1033 ICV_13 $T=274620 334560 0 0 $X=274430 $Y=334320
X1371 1 2 1045 1047 179 1035 171 1045 ICV_13 $T=284740 323680 1 0 $X=284550 $Y=320720
X1372 1 2 1051 1039 199 1030 189 1051 ICV_13 $T=286580 345440 0 0 $X=286390 $Y=345200
X1373 1 2 1052 239 174 1022 161 1052 ICV_13 $T=286580 356320 0 0 $X=286390 $Y=356080
X1374 1 2 1054 245 184 244 168 1054 ICV_13 $T=287500 318240 1 0 $X=287310 $Y=315280
X1375 1 2 1065 1021 176 1008 163 1068 ICV_13 $T=294400 367200 0 0 $X=294210 $Y=366960
X1376 1 2 1063 1021 167 1008 161 1070 ICV_13 $T=295320 361760 0 0 $X=295130 $Y=361520
X1377 1 2 1082 243 176 242 152 1082 ICV_13 $T=300840 378080 1 0 $X=300650 $Y=375120
X1378 1 2 1089 1094 180 1079 158 1089 ICV_13 $T=306360 361760 1 0 $X=306170 $Y=358800
X1379 1 2 1093 1094 193 1079 177 1093 ICV_13 $T=306820 372640 1 0 $X=306630 $Y=369680
X1380 1 2 1097 1076 179 1061 171 1097 ICV_13 $T=309120 350880 1 0 $X=308930 $Y=347920
X1381 1 2 1105 261 267 1095 253 1101 ICV_13 $T=315100 367200 1 0 $X=314910 $Y=364240
X1382 1 2 1128 1094 174 1079 161 1128 ICV_13 $T=328900 361760 1 0 $X=328710 $Y=358800
X1383 1 2 1108 1083 166 1118 273 1135 ICV_13 $T=330740 329120 0 0 $X=330550 $Y=328880
X1384 1 2 1141 1131 263 278 273 1143 ICV_13 $T=334880 318240 1 0 $X=334690 $Y=315280
X1385 1 2 1154 1120 268 1102 253 1149 ICV_13 $T=341320 350880 1 0 $X=341130 $Y=347920
X1386 1 2 1126 1131 296 165 176 290 ICV_13 $T=342240 356320 1 0 $X=342050 $Y=353360
X1387 1 2 1153 1158 269 1146 253 1155 ICV_13 $T=342700 361760 0 0 $X=342510 $Y=361520
X1388 1 2 1163 1131 268 165 193 298 ICV_13 $T=348220 350880 0 0 $X=348030 $Y=350640
X1389 1 2 1195 1186 277 1171 265 1195 ICV_13 $T=365700 334560 1 0 $X=365510 $Y=331600
X1390 1 2 1209 1188 275 1187 266 1209 ICV_13 $T=371680 356320 1 0 $X=371490 $Y=353360
X1391 1 2 1220 1188 267 1187 257 1216 ICV_13 $T=377660 350880 0 0 $X=377470 $Y=350640
X1392 1 2 1228 1223 267 1203 273 1232 ICV_13 $T=385020 340000 1 0 $X=384830 $Y=337040
X1393 1 2 1233 319 267 312 260 1233 ICV_13 $T=385020 372640 1 0 $X=384830 $Y=369680
X1394 1 2 1235 1188 263 1187 253 1235 ICV_13 $T=386400 361760 0 0 $X=386210 $Y=361520
X1395 1 2 1240 328 263 325 253 1240 ICV_13 $T=389160 318240 1 0 $X=388970 $Y=315280
X1396 1 2 1243 1225 275 1205 266 1243 ICV_13 $T=390540 345440 1 0 $X=390350 $Y=342480
X1397 1 2 1244 1250 296 1229 260 1252 ICV_13 $T=393760 323680 1 0 $X=393570 $Y=320720
X1398 1 2 1254 1250 280 1229 273 1254 ICV_13 $T=394220 329120 1 0 $X=394030 $Y=326160
X1399 1 2 1262 1227 277 1230 265 1262 ICV_13 $T=398360 367200 1 0 $X=398170 $Y=364240
X1400 1 2 1264 333 277 329 265 1264 ICV_13 $T=398820 372640 0 0 $X=398630 $Y=372400
X1401 1 2 1265 1256 277 1249 264 1255 ICV_13 $T=399740 334560 1 0 $X=399550 $Y=331600
X1402 1 2 1281 1250 275 1229 253 1267 ICV_13 $T=408020 323680 0 0 $X=407830 $Y=323440
X1403 1 2 1278 1261 275 1257 266 1278 ICV_13 $T=408020 345440 0 0 $X=407830 $Y=345200
X1404 1 2 1288 1256 269 1249 253 1286 ICV_13 $T=413080 340000 1 0 $X=412890 $Y=337040
X1405 1 2 1286 1256 263 1229 265 1283 ICV_13 $T=414460 329120 0 0 $X=414270 $Y=328880
X1406 1 2 346 347 275 339 265 344 ICV_13 $T=416760 378080 1 0 $X=416570 $Y=375120
X1407 1 2 1303 1295 267 1284 260 1303 ICV_13 $T=419520 323680 1 0 $X=419330 $Y=320720
X1408 1 2 1305 1306 275 343 266 1305 ICV_13 $T=420440 372640 1 0 $X=420250 $Y=369680
X1409 1 2 1325 349 296 342 264 1325 ICV_13 $T=431020 312800 0 0 $X=430830 $Y=312560
X1410 1 2 1338 1308 268 1294 257 1338 ICV_13 $T=438380 350880 0 0 $X=438190 $Y=350640
X1411 1 2 1345 1350 275 1331 266 1345 ICV_13 $T=442980 323680 0 0 $X=442790 $Y=323440
X1412 1 2 1349 1342 269 1334 262 1349 ICV_13 $T=442980 361760 0 0 $X=442790 $Y=361520
X1413 1 2 361 358 269 359 257 1365 ICV_13 $T=451260 378080 1 0 $X=451070 $Y=375120
X1414 1 2 1372 1371 275 1360 266 1372 ICV_13 $T=454480 340000 1 0 $X=454290 $Y=337040
X1415 1 2 1376 360 275 356 266 1376 ICV_13 $T=455860 318240 1 0 $X=455670 $Y=315280
X1416 1 2 1403 1400 275 1384 266 1403 ICV_13 $T=469200 356320 1 0 $X=469010 $Y=353360
X1417 1 2 1442 1434 280 1429 264 1432 ICV_13 $T=488980 367200 0 0 $X=488790 $Y=366960
X1418 1 2 1454 381 267 378 260 1454 ICV_13 $T=490360 312800 0 0 $X=490170 $Y=312560
X1419 1 2 1464 382 277 377 265 1464 ICV_13 $T=501400 378080 1 0 $X=501210 $Y=375120
X1420 1 2 1480 1456 275 1431 266 1480 ICV_13 $T=505540 356320 1 0 $X=505350 $Y=353360
X1421 1 2 1498 1503 407 1486 400 1498 ICV_13 $T=518880 345440 0 0 $X=518690 $Y=345200
X1422 1 2 1492 1507 409 1484 400 1499 ICV_13 $T=519340 318240 0 0 $X=519150 $Y=318000
X1423 1 2 1494 1506 409 1485 399 1501 ICV_13 $T=519340 329120 0 0 $X=519150 $Y=328880
X1424 1 2 1510 1509 408 1496 399 1510 ICV_13 $T=525320 356320 1 0 $X=525130 $Y=353360
X1425 1 2 1511 1506 405 1485 398 1511 ICV_13 $T=526700 334560 0 0 $X=526510 $Y=334320
X1426 1 2 1522 1506 422 1485 414 1522 ICV_13 $T=531760 329120 1 0 $X=531570 $Y=326160
X1427 1 2 420 406 418 1484 414 1526 ICV_13 $T=534060 318240 1 0 $X=533870 $Y=315280
X1428 1 2 1521 1503 424 1486 415 1514 ICV_13 $T=539120 345440 1 0 $X=538930 $Y=342480
X1429 1 2 1549 1542 422 1529 398 1553 ICV_13 $T=552920 329120 0 0 $X=552730 $Y=328880
X1430 1 2 1559 1557 408 1551 399 1559 ICV_13 $T=553380 361760 1 0 $X=553190 $Y=358800
X1431 1 2 1567 1542 408 1529 415 1563 ICV_13 $T=555220 329120 1 0 $X=555030 $Y=326160
X1432 1 2 1558 1557 405 1551 410 1576 ICV_13 $T=560740 356320 1 0 $X=560550 $Y=353360
X1433 1 2 1584 1557 407 1551 400 1584 ICV_13 $T=566260 361760 1 0 $X=566070 $Y=358800
X1434 1 2 1592 1557 422 1551 414 1592 ICV_13 $T=567180 356320 0 0 $X=566990 $Y=356080
X1435 1 2 1593 1557 418 1551 415 1593 ICV_13 $T=567180 361760 0 0 $X=566990 $Y=361520
X1436 1 2 1581 426 424 1540 410 433 ICV_13 $T=567180 372640 0 0 $X=566990 $Y=372400
X1437 1 2 1606 1585 405 1575 398 1606 ICV_13 $T=574080 350880 0 0 $X=573890 $Y=350640
X1438 1 2 1613 1599 424 1578 412 1613 ICV_13 $T=578680 318240 0 0 $X=578490 $Y=318000
X1439 1 2 1621 1604 422 1602 415 1619 ICV_13 $T=580520 367200 0 0 $X=580330 $Y=366960
X1440 1 2 1629 1599 408 1578 399 1629 ICV_13 $T=586960 323680 1 0 $X=586770 $Y=320720
X1441 1 2 1634 1633 407 1618 400 1634 ICV_13 $T=589260 334560 1 0 $X=589070 $Y=331600
X1442 1 2 1637 1633 405 1618 398 1637 ICV_13 $T=590640 329120 1 0 $X=590450 $Y=326160
X1443 1 2 1641 1616 408 1612 399 1641 ICV_13 $T=594320 350880 1 0 $X=594130 $Y=347920
X1444 1 2 1646 1616 424 1612 412 1646 ICV_13 $T=595240 345440 0 0 $X=595050 $Y=345200
X1445 1 2 1659 1633 422 1618 414 1659 ICV_13 $T=599840 329120 0 0 $X=599650 $Y=328880
X1446 1 2 1676 1682 405 1663 398 1676 ICV_13 $T=611340 323680 0 0 $X=611150 $Y=323440
X1447 1 2 1677 1682 407 1663 400 1677 ICV_13 $T=611340 329120 0 0 $X=611150 $Y=328880
X1448 1 2 1690 1665 424 1652 412 1690 ICV_13 $T=616860 356320 1 0 $X=616670 $Y=353360
X1449 1 2 1691 1668 409 1655 397 1691 ICV_13 $T=616860 372640 1 0 $X=616670 $Y=369680
X1450 1 2 1698 1682 408 1663 397 1703 ICV_13 $T=623760 329120 1 0 $X=623570 $Y=326160
X1451 1 2 1726 1719 407 1712 400 1726 ICV_13 $T=635260 323680 0 0 $X=635070 $Y=323440
X1452 1 2 1729 1719 408 1712 399 1729 ICV_13 $T=637560 329120 1 0 $X=637370 $Y=326160
X1453 1 2 1727 1722 424 1713 397 1725 ICV_13 $T=637560 350880 1 0 $X=637370 $Y=347920
X1454 1 2 1715 450 417 447 415 1731 ICV_13 $T=637560 372640 1 0 $X=637370 $Y=369680
X1455 1 2 1732 445 424 446 399 1733 ICV_13 $T=638480 318240 0 0 $X=638290 $Y=318000
X1456 1 2 1757 1719 417 1720 399 1755 ICV_13 $T=650900 334560 1 0 $X=650710 $Y=331600
X1457 1 2 1759 453 417 451 410 1759 ICV_13 $T=651360 367200 0 0 $X=651170 $Y=366960
X1458 1 2 1760 453 422 451 414 1760 ICV_13 $T=651360 372640 0 0 $X=651170 $Y=372400
X1459 1 2 1762 453 407 451 400 1762 ICV_13 $T=652280 367200 1 0 $X=652090 $Y=364240
X1460 1 2 1763 1749 407 1747 400 1763 ICV_13 $T=653200 318240 0 0 $X=653010 $Y=318000
X1461 1 2 1769 1749 408 1747 415 1768 ICV_13 $T=655500 312800 0 0 $X=655310 $Y=312560
X1462 1 2 1788 1781 408 1775 399 1788 ICV_13 $T=666540 329120 0 0 $X=666350 $Y=328880
X1463 1 2 1791 1780 417 1756 410 1791 ICV_13 $T=667000 356320 0 0 $X=666810 $Y=356080
X1464 1 2 1789 1749 417 1775 398 1782 ICV_13 $T=667460 329120 1 0 $X=667270 $Y=326160
X1465 1 2 1802 455 407 454 400 1802 ICV_13 $T=672060 372640 1 0 $X=671870 $Y=369680
X1466 1 2 1815 456 409 1801 410 1811 ICV_13 $T=679420 318240 0 0 $X=679230 $Y=318000
X1467 1 2 1817 1780 407 1756 400 1817 ICV_13 $T=679880 356320 1 0 $X=679690 $Y=353360
X1468 1 2 1820 1781 424 1775 397 1813 ICV_13 $T=680340 334560 1 0 $X=680150 $Y=331600
X1469 1 2 1836 1781 422 1775 410 1840 ICV_13 $T=693680 334560 1 0 $X=693490 $Y=331600
X1470 1 2 1841 1818 422 1808 414 1841 ICV_13 $T=693680 350880 0 0 $X=693490 $Y=350640
X1471 1 2 1842 1818 418 1808 415 1842 ICV_13 $T=693680 356320 1 0 $X=693490 $Y=353360
X1472 1 2 1848 462 424 457 412 1848 ICV_13 $T=695520 372640 1 0 $X=695330 $Y=369680
X1473 1 2 1839 1781 418 1850 397 1863 ICV_13 $T=702880 329120 1 0 $X=702690 $Y=326160
X1474 1 2 1866 1871 407 1860 400 1866 ICV_13 $T=707480 356320 0 0 $X=707290 $Y=356080
X1475 1 2 1865 469 407 466 397 1873 ICV_13 $T=709320 312800 0 0 $X=709130 $Y=312560
X1476 1 2 1858 1827 405 1861 400 1874 ICV_13 $T=709320 345440 0 0 $X=709130 $Y=345200
X1477 1 2 1884 1889 422 1859 397 1876 ICV_13 $T=709780 334560 1 0 $X=709590 $Y=331600
X1478 1 2 1878 1871 409 1860 397 1878 ICV_13 $T=709780 361760 1 0 $X=709590 $Y=358800
X1479 1 2 1894 1871 417 1860 410 1894 ICV_13 $T=721740 361760 1 0 $X=721550 $Y=358800
X1480 1 2 1898 1869 418 1850 415 1898 ICV_13 $T=722200 329120 0 0 $X=722010 $Y=328880
X1481 1 2 1899 1871 408 1860 399 1899 ICV_13 $T=722200 356320 0 0 $X=722010 $Y=356080
X1482 1 2 1882 468 409 467 415 1918 ICV_13 $T=731400 378080 1 0 $X=731210 $Y=375120
X1483 1 2 524 18 540 540 545 37 ICV_14 $T=6900 318240 0 0 $X=6710 $Y=318000
X1484 1 2 526 13 542 547 533 37 ICV_14 $T=6900 350880 1 0 $X=6710 $Y=347920
X1485 1 2 41 25 566 566 51 28 ICV_14 $T=20240 318240 1 0 $X=20050 $Y=315280
X1486 1 2 602 11 613 615 609 47 ICV_14 $T=45080 367200 0 0 $X=44890 $Y=366960
X1487 1 2 637 43 676 676 653 52 ICV_14 $T=76360 318240 0 0 $X=76170 $Y=318000
X1488 1 2 672 14 693 693 690 36 ICV_14 $T=81880 340000 1 0 $X=81690 $Y=337040
X1489 1 2 800 156 818 818 821 167 ICV_14 $T=155020 372640 0 0 $X=154830 $Y=372400
X1490 1 2 884 168 901 893 888 197 ICV_14 $T=206540 334560 0 0 $X=206350 $Y=334320
X1491 1 2 884 191 892 896 888 166 ICV_14 $T=206540 340000 0 0 $X=206350 $Y=339760
X1492 1 2 884 190 902 902 888 201 ICV_14 $T=206540 350880 0 0 $X=206350 $Y=350640
X1493 1 2 992 170 1034 1034 1010 166 ICV_14 $T=274160 334560 1 0 $X=273970 $Y=331600
X1494 1 2 1118 266 1130 1135 1138 280 ICV_14 $T=328900 323680 1 0 $X=328710 $Y=320720
X1495 1 2 278 257 1176 1177 289 269 ICV_14 $T=351900 318240 0 0 $X=351710 $Y=318000
X1496 1 2 1169 273 1194 1198 1173 263 ICV_14 $T=364320 350880 1 0 $X=364130 $Y=347920
X1497 1 2 1205 273 1242 1242 1225 280 ICV_14 $T=389160 350880 1 0 $X=388970 $Y=347920
X1498 1 2 1249 266 1287 1287 1256 275 ICV_14 $T=412160 340000 0 0 $X=411970 $Y=339760
X1499 1 2 343 273 1319 1319 1306 280 ICV_14 $T=428260 378080 1 0 $X=428070 $Y=375120
X1500 1 2 1334 253 1340 1329 1306 296 ICV_14 $T=441600 367200 0 0 $X=441410 $Y=366960
X1501 1 2 356 257 1355 1351 360 280 ICV_14 $T=443440 318240 1 0 $X=443250 $Y=315280
X1502 1 2 1331 262 1363 1366 1350 280 ICV_14 $T=450340 329120 1 0 $X=450150 $Y=326160
X1503 1 2 1331 253 1367 1368 1350 267 ICV_14 $T=451260 334560 1 0 $X=451070 $Y=331600
X1504 1 2 356 253 1377 1377 360 263 ICV_14 $T=454940 318240 0 0 $X=454750 $Y=318000
X1505 1 2 378 257 1467 1466 381 275 ICV_14 $T=501400 318240 1 0 $X=501210 $Y=315280
X1506 1 2 1496 414 1532 1532 1509 422 ICV_14 $T=539120 350880 0 0 $X=538930 $Y=350640
X1507 1 2 1578 414 1601 1601 1599 422 ICV_14 $T=571320 312800 0 0 $X=571130 $Y=312560
X1508 1 2 1602 397 1635 1635 1604 409 ICV_14 $T=588800 361760 1 0 $X=588610 $Y=358800
X1509 1 2 1661 414 1705 1705 1678 422 ICV_14 $T=623760 340000 1 0 $X=623570 $Y=337040
X1510 1 2 1712 398 1752 1754 1719 409 ICV_14 $T=649060 329120 1 0 $X=648870 $Y=326160
X1511 1 2 1747 412 1787 1787 1749 424 ICV_14 $T=665620 323680 1 0 $X=665430 $Y=320720
X1512 1 2 1779 412 1790 1790 1797 424 ICV_14 $T=666080 340000 0 0 $X=665890 $Y=339760
X1513 1 2 1801 412 1812 1812 456 424 ICV_14 $T=678040 323680 1 0 $X=677850 $Y=320720
X1514 1 2 1859 414 1884 1863 1869 409 ICV_14 $T=709780 329120 0 0 $X=709590 $Y=328880
X1515 1 2 1860 415 1900 1901 1871 424 ICV_14 $T=721740 356320 1 0 $X=721550 $Y=353360
X1516 1 2 524 13 537 537 545 34 ICV_16 $T=6900 318240 1 0 $X=6710 $Y=315280
X1517 1 2 524 14 538 538 545 36 ICV_16 $T=6900 323680 1 0 $X=6710 $Y=320720
X1518 1 2 524 15 539 539 545 39 ICV_16 $T=6900 329120 1 0 $X=6710 $Y=326160
X1519 1 2 524 25 552 549 553 34 ICV_16 $T=12420 323680 0 0 $X=12230 $Y=323440
X1520 1 2 524 43 560 560 545 52 ICV_16 $T=19320 318240 0 0 $X=19130 $Y=318000
X1521 1 2 41 15 64 65 51 34 ICV_16 $T=32660 318240 1 0 $X=32470 $Y=315280
X1522 1 2 531 18 584 584 553 37 ICV_16 $T=33580 329120 1 0 $X=33390 $Y=326160
X1523 1 2 627 13 665 647 645 36 ICV_16 $T=69460 334560 0 0 $X=69270 $Y=334320
X1524 1 2 118 42 753 753 126 54 ICV_16 $T=118220 312800 0 0 $X=118030 $Y=312560
X1525 1 2 786 43 798 801 783 57 ICV_16 $T=145360 340000 1 0 $X=145170 $Y=337040
X1526 1 2 853 189 869 862 854 166 ICV_16 $T=191820 318240 1 0 $X=191630 $Y=315280
X1527 1 2 855 168 877 867 852 166 ICV_16 $T=192740 340000 1 0 $X=192550 $Y=337040
X1528 1 2 882 168 898 898 887 184 ICV_16 $T=206540 323680 0 0 $X=206350 $Y=323440
X1529 1 2 884 172 899 899 888 186 ICV_16 $T=206540 345440 0 0 $X=206350 $Y=345200
X1530 1 2 882 172 905 908 911 198 ICV_16 $T=210680 318240 0 0 $X=210490 $Y=318000
X1531 1 2 907 181 943 942 924 185 ICV_16 $T=230460 372640 1 0 $X=230270 $Y=369680
X1532 1 2 968 172 988 982 987 197 ICV_16 $T=253000 345440 1 0 $X=252810 $Y=342480
X1533 1 2 992 172 1007 1007 1010 186 ICV_16 $T=262660 329120 0 0 $X=262470 $Y=328880
X1534 1 2 250 189 1106 1106 254 199 ICV_16 $T=316020 318240 0 0 $X=315830 $Y=318000
X1535 1 2 1095 266 1129 1129 261 275 ICV_16 $T=328900 367200 0 0 $X=328710 $Y=366960
X1536 1 2 1146 266 1159 1159 1158 275 ICV_16 $T=343160 367200 1 0 $X=342970 $Y=364240
X1537 1 2 1112 273 1165 1165 1131 280 ICV_16 $T=345000 334560 0 0 $X=344810 $Y=334320
X1538 1 2 1169 262 1196 1192 1173 277 ICV_16 $T=365240 340000 1 0 $X=365050 $Y=337040
X1539 1 2 1205 260 1219 1219 1225 267 ICV_16 $T=378120 345440 0 0 $X=377930 $Y=345200
X1540 1 2 1205 257 1222 1222 1225 268 ICV_16 $T=378580 340000 0 0 $X=378390 $Y=339760
X1541 1 2 325 264 1272 1270 328 269 ICV_16 $T=402960 312800 0 0 $X=402770 $Y=312560
X1542 1 2 1360 264 1369 1373 1371 263 ICV_16 $T=453560 345440 1 0 $X=453370 $Y=342480
X1543 1 2 1385 257 1395 368 370 277 ICV_16 $T=465520 372640 0 0 $X=465330 $Y=372400
X1544 1 2 1378 257 1416 1416 1382 268 ICV_16 $T=476560 323680 1 0 $X=476370 $Y=320720
X1545 1 2 1429 265 1465 1465 1434 277 ICV_16 $T=501400 372640 1 0 $X=501210 $Y=369680
X1546 1 2 1486 410 1524 1516 1509 417 ICV_16 $T=532220 350880 1 0 $X=532030 $Y=347920
X1547 1 2 1496 398 1531 1531 1509 405 ICV_16 $T=539120 356320 0 0 $X=538930 $Y=356080
X1548 1 2 1551 397 1566 1569 426 405 ICV_16 $T=554760 361760 0 0 $X=554570 $Y=361520
X1549 1 2 1540 398 1569 1570 426 409 ICV_16 $T=555680 367200 1 0 $X=555490 $Y=364240
X1550 1 2 1574 414 1582 1582 1580 422 ICV_16 $T=565800 334560 1 0 $X=565610 $Y=331600
X1551 1 2 1602 412 1615 1617 1604 407 ICV_16 $T=578680 361760 0 0 $X=578490 $Y=361520
X1552 1 2 434 400 1647 1647 437 407 ICV_16 $T=595240 378080 1 0 $X=595050 $Y=375120
X1553 1 2 434 399 1648 1648 437 408 ICV_16 $T=595700 372640 1 0 $X=595510 $Y=369680
X1554 1 2 1640 398 1656 1658 439 409 ICV_16 $T=599380 318240 0 0 $X=599190 $Y=318000
X1555 1 2 1640 397 1658 1657 439 408 ICV_16 $T=599380 323680 0 0 $X=599190 $Y=323440
X1556 1 2 1640 400 1681 1680 439 422 ICV_16 $T=611800 318240 1 0 $X=611610 $Y=315280
X1557 1 2 1663 412 1704 1704 1682 424 ICV_16 $T=623300 323680 0 0 $X=623110 $Y=323440
X1558 1 2 1720 414 1736 1736 1740 422 ICV_16 $T=638480 340000 0 0 $X=638290 $Y=339760
X1559 1 2 1756 399 1798 1795 1780 424 ICV_16 $T=667920 361760 1 0 $X=667730 $Y=358800
X1560 1 2 1814 397 1851 1857 1827 424 ICV_16 $T=697820 340000 1 0 $X=697630 $Y=337040
X1561 1 2 1850 412 1895 1895 1869 424 ICV_16 $T=721740 323680 1 0 $X=721550 $Y=320720
X1562 1 2 1850 399 1896 1879 1869 405 ICV_16 $T=721740 323680 0 0 $X=721550 $Y=323440
X1563 1 2 525 15 544 541 548 36 ICV_17 $T=6900 340000 1 0 $X=6710 $Y=337040
X1564 1 2 526 42 558 558 533 54 ICV_17 $T=17480 356320 0 0 $X=17290 $Y=356080
X1565 1 2 580 44 599 599 596 57 ICV_17 $T=36340 340000 0 0 $X=36150 $Y=339760
X1566 1 2 580 25 616 616 596 28 ICV_17 $T=47840 334560 0 0 $X=47650 $Y=334320
X1567 1 2 602 10 639 641 609 55 ICV_17 $T=57040 372640 1 0 $X=56850 $Y=369680
X1568 1 2 637 18 668 668 653 37 ICV_17 $T=70380 323680 0 0 $X=70190 $Y=323440
X1569 1 2 94 42 735 735 96 54 ICV_17 $T=104420 318240 1 0 $X=104230 $Y=315280
X1570 1 2 173 172 183 832 830 166 ICV_17 $T=167900 318240 1 0 $X=167710 $Y=315280
X1571 1 2 195 181 856 856 205 194 ICV_17 $T=183540 367200 0 0 $X=183350 $Y=366960
X1572 1 2 914 168 944 944 911 184 ICV_17 $T=230460 318240 0 0 $X=230270 $Y=318000
X1573 1 2 914 189 946 946 911 199 ICV_17 $T=230460 323680 0 0 $X=230270 $Y=323440
X1574 1 2 963 181 991 991 975 194 ICV_17 $T=253920 367200 1 0 $X=253730 $Y=364240
X1575 1 2 165 75 241 1023 1021 180 ICV_17 $T=269560 356320 0 0 $X=269370 $Y=356080
X1576 1 2 1061 191 1075 1077 1076 184 ICV_17 $T=296700 340000 0 0 $X=296510 $Y=339760
X1577 1 2 1079 175 1142 1142 1094 188 ICV_17 $T=333040 372640 1 0 $X=332850 $Y=369680
X1578 1 2 1203 253 1237 1236 1223 268 ICV_17 $T=385480 329120 0 0 $X=385290 $Y=328880
X1579 1 2 1249 273 1266 1266 1256 280 ICV_17 $T=398820 334560 0 0 $X=398630 $Y=334320
X1580 1 2 1301 257 1311 1314 1313 269 ICV_17 $T=424580 340000 1 0 $X=424390 $Y=337040
X1581 1 2 1331 265 1347 1346 1350 268 ICV_17 $T=441600 329120 0 0 $X=441410 $Y=328880
X1582 1 2 1428 260 1447 1439 1450 296 ICV_17 $T=487600 329120 0 0 $X=487410 $Y=328880
X1583 1 2 1413 253 1479 1472 1456 268 ICV_17 $T=503700 350880 1 0 $X=503510 $Y=347920
X1584 1 2 1551 398 1558 1533 1509 418 ICV_17 $T=551080 356320 0 0 $X=550890 $Y=356080
X1585 1 2 434 414 1622 1622 437 422 ICV_17 $T=580980 372640 0 0 $X=580790 $Y=372400
X1586 1 2 434 397 1650 1650 437 409 ICV_17 $T=595240 372640 0 0 $X=595050 $Y=372400
X1587 1 2 1640 410 438 1656 439 405 ICV_17 $T=599380 312800 0 0 $X=599190 $Y=312560
X1588 1 2 1652 410 1662 1669 1665 405 ICV_17 $T=603520 350880 0 0 $X=603330 $Y=350640
X1589 1 2 1661 400 1675 1675 1678 407 ICV_17 $T=609500 345440 1 0 $X=609310 $Y=342480
X1590 1 2 1663 399 1698 1701 1682 422 ICV_17 $T=620540 334560 1 0 $X=620350 $Y=331600
X1591 1 2 1661 415 1700 1708 1678 409 ICV_17 $T=623300 340000 0 0 $X=623110 $Y=339760
X1592 1 2 1720 398 1735 1735 1740 405 ICV_17 $T=637560 340000 1 0 $X=637370 $Y=337040
X1593 1 2 451 412 1753 1753 453 424 ICV_17 $T=649060 378080 1 0 $X=648870 $Y=375120
X1594 1 2 1747 398 1785 1786 1749 422 ICV_17 $T=664700 318240 0 0 $X=664510 $Y=318000
X1595 1 2 1814 410 1832 1833 1827 422 ICV_17 $T=686780 340000 0 0 $X=686590 $Y=339760
X1596 1 2 1859 412 1902 1902 1889 424 ICV_17 $T=723120 334560 1 0 $X=722930 $Y=331600
X1597 1 2 1862 415 1916 1916 1881 418 ICV_17 $T=725880 367200 1 0 $X=725690 $Y=364240
X1598 1 2 531 13 549 ICV_20 $T=10580 329120 0 0 $X=10390 $Y=328880
X1599 1 2 531 14 550 ICV_20 $T=10580 334560 1 0 $X=10390 $Y=331600
X1600 1 2 9 40 556 ICV_20 $T=17020 367200 0 0 $X=16830 $Y=366960
X1601 1 2 525 18 565 ICV_20 $T=20240 340000 1 0 $X=20050 $Y=337040
X1602 1 2 524 42 579 ICV_20 $T=28520 323680 1 0 $X=28330 $Y=320720
X1603 1 2 591 14 606 ICV_20 $T=41860 318240 0 0 $X=41670 $Y=318000
X1604 1 2 66 18 73 ICV_20 $T=44160 312800 0 0 $X=43970 $Y=312560
X1605 1 2 608 14 622 ICV_20 $T=50140 350880 1 0 $X=49950 $Y=347920
X1606 1 2 608 25 628 ICV_20 $T=52900 345440 0 0 $X=52710 $Y=345200
X1607 1 2 591 42 623 ICV_20 $T=54280 323680 1 0 $X=54090 $Y=320720
X1608 1 2 83 11 666 ICV_20 $T=69460 367200 0 0 $X=69270 $Y=366960
X1609 1 2 644 15 685 ICV_20 $T=79120 356320 1 0 $X=78930 $Y=353360
X1610 1 2 98 20 718 ICV_20 $T=94300 372640 0 0 $X=94110 $Y=372400
X1611 1 2 98 11 719 ICV_20 $T=94760 372640 1 0 $X=94570 $Y=369680
X1612 1 2 94 15 101 ICV_20 $T=96140 318240 1 0 $X=95950 $Y=315280
X1613 1 2 720 43 724 ICV_20 $T=102120 345440 0 0 $X=101930 $Y=345200
X1614 1 2 94 43 115 ICV_20 $T=107640 312800 0 0 $X=107450 $Y=312560
X1615 1 2 744 18 761 ICV_20 $T=120520 345440 0 0 $X=120330 $Y=345200
X1616 1 2 750 44 766 ICV_20 $T=124660 334560 0 0 $X=124470 $Y=334320
X1617 1 2 750 18 784 ICV_20 $T=135240 334560 0 0 $X=135050 $Y=334320
X1618 1 2 772 14 806 ICV_20 $T=148580 318240 1 0 $X=148390 $Y=315280
X1619 1 2 772 15 810 ICV_20 $T=150880 329120 1 0 $X=150690 $Y=326160
X1620 1 2 785 25 813 ICV_20 $T=153180 345440 0 0 $X=152990 $Y=345200
X1621 1 2 785 42 807 ICV_20 $T=153640 356320 0 0 $X=153450 $Y=356080
X1622 1 2 825 191 847 ICV_20 $T=178020 323680 1 0 $X=177830 $Y=320720
X1623 1 2 853 191 864 ICV_20 $T=191360 323680 1 0 $X=191170 $Y=320720
X1624 1 2 859 181 879 ICV_20 $T=194580 367200 1 0 $X=194390 $Y=364240
X1625 1 2 882 190 912 ICV_20 $T=212520 329120 0 0 $X=212330 $Y=328880
X1626 1 2 165 49 221 ICV_20 $T=223100 356320 1 0 $X=222910 $Y=353360
X1627 1 2 165 47 222 ICV_20 $T=235060 361760 1 0 $X=234870 $Y=358800
X1628 1 2 939 190 960 ICV_20 $T=237820 350880 0 0 $X=237630 $Y=350640
X1629 1 2 968 191 983 ICV_20 $T=250240 345440 0 0 $X=250050 $Y=345200
X1630 1 2 950 172 985 ICV_20 $T=252080 329120 1 0 $X=251890 $Y=326160
X1631 1 2 165 33 235 ICV_20 $T=261740 356320 0 0 $X=261550 $Y=356080
X1632 1 2 233 171 1012 ICV_20 $T=264500 318240 1 0 $X=264310 $Y=315280
X1633 1 2 992 190 1025 ICV_20 $T=272780 329120 1 0 $X=272590 $Y=326160
X1634 1 2 1008 156 1063 ICV_20 $T=292560 361760 1 0 $X=292370 $Y=358800
X1635 1 2 1035 189 1067 ICV_20 $T=293940 329120 0 0 $X=293750 $Y=328880
X1636 1 2 242 163 1080 ICV_20 $T=299000 372640 0 0 $X=298810 $Y=372400
X1637 1 2 1061 170 1099 ICV_20 $T=310040 340000 1 0 $X=309850 $Y=337040
X1638 1 2 1095 262 1109 ICV_20 $T=317400 372640 0 0 $X=317210 $Y=372400
X1639 1 2 1102 262 1116 ICV_20 $T=320620 350880 1 0 $X=320430 $Y=347920
X1640 1 2 165 180 302 ICV_20 $T=352820 356320 0 0 $X=352630 $Y=356080
X1641 1 2 1146 260 1174 ICV_20 $T=352820 367200 0 0 $X=352630 $Y=366960
X1642 1 2 1171 260 1182 ICV_20 $T=357420 323680 0 0 $X=357230 $Y=323440
X1643 1 2 1205 253 1215 ICV_20 $T=376740 350880 1 0 $X=376550 $Y=347920
X1644 1 2 1187 260 1220 ICV_20 $T=378120 356320 0 0 $X=377930 $Y=356080
X1645 1 2 165 167 326 ICV_20 $T=386860 356320 1 0 $X=386670 $Y=353360
X1646 1 2 1205 262 1245 ICV_20 $T=390540 340000 0 0 $X=390350 $Y=339760
X1647 1 2 1229 257 1277 ICV_20 $T=406640 329120 0 0 $X=406450 $Y=328880
X1648 1 2 1257 262 1292 ICV_20 $T=415840 350880 1 0 $X=415650 $Y=347920
X1649 1 2 1284 273 1300 ICV_20 $T=418600 318240 0 0 $X=418410 $Y=318000
X1650 1 2 1294 264 1307 ICV_20 $T=422280 361760 1 0 $X=422090 $Y=358800
X1651 1 2 1284 262 1321 ICV_20 $T=429640 318240 0 0 $X=429450 $Y=318000
X1652 1 2 1284 257 1327 ICV_20 $T=431020 323680 1 0 $X=430830 $Y=320720
X1653 1 2 1301 253 1336 ICV_20 $T=437000 334560 0 0 $X=436810 $Y=334320
X1654 1 2 1334 260 1370 ICV_20 $T=453100 372640 1 0 $X=452910 $Y=369680
X1655 1 2 1334 266 1375 ICV_20 $T=454940 361760 0 0 $X=454750 $Y=361520
X1656 1 2 1339 265 1387 ICV_20 $T=459540 350880 1 0 $X=459350 $Y=347920
X1657 1 2 1378 266 1388 ICV_20 $T=462300 323680 0 0 $X=462110 $Y=323440
X1658 1 2 1384 262 1394 ICV_20 $T=465520 356320 0 0 $X=465330 $Y=356080
X1659 1 2 1385 266 1405 ICV_20 $T=469200 367200 1 0 $X=469010 $Y=364240
X1660 1 2 1378 265 1414 ICV_20 $T=476100 329120 1 0 $X=475910 $Y=326160
X1661 1 2 1385 265 1420 ICV_20 $T=477480 378080 1 0 $X=477290 $Y=375120
X1662 1 2 1384 253 1415 ICV_20 $T=478400 350880 1 0 $X=478210 $Y=347920
X1663 1 2 1428 262 1438 ICV_20 $T=487140 334560 0 0 $X=486950 $Y=334320
X1664 1 2 1429 273 1442 ICV_20 $T=488060 367200 1 0 $X=487870 $Y=364240
X1665 1 2 1429 262 1443 ICV_20 $T=488060 372640 1 0 $X=487870 $Y=369680
X1666 1 2 1430 262 1444 ICV_20 $T=488520 323680 1 0 $X=488330 $Y=320720
X1667 1 2 1429 260 1448 ICV_20 $T=488520 372640 0 0 $X=488330 $Y=372400
X1668 1 2 378 266 1466 ICV_20 $T=501860 312800 0 0 $X=501670 $Y=312560
X1669 1 2 1430 265 1468 ICV_20 $T=502780 323680 0 0 $X=502590 $Y=323440
X1670 1 2 1484 398 1493 ICV_20 $T=517040 323680 1 0 $X=516850 $Y=320720
X1671 1 2 1484 410 1513 ICV_20 $T=530840 318240 0 0 $X=530650 $Y=318000
X1672 1 2 1527 410 1539 ICV_20 $T=543260 334560 0 0 $X=543070 $Y=334320
X1673 1 2 1529 400 1537 ICV_20 $T=544640 323680 0 0 $X=544450 $Y=323440
X1674 1 2 1529 399 1567 ICV_20 $T=555220 323680 1 0 $X=555030 $Y=320720
X1675 1 2 1574 410 1588 ICV_20 $T=566720 329120 1 0 $X=566530 $Y=326160
X1676 1 2 1578 415 1627 ICV_20 $T=585580 318240 1 0 $X=585390 $Y=315280
X1677 1 2 1578 397 1630 ICV_20 $T=586500 323680 0 0 $X=586310 $Y=323440
X1678 1 2 1655 399 1671 ICV_20 $T=605360 367200 0 0 $X=605170 $Y=366960
X1679 1 2 1699 400 1714 ICV_20 $T=628360 356320 1 0 $X=628170 $Y=353360
X1680 1 2 1699 415 1721 ICV_20 $T=632040 356320 0 0 $X=631850 $Y=356080
X1681 1 2 1699 412 1723 ICV_20 $T=632960 361760 0 0 $X=632770 $Y=361520
X1682 1 2 1712 412 1738 ICV_20 $T=639400 323680 1 0 $X=639210 $Y=320720
X1683 1 2 1713 399 1737 ICV_20 $T=639400 350880 0 0 $X=639210 $Y=350640
X1684 1 2 1713 414 1761 ICV_20 $T=651360 345440 0 0 $X=651170 $Y=345200
X1685 1 2 1747 414 1786 ICV_20 $T=665620 318240 1 0 $X=665430 $Y=315280
X1686 1 2 1808 398 1822 ICV_20 $T=682180 361760 0 0 $X=681990 $Y=361520
X1687 1 2 457 415 1826 ICV_20 $T=683560 372640 1 0 $X=683370 $Y=369680
X1688 1 2 1814 415 1834 ICV_20 $T=688620 334560 0 0 $X=688430 $Y=334320
X1689 1 2 1801 398 1835 ICV_20 $T=689540 323680 0 0 $X=689350 $Y=323440
X1690 1 2 1814 398 1858 ICV_20 $T=698280 345440 0 0 $X=698090 $Y=345200
X1691 1 2 1862 397 1868 ICV_20 $T=707480 367200 0 0 $X=707290 $Y=366960
X1692 1 2 1850 410 1897 ICV_20 $T=721740 329120 1 0 $X=721550 $Y=326160
X1693 1 2 467 410 470 ICV_20 $T=723580 378080 1 0 $X=723390 $Y=375120
X1694 1 2 466 415 1912 ICV_20 $T=724960 318240 0 0 $X=724770 $Y=318000
X1695 1 2 575 44 593 593 590 57 ICV_22 $T=33120 356320 1 0 $X=32930 $Y=353360
X1696 1 2 580 14 595 595 596 36 ICV_22 $T=34040 334560 0 0 $X=33850 $Y=334320
X1697 1 2 602 46 636 640 609 49 ICV_22 $T=55660 378080 1 0 $X=55470 $Y=375120
X1698 1 2 83 35 683 683 90 49 ICV_22 $T=76360 378080 1 0 $X=76170 $Y=375120
X1699 1 2 720 44 729 729 713 57 ICV_22 $T=100280 334560 0 0 $X=100090 $Y=334320
X1700 1 2 825 189 844 844 830 199 ICV_22 $T=175720 323680 0 0 $X=175530 $Y=323440
X1701 1 2 907 177 920 919 924 176 ICV_22 $T=216660 372640 1 0 $X=216470 $Y=369680
X1702 1 2 1030 172 1042 1042 1039 186 ICV_22 $T=280140 350880 1 0 $X=279950 $Y=347920
X1703 1 2 1061 172 1098 1099 1076 166 ICV_22 $T=307740 345440 1 0 $X=307550 $Y=342480
X1704 1 2 1112 266 1123 1116 1120 269 ICV_22 $T=322920 340000 0 0 $X=322730 $Y=339760
X1705 1 2 1230 266 1275 1275 1227 275 ICV_22 $T=402960 361760 0 0 $X=402770 $Y=361520
X1706 1 2 1484 399 1500 1493 1507 405 ICV_22 $T=517040 323680 0 0 $X=516850 $Y=323440
X1707 1 2 1661 412 1706 1706 1678 424 ICV_22 $T=622380 345440 1 0 $X=622190 $Y=342480
X1708 1 2 447 398 1724 1717 450 407 ICV_22 $T=631120 372640 0 0 $X=630930 $Y=372400
X1709 1 2 1720 400 1764 1764 1740 407 ICV_22 $T=651360 334560 0 0 $X=651170 $Y=334320
X1710 1 2 457 414 1847 1847 462 422 ICV_22 $T=693220 367200 0 0 $X=693030 $Y=366960
X1711 1 2 ICV_23 $T=18400 372640 1 0 $X=18210 $Y=369680
X1712 1 2 ICV_23 $T=74520 318240 1 0 $X=74330 $Y=315280
X1713 1 2 ICV_23 $T=158700 350880 1 0 $X=158510 $Y=347920
X1714 1 2 ICV_23 $T=228620 345440 0 0 $X=228430 $Y=345200
X1715 1 2 ICV_23 $T=312800 329120 0 0 $X=312610 $Y=328880
X1716 1 2 ICV_23 $T=340860 367200 0 0 $X=340670 $Y=366960
X1717 1 2 ICV_23 $T=411240 334560 1 0 $X=411050 $Y=331600
X1718 1 2 ICV_23 $T=439300 372640 1 0 $X=439110 $Y=369680
X1719 1 2 ICV_23 $T=467360 350880 1 0 $X=467170 $Y=347920
X1720 1 2 ICV_23 $T=481160 318240 0 0 $X=480970 $Y=318000
X1721 1 2 ICV_23 $T=523480 356320 1 0 $X=523290 $Y=353360
X1722 1 2 ICV_23 $T=551540 361760 1 0 $X=551350 $Y=358800
X1723 1 2 ICV_23 $T=593400 356320 0 0 $X=593210 $Y=356080
X1724 1 2 ICV_23 $T=635720 334560 1 0 $X=635530 $Y=331600
X1725 1 2 ICV_23 $T=663780 367200 1 0 $X=663590 $Y=364240
X1726 1 2 ICV_23 $T=691840 334560 1 0 $X=691650 $Y=331600
X1727 1 2 ICV_23 $T=719900 318240 1 0 $X=719710 $Y=315280
X1728 1 2 ICV_23 $T=733700 356320 0 0 $X=733510 $Y=356080
X1729 1 2 ICV_24 $T=158240 361760 1 0 $X=158050 $Y=358800
X1730 1 2 ICV_24 $T=200100 312800 0 0 $X=199910 $Y=312560
X1731 1 2 ICV_24 $T=214360 356320 1 0 $X=214170 $Y=353360
X1732 1 2 ICV_24 $T=242420 334560 1 0 $X=242230 $Y=331600
X1733 1 2 ICV_24 $T=242420 372640 1 0 $X=242230 $Y=369680
X1734 1 2 ICV_24 $T=284280 340000 0 0 $X=284090 $Y=339760
X1735 1 2 ICV_24 $T=312340 345440 0 0 $X=312150 $Y=345200
X1736 1 2 ICV_24 $T=326600 323680 1 0 $X=326410 $Y=320720
X1737 1 2 ICV_24 $T=326600 367200 1 0 $X=326410 $Y=364240
X1738 1 2 ICV_24 $T=424580 340000 0 0 $X=424390 $Y=339760
X1739 1 2 ICV_24 $T=438840 350880 1 0 $X=438650 $Y=347920
X1740 1 2 ICV_24 $T=494960 340000 1 0 $X=494770 $Y=337040
X1741 1 2 ICV_24 $T=508760 361760 0 0 $X=508570 $Y=361520
X1742 1 2 ICV_24 $T=551080 367200 1 0 $X=550890 $Y=364240
X1743 1 2 ICV_24 $T=607200 323680 1 0 $X=607010 $Y=320720
X1744 1 2 ICV_24 $T=621000 312800 0 0 $X=620810 $Y=312560
X1745 1 2 ICV_24 $T=635260 329120 1 0 $X=635070 $Y=326160
X1746 1 2 ICV_24 $T=649060 334560 0 0 $X=648870 $Y=334320
X1747 1 2 ICV_24 $T=691380 356320 1 0 $X=691190 $Y=353360
X1748 1 2 ICV_24 $T=705180 350880 0 0 $X=704990 $Y=350640
X1749 1 2 ICV_24 $T=719440 345440 1 0 $X=719250 $Y=342480
X1750 1 2 ICV_24 $T=719440 356320 1 0 $X=719250 $Y=353360
X1751 1 2 ICV_24 $T=719440 372640 1 0 $X=719250 $Y=369680
X1752 1 2 17 2 553 1 sky130_fd_sc_hd__inv_1 $T=20700 329120 1 0 $X=20510 $Y=326160
X1753 1 2 29 2 27 1 sky130_fd_sc_hd__inv_1 $T=24840 367200 0 0 $X=24650 $Y=366960
X1754 1 2 56 2 545 1 sky130_fd_sc_hd__inv_1 $T=31740 318240 0 0 $X=31550 $Y=318000
X1755 1 2 26 2 548 1 sky130_fd_sc_hd__inv_1 $T=31740 340000 0 0 $X=31550 $Y=339760
X1756 1 2 30 2 533 1 sky130_fd_sc_hd__inv_1 $T=31740 356320 1 0 $X=31550 $Y=353360
X1757 1 2 60 2 53 1 sky130_fd_sc_hd__inv_1 $T=42320 372640 1 0 $X=42130 $Y=369680
X1758 1 2 58 2 590 1 sky130_fd_sc_hd__inv_1 $T=48300 356320 1 0 $X=48110 $Y=353360
X1759 1 2 62 2 596 1 sky130_fd_sc_hd__inv_1 $T=56580 340000 1 0 $X=56390 $Y=337040
X1760 1 2 79 2 609 1 sky130_fd_sc_hd__inv_1 $T=60260 372640 0 0 $X=60070 $Y=372400
X1761 1 2 69 2 624 1 sky130_fd_sc_hd__inv_1 $T=64400 356320 1 0 $X=64210 $Y=353360
X1762 1 2 78 2 645 1 sky130_fd_sc_hd__inv_1 $T=80500 340000 1 0 $X=80310 $Y=337040
X1763 1 2 81 2 664 1 sky130_fd_sc_hd__inv_1 $T=86940 356320 1 0 $X=86750 $Y=353360
X1764 1 2 88 2 653 1 sky130_fd_sc_hd__inv_1 $T=87400 329120 0 0 $X=87210 $Y=328880
X1765 1 2 85 2 90 1 sky130_fd_sc_hd__inv_1 $T=87400 361760 0 0 $X=87210 $Y=361520
X1766 1 2 89 2 690 1 sky130_fd_sc_hd__inv_1 $T=102580 340000 1 0 $X=102390 $Y=337040
X1767 1 2 92 2 100 1 sky130_fd_sc_hd__inv_1 $T=102580 367200 1 0 $X=102390 $Y=364240
X1768 1 2 102 2 705 1 sky130_fd_sc_hd__inv_1 $T=113160 356320 0 0 $X=112970 $Y=356080
X1769 1 2 91 2 96 1 sky130_fd_sc_hd__inv_1 $T=115460 312800 0 0 $X=115270 $Y=312560
X1770 1 2 119 2 713 1 sky130_fd_sc_hd__inv_1 $T=119140 345440 1 0 $X=118950 $Y=342480
X1771 1 2 106 2 747 1 sky130_fd_sc_hd__inv_1 $T=136620 323680 1 0 $X=136430 $Y=320720
X1772 1 2 120 2 759 1 sky130_fd_sc_hd__inv_1 $T=139840 356320 1 0 $X=139650 $Y=353360
X1773 1 2 141 2 701 1 sky130_fd_sc_hd__inv_1 $T=143980 340000 1 0 $X=143790 $Y=337040
X1774 1 2 134 2 791 1 sky130_fd_sc_hd__inv_1 $T=158240 323680 1 0 $X=158050 $Y=320720
X1775 1 2 142 2 741 1 sky130_fd_sc_hd__inv_1 $T=160540 356320 1 0 $X=160350 $Y=353360
X1776 1 2 147 2 783 1 sky130_fd_sc_hd__inv_1 $T=164680 340000 1 0 $X=164490 $Y=337040
X1777 1 2 26 2 820 1 sky130_fd_sc_hd__inv_1 $T=169280 345440 1 0 $X=169090 $Y=342480
X1778 1 2 29 2 821 1 sky130_fd_sc_hd__inv_1 $T=170200 367200 0 0 $X=170010 $Y=366960
X1779 1 2 17 2 178 1 sky130_fd_sc_hd__inv_1 $T=171580 312800 0 0 $X=171390 $Y=312560
X1780 1 2 56 2 830 1 sky130_fd_sc_hd__inv_1 $T=174340 323680 0 0 $X=174150 $Y=323440
X1781 1 2 62 2 854 1 sky130_fd_sc_hd__inv_1 $T=190440 334560 0 0 $X=190250 $Y=334320
X1782 1 2 30 2 852 1 sky130_fd_sc_hd__inv_1 $T=190900 356320 1 0 $X=190710 $Y=353360
X1783 1 2 74 2 207 1 sky130_fd_sc_hd__inv_1 $T=198720 312800 0 0 $X=198530 $Y=312560
X1784 1 2 85 2 868 1 sky130_fd_sc_hd__inv_1 $T=203320 361760 1 0 $X=203130 $Y=358800
X1785 1 2 68 2 887 1 sky130_fd_sc_hd__inv_1 $T=209300 329120 1 0 $X=209110 $Y=326160
X1786 1 2 58 2 888 1 sky130_fd_sc_hd__inv_1 $T=209300 350880 1 0 $X=209110 $Y=347920
X1787 1 2 112 2 211 1 sky130_fd_sc_hd__inv_1 $T=214820 378080 1 0 $X=214630 $Y=375120
X1788 1 2 91 2 219 1 sky130_fd_sc_hd__inv_1 $T=221260 312800 0 0 $X=221070 $Y=312560
X1789 1 2 89 2 911 1 sky130_fd_sc_hd__inv_1 $T=224020 334560 1 0 $X=223830 $Y=331600
X1790 1 2 69 2 922 1 sky130_fd_sc_hd__inv_1 $T=230920 356320 1 0 $X=230730 $Y=353360
X1791 1 2 92 2 924 1 sky130_fd_sc_hd__inv_1 $T=233680 361760 1 0 $X=233490 $Y=358800
X1792 1 2 78 2 958 1 sky130_fd_sc_hd__inv_1 $T=244720 334560 1 0 $X=244530 $Y=331600
X1793 1 2 81 2 961 1 sky130_fd_sc_hd__inv_1 $T=245180 356320 0 0 $X=244990 $Y=356080
X1794 1 2 102 2 987 1 sky130_fd_sc_hd__inv_1 $T=260360 356320 0 0 $X=260170 $Y=356080
X1795 1 2 143 2 975 1 sky130_fd_sc_hd__inv_1 $T=262200 367200 0 0 $X=262010 $Y=366960
X1796 1 2 106 2 228 1 sky130_fd_sc_hd__inv_1 $T=263120 318240 1 0 $X=262930 $Y=315280
X1797 1 2 88 2 1010 1 sky130_fd_sc_hd__inv_1 $T=272780 334560 1 0 $X=272590 $Y=331600
X1798 1 2 119 2 1004 1 sky130_fd_sc_hd__inv_1 $T=272780 350880 1 0 $X=272590 $Y=347920
X1799 1 2 117 2 238 1 sky130_fd_sc_hd__inv_1 $T=278760 312800 0 0 $X=278570 $Y=312560
X1800 1 2 117 2 243 1 sky130_fd_sc_hd__inv_1 $T=279220 378080 1 0 $X=279030 $Y=375120
X1801 1 2 147 2 245 1 sky130_fd_sc_hd__inv_1 $T=286120 318240 1 0 $X=285930 $Y=315280
X1802 1 2 120 2 1039 1 sky130_fd_sc_hd__inv_1 $T=286580 350880 0 0 $X=286390 $Y=350640
X1803 1 2 162 2 1021 1 sky130_fd_sc_hd__inv_1 $T=300380 356320 0 0 $X=300190 $Y=356080
X1804 1 2 93 2 1047 1 sky130_fd_sc_hd__inv_1 $T=301760 329120 0 0 $X=301570 $Y=328880
X1805 1 2 142 2 1076 1 sky130_fd_sc_hd__inv_1 $T=303600 350880 0 0 $X=303410 $Y=350640
X1806 1 2 141 2 1083 1 sky130_fd_sc_hd__inv_1 $T=307280 334560 0 0 $X=307090 $Y=334320
X1807 1 2 134 2 254 1 sky130_fd_sc_hd__inv_1 $T=314640 318240 0 0 $X=314450 $Y=318000
X1808 1 2 132 2 1094 1 sky130_fd_sc_hd__inv_1 $T=340400 361760 1 0 $X=340210 $Y=358800
X1809 1 2 281 2 1120 1 sky130_fd_sc_hd__inv_1 $T=342700 350880 0 0 $X=342510 $Y=350640
X1810 1 2 285 2 1138 1 sky130_fd_sc_hd__inv_1 $T=353740 329120 1 0 $X=353550 $Y=326160
X1811 1 2 292 2 289 1 sky130_fd_sc_hd__inv_1 $T=355120 318240 1 0 $X=354930 $Y=315280
X1812 1 2 283 2 1158 1 sky130_fd_sc_hd__inv_1 $T=355120 367200 1 0 $X=354930 $Y=364240
X1813 1 2 297 2 1173 1 sky130_fd_sc_hd__inv_1 $T=368920 345440 0 0 $X=368730 $Y=345200
X1814 1 2 295 2 1186 1 sky130_fd_sc_hd__inv_1 $T=374900 329120 0 0 $X=374710 $Y=328880
X1815 1 2 317 2 1188 1 sky130_fd_sc_hd__inv_1 $T=381800 367200 1 0 $X=381610 $Y=364240
X1816 1 2 316 2 1223 1 sky130_fd_sc_hd__inv_1 $T=390080 334560 1 0 $X=389890 $Y=331600
X1817 1 2 310 2 319 1 sky130_fd_sc_hd__inv_1 $T=390080 378080 1 0 $X=389890 $Y=375120
X1818 1 2 330 2 1250 1 sky130_fd_sc_hd__inv_1 $T=398820 329120 0 0 $X=398630 $Y=328880
X1819 1 2 314 2 1225 1 sky130_fd_sc_hd__inv_1 $T=398820 350880 0 0 $X=398630 $Y=350640
X1820 1 2 331 2 328 1 sky130_fd_sc_hd__inv_1 $T=401120 318240 1 0 $X=400930 $Y=315280
X1821 1 2 321 2 1227 1 sky130_fd_sc_hd__inv_1 $T=411240 356320 0 0 $X=411050 $Y=356080
X1822 1 2 336 2 333 1 sky130_fd_sc_hd__inv_1 $T=413540 378080 1 0 $X=413350 $Y=375120
X1823 1 2 335 2 1256 1 sky130_fd_sc_hd__inv_1 $T=419520 345440 0 0 $X=419330 $Y=345200
X1824 1 2 340 2 1261 1 sky130_fd_sc_hd__inv_1 $T=420900 361760 1 0 $X=420710 $Y=358800
X1825 1 2 345 2 1295 1 sky130_fd_sc_hd__inv_1 $T=432400 334560 1 0 $X=432210 $Y=331600
X1826 1 2 352 2 1308 1 sky130_fd_sc_hd__inv_1 $T=441600 367200 1 0 $X=441410 $Y=364240
X1827 1 2 338 2 349 1 sky130_fd_sc_hd__inv_1 $T=442520 312800 0 0 $X=442330 $Y=312560
X1828 1 2 348 2 1313 1 sky130_fd_sc_hd__inv_1 $T=442980 345440 0 0 $X=442790 $Y=345200
X1829 1 2 353 2 1350 1 sky130_fd_sc_hd__inv_1 $T=449880 334560 1 0 $X=449690 $Y=331600
X1830 1 2 363 2 1356 1 sky130_fd_sc_hd__inv_1 $T=462760 356320 1 0 $X=462570 $Y=353360
X1831 1 2 355 2 1342 1 sky130_fd_sc_hd__inv_1 $T=463680 367200 0 0 $X=463490 $Y=366960
X1832 1 2 375 2 1400 1 sky130_fd_sc_hd__inv_1 $T=481160 361760 0 0 $X=480970 $Y=361520
X1833 1 2 373 2 371 1 sky130_fd_sc_hd__inv_1 $T=483000 318240 0 0 $X=482810 $Y=318000
X1834 1 2 364 2 1391 1 sky130_fd_sc_hd__inv_1 $T=487140 372640 0 0 $X=486950 $Y=372400
X1835 1 2 379 2 1456 1 sky130_fd_sc_hd__inv_1 $T=508760 361760 1 0 $X=508570 $Y=358800
X1836 1 2 388 2 381 1 sky130_fd_sc_hd__inv_1 $T=511060 312800 0 0 $X=510870 $Y=312560
X1837 1 2 389 2 1434 1 sky130_fd_sc_hd__inv_1 $T=511060 372640 0 0 $X=510870 $Y=372400
X1838 1 2 386 2 1457 1 sky130_fd_sc_hd__inv_1 $T=515200 345440 0 0 $X=515010 $Y=345200
X1839 1 2 385 2 1450 1 sky130_fd_sc_hd__inv_1 $T=517040 340000 1 0 $X=516850 $Y=337040
X1840 1 2 310 2 1506 1 sky130_fd_sc_hd__inv_1 $T=527160 340000 1 0 $X=526970 $Y=337040
X1841 1 2 292 2 1507 1 sky130_fd_sc_hd__inv_1 $T=530840 318240 1 0 $X=530650 $Y=315280
X1842 1 2 288 2 1503 1 sky130_fd_sc_hd__inv_1 $T=530840 350880 1 0 $X=530650 $Y=347920
X1843 1 2 321 2 1509 1 sky130_fd_sc_hd__inv_1 $T=531300 356320 0 0 $X=531110 $Y=356080
X1844 1 2 336 2 426 1 sky130_fd_sc_hd__inv_1 $T=544640 372640 0 0 $X=544450 $Y=372400
X1845 1 2 285 2 1542 1 sky130_fd_sc_hd__inv_1 $T=553380 334560 1 0 $X=553190 $Y=331600
X1846 1 2 314 2 1543 1 sky130_fd_sc_hd__inv_1 $T=553380 350880 1 0 $X=553190 $Y=347920
X1847 1 2 317 2 1557 1 sky130_fd_sc_hd__inv_1 $T=564880 361760 1 0 $X=564690 $Y=358800
X1848 1 2 330 2 1580 1 sky130_fd_sc_hd__inv_1 $T=571780 329120 0 0 $X=571590 $Y=328880
X1849 1 2 297 2 1585 1 sky130_fd_sc_hd__inv_1 $T=572700 350880 0 0 $X=572510 $Y=350640
X1850 1 2 392 2 1599 1 sky130_fd_sc_hd__inv_1 $T=577300 323680 1 0 $X=577110 $Y=320720
X1851 1 2 283 2 1604 1 sky130_fd_sc_hd__inv_1 $T=579600 367200 1 0 $X=579410 $Y=364240
X1852 1 2 271 2 437 1 sky130_fd_sc_hd__inv_1 $T=593860 378080 1 0 $X=593670 $Y=375120
X1853 1 2 353 2 1633 1 sky130_fd_sc_hd__inv_1 $T=595240 334560 0 0 $X=595050 $Y=334320
X1854 1 2 335 2 1665 1 sky130_fd_sc_hd__inv_1 $T=612720 356320 0 0 $X=612530 $Y=356080
X1855 1 2 352 2 1668 1 sky130_fd_sc_hd__inv_1 $T=613180 367200 0 0 $X=612990 $Y=366960
X1856 1 2 286 2 1678 1 sky130_fd_sc_hd__inv_1 $T=618700 345440 0 0 $X=618510 $Y=345200
X1857 1 2 340 2 1694 1 sky130_fd_sc_hd__inv_1 $T=625140 361760 1 0 $X=624950 $Y=358800
X1858 1 2 338 2 445 1 sky130_fd_sc_hd__inv_1 $T=626060 318240 1 0 $X=625870 $Y=315280
X1859 1 2 295 2 1719 1 sky130_fd_sc_hd__inv_1 $T=637560 329120 0 0 $X=637370 $Y=328880
X1860 1 2 348 2 1722 1 sky130_fd_sc_hd__inv_1 $T=639400 345440 1 0 $X=639210 $Y=342480
X1861 1 2 345 2 1740 1 sky130_fd_sc_hd__inv_1 $T=647680 334560 0 0 $X=647490 $Y=334320
X1862 1 2 331 2 1749 1 sky130_fd_sc_hd__inv_1 $T=653660 323680 1 0 $X=653470 $Y=320720
X1863 1 2 374 2 1781 1 sky130_fd_sc_hd__inv_1 $T=667460 334560 1 0 $X=667270 $Y=331600
X1864 1 2 354 2 456 1 sky130_fd_sc_hd__inv_1 $T=677580 318240 0 0 $X=677390 $Y=318000
X1865 1 2 366 2 1797 1 sky130_fd_sc_hd__inv_1 $T=678960 345440 1 0 $X=678770 $Y=342480
X1866 1 2 363 2 1780 1 sky130_fd_sc_hd__inv_1 $T=679880 361760 1 0 $X=679690 $Y=358800
X1867 1 2 355 2 1818 1 sky130_fd_sc_hd__inv_1 $T=686320 367200 1 0 $X=686130 $Y=364240
X1868 1 2 385 2 1827 1 sky130_fd_sc_hd__inv_1 $T=691380 340000 1 0 $X=691190 $Y=337040
X1869 1 2 364 2 468 1 sky130_fd_sc_hd__inv_1 $T=708860 378080 1 0 $X=708670 $Y=375120
X1870 1 2 388 2 1869 1 sky130_fd_sc_hd__inv_1 $T=714840 318240 0 0 $X=714650 $Y=318000
X1871 1 2 386 2 1891 1 sky130_fd_sc_hd__inv_1 $T=718060 345440 1 0 $X=717870 $Y=342480
X1872 1 2 379 2 1871 1 sky130_fd_sc_hd__inv_1 $T=718980 356320 0 0 $X=718790 $Y=356080
X1873 1 2 380 2 1889 1 sky130_fd_sc_hd__inv_1 $T=721740 334560 1 0 $X=721550 $Y=331600
X1874 1 2 ICV_25 $T=16560 367200 1 0 $X=16370 $Y=364240
X1875 1 2 ICV_25 $T=30360 356320 0 0 $X=30170 $Y=356080
X1876 1 2 ICV_25 $T=44620 318240 1 0 $X=44430 $Y=315280
X1877 1 2 ICV_25 $T=114540 356320 0 0 $X=114350 $Y=356080
X1878 1 2 ICV_25 $T=142600 350880 0 0 $X=142410 $Y=350640
X1879 1 2 ICV_25 $T=170660 356320 0 0 $X=170470 $Y=356080
X1880 1 2 ICV_25 $T=310960 356320 0 0 $X=310770 $Y=356080
X1881 1 2 ICV_25 $T=339020 345440 0 0 $X=338830 $Y=345200
X1882 1 2 ICV_25 $T=381340 372640 1 0 $X=381150 $Y=369680
X1883 1 2 ICV_25 $T=409400 356320 1 0 $X=409210 $Y=353360
X1884 1 2 ICV_25 $T=409400 378080 1 0 $X=409210 $Y=375120
X1885 1 2 ICV_25 $T=437460 340000 1 0 $X=437270 $Y=337040
X1886 1 2 ICV_25 $T=451260 372640 0 0 $X=451070 $Y=372400
X1887 1 2 ICV_25 $T=535440 367200 0 0 $X=535250 $Y=366960
X1888 1 2 ICV_25 $T=535440 372640 0 0 $X=535250 $Y=372400
X1889 1 2 ICV_25 $T=577760 334560 1 0 $X=577570 $Y=331600
X1890 1 2 ICV_25 $T=605820 340000 1 0 $X=605630 $Y=337040
X1891 1 2 ICV_25 $T=605820 350880 1 0 $X=605630 $Y=347920
X1892 1 2 ICV_25 $T=661940 340000 1 0 $X=661750 $Y=337040
X1893 1 2 ICV_25 $T=661940 378080 1 0 $X=661750 $Y=375120
X1894 1 2 ICV_25 $T=718060 323680 1 0 $X=717870 $Y=320720
X1895 1 2 569 548 54 ICV_26 $T=28060 340000 1 0 $X=27870 $Y=337040
X1896 1 2 623 72 54 ICV_26 $T=57040 318240 0 0 $X=56850 $Y=318000
X1897 1 2 642 645 57 ICV_26 $T=66240 340000 0 0 $X=66050 $Y=339760
X1898 1 2 86 87 52 ICV_26 $T=74520 312800 0 0 $X=74330 $Y=312560
X1899 1 2 700 699 52 ICV_26 $T=94300 334560 1 0 $X=94110 $Y=331600
X1900 1 2 739 741 39 ICV_26 $T=115920 356320 1 0 $X=115730 $Y=353360
X1901 1 2 774 701 34 ICV_26 $T=138000 323680 1 0 $X=137810 $Y=320720
X1902 1 2 182 178 184 ICV_26 $T=174340 312800 0 0 $X=174150 $Y=312560
X1903 1 2 836 820 186 ICV_26 $T=174340 340000 0 0 $X=174150 $Y=339760
X1904 1 2 870 854 184 ICV_26 $T=199180 323680 1 0 $X=198990 $Y=320720
X1905 1 2 921 922 197 ICV_26 $T=225400 334560 0 0 $X=225210 $Y=334320
X1906 1 2 931 922 201 ICV_26 $T=230000 350880 1 0 $X=229810 $Y=347920
X1907 1 2 954 961 166 ICV_26 $T=244720 340000 0 0 $X=244530 $Y=339760
X1908 1 2 972 975 185 ICV_26 $T=252540 367200 0 0 $X=252350 $Y=366960
X1909 1 2 979 228 198 ICV_26 $T=256220 323680 1 0 $X=256030 $Y=320720
X1910 1 2 1043 239 188 ICV_26 $T=290720 361760 0 0 $X=290530 $Y=361520
X1911 1 2 1058 1039 201 ICV_26 $T=294860 356320 1 0 $X=294670 $Y=353360
X1912 1 2 1060 1047 186 ICV_26 $T=296240 334560 0 0 $X=296050 $Y=334320
X1913 1 2 1080 243 185 ICV_26 $T=306820 372640 0 0 $X=306630 $Y=372400
X1914 1 2 1086 1083 198 ICV_26 $T=309580 340000 0 0 $X=309390 $Y=339760
X1915 1 2 1321 1295 269 ICV_26 $T=436080 318240 1 0 $X=435890 $Y=315280
X1916 1 2 1337 1313 280 ICV_26 $T=445740 340000 0 0 $X=445550 $Y=339760
X1917 1 2 1353 1356 296 ICV_26 $T=449880 350880 0 0 $X=449690 $Y=350640
X1918 1 2 1417 1382 267 ICV_26 $T=483000 329120 0 0 $X=482810 $Y=328880
X1919 1 2 1475 1450 275 ICV_26 $T=511060 334560 0 0 $X=510870 $Y=334320
X1920 1 2 1514 1503 418 ICV_26 $T=534060 345440 0 0 $X=533870 $Y=345200
X1921 1 2 1537 1542 407 ICV_26 $T=548320 323680 1 0 $X=548130 $Y=320720
X1922 1 2 1554 426 407 ICV_26 $T=554760 372640 0 0 $X=554570 $Y=372400
X1923 1 2 1586 1580 409 ICV_26 $T=572700 323680 1 0 $X=572510 $Y=320720
X1924 1 2 1631 1633 408 ICV_26 $T=595240 329120 0 0 $X=595050 $Y=328880
X1925 1 2 1716 1694 409 ICV_26 $T=637560 361760 1 0 $X=637370 $Y=358800
X1926 1 2 1796 455 424 ICV_26 $T=675280 378080 1 0 $X=675090 $Y=375120
X1927 1 2 1886 1891 422 ICV_26 $T=716680 350880 1 0 $X=716490 $Y=347920
X1928 1 2 591 43 635 68 72 ICV_27 $T=55660 329120 1 0 $X=55470 $Y=326160
X1929 1 2 687 42 722 93 699 ICV_27 $T=97520 329120 0 0 $X=97330 $Y=328880
X1930 1 2 118 44 771 117 126 ICV_27 $T=132480 318240 1 0 $X=132290 $Y=315280
X1931 1 2 859 177 881 60 205 ICV_27 $T=195960 372640 1 0 $X=195770 $Y=369680
X1932 1 2 1022 175 1043 141 239 ICV_27 $T=283820 361760 1 0 $X=283630 $Y=358800
X1933 1 2 1112 257 1163 286 1131 ICV_27 $T=345000 340000 0 0 $X=344810 $Y=339760
X1934 1 2 309 273 322 324 315 ICV_27 $T=378120 312800 0 0 $X=377930 $Y=312560
X1935 1 2 343 260 1332 350 1306 ICV_27 $T=433780 372640 0 0 $X=433590 $Y=372400
X1936 1 2 356 265 362 354 360 ICV_27 $T=454940 312800 0 0 $X=454750 $Y=312560
X1937 1 2 1360 260 1408 366 1371 ICV_27 $T=471500 340000 0 0 $X=471310 $Y=339760
X1938 1 2 1378 260 1417 374 1382 ICV_27 $T=477940 334560 1 0 $X=477750 $Y=331600
X1939 1 2 1430 266 1481 380 1425 ICV_27 $T=506460 329120 1 0 $X=506270 $Y=326160
X1940 1 2 1612 397 1626 281 1616 ICV_27 $T=585580 350880 0 0 $X=585390 $Y=350640
X1941 1 2 1663 415 1679 316 1682 ICV_27 $T=611800 334560 1 0 $X=611610 $Y=331600
X1942 1 2 1640 414 1680 419 439 ICV_27 $T=612260 312800 0 0 $X=612070 $Y=312560
X1943 1 2 1862 398 1887 375 1881 ICV_27 $T=710700 372640 1 0 $X=710510 $Y=369680
X1944 1 2 466 414 1888 373 469 ICV_27 $T=711160 318240 1 0 $X=710970 $Y=315280
X1945 1 2 525 13 546 ICV_28 $T=6900 345440 1 0 $X=6710 $Y=342480
X1946 1 2 9 20 32 ICV_28 $T=6900 378080 1 0 $X=6710 $Y=375120
X1947 1 2 608 43 630 ICV_28 $T=51980 361760 0 0 $X=51790 $Y=361520
X1948 1 2 644 18 658 ICV_28 $T=65780 356320 1 0 $X=65590 $Y=353360
X1949 1 2 637 44 677 ICV_28 $T=76360 323680 1 0 $X=76170 $Y=320720
X1950 1 2 720 18 749 ICV_28 $T=111780 334560 1 0 $X=111590 $Y=331600
X1951 1 2 720 13 743 ICV_28 $T=111780 340000 1 0 $X=111590 $Y=337040
X1952 1 2 785 15 739 ICV_28 $T=141220 356320 1 0 $X=141030 $Y=353360
X1953 1 2 785 43 803 ICV_28 $T=144900 361760 1 0 $X=144710 $Y=358800
X1954 1 2 826 172 836 ICV_28 $T=166060 340000 1 0 $X=165870 $Y=337040
X1955 1 2 884 187 893 ICV_28 $T=204240 334560 1 0 $X=204050 $Y=331600
X1956 1 2 884 170 896 ICV_28 $T=204700 340000 1 0 $X=204510 $Y=337040
X1957 1 2 859 163 863 ICV_28 $T=204700 372640 1 0 $X=204510 $Y=369680
X1958 1 2 913 172 930 ICV_28 $T=220800 350880 1 0 $X=220610 $Y=347920
X1959 1 2 218 170 947 ICV_28 $T=230460 312800 0 0 $X=230270 $Y=312560
X1960 1 2 963 175 973 ICV_28 $T=244720 367200 1 0 $X=244530 $Y=364240
X1961 1 2 963 156 974 ICV_28 $T=244720 372640 1 0 $X=244530 $Y=369680
X1962 1 2 250 187 1096 ICV_28 $T=308200 318240 1 0 $X=308010 $Y=315280
X1963 1 2 1112 260 1145 ICV_28 $T=333040 340000 1 0 $X=332850 $Y=337040
X1964 1 2 1118 253 1161 ICV_28 $T=342700 329120 0 0 $X=342510 $Y=328880
X1965 1 2 1171 253 1190 ICV_28 $T=361100 329120 1 0 $X=360910 $Y=326160
X1966 1 2 312 273 1211 ICV_28 $T=372140 372640 1 0 $X=371950 $Y=369680
X1967 1 2 1203 264 1217 ICV_28 $T=376280 329120 0 0 $X=376090 $Y=328880
X1968 1 2 1203 257 1236 ICV_28 $T=385020 329120 1 0 $X=384830 $Y=326160
X1969 1 2 1230 257 1247 ICV_28 $T=389160 367200 1 0 $X=388970 $Y=364240
X1970 1 2 1257 257 1259 ICV_28 $T=400200 350880 0 0 $X=400010 $Y=350640
X1971 1 2 1230 253 1274 ICV_28 $T=403420 361760 1 0 $X=403230 $Y=358800
X1972 1 2 1331 257 1346 ICV_28 $T=441140 329120 1 0 $X=440950 $Y=326160
X1973 1 2 1384 257 1406 ICV_28 $T=469200 350880 1 0 $X=469010 $Y=347920
X1974 1 2 1430 273 1445 ICV_28 $T=487140 323680 0 0 $X=486950 $Y=323440
X1975 1 2 1661 397 1708 ICV_28 $T=623300 345440 0 0 $X=623110 $Y=345200
X1976 1 2 1775 414 1836 ICV_28 $T=689080 329120 0 0 $X=688890 $Y=328880
X1977 1 2 1861 414 1886 ICV_28 $T=708860 345440 1 0 $X=708670 $Y=342480
X1978 1 2 48 46 571 ICV_29 $T=23920 372640 0 0 $X=23730 $Y=372400
X1979 1 2 575 42 601 ICV_29 $T=35420 361760 1 0 $X=35230 $Y=358800
X1980 1 2 83 20 669 ICV_29 $T=69460 372640 0 0 $X=69270 $Y=372400
X1981 1 2 786 13 817 ICV_29 $T=153640 340000 0 0 $X=153450 $Y=339760
X1982 1 2 825 168 831 ICV_29 $T=163760 318240 0 0 $X=163570 $Y=318000
X1983 1 2 853 190 865 ICV_29 $T=189520 323680 0 0 $X=189330 $Y=323440
X1984 1 2 223 187 227 ICV_29 $T=248400 312800 0 0 $X=248210 $Y=312560
X1985 1 2 1073 187 1088 ICV_29 $T=303140 329120 0 0 $X=302950 $Y=328880
X1986 1 2 1095 257 1103 ICV_29 $T=312340 378080 1 0 $X=312150 $Y=375120
X1987 1 2 1102 264 1150 ICV_29 $T=336260 345440 1 0 $X=336070 $Y=342480
X1988 1 2 325 266 1239 ICV_29 $T=386860 312800 0 0 $X=386670 $Y=312560
X1989 1 2 1339 262 1358 ICV_29 $T=444360 345440 0 0 $X=444170 $Y=345200
X1990 1 2 377 262 1440 ICV_29 $T=485300 378080 1 0 $X=485110 $Y=375120
X1991 1 2 1485 397 1494 ICV_29 $T=515200 329120 1 0 $X=515010 $Y=326160
X1992 1 2 1529 412 1548 ICV_29 $T=543260 329120 1 0 $X=543070 $Y=326160
X1993 1 2 1527 397 1573 ICV_29 $T=554760 350880 1 0 $X=554570 $Y=347920
X1994 1 2 1574 398 1611 ICV_29 $T=574540 334560 0 0 $X=574350 $Y=334320
X1995 1 2 1612 415 1643 ICV_29 $T=592480 356320 1 0 $X=592290 $Y=353360
X1996 1 2 1618 410 1653 ICV_29 $T=596620 334560 0 0 $X=596430 $Y=334320
X1997 1 2 1661 398 1685 ICV_29 $T=612260 340000 0 0 $X=612070 $Y=339760
X1998 1 2 1652 397 1688 ICV_29 $T=613640 361760 1 0 $X=613450 $Y=358800
X1999 1 2 447 400 1717 ICV_29 $T=627440 367200 0 0 $X=627250 $Y=366960
X2000 1 2 1779 397 1792 ICV_29 $T=665620 340000 1 0 $X=665430 $Y=337040
X2001 1 2 454 412 1796 ICV_29 $T=665620 378080 1 0 $X=665430 $Y=375120
X2002 1 2 1775 412 1820 ICV_29 $T=679420 329120 0 0 $X=679230 $Y=328880
X2003 1 2 1808 412 1824 ICV_29 $T=681260 361760 1 0 $X=681070 $Y=358800
X2004 1 2 457 399 1830 ICV_29 $T=683560 367200 0 0 $X=683370 $Y=366960
X2005 1 2 1814 412 1857 ICV_29 $T=696440 334560 0 0 $X=696250 $Y=334320
X2006 1 2 532 533 28 542 533 34 ICV_30 $T=10580 356320 1 0 $X=10390 $Y=353360
X2007 1 2 546 548 34 551 548 28 ICV_30 $T=15640 340000 0 0 $X=15450 $Y=339760
X2008 1 2 552 545 28 557 553 28 ICV_30 $T=20240 323680 1 0 $X=20050 $Y=320720
X2009 1 2 554 27 47 556 27 55 ICV_30 $T=23000 361760 0 0 $X=22810 $Y=361520
X2010 1 2 578 53 55 582 53 38 ICV_30 $T=37720 367200 1 0 $X=37530 $Y=364240
X2011 1 2 600 596 52 612 596 37 ICV_30 $T=48300 340000 1 0 $X=48110 $Y=337040
X2012 1 2 607 609 75 614 609 63 ICV_30 $T=48760 372640 1 0 $X=48570 $Y=369680
X2013 1 2 622 624 36 628 624 28 ICV_30 $T=59340 350880 1 0 $X=59150 $Y=347920
X2014 1 2 635 72 52 632 72 39 ICV_30 $T=62100 323680 0 0 $X=61910 $Y=323440
X2015 1 2 633 624 57 638 624 39 ICV_30 $T=62100 356320 0 0 $X=61910 $Y=356080
X2016 1 2 643 645 52 651 653 39 ICV_30 $T=67620 334560 1 0 $X=67430 $Y=331600
X2017 1 2 656 87 37 657 87 39 ICV_30 $T=76360 318240 1 0 $X=76170 $Y=315280
X2018 1 2 678 664 36 688 690 52 ICV_30 $T=83720 350880 1 0 $X=83530 $Y=347920
X2019 1 2 695 96 37 696 699 28 ICV_30 $T=90160 318240 0 0 $X=89970 $Y=318000
X2020 1 2 685 664 39 703 705 28 ICV_30 $T=92000 350880 1 0 $X=91810 $Y=347920
X2021 1 2 692 690 37 708 690 39 ICV_30 $T=94300 340000 1 0 $X=94110 $Y=337040
X2022 1 2 717 100 47 716 100 38 ICV_30 $T=103040 367200 0 0 $X=102850 $Y=366960
X2023 1 2 724 713 52 730 713 54 ICV_30 $T=104880 340000 0 0 $X=104690 $Y=339760
X2024 1 2 725 705 36 706 705 39 ICV_30 $T=105800 350880 1 0 $X=105610 $Y=347920
X2025 1 2 746 747 54 751 747 36 ICV_30 $T=119140 329120 0 0 $X=118950 $Y=328880
X2026 1 2 768 126 37 771 126 57 ICV_30 $T=132940 312800 0 0 $X=132750 $Y=312560
X2027 1 2 770 759 34 777 759 52 ICV_30 $T=134320 350880 0 0 $X=134130 $Y=350640
X2028 1 2 797 741 57 807 741 54 ICV_30 $T=151800 356320 1 0 $X=151610 $Y=353360
X2029 1 2 153 155 34 811 791 34 ICV_30 $T=154100 312800 0 0 $X=153910 $Y=312560
X2030 1 2 837 821 188 839 821 194 ICV_30 $T=175260 367200 0 0 $X=175070 $Y=366960
X2031 1 2 838 821 193 828 821 185 ICV_30 $T=176640 372640 0 0 $X=176450 $Y=372400
X2032 1 2 857 205 188 860 205 193 ICV_30 $T=192740 372640 0 0 $X=192550 $Y=372400
X2033 1 2 869 854 199 864 854 198 ICV_30 $T=202400 318240 0 0 $X=202210 $Y=318000
X2034 1 2 905 887 186 904 887 179 ICV_30 $T=218500 318240 1 0 $X=218310 $Y=315280
X2035 1 2 215 211 193 915 211 188 ICV_30 $T=218500 372640 0 0 $X=218310 $Y=372400
X2036 1 2 912 887 201 916 887 198 ICV_30 $T=219420 329120 1 0 $X=219230 $Y=326160
X2037 1 2 926 219 199 928 911 166 ICV_30 $T=228620 318240 1 0 $X=228430 $Y=315280
X2038 1 2 925 922 199 932 922 198 ICV_30 $T=230460 345440 0 0 $X=230270 $Y=345200
X2039 1 2 929 911 201 936 911 186 ICV_30 $T=230920 329120 1 0 $X=230730 $Y=326160
X2040 1 2 943 924 194 949 211 180 ICV_30 $T=237820 372640 0 0 $X=237630 $Y=372400
X2041 1 2 955 961 186 952 961 198 ICV_30 $T=244720 345440 1 0 $X=244530 $Y=342480
X2042 1 2 978 228 199 232 217 198 ICV_30 $T=258520 318240 0 0 $X=258330 $Y=318000
X2043 1 2 237 238 197 1012 238 179 ICV_30 $T=269100 312800 0 0 $X=268910 $Y=312560
X2044 1 2 1009 230 194 1018 239 193 ICV_30 $T=270480 372640 0 0 $X=270290 $Y=372400
X2045 1 2 1015 239 194 1020 1021 188 ICV_30 $T=272780 361760 1 0 $X=272590 $Y=358800
X2046 1 2 1006 1010 179 1013 1010 198 ICV_30 $T=274620 329120 0 0 $X=274430 $Y=328880
X2047 1 2 1017 1004 166 1026 1004 197 ICV_30 $T=276000 340000 0 0 $X=275810 $Y=339760
X2048 1 2 1040 1039 184 1048 1039 166 ICV_30 $T=287960 334560 0 0 $X=287770 $Y=334320
X2049 1 2 1046 1047 201 1050 1047 184 ICV_30 $T=291640 329120 1 0 $X=291450 $Y=326160
X2050 1 2 1066 245 186 249 245 199 ICV_30 $T=299920 312800 0 0 $X=299730 $Y=312560
X2051 1 2 1092 1094 194 1103 261 268 ICV_30 $T=318320 372640 1 0 $X=318130 $Y=369680
X2052 1 2 287 284 263 1160 1158 277 ICV_30 $T=345920 372640 1 0 $X=345730 $Y=369680
X2053 1 2 1143 289 280 1144 289 275 ICV_30 $T=346380 318240 1 0 $X=346190 $Y=315280
X2054 1 2 1133 1138 277 1161 1138 263 ICV_30 $T=347760 334560 1 0 $X=347570 $Y=331600
X2055 1 2 1170 1158 268 1178 1158 296 ICV_30 $T=356500 361760 0 0 $X=356310 $Y=361520
X2056 1 2 1172 1173 296 1179 1173 268 ICV_30 $T=357880 345440 1 0 $X=357690 $Y=342480
X2057 1 2 1182 1186 267 1197 1186 275 ICV_30 $T=370760 323680 0 0 $X=370570 $Y=323440
X2058 1 2 1201 315 275 1208 315 296 ICV_30 $T=375360 323680 1 0 $X=375170 $Y=320720
X2059 1 2 1217 1223 296 1156 289 263 ICV_30 $T=385480 323680 1 0 $X=385290 $Y=320720
X2060 1 2 1215 1225 263 1238 1225 296 ICV_30 $T=390080 345440 0 0 $X=389890 $Y=345200
X2061 1 2 1232 1223 280 1241 1223 277 ICV_30 $T=391460 334560 1 0 $X=391270 $Y=331600
X2062 1 2 332 333 269 334 333 280 ICV_30 $T=401120 378080 1 0 $X=400930 $Y=375120
X2063 1 2 1263 333 263 337 333 296 ICV_30 $T=410320 372640 0 0 $X=410130 $Y=372400
X2064 1 2 1269 1261 267 1273 1261 263 ICV_30 $T=413080 356320 1 0 $X=412890 $Y=353360
X2065 1 2 1277 1250 268 1283 1250 277 ICV_30 $T=414000 334560 1 0 $X=413810 $Y=331600
X2066 1 2 1302 1306 268 1309 1306 277 ICV_30 $T=427340 367200 1 0 $X=427150 $Y=364240
X2067 1 2 1307 1308 296 1312 1308 263 ICV_30 $T=428260 361760 0 0 $X=428070 $Y=361520
X2068 1 2 1348 1342 268 1359 1356 275 ICV_30 $T=449420 361760 1 0 $X=449230 $Y=358800
X2069 1 2 1355 360 268 1352 360 296 ICV_30 $T=450800 323680 1 0 $X=450610 $Y=320720
X2070 1 2 1361 1356 267 1341 1308 277 ICV_30 $T=454940 356320 0 0 $X=454750 $Y=356080
X2071 1 2 1362 1342 280 1370 1342 267 ICV_30 $T=455400 367200 0 0 $X=455210 $Y=366960
X2072 1 2 1354 1342 277 1374 1342 296 ICV_30 $T=457700 361760 1 0 $X=457510 $Y=358800
X2073 1 2 1389 1391 269 1394 1400 269 ICV_30 $T=469200 361760 1 0 $X=469010 $Y=358800
X2074 1 2 1398 1400 277 1410 1400 296 ICV_30 $T=473800 356320 0 0 $X=473610 $Y=356080
X2075 1 2 1399 1391 267 1404 1391 280 ICV_30 $T=474260 367200 0 0 $X=474070 $Y=366960
X2076 1 2 1432 1434 296 1453 1456 269 ICV_30 $T=492200 361760 0 0 $X=492010 $Y=361520
X2077 1 2 1438 1450 269 1436 1457 280 ICV_30 $T=495420 340000 0 0 $X=495230 $Y=339760
X2078 1 2 1445 1425 280 1444 1425 269 ICV_30 $T=497260 323680 1 0 $X=497070 $Y=320720
X2079 1 2 1424 1391 263 1421 1391 296 ICV_30 $T=500480 361760 0 0 $X=500290 $Y=361520
X2080 1 2 1467 381 268 1463 1425 268 ICV_30 $T=511060 318240 0 0 $X=510870 $Y=318000
X2081 1 2 1469 1450 277 1468 1425 277 ICV_30 $T=511060 329120 0 0 $X=510870 $Y=328880
X2082 1 2 1473 1456 277 1479 1457 263 ICV_30 $T=511060 356320 0 0 $X=510870 $Y=356080
X2083 1 2 1505 406 408 413 406 405 ICV_30 $T=528080 312800 0 0 $X=527890 $Y=312560
X2084 1 2 1545 430 408 1552 430 424 ICV_30 $T=549700 312800 0 0 $X=549510 $Y=312560
X2085 1 2 1550 1543 418 1556 1557 424 ICV_30 $T=552000 350880 0 0 $X=551810 $Y=350640
X2086 1 2 1587 1580 408 1588 1580 417 ICV_30 $T=573160 329120 0 0 $X=572970 $Y=328880
X2087 1 2 1626 1616 409 1625 1616 405 ICV_30 $T=595240 350880 0 0 $X=595050 $Y=350640
X2088 1 2 1638 1604 408 1644 1604 417 ICV_30 $T=597080 367200 0 0 $X=596890 $Y=366960
X2089 1 2 1632 1633 409 1654 1633 424 ICV_30 $T=600760 334560 1 0 $X=600570 $Y=331600
X2090 1 2 1662 1665 417 1645 1633 418 ICV_30 $T=610420 345440 0 0 $X=610230 $Y=345200
X2091 1 2 1672 439 424 1681 439 407 ICV_30 $T=614560 318240 0 0 $X=614370 $Y=318000
X2092 1 2 1673 1668 424 1671 1668 408 ICV_30 $T=614560 367200 0 0 $X=614370 $Y=366960
X2093 1 2 1684 1665 422 1696 1665 407 ICV_30 $T=623300 350880 0 0 $X=623110 $Y=350640
X2094 1 2 1686 1665 408 1688 1665 409 ICV_30 $T=623760 356320 0 0 $X=623570 $Y=356080
X2095 1 2 1714 1694 407 1721 1694 418 ICV_30 $T=637560 356320 1 0 $X=637370 $Y=353360
X2096 1 2 449 450 408 1731 450 418 ICV_30 $T=640780 378080 1 0 $X=640590 $Y=375120
X2097 1 2 1743 1694 422 1745 1694 417 ICV_30 $T=651360 356320 0 0 $X=651170 $Y=356080
X2098 1 2 1744 1694 408 1746 1694 405 ICV_30 $T=651360 361760 0 0 $X=651170 $Y=361520
X2099 1 2 1750 1740 409 1758 1722 405 ICV_30 $T=654120 345440 1 0 $X=653930 $Y=342480
X2100 1 2 1766 1740 424 1755 1740 408 ICV_30 $T=665160 334560 0 0 $X=664970 $Y=334320
X2101 1 2 1771 1780 418 1774 1722 418 ICV_30 $T=666540 350880 0 0 $X=666350 $Y=350640
X2102 1 2 1778 1780 409 1783 455 417 ICV_30 $T=666540 367200 1 0 $X=666350 $Y=364240
X2103 1 2 1821 1818 407 1824 1818 424 ICV_30 $T=687700 356320 0 0 $X=687510 $Y=356080
X2104 1 2 1831 456 408 1837 456 407 ICV_30 $T=693680 318240 0 0 $X=693490 $Y=318000
X2105 1 2 1830 462 408 1825 462 417 ICV_30 $T=693680 367200 1 0 $X=693490 $Y=364240
X2106 1 2 1868 1881 409 1887 1881 405 ICV_30 $T=716220 367200 0 0 $X=716030 $Y=366960
X2107 1 2 16 19 2 21 1 sky130_fd_sc_hd__and2_1 $T=8280 312800 0 0 $X=8090 $Y=312560
X2108 1 2 17 19 2 529 1 sky130_fd_sc_hd__and2_1 $T=8280 329120 0 0 $X=8090 $Y=328880
X2109 1 2 26 19 2 527 1 sky130_fd_sc_hd__and2_1 $T=13340 340000 0 0 $X=13150 $Y=339760
X2110 1 2 29 31 2 528 1 sky130_fd_sc_hd__and2_1 $T=14260 367200 1 0 $X=14070 $Y=364240
X2111 1 2 30 19 2 530 1 sky130_fd_sc_hd__and2_1 $T=15180 356320 0 0 $X=14990 $Y=356080
X2112 1 2 56 19 2 559 1 sky130_fd_sc_hd__and2_1 $T=30820 323680 0 0 $X=30630 $Y=323440
X2113 1 2 58 19 2 573 1 sky130_fd_sc_hd__and2_1 $T=31280 361760 0 0 $X=31090 $Y=361520
X2114 1 2 62 19 2 576 1 sky130_fd_sc_hd__and2_1 $T=34040 340000 0 0 $X=33850 $Y=339760
X2115 1 2 60 31 2 577 1 sky130_fd_sc_hd__and2_1 $T=34040 367200 0 0 $X=33850 $Y=366960
X2116 1 2 68 19 2 603 1 sky130_fd_sc_hd__and2_1 $T=45540 329120 1 0 $X=45350 $Y=326160
X2117 1 2 69 19 2 604 1 sky130_fd_sc_hd__and2_1 $T=45540 361760 1 0 $X=45350 $Y=358800
X2118 1 2 74 19 2 610 1 sky130_fd_sc_hd__and2_1 $T=51980 312800 0 0 $X=51790 $Y=312560
X2119 1 2 78 19 2 626 1 sky130_fd_sc_hd__and2_1 $T=57960 340000 1 0 $X=57770 $Y=337040
X2120 1 2 81 19 2 646 1 sky130_fd_sc_hd__and2_1 $T=66240 361760 1 0 $X=66050 $Y=358800
X2121 1 2 79 31 2 625 1 sky130_fd_sc_hd__and2_1 $T=66240 361760 0 0 $X=66050 $Y=361520
X2122 1 2 85 31 2 649 1 sky130_fd_sc_hd__and2_1 $T=73600 367200 1 0 $X=73410 $Y=364240
X2123 1 2 88 19 2 671 1 sky130_fd_sc_hd__and2_1 $T=80500 334560 1 0 $X=80310 $Y=331600
X2124 1 2 89 19 2 670 1 sky130_fd_sc_hd__and2_1 $T=80500 350880 1 0 $X=80310 $Y=347920
X2125 1 2 91 19 2 681 1 sky130_fd_sc_hd__and2_1 $T=84640 318240 1 0 $X=84450 $Y=315280
X2126 1 2 93 19 2 673 1 sky130_fd_sc_hd__and2_1 $T=85100 329120 0 0 $X=84910 $Y=328880
X2127 1 2 102 19 2 711 1 sky130_fd_sc_hd__and2_1 $T=104420 367200 1 0 $X=104230 $Y=364240
X2128 1 2 106 19 2 728 1 sky130_fd_sc_hd__and2_1 $T=108100 323680 0 0 $X=107910 $Y=323440
X2129 1 2 117 19 2 745 1 sky130_fd_sc_hd__and2_1 $T=117760 318240 1 0 $X=117570 $Y=315280
X2130 1 2 119 19 2 737 1 sky130_fd_sc_hd__and2_1 $T=118220 345440 0 0 $X=118030 $Y=345200
X2131 1 2 120 19 2 748 1 sky130_fd_sc_hd__and2_1 $T=118220 356320 0 0 $X=118030 $Y=356080
X2132 1 2 134 19 2 775 1 sky130_fd_sc_hd__and2_1 $T=138000 329120 1 0 $X=137810 $Y=326160
X2133 1 2 141 19 2 776 1 sky130_fd_sc_hd__and2_1 $T=143520 345440 1 0 $X=143330 $Y=342480
X2134 1 2 142 19 2 788 1 sky130_fd_sc_hd__and2_1 $T=143520 356320 0 0 $X=143330 $Y=356080
X2135 1 2 29 144 2 789 1 sky130_fd_sc_hd__and2_1 $T=143520 361760 0 0 $X=143330 $Y=361520
X2136 1 2 147 19 2 793 1 sky130_fd_sc_hd__and2_1 $T=148580 329120 1 0 $X=148390 $Y=326160
X2137 1 2 26 164 2 822 1 sky130_fd_sc_hd__and2_1 $T=163300 340000 0 0 $X=163110 $Y=339760
X2138 1 2 56 164 2 815 1 sky130_fd_sc_hd__and2_1 $T=164680 329120 1 0 $X=164490 $Y=326160
X2139 1 2 17 164 2 824 1 sky130_fd_sc_hd__and2_1 $T=165600 318240 1 0 $X=165410 $Y=315280
X2140 1 2 60 144 2 840 1 sky130_fd_sc_hd__and2_1 $T=184460 372640 1 0 $X=184270 $Y=369680
X2141 1 2 62 164 2 849 1 sky130_fd_sc_hd__and2_1 $T=185380 334560 1 0 $X=185190 $Y=331600
X2142 1 2 30 164 2 850 1 sky130_fd_sc_hd__and2_1 $T=188600 356320 1 0 $X=188410 $Y=353360
X2143 1 2 74 164 2 204 1 sky130_fd_sc_hd__and2_1 $T=189520 318240 1 0 $X=189330 $Y=315280
X2144 1 2 85 144 2 858 1 sky130_fd_sc_hd__and2_1 $T=198720 361760 0 0 $X=198530 $Y=361520
X2145 1 2 68 164 2 883 1 sky130_fd_sc_hd__and2_1 $T=202860 329120 0 0 $X=202670 $Y=328880
X2146 1 2 112 144 2 212 1 sky130_fd_sc_hd__and2_1 $T=213900 372640 1 0 $X=213710 $Y=369680
X2147 1 2 69 164 2 906 1 sky130_fd_sc_hd__and2_1 $T=218960 350880 0 0 $X=218770 $Y=350640
X2148 1 2 89 164 2 917 1 sky130_fd_sc_hd__and2_1 $T=223100 334560 0 0 $X=222910 $Y=334320
X2149 1 2 81 164 2 938 1 sky130_fd_sc_hd__and2_1 $T=234600 356320 0 0 $X=234410 $Y=356080
X2150 1 2 143 144 2 951 1 sky130_fd_sc_hd__and2_1 $T=241040 367200 1 0 $X=240850 $Y=364240
X2151 1 2 106 164 2 953 1 sky130_fd_sc_hd__and2_1 $T=244720 318240 1 0 $X=244530 $Y=315280
X2152 1 2 88 164 2 990 1 sky130_fd_sc_hd__and2_1 $T=262660 334560 1 0 $X=262470 $Y=331600
X2153 1 2 119 164 2 999 1 sky130_fd_sc_hd__and2_1 $T=264040 350880 1 0 $X=263850 $Y=347920
X2154 1 2 141 144 2 1014 1 sky130_fd_sc_hd__and2_1 $T=270020 372640 1 0 $X=269830 $Y=369680
X2155 1 2 147 164 2 1032 1 sky130_fd_sc_hd__and2_1 $T=283820 318240 1 0 $X=283630 $Y=315280
X2156 1 2 93 164 2 1038 1 sky130_fd_sc_hd__and2_1 $T=283820 329120 0 0 $X=283630 $Y=328880
X2157 1 2 120 164 2 1031 1 sky130_fd_sc_hd__and2_1 $T=284280 356320 1 0 $X=284090 $Y=353360
X2158 1 2 142 164 2 1062 1 sky130_fd_sc_hd__and2_1 $T=298080 350880 1 0 $X=297890 $Y=347920
X2159 1 2 141 164 2 1071 1 sky130_fd_sc_hd__and2_1 $T=301300 334560 1 0 $X=301110 $Y=331600
X2160 1 2 134 164 2 1078 1 sky130_fd_sc_hd__and2_1 $T=304520 318240 0 0 $X=304330 $Y=318000
X2161 1 2 281 272 2 1136 1 sky130_fd_sc_hd__and2_1 $T=339020 350880 0 0 $X=338830 $Y=350640
X2162 1 2 283 272 2 1137 1 sky130_fd_sc_hd__and2_1 $T=339940 356320 0 0 $X=339750 $Y=356080
X2163 1 2 285 272 2 1147 1 sky130_fd_sc_hd__and2_1 $T=342700 334560 0 0 $X=342510 $Y=334320
X2164 1 2 286 272 2 1148 1 sky130_fd_sc_hd__and2_1 $T=342700 340000 0 0 $X=342510 $Y=339760
X2165 1 2 288 272 2 1152 1 sky130_fd_sc_hd__and2_1 $T=346840 372640 0 0 $X=346650 $Y=372400
X2166 1 2 292 272 2 1157 1 sky130_fd_sc_hd__and2_1 $T=349600 318240 0 0 $X=349410 $Y=318000
X2167 1 2 297 272 2 1164 1 sky130_fd_sc_hd__and2_1 $T=354200 350880 1 0 $X=354010 $Y=347920
X2168 1 2 310 272 2 1193 1 sky130_fd_sc_hd__and2_1 $T=368000 372640 0 0 $X=367810 $Y=372400
X2169 1 2 314 272 2 1199 1 sky130_fd_sc_hd__and2_1 $T=375820 345440 0 0 $X=375630 $Y=345200
X2170 1 2 316 272 2 1204 1 sky130_fd_sc_hd__and2_1 $T=376280 340000 0 0 $X=376090 $Y=339760
X2171 1 2 317 272 2 1206 1 sky130_fd_sc_hd__and2_1 $T=377200 367200 0 0 $X=377010 $Y=366960
X2172 1 2 330 272 2 1253 1 sky130_fd_sc_hd__and2_1 $T=398820 323680 0 0 $X=398630 $Y=323440
X2173 1 2 331 272 2 1251 1 sky130_fd_sc_hd__and2_1 $T=405260 318240 0 0 $X=405070 $Y=318000
X2174 1 2 335 272 2 1258 1 sky130_fd_sc_hd__and2_1 $T=408940 345440 1 0 $X=408750 $Y=342480
X2175 1 2 338 272 2 1282 1 sky130_fd_sc_hd__and2_1 $T=416300 312800 0 0 $X=416110 $Y=312560
X2176 1 2 340 272 2 1289 1 sky130_fd_sc_hd__and2_1 $T=418140 361760 1 0 $X=417950 $Y=358800
X2177 1 2 348 272 2 1291 1 sky130_fd_sc_hd__and2_1 $T=426880 340000 0 0 $X=426690 $Y=339760
X2178 1 2 350 272 2 351 1 sky130_fd_sc_hd__and2_1 $T=431480 372640 0 0 $X=431290 $Y=372400
X2179 1 2 352 272 2 1328 1 sky130_fd_sc_hd__and2_1 $T=438380 361760 1 0 $X=438190 $Y=358800
X2180 1 2 353 272 2 1318 1 sky130_fd_sc_hd__and2_1 $T=439300 329120 0 0 $X=439110 $Y=328880
X2181 1 2 354 272 2 1330 1 sky130_fd_sc_hd__and2_1 $T=441140 318240 1 0 $X=440950 $Y=315280
X2182 1 2 355 272 2 1335 1 sky130_fd_sc_hd__and2_1 $T=441600 372640 1 0 $X=441410 $Y=369680
X2183 1 2 363 272 2 1364 1 sky130_fd_sc_hd__and2_1 $T=463220 356320 0 0 $X=463030 $Y=356080
X2184 1 2 364 272 2 1379 1 sky130_fd_sc_hd__and2_1 $T=463220 372640 0 0 $X=463030 $Y=372400
X2185 1 2 366 272 2 1386 1 sky130_fd_sc_hd__and2_1 $T=466440 345440 1 0 $X=466250 $Y=342480
X2186 1 2 373 272 2 1407 1 sky130_fd_sc_hd__and2_1 $T=478860 318240 0 0 $X=478670 $Y=318000
X2187 1 2 374 272 2 1397 1 sky130_fd_sc_hd__and2_1 $T=479780 334560 0 0 $X=479590 $Y=334320
X2188 1 2 375 272 2 1419 1 sky130_fd_sc_hd__and2_1 $T=485760 367200 1 0 $X=485570 $Y=364240
X2189 1 2 379 272 2 1459 1 sky130_fd_sc_hd__and2_1 $T=497260 361760 1 0 $X=497070 $Y=358800
X2190 1 2 385 272 2 1461 1 sky130_fd_sc_hd__and2_1 $T=500940 334560 0 0 $X=500750 $Y=334320
X2191 1 2 386 272 2 1458 1 sky130_fd_sc_hd__and2_1 $T=501400 350880 1 0 $X=501210 $Y=347920
X2192 1 2 292 387 2 1483 1 sky130_fd_sc_hd__and2_1 $T=513820 318240 1 0 $X=513630 $Y=315280
X2193 1 2 288 387 2 1489 1 sky130_fd_sc_hd__and2_1 $T=516580 345440 0 0 $X=516390 $Y=345200
X2194 1 2 310 387 2 1490 1 sky130_fd_sc_hd__and2_1 $T=517040 334560 0 0 $X=516850 $Y=334320
X2195 1 2 321 387 2 1491 1 sky130_fd_sc_hd__and2_1 $T=521180 356320 1 0 $X=520990 $Y=353360
X2196 1 2 285 387 2 1528 1 sky130_fd_sc_hd__and2_1 $T=543260 329120 0 0 $X=543070 $Y=328880
X2197 1 2 314 387 2 1530 1 sky130_fd_sc_hd__and2_1 $T=550620 345440 1 0 $X=550430 $Y=342480
X2198 1 2 336 387 2 1536 1 sky130_fd_sc_hd__and2_1 $T=552460 372640 0 0 $X=552270 $Y=372400
X2199 1 2 317 387 2 1546 1 sky130_fd_sc_hd__and2_1 $T=553380 367200 1 0 $X=553190 $Y=364240
X2200 1 2 330 387 2 1560 1 sky130_fd_sc_hd__and2_1 $T=563500 334560 1 0 $X=563310 $Y=331600
X2201 1 2 297 387 2 1565 1 sky130_fd_sc_hd__and2_1 $T=564420 345440 0 0 $X=564230 $Y=345200
X2202 1 2 392 387 2 1577 1 sky130_fd_sc_hd__and2_1 $T=568560 318240 1 0 $X=568370 $Y=315280
X2203 1 2 283 387 2 1595 1 sky130_fd_sc_hd__and2_1 $T=577760 361760 1 0 $X=577570 $Y=358800
X2204 1 2 271 387 2 1596 1 sky130_fd_sc_hd__and2_1 $T=578680 372640 0 0 $X=578490 $Y=372400
X2205 1 2 281 387 2 1607 1 sky130_fd_sc_hd__and2_1 $T=581440 356320 1 0 $X=581250 $Y=353360
X2206 1 2 324 387 2 435 1 sky130_fd_sc_hd__and2_1 $T=584200 312800 0 0 $X=584010 $Y=312560
X2207 1 2 353 387 2 1620 1 sky130_fd_sc_hd__and2_1 $T=594780 340000 1 0 $X=594590 $Y=337040
X2208 1 2 335 387 2 1649 1 sky130_fd_sc_hd__and2_1 $T=601680 356320 0 0 $X=601490 $Y=356080
X2209 1 2 352 387 2 1651 1 sky130_fd_sc_hd__and2_1 $T=603520 361760 0 0 $X=603330 $Y=361520
X2210 1 2 286 387 2 1660 1 sky130_fd_sc_hd__and2_1 $T=606280 345440 1 0 $X=606090 $Y=342480
X2211 1 2 419 387 2 1636 1 sky130_fd_sc_hd__and2_1 $T=609500 318240 1 0 $X=609310 $Y=315280
X2212 1 2 316 387 2 1664 1 sky130_fd_sc_hd__and2_1 $T=609500 334560 1 0 $X=609310 $Y=331600
X2213 1 2 338 387 2 1692 1 sky130_fd_sc_hd__and2_1 $T=623760 318240 1 0 $X=623570 $Y=315280
X2214 1 2 350 387 2 448 1 sky130_fd_sc_hd__and2_1 $T=628820 372640 0 0 $X=628630 $Y=372400
X2215 1 2 340 387 2 1697 1 sky130_fd_sc_hd__and2_1 $T=630660 361760 0 0 $X=630470 $Y=361520
X2216 1 2 348 387 2 1707 1 sky130_fd_sc_hd__and2_1 $T=631580 350880 0 0 $X=631390 $Y=350640
X2217 1 2 295 387 2 1709 1 sky130_fd_sc_hd__and2_1 $T=633420 334560 1 0 $X=633230 $Y=331600
X2218 1 2 345 387 2 1711 1 sky130_fd_sc_hd__and2_1 $T=636180 340000 0 0 $X=635990 $Y=339760
X2219 1 2 374 387 2 1767 1 sky130_fd_sc_hd__and2_1 $T=662400 334560 1 0 $X=662210 $Y=331600
X2220 1 2 366 387 2 1770 1 sky130_fd_sc_hd__and2_1 $T=665620 350880 1 0 $X=665430 $Y=347920
X2221 1 2 363 387 2 1765 1 sky130_fd_sc_hd__and2_1 $T=665620 361760 1 0 $X=665430 $Y=358800
X2222 1 2 354 387 2 1799 1 sky130_fd_sc_hd__and2_1 $T=676660 312800 0 0 $X=676470 $Y=312560
X2223 1 2 355 387 2 1805 1 sky130_fd_sc_hd__and2_1 $T=679880 361760 0 0 $X=679690 $Y=361520
X2224 1 2 460 387 2 461 1 sky130_fd_sc_hd__and2_1 $T=690920 378080 1 0 $X=690730 $Y=375120
X2225 1 2 388 387 2 1845 1 sky130_fd_sc_hd__and2_1 $T=701040 323680 1 0 $X=700850 $Y=320720
X2226 1 2 379 387 2 1852 1 sky130_fd_sc_hd__and2_1 $T=703800 356320 0 0 $X=703610 $Y=356080
X2227 1 2 364 387 2 1854 1 sky130_fd_sc_hd__and2_1 $T=704260 372640 0 0 $X=704070 $Y=372400
X2228 1 2 373 387 2 1849 1 sky130_fd_sc_hd__and2_1 $T=704720 312800 0 0 $X=704530 $Y=312560
X2229 1 2 375 387 2 1856 1 sky130_fd_sc_hd__and2_1 $T=704720 361760 0 0 $X=704530 $Y=361520
X2230 1 2 380 387 2 1846 1 sky130_fd_sc_hd__and2_1 $T=707480 329120 0 0 $X=707290 $Y=328880
X2231 1 2 386 387 2 1853 1 sky130_fd_sc_hd__and2_1 $T=707480 350880 0 0 $X=707290 $Y=350640
X2232 1 2 200 527 2 525 1 sky130_fd_sc_hd__dlclkp_1 $T=6900 340000 0 0 $X=6710 $Y=339760
X2233 1 2 200 528 2 9 1 sky130_fd_sc_hd__dlclkp_1 $T=7820 367200 1 0 $X=7630 $Y=364240
X2234 1 2 200 530 2 526 1 sky130_fd_sc_hd__dlclkp_1 $T=8280 361760 1 0 $X=8090 $Y=358800
X2235 1 2 200 529 2 531 1 sky130_fd_sc_hd__dlclkp_1 $T=15180 334560 0 0 $X=14990 $Y=334320
X2236 1 2 200 559 2 524 1 sky130_fd_sc_hd__dlclkp_1 $T=24380 323680 0 0 $X=24190 $Y=323440
X2237 1 2 200 573 2 575 1 sky130_fd_sc_hd__dlclkp_1 $T=28980 361760 1 0 $X=28790 $Y=358800
X2238 1 2 200 576 2 580 1 sky130_fd_sc_hd__dlclkp_1 $T=31280 345440 1 0 $X=31090 $Y=342480
X2239 1 2 200 577 2 48 1 sky130_fd_sc_hd__dlclkp_1 $T=31280 367200 1 0 $X=31090 $Y=364240
X2240 1 2 200 604 2 608 1 sky130_fd_sc_hd__dlclkp_1 $T=45540 361760 0 0 $X=45350 $Y=361520
X2241 1 2 200 610 2 66 1 sky130_fd_sc_hd__dlclkp_1 $T=48300 318240 1 0 $X=48110 $Y=315280
X2242 1 2 200 603 2 591 1 sky130_fd_sc_hd__dlclkp_1 $T=50140 323680 0 0 $X=49950 $Y=323440
X2243 1 2 200 625 2 602 1 sky130_fd_sc_hd__dlclkp_1 $T=56580 367200 1 0 $X=56390 $Y=364240
X2244 1 2 200 626 2 627 1 sky130_fd_sc_hd__dlclkp_1 $T=59340 334560 1 0 $X=59150 $Y=331600
X2245 1 2 200 649 2 83 1 sky130_fd_sc_hd__dlclkp_1 $T=67160 367200 1 0 $X=66970 $Y=364240
X2246 1 2 200 646 2 644 1 sky130_fd_sc_hd__dlclkp_1 $T=69460 361760 0 0 $X=69270 $Y=361520
X2247 1 2 200 670 2 672 1 sky130_fd_sc_hd__dlclkp_1 $T=77280 340000 0 0 $X=77090 $Y=339760
X2248 1 2 200 671 2 637 1 sky130_fd_sc_hd__dlclkp_1 $T=78660 329120 0 0 $X=78470 $Y=328880
X2249 1 2 200 673 2 687 1 sky130_fd_sc_hd__dlclkp_1 $T=81420 329120 1 0 $X=81230 $Y=326160
X2250 1 2 200 681 2 94 1 sky130_fd_sc_hd__dlclkp_1 $T=82800 312800 0 0 $X=82610 $Y=312560
X2251 1 2 200 711 2 694 1 sky130_fd_sc_hd__dlclkp_1 $T=97520 361760 1 0 $X=97330 $Y=358800
X2252 1 2 200 728 2 732 1 sky130_fd_sc_hd__dlclkp_1 $T=107640 329120 0 0 $X=107450 $Y=328880
X2253 1 2 200 737 2 720 1 sky130_fd_sc_hd__dlclkp_1 $T=111320 345440 0 0 $X=111130 $Y=345200
X2254 1 2 200 748 2 744 1 sky130_fd_sc_hd__dlclkp_1 $T=118220 350880 0 0 $X=118030 $Y=350640
X2255 1 2 200 745 2 118 1 sky130_fd_sc_hd__dlclkp_1 $T=120520 318240 0 0 $X=120330 $Y=318000
X2256 1 2 200 775 2 772 1 sky130_fd_sc_hd__dlclkp_1 $T=137080 323680 0 0 $X=136890 $Y=323440
X2257 1 2 200 776 2 750 1 sky130_fd_sc_hd__dlclkp_1 $T=137080 345440 1 0 $X=136890 $Y=342480
X2258 1 2 200 788 2 785 1 sky130_fd_sc_hd__dlclkp_1 $T=146280 361760 0 0 $X=146090 $Y=361520
X2259 1 2 200 793 2 786 1 sky130_fd_sc_hd__dlclkp_1 $T=147200 329120 0 0 $X=147010 $Y=328880
X2260 1 2 200 789 2 800 1 sky130_fd_sc_hd__dlclkp_1 $T=153180 361760 0 0 $X=152990 $Y=361520
X2261 1 2 200 815 2 825 1 sky130_fd_sc_hd__dlclkp_1 $T=160080 323680 0 0 $X=159890 $Y=323440
X2262 1 2 200 822 2 826 1 sky130_fd_sc_hd__dlclkp_1 $T=162840 345440 1 0 $X=162650 $Y=342480
X2263 1 2 200 824 2 173 1 sky130_fd_sc_hd__dlclkp_1 $T=164220 312800 0 0 $X=164030 $Y=312560
X2264 1 2 200 840 2 195 1 sky130_fd_sc_hd__dlclkp_1 $T=181240 378080 1 0 $X=181050 $Y=375120
X2265 1 2 200 849 2 853 1 sky130_fd_sc_hd__dlclkp_1 $T=185840 329120 0 0 $X=185650 $Y=328880
X2266 1 2 200 850 2 855 1 sky130_fd_sc_hd__dlclkp_1 $T=186300 356320 0 0 $X=186110 $Y=356080
X2267 1 2 200 858 2 859 1 sky130_fd_sc_hd__dlclkp_1 $T=192280 361760 0 0 $X=192090 $Y=361520
X2268 1 2 200 883 2 882 1 sky130_fd_sc_hd__dlclkp_1 $T=202860 329120 1 0 $X=202670 $Y=326160
X2269 1 2 200 213 2 218 1 sky130_fd_sc_hd__dlclkp_1 $T=214360 312800 0 0 $X=214170 $Y=312560
X2270 1 2 200 906 2 913 1 sky130_fd_sc_hd__dlclkp_1 $T=216660 356320 1 0 $X=216470 $Y=353360
X2271 1 2 200 917 2 914 1 sky130_fd_sc_hd__dlclkp_1 $T=222180 329120 0 0 $X=221990 $Y=328880
X2272 1 2 200 938 2 939 1 sky130_fd_sc_hd__dlclkp_1 $T=233680 356320 1 0 $X=233490 $Y=353360
X2273 1 2 200 951 2 963 1 sky130_fd_sc_hd__dlclkp_1 $T=240580 367200 0 0 $X=240390 $Y=366960
X2274 1 2 200 953 2 223 1 sky130_fd_sc_hd__dlclkp_1 $T=241960 312800 0 0 $X=241770 $Y=312560
X2275 1 2 200 990 2 992 1 sky130_fd_sc_hd__dlclkp_1 $T=259440 334560 0 0 $X=259250 $Y=334320
X2276 1 2 200 999 2 995 1 sky130_fd_sc_hd__dlclkp_1 $T=264040 350880 0 0 $X=263850 $Y=350640
X2277 1 2 200 1014 2 1022 1 sky130_fd_sc_hd__dlclkp_1 $T=272320 367200 0 0 $X=272130 $Y=366960
X2278 1 2 200 240 2 242 1 sky130_fd_sc_hd__dlclkp_1 $T=272780 378080 1 0 $X=272590 $Y=375120
X2279 1 2 200 1031 2 1030 1 sky130_fd_sc_hd__dlclkp_1 $T=279220 350880 0 0 $X=279030 $Y=350640
X2280 1 2 200 1032 2 244 1 sky130_fd_sc_hd__dlclkp_1 $T=279680 318240 0 0 $X=279490 $Y=318000
X2281 1 2 200 1038 2 1035 1 sky130_fd_sc_hd__dlclkp_1 $T=286580 334560 1 0 $X=286390 $Y=331600
X2282 1 2 200 1062 2 1061 1 sky130_fd_sc_hd__dlclkp_1 $T=297160 350880 0 0 $X=296970 $Y=350640
X2283 1 2 200 1071 2 1073 1 sky130_fd_sc_hd__dlclkp_1 $T=300840 334560 0 0 $X=300650 $Y=334320
X2284 1 2 200 1078 2 250 1 sky130_fd_sc_hd__dlclkp_1 $T=307280 323680 1 0 $X=307090 $Y=320720
X2285 1 2 276 1136 2 1102 1 sky130_fd_sc_hd__dlclkp_1 $T=335800 356320 1 0 $X=335610 $Y=353360
X2286 1 2 276 1137 2 1146 1 sky130_fd_sc_hd__dlclkp_1 $T=335800 361760 0 0 $X=335610 $Y=361520
X2287 1 2 276 1147 2 1118 1 sky130_fd_sc_hd__dlclkp_1 $T=341320 334560 1 0 $X=341130 $Y=331600
X2288 1 2 276 1152 2 293 1 sky130_fd_sc_hd__dlclkp_1 $T=344080 378080 1 0 $X=343890 $Y=375120
X2289 1 2 276 1148 2 1112 1 sky130_fd_sc_hd__dlclkp_1 $T=345920 345440 1 0 $X=345730 $Y=342480
X2290 1 2 276 1157 2 278 1 sky130_fd_sc_hd__dlclkp_1 $T=347760 323680 1 0 $X=347570 $Y=320720
X2291 1 2 276 1164 2 1169 1 sky130_fd_sc_hd__dlclkp_1 $T=350060 345440 0 0 $X=349870 $Y=345200
X2292 1 2 276 307 2 309 1 sky130_fd_sc_hd__dlclkp_1 $T=362480 312800 0 0 $X=362290 $Y=312560
X2293 1 2 276 1193 2 312 1 sky130_fd_sc_hd__dlclkp_1 $T=370760 367200 0 0 $X=370570 $Y=366960
X2294 1 2 276 1199 2 1205 1 sky130_fd_sc_hd__dlclkp_1 $T=371220 350880 0 0 $X=371030 $Y=350640
X2295 1 2 276 1204 2 1203 1 sky130_fd_sc_hd__dlclkp_1 $T=375360 334560 0 0 $X=375170 $Y=334320
X2296 1 2 276 1206 2 1187 1 sky130_fd_sc_hd__dlclkp_1 $T=375360 367200 1 0 $X=375170 $Y=364240
X2297 1 2 276 327 2 329 1 sky130_fd_sc_hd__dlclkp_1 $T=393760 378080 1 0 $X=393570 $Y=375120
X2298 1 2 276 1251 2 325 1 sky130_fd_sc_hd__dlclkp_1 $T=398820 318240 0 0 $X=398630 $Y=318000
X2299 1 2 276 1253 2 1229 1 sky130_fd_sc_hd__dlclkp_1 $T=400200 329120 0 0 $X=400010 $Y=328880
X2300 1 2 276 1258 2 1249 1 sky130_fd_sc_hd__dlclkp_1 $T=402500 345440 1 0 $X=402310 $Y=342480
X2301 1 2 276 1282 2 342 1 sky130_fd_sc_hd__dlclkp_1 $T=414920 318240 1 0 $X=414730 $Y=315280
X2302 1 2 276 1289 2 1257 1 sky130_fd_sc_hd__dlclkp_1 $T=419980 356320 0 0 $X=419790 $Y=356080
X2303 1 2 276 1291 2 1301 1 sky130_fd_sc_hd__dlclkp_1 $T=420440 345440 1 0 $X=420250 $Y=342480
X2304 1 2 276 1318 2 1331 1 sky130_fd_sc_hd__dlclkp_1 $T=434240 334560 1 0 $X=434050 $Y=331600
X2305 1 2 276 1328 2 1294 1 sky130_fd_sc_hd__dlclkp_1 $T=436540 361760 0 0 $X=436350 $Y=361520
X2306 1 2 276 1330 2 356 1 sky130_fd_sc_hd__dlclkp_1 $T=437460 318240 0 0 $X=437270 $Y=318000
X2307 1 2 276 1335 2 1334 1 sky130_fd_sc_hd__dlclkp_1 $T=444820 372640 0 0 $X=444630 $Y=372400
X2308 1 2 276 1364 2 1339 1 sky130_fd_sc_hd__dlclkp_1 $T=456320 356320 1 0 $X=456130 $Y=353360
X2309 1 2 276 1379 2 1385 1 sky130_fd_sc_hd__dlclkp_1 $T=462300 372640 1 0 $X=462110 $Y=369680
X2310 1 2 276 1386 2 1360 1 sky130_fd_sc_hd__dlclkp_1 $T=465060 340000 0 0 $X=464870 $Y=339760
X2311 1 2 276 1397 2 1378 1 sky130_fd_sc_hd__dlclkp_1 $T=471500 334560 1 0 $X=471310 $Y=331600
X2312 1 2 276 1407 2 365 1 sky130_fd_sc_hd__dlclkp_1 $T=476560 318240 1 0 $X=476370 $Y=315280
X2313 1 2 276 376 2 378 1 sky130_fd_sc_hd__dlclkp_1 $T=483000 318240 1 0 $X=482810 $Y=315280
X2314 1 2 276 1419 2 1384 1 sky130_fd_sc_hd__dlclkp_1 $T=483000 361760 0 0 $X=482810 $Y=361520
X2315 1 2 276 1458 2 1413 1 sky130_fd_sc_hd__dlclkp_1 $T=496800 345440 0 0 $X=496610 $Y=345200
X2316 1 2 276 1459 2 1431 1 sky130_fd_sc_hd__dlclkp_1 $T=496800 356320 0 0 $X=496610 $Y=356080
X2317 1 2 276 383 2 1429 1 sky130_fd_sc_hd__dlclkp_1 $T=496800 372640 0 0 $X=496610 $Y=372400
X2318 1 2 276 1461 2 1428 1 sky130_fd_sc_hd__dlclkp_1 $T=498180 340000 1 0 $X=497990 $Y=337040
X2319 1 2 276 1483 2 1484 1 sky130_fd_sc_hd__dlclkp_1 $T=513820 312800 0 0 $X=513630 $Y=312560
X2320 1 2 276 1490 2 1485 1 sky130_fd_sc_hd__dlclkp_1 $T=518420 340000 1 0 $X=518230 $Y=337040
X2321 1 2 276 1489 2 1486 1 sky130_fd_sc_hd__dlclkp_1 $T=518420 350880 1 0 $X=518230 $Y=347920
X2322 1 2 276 1491 2 1496 1 sky130_fd_sc_hd__dlclkp_1 $T=519800 356320 0 0 $X=519610 $Y=356080
X2323 1 2 276 423 2 427 1 sky130_fd_sc_hd__dlclkp_1 $T=540960 312800 0 0 $X=540770 $Y=312560
X2324 1 2 276 1528 2 1529 1 sky130_fd_sc_hd__dlclkp_1 $T=542340 334560 1 0 $X=542150 $Y=331600
X2325 1 2 276 1530 2 1527 1 sky130_fd_sc_hd__dlclkp_1 $T=543260 345440 0 0 $X=543070 $Y=345200
X2326 1 2 276 1536 2 1540 1 sky130_fd_sc_hd__dlclkp_1 $T=546020 372640 0 0 $X=545830 $Y=372400
X2327 1 2 276 1546 2 1551 1 sky130_fd_sc_hd__dlclkp_1 $T=548320 361760 0 0 $X=548130 $Y=361520
X2328 1 2 276 1560 2 1574 1 sky130_fd_sc_hd__dlclkp_1 $T=559360 334560 0 0 $X=559170 $Y=334320
X2329 1 2 276 1565 2 1575 1 sky130_fd_sc_hd__dlclkp_1 $T=560280 350880 0 0 $X=560090 $Y=350640
X2330 1 2 276 1577 2 1578 1 sky130_fd_sc_hd__dlclkp_1 $T=566260 323680 1 0 $X=566070 $Y=320720
X2331 1 2 276 1595 2 1602 1 sky130_fd_sc_hd__dlclkp_1 $T=573160 367200 1 0 $X=572970 $Y=364240
X2332 1 2 276 1596 2 434 1 sky130_fd_sc_hd__dlclkp_1 $T=574540 378080 1 0 $X=574350 $Y=375120
X2333 1 2 276 1607 2 1612 1 sky130_fd_sc_hd__dlclkp_1 $T=579140 356320 0 0 $X=578950 $Y=356080
X2334 1 2 276 1620 2 1618 1 sky130_fd_sc_hd__dlclkp_1 $T=586040 334560 0 0 $X=585850 $Y=334320
X2335 1 2 276 1636 2 1640 1 sky130_fd_sc_hd__dlclkp_1 $T=595240 318240 1 0 $X=595050 $Y=315280
X2336 1 2 276 1649 2 1652 1 sky130_fd_sc_hd__dlclkp_1 $T=602140 356320 1 0 $X=601950 $Y=353360
X2337 1 2 276 1651 2 1655 1 sky130_fd_sc_hd__dlclkp_1 $T=602600 361760 1 0 $X=602410 $Y=358800
X2338 1 2 276 1660 2 1661 1 sky130_fd_sc_hd__dlclkp_1 $T=605820 340000 0 0 $X=605630 $Y=339760
X2339 1 2 276 1664 2 1663 1 sky130_fd_sc_hd__dlclkp_1 $T=609500 329120 1 0 $X=609310 $Y=326160
X2340 1 2 276 1692 2 446 1 sky130_fd_sc_hd__dlclkp_1 $T=623300 312800 0 0 $X=623110 $Y=312560
X2341 1 2 276 1697 2 1699 1 sky130_fd_sc_hd__dlclkp_1 $T=626520 361760 1 0 $X=626330 $Y=358800
X2342 1 2 276 1707 2 1713 1 sky130_fd_sc_hd__dlclkp_1 $T=629740 350880 1 0 $X=629550 $Y=347920
X2343 1 2 276 1709 2 1712 1 sky130_fd_sc_hd__dlclkp_1 $T=630660 329120 0 0 $X=630470 $Y=328880
X2344 1 2 276 1711 2 1720 1 sky130_fd_sc_hd__dlclkp_1 $T=632960 334560 0 0 $X=632770 $Y=334320
X2345 1 2 276 1765 2 1756 1 sky130_fd_sc_hd__dlclkp_1 $T=658720 361760 1 0 $X=658530 $Y=358800
X2346 1 2 276 1767 2 1775 1 sky130_fd_sc_hd__dlclkp_1 $T=660100 329120 0 0 $X=659910 $Y=328880
X2347 1 2 276 1770 2 1779 1 sky130_fd_sc_hd__dlclkp_1 $T=661480 345440 0 0 $X=661290 $Y=345200
X2348 1 2 276 1799 2 1801 1 sky130_fd_sc_hd__dlclkp_1 $T=674360 318240 1 0 $X=674170 $Y=315280
X2349 1 2 276 1805 2 1808 1 sky130_fd_sc_hd__dlclkp_1 $T=679880 367200 1 0 $X=679690 $Y=364240
X2350 1 2 276 464 2 465 1 sky130_fd_sc_hd__dlclkp_1 $T=698280 312800 0 0 $X=698090 $Y=312560
X2351 1 2 276 1845 2 1850 1 sky130_fd_sc_hd__dlclkp_1 $T=699660 323680 0 0 $X=699470 $Y=323440
X2352 1 2 276 1846 2 1859 1 sky130_fd_sc_hd__dlclkp_1 $T=700580 329120 0 0 $X=700390 $Y=328880
X2353 1 2 276 1849 2 466 1 sky130_fd_sc_hd__dlclkp_1 $T=701040 318240 1 0 $X=700850 $Y=315280
X2354 1 2 276 1852 2 1860 1 sky130_fd_sc_hd__dlclkp_1 $T=701500 361760 1 0 $X=701310 $Y=358800
X2355 1 2 276 1853 2 1861 1 sky130_fd_sc_hd__dlclkp_1 $T=701960 350880 1 0 $X=701770 $Y=347920
X2356 1 2 276 1854 2 467 1 sky130_fd_sc_hd__dlclkp_1 $T=701960 378080 1 0 $X=701770 $Y=375120
X2357 1 2 276 1856 2 1862 1 sky130_fd_sc_hd__dlclkp_1 $T=702420 367200 1 0 $X=702230 $Y=364240
X2358 1 2 525 14 541 ICV_35 $T=6900 334560 0 0 $X=6710 $Y=334320
X2359 1 2 526 15 543 ICV_35 $T=6900 356320 0 0 $X=6710 $Y=356080
X2360 1 2 525 44 568 ICV_35 $T=20240 345440 1 0 $X=20050 $Y=342480
X2361 1 2 602 20 614 ICV_35 $T=45540 372640 0 0 $X=45350 $Y=372400
X2362 1 2 82 18 656 ICV_35 $T=66240 312800 0 0 $X=66050 $Y=312560
X2363 1 2 82 15 657 ICV_35 $T=66240 318240 1 0 $X=66050 $Y=315280
X2364 1 2 627 18 655 ICV_35 $T=67620 340000 1 0 $X=67430 $Y=337040
X2365 1 2 644 25 661 ICV_35 $T=67620 350880 1 0 $X=67430 $Y=347920
X2366 1 2 672 43 688 ICV_35 $T=80960 345440 0 0 $X=80770 $Y=345200
X2367 1 2 672 13 691 ICV_35 $T=81420 334560 0 0 $X=81230 $Y=334320
X2368 1 2 98 10 716 ICV_35 $T=93840 361760 0 0 $X=93650 $Y=361520
X2369 1 2 694 14 725 ICV_35 $T=97520 350880 0 0 $X=97330 $Y=350640
X2370 1 2 772 44 790 ICV_35 $T=140300 329120 1 0 $X=140110 $Y=326160
X2371 1 2 826 170 819 ICV_35 $T=165600 334560 0 0 $X=165410 $Y=334320
X2372 1 2 826 171 833 ICV_35 $T=165600 340000 0 0 $X=165410 $Y=339760
X2373 1 2 800 175 837 ICV_35 $T=167900 367200 1 0 $X=167710 $Y=364240
X2374 1 2 160 181 192 ICV_35 $T=172040 378080 1 0 $X=171850 $Y=375120
X2375 1 2 853 170 862 ICV_35 $T=190440 312800 0 0 $X=190250 $Y=312560
X2376 1 2 859 161 880 ICV_35 $T=194580 361760 1 0 $X=194390 $Y=358800
X2377 1 2 859 158 903 ICV_35 $T=206540 361760 0 0 $X=206350 $Y=361520
X2378 1 2 882 171 904 ICV_35 $T=207920 318240 1 0 $X=207730 $Y=315280
X2379 1 2 907 152 919 ICV_35 $T=218040 367200 0 0 $X=217850 $Y=366960
X2380 1 2 214 161 935 ICV_35 $T=224020 378080 1 0 $X=223830 $Y=375120
X2381 1 2 165 38 236 ICV_35 $T=261280 361760 1 0 $X=261090 $Y=358800
X2382 1 2 1022 158 1037 ICV_35 $T=277380 361760 0 0 $X=277190 $Y=361520
X2383 1 2 1030 168 1040 ICV_35 $T=280140 340000 1 0 $X=279950 $Y=337040
X2384 1 2 1030 171 1055 ICV_35 $T=286580 356320 1 0 $X=286390 $Y=353360
X2385 1 2 1030 190 1058 ICV_35 $T=287960 350880 0 0 $X=287770 $Y=350640
X2386 1 2 1061 190 1084 ICV_35 $T=300840 350880 1 0 $X=300650 $Y=347920
X2387 1 2 1079 181 1092 ICV_35 $T=305900 367200 0 0 $X=305710 $Y=366960
X2388 1 2 1079 152 1140 ICV_35 $T=332580 372640 0 0 $X=332390 $Y=372400
X2389 1 2 1169 264 1172 ICV_35 $T=356960 340000 1 0 $X=356770 $Y=337040
X2390 1 2 309 260 1218 ICV_35 $T=378120 318240 0 0 $X=377930 $Y=318000
X2391 1 2 1187 262 1221 ICV_35 $T=378120 361760 0 0 $X=377930 $Y=361520
X2392 1 2 329 257 1260 ICV_35 $T=396520 372640 1 0 $X=396330 $Y=369680
X2393 1 2 1229 262 1279 ICV_35 $T=407560 318240 0 0 $X=407370 $Y=318000
X2394 1 2 1284 265 1322 ICV_35 $T=431020 329120 0 0 $X=430830 $Y=328880
X2395 1 2 1334 257 1348 ICV_35 $T=442980 367200 1 0 $X=442790 $Y=364240
X2396 1 2 1339 257 1357 ICV_35 $T=444820 350880 1 0 $X=444630 $Y=347920
X2397 1 2 1378 273 1390 ICV_35 $T=462300 329120 0 0 $X=462110 $Y=328880
X2398 1 2 1385 262 1389 ICV_35 $T=465060 367200 0 0 $X=464870 $Y=366960
X2399 1 2 1413 260 1441 ICV_35 $T=487140 345440 0 0 $X=486950 $Y=345200
X2400 1 2 1431 273 1452 ICV_35 $T=488520 356320 0 0 $X=488330 $Y=356080
X2401 1 2 1486 412 1521 ICV_35 $T=530380 340000 0 0 $X=530190 $Y=339760
X2402 1 2 1575 400 1608 ICV_35 $T=574540 340000 0 0 $X=574350 $Y=339760
X2403 1 2 447 410 1715 ICV_35 $T=628360 372640 1 0 $X=628170 $Y=369680
X2404 1 2 446 412 1732 ICV_35 $T=637560 318240 1 0 $X=637370 $Y=315280
X2405 1 2 1720 415 1739 ICV_35 $T=639400 334560 0 0 $X=639210 $Y=334320
X2406 1 2 1699 398 1746 ICV_35 $T=644000 367200 1 0 $X=643810 $Y=364240
X2407 1 2 1747 397 1776 ICV_35 $T=658720 323680 0 0 $X=658530 $Y=323440
X2408 1 2 1756 412 1795 ICV_35 $T=667000 361760 0 0 $X=666810 $Y=361520
X2409 1 2 1861 397 1875 ICV_35 $T=708400 350880 1 0 $X=708210 $Y=347920
X2410 1 2 526 44 563 ICV_37 $T=19780 361760 1 0 $X=19590 $Y=358800
X2411 1 2 41 18 572 ICV_37 $T=33580 312800 0 0 $X=33390 $Y=312560
X2412 1 2 575 14 586 ICV_37 $T=33580 345440 0 0 $X=33390 $Y=345200
X2413 1 2 591 44 611 ICV_37 $T=47840 329120 1 0 $X=47650 $Y=326160
X2414 1 2 602 45 615 ICV_37 $T=47840 367200 1 0 $X=47650 $Y=364240
X2415 1 2 602 70 607 ICV_37 $T=47840 378080 1 0 $X=47650 $Y=375120
X2416 1 2 627 14 647 ICV_37 $T=61640 334560 0 0 $X=61450 $Y=334320
X2417 1 2 627 15 648 ICV_37 $T=61640 345440 0 0 $X=61450 $Y=345200
X2418 1 2 602 40 641 ICV_37 $T=61640 367200 0 0 $X=61450 $Y=366960
X2419 1 2 602 35 640 ICV_37 $T=61640 372640 0 0 $X=61450 $Y=372400
X2420 1 2 83 45 674 ICV_37 $T=75900 367200 1 0 $X=75710 $Y=364240
X2421 1 2 687 43 700 ICV_37 $T=89700 329120 0 0 $X=89510 $Y=328880
X2422 1 2 694 25 703 ICV_37 $T=89700 350880 0 0 $X=89510 $Y=350640
X2423 1 2 720 25 712 ICV_37 $T=103960 334560 1 0 $X=103770 $Y=331600
X2424 1 2 720 14 733 ICV_37 $T=103960 340000 1 0 $X=103770 $Y=337040
X2425 1 2 732 43 752 ICV_37 $T=117760 323680 0 0 $X=117570 $Y=323440
X2426 1 2 744 13 770 ICV_37 $T=132020 350880 1 0 $X=131830 $Y=347920
X2427 1 2 744 42 778 ICV_37 $T=132020 356320 1 0 $X=131830 $Y=353360
X2428 1 2 786 44 801 ICV_37 $T=145820 340000 0 0 $X=145630 $Y=339760
X2429 1 2 785 44 797 ICV_37 $T=145820 356320 0 0 $X=145630 $Y=356080
X2430 1 2 195 177 860 ICV_37 $T=188140 372640 1 0 $X=187950 $Y=369680
X2431 1 2 882 189 909 ICV_37 $T=216200 323680 1 0 $X=216010 $Y=320720
X2432 1 2 882 191 916 ICV_37 $T=216200 334560 1 0 $X=216010 $Y=331600
X2433 1 2 214 175 915 ICV_37 $T=216200 378080 1 0 $X=216010 $Y=375120
X2434 1 2 914 171 941 ICV_37 $T=230000 329120 0 0 $X=229810 $Y=328880
X2435 1 2 913 171 934 ICV_37 $T=230000 350880 0 0 $X=229810 $Y=350640
X2436 1 2 907 163 942 ICV_37 $T=230000 367200 0 0 $X=229810 $Y=366960
X2437 1 2 950 187 966 ICV_37 $T=244260 329120 1 0 $X=244070 $Y=326160
X2438 1 2 165 55 224 ICV_37 $T=244260 361760 1 0 $X=244070 $Y=358800
X2439 1 2 995 187 1026 ICV_37 $T=272320 340000 1 0 $X=272130 $Y=337040
X2440 1 2 1008 158 1023 ICV_37 $T=272320 367200 1 0 $X=272130 $Y=364240
X2441 1 2 1035 190 1046 ICV_37 $T=286120 329120 0 0 $X=285930 $Y=328880
X2442 1 2 244 172 1066 ICV_37 $T=300380 318240 1 0 $X=300190 $Y=315280
X2443 1 2 1112 264 1126 ICV_37 $T=328440 345440 1 0 $X=328250 $Y=342480
X2444 1 2 278 262 1177 ICV_37 $T=356500 318240 1 0 $X=356310 $Y=315280
X2445 1 2 1169 266 1181 ICV_37 $T=356500 350880 1 0 $X=356310 $Y=347920
X2446 1 2 165 174 306 ICV_37 $T=356500 356320 1 0 $X=356310 $Y=353360
X2447 1 2 1146 264 1178 ICV_37 $T=356500 361760 1 0 $X=356310 $Y=358800
X2448 1 2 309 253 1207 ICV_37 $T=370300 312800 0 0 $X=370110 $Y=312560
X2449 1 2 309 264 1208 ICV_37 $T=370300 318240 0 0 $X=370110 $Y=318000
X2450 1 2 1187 273 1202 ICV_37 $T=370300 361760 0 0 $X=370110 $Y=361520
X2451 1 2 329 253 1263 ICV_37 $T=398360 367200 0 0 $X=398170 $Y=366960
X2452 1 2 1229 266 1281 ICV_37 $T=412620 329120 1 0 $X=412430 $Y=326160
X2453 1 2 1249 262 1288 ICV_37 $T=412620 345440 1 0 $X=412430 $Y=342480
X2454 1 2 329 260 1280 ICV_37 $T=412620 372640 1 0 $X=412430 $Y=369680
X2455 1 2 1301 262 1314 ICV_37 $T=426420 334560 0 0 $X=426230 $Y=334320
X2456 1 2 343 265 1309 ICV_37 $T=426420 367200 0 0 $X=426230 $Y=366960
X2457 1 2 1331 273 1366 ICV_37 $T=454480 323680 0 0 $X=454290 $Y=323440
X2458 1 2 1331 260 1368 ICV_37 $T=454480 329120 0 0 $X=454290 $Y=328880
X2459 1 2 365 266 1402 ICV_37 $T=468740 318240 1 0 $X=468550 $Y=315280
X2460 1 2 1378 253 1401 ICV_37 $T=468740 323680 1 0 $X=468550 $Y=320720
X2461 1 2 1385 273 1404 ICV_37 $T=468740 372640 1 0 $X=468550 $Y=369680
X2462 1 2 1431 253 1487 ICV_37 $T=510600 350880 0 0 $X=510410 $Y=350640
X2463 1 2 1551 412 1556 ICV_37 $T=552920 356320 1 0 $X=552730 $Y=353360
X2464 1 2 431 400 1541 ICV_37 $T=552920 378080 1 0 $X=552730 $Y=375120
X2465 1 2 1574 397 1586 ICV_37 $T=566720 323680 0 0 $X=566530 $Y=323440
X2466 1 2 1574 399 1587 ICV_37 $T=566720 334560 0 0 $X=566530 $Y=334320
X2467 1 2 1575 414 1589 ICV_37 $T=566720 340000 0 0 $X=566530 $Y=339760
X2468 1 2 1574 415 1609 ICV_37 $T=580980 329120 1 0 $X=580790 $Y=326160
X2469 1 2 1602 400 1617 ICV_37 $T=580980 361760 1 0 $X=580790 $Y=358800
X2470 1 2 1602 414 1621 ICV_37 $T=580980 367200 1 0 $X=580790 $Y=364240
X2471 1 2 434 410 436 ICV_37 $T=580980 378080 1 0 $X=580790 $Y=375120
X2472 1 2 1602 398 1639 ICV_37 $T=594780 361760 0 0 $X=594590 $Y=361520
X2473 1 2 1655 412 1673 ICV_37 $T=609040 372640 1 0 $X=608850 $Y=369680
X2474 1 2 441 400 442 ICV_37 $T=609040 378080 1 0 $X=608850 $Y=375120
X2475 1 2 1663 414 1701 ICV_37 $T=622840 329120 0 0 $X=622650 $Y=328880
X2476 1 2 1712 397 1754 ICV_37 $T=650900 323680 0 0 $X=650710 $Y=323440
X2477 1 2 1713 400 1748 ICV_37 $T=650900 350880 0 0 $X=650710 $Y=350640
X2478 1 2 1779 414 1807 ICV_37 $T=678960 345440 0 0 $X=678770 $Y=345200
X2479 1 2 1801 400 1837 ICV_37 $T=693220 318240 1 0 $X=693030 $Y=315280
X2480 1 2 1801 399 1831 ICV_37 $T=693220 323680 1 0 $X=693030 $Y=320720
X2481 1 2 1775 415 1839 ICV_37 $T=693220 329120 1 0 $X=693030 $Y=326160
X2482 1 2 457 400 1844 ICV_37 $T=693220 378080 1 0 $X=693030 $Y=375120
X2483 1 2 466 400 1865 ICV_37 $T=707020 318240 0 0 $X=706830 $Y=318000
X2484 1 2 608 18 620 608 15 638 ICV_38 $T=49680 356320 1 0 $X=49490 $Y=353360
X2485 1 2 637 15 651 637 42 667 ICV_38 $T=63940 329120 0 0 $X=63750 $Y=328880
X2486 1 2 687 13 723 687 15 727 ICV_38 $T=98440 318240 0 0 $X=98250 $Y=318000
X2487 1 2 720 42 730 720 15 738 ICV_38 $T=104420 345440 1 0 $X=104230 $Y=342480
X2488 1 2 118 18 768 772 43 787 ICV_38 $T=131100 318240 0 0 $X=130910 $Y=318000
X2489 1 2 800 163 828 800 177 838 ICV_38 $T=162380 372640 1 0 $X=162190 $Y=369680
X2490 1 2 913 168 927 913 170 933 ICV_38 $T=222180 340000 1 0 $X=221990 $Y=337040
X2491 1 2 950 168 967 950 171 980 ICV_38 $T=243340 323680 0 0 $X=243150 $Y=323440
X2492 1 2 223 189 978 223 191 979 ICV_38 $T=248400 318240 1 0 $X=248210 $Y=315280
X2493 1 2 995 189 1019 995 191 1002 ICV_38 $T=268640 345440 0 0 $X=268450 $Y=345200
X2494 1 2 1022 152 1049 1008 152 1065 ICV_38 $T=285660 372640 1 0 $X=285470 $Y=369680
X2495 1 2 1035 170 1069 1035 187 1085 ICV_38 $T=295780 323680 0 0 $X=295590 $Y=323440
X2496 1 2 1073 191 1086 1073 189 1100 ICV_38 $T=303600 334560 1 0 $X=303410 $Y=331600
X2497 1 2 1102 260 1121 1102 273 1127 ICV_38 $T=323840 350880 0 0 $X=323650 $Y=350640
X2498 1 2 1102 266 1119 1102 265 1134 ICV_38 $T=324300 345440 0 0 $X=324110 $Y=345200
X2499 1 2 1112 265 1125 1112 253 1141 ICV_38 $T=327060 334560 0 0 $X=326870 $Y=334320
X2500 1 2 1118 257 1151 1118 264 1167 ICV_38 $T=339020 329120 1 0 $X=338830 $Y=326160
X2501 1 2 1146 262 1153 1146 257 1170 ICV_38 $T=341780 361760 1 0 $X=341590 $Y=358800
X2502 1 2 1169 257 1179 1169 265 1192 ICV_38 $T=355580 340000 0 0 $X=355390 $Y=339760
X2503 1 2 1171 273 1184 1171 266 1197 ICV_38 $T=358800 323680 1 0 $X=358610 $Y=320720
X2504 1 2 1203 260 1228 1203 265 1241 ICV_38 $T=382720 334560 0 0 $X=382530 $Y=334320
X2505 1 2 1230 264 1226 1257 260 1269 ICV_38 $T=394680 356320 1 0 $X=394490 $Y=353360
X2506 1 2 1284 253 1304 1284 264 1293 ICV_38 $T=420440 329120 1 0 $X=420250 $Y=326160
X2507 1 2 1301 264 1317 1301 265 1333 ICV_38 $T=428260 345440 0 0 $X=428070 $Y=345200
X2508 1 2 1294 265 1341 1339 266 1359 ICV_38 $T=439300 356320 0 0 $X=439110 $Y=356080
X2509 1 2 1384 265 1398 1384 264 1410 ICV_38 $T=466440 350880 0 0 $X=466250 $Y=350640
X2510 1 2 1360 257 1409 1413 264 1427 ICV_38 $T=471960 345440 1 0 $X=471770 $Y=342480
X2511 1 2 1429 266 1462 1429 257 1477 ICV_38 $T=499100 367200 1 0 $X=498910 $Y=364240
X2512 1 2 1484 412 1525 1484 415 1535 ICV_38 $T=533600 323680 1 0 $X=533410 $Y=320720
X2513 1 2 1540 400 1554 1540 397 1570 ICV_38 $T=549240 367200 0 0 $X=549050 $Y=366960
X2514 1 2 1527 412 1555 1527 399 1564 ICV_38 $T=549700 345440 0 0 $X=549510 $Y=345200
X2515 1 2 1540 412 1581 1540 415 1579 ICV_38 $T=565800 372640 1 0 $X=565610 $Y=369680
X2516 1 2 1575 415 1583 1575 399 1605 ICV_38 $T=566260 350880 1 0 $X=566070 $Y=347920
X2517 1 2 1602 399 1638 1602 410 1644 ICV_38 $T=590640 367200 1 0 $X=590450 $Y=364240
X2518 1 2 1655 400 1670 1655 410 1666 ICV_38 $T=605820 361760 0 0 $X=605630 $Y=361520
X2519 1 2 1652 414 1684 1652 400 1696 ICV_38 $T=613180 350880 1 0 $X=612990 $Y=347920
X2520 1 2 441 414 443 441 410 1693 ICV_38 $T=616860 378080 1 0 $X=616670 $Y=375120
X2521 1 2 1713 412 1727 1713 410 1742 ICV_38 $T=636180 345440 0 0 $X=635990 $Y=345200
X2522 1 2 1720 397 1750 1720 410 1773 ICV_38 $T=651360 340000 0 0 $X=651170 $Y=339760
X2523 1 2 1850 400 1864 1850 414 1883 ICV_38 $T=703340 323680 1 0 $X=703150 $Y=320720
X2524 1 2 467 400 1870 467 398 1893 ICV_38 $T=708400 372640 0 0 $X=708210 $Y=372400
X2525 1 2 76 77 38 ICV_40 $T=54280 372640 0 0 $X=54090 $Y=372400
X2526 1 2 639 609 38 ICV_40 $T=69920 372640 1 0 $X=69730 $Y=369680
X2527 1 2 677 653 57 ICV_40 $T=83720 323680 0 0 $X=83530 $Y=323440
X2528 1 2 663 645 28 ICV_40 $T=83720 340000 0 0 $X=83530 $Y=339760
X2529 1 2 743 713 34 ICV_40 $T=118680 334560 0 0 $X=118490 $Y=334320
X2530 1 2 812 821 176 ICV_40 $T=167440 372640 0 0 $X=167250 $Y=372400
X2531 1 2 252 245 166 ICV_40 $T=308200 312800 0 0 $X=308010 $Y=312560
X2532 1 2 1084 1076 201 ICV_40 $T=308200 350880 0 0 $X=308010 $Y=350640
X2533 1 2 1119 1120 275 ICV_40 $T=329360 350880 1 0 $X=329170 $Y=347920
X2534 1 2 1121 1120 267 ICV_40 $T=329820 356320 1 0 $X=329630 $Y=353360
X2535 1 2 1127 1120 280 ICV_40 $T=335340 350880 1 0 $X=335150 $Y=347920
X2536 1 2 1113 254 166 ICV_40 $T=335800 312800 0 0 $X=335610 $Y=312560
X2537 1 2 294 284 277 ICV_40 $T=350520 378080 1 0 $X=350330 $Y=375120
X2538 1 2 1162 1131 269 ICV_40 $T=356960 334560 0 0 $X=356770 $Y=334320
X2539 1 2 1176 289 268 ICV_40 $T=364320 318240 0 0 $X=364130 $Y=318000
X2540 1 2 1190 1186 263 ICV_40 $T=371220 329120 1 0 $X=371030 $Y=326160
X2541 1 2 1200 1188 277 ICV_40 $T=378580 361760 1 0 $X=378390 $Y=358800
X2542 1 2 1311 1313 268 ICV_40 $T=432400 340000 0 0 $X=432210 $Y=339760
X2543 1 2 1358 1356 269 ICV_40 $T=453560 350880 1 0 $X=453370 $Y=347920
X2544 1 2 1367 1350 263 ICV_40 $T=462760 329120 1 0 $X=462570 $Y=326160
X2545 1 2 1365 358 268 ICV_40 $T=462760 378080 1 0 $X=462570 $Y=375120
X2546 1 2 1393 1371 269 ICV_40 $T=470120 329120 1 0 $X=469930 $Y=326160
X2547 1 2 1446 1425 267 ICV_40 $T=496800 323680 0 0 $X=496610 $Y=323440
X2548 1 2 1495 1503 405 ICV_40 $T=525780 345440 1 0 $X=525590 $Y=342480
X2549 1 2 1561 426 408 ICV_40 $T=560740 372640 0 0 $X=560550 $Y=372400
X2550 1 2 1667 1665 418 ICV_40 $T=616400 350880 0 0 $X=616210 $Y=350640
X2551 1 2 1724 450 405 ICV_40 $T=644920 372640 0 0 $X=644730 $Y=372400
X2552 1 2 1777 1780 405 ICV_40 $T=666540 356320 1 0 $X=666350 $Y=353360
X2553 1 2 1784 455 405 ICV_40 $T=672520 372640 0 0 $X=672330 $Y=372400
X2554 1 2 1893 468 405 ICV_40 $T=736920 372640 1 0 $X=736730 $Y=369680
X2555 1 2 580 43 600 ICV_41 $T=37720 345440 1 0 $X=37530 $Y=342480
X2556 1 2 644 14 678 ICV_41 $T=79580 350880 0 0 $X=79390 $Y=350640
X2557 1 2 94 44 99 ICV_41 $T=90160 312800 0 0 $X=89970 $Y=312560
X2558 1 2 825 190 845 ICV_41 $T=178020 329120 1 0 $X=177830 $Y=326160
X2559 1 2 855 187 866 ICV_41 $T=191820 334560 0 0 $X=191630 $Y=334320
X2560 1 2 859 156 895 ICV_41 $T=206080 367200 1 0 $X=205890 $Y=364240
X2561 1 2 950 190 965 ICV_41 $T=240580 329120 0 0 $X=240390 $Y=328880
X2562 1 2 1073 190 1110 ICV_41 $T=318320 334560 1 0 $X=318130 $Y=331600
X2563 1 2 325 262 1270 ICV_41 $T=402500 318240 1 0 $X=402310 $Y=315280
X2564 1 2 356 273 1351 ICV_41 $T=443900 312800 0 0 $X=443710 $Y=312560
X2565 1 2 356 264 1352 ICV_41 $T=443900 318240 0 0 $X=443710 $Y=318000
X2566 1 2 1360 253 1373 ICV_41 $T=454940 340000 0 0 $X=454750 $Y=339760
X2567 1 2 1413 266 1435 ICV_41 $T=486680 345440 1 0 $X=486490 $Y=342480
X2568 1 2 1430 257 1463 ICV_41 $T=500020 318240 0 0 $X=499830 $Y=318000
X2569 1 2 1578 410 1598 ICV_41 $T=570860 318240 1 0 $X=570670 $Y=315280
X2570 1 2 1801 397 1815 ICV_41 $T=679420 323680 0 0 $X=679230 $Y=323440
X2571 1 2 1859 410 1910 ICV_41 $T=724960 334560 0 0 $X=724770 $Y=334320
X2572 1 2 9 10 536 ICV_47 $T=5520 367200 0 0 $X=5330 $Y=366960
X2573 1 2 48 45 598 ICV_47 $T=36340 367200 0 0 $X=36150 $Y=366960
X2574 1 2 591 18 71 ICV_47 $T=41400 323680 0 0 $X=41210 $Y=323440
X2575 1 2 580 15 619 ICV_47 $T=48300 345440 1 0 $X=48110 $Y=342480
X2576 1 2 608 42 629 ICV_47 $T=52440 361760 1 0 $X=52250 $Y=358800
X2577 1 2 637 14 654 ICV_47 $T=64400 329120 1 0 $X=64210 $Y=326160
X2578 1 2 627 42 660 ICV_47 $T=67160 345440 1 0 $X=66970 $Y=342480
X2579 1 2 672 44 689 ICV_47 $T=80500 345440 1 0 $X=80310 $Y=342480
X2580 1 2 98 45 717 ICV_47 $T=93380 367200 1 0 $X=93190 $Y=364240
X2581 1 2 687 14 721 ICV_47 $T=95220 329120 1 0 $X=95030 $Y=326160
X2582 1 2 732 18 764 ICV_47 $T=123280 323680 1 0 $X=123090 $Y=320720
X2583 1 2 785 18 808 ICV_47 $T=149960 350880 1 0 $X=149770 $Y=347920
X2584 1 2 800 152 812 ICV_47 $T=151340 372640 1 0 $X=151150 $Y=369680
X2585 1 2 786 25 816 ICV_47 $T=153640 329120 0 0 $X=153450 $Y=328880
X2586 1 2 853 187 861 ICV_47 $T=188600 329120 1 0 $X=188410 $Y=326160
X2587 1 2 855 170 867 ICV_47 $T=190440 340000 0 0 $X=190250 $Y=339760
X2588 1 2 208 187 209 ICV_47 $T=202400 312800 0 0 $X=202210 $Y=312560
X2589 1 2 884 189 894 ICV_47 $T=204700 345440 1 0 $X=204510 $Y=342480
X2590 1 2 884 171 900 ICV_47 $T=205620 356320 1 0 $X=205430 $Y=353360
X2591 1 2 913 190 931 ICV_47 $T=221260 350880 0 0 $X=221070 $Y=350640
X2592 1 2 939 191 952 ICV_47 $T=234600 350880 1 0 $X=234410 $Y=347920
X2593 1 2 165 59 226 ICV_47 $T=246560 356320 0 0 $X=246370 $Y=356080
X2594 1 2 968 187 982 ICV_47 $T=249320 340000 0 0 $X=249130 $Y=339760
X2595 1 2 995 170 1017 ICV_47 $T=265880 334560 0 0 $X=265690 $Y=334320
X2596 1 2 1073 172 1087 ICV_47 $T=304980 329120 1 0 $X=304790 $Y=326160
X2597 1 2 1095 260 1105 ICV_47 $T=314640 361760 0 0 $X=314450 $Y=361520
X2598 1 2 250 191 1114 ICV_47 $T=317400 318240 1 0 $X=317210 $Y=315280
X2599 1 2 250 168 1115 ICV_47 $T=317860 323680 1 0 $X=317670 $Y=320720
X2600 1 2 1118 265 1133 ICV_47 $T=328900 334560 1 0 $X=328710 $Y=331600
X2601 1 2 1171 262 1183 ICV_47 $T=356960 334560 1 0 $X=356770 $Y=331600
X2602 1 2 312 265 320 ICV_47 $T=373520 378080 1 0 $X=373330 $Y=375120
X2603 1 2 1205 264 1238 ICV_47 $T=389160 350880 0 0 $X=388970 $Y=350640
X2604 1 2 1229 264 1244 ICV_47 $T=389620 323680 0 0 $X=389430 $Y=323440
X2605 1 2 1257 273 1271 ICV_47 $T=401580 350880 1 0 $X=401390 $Y=347920
X2606 1 2 1331 264 1344 ICV_47 $T=441140 334560 1 0 $X=440950 $Y=331600
X2607 1 2 1360 273 1412 ICV_47 $T=471040 334560 0 0 $X=470850 $Y=334320
X2608 1 2 1385 264 1421 ICV_47 $T=476560 372640 1 0 $X=476370 $Y=369680
X2609 1 2 1385 253 1424 ICV_47 $T=477020 367200 1 0 $X=476830 $Y=364240
X2610 1 2 1431 264 1451 ICV_47 $T=488060 356320 1 0 $X=487870 $Y=353360
X2611 1 2 1431 257 1472 ICV_47 $T=501860 350880 0 0 $X=501670 $Y=350640
X2612 1 2 1430 253 1482 ICV_47 $T=505540 323680 1 0 $X=505350 $Y=320720
X2613 1 2 1484 397 1492 ICV_47 $T=516120 318240 1 0 $X=515930 $Y=315280
X2614 1 2 1486 398 1495 ICV_47 $T=516120 345440 1 0 $X=515930 $Y=342480
X2615 1 2 1486 397 1504 ICV_47 $T=518420 350880 0 0 $X=518230 $Y=350640
X2616 1 2 1485 415 1520 ICV_47 $T=530380 334560 1 0 $X=530190 $Y=331600
X2617 1 2 1540 399 1561 ICV_47 $T=553380 372640 1 0 $X=553190 $Y=369680
X2618 1 2 1529 410 1568 ICV_47 $T=554760 334560 1 0 $X=554570 $Y=331600
X2619 1 2 1527 415 1550 ICV_47 $T=555220 340000 0 0 $X=555030 $Y=339760
X2620 1 2 434 412 1623 ICV_47 $T=581440 372640 1 0 $X=581250 $Y=369680
X2621 1 2 1612 398 1625 ICV_47 $T=583740 356320 1 0 $X=583550 $Y=353360
X2622 1 2 1618 412 1654 ICV_47 $T=597080 340000 1 0 $X=596890 $Y=337040
X2623 1 2 1640 399 1657 ICV_47 $T=598460 323680 1 0 $X=598270 $Y=320720
X2624 1 2 1652 415 1667 ICV_47 $T=603980 356320 0 0 $X=603790 $Y=356080
X2625 1 2 1652 399 1686 ICV_47 $T=614100 356320 0 0 $X=613910 $Y=356080
X2626 1 2 454 415 1772 ICV_47 $T=656420 372640 1 0 $X=656230 $Y=369680
X2627 1 2 454 398 1784 ICV_47 $T=662860 372640 0 0 $X=662670 $Y=372400
X2628 1 2 454 414 1800 ICV_47 $T=670220 367200 0 0 $X=670030 $Y=366960
X2629 1 2 1808 410 1829 ICV_47 $T=684480 350880 1 0 $X=684290 $Y=347920
X2630 1 2 1814 414 1833 ICV_47 $T=686780 345440 0 0 $X=686590 $Y=345200
X2631 1 2 1859 398 1890 ICV_47 $T=709780 340000 1 0 $X=709590 $Y=337040
X2632 1 2 467 412 1907 ICV_47 $T=723120 372640 0 0 $X=722930 $Y=372400
X2633 1 2 1862 412 1915 ICV_47 $T=724500 367200 0 0 $X=724310 $Y=366960
X2634 1 2 598 53 47 ICV_48 $T=43700 372640 1 0 $X=43510 $Y=369680
X2635 1 2 84 77 75 ICV_48 $T=71760 378080 1 0 $X=71570 $Y=375120
X2636 1 2 781 783 39 ICV_48 $T=141680 329120 0 0 $X=141490 $Y=328880
X2637 1 2 808 741 37 ICV_48 $T=155940 378080 1 0 $X=155750 $Y=375120
X2638 1 2 816 783 28 ICV_48 $T=169740 345440 0 0 $X=169550 $Y=345200
X2639 1 2 841 830 197 ICV_48 $T=184000 318240 1 0 $X=183810 $Y=315280
X2640 1 2 843 820 198 ICV_48 $T=184000 345440 1 0 $X=183810 $Y=342480
X2641 1 2 976 958 166 ICV_48 $T=253920 334560 0 0 $X=253730 $Y=334320
X2642 1 2 1002 1004 198 ICV_48 $T=268180 345440 1 0 $X=267990 $Y=342480
X2643 1 2 1003 1004 179 ICV_48 $T=268180 350880 1 0 $X=267990 $Y=347920
X2644 1 2 1041 1047 198 ICV_48 $T=296240 323680 1 0 $X=296050 $Y=320720
X2645 1 2 1087 1083 186 ICV_48 $T=310040 334560 0 0 $X=309850 $Y=334320
X2646 1 2 1109 261 269 ICV_48 $T=324300 378080 1 0 $X=324110 $Y=375120
X2647 1 2 1150 1120 296 ICV_48 $T=352360 345440 1 0 $X=352170 $Y=342480
X2648 1 2 1184 1186 280 ICV_48 $T=366160 323680 0 0 $X=365970 $Y=323440
X2649 1 2 1267 1250 263 ICV_48 $T=408480 323680 1 0 $X=408290 $Y=320720
X2650 1 2 1268 1256 267 ICV_48 $T=408480 340000 1 0 $X=408290 $Y=337040
X2651 1 2 1293 1295 296 ICV_48 $T=422280 323680 0 0 $X=422090 $Y=323440
X2652 1 2 1322 1295 277 ICV_48 $T=436540 329120 1 0 $X=436350 $Y=326160
X2653 1 2 1324 1306 263 ICV_48 $T=436540 367200 1 0 $X=436350 $Y=364240
X2654 1 2 1381 1382 269 ICV_48 $T=464600 334560 1 0 $X=464410 $Y=331600
X2655 1 2 1513 1507 417 ICV_48 $T=534520 323680 0 0 $X=534330 $Y=323440
X2656 1 2 1515 1509 407 ICV_48 $T=534520 356320 0 0 $X=534330 $Y=356080
X2657 1 2 1538 1543 405 ICV_48 $T=548780 334560 1 0 $X=548590 $Y=331600
X2658 1 2 1539 1543 417 ICV_48 $T=548780 350880 1 0 $X=548590 $Y=347920
X2659 1 2 428 429 408 ICV_48 $T=548780 372640 1 0 $X=548590 $Y=369680
X2660 1 2 1653 1633 417 ICV_48 $T=604900 329120 1 0 $X=604710 $Y=326160
X2661 1 2 1702 1668 418 ICV_48 $T=632960 361760 1 0 $X=632770 $Y=358800
X2662 1 2 1792 1797 409 ICV_48 $T=674820 334560 0 0 $X=674630 $Y=334320
X2663 1 2 1794 1797 417 ICV_48 $T=674820 350880 0 0 $X=674630 $Y=350640
X2664 1 2 1822 1818 405 ICV_48 $T=689080 367200 1 0 $X=688890 $Y=364240
X2665 1 2 1851 1827 409 ICV_48 $T=702880 340000 0 0 $X=702690 $Y=339760
X2666 1 2 580 13 592 592 596 34 ICV_49 $T=32660 340000 1 0 $X=32470 $Y=337040
X2667 1 2 637 13 652 652 653 34 ICV_49 $T=62100 318240 0 0 $X=61910 $Y=318000
X2668 1 2 1061 189 1081 1081 1076 199 ICV_49 $T=298080 345440 0 0 $X=297890 $Y=345200
X2669 1 2 1095 273 1139 1139 261 280 ICV_49 $T=328900 367200 1 0 $X=328710 $Y=364240
X2670 1 2 1112 262 1162 1145 1131 267 ICV_49 $T=342240 340000 1 0 $X=342050 $Y=337040
X2671 1 2 1187 265 1200 1202 1188 280 ICV_49 $T=364320 361760 1 0 $X=364130 $Y=358800
X2672 1 2 1230 260 1248 1248 1227 267 ICV_49 $T=389160 361760 1 0 $X=388970 $Y=358800
X2673 1 2 365 260 1396 1396 371 267 ICV_49 $T=463680 312800 0 0 $X=463490 $Y=312560
X2674 1 2 1360 265 1411 1408 1371 267 ICV_49 $T=469200 340000 1 0 $X=469010 $Y=337040
X2675 1 2 1529 397 1562 1548 1542 424 ICV_49 $T=552460 323680 0 0 $X=552270 $Y=323440
X2676 1 2 1527 398 1538 1563 1542 418 ICV_49 $T=553380 340000 1 0 $X=553190 $Y=337040
X2677 1 2 1661 399 1683 1683 1678 408 ICV_49 $T=609500 340000 1 0 $X=609310 $Y=337040
X2678 1 2 1808 400 1821 1809 1797 418 ICV_49 $T=679420 350880 0 0 $X=679230 $Y=350640
X2679 1 2 1860 398 1867 1867 1871 405 ICV_49 $T=705180 356320 1 0 $X=704990 $Y=353360
X2680 1 2 1850 398 1879 1883 1869 422 ICV_49 $T=707480 323680 0 0 $X=707290 $Y=323440
X2681 1 2 1861 398 1880 1832 1827 417 ICV_49 $T=707480 340000 0 0 $X=707290 $Y=339760
X2682 1 2 1861 410 1904 1880 1891 405 ICV_49 $T=721740 345440 1 0 $X=721550 $Y=342480
X2683 1 2 1861 399 1906 1874 1891 407 ICV_49 $T=721740 350880 1 0 $X=721550 $Y=347920
X2684 1 2 687 18 702 702 699 37 ICV_50 $T=85560 323680 1 0 $X=85370 $Y=320720
X2685 1 2 750 43 762 749 713 37 ICV_50 $T=118220 340000 0 0 $X=118030 $Y=339760
X2686 1 2 744 43 777 778 759 54 ICV_50 $T=128340 356320 0 0 $X=128150 $Y=356080
X2687 1 2 825 187 841 845 830 201 ICV_50 $T=174340 318240 0 0 $X=174150 $Y=318000
X2688 1 2 907 158 918 918 924 180 ICV_50 $T=214820 361760 0 0 $X=214630 $Y=361520
X2689 1 2 907 156 940 940 924 167 ICV_50 $T=225860 367200 1 0 $X=225670 $Y=364240
X2690 1 2 1030 191 1056 1056 1039 198 ICV_50 $T=284280 345440 1 0 $X=284090 $Y=342480
X2691 1 2 309 266 1201 313 315 277 ICV_50 $T=364320 318240 1 0 $X=364130 $Y=315280
X2692 1 2 1294 266 1316 1317 1313 296 ICV_50 $T=423660 350880 1 0 $X=423470 $Y=347920
X2693 1 2 1339 253 1383 1357 1356 268 ICV_50 $T=454940 345440 0 0 $X=454750 $Y=345200
X2694 1 2 1428 257 1478 1478 1450 268 ICV_50 $T=501400 334560 1 0 $X=501210 $Y=331600
X2695 1 2 1486 399 1497 1497 1503 408 ICV_50 $T=515200 340000 0 0 $X=515010 $Y=339760
X2696 1 2 1496 415 1533 1517 1509 409 ICV_50 $T=536360 361760 1 0 $X=536170 $Y=358800
X2697 1 2 427 397 1571 1572 430 405 ICV_50 $T=553380 318240 1 0 $X=553190 $Y=315280
X2698 1 2 1661 410 1674 1674 1678 417 ICV_50 $T=606280 334560 0 0 $X=606090 $Y=334320
X2699 1 2 457 397 1823 458 459 417 ICV_50 $T=679420 372640 0 0 $X=679230 $Y=372400
X2700 1 2 1814 399 1855 1855 1827 408 ICV_50 $T=693680 345440 1 0 $X=693490 $Y=342480
X2701 1 2 1862 399 1913 1913 1881 408 ICV_50 $T=721740 372640 1 0 $X=721550 $Y=369680
X2702 1 2 535 27 33 9 35 555 ICV_51 $T=12420 372640 0 0 $X=12230 $Y=372400
X2703 1 2 571 53 59 48 10 582 ICV_51 $T=28520 372640 1 0 $X=28330 $Y=369680
X2704 1 2 61 53 63 48 35 67 ICV_51 $T=33580 378080 1 0 $X=33390 $Y=375120
X2705 1 2 611 72 57 591 15 632 ICV_51 $T=50140 329120 0 0 $X=49950 $Y=328880
X2706 1 2 95 97 75 98 35 715 ICV_51 $T=90160 378080 1 0 $X=89970 $Y=375120
X2707 1 2 738 713 39 744 25 754 ICV_51 $T=115000 350880 1 0 $X=114810 $Y=347920
X2708 1 2 790 791 57 772 18 809 ICV_51 $T=146740 323680 0 0 $X=146550 $Y=323440
X2709 1 2 819 820 166 826 168 835 ICV_51 $T=162840 334560 1 0 $X=162650 $Y=331600
X2710 1 2 851 852 198 855 189 872 ICV_51 $T=188140 345440 0 0 $X=187950 $Y=345200
X2711 1 2 903 868 180 165 63 220 ICV_51 $T=213900 356320 0 0 $X=213710 $Y=356080
X2712 1 2 909 887 199 914 190 929 ICV_51 $T=218500 323680 0 0 $X=218310 $Y=323440
X2713 1 2 956 958 198 223 190 977 ICV_51 $T=243800 318240 0 0 $X=243610 $Y=318000
X2714 1 2 229 230 185 234 181 1009 ICV_51 $T=260820 378080 1 0 $X=260630 $Y=375120
X2715 1 2 1101 261 263 1079 163 1117 ICV_51 $T=317400 367200 0 0 $X=317210 $Y=366960
X2716 1 2 1226 1227 296 1230 273 1246 ICV_51 $T=386860 356320 0 0 $X=386670 $Y=356080
X2717 1 2 1246 1227 280 1257 253 1273 ICV_51 $T=399740 356320 0 0 $X=399550 $Y=356080
X2718 1 2 1255 1256 296 1249 260 1268 ICV_51 $T=400660 340000 0 0 $X=400470 $Y=339760
X2719 1 2 1280 333 267 343 257 1302 ICV_51 $T=414920 367200 0 0 $X=414730 $Y=366960
X2720 1 2 1285 1261 296 1294 262 1310 ICV_51 $T=421360 356320 1 0 $X=421170 $Y=353360
X2721 1 2 1333 1313 277 1339 264 1353 ICV_51 $T=442060 345440 1 0 $X=441870 $Y=342480
X2722 1 2 1369 1371 296 1360 262 1393 ICV_51 $T=459540 334560 0 0 $X=459350 $Y=334320
X2723 1 2 1411 1371 277 1428 264 1439 ICV_51 $T=483460 340000 1 0 $X=483270 $Y=337040
X2724 1 2 1422 371 296 1430 264 1423 ICV_51 $T=484840 318240 0 0 $X=484650 $Y=318000
X2725 1 2 1423 1425 296 1430 260 1446 ICV_51 $T=484840 329120 1 0 $X=484650 $Y=326160
X2726 1 2 1426 1400 280 1431 262 1453 ICV_51 $T=485300 361760 1 0 $X=485110 $Y=358800
X2727 1 2 1603 1585 417 1612 414 1624 ICV_51 $T=579600 345440 0 0 $X=579410 $Y=345200
X2728 1 2 1610 1580 407 1618 399 1631 ICV_51 $T=583280 329120 0 0 $X=583090 $Y=328880
X2729 1 2 1611 1580 405 1618 397 1632 ICV_51 $T=583280 340000 1 0 $X=583090 $Y=337040
X2730 1 2 1666 1668 417 1655 398 1687 ICV_51 $T=611340 372640 0 0 $X=611150 $Y=372400
X2731 1 2 1695 1682 417 446 397 1718 ICV_51 $T=626980 318240 0 0 $X=626790 $Y=318000
X2732 1 2 1739 1740 418 1720 412 1766 ICV_51 $T=650440 340000 1 0 $X=650250 $Y=337040
X2733 1 2 1748 1722 407 1756 415 1771 ICV_51 $T=653660 356320 1 0 $X=653470 $Y=353360
X2734 1 2 1782 1781 405 1775 400 1803 ICV_51 $T=668840 334560 1 0 $X=668650 $Y=331600
X2735 1 2 1807 1797 422 1814 400 1828 ICV_51 $T=681720 345440 1 0 $X=681530 $Y=342480
X2736 1 2 1811 456 417 1801 415 463 ICV_51 $T=684940 312800 0 0 $X=684750 $Y=312560
X2737 1 2 1873 469 409 466 399 1908 ICV_51 $T=720820 312800 0 0 $X=720630 $Y=312560
X2738 1 2 555 27 49 ICV_52 $T=23000 372640 1 0 $X=22810 $Y=369680
X2739 1 2 890 887 197 ICV_52 $T=210680 329120 1 0 $X=210490 $Y=326160
X2740 1 2 947 219 166 ICV_52 $T=238740 318240 1 0 $X=238550 $Y=315280
X2741 1 2 1025 1010 201 ICV_52 $T=279220 323680 1 0 $X=279030 $Y=320720
X2742 1 2 1069 1047 166 ICV_52 $T=301760 323680 1 0 $X=301570 $Y=320720
X2743 1 2 1134 1120 277 ICV_52 $T=336720 340000 0 0 $X=336530 $Y=339760
X2744 1 2 1443 1434 269 ICV_52 $T=500480 367200 0 0 $X=500290 $Y=366960
X2745 1 2 1501 1506 408 ICV_52 $T=526240 329120 1 0 $X=526050 $Y=326160
X2746 1 2 1553 1542 405 ICV_52 $T=553840 334560 0 0 $X=553650 $Y=334320
X2747 1 2 1564 1543 408 ICV_52 $T=561660 345440 1 0 $X=561470 $Y=342480
X2748 1 2 1566 1557 409 ICV_52 $T=567640 367200 1 0 $X=567450 $Y=364240
X2749 1 2 1679 1682 418 ICV_52 $T=618240 329120 1 0 $X=618050 $Y=326160
X2750 1 2 1710 445 405 ICV_52 $T=632960 312800 0 0 $X=632770 $Y=312560
X2751 1 2 1733 445 408 ICV_52 $T=645380 312800 0 0 $X=645190 $Y=312560
X2752 1 2 1742 1722 417 ICV_52 $T=648600 345440 1 0 $X=648410 $Y=342480
X2753 1 2 1768 1749 418 ICV_52 $T=667000 312800 0 0 $X=666810 $Y=312560
X2754 1 2 1823 462 409 ICV_52 $T=694600 372640 0 0 $X=694410 $Y=372400
X2755 1 2 718 100 63 ICV_53 $T=102120 372640 0 0 $X=101930 $Y=372400
X2756 1 2 761 759 37 ICV_53 $T=126500 350880 1 0 $X=126310 $Y=347920
X2757 1 2 769 747 34 ICV_53 $T=132480 329120 1 0 $X=132290 $Y=326160
X2758 1 2 817 783 34 ICV_53 $T=160540 350880 1 0 $X=160350 $Y=347920
X2759 1 2 863 868 185 ICV_53 $T=196420 367200 0 0 $X=196230 $Y=366960
X2760 1 2 871 854 179 ICV_53 $T=197340 329120 1 0 $X=197150 $Y=326160
X2761 1 2 892 888 198 ICV_53 $T=210680 350880 1 0 $X=210490 $Y=347920
X2762 1 2 973 975 188 ICV_53 $T=252080 361760 1 0 $X=251890 $Y=358800
X2763 1 2 989 987 201 ICV_53 $T=258520 350880 0 0 $X=258330 $Y=350640
X2764 1 2 1174 1158 267 ICV_53 $T=356960 367200 1 0 $X=356770 $Y=364240
X2765 1 2 1185 1188 296 ICV_53 $T=364780 361760 0 0 $X=364590 $Y=361520
X2766 1 2 1196 1173 269 ICV_53 $T=370760 340000 0 0 $X=370570 $Y=339760
X2767 1 2 1316 1308 275 ICV_53 $T=432860 356320 1 0 $X=432670 $Y=353360
X2768 1 2 1418 1400 267 ICV_53 $T=483000 356320 0 0 $X=482810 $Y=356080
X2769 1 2 1499 1507 407 ICV_53 $T=525320 318240 1 0 $X=525130 $Y=315280
X2770 1 2 1504 1503 409 ICV_53 $T=525320 350880 1 0 $X=525130 $Y=347920
X2771 1 2 1525 1507 424 ICV_53 $T=539120 323680 0 0 $X=538930 $Y=323440
X2772 1 2 1541 429 407 ICV_53 $T=547400 378080 1 0 $X=547210 $Y=375120
X2773 1 2 1609 1580 418 ICV_53 $T=581440 323680 1 0 $X=581250 $Y=320720
X2774 1 2 1693 444 417 ICV_53 $T=623300 372640 0 0 $X=623110 $Y=372400
X2775 1 2 1700 1678 418 ICV_53 $T=627440 334560 0 0 $X=627250 $Y=334320
X2776 1 2 1752 1719 405 ICV_53 $T=655040 323680 1 0 $X=654850 $Y=320720
X2777 1 2 1793 1797 407 ICV_53 $T=673440 345440 1 0 $X=673250 $Y=342480
X2778 1 2 ICV_54 $T=47840 323680 1 0 $X=47650 $Y=320720
X2779 1 2 ICV_54 $T=47840 350880 1 0 $X=47650 $Y=347920
X2780 1 2 ICV_54 $T=61640 329120 0 0 $X=61450 $Y=328880
X2781 1 2 ICV_54 $T=145820 318240 0 0 $X=145630 $Y=318000
X2782 1 2 ICV_54 $T=160080 372640 1 0 $X=159890 $Y=369680
X2783 1 2 ICV_54 $T=216200 318240 1 0 $X=216010 $Y=315280
X2784 1 2 ICV_54 $T=230000 361760 0 0 $X=229810 $Y=361520
X2785 1 2 ICV_54 $T=258060 356320 0 0 $X=257870 $Y=356080
X2786 1 2 ICV_54 $T=384560 356320 1 0 $X=384370 $Y=353360
X2787 1 2 ICV_54 $T=398360 340000 0 0 $X=398170 $Y=339760
X2788 1 2 ICV_54 $T=412620 318240 1 0 $X=412430 $Y=315280
X2789 1 2 ICV_54 $T=510600 323680 0 0 $X=510410 $Y=323440
X2790 1 2 ICV_54 $T=524860 340000 1 0 $X=524670 $Y=337040
X2791 1 2 ICV_54 $T=538660 318240 0 0 $X=538470 $Y=318000
X2792 1 2 ICV_54 $T=552920 323680 1 0 $X=552730 $Y=320720
X2793 1 2 ICV_54 $T=552920 329120 1 0 $X=552730 $Y=326160
X2794 1 2 ICV_54 $T=580980 340000 1 0 $X=580790 $Y=337040
X2795 1 2 ICV_54 $T=594780 367200 0 0 $X=594590 $Y=366960
X2796 1 2 ICV_54 $T=637100 323680 1 0 $X=636910 $Y=320720
X2797 1 2 ICV_54 $T=665160 329120 1 0 $X=664970 $Y=326160
X2798 1 2 ICV_54 $T=693220 372640 1 0 $X=693030 $Y=369680
X2799 1 2 ICV_54 $T=707020 312800 0 0 $X=706830 $Y=312560
X2800 1 2 ICV_54 $T=721280 378080 1 0 $X=721090 $Y=375120
X2801 1 2 22 2 31 1 sky130_fd_sc_hd__clkbuf_16 $T=10580 361760 0 0 $X=10390 $Y=361520
X2802 1 2 103 2 105 1 sky130_fd_sc_hd__clkbuf_16 $T=105340 361760 1 0 $X=105150 $Y=358800
X2803 1 2 111 2 108 1 sky130_fd_sc_hd__clkbuf_16 $T=111780 367200 1 0 $X=111590 $Y=364240
X2804 1 2 114 2 107 1 sky130_fd_sc_hd__clkbuf_16 $T=114540 361760 1 0 $X=114350 $Y=358800
X2805 1 2 248 2 253 1 sky130_fd_sc_hd__clkbuf_16 $T=301760 356320 0 0 $X=301570 $Y=356080
X2806 1 2 251 2 257 1 sky130_fd_sc_hd__clkbuf_16 $T=307740 356320 1 0 $X=307550 $Y=353360
X2807 1 2 255 2 264 1 sky130_fd_sc_hd__clkbuf_16 $T=314640 350880 0 0 $X=314450 $Y=350640
X2808 1 2 256 2 265 1 sky130_fd_sc_hd__clkbuf_16 $T=315100 345440 0 0 $X=314910 $Y=345200
X2809 1 2 258 2 262 1 sky130_fd_sc_hd__clkbuf_16 $T=316020 356320 0 0 $X=315830 $Y=356080
X2810 1 2 259 2 266 1 sky130_fd_sc_hd__clkbuf_16 $T=316940 356320 1 0 $X=316750 $Y=353360
X2811 1 2 165 2 276 1 sky130_fd_sc_hd__clkbuf_16 $T=326600 312800 0 0 $X=326410 $Y=312560
X2812 1 2 291 2 158 1 sky130_fd_sc_hd__clkbuf_16 $T=349600 372640 0 0 $X=349410 $Y=372400
X2813 1 2 301 2 152 1 sky130_fd_sc_hd__clkbuf_16 $T=358800 372640 0 0 $X=358610 $Y=372400
X2814 1 2 303 2 181 1 sky130_fd_sc_hd__clkbuf_16 $T=360640 378080 1 0 $X=360450 $Y=375120
X2815 1 2 304 2 175 1 sky130_fd_sc_hd__clkbuf_16 $T=362480 367200 1 0 $X=362290 $Y=364240
X2816 1 2 305 2 163 1 sky130_fd_sc_hd__clkbuf_16 $T=362940 372640 1 0 $X=362750 $Y=369680
X2817 1 2 341 2 156 1 sky130_fd_sc_hd__clkbuf_16 $T=418140 367200 1 0 $X=417950 $Y=364240
X2818 1 2 384 2 387 1 sky130_fd_sc_hd__clkbuf_16 $T=499560 361760 1 0 $X=499370 $Y=358800
X2819 1 2 111 2 394 1 sky130_fd_sc_hd__clkbuf_16 $T=510140 361760 1 0 $X=509950 $Y=358800
X2820 1 2 103 2 390 1 sky130_fd_sc_hd__clkbuf_16 $T=511060 361760 0 0 $X=510870 $Y=361520
X2821 1 2 114 2 396 1 sky130_fd_sc_hd__clkbuf_16 $T=520260 361760 0 0 $X=520070 $Y=361520
X2822 1 2 561 533 52 ICV_56 $T=26220 350880 0 0 $X=26030 $Y=350640
X2823 1 2 579 545 54 ICV_56 $T=34960 318240 0 0 $X=34770 $Y=318000
X2824 1 2 583 553 39 ICV_56 $T=40480 334560 1 0 $X=40290 $Y=331600
X2825 1 2 586 590 36 ICV_56 $T=40940 350880 1 0 $X=40750 $Y=347920
X2826 1 2 648 645 39 ICV_56 $T=70380 356320 0 0 $X=70190 $Y=356080
X2827 1 2 680 90 55 ICV_56 $T=87860 372640 1 0 $X=87670 $Y=369680
X2828 1 2 798 783 52 ICV_56 $T=152720 334560 1 0 $X=152530 $Y=331600
X2829 1 2 1049 239 176 ICV_56 $T=292100 372640 0 0 $X=291910 $Y=372400
X2830 1 2 1104 1076 197 ICV_56 $T=321540 345440 1 0 $X=321350 $Y=342480
X2831 1 2 1115 254 184 ICV_56 $T=327980 318240 0 0 $X=327790 $Y=318000
X2832 1 2 1181 1173 275 ICV_56 $T=363400 350880 0 0 $X=363210 $Y=350640
X2833 1 2 1191 1186 296 ICV_56 $T=377200 340000 1 0 $X=377010 $Y=337040
X2834 1 2 1252 1250 267 ICV_56 $T=401120 323680 0 0 $X=400930 $Y=323440
X2835 1 2 1237 1223 263 ICV_56 $T=405720 329120 1 0 $X=405530 $Y=326160
X2836 1 2 1260 333 268 ICV_56 $T=405720 372640 1 0 $X=405530 $Y=369680
X2837 1 2 1271 1261 280 ICV_56 $T=410320 350880 0 0 $X=410130 $Y=350640
X2838 1 2 1435 1457 275 ICV_56 $T=503700 340000 0 0 $X=503510 $Y=339760
X2839 1 2 1526 1507 422 ICV_56 $T=540960 318240 0 0 $X=540770 $Y=318000
X2840 1 2 1583 1585 418 ICV_56 $T=573620 356320 1 0 $X=573430 $Y=353360
X2841 1 2 1590 1585 424 ICV_56 $T=574080 340000 1 0 $X=573890 $Y=337040
X2842 1 2 1703 1682 409 ICV_56 $T=630200 323680 1 0 $X=630010 $Y=320720
X2843 1 2 1718 445 409 ICV_56 $T=638480 312800 0 0 $X=638290 $Y=312560
X2844 1 2 1806 1797 408 ICV_56 $T=681720 334560 0 0 $X=681530 $Y=334320
X2845 1 2 1864 1869 407 ICV_56 $T=714380 329120 1 0 $X=714190 $Y=326160
X2846 1 2 1888 469 422 ICV_56 $T=718060 318240 0 0 $X=717870 $Y=318000
X2847 1 2 1890 1889 405 ICV_56 $T=736000 334560 1 0 $X=735810 $Y=331600
X2848 1 2 1904 1891 417 ICV_56 $T=736000 345440 1 0 $X=735810 $Y=342480
X2849 1 2 1906 1891 408 ICV_56 $T=736000 350880 1 0 $X=735810 $Y=347920
X2850 1 2 575 15 597 597 590 39 ICV_58 $T=34040 356320 0 0 $X=33850 $Y=356080
X2851 1 2 732 25 742 742 747 28 ICV_58 $T=108560 323680 1 0 $X=108370 $Y=320720
X2852 1 2 744 14 773 773 759 36 ICV_58 $T=128340 345440 0 0 $X=128150 $Y=345200
X2853 1 2 826 187 842 842 820 197 ICV_58 $T=174340 334560 0 0 $X=174150 $Y=334320
X2854 1 2 907 175 923 923 924 188 ICV_58 $T=216660 361760 1 0 $X=216470 $Y=358800
X2855 1 2 939 187 959 959 961 197 ICV_58 $T=234600 334560 0 0 $X=234410 $Y=334320
X2856 1 2 963 152 994 994 975 176 ICV_58 $T=253920 372640 1 0 $X=253730 $Y=369680
X2857 1 2 165 194 279 1123 1131 275 ICV_58 $T=325220 356320 0 0 $X=325030 $Y=356080
X2858 1 2 1118 262 1166 1166 1138 269 ICV_58 $T=342700 323680 0 0 $X=342510 $Y=323440
X2859 1 2 312 264 1231 1231 319 296 ICV_58 $T=380880 372640 0 0 $X=380690 $Y=372400
X2860 1 2 1431 260 1455 1455 1456 267 ICV_58 $T=487140 350880 0 0 $X=486950 $Y=350640
X2861 1 2 1413 257 1476 1471 1457 277 ICV_58 $T=501400 345440 1 0 $X=501210 $Y=342480
X2862 1 2 1612 410 1642 1642 1616 417 ICV_58 $T=591560 345440 1 0 $X=591370 $Y=342480
X2863 1 2 1808 397 1838 1843 1818 408 ICV_58 $T=690000 361760 0 0 $X=689810 $Y=361520
X2864 1 2 1859 400 1885 1834 1827 418 ICV_58 $T=707480 334560 0 0 $X=707290 $Y=334320
X2865 1 2 466 410 1909 1909 469 417 ICV_58 $T=721740 318240 1 0 $X=721550 $Y=315280
X2866 1 2 1859 399 1911 1911 1889 408 ICV_58 $T=721740 340000 1 0 $X=721550 $Y=337040
X2867 1 2 587 590 37 ICV_62 $T=45540 350880 0 0 $X=45350 $Y=350640
X2868 1 2 629 624 54 ICV_62 $T=61640 361760 1 0 $X=61450 $Y=358800
X2869 1 2 795 741 36 ICV_62 $T=157780 350880 0 0 $X=157590 $Y=350640
X2870 1 2 897 868 176 ICV_62 $T=213900 372640 0 0 $X=213710 $Y=372400
X2871 1 2 965 958 201 ICV_62 $T=246560 334560 1 0 $X=246370 $Y=331600
X2872 1 2 966 958 197 ICV_62 $T=249320 334560 0 0 $X=249130 $Y=334320
X2873 1 2 969 211 185 ICV_62 $T=256220 378080 1 0 $X=256030 $Y=375120
X2874 1 2 986 987 184 ICV_62 $T=259900 340000 0 0 $X=259710 $Y=339760
X2875 1 2 1070 1021 174 ICV_62 $T=301760 361760 1 0 $X=301570 $Y=358800
X2876 1 2 1064 1021 194 ICV_62 $T=310500 367200 1 0 $X=310310 $Y=364240
X2877 1 2 1114 254 198 ICV_62 $T=325680 323680 0 0 $X=325490 $Y=323440
X2878 1 2 1214 1225 277 ICV_62 $T=385940 345440 1 0 $X=385750 $Y=342480
X2879 1 2 1279 1250 269 ICV_62 $T=414920 323680 1 0 $X=414730 $Y=320720
X2880 1 2 1336 1313 263 ICV_62 $T=445280 334560 0 0 $X=445090 $Y=334320
X2881 1 2 1347 1350 277 ICV_62 $T=449880 334560 0 0 $X=449690 $Y=334320
X2882 1 2 1392 1382 296 ICV_62 $T=470120 318240 0 0 $X=469930 $Y=318000
X2883 1 2 1409 1371 268 ICV_62 $T=477940 345440 0 0 $X=477750 $Y=345200
X2884 1 2 1420 1391 277 ICV_62 $T=484380 367200 0 0 $X=484190 $Y=366960
X2885 1 2 1462 1434 275 ICV_62 $T=506000 367200 0 0 $X=505810 $Y=366960
X2886 1 2 391 393 263 ICV_62 $T=512900 378080 1 0 $X=512710 $Y=375120
X2887 1 2 1524 1503 417 ICV_62 $T=544180 350880 1 0 $X=543990 $Y=347920
X2888 1 2 1624 1616 422 ICV_62 $T=589720 350880 1 0 $X=589530 $Y=347920
X2889 1 2 1598 1599 417 ICV_62 $T=590180 318240 0 0 $X=589990 $Y=318000
X2890 1 2 1798 1780 408 ICV_62 $T=675280 367200 1 0 $X=675090 $Y=364240
X2891 1 2 1840 1781 417 ICV_62 $T=705180 334560 1 0 $X=704990 $Y=331600
X2892 1 2 48 40 578 ICV_66 $T=26220 367200 0 0 $X=26030 $Y=366960
X2893 1 2 608 44 633 ICV_66 $T=54280 356320 0 0 $X=54090 $Y=356080
X2894 1 2 644 42 662 ICV_66 $T=68540 361760 1 0 $X=68350 $Y=358800
X2895 1 2 750 25 765 ICV_66 $T=124660 340000 1 0 $X=124470 $Y=337040
X2896 1 2 825 171 829 ICV_66 $T=166520 323680 0 0 $X=166330 $Y=323440
X2897 1 2 218 189 926 ICV_66 $T=222640 312800 0 0 $X=222450 $Y=312560
X2898 1 2 914 170 928 ICV_66 $T=222640 318240 0 0 $X=222450 $Y=318000
X2899 1 2 939 172 955 ICV_66 $T=236900 345440 1 0 $X=236710 $Y=342480
X2900 1 2 992 191 1013 ICV_66 $T=264960 334560 1 0 $X=264770 $Y=331600
X2901 1 2 1022 181 1015 ICV_66 $T=278760 367200 0 0 $X=278570 $Y=366960
X2902 1 2 1035 172 1060 ICV_66 $T=293020 334560 1 0 $X=292830 $Y=331600
X2903 1 2 1008 181 1064 ICV_66 $T=293020 367200 1 0 $X=292830 $Y=364240
X2904 1 2 250 190 1090 ICV_66 $T=306820 318240 0 0 $X=306630 $Y=318000
X2905 1 2 1079 156 1091 ICV_66 $T=306820 361760 0 0 $X=306630 $Y=361520
X2906 1 2 278 266 1144 ICV_66 $T=334880 318240 0 0 $X=334690 $Y=318000
X2907 1 2 1203 266 1212 ICV_66 $T=377200 329120 1 0 $X=377010 $Y=326160
X2908 1 2 1205 265 1214 ICV_66 $T=377200 345440 1 0 $X=377010 $Y=342480
X2909 1 2 1428 265 1469 ICV_66 $T=503240 329120 0 0 $X=503050 $Y=328880
X2910 1 2 1428 253 1470 ICV_66 $T=503240 334560 0 0 $X=503050 $Y=334320
X2911 1 2 1431 265 1473 ICV_66 $T=503240 356320 0 0 $X=503050 $Y=356080
X2912 1 2 1429 253 1474 ICV_66 $T=503240 372640 0 0 $X=503050 $Y=372400
X2913 1 2 427 399 1545 ICV_66 $T=545560 318240 1 0 $X=545370 $Y=315280
X2914 1 2 1640 415 440 ICV_66 $T=601680 318240 1 0 $X=601490 $Y=315280
X2915 1 2 1699 397 1716 ICV_66 $T=629740 367200 1 0 $X=629550 $Y=364240
X2916 1 2 1699 414 1743 ICV_66 $T=643540 356320 0 0 $X=643350 $Y=356080
X2917 1 2 1699 399 1744 ICV_66 $T=643540 361760 0 0 $X=643350 $Y=361520
X2918 1 2 105 107 108 731 2 109 1 sky130_fd_sc_hd__and4b_2 $T=107640 367200 1 0 $X=107450 $Y=364240
X2919 1 2 105 107 108 110 2 78 1 sky130_fd_sc_hd__and4b_2 $T=108560 378080 1 0 $X=108370 $Y=375120
X2920 1 2 107 105 108 110 2 74 1 sky130_fd_sc_hd__and4b_2 $T=118220 372640 1 0 $X=118030 $Y=369680
X2921 1 2 108 107 105 110 2 17 1 sky130_fd_sc_hd__and4b_2 $T=118220 372640 0 0 $X=118030 $Y=372400
X2922 1 2 108 107 105 731 2 117 1 sky130_fd_sc_hd__and4b_2 $T=119600 361760 0 0 $X=119410 $Y=361520
X2923 1 2 107 105 108 731 2 125 1 sky130_fd_sc_hd__and4b_2 $T=122360 372640 1 0 $X=122170 $Y=369680
X2924 1 2 107 105 108 755 2 102 1 sky130_fd_sc_hd__and4b_2 $T=123740 372640 0 0 $X=123550 $Y=372400
X2925 1 2 121 122 123 6 2 755 1 sky130_fd_sc_hd__and4b_2 $T=127880 372640 1 0 $X=127690 $Y=369680
X2926 1 2 108 107 105 757 2 130 1 sky130_fd_sc_hd__and4b_2 $T=130180 361760 0 0 $X=129990 $Y=361520
X2927 1 2 105 107 108 757 2 133 1 sky130_fd_sc_hd__and4b_2 $T=132480 367200 1 0 $X=132290 $Y=364240
X2928 1 2 108 107 105 755 2 81 1 sky130_fd_sc_hd__and4b_2 $T=132480 372640 0 0 $X=132290 $Y=372400
X2929 1 2 105 107 108 755 2 119 1 sky130_fd_sc_hd__and4b_2 $T=132480 378080 1 0 $X=132290 $Y=375120
X2930 1 2 107 105 108 757 2 143 1 sky130_fd_sc_hd__and4b_2 $T=140760 361760 1 0 $X=140570 $Y=358800
X2931 1 2 105 107 108 782 2 149 1 sky130_fd_sc_hd__and4b_2 $T=146280 372640 0 0 $X=146090 $Y=372400
X2932 1 2 107 105 108 148 2 142 1 sky130_fd_sc_hd__and4b_2 $T=146280 378080 1 0 $X=146090 $Y=375120
X2933 1 2 122 121 123 6 2 780 1 sky130_fd_sc_hd__and4b_2 $T=146740 367200 0 0 $X=146550 $Y=366960
X2934 1 2 108 107 105 782 2 88 1 sky130_fd_sc_hd__and4b_2 $T=147200 372640 1 0 $X=147010 $Y=369680
X2935 1 2 105 107 108 148 2 151 1 sky130_fd_sc_hd__and4b_2 $T=150420 378080 1 0 $X=150230 $Y=375120
X2936 1 2 107 105 108 782 2 154 1 sky130_fd_sc_hd__and4b_2 $T=150880 367200 0 0 $X=150690 $Y=366960
X2937 1 2 108 107 105 780 2 147 1 sky130_fd_sc_hd__and4b_2 $T=151340 367200 1 0 $X=151150 $Y=364240
X2938 1 2 105 107 108 780 2 91 1 sky130_fd_sc_hd__and4b_2 $T=154100 361760 1 0 $X=153910 $Y=358800
X2939 1 2 107 105 108 780 2 106 1 sky130_fd_sc_hd__and4b_2 $T=155480 367200 1 0 $X=155290 $Y=364240
X2940 1 2 394 396 390 1488 2 373 1 sky130_fd_sc_hd__and4b_2 $T=515660 367200 1 0 $X=515470 $Y=364240
X2941 1 2 396 390 394 1488 2 331 1 sky130_fd_sc_hd__and4b_2 $T=520720 361760 1 0 $X=520530 $Y=358800
X2942 1 2 390 396 394 1488 2 411 1 sky130_fd_sc_hd__and4b_2 $T=527160 367200 0 0 $X=526970 $Y=366960
X2943 1 2 396 390 394 1508 2 425 1 sky130_fd_sc_hd__and4b_2 $T=540040 372640 1 0 $X=539850 $Y=369680
X2944 1 2 394 396 390 1508 2 338 1 sky130_fd_sc_hd__and4b_2 $T=540040 372640 0 0 $X=539850 $Y=372400
X2945 1 2 394 396 390 1512 2 385 1 sky130_fd_sc_hd__and4b_2 $T=543260 367200 1 0 $X=543070 $Y=364240
X2946 1 2 390 396 394 1508 2 354 1 sky130_fd_sc_hd__and4b_2 $T=543260 378080 1 0 $X=543070 $Y=375120
X2947 1 2 390 396 394 1512 2 380 1 sky130_fd_sc_hd__and4b_2 $T=543720 361760 0 0 $X=543530 $Y=361520
X2948 1 2 396 390 394 1512 2 386 1 sky130_fd_sc_hd__and4b_2 $T=543720 367200 0 0 $X=543530 $Y=366960
X2949 1 2 105 107 108 731 2 129 1 sky130_fd_sc_hd__and4_2 $T=128340 367200 1 0 $X=128150 $Y=364240
X2950 1 2 105 107 108 757 2 131 1 sky130_fd_sc_hd__and4_2 $T=132480 361760 1 0 $X=132290 $Y=358800
X2951 1 2 105 107 108 755 2 132 1 sky130_fd_sc_hd__and4_2 $T=132480 372640 1 0 $X=132290 $Y=369680
X2952 1 2 105 107 108 782 2 157 1 sky130_fd_sc_hd__and4_2 $T=155020 367200 0 0 $X=154830 $Y=366960
X2953 1 2 105 107 108 780 2 162 1 sky130_fd_sc_hd__and4_2 $T=159620 361760 0 0 $X=159430 $Y=361520
X2954 1 2 390 396 394 1488 2 297 1 sky130_fd_sc_hd__and4_2 $T=525320 372640 1 0 $X=525130 $Y=369680
X2955 1 2 121 122 123 7 2 1512 1 sky130_fd_sc_hd__and4_2 $T=531760 367200 0 0 $X=531570 $Y=366960
X2956 1 2 390 396 394 1508 2 336 1 sky130_fd_sc_hd__and4_2 $T=544180 372640 1 0 $X=543990 $Y=369680
X2957 1 2 390 396 394 1512 2 352 1 sky130_fd_sc_hd__and4_2 $T=547400 367200 1 0 $X=547210 $Y=364240
X2958 1 2 804 805 2 28 1 sky130_fd_sc_hd__ebufn_4 $T=154100 345440 1 0 $X=153910 $Y=342480
X2959 1 2 804 805 2 37 1 sky130_fd_sc_hd__ebufn_4 $T=162380 350880 0 0 $X=162190 $Y=350640
X2960 1 2 804 805 2 52 1 sky130_fd_sc_hd__ebufn_4 $T=162380 356320 1 0 $X=162190 $Y=353360
X2961 1 2 804 805 2 63 1 sky130_fd_sc_hd__ebufn_4 $T=163300 361760 1 0 $X=163110 $Y=358800
X2962 1 2 804 805 2 38 1 sky130_fd_sc_hd__ebufn_4 $T=163300 361760 0 0 $X=163110 $Y=361520
X2963 1 2 804 805 2 36 1 sky130_fd_sc_hd__ebufn_4 $T=163760 345440 0 0 $X=163570 $Y=345200
X2964 1 2 804 805 2 176 1 sky130_fd_sc_hd__ebufn_4 $T=164680 356320 0 0 $X=164490 $Y=356080
X2965 1 2 804 805 2 34 1 sky130_fd_sc_hd__ebufn_4 $T=166060 350880 1 0 $X=165870 $Y=347920
X2966 1 2 804 805 2 57 1 sky130_fd_sc_hd__ebufn_4 $T=168360 356320 1 0 $X=168170 $Y=353360
X2967 1 2 804 805 2 180 1 sky130_fd_sc_hd__ebufn_4 $T=169280 361760 1 0 $X=169090 $Y=358800
X2968 1 2 804 805 2 184 1 sky130_fd_sc_hd__ebufn_4 $T=172040 345440 1 0 $X=171850 $Y=342480
X2969 1 2 804 805 2 185 1 sky130_fd_sc_hd__ebufn_4 $T=172040 350880 1 0 $X=171850 $Y=347920
X2970 1 2 804 805 2 193 1 sky130_fd_sc_hd__ebufn_4 $T=174800 350880 0 0 $X=174610 $Y=350640
X2971 1 2 804 805 2 59 1 sky130_fd_sc_hd__ebufn_4 $T=175260 361760 1 0 $X=175070 $Y=358800
X2972 1 2 804 805 2 54 1 sky130_fd_sc_hd__ebufn_4 $T=175720 356320 1 0 $X=175530 $Y=353360
X2973 1 2 804 805 2 186 1 sky130_fd_sc_hd__ebufn_4 $T=176180 345440 0 0 $X=175990 $Y=345200
X2974 1 2 804 805 2 33 1 sky130_fd_sc_hd__ebufn_4 $T=176180 367200 1 0 $X=175990 $Y=364240
X2975 1 2 804 805 2 174 1 sky130_fd_sc_hd__ebufn_4 $T=177100 356320 0 0 $X=176910 $Y=356080
X2976 1 2 804 805 2 47 1 sky130_fd_sc_hd__ebufn_4 $T=177560 361760 0 0 $X=177370 $Y=361520
X2977 1 2 804 805 2 179 1 sky130_fd_sc_hd__ebufn_4 $T=178020 345440 1 0 $X=177830 $Y=342480
X2978 1 2 804 805 2 39 1 sky130_fd_sc_hd__ebufn_4 $T=181700 356320 1 0 $X=181510 $Y=353360
X2979 1 2 804 805 2 166 1 sky130_fd_sc_hd__ebufn_4 $T=182160 345440 0 0 $X=181970 $Y=345200
X2980 1 2 804 805 2 199 1 sky130_fd_sc_hd__ebufn_4 $T=182160 350880 1 0 $X=181970 $Y=347920
X2981 1 2 804 805 2 188 1 sky130_fd_sc_hd__ebufn_4 $T=182160 361760 1 0 $X=181970 $Y=358800
X2982 1 2 804 805 2 167 1 sky130_fd_sc_hd__ebufn_4 $T=182160 367200 1 0 $X=181970 $Y=364240
X2983 1 2 804 805 2 201 1 sky130_fd_sc_hd__ebufn_4 $T=184000 350880 0 0 $X=183810 $Y=350640
X2984 1 2 804 805 2 55 1 sky130_fd_sc_hd__ebufn_4 $T=185380 361760 0 0 $X=185190 $Y=361520
X2985 1 2 804 805 2 197 1 sky130_fd_sc_hd__ebufn_4 $T=188600 345440 1 0 $X=188410 $Y=342480
X2986 1 2 804 805 2 194 1 sky130_fd_sc_hd__ebufn_4 $T=188600 361760 1 0 $X=188410 $Y=358800
X2987 1 2 804 805 2 75 1 sky130_fd_sc_hd__ebufn_4 $T=188600 367200 1 0 $X=188410 $Y=364240
X2988 1 2 804 805 2 198 1 sky130_fd_sc_hd__ebufn_4 $T=194580 345440 1 0 $X=194390 $Y=342480
X2989 1 2 804 805 2 49 1 sky130_fd_sc_hd__ebufn_4 $T=199640 356320 1 0 $X=199450 $Y=353360
X2990 1 2 105 107 108 731 2 116 1 sky130_fd_sc_hd__nor4b_2 $T=112240 367200 0 0 $X=112050 $Y=366960
X2991 1 2 105 107 108 110 2 56 1 sky130_fd_sc_hd__nor4b_2 $T=112700 378080 1 0 $X=112510 $Y=375120
X2992 1 2 121 122 123 6 2 110 1 sky130_fd_sc_hd__nor4b_2 $T=119600 378080 1 0 $X=119410 $Y=375120
X2993 1 2 105 107 108 757 2 16 1 sky130_fd_sc_hd__nor4b_2 $T=123740 361760 1 0 $X=123550 $Y=358800
X2994 1 2 105 107 108 755 2 89 1 sky130_fd_sc_hd__nor4b_2 $T=126040 367200 0 0 $X=125850 $Y=366960
X2995 1 2 105 107 108 780 2 68 1 sky130_fd_sc_hd__nor4b_2 $T=136620 367200 1 0 $X=136430 $Y=364240
X2996 1 2 105 107 108 782 2 23 1 sky130_fd_sc_hd__nor4b_2 $T=138000 372640 0 0 $X=137810 $Y=372400
X2997 1 2 390 396 394 1488 2 283 1 sky130_fd_sc_hd__nor4b_2 $T=517040 367200 0 0 $X=516850 $Y=366960
X2998 1 2 390 396 394 395 2 403 1 sky130_fd_sc_hd__nor4b_2 $T=517500 372640 0 0 $X=517310 $Y=372400
X2999 1 2 390 396 394 1512 2 286 1 sky130_fd_sc_hd__nor4b_2 $T=529920 367200 1 0 $X=529730 $Y=364240
X3000 1 2 390 396 394 1508 2 314 1 sky130_fd_sc_hd__nor4b_2 $T=530380 372640 1 0 $X=530190 $Y=369680
X3001 1 2 105 108 731 107 2 79 1 sky130_fd_sc_hd__and4bb_2 $T=109020 372640 1 0 $X=108830 $Y=369680
X3002 1 2 108 107 731 105 2 112 1 sky130_fd_sc_hd__and4bb_2 $T=113160 361760 0 0 $X=112970 $Y=361520
X3003 1 2 105 108 110 107 2 113 1 sky130_fd_sc_hd__and4bb_2 $T=113160 372640 0 0 $X=112970 $Y=372400
X3004 1 2 108 105 731 107 2 60 1 sky130_fd_sc_hd__and4bb_2 $T=113620 372640 1 0 $X=113430 $Y=369680
X3005 1 2 121 123 6 122 2 731 1 sky130_fd_sc_hd__and4bb_2 $T=121440 367200 0 0 $X=121250 $Y=366960
X3006 1 2 105 108 757 107 2 29 1 sky130_fd_sc_hd__and4bb_2 $T=123740 367200 1 0 $X=123550 $Y=364240
X3007 1 2 108 105 757 107 2 124 1 sky130_fd_sc_hd__and4bb_2 $T=124200 361760 0 0 $X=124010 $Y=361520
X3008 1 2 105 108 755 107 2 127 1 sky130_fd_sc_hd__and4bb_2 $T=126960 378080 1 0 $X=126770 $Y=375120
X3009 1 2 108 105 755 107 2 128 1 sky130_fd_sc_hd__and4bb_2 $T=127880 372640 0 0 $X=127690 $Y=372400
X3010 1 2 108 107 755 105 2 85 1 sky130_fd_sc_hd__and4bb_2 $T=131560 367200 0 0 $X=131370 $Y=366960
X3011 1 2 108 107 757 105 2 92 1 sky130_fd_sc_hd__and4bb_2 $T=134320 361760 0 0 $X=134130 $Y=361520
X3012 1 2 123 122 6 121 2 757 1 sky130_fd_sc_hd__and4bb_2 $T=136160 361760 1 0 $X=135970 $Y=358800
X3013 1 2 108 107 780 105 2 135 1 sky130_fd_sc_hd__and4bb_2 $T=138920 361760 0 0 $X=138730 $Y=361520
X3014 1 2 105 108 782 107 2 136 1 sky130_fd_sc_hd__and4bb_2 $T=138920 367200 0 0 $X=138730 $Y=366960
X3015 1 2 108 107 782 105 2 137 1 sky130_fd_sc_hd__and4bb_2 $T=139380 372640 1 0 $X=139190 $Y=369680
X3016 1 2 108 105 782 107 2 138 1 sky130_fd_sc_hd__and4bb_2 $T=139380 378080 1 0 $X=139190 $Y=375120
X3017 1 2 108 105 780 107 2 140 1 sky130_fd_sc_hd__and4bb_2 $T=142140 367200 1 0 $X=141950 $Y=364240
X3018 1 2 105 108 780 107 2 146 1 sky130_fd_sc_hd__and4bb_2 $T=146740 367200 1 0 $X=146550 $Y=364240
X3019 1 2 123 121 6 122 2 782 1 sky130_fd_sc_hd__and4bb_2 $T=150420 372640 0 0 $X=150230 $Y=372400
X3020 1 2 390 394 395 396 2 392 1 sky130_fd_sc_hd__and4bb_2 $T=512900 372640 0 0 $X=512710 $Y=372400
X3021 1 2 394 390 395 396 2 285 1 sky130_fd_sc_hd__and4bb_2 $T=517500 378080 1 0 $X=517310 $Y=375120
X3022 1 2 390 394 1488 396 2 330 1 sky130_fd_sc_hd__and4bb_2 $T=519800 367200 1 0 $X=519610 $Y=364240
X3023 1 2 394 396 1488 390 2 402 1 sky130_fd_sc_hd__and4bb_2 $T=519800 372640 1 0 $X=519610 $Y=369680
X3024 1 2 394 390 1488 396 2 310 1 sky130_fd_sc_hd__and4bb_2 $T=522560 367200 0 0 $X=522370 $Y=366960
X3025 1 2 123 122 7 121 2 1488 1 sky130_fd_sc_hd__and4bb_2 $T=525320 367200 1 0 $X=525130 $Y=364240
X3026 1 2 394 396 1508 390 2 404 1 sky130_fd_sc_hd__and4bb_2 $T=526240 372640 0 0 $X=526050 $Y=372400
X3027 1 2 394 390 1508 396 2 292 1 sky130_fd_sc_hd__and4bb_2 $T=529000 378080 1 0 $X=528810 $Y=375120
X3028 1 2 123 121 7 122 2 1508 1 sky130_fd_sc_hd__and4bb_2 $T=530840 372640 0 0 $X=530650 $Y=372400
X3029 1 2 390 394 1508 396 2 416 1 sky130_fd_sc_hd__and4bb_2 $T=533600 378080 1 0 $X=533410 $Y=375120
X3030 1 2 394 390 1512 396 2 388 1 sky130_fd_sc_hd__and4bb_2 $T=538660 367200 1 0 $X=538470 $Y=364240
X3031 1 2 390 394 421 396 2 316 1 sky130_fd_sc_hd__and4bb_2 $T=538660 378080 1 0 $X=538470 $Y=375120
X3032 1 2 390 394 1512 396 2 419 1 sky130_fd_sc_hd__and4bb_2 $T=539120 361760 0 0 $X=538930 $Y=361520
X3033 1 2 394 396 1512 390 2 353 1 sky130_fd_sc_hd__and4bb_2 $T=539120 367200 0 0 $X=538930 $Y=366960
X3034 1 2 12 2 3 1 sky130_fd_sc_hd__clkbuf_4 $T=7820 361760 0 0 $X=7630 $Y=361520
X3035 1 2 6 2 805 1 sky130_fd_sc_hd__clkbuf_4 $T=160540 361760 1 0 $X=160350 $Y=358800
X3036 2 1 804 sky130_fd_sc_hd__conb_1 $T=172500 350880 0 0 $X=172310 $Y=350640
X3037 1 2 9 46 564 564 27 59 ICV_68 $T=20240 378080 1 0 $X=20050 $Y=375120
X3038 1 2 694 15 706 704 705 52 ICV_68 $T=90160 356320 1 0 $X=89970 $Y=353360
X3039 1 2 913 191 932 930 922 186 ICV_68 $T=223560 345440 1 0 $X=223370 $Y=342480
X3040 1 2 992 189 1024 1024 1010 199 ICV_68 $T=272320 323680 0 0 $X=272130 $Y=323440
X3041 1 2 1073 170 1108 1100 1083 199 ICV_68 $T=317400 329120 0 0 $X=317210 $Y=328880
X3042 1 2 1301 266 1315 1315 1313 275 ICV_68 $T=426880 345440 1 0 $X=426690 $Y=342480
X3043 1 2 1284 266 1320 1320 1295 275 ICV_68 $T=429640 323680 0 0 $X=429450 $Y=323440
X3044 1 2 1301 260 1343 1343 1313 267 ICV_68 $T=441140 340000 1 0 $X=440950 $Y=337040
X3045 1 2 1334 264 1374 1375 1342 275 ICV_68 $T=454940 367200 1 0 $X=454750 $Y=364240
X3046 1 2 1485 410 1518 1520 1506 418 ICV_68 $T=530380 340000 1 0 $X=530190 $Y=337040
X3047 1 2 1575 412 1590 1589 1585 422 ICV_68 $T=567180 345440 1 0 $X=566990 $Y=342480
X3048 1 2 1540 414 1594 1594 426 422 ICV_68 $T=567180 367200 0 0 $X=566990 $Y=366960
X3049 1 2 1655 414 1689 1689 1668 422 ICV_68 $T=616400 367200 1 0 $X=616210 $Y=364240
X3050 1 2 447 414 1728 1728 450 422 ICV_68 $T=637100 367200 0 0 $X=636910 $Y=366960
X3051 1 2 1712 415 1730 1730 1719 418 ICV_68 $T=637560 334560 1 0 $X=637370 $Y=331600
X3052 1 2 1713 398 1758 1761 1722 422 ICV_68 $T=651360 350880 1 0 $X=651170 $Y=347920
X3053 1 2 1860 414 1877 1877 1871 422 ICV_68 $T=709780 350880 0 0 $X=709590 $Y=350640
X3054 1 2 1859 415 1917 1917 1889 418 ICV_68 $T=729560 329120 1 0 $X=729370 $Y=326160
X3055 1 2 526 18 547 ICV_69 $T=8740 350880 0 0 $X=8550 $Y=350640
X3056 1 2 525 25 551 ICV_69 $T=11960 345440 0 0 $X=11770 $Y=345200
X3057 1 2 41 14 50 ICV_69 $T=20240 312800 0 0 $X=20050 $Y=312560
X3058 1 2 575 13 581 ICV_69 $T=31740 350880 1 0 $X=31550 $Y=347920
X3059 1 2 94 18 695 ICV_69 $T=86940 318240 1 0 $X=86750 $Y=315280
X3060 1 2 672 25 709 ICV_69 $T=92920 345440 0 0 $X=92730 $Y=345200
X3061 1 2 750 13 774 ICV_69 $T=135240 334560 1 0 $X=135050 $Y=331600
X3062 1 2 826 190 848 ICV_69 $T=178940 340000 1 0 $X=178750 $Y=337040
X3063 1 2 853 168 870 ICV_69 $T=192280 318240 0 0 $X=192090 $Y=318000
X3064 1 2 853 171 871 ICV_69 $T=192280 329120 0 0 $X=192090 $Y=328880
X3065 1 2 855 191 851 ICV_69 $T=192740 350880 0 0 $X=192550 $Y=350640
X3066 1 2 855 171 876 ICV_69 $T=192740 356320 0 0 $X=192550 $Y=356080
X3067 1 2 992 171 1006 ICV_69 $T=262660 329120 1 0 $X=262470 $Y=326160
X3068 1 2 1035 191 1041 ICV_69 $T=282440 329120 1 0 $X=282250 $Y=326160
X3069 1 2 1022 156 1044 ICV_69 $T=283820 367200 1 0 $X=283630 $Y=364240
X3070 1 2 1035 168 1050 ICV_69 $T=286580 323680 0 0 $X=286390 $Y=323440
X3071 1 2 244 171 1053 ICV_69 $T=287500 318240 0 0 $X=287310 $Y=318000
X3072 1 2 1061 168 1077 ICV_69 $T=300840 340000 1 0 $X=300650 $Y=337040
X3073 1 2 1146 265 1160 ICV_69 $T=343620 367200 0 0 $X=343430 $Y=366960
X3074 1 2 165 185 308 ICV_69 $T=360640 356320 0 0 $X=360450 $Y=356080
X3075 1 2 1146 273 1175 ICV_69 $T=360640 367200 0 0 $X=360450 $Y=366960
X3076 1 2 1171 257 1189 ICV_69 $T=361100 329120 0 0 $X=360910 $Y=328880
X3077 1 2 1249 265 1265 ICV_69 $T=399280 340000 1 0 $X=399090 $Y=337040
X3078 1 2 1257 265 1296 ICV_69 $T=417220 350880 0 0 $X=417030 $Y=350640
X3079 1 2 1334 265 1354 ICV_69 $T=443900 372640 1 0 $X=443710 $Y=369680
X3080 1 2 1428 273 1437 ICV_69 $T=487600 334560 1 0 $X=487410 $Y=331600
X3081 1 2 1496 410 1516 ICV_69 $T=529000 350880 0 0 $X=528810 $Y=350640
X3082 1 2 1496 397 1517 ICV_69 $T=529460 361760 0 0 $X=529270 $Y=361520
X3083 1 2 1527 414 1547 ICV_69 $T=543720 340000 1 0 $X=543530 $Y=337040
X3084 1 2 427 412 1552 ICV_69 $T=547860 318240 0 0 $X=547670 $Y=318000
X3085 1 2 1574 412 1597 ICV_69 $T=577300 323680 0 0 $X=577110 $Y=323440
X3086 1 2 1640 412 1672 ICV_69 $T=612260 323680 1 0 $X=612070 $Y=320720
X3087 1 2 446 398 1710 ICV_69 $T=627440 318240 1 0 $X=627250 $Y=315280
X3088 1 2 1747 399 1769 ICV_69 $T=655960 318240 1 0 $X=655770 $Y=315280
X3089 1 2 1779 410 1794 ICV_69 $T=667920 350880 1 0 $X=667730 $Y=347920
X3090 1 2 1862 410 1914 ICV_69 $T=725880 361760 0 0 $X=725690 $Y=361520
X3091 1 2 525 42 569 565 548 37 ICV_70 $T=21620 334560 0 0 $X=21430 $Y=334320
X3092 1 2 637 25 650 650 653 28 ICV_70 $T=63940 323680 1 0 $X=63750 $Y=320720
X3093 1 2 672 42 710 710 690 54 ICV_70 $T=92000 345440 1 0 $X=91810 $Y=342480
X3094 1 2 694 13 736 736 705 34 ICV_70 $T=105800 350880 0 0 $X=105610 $Y=350640
X3095 1 2 118 25 756 756 126 28 ICV_70 $T=120060 318240 1 0 $X=119870 $Y=315280
X3096 1 2 732 14 751 752 747 52 ICV_70 $T=120060 329120 1 0 $X=119870 $Y=326160
X3097 1 2 214 158 949 935 211 174 ICV_70 $T=232300 378080 1 0 $X=232110 $Y=375120
X3098 1 2 963 161 971 971 975 174 ICV_70 $T=246100 361760 0 0 $X=245910 $Y=361520
X3099 1 2 963 163 972 974 975 167 ICV_70 $T=246100 372640 0 0 $X=245910 $Y=372400
X3100 1 2 1030 170 1048 1059 1039 197 ICV_70 $T=288420 340000 1 0 $X=288230 $Y=337040
X3101 1 2 242 161 1057 1057 243 174 ICV_70 $T=288420 378080 1 0 $X=288230 $Y=375120
X3102 1 2 1118 260 1132 1132 1138 267 ICV_70 $T=330280 323680 0 0 $X=330090 $Y=323440
X3103 1 2 309 257 1234 1234 315 268 ICV_70 $T=386400 318240 0 0 $X=386210 $Y=318000
X3104 1 2 1378 262 1381 1390 1382 280 ICV_70 $T=470580 329120 0 0 $X=470390 $Y=328880
X3105 1 2 1575 410 1603 1608 1585 407 ICV_70 $T=582820 340000 0 0 $X=582630 $Y=339760
X3106 1 2 1712 414 1734 1734 1719 422 ICV_70 $T=638940 329120 0 0 $X=638750 $Y=328880
X3107 1 2 1747 410 1789 1776 1749 409 ICV_70 $T=667000 323680 0 0 $X=666810 $Y=323440
X3108 1 2 1860 412 1901 1875 1891 409 ICV_70 $T=723120 350880 0 0 $X=722930 $Y=350640
X3109 1 2 525 43 567 568 548 57 ICV_71 $T=21160 345440 0 0 $X=20970 $Y=345200
X3110 1 2 580 42 617 617 596 54 ICV_71 $T=49220 340000 0 0 $X=49030 $Y=339760
X3111 1 2 83 40 680 674 90 47 ICV_71 $T=77280 367200 0 0 $X=77090 $Y=366960
X3112 1 2 750 14 779 779 701 36 ICV_71 $T=133400 340000 0 0 $X=133210 $Y=339760
X3113 1 2 882 170 889 889 887 166 ICV_71 $T=203780 323680 1 0 $X=203590 $Y=320720
X3114 1 2 968 170 1000 1000 987 166 ICV_71 $T=259900 340000 1 0 $X=259710 $Y=337040
X3115 1 2 1095 265 1122 1122 261 277 ICV_71 $T=323380 361760 0 0 $X=323190 $Y=361520
X3116 1 2 278 264 299 300 289 267 ICV_71 $T=350060 312800 0 0 $X=349870 $Y=312560
X3117 1 2 1169 260 1180 1180 1173 267 ICV_71 $T=356500 345440 0 0 $X=356310 $Y=345200
X3118 1 2 1249 257 1290 1290 1256 268 ICV_71 $T=414000 334560 0 0 $X=413810 $Y=334320
X3119 1 2 1294 253 1312 1310 1308 269 ICV_71 $T=426880 356320 0 0 $X=426690 $Y=356080
X3120 1 2 1378 264 1392 1388 1382 275 ICV_71 $T=470120 323680 0 0 $X=469930 $Y=323440
X3121 1 2 1496 412 1534 1534 1509 424 ICV_71 $T=540500 356320 1 0 $X=540310 $Y=353360
X3122 1 2 1575 397 1591 1591 1585 409 ICV_71 $T=567180 345440 0 0 $X=566990 $Y=345200
X3123 1 2 1801 414 1819 1819 456 422 ICV_71 $T=680800 318240 1 0 $X=680610 $Y=315280
X3124 1 2 1862 414 1892 1892 1881 422 ICV_71 $T=713460 361760 0 0 $X=713270 $Y=361520
X3125 1 2 694 43 704 ICV_72 $T=89700 361760 1 0 $X=89510 $Y=358800
X3126 1 2 145 18 150 ICV_72 $T=146280 312800 0 0 $X=146090 $Y=312560
X3127 1 2 195 175 857 ICV_72 $T=184920 372640 0 0 $X=184730 $Y=372400
X3128 1 2 855 172 873 ICV_72 $T=192280 350880 1 0 $X=192090 $Y=347920
X3129 1 2 914 191 908 ICV_72 $T=224020 323680 1 0 $X=223830 $Y=320720
X3130 1 2 1022 163 247 ICV_72 $T=280600 378080 1 0 $X=280410 $Y=375120
X3131 1 2 244 191 1072 ICV_72 $T=296700 318240 0 0 $X=296510 $Y=318000
X3132 1 2 250 170 1113 ICV_72 $T=318780 312800 0 0 $X=318590 $Y=312560
X3133 1 2 342 260 1297 ICV_72 $T=418600 312800 0 0 $X=418410 $Y=312560
X3134 1 2 343 262 1299 ICV_72 $T=418600 372640 0 0 $X=418410 $Y=372400
X3135 1 2 1384 260 1418 ICV_72 $T=477480 361760 1 0 $X=477290 $Y=358800
X3136 1 2 401 399 1505 ICV_72 $T=520260 312800 0 0 $X=520070 $Y=312560
X3137 1 2 1485 412 1519 ICV_72 $T=530840 329120 0 0 $X=530650 $Y=328880
X3138 1 2 1574 400 1610 ICV_72 $T=581440 334560 1 0 $X=581250 $Y=331600
X3139 1 2 1713 415 1774 ICV_72 $T=658720 350880 0 0 $X=658530 $Y=350640
X3140 1 2 1808 399 1843 ICV_72 $T=693680 361760 1 0 $X=693490 $Y=358800
X3141 1 2 689 690 57 698 701 39 ICV_73 $T=89700 340000 0 0 $X=89510 $Y=339760
X3142 1 2 722 699 54 727 699 39 ICV_73 $T=103960 329120 1 0 $X=103770 $Y=326160
X3143 1 2 834 830 186 835 820 184 ICV_73 $T=173880 329120 0 0 $X=173690 $Y=328880
X3144 1 2 874 852 201 879 868 194 ICV_73 $T=201940 356320 0 0 $X=201750 $Y=356080
X3145 1 2 977 228 201 231 228 166 ICV_73 $T=258060 312800 0 0 $X=257870 $Y=312560
X3146 1 2 984 987 199 988 987 186 ICV_73 $T=258060 345440 0 0 $X=257870 $Y=345200
X3147 1 2 1085 1047 197 1072 245 198 ICV_73 $T=314180 323680 0 0 $X=313990 $Y=323440
X3148 1 2 1088 1083 197 1098 1076 186 ICV_73 $T=314180 340000 0 0 $X=313990 $Y=339760
X3149 1 2 1111 1083 184 1107 1083 179 ICV_73 $T=328440 329120 1 0 $X=328250 $Y=326160
X3150 1 2 1323 1308 280 1340 1342 263 ICV_73 $T=440680 361760 1 0 $X=440490 $Y=358800
X3151 1 2 367 358 296 369 370 268 ICV_73 $T=468740 378080 1 0 $X=468550 $Y=375120
X3152 1 2 1452 1456 280 1427 1457 296 ICV_73 $T=496800 356320 1 0 $X=496610 $Y=353360
X3153 1 2 1482 1425 263 1500 1507 408 ICV_73 $T=524860 323680 1 0 $X=524670 $Y=320720
X3154 1 2 1544 1543 407 1555 1543 424 ICV_73 $T=552920 345440 1 0 $X=552730 $Y=342480
X3155 1 2 1605 1585 408 1614 1616 407 ICV_73 $T=580980 350880 1 0 $X=580790 $Y=347920
X3156 1 2 1829 1818 417 1828 1827 407 ICV_73 $T=693220 350880 1 0 $X=693030 $Y=347920
X3157 1 2 23 19 534 534 41 200 ICV_74 $T=10580 312800 0 0 $X=10390 $Y=312560
X3158 1 2 92 31 686 686 98 200 ICV_74 $T=84640 367200 1 0 $X=84450 $Y=364240
X3159 1 2 58 164 878 878 884 200 ICV_74 $T=200100 350880 1 0 $X=199910 $Y=347920
X3160 1 2 92 144 910 910 907 200 ICV_74 $T=217120 367200 1 0 $X=216930 $Y=364240
X3161 1 2 78 164 937 937 950 200 ICV_74 $T=233680 334560 1 0 $X=233490 $Y=331600
X3162 1 2 102 164 964 964 968 200 ICV_74 $T=244720 356320 1 0 $X=244530 $Y=353360
X3163 1 2 117 164 993 993 233 200 ICV_74 $T=262200 323680 1 0 $X=262010 $Y=320720
X3164 1 2 162 144 997 997 1008 200 ICV_74 $T=263580 367200 0 0 $X=263390 $Y=366960
X3165 1 2 132 144 1074 1074 1079 200 ICV_74 $T=301760 367200 1 0 $X=301570 $Y=364240
X3166 1 2 271 272 1124 1124 1095 276 ICV_74 $T=330280 378080 1 0 $X=330090 $Y=375120
X3167 1 2 295 272 1168 1168 1171 276 ICV_74 $T=352360 329120 0 0 $X=352170 $Y=328880
X3168 1 2 321 272 1224 1224 1230 276 ICV_74 $T=384560 367200 0 0 $X=384370 $Y=366960
X3169 1 2 345 272 1298 1298 1284 276 ICV_74 $T=423660 334560 1 0 $X=423470 $Y=331600
X3170 1 2 380 272 1460 1460 1430 276 ICV_74 $T=497720 329120 1 0 $X=497530 $Y=326160
X3171 1 2 331 387 1741 1741 1747 276 ICV_74 $T=646300 318240 1 0 $X=646110 $Y=315280
X3172 1 2 385 387 1810 1810 1814 276 ICV_74 $T=682640 340000 1 0 $X=682450 $Y=337040
.ENDS
***************************************
.SUBCKT ICV_76 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=26
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 3 4 5 ICV_37 $T=1380 0 0 0 $X=1190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_77 1 2 3 4 5 6 7 8 9 10 11 12 13
** N=13 EP=13 IP=16 FDC=72
*.SEEDPROM
X0 1 2 6 7 8 3 4 5 ICV_13 $T=0 0 1 0 $X=-190 $Y=-2960
X1 1 2 11 12 13 3 9 10 ICV_13 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__mux4_1 VNB VPB A1 A0 S0 A3 A2 S1 VPWR X VGND
** N=161 EP=11 IP=0 FDC=26
*.SEEDPROM
M0 VGND A1 21 VNB nshort L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75001.3 a=0.063 p=1.14 mult=1 $X=395 $Y=235 $D=9
M1 22 A0 VGND VNB nshort L=0.15 W=0.42 AD=0.0567 AS=0.0567 PD=0.69 PS=0.69 NRD=22.848 NRS=0 m=1 r=2.8 sa=75000.6 sb=75000.9 a=0.063 p=1.14 mult=1 $X=815 $Y=235 $D=9
M2 17 12 22 VNB nshort L=0.15 W=0.42 AD=0.085225 AS=0.0567 PD=0.925 PS=0.69 NRD=18.564 NRS=22.848 m=1 r=2.8 sa=75001 sb=75000.5 a=0.063 p=1.14 mult=1 $X=1235 $Y=235 $D=9
M3 21 S0 17 VNB nshort L=0.15 W=0.42 AD=0.1092 AS=0.085225 PD=1.36 PS=0.925 NRD=0 NRS=0 m=1 r=2.8 sa=75001 sb=75000.2 a=0.063 p=1.14 mult=1 $X=1720 $Y=405 $D=9
M4 VGND S0 12 VNB nshort L=0.15 W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75000.2 a=0.063 p=1.14 mult=1 $X=2660 $Y=450 $D=9
M5 19 S0 23 VNB nshort L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75000.6 a=0.063 p=1.14 mult=1 $X=3600 $Y=485 $D=9
M6 24 12 19 VNB nshort L=0.15 W=0.42 AD=0.10795 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 m=1 r=2.8 sa=75000.6 sb=75000.2 a=0.063 p=1.14 mult=1 $X=4020 $Y=485 $D=9
M7 VGND A3 23 VNB nshort L=0.15 W=0.42 AD=0.0567 AS=0.1079 PD=0.69 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75000.6 a=0.063 p=1.14 mult=1 $X=4950 $Y=235 $D=9
M8 24 A2 VGND VNB nshort L=0.15 W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 m=1 r=2.8 sa=75000.6 sb=75000.2 a=0.063 p=1.14 mult=1 $X=5370 $Y=235 $D=9
M9 13 S1 VGND VNB nshort L=0.15 W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75000.2 a=0.063 p=1.14 mult=1 $X=6310 $Y=235 $D=9
M10 14 S1 19 VNB nshort L=0.15 W=0.42 AD=0.151025 AS=0.1092 PD=1.285 PS=1.36 NRD=78.564 NRS=0 m=1 r=2.8 sa=75000.2 sb=75000.7 a=0.063 p=1.14 mult=1 $X=7250 $Y=235 $D=9
M11 17 13 14 VNB nshort L=0.15 W=0.42 AD=0.1092 AS=0.151025 PD=1.36 PS=1.285 NRD=0 NRS=87.012 m=1 r=2.8 sa=75000.5 sb=75000.2 a=0.063 p=1.14 mult=1 $X=8015 $Y=485 $D=9
M12 X 14 VGND VNB nshort L=0.15 W=0.65 AD=0.169 AS=0.169 PD=1.82 PS=1.82 NRD=0 NRS=0 m=1 r=4.33333 sa=75000.2 sb=75000.2 a=0.0975 p=1.6 mult=1 $X=9115 $Y=235 $D=9
M13 VPWR A1 15 VPB phighvt L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75000.6 a=0.063 p=1.14 mult=1 $X=395 $Y=2065 $D=89
M14 16 A0 VPWR VPB phighvt L=0.15 W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 m=1 r=2.8 sa=75000.6 sb=75000.2 a=0.063 p=1.14 mult=1 $X=815 $Y=2065 $D=89
M15 17 12 15 VPB phighvt L=0.15 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75000.6 a=0.063 p=1.14 mult=1 $X=1755 $Y=1815 $D=89
M16 16 S0 17 VPB phighvt L=0.15 W=0.42 AD=0.1079 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 m=1 r=2.8 sa=75000.6 sb=75000.2 a=0.063 p=1.14 mult=1 $X=2175 $Y=1815 $D=89
M17 VPWR S0 12 VPB phighvt L=0.15 W=0.42 AD=0.1079 AS=0.1083 PD=1.36 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75000.2 a=0.063 p=1.14 mult=1 $X=3115 $Y=2065 $D=89
M18 19 S0 18 VPB phighvt L=0.15 W=0.42 AD=0.0567 AS=0.1079 PD=0.69 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75001 a=0.063 p=1.14 mult=1 $X=4045 $Y=1815 $D=89
M19 20 12 19 VPB phighvt L=0.15 W=0.42 AD=0.090125 AS=0.0567 PD=0.995 PS=0.69 NRD=74.8403 NRS=0 m=1 r=2.8 sa=75000.6 sb=75000.5 a=0.063 p=1.14 mult=1 $X=4465 $Y=1815 $D=89
M20 VPWR A3 20 VPB phighvt L=0.15 W=0.42 AD=0.0567 AS=0.090125 PD=0.69 PS=0.995 NRD=0 NRS=74.8403 m=1 r=2.8 sa=75000.5 sb=75000.6 a=0.063 p=1.14 mult=1 $X=4940 $Y=2065 $D=89
M21 18 A2 VPWR VPB phighvt L=0.15 W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 m=1 r=2.8 sa=75001 sb=75000.2 a=0.063 p=1.14 mult=1 $X=5360 $Y=2065 $D=89
M22 13 S1 VPWR VPB phighvt L=0.15 W=0.42 AD=0.1092 AS=0.1092 PD=1.36 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75000.2 a=0.063 p=1.14 mult=1 $X=6300 $Y=2065 $D=89
M23 14 S1 17 VPB phighvt L=0.15 W=0.42 AD=0.0920875 AS=0.1092 PD=0.99 PS=1.36 NRD=0 NRS=0 m=1 r=2.8 sa=75000.2 sb=75000.6 a=0.063 p=1.14 mult=1 $X=7240 $Y=2065 $D=89
M24 19 13 14 VPB phighvt L=0.15 W=0.42 AD=0.2688 AS=0.0920875 PD=2.12 PS=0.99 NRD=0 NRS=77.027 m=1 r=2.8 sa=75000.4 sb=75000.6 a=0.063 p=1.14 mult=1 $X=7725 $Y=1830 $D=89
M25 X 14 VPWR VPB phighvt L=0.15 W=1 AD=0.26 AS=0.26 PD=2.52 PS=2.52 NRD=0 NRS=0 m=1 r=6.66667 sa=75000.2 sb=75000.2 a=0.15 p=2.3 mult=1 $X=9115 $Y=1485 $D=89
.ENDS
***************************************
.SUBCKT ICV_78 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221
+ 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241
+ 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260 261
+ 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280 281
+ 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300 301
+ 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320 321
+ 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340 341
+ 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360 361
+ 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380 381
+ 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400 401
+ 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420 421
+ 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440 441
+ 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460 461
+ 462 463 464 465 466 467 468 469 470 471 479
** N=1989 EP=471 IP=16673 FDC=49046
*.SEEDPROM
X0 1 2 Dpar a=2090.79 p=1485.14 m=1 $[nwdiode] $X=5330 $Y=248825 $D=191
X1 1 2 Dpar a=2090.87 p=1485.04 m=1 $[nwdiode] $X=5330 $Y=254265 $D=191
X2 1 2 Dpar a=2091.03 p=1484.84 m=1 $[nwdiode] $X=5330 $Y=259705 $D=191
X3 1 2 Dpar a=2090.63 p=1485.34 m=1 $[nwdiode] $X=5330 $Y=265145 $D=191
X4 1 2 Dpar a=2090.87 p=1485.04 m=1 $[nwdiode] $X=5330 $Y=270585 $D=191
X5 1 2 Dpar a=2090.63 p=1485.34 m=1 $[nwdiode] $X=5330 $Y=276025 $D=191
X6 1 2 Dpar a=2090.71 p=1485.24 m=1 $[nwdiode] $X=5330 $Y=281465 $D=191
X7 1 2 Dpar a=2091.28 p=1484.54 m=1 $[nwdiode] $X=5330 $Y=286905 $D=191
X8 1 2 Dpar a=2091.36 p=1484.44 m=1 $[nwdiode] $X=5330 $Y=292345 $D=191
X9 1 2 Dpar a=2091.2 p=1484.64 m=1 $[nwdiode] $X=5330 $Y=297785 $D=191
X10 1 2 Dpar a=2090.47 p=1485.54 m=1 $[nwdiode] $X=5330 $Y=303225 $D=191
X11 1 2 Dpar a=2091.12 p=1484.74 m=1 $[nwdiode] $X=5330 $Y=308665 $D=191
X12 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 247520 1 0 $X=5330 $Y=244560
X13 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 247520 0 0 $X=5330 $Y=247280
X14 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 258400 1 0 $X=5330 $Y=255440
X15 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 258400 0 0 $X=5330 $Y=258160
X16 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 301920 1 0 $X=5330 $Y=298960
X17 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 301920 0 0 $X=5330 $Y=301680
X18 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 312800 1 0 $X=5330 $Y=309840
X19 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=6900 247520 1 0 $X=6710 $Y=244560
X20 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=6900 258400 1 0 $X=6710 $Y=255440
X21 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=6900 291040 1 0 $X=6710 $Y=288080
X22 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=19780 263840 0 0 $X=19590 $Y=263600
X23 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=20240 296480 1 0 $X=20050 $Y=293520
X24 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=24380 247520 1 0 $X=24190 $Y=244560
X25 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=27140 247520 1 0 $X=26950 $Y=244560
X26 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=32660 280160 1 0 $X=32470 $Y=277200
X27 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=42320 312800 1 0 $X=42130 $Y=309840
X28 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=48300 301920 1 0 $X=48110 $Y=298960
X29 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=69000 280160 1 0 $X=68810 $Y=277200
X30 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=71760 296480 1 0 $X=71570 $Y=293520
X31 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=93380 291040 1 0 $X=93190 $Y=288080
X32 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=95220 312800 1 0 $X=95030 $Y=309840
X33 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=104420 280160 1 0 $X=104230 $Y=277200
X34 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=119140 252960 1 0 $X=118950 $Y=250000
X35 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=130640 307360 0 0 $X=130450 $Y=307120
X36 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=147200 280160 1 0 $X=147010 $Y=277200
X37 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=160540 291040 1 0 $X=160350 $Y=288080
X38 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=160540 307360 1 0 $X=160350 $Y=304400
X39 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=164680 263840 0 0 $X=164490 $Y=263600
X40 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=175720 252960 0 0 $X=175530 $Y=252720
X41 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=188600 258400 1 0 $X=188410 $Y=255440
X42 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=196420 269280 0 0 $X=196230 $Y=269040
X43 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=201480 258400 1 0 $X=201290 $Y=255440
X44 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=218500 291040 0 0 $X=218310 $Y=290800
X45 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=223100 252960 0 0 $X=222910 $Y=252720
X46 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=224940 258400 1 0 $X=224750 $Y=255440
X47 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=230460 258400 0 0 $X=230270 $Y=258160
X48 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=234600 291040 0 0 $X=234410 $Y=290800
X49 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=239200 307360 0 0 $X=239010 $Y=307120
X50 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=252540 296480 0 0 $X=252350 $Y=296240
X51 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=256680 274720 0 0 $X=256490 $Y=274480
X52 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=285200 307360 1 0 $X=285010 $Y=304400
X53 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=300840 252960 1 0 $X=300650 $Y=250000
X54 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=300840 285600 1 0 $X=300650 $Y=282640
X55 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=314640 301920 0 0 $X=314450 $Y=301680
X56 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=315560 307360 1 0 $X=315370 $Y=304400
X57 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=328900 247520 1 0 $X=328710 $Y=244560
X58 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=336260 307360 1 0 $X=336070 $Y=304400
X59 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=355120 274720 1 0 $X=354930 $Y=271760
X60 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=380880 280160 1 0 $X=380690 $Y=277200
X61 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=387780 247520 0 0 $X=387590 $Y=247280
X62 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=396520 263840 1 0 $X=396330 $Y=260880
X63 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=407100 285600 1 0 $X=406910 $Y=282640
X64 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=408940 247520 1 0 $X=408750 $Y=244560
X65 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=412160 247520 0 0 $X=411970 $Y=247280
X66 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=417220 301920 0 0 $X=417030 $Y=301680
X67 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=451720 301920 0 0 $X=451530 $Y=301680
X68 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=488980 252960 1 0 $X=488790 $Y=250000
X69 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=497720 247520 0 0 $X=497530 $Y=247280
X70 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=511060 263840 0 0 $X=510870 $Y=263600
X71 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=515200 247520 0 0 $X=515010 $Y=247280
X72 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=537280 263840 0 0 $X=537090 $Y=263600
X73 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=553380 291040 1 0 $X=553190 $Y=288080
X74 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=553380 301920 1 0 $X=553190 $Y=298960
X75 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=603520 307360 1 0 $X=603330 $Y=304400
X76 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=630660 252960 0 0 $X=630470 $Y=252720
X77 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=637560 258400 1 0 $X=637370 $Y=255440
X78 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=642160 291040 0 0 $X=641970 $Y=290800
X79 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=645380 269280 0 0 $X=645190 $Y=269040
X80 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=657340 263840 1 0 $X=657150 $Y=260880
X81 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=669300 307360 0 0 $X=669110 $Y=307120
X82 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=679420 274720 0 0 $X=679230 $Y=274480
X83 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=690460 291040 0 0 $X=690270 $Y=290800
X84 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=705640 285600 1 0 $X=705450 $Y=282640
X85 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=715760 285600 1 0 $X=715570 $Y=282640
X86 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=735540 263840 0 0 $X=735350 $Y=263600
X87 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=741520 269280 1 0 $X=741330 $Y=266320
X88 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 312800 0 180 $X=742710 $Y=309840
X89 1 2 ICV_1 $T=5520 252960 1 0 $X=5330 $Y=250000
X90 1 2 ICV_1 $T=5520 263840 1 0 $X=5330 $Y=260880
X91 1 2 ICV_1 $T=5520 274720 1 0 $X=5330 $Y=271760
X92 1 2 ICV_1 $T=5520 280160 1 0 $X=5330 $Y=277200
X93 1 2 ICV_1 $T=5520 285600 1 0 $X=5330 $Y=282640
X94 1 2 ICV_1 $T=5520 291040 1 0 $X=5330 $Y=288080
X95 1 2 ICV_1 $T=5520 296480 1 0 $X=5330 $Y=293520
X96 1 2 ICV_1 $T=5520 307360 1 0 $X=5330 $Y=304400
X97 1 2 ICV_1 $T=744280 247520 0 180 $X=742710 $Y=244560
X98 1 2 ICV_1 $T=744280 252960 0 180 $X=742710 $Y=250000
X99 1 2 ICV_1 $T=744280 258400 0 180 $X=742710 $Y=255440
X100 1 2 ICV_1 $T=744280 263840 0 180 $X=742710 $Y=260880
X101 1 2 ICV_1 $T=744280 269280 0 180 $X=742710 $Y=266320
X102 1 2 ICV_1 $T=744280 274720 0 180 $X=742710 $Y=271760
X103 1 2 ICV_1 $T=744280 280160 0 180 $X=742710 $Y=277200
X104 1 2 ICV_1 $T=744280 285600 0 180 $X=742710 $Y=282640
X105 1 2 ICV_1 $T=744280 291040 0 180 $X=742710 $Y=288080
X106 1 2 ICV_1 $T=744280 296480 0 180 $X=742710 $Y=293520
X107 1 2 ICV_1 $T=744280 301920 0 180 $X=742710 $Y=298960
X108 1 2 ICV_1 $T=744280 307360 0 180 $X=742710 $Y=304400
X278 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17480 263840 1 0 $X=17290 $Y=260880
X279 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=20240 301920 1 0 $X=20050 $Y=298960
X280 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=34040 301920 0 0 $X=33850 $Y=301680
X281 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=45540 280160 1 0 $X=45350 $Y=277200
X282 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=48300 307360 1 0 $X=48110 $Y=304400
X283 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=48300 312800 1 0 $X=48110 $Y=309840
X284 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=69460 258400 0 0 $X=69270 $Y=258160
X285 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=73600 247520 1 0 $X=73410 $Y=244560
X286 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=74060 307360 1 0 $X=73870 $Y=304400
X287 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=90160 307360 0 0 $X=89970 $Y=307120
X288 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=104420 291040 1 0 $X=104230 $Y=288080
X289 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=118220 252960 0 0 $X=118030 $Y=252720
X290 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=143520 269280 0 0 $X=143330 $Y=269040
X291 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=153640 301920 0 0 $X=153450 $Y=301680
X292 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=160540 285600 1 0 $X=160350 $Y=282640
X293 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=160540 312800 1 0 $X=160350 $Y=309840
X294 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=171580 296480 0 0 $X=171390 $Y=296240
X295 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=178480 269280 1 0 $X=178290 $Y=266320
X296 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=185840 301920 1 0 $X=185650 $Y=298960
X297 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=216660 274720 1 0 $X=216470 $Y=271760
X298 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=216660 312800 1 0 $X=216470 $Y=309840
X299 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=226780 274720 1 0 $X=226590 $Y=271760
X300 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=242420 269280 1 0 $X=242230 $Y=266320
X301 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=242420 269280 0 0 $X=242230 $Y=269040
X302 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=255300 307360 1 0 $X=255110 $Y=304400
X303 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=272780 263840 1 0 $X=272590 $Y=260880
X304 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=286580 263840 0 0 $X=286390 $Y=263600
X305 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=293020 269280 1 0 $X=292830 $Y=266320
X306 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=298080 296480 1 0 $X=297890 $Y=293520
X307 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=328440 258400 0 0 $X=328250 $Y=258160
X308 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=351440 258400 0 0 $X=351250 $Y=258160
X309 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=356960 285600 1 0 $X=356770 $Y=282640
X310 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=382260 301920 1 0 $X=382070 $Y=298960
X311 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=385020 307360 1 0 $X=384830 $Y=304400
X312 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=396060 269280 0 0 $X=395870 $Y=269040
X313 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=410320 312800 1 0 $X=410130 $Y=309840
X314 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=413540 285600 0 0 $X=413350 $Y=285360
X315 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=424120 296480 0 0 $X=423930 $Y=296240
X316 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=438380 274720 1 0 $X=438190 $Y=271760
X317 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=448500 307360 0 0 $X=448310 $Y=307120
X318 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=469200 258400 1 0 $X=469010 $Y=255440
X319 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=480700 280160 0 0 $X=480510 $Y=279920
X320 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=483000 307360 0 0 $X=482810 $Y=307120
X321 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=490360 263840 0 0 $X=490170 $Y=263600
X322 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=508760 291040 0 0 $X=508570 $Y=290800
X323 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=522560 296480 1 0 $X=522370 $Y=293520
X324 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=532680 285600 1 0 $X=532490 $Y=282640
X325 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=533600 280160 1 0 $X=533410 $Y=277200
X326 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=539120 285600 0 0 $X=538930 $Y=285360
X327 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=539120 301920 0 0 $X=538930 $Y=301680
X328 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=581440 312800 1 0 $X=581250 $Y=309840
X329 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=592940 274720 0 0 $X=592750 $Y=274480
X330 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=611800 291040 1 0 $X=611610 $Y=288080
X331 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=616860 274720 0 0 $X=616670 $Y=274480
X332 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=621000 285600 0 0 $X=620810 $Y=285360
X333 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=637100 258400 0 0 $X=636910 $Y=258160
X334 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=644000 280160 1 0 $X=643810 $Y=277200
X335 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=644920 269280 1 0 $X=644730 $Y=266320
X336 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=648600 285600 0 0 $X=648410 $Y=285360
X337 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=658720 274720 0 0 $X=658530 $Y=274480
X338 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=676660 258400 0 0 $X=676470 $Y=258160
X339 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=677120 307360 0 0 $X=676930 $Y=307120
X340 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=695520 280160 0 0 $X=695330 $Y=279920
X341 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=707480 296480 0 0 $X=707290 $Y=296240
X342 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 296480 0 0 $X=740870 $Y=296240
X343 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 301920 1 0 $X=740870 $Y=298960
X344 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 301920 0 0 $X=740870 $Y=301680
X345 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 307360 0 0 $X=740870 $Y=307120
X346 1 2 ICV_3 $T=48300 285600 1 0 $X=48110 $Y=282640
X347 1 2 ICV_3 $T=59800 291040 1 0 $X=59610 $Y=288080
X348 1 2 ICV_3 $T=70380 269280 0 0 $X=70190 $Y=269040
X349 1 2 ICV_3 $T=87400 280160 0 0 $X=87210 $Y=279920
X350 1 2 ICV_3 $T=111320 307360 0 0 $X=111130 $Y=307120
X351 1 2 ICV_3 $T=129720 285600 0 0 $X=129530 $Y=285360
X352 1 2 ICV_3 $T=132480 247520 1 0 $X=132290 $Y=244560
X353 1 2 ICV_3 $T=146280 258400 1 0 $X=146090 $Y=255440
X354 1 2 ICV_3 $T=162840 296480 0 0 $X=162650 $Y=296240
X355 1 2 ICV_3 $T=187680 258400 0 0 $X=187490 $Y=258160
X356 1 2 ICV_3 $T=209760 291040 0 0 $X=209570 $Y=290800
X357 1 2 ICV_3 $T=241960 296480 0 0 $X=241770 $Y=296240
X358 1 2 ICV_3 $T=280140 252960 1 0 $X=279950 $Y=250000
X359 1 2 ICV_3 $T=340860 291040 1 0 $X=340670 $Y=288080
X360 1 2 ICV_3 $T=344080 269280 1 0 $X=343890 $Y=266320
X361 1 2 ICV_3 $T=368000 258400 0 0 $X=367810 $Y=258160
X362 1 2 ICV_3 $T=385020 291040 1 0 $X=384830 $Y=288080
X363 1 2 ICV_3 $T=391920 258400 0 0 $X=391730 $Y=258160
X364 1 2 ICV_3 $T=398820 269280 0 0 $X=398630 $Y=269040
X365 1 2 ICV_3 $T=412160 252960 0 0 $X=411970 $Y=252720
X366 1 2 ICV_3 $T=432400 291040 1 0 $X=432210 $Y=288080
X367 1 2 ICV_3 $T=438380 263840 1 0 $X=438190 $Y=260880
X368 1 2 ICV_3 $T=441140 274720 1 0 $X=440950 $Y=271760
X369 1 2 ICV_3 $T=450800 252960 1 0 $X=450610 $Y=250000
X370 1 2 ICV_3 $T=454940 307360 0 0 $X=454750 $Y=307120
X371 1 2 ICV_3 $T=466440 312800 1 0 $X=466250 $Y=309840
X372 1 2 ICV_3 $T=494960 291040 0 0 $X=494770 $Y=290800
X373 1 2 ICV_3 $T=501860 280160 0 0 $X=501670 $Y=279920
X374 1 2 ICV_3 $T=505080 307360 1 0 $X=504890 $Y=304400
X375 1 2 ICV_3 $T=508300 252960 0 0 $X=508110 $Y=252720
X376 1 2 ICV_3 $T=536360 307360 0 0 $X=536170 $Y=307120
X377 1 2 ICV_3 $T=546940 252960 1 0 $X=546750 $Y=250000
X378 1 2 ICV_3 $T=561200 252960 1 0 $X=561010 $Y=250000
X379 1 2 ICV_3 $T=564420 247520 0 0 $X=564230 $Y=247280
X380 1 2 ICV_3 $T=565340 263840 1 0 $X=565150 $Y=260880
X381 1 2 ICV_3 $T=574540 258400 1 0 $X=574350 $Y=255440
X382 1 2 ICV_3 $T=580060 291040 0 0 $X=579870 $Y=290800
X383 1 2 ICV_3 $T=609500 263840 1 0 $X=609310 $Y=260880
X384 1 2 ICV_3 $T=614100 301920 0 0 $X=613910 $Y=301680
X385 1 2 ICV_3 $T=623300 263840 0 0 $X=623110 $Y=263600
X386 1 2 ICV_3 $T=623300 291040 0 0 $X=623110 $Y=290800
X387 1 2 ICV_3 $T=644920 291040 1 0 $X=644730 $Y=288080
X388 1 2 ICV_3 $T=676660 291040 0 0 $X=676470 $Y=290800
X389 1 2 ICV_3 $T=693680 312800 1 0 $X=693490 $Y=309840
X390 1 2 ICV_3 $T=702420 301920 0 0 $X=702230 $Y=301680
X391 1 2 ICV_3 $T=707480 263840 0 0 $X=707290 $Y=263600
X392 1 2 ICV_3 $T=709780 301920 1 0 $X=709590 $Y=298960
X393 1 2 ICV_3 $T=718980 258400 1 0 $X=718790 $Y=255440
X394 1 2 ICV_3 $T=721740 307360 1 0 $X=721550 $Y=304400
X395 1 2 ICV_3 $T=724960 274720 0 0 $X=724770 $Y=274480
X396 1 2 ICV_3 $T=735540 258400 0 0 $X=735350 $Y=258160
X397 1 2 ICV_3 $T=735540 274720 0 0 $X=735350 $Y=274480
X398 1 2 ICV_3 $T=735540 280160 0 0 $X=735350 $Y=279920
X399 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=27140 274720 1 0 $X=26950 $Y=271760
X400 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=71300 301920 0 0 $X=71110 $Y=301680
X401 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=78660 291040 0 0 $X=78470 $Y=290800
X402 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=90160 269280 0 0 $X=89970 $Y=269040
X403 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=92920 263840 1 0 $X=92730 $Y=260880
X404 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=104420 263840 1 0 $X=104230 $Y=260880
X405 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=111780 296480 0 0 $X=111590 $Y=296240
X406 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=118220 269280 0 0 $X=118030 $Y=269040
X407 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=122360 307360 1 0 $X=122170 $Y=304400
X408 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=132480 291040 1 0 $X=132290 $Y=288080
X409 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=132480 301920 1 0 $X=132290 $Y=298960
X410 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=143060 263840 0 0 $X=142870 $Y=263600
X411 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=155020 247520 0 0 $X=154830 $Y=247280
X412 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=157320 274720 1 0 $X=157130 $Y=271760
X413 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=176180 312800 1 0 $X=175990 $Y=309840
X414 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=205620 274720 1 0 $X=205430 $Y=271760
X415 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=224020 301920 1 0 $X=223830 $Y=298960
X416 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=260820 274720 1 0 $X=260630 $Y=271760
X417 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=272780 258400 1 0 $X=272590 $Y=255440
X418 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=283360 280160 0 0 $X=283170 $Y=279920
X419 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=284280 274720 1 0 $X=284090 $Y=271760
X420 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=287040 280160 1 0 $X=286850 $Y=277200
X421 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=300840 312800 1 0 $X=300650 $Y=309840
X422 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=308200 291040 1 0 $X=308010 $Y=288080
X423 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=310500 258400 1 0 $X=310310 $Y=255440
X424 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=325680 296480 1 0 $X=325490 $Y=293520
X425 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=325680 312800 1 0 $X=325490 $Y=309840
X426 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=335340 285600 0 0 $X=335150 $Y=285360
X427 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=337640 274720 1 0 $X=337450 $Y=271760
X428 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=340860 296480 1 0 $X=340670 $Y=293520
X429 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=344540 263840 1 0 $X=344350 $Y=260880
X430 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=361100 274720 1 0 $X=360910 $Y=271760
X431 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=364780 269280 1 0 $X=364590 $Y=266320
X432 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=370760 285600 0 0 $X=370570 $Y=285360
X433 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=385020 247520 1 0 $X=384830 $Y=244560
X434 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=395600 263840 0 0 $X=395410 $Y=263600
X435 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=398820 274720 0 0 $X=398630 $Y=274480
X436 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=418600 274720 1 0 $X=418410 $Y=271760
X437 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=426880 247520 0 0 $X=426690 $Y=247280
X438 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=448500 263840 1 0 $X=448310 $Y=260880
X439 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=473340 252960 1 0 $X=473150 $Y=250000
X440 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=489900 291040 1 0 $X=489710 $Y=288080
X441 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=494040 296480 1 0 $X=493850 $Y=293520
X442 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=511060 280160 0 0 $X=510870 $Y=279920
X443 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=511060 285600 0 0 $X=510870 $Y=285360
X444 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=525320 258400 1 0 $X=525130 $Y=255440
X445 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=554300 301920 0 0 $X=554110 $Y=301680
X446 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=559820 307360 1 0 $X=559630 $Y=304400
X447 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=569940 269280 1 0 $X=569750 $Y=266320
X448 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=578680 285600 0 0 $X=578490 $Y=285360
X449 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=581440 247520 1 0 $X=581250 $Y=244560
X450 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=587880 301920 0 0 $X=587690 $Y=301680
X451 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=592020 258400 0 0 $X=591830 $Y=258160
X452 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=601680 269280 1 0 $X=601490 $Y=266320
X453 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=607660 269280 0 0 $X=607470 $Y=269040
X454 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=637560 285600 1 0 $X=637370 $Y=282640
X455 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=647680 274720 1 0 $X=647490 $Y=271760
X456 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=648140 280160 0 0 $X=647950 $Y=279920
X457 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=649060 312800 1 0 $X=648870 $Y=309840
X458 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=656880 296480 0 0 $X=656690 $Y=296240
X459 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=662400 301920 1 0 $X=662210 $Y=298960
X460 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=665620 307360 1 0 $X=665430 $Y=304400
X461 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=679420 269280 0 0 $X=679230 $Y=269040
X462 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=686320 307360 1 0 $X=686130 $Y=304400
X463 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=722200 296480 0 0 $X=722010 $Y=296240
X464 1 2 ICV_4 $T=18860 301920 0 0 $X=18670 $Y=301680
X465 1 2 ICV_4 $T=22540 274720 1 0 $X=22350 $Y=271760
X466 1 2 ICV_4 $T=33120 285600 1 0 $X=32930 $Y=282640
X467 1 2 ICV_4 $T=57040 307360 0 0 $X=56850 $Y=307120
X468 1 2 ICV_4 $T=86480 263840 0 0 $X=86290 $Y=263600
X469 1 2 ICV_4 $T=114540 247520 1 0 $X=114350 $Y=244560
X470 1 2 ICV_4 $T=142600 301920 0 0 $X=142410 $Y=301680
X471 1 2 ICV_4 $T=170660 285600 0 0 $X=170470 $Y=285360
X472 1 2 ICV_4 $T=269100 247520 1 0 $X=268910 $Y=244560
X473 1 2 ICV_4 $T=280140 258400 1 0 $X=279950 $Y=255440
X474 1 2 ICV_4 $T=297160 307360 1 0 $X=296970 $Y=304400
X475 1 2 ICV_4 $T=350060 307360 0 0 $X=349870 $Y=307120
X476 1 2 ICV_4 $T=361100 291040 1 0 $X=360910 $Y=288080
X477 1 2 ICV_4 $T=385020 285600 1 0 $X=384830 $Y=282640
X478 1 2 ICV_4 $T=395600 291040 1 0 $X=395410 $Y=288080
X479 1 2 ICV_4 $T=442980 307360 0 0 $X=442790 $Y=307120
X480 1 2 ICV_4 $T=465980 263840 0 0 $X=465790 $Y=263600
X481 1 2 ICV_4 $T=493580 274720 1 0 $X=493390 $Y=271760
X482 1 2 ICV_4 $T=548780 296480 0 0 $X=548590 $Y=296240
X483 1 2 ICV_4 $T=563500 301920 0 0 $X=563310 $Y=301680
X484 1 2 ICV_4 $T=563500 307360 0 0 $X=563310 $Y=307120
X485 1 2 ICV_4 $T=647680 274720 0 0 $X=647490 $Y=274480
X486 1 2 ICV_4 $T=690000 258400 1 0 $X=689810 $Y=255440
X487 1 2 ICV_4 $T=700120 280160 1 0 $X=699930 $Y=277200
X488 1 2 ICV_4 $T=703800 258400 0 0 $X=703610 $Y=258160
X489 1 2 ICV_4 $T=704260 252960 1 0 $X=704070 $Y=250000
X490 1 2 ICV_4 $T=726340 247520 1 0 $X=726150 $Y=244560
X491 1 2 ICV_4 $T=739680 285600 0 0 $X=739490 $Y=285360
X492 1 2 ICV_4 $T=739680 291040 0 0 $X=739490 $Y=290800
X493 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=28520 258400 1 0 $X=28330 $Y=255440
X494 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=42320 274720 0 0 $X=42130 $Y=274480
X495 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=45540 258400 0 0 $X=45350 $Y=258160
X496 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=46460 296480 0 0 $X=46270 $Y=296240
X497 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=57500 274720 0 0 $X=57310 $Y=274480
X498 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=59800 280160 1 0 $X=59610 $Y=277200
X499 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=72220 274720 0 0 $X=72030 $Y=274480
X500 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=81880 296480 1 0 $X=81690 $Y=293520
X501 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=90160 291040 0 0 $X=89970 $Y=290800
X502 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=100280 296480 1 0 $X=100090 $Y=293520
X503 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=108560 296480 1 0 $X=108370 $Y=293520
X504 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=109940 247520 0 0 $X=109750 $Y=247280
X505 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=128340 258400 1 0 $X=128150 $Y=255440
X506 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=128340 285600 1 0 $X=128150 $Y=282640
X507 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=132480 263840 1 0 $X=132290 $Y=260880
X508 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=132480 307360 1 0 $X=132290 $Y=304400
X509 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=134780 252960 0 0 $X=134590 $Y=252720
X510 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=139840 252960 1 0 $X=139650 $Y=250000
X511 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=139840 312800 1 0 $X=139650 $Y=309840
X512 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=162840 291040 0 0 $X=162650 $Y=290800
X513 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=170200 301920 0 0 $X=170010 $Y=301680
X514 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=176180 280160 1 0 $X=175990 $Y=277200
X515 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=184460 269280 1 0 $X=184270 $Y=266320
X516 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=184460 274720 1 0 $X=184270 $Y=271760
X517 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=188600 280160 1 0 $X=188410 $Y=277200
X518 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=198260 307360 0 0 $X=198070 $Y=307120
X519 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=200100 263840 1 0 $X=199910 $Y=260880
X520 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=206540 301920 1 0 $X=206350 $Y=298960
X521 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=212520 263840 0 0 $X=212330 $Y=263600
X522 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=212520 274720 1 0 $X=212330 $Y=271760
X523 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=226320 307360 0 0 $X=226130 $Y=307120
X524 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=244720 258400 1 0 $X=244530 $Y=255440
X525 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=250240 280160 0 0 $X=250050 $Y=279920
X526 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=254380 307360 0 0 $X=254190 $Y=307120
X527 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=258520 252960 0 0 $X=258330 $Y=252720
X528 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=258520 280160 0 0 $X=258330 $Y=279920
X529 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=262660 274720 0 0 $X=262470 $Y=274480
X530 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=270940 291040 0 0 $X=270750 $Y=290800
X531 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=278300 296480 0 0 $X=278110 $Y=296240
X532 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=282440 269280 0 0 $X=282250 $Y=269040
X533 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=282900 296480 1 0 $X=282710 $Y=293520
X534 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=296700 252960 1 0 $X=296510 $Y=250000
X535 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=300840 296480 1 0 $X=300650 $Y=293520
X536 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=309580 296480 1 0 $X=309390 $Y=293520
X537 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=314640 274720 0 0 $X=314450 $Y=274480
X538 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=320160 269280 0 0 $X=319970 $Y=269040
X539 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=329820 301920 0 0 $X=329630 $Y=301680
X540 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=352820 247520 0 0 $X=352630 $Y=247280
X541 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=352820 252960 1 0 $X=352630 $Y=250000
X542 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=365700 258400 1 0 $X=365510 $Y=255440
X543 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=366620 301920 0 0 $X=366430 $Y=301680
X544 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=401580 296480 1 0 $X=401390 $Y=293520
X545 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=408480 263840 1 0 $X=408290 $Y=260880
X546 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=413080 307360 1 0 $X=412890 $Y=304400
X547 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=421360 291040 1 0 $X=421170 $Y=288080
X548 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=422740 307360 0 0 $X=422550 $Y=307120
X549 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=440220 263840 0 0 $X=440030 $Y=263600
X550 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=445280 296480 1 0 $X=445090 $Y=293520
X551 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=448040 301920 0 0 $X=447850 $Y=301680
X552 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=449420 291040 0 0 $X=449230 $Y=290800
X553 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=451260 312800 1 0 $X=451070 $Y=309840
X554 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=454940 263840 0 0 $X=454750 $Y=263600
X555 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=459540 291040 0 0 $X=459350 $Y=290800
X556 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=477480 274720 1 0 $X=477290 $Y=271760
X557 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=478860 252960 0 0 $X=478670 $Y=252720
X558 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=478860 291040 1 0 $X=478670 $Y=288080
X559 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=497260 280160 1 0 $X=497070 $Y=277200
X560 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=519800 307360 1 0 $X=519610 $Y=304400
X561 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=521640 301920 0 0 $X=521450 $Y=301680
X562 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=536820 291040 1 0 $X=536630 $Y=288080
X563 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=548780 291040 1 0 $X=548590 $Y=288080
X564 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=549240 247520 0 0 $X=549050 $Y=247280
X565 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=549240 285600 1 0 $X=549050 $Y=282640
X566 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=552460 274720 0 0 $X=552270 $Y=274480
X567 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=553380 258400 1 0 $X=553190 $Y=255440
X568 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=557520 274720 0 0 $X=557330 $Y=274480
X569 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=582820 252960 0 0 $X=582630 $Y=252720
X570 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=591100 269280 0 0 $X=590910 $Y=269040
X571 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=593860 280160 1 0 $X=593670 $Y=277200
X572 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=599840 307360 1 0 $X=599650 $Y=304400
X573 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=600760 247520 1 0 $X=600570 $Y=244560
X574 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=604900 291040 1 0 $X=604710 $Y=288080
X575 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=605360 296480 1 0 $X=605170 $Y=293520
X576 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=609960 296480 0 0 $X=609770 $Y=296240
X577 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=617780 296480 0 0 $X=617590 $Y=296240
X578 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=629740 263840 0 0 $X=629550 $Y=263600
X579 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=629740 291040 0 0 $X=629550 $Y=290800
X580 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=630660 285600 0 0 $X=630470 $Y=285360
X581 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=631120 247520 0 0 $X=630930 $Y=247280
X582 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=632960 252960 1 0 $X=632770 $Y=250000
X583 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=636180 296480 0 0 $X=635990 $Y=296240
X584 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=645840 301920 0 0 $X=645650 $Y=301680
X585 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=657340 280160 1 0 $X=657150 $Y=277200
X586 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=664240 296480 0 0 $X=664050 $Y=296240
X587 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=673900 301920 0 0 $X=673710 $Y=301680
X588 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=675280 274720 0 0 $X=675090 $Y=274480
X589 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=683560 247520 0 0 $X=683370 $Y=247280
X590 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=686780 291040 0 0 $X=686590 $Y=290800
X591 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=694140 263840 0 0 $X=693950 $Y=263600
X592 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=698280 301920 1 0 $X=698090 $Y=298960
X593 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=703340 269280 0 0 $X=703150 $Y=269040
X594 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=707480 291040 0 0 $X=707290 $Y=290800
X595 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=717600 312800 1 0 $X=717410 $Y=309840
X596 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=725880 252960 1 0 $X=725690 $Y=250000
X597 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=730020 307360 0 0 $X=729830 $Y=307120
X598 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=731400 274720 0 0 $X=731210 $Y=274480
X599 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=738300 291040 1 0 $X=738110 $Y=288080
X600 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=738300 296480 1 0 $X=738110 $Y=293520
X601 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=738760 307360 1 0 $X=738570 $Y=304400
X602 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 274720 1 0 $X=6710 $Y=271760
X603 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=12420 274720 1 0 $X=12230 $Y=271760
X604 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=13340 312800 1 0 $X=13150 $Y=309840
X605 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=25300 258400 0 0 $X=25110 $Y=258160
X606 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=76360 291040 1 0 $X=76170 $Y=288080
X607 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=81420 258400 1 0 $X=81230 $Y=255440
X608 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=322000 263840 1 0 $X=321810 $Y=260880
X609 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=339940 247520 1 0 $X=339750 $Y=244560
X610 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=350520 269280 1 0 $X=350330 $Y=266320
X611 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=370760 247520 0 0 $X=370570 $Y=247280
X612 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=406640 269280 1 0 $X=406450 $Y=266320
X613 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=432860 274720 1 0 $X=432670 $Y=271760
X614 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=434240 285600 1 0 $X=434050 $Y=282640
X615 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=447580 280160 0 0 $X=447390 $Y=279920
X616 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=462300 291040 1 0 $X=462110 $Y=288080
X617 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=518880 301920 1 0 $X=518690 $Y=298960
X618 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=523480 291040 0 0 $X=523290 $Y=290800
X619 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=543260 296480 0 0 $X=543070 $Y=296240
X620 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=560280 296480 0 0 $X=560090 $Y=296240
X621 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=574540 291040 0 0 $X=574350 $Y=290800
X622 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=582820 296480 0 0 $X=582630 $Y=296240
X623 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=588340 296480 0 0 $X=588150 $Y=296240
X624 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=593860 291040 1 0 $X=593670 $Y=288080
X625 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=609960 274720 0 0 $X=609770 $Y=274480
X626 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=630200 296480 1 0 $X=630010 $Y=293520
X627 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=630660 296480 0 0 $X=630470 $Y=296240
X628 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=634800 301920 0 0 $X=634610 $Y=301680
X629 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=637560 301920 1 0 $X=637370 $Y=298960
X630 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=637560 307360 1 0 $X=637370 $Y=304400
X631 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=640320 301920 0 0 $X=640130 $Y=301680
X632 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=643080 301920 1 0 $X=642890 $Y=298960
X633 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=651360 296480 0 0 $X=651170 $Y=296240
X634 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=653200 296480 1 0 $X=653010 $Y=293520
X635 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=658720 296480 1 0 $X=658530 $Y=293520
X636 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=665620 291040 1 0 $X=665430 $Y=288080
X637 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=672980 296480 0 0 $X=672790 $Y=296240
X638 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=679420 296480 0 0 $X=679230 $Y=296240
X639 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=684940 296480 0 0 $X=684750 $Y=296240
X640 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=686320 296480 1 0 $X=686130 $Y=293520
X641 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=690460 296480 0 0 $X=690270 $Y=296240
X642 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=693680 296480 1 0 $X=693490 $Y=293520
X643 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=695980 296480 0 0 $X=695790 $Y=296240
X644 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=699200 296480 1 0 $X=699010 $Y=293520
X645 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=701500 296480 0 0 $X=701310 $Y=296240
X646 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=704720 296480 1 0 $X=704530 $Y=293520
X647 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=710240 296480 1 0 $X=710050 $Y=293520
X648 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=715760 296480 1 0 $X=715570 $Y=293520
X649 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=726340 301920 0 0 $X=726150 $Y=301680
X650 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=729100 296480 0 0 $X=728910 $Y=296240
X651 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=730020 301920 1 0 $X=729830 $Y=298960
X652 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=733240 307360 1 0 $X=733050 $Y=304400
X653 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 296480 0 0 $X=735350 $Y=296240
X654 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 301920 1 0 $X=735350 $Y=298960
X655 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 301920 0 0 $X=735350 $Y=301680
X656 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 307360 0 0 $X=735350 $Y=307120
X657 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=736460 312800 1 0 $X=736270 $Y=309840
X658 1 2 590 585 2 16 1 sky130_fd_sc_hd__ebufn_2 $T=46460 291040 0 0 $X=46270 $Y=290800
X659 1 2 591 45 2 30 1 sky130_fd_sc_hd__ebufn_2 $T=48300 252960 1 0 $X=48110 $Y=250000
X660 1 2 611 47 2 33 1 sky130_fd_sc_hd__ebufn_2 $T=50140 307360 1 0 $X=49950 $Y=304400
X661 1 2 632 641 2 13 1 sky130_fd_sc_hd__ebufn_2 $T=63480 280160 1 0 $X=63290 $Y=277200
X662 1 2 671 676 2 18 1 sky130_fd_sc_hd__ebufn_2 $T=82340 263840 0 0 $X=82150 $Y=263600
X663 1 2 681 642 2 18 1 sky130_fd_sc_hd__ebufn_2 $T=85100 296480 0 0 $X=84910 $Y=296240
X664 1 2 698 693 2 19 1 sky130_fd_sc_hd__ebufn_2 $T=92000 301920 0 0 $X=91810 $Y=301680
X665 1 2 703 684 2 34 1 sky130_fd_sc_hd__ebufn_2 $T=93840 291040 0 0 $X=93650 $Y=290800
X666 1 2 716 74 2 16 1 sky130_fd_sc_hd__ebufn_2 $T=98900 258400 0 0 $X=98710 $Y=258160
X667 1 2 725 693 2 34 1 sky130_fd_sc_hd__ebufn_2 $T=104420 301920 1 0 $X=104230 $Y=298960
X668 1 2 82 77 2 13 1 sky130_fd_sc_hd__ebufn_2 $T=104420 312800 1 0 $X=104230 $Y=309840
X669 1 2 758 718 2 17 1 sky130_fd_sc_hd__ebufn_2 $T=120060 252960 0 0 $X=119870 $Y=252720
X670 1 2 93 77 2 34 1 sky130_fd_sc_hd__ebufn_2 $T=120060 312800 1 0 $X=119870 $Y=309840
X671 1 2 756 757 2 13 1 sky130_fd_sc_hd__ebufn_2 $T=124660 296480 0 0 $X=124470 $Y=296240
X672 1 2 781 772 2 17 1 sky130_fd_sc_hd__ebufn_2 $T=132020 285600 0 0 $X=131830 $Y=285360
X673 1 2 786 757 2 33 1 sky130_fd_sc_hd__ebufn_2 $T=135240 301920 1 0 $X=135050 $Y=298960
X674 1 2 774 779 2 34 1 sky130_fd_sc_hd__ebufn_2 $T=139840 285600 1 0 $X=139650 $Y=282640
X675 1 2 800 779 2 19 1 sky130_fd_sc_hd__ebufn_2 $T=141680 274720 1 0 $X=141490 $Y=271760
X676 1 2 802 811 2 34 1 sky130_fd_sc_hd__ebufn_2 $T=146280 258400 0 0 $X=146090 $Y=258160
X677 1 2 820 824 2 18 1 sky130_fd_sc_hd__ebufn_2 $T=151800 285600 0 0 $X=151610 $Y=285360
X678 1 2 844 89 2 33 1 sky130_fd_sc_hd__ebufn_2 $T=162380 312800 1 0 $X=162190 $Y=309840
X679 1 2 878 862 2 123 1 sky130_fd_sc_hd__ebufn_2 $T=180320 269280 1 0 $X=180130 $Y=266320
X680 1 2 901 139 2 123 1 sky130_fd_sc_hd__ebufn_2 $T=191360 263840 0 0 $X=191170 $Y=263600
X681 1 2 890 119 2 131 1 sky130_fd_sc_hd__ebufn_2 $T=195960 301920 0 0 $X=195770 $Y=301680
X682 1 2 931 921 2 122 1 sky130_fd_sc_hd__ebufn_2 $T=208380 274720 1 0 $X=208190 $Y=271760
X683 1 2 959 139 2 122 1 sky130_fd_sc_hd__ebufn_2 $T=222640 301920 0 0 $X=222450 $Y=301680
X684 1 2 961 954 2 123 1 sky130_fd_sc_hd__ebufn_2 $T=225860 280160 0 0 $X=225670 $Y=279920
X685 1 2 974 975 2 131 1 sky130_fd_sc_hd__ebufn_2 $T=226780 301920 1 0 $X=226590 $Y=298960
X686 1 2 981 973 2 122 1 sky130_fd_sc_hd__ebufn_2 $T=228620 274720 1 0 $X=228430 $Y=271760
X687 1 2 972 154 2 121 1 sky130_fd_sc_hd__ebufn_2 $T=230460 307360 1 0 $X=230270 $Y=304400
X688 1 2 996 954 2 121 1 sky130_fd_sc_hd__ebufn_2 $T=237820 285600 1 0 $X=237630 $Y=282640
X689 1 2 1006 975 2 117 1 sky130_fd_sc_hd__ebufn_2 $T=240120 296480 1 0 $X=239930 $Y=293520
X690 1 2 1004 986 2 123 1 sky130_fd_sc_hd__ebufn_2 $T=244720 258400 0 0 $X=244530 $Y=258160
X691 1 2 165 164 2 135 1 sky130_fd_sc_hd__ebufn_2 $T=258520 301920 0 0 $X=258330 $Y=301680
X692 1 2 1038 986 2 131 1 sky130_fd_sc_hd__ebufn_2 $T=260820 258400 1 0 $X=260630 $Y=255440
X693 1 2 1058 1059 2 136 1 sky130_fd_sc_hd__ebufn_2 $T=266340 274720 0 0 $X=266150 $Y=274480
X694 1 2 1072 1053 2 122 1 sky130_fd_sc_hd__ebufn_2 $T=274620 263840 1 0 $X=274430 $Y=260880
X695 1 2 1091 168 2 131 1 sky130_fd_sc_hd__ebufn_2 $T=281980 307360 0 0 $X=281790 $Y=307120
X696 1 2 1119 1123 2 131 1 sky130_fd_sc_hd__ebufn_2 $T=296240 280160 1 0 $X=296050 $Y=277200
X697 1 2 1121 1105 2 131 1 sky130_fd_sc_hd__ebufn_2 $T=296240 291040 1 0 $X=296050 $Y=288080
X698 1 2 1125 159 2 122 1 sky130_fd_sc_hd__ebufn_2 $T=301760 252960 0 0 $X=301570 $Y=252720
X699 1 2 1151 1124 2 134 1 sky130_fd_sc_hd__ebufn_2 $T=313260 296480 1 0 $X=313070 $Y=293520
X700 1 2 1164 1146 2 131 1 sky130_fd_sc_hd__ebufn_2 $T=324300 269280 1 0 $X=324110 $Y=266320
X701 1 2 1212 1183 2 121 1 sky130_fd_sc_hd__ebufn_2 $T=346380 269280 1 0 $X=346190 $Y=266320
X702 1 2 1235 1240 2 257 1 sky130_fd_sc_hd__ebufn_2 $T=363860 274720 1 0 $X=363670 $Y=271760
X703 1 2 1276 1277 2 257 1 sky130_fd_sc_hd__ebufn_2 $T=380420 269280 1 0 $X=380230 $Y=266320
X704 1 2 1295 1299 2 178 1 sky130_fd_sc_hd__ebufn_2 $T=391000 301920 1 0 $X=390810 $Y=298960
X705 1 2 1300 1273 2 257 1 sky130_fd_sc_hd__ebufn_2 $T=394220 258400 0 0 $X=394030 $Y=258160
X706 1 2 1324 1299 2 186 1 sky130_fd_sc_hd__ebufn_2 $T=408020 291040 1 0 $X=407830 $Y=288080
X707 1 2 1337 1312 2 229 1 sky130_fd_sc_hd__ebufn_2 $T=413080 274720 0 0 $X=412890 $Y=274480
X708 1 2 1398 1387 2 186 1 sky130_fd_sc_hd__ebufn_2 $T=441140 296480 1 0 $X=440950 $Y=293520
X709 1 2 1419 319 2 257 1 sky130_fd_sc_hd__ebufn_2 $T=453100 252960 1 0 $X=452910 $Y=250000
X710 1 2 1424 1375 2 262 1 sky130_fd_sc_hd__ebufn_2 $T=454940 258400 0 0 $X=454750 $Y=258160
X711 1 2 1446 1449 2 178 1 sky130_fd_sc_hd__ebufn_2 $T=464600 307360 1 0 $X=464410 $Y=304400
X712 1 2 1469 1470 2 201 1 sky130_fd_sc_hd__ebufn_2 $T=476100 252960 1 0 $X=475910 $Y=250000
X713 1 2 1480 1449 2 199 1 sky130_fd_sc_hd__ebufn_2 $T=483000 301920 0 0 $X=482810 $Y=301680
X714 1 2 1489 334 2 188 1 sky130_fd_sc_hd__ebufn_2 $T=484840 307360 0 0 $X=484650 $Y=307120
X715 1 2 1493 1470 2 257 1 sky130_fd_sc_hd__ebufn_2 $T=488980 258400 0 0 $X=488790 $Y=258160
X716 1 2 1494 1484 2 233 1 sky130_fd_sc_hd__ebufn_2 $T=489440 274720 1 0 $X=489250 $Y=271760
X717 1 2 1495 1484 2 229 1 sky130_fd_sc_hd__ebufn_2 $T=497720 280160 0 0 $X=497530 $Y=279920
X718 1 2 1516 1484 2 262 1 sky130_fd_sc_hd__ebufn_2 $T=498640 269280 1 0 $X=498450 $Y=266320
X719 1 2 1536 1504 2 180 1 sky130_fd_sc_hd__ebufn_2 $T=507380 307360 1 0 $X=507190 $Y=304400
X720 1 2 1586 1583 2 382 1 sky130_fd_sc_hd__ebufn_2 $T=539120 296480 0 0 $X=538930 $Y=296240
X721 1 2 1598 1583 2 328 1 sky130_fd_sc_hd__ebufn_2 $T=540960 285600 0 0 $X=540770 $Y=285360
X722 1 2 1596 394 2 370 1 sky130_fd_sc_hd__ebufn_2 $T=540960 301920 0 0 $X=540770 $Y=301680
X723 1 2 1593 1576 2 306 1 sky130_fd_sc_hd__ebufn_2 $T=542800 252960 1 0 $X=542610 $Y=250000
X724 1 2 1634 1620 2 341 1 sky130_fd_sc_hd__ebufn_2 $T=559820 280160 0 0 $X=559630 $Y=279920
X725 1 2 1670 415 2 263 1 sky130_fd_sc_hd__ebufn_2 $T=576840 252960 1 0 $X=576650 $Y=250000
X726 1 2 419 415 2 201 1 sky130_fd_sc_hd__ebufn_2 $T=576840 258400 1 0 $X=576650 $Y=255440
X727 1 2 1661 1635 2 341 1 sky130_fd_sc_hd__ebufn_2 $T=578680 252960 0 0 $X=578490 $Y=252720
X728 1 2 1666 1656 2 400 1 sky130_fd_sc_hd__ebufn_2 $T=578680 296480 0 0 $X=578490 $Y=296240
X729 1 2 1680 1681 2 201 1 sky130_fd_sc_hd__ebufn_2 $T=586960 269280 0 0 $X=586770 $Y=269040
X730 1 2 1673 1681 2 229 1 sky130_fd_sc_hd__ebufn_2 $T=589720 280160 1 0 $X=589530 $Y=277200
X731 1 2 1709 1688 2 260 1 sky130_fd_sc_hd__ebufn_2 $T=596160 263840 1 0 $X=595970 $Y=260880
X732 1 2 432 430 2 400 1 sky130_fd_sc_hd__ebufn_2 $T=609960 301920 0 0 $X=609770 $Y=301680
X733 1 2 1742 1739 2 382 1 sky130_fd_sc_hd__ebufn_2 $T=613640 296480 0 0 $X=613450 $Y=296240
X734 1 2 1762 1730 2 260 1 sky130_fd_sc_hd__ebufn_2 $T=625600 263840 0 0 $X=625410 $Y=263600
X735 1 2 1766 1739 2 337 1 sky130_fd_sc_hd__ebufn_2 $T=625600 291040 0 0 $X=625410 $Y=290800
X736 1 2 1771 435 2 201 1 sky130_fd_sc_hd__ebufn_2 $T=628820 252960 1 0 $X=628630 $Y=250000
X737 1 2 1798 440 2 361 1 sky130_fd_sc_hd__ebufn_2 $T=643080 307360 1 0 $X=642890 $Y=304400
X738 1 2 1815 1813 2 229 1 sky130_fd_sc_hd__ebufn_2 $T=646760 269280 1 0 $X=646570 $Y=266320
X739 1 2 1814 1804 2 382 1 sky130_fd_sc_hd__ebufn_2 $T=649060 296480 1 0 $X=648870 $Y=293520
X740 1 2 1823 1813 2 201 1 sky130_fd_sc_hd__ebufn_2 $T=656420 269280 0 0 $X=656230 $Y=269040
X741 1 2 1843 1844 2 382 1 sky130_fd_sc_hd__ebufn_2 $T=661020 280160 1 0 $X=660830 $Y=277200
X742 1 2 1833 1812 2 260 1 sky130_fd_sc_hd__ebufn_2 $T=662860 258400 0 0 $X=662670 $Y=258160
X743 1 2 1871 1844 2 337 1 sky130_fd_sc_hd__ebufn_2 $T=674820 280160 0 0 $X=674630 $Y=279920
X744 1 2 1883 1844 2 306 1 sky130_fd_sc_hd__ebufn_2 $T=682180 269280 0 0 $X=681990 $Y=269040
X745 1 2 1887 1859 2 372 1 sky130_fd_sc_hd__ebufn_2 $T=685860 258400 1 0 $X=685670 $Y=255440
X746 1 2 1888 1844 2 348 1 sky130_fd_sc_hd__ebufn_2 $T=686780 280160 1 0 $X=686590 $Y=277200
X747 1 2 1924 1904 2 328 1 sky130_fd_sc_hd__ebufn_2 $T=707480 280160 0 0 $X=707290 $Y=279920
X748 1 2 1938 1926 2 361 1 sky130_fd_sc_hd__ebufn_2 $T=709320 296480 0 0 $X=709130 $Y=296240
X749 1 2 1968 1950 2 372 1 sky130_fd_sc_hd__ebufn_2 $T=724960 296480 0 0 $X=724770 $Y=296240
X750 1 2 1958 1926 2 373 1 sky130_fd_sc_hd__ebufn_2 $T=725880 307360 0 0 $X=725690 $Y=307120
X751 1 2 1971 1965 2 341 1 sky130_fd_sc_hd__ebufn_2 $T=727260 274720 0 0 $X=727070 $Y=274480
X877 1 2 22 23 19 ICV_6 $T=19780 247520 1 0 $X=19590 $Y=244560
X878 1 2 635 47 16 ICV_6 $T=61640 307360 0 0 $X=61450 $Y=307120
X879 1 2 726 693 18 ICV_6 $T=103960 296480 1 0 $X=103770 $Y=293520
X880 1 2 804 811 30 ICV_6 $T=145820 263840 0 0 $X=145630 $Y=263600
X881 1 2 118 119 123 ICV_6 $T=173880 307360 0 0 $X=173690 $Y=307120
X882 1 2 896 116 136 ICV_6 $T=188140 252960 1 0 $X=187950 $Y=250000
X883 1 2 891 119 136 ICV_6 $T=188140 312800 1 0 $X=187950 $Y=309840
X884 1 2 920 923 135 ICV_6 $T=201940 296480 0 0 $X=201750 $Y=296240
X885 1 2 977 973 123 ICV_6 $T=230000 269280 0 0 $X=229810 $Y=269040
X886 1 2 978 954 131 ICV_6 $T=230000 291040 0 0 $X=229810 $Y=290800
X887 1 2 1010 973 117 ICV_6 $T=244260 269280 1 0 $X=244070 $Y=266320
X888 1 2 1001 154 131 ICV_6 $T=244260 312800 1 0 $X=244070 $Y=309840
X889 1 2 1039 986 121 ICV_6 $T=258060 263840 0 0 $X=257870 $Y=263600
X890 1 2 1037 1012 122 ICV_6 $T=258060 274720 0 0 $X=257870 $Y=274480
X891 1 2 1034 164 122 ICV_6 $T=258060 307360 0 0 $X=257870 $Y=307120
X892 1 2 1068 168 136 ICV_6 $T=272320 312800 1 0 $X=272130 $Y=309840
X893 1 2 1090 1086 121 ICV_6 $T=286120 291040 0 0 $X=285930 $Y=290800
X894 1 2 1130 1105 122 ICV_6 $T=300380 280160 1 0 $X=300190 $Y=277200
X895 1 2 1192 1184 123 ICV_6 $T=342240 252960 0 0 $X=342050 $Y=252720
X896 1 2 1190 1184 135 ICV_6 $T=342240 263840 0 0 $X=342050 $Y=263600
X897 1 2 245 248 178 ICV_6 $T=356500 274720 1 0 $X=356310 $Y=271760
X898 1 2 1224 1199 131 ICV_6 $T=356500 291040 1 0 $X=356310 $Y=288080
X899 1 2 271 270 202 ICV_6 $T=384560 312800 1 0 $X=384370 $Y=309840
X900 1 2 1309 280 188 ICV_6 $T=398360 307360 0 0 $X=398170 $Y=307120
X901 1 2 1336 1312 262 ICV_6 $T=412620 274720 1 0 $X=412430 $Y=271760
X902 1 2 1365 1348 201 ICV_6 $T=426420 269280 0 0 $X=426230 $Y=269040
X903 1 2 1453 319 262 ICV_6 $T=468740 252960 1 0 $X=468550 $Y=250000
X904 1 2 1486 1449 186 ICV_6 $T=482540 291040 0 0 $X=482350 $Y=290800
X905 1 2 1509 1504 202 ICV_6 $T=496800 296480 1 0 $X=496610 $Y=293520
X906 1 2 1510 355 178 ICV_6 $T=496800 312800 1 0 $X=496610 $Y=309840
X907 1 2 1542 369 348 ICV_6 $T=510600 247520 0 0 $X=510410 $Y=247280
X908 1 2 1540 1504 188 ICV_6 $T=510600 307360 0 0 $X=510410 $Y=307120
X909 1 2 1569 369 303 ICV_6 $T=524860 247520 1 0 $X=524670 $Y=244560
X910 1 2 1591 1576 372 ICV_6 $T=538660 263840 0 0 $X=538470 $Y=263600
X911 1 2 1623 411 370 ICV_6 $T=552920 307360 1 0 $X=552730 $Y=304400
X912 1 2 1703 1681 263 ICV_6 $T=594780 269280 0 0 $X=594590 $Y=269040
X913 1 2 1707 1701 376 ICV_6 $T=594780 307360 0 0 $X=594590 $Y=307120
X914 1 2 1876 1859 341 ICV_6 $T=678960 247520 0 0 $X=678770 $Y=247280
X915 1 2 1908 1904 341 ICV_6 $T=693220 285600 1 0 $X=693030 $Y=282640
X916 1 2 1903 1904 337 ICV_6 $T=693220 291040 1 0 $X=693030 $Y=288080
X917 1 2 1922 453 328 ICV_6 $T=707020 247520 0 0 $X=706830 $Y=247280
X918 1 2 1959 463 348 ICV_6 $T=721280 252960 1 0 $X=721090 $Y=250000
X919 1 2 1975 1950 328 ICV_6 $T=735080 285600 0 0 $X=734890 $Y=285360
X920 1 2 1981 1950 337 ICV_6 $T=735080 291040 0 0 $X=734890 $Y=290800
X1086 1 2 ICV_10 $T=17020 285600 1 0 $X=16830 $Y=282640
X1087 1 2 ICV_10 $T=17020 296480 1 0 $X=16830 $Y=293520
X1088 1 2 ICV_10 $T=30820 258400 0 0 $X=30630 $Y=258160
X1089 1 2 ICV_10 $T=45080 258400 1 0 $X=44890 $Y=255440
X1090 1 2 ICV_10 $T=45080 285600 1 0 $X=44890 $Y=282640
X1091 1 2 ICV_10 $T=101200 247520 1 0 $X=101010 $Y=244560
X1092 1 2 ICV_10 $T=241500 274720 1 0 $X=241310 $Y=271760
X1093 1 2 ICV_10 $T=241500 291040 1 0 $X=241310 $Y=288080
X1094 1 2 ICV_10 $T=255300 252960 0 0 $X=255110 $Y=252720
X1095 1 2 ICV_10 $T=269560 269280 1 0 $X=269370 $Y=266320
X1096 1 2 ICV_10 $T=325680 274720 1 0 $X=325490 $Y=271760
X1097 1 2 ICV_10 $T=339480 269280 0 0 $X=339290 $Y=269040
X1098 1 2 ICV_10 $T=339480 296480 0 0 $X=339290 $Y=296240
X1099 1 2 ICV_10 $T=353740 312800 1 0 $X=353550 $Y=309840
X1100 1 2 ICV_10 $T=395600 252960 0 0 $X=395410 $Y=252720
X1101 1 2 ICV_10 $T=522100 291040 1 0 $X=521910 $Y=288080
X1102 1 2 ICV_10 $T=535900 269280 0 0 $X=535710 $Y=269040
X1103 1 2 ICV_10 $T=535900 274720 0 0 $X=535710 $Y=274480
X1104 1 2 ICV_10 $T=563960 252960 0 0 $X=563770 $Y=252720
X1105 1 2 ICV_10 $T=563960 269280 0 0 $X=563770 $Y=269040
X1106 1 2 ICV_10 $T=662400 269280 1 0 $X=662210 $Y=266320
X1107 1 2 ICV_10 $T=662400 307360 1 0 $X=662210 $Y=304400
X1108 1 2 ICV_10 $T=718520 285600 1 0 $X=718330 $Y=282640
X1109 1 2 525 10 2 548 1 sky130_fd_sc_hd__dfxtp_1 $T=9660 285600 1 0 $X=9470 $Y=282640
X1110 1 2 628 14 2 626 1 sky130_fd_sc_hd__dfxtp_1 $T=67160 269280 1 0 $X=66970 $Y=266320
X1111 1 2 70 14 2 705 1 sky130_fd_sc_hd__dfxtp_1 $T=87860 312800 1 0 $X=87670 $Y=309840
X1112 1 2 708 26 2 731 1 sky130_fd_sc_hd__dfxtp_1 $T=99820 280160 0 0 $X=99630 $Y=279920
X1113 1 2 707 11 2 734 1 sky130_fd_sc_hd__dfxtp_1 $T=101200 269280 0 0 $X=101010 $Y=269040
X1114 1 2 685 11 2 726 1 sky130_fd_sc_hd__dfxtp_1 $T=104420 296480 0 0 $X=104230 $Y=296240
X1115 1 2 84 25 2 745 1 sky130_fd_sc_hd__dfxtp_1 $T=111780 252960 1 0 $X=111590 $Y=250000
X1116 1 2 738 10 2 756 1 sky130_fd_sc_hd__dfxtp_1 $T=112240 296480 1 0 $X=112050 $Y=293520
X1117 1 2 738 4 2 796 1 sky130_fd_sc_hd__dfxtp_1 $T=135240 301920 0 0 $X=135050 $Y=301680
X1118 1 2 789 26 2 802 1 sky130_fd_sc_hd__dfxtp_1 $T=135700 263840 0 0 $X=135510 $Y=263600
X1119 1 2 761 14 2 800 1 sky130_fd_sc_hd__dfxtp_1 $T=137540 274720 0 0 $X=137350 $Y=274480
X1120 1 2 101 26 2 815 1 sky130_fd_sc_hd__dfxtp_1 $T=143060 307360 1 0 $X=142870 $Y=304400
X1121 1 2 789 11 2 830 1 sky130_fd_sc_hd__dfxtp_1 $T=147200 263840 1 0 $X=147010 $Y=260880
X1122 1 2 854 112 2 869 1 sky130_fd_sc_hd__dfxtp_1 $T=168360 301920 1 0 $X=168170 $Y=298960
X1123 1 2 853 112 2 872 1 sky130_fd_sc_hd__dfxtp_1 $T=168820 285600 1 0 $X=168630 $Y=282640
X1124 1 2 859 111 2 883 1 sky130_fd_sc_hd__dfxtp_1 $T=176180 263840 1 0 $X=175990 $Y=260880
X1125 1 2 109 128 2 890 1 sky130_fd_sc_hd__dfxtp_1 $T=178940 301920 0 0 $X=178750 $Y=301680
X1126 1 2 853 127 2 892 1 sky130_fd_sc_hd__dfxtp_1 $T=179860 280160 1 0 $X=179670 $Y=277200
X1127 1 2 906 112 2 901 1 sky130_fd_sc_hd__dfxtp_1 $T=194580 296480 1 0 $X=194390 $Y=293520
X1128 1 2 153 125 2 1000 1 sky130_fd_sc_hd__dfxtp_1 $T=231840 307360 0 0 $X=231650 $Y=307120
X1129 1 2 987 111 2 1009 1 sky130_fd_sc_hd__dfxtp_1 $T=235980 263840 1 0 $X=235790 $Y=260880
X1130 1 2 987 108 2 1039 1 sky130_fd_sc_hd__dfxtp_1 $T=249780 263840 0 0 $X=249590 $Y=263600
X1131 1 2 1020 128 2 1040 1 sky130_fd_sc_hd__dfxtp_1 $T=250700 269280 0 0 $X=250510 $Y=269040
X1132 1 2 990 128 2 1043 1 sky130_fd_sc_hd__dfxtp_1 $T=252080 285600 1 0 $X=251890 $Y=282640
X1133 1 2 1045 125 2 1061 1 sky130_fd_sc_hd__dfxtp_1 $T=262200 280160 0 0 $X=262010 $Y=279920
X1134 1 2 1020 112 2 1074 1 sky130_fd_sc_hd__dfxtp_1 $T=270480 269280 0 0 $X=270290 $Y=269040
X1135 1 2 1054 108 2 1078 1 sky130_fd_sc_hd__dfxtp_1 $T=275540 258400 0 0 $X=275350 $Y=258160
X1136 1 2 1070 110 2 1113 1 sky130_fd_sc_hd__dfxtp_1 $T=289340 301920 1 0 $X=289150 $Y=298960
X1137 1 2 1096 110 2 1130 1 sky130_fd_sc_hd__dfxtp_1 $T=293940 280160 0 0 $X=293750 $Y=279920
X1138 1 2 1116 128 2 1155 1 sky130_fd_sc_hd__dfxtp_1 $T=308200 307360 1 0 $X=308010 $Y=304400
X1139 1 2 179 112 2 1158 1 sky130_fd_sc_hd__dfxtp_1 $T=309580 312800 1 0 $X=309390 $Y=309840
X1140 1 2 1180 111 2 1188 1 sky130_fd_sc_hd__dfxtp_1 $T=327980 285600 0 0 $X=327790 $Y=285360
X1141 1 2 1182 127 2 1204 1 sky130_fd_sc_hd__dfxtp_1 $T=332120 269280 0 0 $X=331930 $Y=269040
X1142 1 2 177 202 2 211 1 sky130_fd_sc_hd__dfxtp_1 $T=333500 291040 0 0 $X=333310 $Y=290800
X1143 1 2 1182 126 2 1207 1 sky130_fd_sc_hd__dfxtp_1 $T=335340 280160 1 0 $X=335150 $Y=277200
X1144 1 2 220 253 2 1246 1 sky130_fd_sc_hd__dfxtp_1 $T=359720 247520 1 0 $X=359530 $Y=244560
X1145 1 2 1231 213 2 1251 1 sky130_fd_sc_hd__dfxtp_1 $T=359720 307360 0 0 $X=359530 $Y=307120
X1146 1 2 1258 218 2 1280 1 sky130_fd_sc_hd__dfxtp_1 $T=374900 307360 1 0 $X=374710 $Y=304400
X1147 1 2 1258 210 2 1288 1 sky130_fd_sc_hd__dfxtp_1 $T=379500 291040 0 0 $X=379310 $Y=290800
X1148 1 2 1256 251 2 1303 1 sky130_fd_sc_hd__dfxtp_1 $T=391000 258400 1 0 $X=390810 $Y=255440
X1149 1 2 284 224 2 1325 1 sky130_fd_sc_hd__dfxtp_1 $T=400200 247520 0 0 $X=400010 $Y=247280
X1150 1 2 1290 250 2 1336 1 sky130_fd_sc_hd__dfxtp_1 $T=405260 274720 1 0 $X=405070 $Y=271760
X1151 1 2 1322 222 2 1347 1 sky130_fd_sc_hd__dfxtp_1 $T=409860 301920 0 0 $X=409670 $Y=301680
X1152 1 2 1338 238 2 1365 1 sky130_fd_sc_hd__dfxtp_1 $T=418140 269280 0 0 $X=417950 $Y=269040
X1153 1 2 177 303 2 1332 1 sky130_fd_sc_hd__dfxtp_1 $T=425040 291040 1 0 $X=424850 $Y=288080
X1154 1 2 1380 223 2 1403 1 sky130_fd_sc_hd__dfxtp_1 $T=443440 274720 0 0 $X=443250 $Y=274480
X1155 1 2 1396 227 2 1416 1 sky130_fd_sc_hd__dfxtp_1 $T=443900 263840 0 0 $X=443710 $Y=263600
X1156 1 2 1412 214 2 1425 1 sky130_fd_sc_hd__dfxtp_1 $T=448500 307360 1 0 $X=448310 $Y=304400
X1157 1 2 1396 251 2 1447 1 sky130_fd_sc_hd__dfxtp_1 $T=458620 263840 0 0 $X=458430 $Y=263600
X1158 1 2 1396 224 2 1426 1 sky130_fd_sc_hd__dfxtp_1 $T=459540 263840 1 0 $X=459350 $Y=260880
X1159 1 2 316 238 2 1450 1 sky130_fd_sc_hd__dfxtp_1 $T=460000 258400 1 0 $X=459810 $Y=255440
X1160 1 2 316 224 2 1452 1 sky130_fd_sc_hd__dfxtp_1 $T=460460 247520 1 0 $X=460270 $Y=244560
X1161 1 2 177 328 2 1318 1 sky130_fd_sc_hd__dfxtp_1 $T=465520 285600 0 0 $X=465330 $Y=285360
X1162 1 2 177 337 2 1463 1 sky130_fd_sc_hd__dfxtp_1 $T=474260 291040 0 0 $X=474070 $Y=290800
X1163 1 2 1441 222 2 1481 1 sky130_fd_sc_hd__dfxtp_1 $T=474720 301920 0 0 $X=474530 $Y=301680
X1164 1 2 1441 216 2 1486 1 sky130_fd_sc_hd__dfxtp_1 $T=476100 296480 1 0 $X=475910 $Y=293520
X1165 1 2 336 223 2 1487 1 sky130_fd_sc_hd__dfxtp_1 $T=477020 247520 1 0 $X=476830 $Y=244560
X1166 1 2 1483 251 2 1490 1 sky130_fd_sc_hd__dfxtp_1 $T=482080 269280 1 0 $X=481890 $Y=266320
X1167 1 2 177 341 2 1440 1 sky130_fd_sc_hd__dfxtp_1 $T=482540 291040 1 0 $X=482350 $Y=288080
X1168 1 2 1483 250 2 1516 1 sky130_fd_sc_hd__dfxtp_1 $T=492660 269280 0 0 $X=492470 $Y=269040
X1169 1 2 1521 359 2 1535 1 sky130_fd_sc_hd__dfxtp_1 $T=500940 280160 1 0 $X=500750 $Y=277200
X1170 1 2 1515 368 2 1550 1 sky130_fd_sc_hd__dfxtp_1 $T=509220 263840 1 0 $X=509030 $Y=260880
X1171 1 2 362 363 2 1569 1 sky130_fd_sc_hd__dfxtp_1 $T=517960 247520 0 0 $X=517770 $Y=247280
X1172 1 2 1572 368 2 1586 1 sky130_fd_sc_hd__dfxtp_1 $T=528080 296480 0 0 $X=527890 $Y=296240
X1173 1 2 1574 364 2 1594 1 sky130_fd_sc_hd__dfxtp_1 $T=531300 269280 1 0 $X=531110 $Y=266320
X1174 1 2 1574 358 2 1609 1 sky130_fd_sc_hd__dfxtp_1 $T=540500 269280 1 0 $X=540310 $Y=266320
X1175 1 2 1601 356 2 1622 1 sky130_fd_sc_hd__dfxtp_1 $T=546480 291040 0 0 $X=546290 $Y=290800
X1176 1 2 393 368 2 413 1 sky130_fd_sc_hd__dfxtp_1 $T=560740 247520 1 0 $X=560550 $Y=244560
X1177 1 2 1641 418 2 1682 1 sky130_fd_sc_hd__dfxtp_1 $T=575920 307360 0 0 $X=575730 $Y=307120
X1178 1 2 412 253 2 1678 1 sky130_fd_sc_hd__dfxtp_1 $T=584200 247520 0 0 $X=584010 $Y=247280
X1179 1 2 1659 223 2 1705 1 sky130_fd_sc_hd__dfxtp_1 $T=587880 285600 1 0 $X=587690 $Y=282640
X1180 1 2 1690 390 2 1707 1 sky130_fd_sc_hd__dfxtp_1 $T=589720 312800 1 0 $X=589530 $Y=309840
X1181 1 2 1763 253 2 1760 1 sky130_fd_sc_hd__dfxtp_1 $T=632040 274720 0 0 $X=631850 $Y=274480
X1182 1 2 441 253 2 1794 1 sky130_fd_sc_hd__dfxtp_1 $T=634800 247520 0 0 $X=634610 $Y=247280
X1183 1 2 437 404 2 445 1 sky130_fd_sc_hd__dfxtp_1 $T=643080 307360 0 0 $X=642890 $Y=307120
X1184 1 2 1848 363 2 1879 1 sky130_fd_sc_hd__dfxtp_1 $T=674360 285600 1 0 $X=674170 $Y=282640
X1185 1 2 1873 418 2 1877 1 sky130_fd_sc_hd__dfxtp_1 $T=675280 312800 1 0 $X=675090 $Y=309840
X1186 1 2 1893 363 2 1907 1 sky130_fd_sc_hd__dfxtp_1 $T=686780 274720 0 0 $X=686590 $Y=274480
X1187 1 2 1886 359 2 1908 1 sky130_fd_sc_hd__dfxtp_1 $T=686780 280160 0 0 $X=686590 $Y=279920
X1188 1 2 1873 388 2 1911 1 sky130_fd_sc_hd__dfxtp_1 $T=695060 301920 0 0 $X=694870 $Y=301680
X1189 1 2 1893 358 2 1931 1 sky130_fd_sc_hd__dfxtp_1 $T=701960 274720 1 0 $X=701770 $Y=271760
X1190 1 2 456 385 2 1934 1 sky130_fd_sc_hd__dfxtp_1 $T=701960 312800 1 0 $X=701770 $Y=309840
X1191 1 2 450 367 2 1929 1 sky130_fd_sc_hd__dfxtp_1 $T=704260 247520 1 0 $X=704070 $Y=244560
X1192 1 2 1946 364 2 1967 1 sky130_fd_sc_hd__dfxtp_1 $T=716220 274720 0 0 $X=716030 $Y=274480
X1193 1 2 1951 359 2 465 1 sky130_fd_sc_hd__dfxtp_1 $T=718980 252960 0 0 $X=718790 $Y=252720
X1194 1 2 1943 364 2 1970 1 sky130_fd_sc_hd__dfxtp_1 $T=719440 280160 0 0 $X=719250 $Y=279920
X1195 1 2 1944 364 2 1968 1 sky130_fd_sc_hd__dfxtp_1 $T=719900 291040 0 0 $X=719710 $Y=290800
X1196 1 2 1951 368 2 468 1 sky130_fd_sc_hd__dfxtp_1 $T=727720 252960 0 0 $X=727530 $Y=252720
X1197 1 2 557 542 33 522 24 557 ICV_13 $T=20240 269280 1 0 $X=20050 $Y=266320
X1198 1 2 27 29 17 524 14 558 ICV_13 $T=20240 307360 1 0 $X=20050 $Y=304400
X1199 1 2 559 29 30 21 25 559 ICV_13 $T=20240 312800 1 0 $X=20050 $Y=309840
X1200 1 2 560 527 34 523 26 560 ICV_13 $T=20700 247520 0 0 $X=20510 $Y=247280
X1201 1 2 562 527 33 523 24 562 ICV_13 $T=21160 252960 0 0 $X=20970 $Y=252720
X1202 1 2 565 545 30 525 25 565 ICV_13 $T=21160 274720 0 0 $X=20970 $Y=274480
X1203 1 2 570 542 19 522 14 570 ICV_13 $T=21620 269280 0 0 $X=21430 $Y=269040
X1204 1 2 586 45 33 32 24 586 ICV_13 $T=33120 252960 1 0 $X=32930 $Y=250000
X1205 1 2 592 578 30 579 25 592 ICV_13 $T=34040 258400 0 0 $X=33850 $Y=258160
X1206 1 2 596 29 33 21 24 596 ICV_13 $T=34040 307360 0 0 $X=33850 $Y=307120
X1207 1 2 614 47 17 42 4 614 ICV_13 $T=45540 307360 0 0 $X=45350 $Y=307120
X1208 1 2 615 602 17 582 4 615 ICV_13 $T=46000 274720 0 0 $X=45810 $Y=274480
X1209 1 2 621 578 17 579 4 621 ICV_13 $T=48300 263840 1 0 $X=48110 $Y=260880
X1210 1 2 622 602 18 582 11 622 ICV_13 $T=48300 280160 1 0 $X=48110 $Y=277200
X1211 1 2 613 585 33 581 14 623 ICV_13 $T=48300 291040 1 0 $X=48110 $Y=288080
X1212 1 2 624 578 33 579 24 624 ICV_13 $T=49220 258400 0 0 $X=49030 $Y=258160
X1213 1 2 629 47 30 42 5 635 ICV_13 $T=54280 307360 1 0 $X=54090 $Y=304400
X1214 1 2 638 47 34 42 26 638 ICV_13 $T=55200 312800 1 0 $X=55010 $Y=309840
X1215 1 2 640 642 34 618 26 640 ICV_13 $T=55660 296480 1 0 $X=55470 $Y=293520
X1216 1 2 645 627 17 617 14 646 ICV_13 $T=62100 274720 1 0 $X=61910 $Y=271760
X1217 1 2 652 641 30 617 25 652 ICV_13 $T=63020 280160 0 0 $X=62830 $Y=279920
X1218 1 2 662 56 13 619 10 662 ICV_13 $T=68540 252960 0 0 $X=68350 $Y=252720
X1219 1 2 650 627 30 628 10 625 ICV_13 $T=69460 263840 0 0 $X=69270 $Y=263600
X1220 1 2 651 56 19 619 5 666 ICV_13 $T=69920 247520 0 0 $X=69730 $Y=247280
X1221 1 2 677 676 17 664 5 672 ICV_13 $T=75900 274720 0 0 $X=75710 $Y=274480
X1222 1 2 672 676 16 665 14 678 ICV_13 $T=76360 280160 1 0 $X=76170 $Y=277200
X1223 1 2 679 684 18 665 11 679 ICV_13 $T=76360 285600 1 0 $X=76170 $Y=282640
X1224 1 2 683 66 30 62 25 683 ICV_13 $T=76360 312800 1 0 $X=76170 $Y=309840
X1225 1 2 688 690 33 670 14 687 ICV_13 $T=81420 263840 1 0 $X=81230 $Y=260880
X1226 1 2 710 78 19 71 14 710 ICV_13 $T=90160 247520 0 0 $X=89970 $Y=247280
X1227 1 2 712 684 33 665 26 703 ICV_13 $T=90160 285600 0 0 $X=89970 $Y=285360
X1228 1 2 715 690 13 670 10 715 ICV_13 $T=91540 258400 1 0 $X=91350 $Y=255440
X1229 1 2 719 690 17 670 26 720 ICV_13 $T=94760 252960 0 0 $X=94570 $Y=252720
X1230 1 2 721 693 16 685 5 721 ICV_13 $T=96140 301920 0 0 $X=95950 $Y=301680
X1231 1 2 739 730 30 707 4 736 ICV_13 $T=103040 258400 0 0 $X=102850 $Y=258160
X1232 1 2 737 730 19 707 14 737 ICV_13 $T=103500 274720 0 0 $X=103310 $Y=274480
X1233 1 2 749 77 17 70 4 749 ICV_13 $T=108560 312800 1 0 $X=108370 $Y=309840
X1234 1 2 748 740 18 708 14 747 ICV_13 $T=109020 285600 1 0 $X=108830 $Y=282640
X1235 1 2 754 757 34 738 26 754 ICV_13 $T=110860 307360 1 0 $X=110670 $Y=304400
X1236 1 2 767 771 13 84 14 95 ICV_13 $T=118220 247520 0 0 $X=118030 $Y=247280
X1237 1 2 765 772 18 755 11 765 ICV_13 $T=118220 285600 0 0 $X=118030 $Y=285360
X1238 1 2 769 772 30 755 25 769 ICV_13 $T=119140 291040 0 0 $X=118950 $Y=290800
X1239 1 2 773 772 16 755 5 773 ICV_13 $T=119600 296480 1 0 $X=119410 $Y=293520
X1240 1 2 775 718 30 744 25 775 ICV_13 $T=120980 269280 0 0 $X=120790 $Y=269040
X1241 1 2 791 771 34 764 26 791 ICV_13 $T=129720 247520 0 0 $X=129530 $Y=247280
X1242 1 2 801 772 34 755 26 801 ICV_13 $T=135240 291040 1 0 $X=135050 $Y=288080
X1243 1 2 818 89 17 101 4 818 ICV_13 $T=143520 312800 1 0 $X=143330 $Y=309840
X1244 1 2 823 822 34 809 26 823 ICV_13 $T=145820 274720 1 0 $X=145630 $Y=271760
X1245 1 2 829 824 30 810 25 829 ICV_13 $T=146740 291040 1 0 $X=146550 $Y=288080
X1246 1 2 850 835 16 813 5 850 ICV_13 $T=157780 247520 0 0 $X=157590 $Y=247280
X1247 1 2 857 835 33 813 24 857 ICV_13 $T=160540 258400 1 0 $X=160350 $Y=255440
X1248 1 2 867 873 117 854 111 867 ICV_13 $T=167900 291040 1 0 $X=167710 $Y=288080
X1249 1 2 876 862 121 861 112 878 ICV_13 $T=174340 263840 0 0 $X=174150 $Y=263600
X1250 1 2 882 119 117 109 111 882 ICV_13 $T=175720 307360 1 0 $X=175530 $Y=304400
X1251 1 2 130 119 134 109 125 887 ICV_13 $T=178480 307360 0 0 $X=178290 $Y=307120
X1252 1 2 889 873 134 854 127 889 ICV_13 $T=178940 296480 0 0 $X=178750 $Y=296240
X1253 1 2 888 874 136 853 125 893 ICV_13 $T=179860 280160 0 0 $X=179670 $Y=279920
X1254 1 2 894 873 136 854 126 894 ICV_13 $T=179860 291040 0 0 $X=179670 $Y=290800
X1255 1 2 909 863 136 859 126 909 ICV_13 $T=188600 263840 1 0 $X=188410 $Y=260880
X1256 1 2 910 862 136 861 126 910 ICV_13 $T=188600 269280 1 0 $X=188410 $Y=266320
X1257 1 2 916 144 123 906 108 142 ICV_13 $T=195040 301920 1 0 $X=194850 $Y=298960
X1258 1 2 926 145 135 140 108 143 ICV_13 $T=195960 247520 1 0 $X=195770 $Y=244560
X1259 1 2 930 146 117 141 128 928 ICV_13 $T=202400 252960 0 0 $X=202210 $Y=252720
X1260 1 2 935 144 122 137 111 941 ICV_13 $T=203320 307360 0 0 $X=203130 $Y=307120
X1261 1 2 942 933 135 927 125 942 ICV_13 $T=203780 263840 1 0 $X=203590 $Y=260880
X1262 1 2 957 139 136 906 111 955 ICV_13 $T=214360 296480 0 0 $X=214170 $Y=296240
X1263 1 2 960 146 123 141 112 960 ICV_13 $T=216660 252960 1 0 $X=216470 $Y=250000
X1264 1 2 962 954 135 906 126 957 ICV_13 $T=216660 296480 1 0 $X=216470 $Y=293520
X1265 1 2 967 921 135 919 125 967 ICV_13 $T=217580 274720 0 0 $X=217390 $Y=274480
X1266 1 2 982 973 134 956 127 982 ICV_13 $T=223100 269280 1 0 $X=222910 $Y=266320
X1267 1 2 992 954 134 950 127 992 ICV_13 $T=230000 291040 1 0 $X=229810 $Y=288080
X1268 1 2 994 973 121 956 108 994 ICV_13 $T=230460 274720 0 0 $X=230270 $Y=274480
X1269 1 2 995 954 117 950 108 996 ICV_13 $T=230460 285600 0 0 $X=230270 $Y=285360
X1270 1 2 997 975 121 979 108 997 ICV_13 $T=230460 296480 0 0 $X=230270 $Y=296240
X1271 1 2 1000 154 135 153 128 1001 ICV_13 $T=231840 312800 1 0 $X=231650 $Y=309840
X1272 1 2 1003 155 131 987 110 1002 ICV_13 $T=232760 258400 1 0 $X=232570 $Y=255440
X1273 1 2 1002 986 122 987 112 1004 ICV_13 $T=233220 258400 0 0 $X=233030 $Y=258160
X1274 1 2 1024 155 134 983 127 1024 ICV_13 $T=244720 247520 1 0 $X=244530 $Y=244560
X1275 1 2 1025 155 122 983 110 1025 ICV_13 $T=244720 252960 1 0 $X=244530 $Y=250000
X1276 1 2 1023 1012 135 979 125 991 ICV_13 $T=244720 291040 1 0 $X=244530 $Y=288080
X1277 1 2 1005 973 131 990 112 1030 ICV_13 $T=249320 274720 1 0 $X=249130 $Y=271760
X1278 1 2 1042 986 134 987 127 1042 ICV_13 $T=252080 263840 1 0 $X=251890 $Y=260880
X1279 1 2 1052 161 135 163 125 1052 ICV_13 $T=258520 247520 0 0 $X=258330 $Y=247280
X1280 1 2 1056 1032 121 1022 128 1051 ICV_13 $T=258520 296480 0 0 $X=258330 $Y=296240
X1281 1 2 1063 1032 122 1022 108 1056 ICV_13 $T=260820 296480 1 0 $X=260630 $Y=293520
X1282 1 2 1077 161 123 163 111 169 ICV_13 $T=270020 247520 0 0 $X=269830 $Y=247280
X1283 1 2 1064 1059 123 1020 111 1075 ICV_13 $T=270480 274720 0 0 $X=270290 $Y=274480
X1284 1 2 1079 1059 122 1045 128 1076 ICV_13 $T=270480 285600 0 0 $X=270290 $Y=285360
X1285 1 2 1082 1027 136 1020 126 1082 ICV_13 $T=272780 269280 1 0 $X=272590 $Y=266320
X1286 1 2 1083 1027 121 1020 108 1083 ICV_13 $T=272780 274720 1 0 $X=272590 $Y=271760
X1287 1 2 1062 1059 134 1045 110 1079 ICV_13 $T=272780 285600 1 0 $X=272590 $Y=282640
X1288 1 2 1088 1086 117 1070 111 1088 ICV_13 $T=274620 291040 0 0 $X=274430 $Y=290800
X1289 1 2 1093 168 117 166 111 1093 ICV_13 $T=276920 312800 1 0 $X=276730 $Y=309840
X1290 1 2 1107 1105 117 1096 111 1107 ICV_13 $T=284740 291040 1 0 $X=284550 $Y=288080
X1291 1 2 1110 1053 131 1054 128 1110 ICV_13 $T=286580 258400 0 0 $X=286390 $Y=258160
X1292 1 2 1099 1053 136 1054 125 1100 ICV_13 $T=287500 263840 1 0 $X=287310 $Y=260880
X1293 1 2 1115 1104 122 1097 110 1115 ICV_13 $T=287500 269280 0 0 $X=287310 $Y=269040
X1294 1 2 1122 159 136 170 126 1122 ICV_13 $T=290260 252960 0 0 $X=290070 $Y=252720
X1295 1 2 1133 1124 123 1116 112 1133 ICV_13 $T=294860 301920 0 0 $X=294670 $Y=301680
X1296 1 2 1144 1104 121 1097 108 1144 ICV_13 $T=300840 269280 1 0 $X=300650 $Y=266320
X1297 1 2 1128 1105 123 1096 125 1134 ICV_13 $T=300840 285600 0 0 $X=300650 $Y=285360
X1298 1 2 1145 1105 121 1096 108 1145 ICV_13 $T=301300 280160 0 0 $X=301110 $Y=279920
X1299 1 2 1148 1146 121 1129 125 1147 ICV_13 $T=302680 258400 0 0 $X=302490 $Y=258160
X1300 1 2 1152 1124 136 1116 127 1151 ICV_13 $T=306820 301920 1 0 $X=306630 $Y=298960
X1301 1 2 1163 1146 122 1129 110 1163 ICV_13 $T=313260 258400 1 0 $X=313070 $Y=255440
X1302 1 2 1172 1123 136 1142 108 1170 ICV_13 $T=318320 274720 0 0 $X=318130 $Y=274480
X1303 1 2 1175 1166 122 1159 110 1175 ICV_13 $T=318320 301920 0 0 $X=318130 $Y=301680
X1304 1 2 1179 184 122 176 110 1179 ICV_13 $T=321080 247520 0 0 $X=320890 $Y=247280
X1305 1 2 1185 1166 123 1159 112 1185 ICV_13 $T=324300 307360 0 0 $X=324110 $Y=307120
X1306 1 2 1195 1166 121 1159 108 1195 ICV_13 $T=328900 301920 1 0 $X=328710 $Y=298960
X1307 1 2 1201 1183 131 1180 125 1197 ICV_13 $T=330280 280160 0 0 $X=330090 $Y=279920
X1308 1 2 1216 1203 186 1206 216 1216 ICV_13 $T=342700 291040 0 0 $X=342510 $Y=290800
X1309 1 2 1217 1203 192 1206 217 1217 ICV_13 $T=342700 296480 0 0 $X=342510 $Y=296240
X1310 1 2 1189 1166 131 1206 219 1220 ICV_13 $T=343620 296480 1 0 $X=343430 $Y=293520
X1311 1 2 1218 1203 188 1206 222 1221 ICV_13 $T=345000 301920 0 0 $X=344810 $Y=301680
X1312 1 2 1225 1199 136 1180 126 1225 ICV_13 $T=347760 285600 0 0 $X=347570 $Y=285360
X1313 1 2 1229 1199 134 1180 108 1233 ICV_13 $T=357420 280160 0 0 $X=357230 $Y=279920
X1314 1 2 1239 247 262 220 250 1239 ICV_13 $T=357880 252960 0 0 $X=357690 $Y=252720
X1315 1 2 1263 1240 252 1230 227 1263 ICV_13 $T=367540 269280 1 0 $X=367350 $Y=266320
X1316 1 2 1259 1252 260 1247 251 1264 ICV_13 $T=368000 274720 1 0 $X=367810 $Y=271760
X1317 1 2 1270 1273 201 1256 238 1270 ICV_13 $T=372140 252960 1 0 $X=371950 $Y=250000
X1318 1 2 1281 1253 180 1258 214 1281 ICV_13 $T=375360 301920 0 0 $X=375170 $Y=301680
X1319 1 2 1282 1273 233 1256 224 1282 ICV_13 $T=376280 247520 0 0 $X=376090 $Y=247280
X1320 1 2 1294 1273 260 1256 223 1294 ICV_13 $T=384100 252960 0 0 $X=383910 $Y=252720
X1321 1 2 1296 1277 229 1274 253 1296 ICV_13 $T=385020 263840 1 0 $X=384830 $Y=260880
X1322 1 2 1302 280 202 275 219 1302 ICV_13 $T=389160 312800 1 0 $X=388970 $Y=309840
X1323 1 2 1305 1299 192 1292 222 1317 ICV_13 $T=395140 301920 1 0 $X=394950 $Y=298960
X1324 1 2 1306 1312 257 1290 238 1329 ICV_13 $T=401580 274720 0 0 $X=401390 $Y=274480
X1325 1 2 1334 280 186 275 216 1334 ICV_13 $T=402960 307360 0 0 $X=402770 $Y=307120
X1326 1 2 1279 1253 185 1322 218 1352 ICV_13 $T=413080 301920 1 0 $X=412890 $Y=298960
X1327 1 2 1339 1343 262 1321 223 1356 ICV_13 $T=414460 263840 0 0 $X=414270 $Y=263600
X1328 1 2 1355 1333 186 1322 219 1357 ICV_13 $T=414920 291040 0 0 $X=414730 $Y=290800
X1329 1 2 1360 302 185 298 210 1363 ICV_13 $T=416760 307360 1 0 $X=416570 $Y=304400
X1330 1 2 1372 1348 262 1338 250 1372 ICV_13 $T=421360 274720 1 0 $X=421170 $Y=271760
X1331 1 2 1381 1343 263 1321 251 1381 ICV_13 $T=426880 263840 1 0 $X=426690 $Y=260880
X1332 1 2 1385 1343 229 1321 253 1385 ICV_13 $T=427800 258400 0 0 $X=427610 $Y=258160
X1333 1 2 1392 302 202 298 219 1392 ICV_13 $T=431480 307360 0 0 $X=431290 $Y=307120
X1334 1 2 1399 1370 252 1349 227 1399 ICV_13 $T=435160 252960 0 0 $X=434970 $Y=252720
X1335 1 2 1401 1387 180 1369 214 1401 ICV_13 $T=435160 296480 0 0 $X=434970 $Y=296240
X1336 1 2 1402 1387 188 1369 218 1402 ICV_13 $T=435160 301920 0 0 $X=434970 $Y=301680
X1337 1 2 1408 1406 252 1380 227 1408 ICV_13 $T=436540 285600 0 0 $X=436350 $Y=285360
X1338 1 2 1410 1406 263 1380 251 1410 ICV_13 $T=437460 269280 0 0 $X=437270 $Y=269040
X1339 1 2 1422 1420 192 1412 222 1430 ICV_13 $T=449420 301920 1 0 $X=449230 $Y=298960
X1340 1 2 1442 1437 262 1418 250 1442 ICV_13 $T=454940 269280 0 0 $X=454750 $Y=269040
X1341 1 2 1432 1437 252 1418 224 1436 ICV_13 $T=454940 280160 0 0 $X=454750 $Y=279920
X1342 1 2 1445 318 192 314 217 1445 ICV_13 $T=454940 312800 1 0 $X=454750 $Y=309840
X1343 1 2 1450 319 201 1396 250 1424 ICV_13 $T=459080 258400 0 0 $X=458890 $Y=258160
X1344 1 2 1444 1420 178 1441 214 1457 ICV_13 $T=462300 296480 0 0 $X=462110 $Y=296240
X1345 1 2 1452 319 233 316 223 332 ICV_13 $T=462760 247520 0 0 $X=462570 $Y=247280
X1346 1 2 1466 1467 229 1454 253 1466 ICV_13 $T=469200 280160 1 0 $X=469010 $Y=277200
X1347 1 2 1471 1467 260 1454 223 1471 ICV_13 $T=470120 274720 0 0 $X=469930 $Y=274480
X1348 1 2 1474 1467 263 1454 251 1474 ICV_13 $T=471040 269280 0 0 $X=470850 $Y=269040
X1349 1 2 1485 1449 188 1441 218 1485 ICV_13 $T=475640 301920 1 0 $X=475450 $Y=298960
X1350 1 2 1498 1470 252 1459 227 1498 ICV_13 $T=484380 252960 0 0 $X=484190 $Y=252720
X1351 1 2 1507 1504 192 1491 217 1507 ICV_13 $T=487140 301920 0 0 $X=486950 $Y=301680
X1352 1 2 1511 1504 185 1491 222 1511 ICV_13 $T=488980 296480 0 0 $X=488790 $Y=296240
X1353 1 2 1512 355 202 347 219 1512 ICV_13 $T=488980 307360 0 0 $X=488790 $Y=307120
X1354 1 2 1520 1484 260 1483 223 1520 ICV_13 $T=494040 274720 0 0 $X=493850 $Y=274480
X1355 1 2 1527 1532 328 1514 359 1531 ICV_13 $T=497720 285600 0 0 $X=497530 $Y=285360
X1356 1 2 1533 1534 341 1515 359 1533 ICV_13 $T=498640 263840 0 0 $X=498450 $Y=263600
X1357 1 2 1538 1504 199 177 361 365 ICV_13 $T=501400 296480 1 0 $X=501210 $Y=293520
X1358 1 2 1537 355 199 347 222 1539 ICV_13 $T=501400 312800 1 0 $X=501210 $Y=309840
X1359 1 2 1541 369 341 362 359 1541 ICV_13 $T=503240 247520 1 0 $X=503050 $Y=244560
X1360 1 2 1551 1519 372 1513 364 1551 ICV_13 $T=510600 252960 1 0 $X=510410 $Y=250000
X1361 1 2 1556 1532 382 1514 368 1556 ICV_13 $T=511980 291040 0 0 $X=511790 $Y=290800
X1362 1 2 1553 1519 306 1513 368 1557 ICV_13 $T=512440 258400 1 0 $X=512250 $Y=255440
X1363 1 2 1558 1547 303 1521 363 1558 ICV_13 $T=513360 274720 1 0 $X=513170 $Y=271760
X1364 1 2 1549 1547 306 1521 368 1559 ICV_13 $T=513820 280160 0 0 $X=513630 $Y=279920
X1365 1 2 1561 1547 337 1521 356 1561 ICV_13 $T=516580 274720 0 0 $X=516390 $Y=274480
X1366 1 2 1575 394 391 379 385 1575 ICV_13 $T=523480 307360 0 0 $X=523290 $Y=307120
X1367 1 2 1577 1583 341 1572 356 1578 ICV_13 $T=525320 291040 1 0 $X=525130 $Y=288080
X1368 1 2 1580 1576 341 1570 359 1580 ICV_13 $T=525780 252960 0 0 $X=525590 $Y=252720
X1369 1 2 1584 1576 382 1570 368 1584 ICV_13 $T=528080 258400 1 0 $X=527890 $Y=255440
X1370 1 2 1592 403 341 1570 367 1593 ICV_13 $T=531300 252960 1 0 $X=531110 $Y=250000
X1371 1 2 1606 1576 337 1570 356 1606 ICV_13 $T=539580 263840 1 0 $X=539390 $Y=260880
X1372 1 2 1612 1589 348 1574 357 1612 ICV_13 $T=540960 280160 1 0 $X=540770 $Y=277200
X1373 1 2 1614 411 389 379 407 1599 ICV_13 $T=541420 307360 1 0 $X=541230 $Y=304400
X1374 1 2 1624 1620 303 1601 363 1624 ICV_13 $T=548320 280160 0 0 $X=548130 $Y=279920
X1375 1 2 1629 1615 348 1617 364 1613 ICV_13 $T=552000 263840 0 0 $X=551810 $Y=263600
X1376 1 2 1632 403 348 393 364 1631 ICV_13 $T=552920 247520 0 0 $X=552730 $Y=247280
X1377 1 2 1638 1620 348 1601 357 1638 ICV_13 $T=553840 291040 0 0 $X=553650 $Y=290800
X1378 1 2 1660 1635 306 1618 367 1660 ICV_13 $T=567180 252960 0 0 $X=566990 $Y=252720
X1379 1 2 1646 1615 328 1617 359 1662 ICV_13 $T=567180 263840 0 0 $X=566990 $Y=263600
X1380 1 2 1663 1650 328 1630 358 1663 ICV_13 $T=567180 285600 0 0 $X=566990 $Y=285360
X1381 1 2 1664 1650 382 1630 364 1665 ICV_13 $T=567180 296480 0 0 $X=566990 $Y=296240
X1382 1 2 417 415 233 412 232 416 ICV_13 $T=568100 247520 1 0 $X=567910 $Y=244560
X1383 1 2 1669 1635 382 1618 368 1669 ICV_13 $T=569020 263840 1 0 $X=568830 $Y=260880
X1384 1 2 1691 1688 262 1672 238 1689 ICV_13 $T=580520 258400 0 0 $X=580330 $Y=258160
X1385 1 2 1693 1685 382 1677 368 1693 ICV_13 $T=581440 296480 1 0 $X=581250 $Y=293520
X1386 1 2 1697 1656 391 1641 385 1697 ICV_13 $T=583280 307360 0 0 $X=583090 $Y=307120
X1387 1 2 1706 1701 375 1690 407 1706 ICV_13 $T=588340 307360 1 0 $X=588150 $Y=304400
X1388 1 2 426 423 260 424 232 1704 ICV_13 $T=595240 247520 0 0 $X=595050 $Y=247280
X1389 1 2 1716 1685 303 1677 363 1716 ICV_13 $T=595240 285600 1 0 $X=595050 $Y=282640
X1390 1 2 1717 1685 337 1677 356 1717 ICV_13 $T=595240 291040 0 0 $X=595050 $Y=290800
X1391 1 2 1720 1701 370 1690 399 1720 ICV_13 $T=597080 301920 1 0 $X=596890 $Y=298960
X1392 1 2 1724 1723 229 1708 253 1724 ICV_13 $T=597540 280160 1 0 $X=597350 $Y=277200
X1393 1 2 1732 1701 373 1690 418 1732 ICV_13 $T=599380 307360 0 0 $X=599190 $Y=307120
X1394 1 2 1752 1723 262 1708 250 1752 ICV_13 $T=610420 269280 0 0 $X=610230 $Y=269040
X1395 1 2 1755 1730 201 1714 238 1755 ICV_13 $T=611340 263840 0 0 $X=611150 $Y=263600
X1396 1 2 1765 1730 252 1714 227 1765 ICV_13 $T=617320 263840 1 0 $X=617130 $Y=260880
X1397 1 2 1768 1739 328 1734 363 1767 ICV_13 $T=619620 291040 1 0 $X=619430 $Y=288080
X1398 1 2 1769 1747 373 1738 418 1769 ICV_13 $T=621000 312800 1 0 $X=620810 $Y=309840
X1399 1 2 1773 1747 375 1738 407 1773 ICV_13 $T=622380 307360 1 0 $X=622190 $Y=304400
X1400 1 2 1775 1730 233 1714 224 1775 ICV_13 $T=623300 258400 0 0 $X=623110 $Y=258160
X1401 1 2 1778 1747 361 1738 388 1778 ICV_13 $T=623300 301920 0 0 $X=623110 $Y=301680
X1402 1 2 1779 435 252 1735 227 1779 ICV_13 $T=623760 247520 1 0 $X=623570 $Y=244560
X1403 1 2 1780 1761 263 1763 251 1780 ICV_13 $T=623760 274720 1 0 $X=623570 $Y=271760
X1404 1 2 1800 444 233 441 224 1800 ICV_13 $T=637560 247520 1 0 $X=637370 $Y=244560
X1405 1 2 1801 1802 233 1788 224 1801 ICV_13 $T=637560 263840 1 0 $X=637370 $Y=260880
X1406 1 2 1805 1804 372 1789 364 1805 ICV_13 $T=637560 296480 1 0 $X=637370 $Y=293520
X1407 1 2 1797 440 370 437 388 1798 ICV_13 $T=637560 312800 1 0 $X=637370 $Y=309840
X1408 1 2 1803 1804 306 1793 224 1817 ICV_13 $T=640320 285600 1 0 $X=640130 $Y=282640
X1409 1 2 1825 1813 262 1793 250 1825 ICV_13 $T=650440 274720 1 0 $X=650250 $Y=271760
X1410 1 2 1826 1802 260 1788 223 1826 ICV_13 $T=650900 269280 1 0 $X=650710 $Y=266320
X1411 1 2 1830 1802 201 1788 238 1830 ICV_13 $T=651360 258400 0 0 $X=651170 $Y=258160
X1412 1 2 1822 1802 262 1788 232 1831 ICV_13 $T=651360 263840 0 0 $X=651170 $Y=263600
X1413 1 2 1849 1812 201 1791 238 1849 ICV_13 $T=658720 247520 0 0 $X=658530 $Y=247280
X1414 1 2 1869 1853 328 1847 363 1870 ICV_13 $T=667920 263840 1 0 $X=667730 $Y=260880
X1415 1 2 1890 1859 306 1846 367 1890 ICV_13 $T=679880 247520 1 0 $X=679690 $Y=244560
X1416 1 2 1898 1866 341 1848 359 1898 ICV_13 $T=681720 285600 1 0 $X=681530 $Y=282640
X1417 1 2 1909 1875 391 1873 385 1909 ICV_13 $T=686780 307360 0 0 $X=686590 $Y=307120
X1418 1 2 1919 1910 372 1893 364 1919 ICV_13 $T=694140 274720 0 0 $X=693950 $Y=274480
X1419 1 2 1945 1916 341 1900 359 1945 ICV_13 $T=707480 252960 0 0 $X=707290 $Y=252720
X1420 1 2 1947 1910 382 1893 356 1930 ICV_13 $T=709320 274720 1 0 $X=709130 $Y=271760
X1421 1 2 1936 1910 306 1893 368 1947 ICV_13 $T=709780 269280 1 0 $X=709590 $Y=266320
X1422 1 2 1960 1950 306 1944 367 1960 ICV_13 $T=714380 285600 0 0 $X=714190 $Y=285360
X1423 1 2 1948 464 376 456 407 1961 ICV_13 $T=714380 307360 0 0 $X=714190 $Y=307120
X1424 1 2 1966 1955 341 1946 359 1966 ICV_13 $T=716220 263840 0 0 $X=716030 $Y=263600
X1425 1 2 1976 1950 303 1944 363 1976 ICV_13 $T=726800 291040 1 0 $X=726610 $Y=288080
X1426 1 2 1977 1950 382 1944 368 1977 ICV_13 $T=726800 296480 1 0 $X=726610 $Y=293520
X1427 1 2 525 5 539 539 545 16 ICV_14 $T=6900 280160 1 0 $X=6710 $Y=277200
X1428 1 2 524 10 540 540 543 13 ICV_14 $T=6900 307360 1 0 $X=6710 $Y=304400
X1429 1 2 525 14 566 566 545 19 ICV_14 $T=20240 280160 1 0 $X=20050 $Y=277200
X1430 1 2 524 25 569 569 543 30 ICV_14 $T=20240 307360 0 0 $X=20050 $Y=307120
X1431 1 2 525 24 571 571 545 33 ICV_14 $T=20700 280160 0 0 $X=20510 $Y=279920
X1432 1 2 581 10 584 595 585 17 ICV_14 $T=34040 291040 0 0 $X=33850 $Y=290800
X1433 1 2 618 4 669 669 642 17 ICV_14 $T=72680 296480 0 0 $X=72490 $Y=296240
X1434 1 2 92 26 770 770 96 34 ICV_14 $T=118220 307360 0 0 $X=118030 $Y=307120
X1435 1 2 755 14 793 793 772 19 ICV_14 $T=130640 291040 0 0 $X=130450 $Y=290800
X1436 1 2 859 127 911 912 863 131 ICV_14 $T=188600 252960 0 0 $X=188410 $Y=252720
X1437 1 2 899 110 932 932 923 122 ICV_14 $T=200100 291040 1 0 $X=199910 $Y=288080
X1438 1 2 137 110 935 925 144 134 ICV_14 $T=201480 312800 1 0 $X=201290 $Y=309840
X1439 1 2 899 127 943 943 923 134 ICV_14 $T=203320 285600 1 0 $X=203130 $Y=282640
X1440 1 2 983 126 998 998 155 136 ICV_14 $T=230000 247520 1 0 $X=229810 $Y=244560
X1441 1 2 990 108 1015 1015 1012 121 ICV_14 $T=237820 280160 0 0 $X=237630 $Y=279920
X1442 1 2 987 125 1035 1035 986 135 ICV_14 $T=248400 258400 1 0 $X=248210 $Y=255440
X1443 1 2 1231 222 1242 1248 1245 188 ICV_14 $T=359260 307360 1 0 $X=359070 $Y=304400
X1444 1 2 1230 253 1266 1254 1240 201 ICV_14 $T=368000 263840 1 0 $X=367810 $Y=260880
X1445 1 2 1292 218 1315 1315 1299 188 ICV_14 $T=393300 307360 1 0 $X=393110 $Y=304400
X1446 1 2 1349 232 1371 1371 1370 257 ICV_14 $T=420440 252960 1 0 $X=420250 $Y=250000
X1447 1 2 1418 238 1438 1435 1437 263 ICV_14 $T=453100 269280 1 0 $X=452910 $Y=266320
X1448 1 2 1513 357 1518 1523 1519 337 ICV_14 $T=495880 252960 0 0 $X=495690 $Y=252720
X1449 1 2 177 391 397 1579 394 361 ICV_14 $T=525320 301920 0 0 $X=525130 $Y=301680
X1450 1 2 1677 364 1712 1712 1685 372 ICV_14 $T=592940 296480 1 0 $X=592750 $Y=293520
X1451 1 2 1735 224 1751 1715 423 229 ICV_14 $T=609500 252960 1 0 $X=609310 $Y=250000
X1452 1 2 1735 238 1771 1774 435 262 ICV_14 $T=621460 258400 1 0 $X=621270 $Y=255440
X1453 1 2 1791 224 1807 1807 1812 233 ICV_14 $T=637560 252960 1 0 $X=637370 $Y=250000
X1454 1 2 1789 363 1838 1838 1804 303 ICV_14 $T=651360 285600 0 0 $X=651170 $Y=285360
X1455 1 2 1847 368 1896 1896 1853 382 ICV_14 $T=679420 269280 1 0 $X=679230 $Y=266320
X1456 1 2 1900 356 1915 1915 1916 337 ICV_14 $T=691380 258400 0 0 $X=691190 $Y=258160
X1457 1 2 456 399 1933 1928 1926 376 ICV_14 $T=701040 307360 1 0 $X=700850 $Y=304400
X1458 1 2 1946 358 1983 1983 1955 328 ICV_14 $T=729100 269280 1 0 $X=728910 $Y=266320
X1459 1 2 1943 356 1984 1979 1955 337 ICV_14 $T=730020 274720 1 0 $X=729830 $Y=271760
X1460 1 2 1943 358 1986 1986 1965 328 ICV_14 $T=730020 285600 1 0 $X=729830 $Y=282640
X1461 1 2 523 5 535 535 527 16 ICV_16 $T=6900 252960 1 0 $X=6710 $Y=250000
X1462 1 2 764 4 783 783 771 17 ICV_16 $T=126500 258400 0 0 $X=126310 $Y=258160
X1463 1 2 115 125 133 895 116 134 ICV_16 $T=181700 247520 0 0 $X=181510 $Y=247280
X1464 1 2 137 128 939 917 144 121 ICV_16 $T=202400 301920 0 0 $X=202210 $Y=301680
X1465 1 2 137 126 940 940 144 136 ICV_16 $T=202400 307360 1 0 $X=202210 $Y=304400
X1466 1 2 950 125 962 915 923 131 ICV_16 $T=216200 285600 0 0 $X=216010 $Y=285360
X1467 1 2 927 127 963 963 933 134 ICV_16 $T=216660 263840 1 0 $X=216470 $Y=260880
X1468 1 2 979 127 989 989 975 134 ICV_16 $T=228160 296480 1 0 $X=227970 $Y=293520
X1469 1 2 1022 126 1055 1055 1032 136 ICV_16 $T=258520 301920 1 0 $X=258330 $Y=298960
X1470 1 2 1045 126 1058 1043 1012 131 ICV_16 $T=259440 285600 1 0 $X=259250 $Y=282640
X1471 1 2 1045 108 1084 1084 1059 121 ICV_16 $T=272780 280160 1 0 $X=272590 $Y=277200
X1472 1 2 1096 127 1106 1109 1105 136 ICV_16 $T=284280 285600 1 0 $X=284090 $Y=282640
X1473 1 2 1129 112 1161 1161 1146 123 ICV_16 $T=312340 269280 1 0 $X=312150 $Y=266320
X1474 1 2 177 199 206 1188 1199 117 ICV_16 $T=328900 291040 1 0 $X=328710 $Y=288080
X1475 1 2 1230 232 1235 1234 1240 260 ICV_16 $T=356960 269280 0 0 $X=356770 $Y=269040
X1476 1 2 1231 219 1237 1237 1245 202 ICV_16 $T=356960 296480 1 0 $X=356770 $Y=293520
X1477 1 2 258 223 1262 265 267 233 ICV_16 $T=367080 247520 1 0 $X=366890 $Y=244560
X1478 1 2 1369 222 1384 1384 1387 185 ICV_16 $T=426880 301920 1 0 $X=426690 $Y=298960
X1479 1 2 298 214 1388 1388 302 180 ICV_16 $T=427800 312800 1 0 $X=427610 $Y=309840
X1480 1 2 298 218 1390 1390 302 188 ICV_16 $T=428260 307360 1 0 $X=428070 $Y=304400
X1481 1 2 1412 210 1429 1431 1420 202 ICV_16 $T=448960 296480 1 0 $X=448770 $Y=293520
X1482 1 2 326 219 1462 1462 334 202 ICV_16 $T=465520 307360 0 0 $X=465330 $Y=307120
X1483 1 2 1515 356 1530 1530 1534 337 ICV_16 $T=497260 263840 1 0 $X=497070 $Y=260880
X1484 1 2 1570 358 1603 1603 1576 328 ICV_16 $T=539120 252960 0 0 $X=538930 $Y=252720
X1485 1 2 393 358 1607 1607 403 328 ICV_16 $T=539580 247520 1 0 $X=539390 $Y=244560
X1486 1 2 1617 357 1629 1633 1615 337 ICV_16 $T=552000 269280 0 0 $X=551810 $Y=269040
X1487 1 2 1618 358 1636 1636 1635 328 ICV_16 $T=553380 258400 0 0 $X=553190 $Y=258160
X1488 1 2 1618 364 1637 1637 1635 372 ICV_16 $T=553380 263840 1 0 $X=553190 $Y=260880
X1489 1 2 1659 250 1700 1700 1681 262 ICV_16 $T=584200 274720 1 0 $X=584010 $Y=271760
X1490 1 2 1690 385 1725 1725 1701 391 ICV_16 $T=597080 312800 1 0 $X=596890 $Y=309840
X1491 1 2 1714 250 1736 1736 1730 262 ICV_16 $T=602600 258400 0 0 $X=602410 $Y=258160
X1492 1 2 1714 251 1748 1748 1730 263 ICV_16 $T=609500 258400 1 0 $X=609310 $Y=255440
X1493 1 2 1708 224 1749 1749 1723 233 ICV_16 $T=609500 280160 1 0 $X=609310 $Y=277200
X1494 1 2 1708 232 1756 1756 1723 257 ICV_16 $T=610880 280160 0 0 $X=610690 $Y=279920
X1495 1 2 1791 253 1808 1810 1812 263 ICV_16 $T=638480 252960 0 0 $X=638290 $Y=252720
X1496 1 2 1847 367 1892 1892 1853 306 ICV_16 $T=679420 258400 0 0 $X=679230 $Y=258160
X1497 1 2 522 4 532 532 542 17 ICV_17 $T=5520 269280 1 0 $X=5330 $Y=266320
X1498 1 2 522 10 541 533 542 16 ICV_17 $T=6900 263840 0 0 $X=6710 $Y=263600
X1499 1 2 525 26 572 572 545 34 ICV_17 $T=20240 285600 1 0 $X=20050 $Y=282640
X1500 1 2 665 5 673 673 684 16 ICV_17 $T=74520 280160 0 0 $X=74330 $Y=279920
X1501 1 2 708 25 741 741 740 30 ICV_17 $T=103040 285600 0 0 $X=102850 $Y=285360
X1502 1 2 755 24 797 797 772 33 ICV_17 $T=132480 296480 1 0 $X=132290 $Y=293520
X1503 1 2 789 4 812 812 811 17 ICV_17 $T=138920 269280 1 0 $X=138730 $Y=266320
X1504 1 2 809 4 828 827 822 30 ICV_17 $T=145360 285600 1 0 $X=145170 $Y=282640
X1505 1 2 789 24 836 836 811 33 ICV_17 $T=150420 263840 0 0 $X=150230 $Y=263600
X1506 1 2 983 108 1019 1019 155 121 ICV_17 $T=240580 247520 0 0 $X=240390 $Y=247280
X1507 1 2 157 111 162 1029 164 123 ICV_17 $T=248860 312800 1 0 $X=248670 $Y=309840
X1508 1 2 163 127 1050 1050 161 134 ICV_17 $T=256220 247520 1 0 $X=256030 $Y=244560
X1509 1 2 170 127 1132 1126 159 121 ICV_17 $T=293940 247520 0 0 $X=293750 $Y=247280
X1510 1 2 1176 110 1211 1211 1184 122 ICV_17 $T=336260 258400 1 0 $X=336070 $Y=255440
X1511 1 2 1274 223 1313 1316 1277 233 ICV_17 $T=392380 269280 1 0 $X=392190 $Y=266320
X1512 1 2 1321 224 1340 1340 1343 233 ICV_17 $T=406180 258400 0 0 $X=405990 $Y=258160
X1513 1 2 1338 227 1353 1353 1348 252 ICV_17 $T=412620 280160 0 0 $X=412430 $Y=279920
X1514 1 2 299 223 307 1367 1370 201 ICV_17 $T=420440 247520 1 0 $X=420250 $Y=244560
X1515 1 2 1338 223 1373 1373 1348 260 ICV_17 $T=420440 280160 1 0 $X=420250 $Y=277200
X1516 1 2 1349 224 1391 1391 1370 233 ICV_17 $T=427800 258400 1 0 $X=427610 $Y=255440
X1517 1 2 1454 227 1464 1464 1467 252 ICV_17 $T=466440 280160 0 0 $X=466250 $Y=279920
X1518 1 2 1454 250 1472 1472 1467 262 ICV_17 $T=469200 269280 1 0 $X=469010 $Y=266320
X1519 1 2 1459 253 1496 1496 1470 229 ICV_17 $T=482540 258400 1 0 $X=482350 $Y=255440
X1520 1 2 1574 363 1610 1609 1589 328 ICV_17 $T=539120 269280 0 0 $X=538930 $Y=269040
X1521 1 2 1618 363 1628 1628 1635 303 ICV_17 $T=551080 252960 0 0 $X=550890 $Y=252720
X1522 1 2 1672 223 1709 1710 1688 233 ICV_17 $T=588800 269280 1 0 $X=588610 $Y=266320
X1523 1 2 1763 224 1772 1767 1739 303 ICV_17 $T=621000 285600 1 0 $X=620810 $Y=282640
X1524 1 2 1763 238 1782 1782 1761 201 ICV_17 $T=623300 269280 1 0 $X=623110 $Y=266320
X1525 1 2 1791 250 1829 1828 444 257 ICV_17 $T=649980 252960 1 0 $X=649790 $Y=250000
X1526 1 2 1791 223 1833 1829 1812 262 ICV_17 $T=650440 258400 1 0 $X=650250 $Y=255440
X1527 1 2 1820 388 1857 1858 1824 370 ICV_17 $T=661020 301920 0 0 $X=660830 $Y=301680
X1528 1 2 1846 358 1867 1867 1859 328 ICV_17 $T=665620 247520 1 0 $X=665430 $Y=244560
X1529 1 2 1846 356 1868 1868 1859 337 ICV_17 $T=665620 252960 1 0 $X=665430 $Y=250000
X1530 1 2 1846 363 1891 1891 1859 303 ICV_17 $T=678500 252960 1 0 $X=678310 $Y=250000
X1531 1 2 450 363 1913 1913 453 303 ICV_17 $T=687240 247520 0 0 $X=687050 $Y=247280
X1532 1 2 1886 357 1927 1925 1904 372 ICV_17 $T=697820 291040 1 0 $X=697630 $Y=288080
X1533 1 2 1951 367 1949 1967 1955 372 ICV_17 $T=717140 258400 0 0 $X=716950 $Y=258160
X1556 1 2 524 11 544 544 543 18 ICV_19 $T=6900 307360 0 0 $X=6710 $Y=307120
X1557 1 2 582 26 612 608 578 19 ICV_19 $T=43240 269280 0 0 $X=43050 $Y=269040
X1558 1 2 617 5 655 655 641 16 ICV_19 $T=62100 285600 0 0 $X=61910 $Y=285360
X1559 1 2 861 111 877 879 862 122 ICV_19 $T=171120 274720 1 0 $X=170930 $Y=271760
X1560 1 2 141 110 968 968 146 122 ICV_19 $T=216660 247520 1 0 $X=216470 $Y=244560
X1561 1 2 950 126 969 969 954 136 ICV_19 $T=216660 291040 1 0 $X=216470 $Y=288080
X1562 1 2 177 186 191 1171 1123 123 ICV_19 $T=314640 285600 0 0 $X=314450 $Y=285360
X1563 1 2 1256 250 1272 1272 1273 262 ICV_19 $T=370760 252960 0 0 $X=370570 $Y=252720
X1564 1 2 284 223 1327 1325 293 233 ICV_19 $T=398820 252960 0 0 $X=398630 $Y=252720
X1565 1 2 1321 238 1389 1389 1343 201 ICV_19 $T=426880 263840 0 0 $X=426690 $Y=263600
X1566 1 2 1380 224 1407 1407 1406 233 ICV_19 $T=434240 280160 0 0 $X=434050 $Y=279920
X1567 1 2 326 210 1488 1488 334 199 ICV_19 $T=476560 307360 1 0 $X=476370 $Y=304400
X1568 1 2 1514 364 1552 1552 1532 372 ICV_19 $T=508760 291040 1 0 $X=508570 $Y=288080
X1569 1 2 177 400 405 1599 394 375 ICV_19 $T=532680 301920 1 0 $X=532490 $Y=298960
X1570 1 2 1574 356 1611 1611 1589 337 ICV_19 $T=539120 274720 0 0 $X=538930 $Y=274480
X1571 1 2 1618 356 1668 1668 1635 337 ICV_19 $T=567180 258400 0 0 $X=566990 $Y=258160
X1572 1 2 1641 399 1683 1683 1656 370 ICV_19 $T=574540 301920 0 0 $X=574350 $Y=301680
X1573 1 2 1690 388 1729 1729 1701 361 ICV_19 $T=596620 301920 0 0 $X=596430 $Y=301680
X1574 1 2 1734 356 1766 1764 1739 372 ICV_19 $T=616860 296480 1 0 $X=616670 $Y=293520
X1575 1 2 1848 357 1861 1861 1866 348 ICV_19 $T=663320 291040 0 0 $X=663130 $Y=290800
X1576 1 2 1848 364 1880 1884 1866 337 ICV_19 $T=672980 296480 1 0 $X=672790 $Y=293520
X1577 1 2 1886 367 1920 1920 1904 306 ICV_19 $T=693220 285600 0 0 $X=693030 $Y=285360
X1578 1 2 1951 356 471 1988 463 382 ICV_19 $T=729100 258400 1 0 $X=728910 $Y=255440
X1579 1 2 1951 363 1973 1989 1955 382 ICV_19 $T=729100 263840 1 0 $X=728910 $Y=260880
X1580 1 2 1943 363 1985 1985 1965 303 ICV_19 $T=729100 280160 1 0 $X=728910 $Y=277200
X1581 1 2 32 26 603 ICV_20 $T=40020 247520 1 0 $X=39830 $Y=244560
X1582 1 2 42 24 611 ICV_20 $T=44160 301920 0 0 $X=43970 $Y=301680
X1583 1 2 582 10 616 ICV_20 $T=45540 280160 0 0 $X=45350 $Y=279920
X1584 1 2 619 11 55 ICV_20 $T=53820 247520 0 0 $X=53630 $Y=247280
X1585 1 2 619 4 59 ICV_20 $T=56120 247520 1 0 $X=55930 $Y=244560
X1586 1 2 628 4 645 ICV_20 $T=59340 269280 1 0 $X=59150 $Y=266320
X1587 1 2 628 11 647 ICV_20 $T=59800 263840 1 0 $X=59610 $Y=260880
X1588 1 2 619 14 651 ICV_20 $T=62100 247520 0 0 $X=61910 $Y=247280
X1589 1 2 62 14 660 ICV_20 $T=66240 307360 0 0 $X=66050 $Y=307120
X1590 1 2 62 26 65 ICV_20 $T=66700 312800 1 0 $X=66510 $Y=309840
X1591 1 2 670 24 688 ICV_20 $T=80500 258400 0 0 $X=80310 $Y=258160
X1592 1 2 670 25 692 ICV_20 $T=81420 247520 0 0 $X=81230 $Y=247280
X1593 1 2 665 4 696 ICV_20 $T=87860 285600 1 0 $X=87670 $Y=282640
X1594 1 2 685 10 722 ICV_20 $T=95680 307360 1 0 $X=95490 $Y=304400
X1595 1 2 738 14 752 ICV_20 $T=109940 301920 0 0 $X=109750 $Y=301680
X1596 1 2 744 24 759 ICV_20 $T=113160 263840 1 0 $X=112970 $Y=260880
X1597 1 2 744 26 760 ICV_20 $T=113160 269280 1 0 $X=112970 $Y=266320
X1598 1 2 761 24 777 ICV_20 $T=120520 285600 1 0 $X=120330 $Y=282640
X1599 1 2 92 10 782 ICV_20 $T=124200 312800 1 0 $X=124010 $Y=309840
X1600 1 2 761 11 806 ICV_20 $T=136620 280160 0 0 $X=136430 $Y=279920
X1601 1 2 809 25 827 ICV_20 $T=146280 280160 0 0 $X=146090 $Y=279920
X1602 1 2 810 11 820 ICV_20 $T=146280 291040 0 0 $X=146090 $Y=290800
X1603 1 2 809 10 848 ICV_20 $T=156400 280160 0 0 $X=156210 $Y=279920
X1604 1 2 109 108 870 ICV_20 $T=167900 307360 1 0 $X=167710 $Y=304400
X1605 1 2 859 110 868 ICV_20 $T=168360 263840 1 0 $X=168170 $Y=260880
X1606 1 2 919 112 938 ICV_20 $T=202400 269280 0 0 $X=202210 $Y=269040
X1607 1 2 927 128 946 ICV_20 $T=204700 263840 0 0 $X=204510 $Y=263600
X1608 1 2 906 128 148 ICV_20 $T=206540 296480 0 0 $X=206350 $Y=296240
X1609 1 2 919 126 951 ICV_20 $T=209760 274720 0 0 $X=209570 $Y=274480
X1610 1 2 950 128 978 ICV_20 $T=221260 291040 0 0 $X=221070 $Y=290800
X1611 1 2 983 128 1003 ICV_20 $T=232760 252960 0 0 $X=232570 $Y=252720
X1612 1 2 956 128 1005 ICV_20 $T=232760 263840 0 0 $X=232570 $Y=263600
X1613 1 2 956 111 1010 ICV_20 $T=234600 269280 1 0 $X=234410 $Y=266320
X1614 1 2 956 125 1011 ICV_20 $T=234600 269280 0 0 $X=234410 $Y=269040
X1615 1 2 153 110 1008 ICV_20 $T=234600 307360 1 0 $X=234410 $Y=304400
X1616 1 2 157 112 1029 ICV_20 $T=246560 307360 0 0 $X=246370 $Y=307120
X1617 1 2 1020 127 1057 ICV_20 $T=261740 269280 1 0 $X=261550 $Y=266320
X1618 1 2 1022 112 1065 ICV_20 $T=262660 301920 0 0 $X=262470 $Y=301680
X1619 1 2 1054 110 1072 ICV_20 $T=267720 258400 0 0 $X=267530 $Y=258160
X1620 1 2 1054 111 1092 ICV_20 $T=276460 252960 0 0 $X=276270 $Y=252720
X1621 1 2 166 128 1091 ICV_20 $T=277380 307360 1 0 $X=277190 $Y=304400
X1622 1 2 170 112 1118 ICV_20 $T=288880 252960 1 0 $X=288690 $Y=250000
X1623 1 2 170 110 1125 ICV_20 $T=291640 258400 1 0 $X=291450 $Y=255440
X1624 1 2 1096 112 1128 ICV_20 $T=293020 285600 0 0 $X=292830 $Y=285360
X1625 1 2 1097 125 1139 ICV_20 $T=297620 274720 0 0 $X=297430 $Y=274480
X1626 1 2 1116 126 1152 ICV_20 $T=306360 296480 0 0 $X=306170 $Y=296240
X1627 1 2 1116 111 1153 ICV_20 $T=306360 301920 0 0 $X=306170 $Y=301680
X1628 1 2 1129 128 1164 ICV_20 $T=314180 263840 1 0 $X=313990 $Y=260880
X1629 1 2 177 185 190 ICV_20 $T=314640 291040 0 0 $X=314450 $Y=290800
X1630 1 2 1176 125 1190 ICV_20 $T=327980 263840 0 0 $X=327790 $Y=263600
X1631 1 2 1176 128 1209 ICV_20 $T=336260 269280 1 0 $X=336070 $Y=266320
X1632 1 2 1180 110 1210 ICV_20 $T=339480 285600 1 0 $X=339290 $Y=282640
X1633 1 2 1180 127 1229 ICV_20 $T=349600 280160 0 0 $X=349410 $Y=279920
X1634 1 2 1230 223 1234 ICV_20 $T=356960 269280 1 0 $X=356770 $Y=266320
X1635 1 2 1258 222 1279 ICV_20 $T=374440 301920 1 0 $X=374250 $Y=298960
X1636 1 2 1274 238 1287 ICV_20 $T=379040 263840 0 0 $X=378850 $Y=263600
X1637 1 2 1290 251 1301 ICV_20 $T=388240 269280 0 0 $X=388050 $Y=269040
X1638 1 2 1292 217 1305 ICV_20 $T=389160 296480 0 0 $X=388970 $Y=296240
X1639 1 2 275 218 1309 ICV_20 $T=390540 307360 0 0 $X=390350 $Y=307120
X1640 1 2 284 232 291 ICV_20 $T=401120 247520 1 0 $X=400930 $Y=244560
X1641 1 2 275 210 1331 ICV_20 $T=402500 312800 1 0 $X=402310 $Y=309840
X1642 1 2 1290 253 1337 ICV_20 $T=404800 280160 1 0 $X=404610 $Y=277200
X1643 1 2 1322 214 1362 ICV_20 $T=416300 296480 0 0 $X=416110 $Y=296240
X1644 1 2 1369 210 1383 ICV_20 $T=426880 291040 0 0 $X=426690 $Y=290800
X1645 1 2 1349 251 1393 ICV_20 $T=432860 252960 1 0 $X=432670 $Y=250000
X1646 1 2 1396 253 1397 ICV_20 $T=441140 258400 1 0 $X=440950 $Y=255440
X1647 1 2 316 232 1419 ICV_20 $T=446660 252960 0 0 $X=446470 $Y=252720
X1648 1 2 1412 217 1422 ICV_20 $T=446660 296480 0 0 $X=446470 $Y=296240
X1649 1 2 316 251 1428 ICV_20 $T=448960 258400 1 0 $X=448770 $Y=255440
X1650 1 2 1441 217 1455 ICV_20 $T=460920 296480 1 0 $X=460730 $Y=293520
X1651 1 2 1441 213 1446 ICV_20 $T=462300 301920 0 0 $X=462110 $Y=301680
X1652 1 2 336 238 339 ICV_20 $T=474260 247520 0 0 $X=474070 $Y=247280
X1653 1 2 1491 219 1509 ICV_20 $T=487140 291040 0 0 $X=486950 $Y=290800
X1654 1 2 336 227 353 ICV_20 $T=487600 247520 0 0 $X=487410 $Y=247280
X1655 1 2 347 213 1510 ICV_20 $T=488060 312800 1 0 $X=487870 $Y=309840
X1656 1 2 347 210 1537 ICV_20 $T=500480 307360 0 0 $X=500290 $Y=307120
X1657 1 2 1513 363 1544 ICV_20 $T=504620 258400 1 0 $X=504430 $Y=255440
X1658 1 2 1515 357 1562 ICV_20 $T=516580 263840 1 0 $X=516390 $Y=260880
X1659 1 2 1572 367 1582 ICV_20 $T=525320 280160 0 0 $X=525130 $Y=279920
X1660 1 2 1574 367 1588 ICV_20 $T=528080 274720 0 0 $X=527890 $Y=274480
X1661 1 2 1570 364 1591 ICV_20 $T=529920 258400 0 0 $X=529730 $Y=258160
X1662 1 2 409 388 1642 ICV_20 $T=555680 307360 0 0 $X=555490 $Y=307120
X1663 1 2 1618 357 1644 ICV_20 $T=557060 258400 1 0 $X=556870 $Y=255440
X1664 1 2 424 251 1721 ICV_20 $T=597540 252960 1 0 $X=597350 $Y=250000
X1665 1 2 1734 357 1741 ICV_20 $T=606740 291040 0 0 $X=606550 $Y=290800
X1666 1 2 1735 253 438 ICV_20 $T=623300 247520 0 0 $X=623110 $Y=247280
X1667 1 2 1788 253 1806 ICV_20 $T=637560 269280 0 0 $X=637370 $Y=269040
X1668 1 2 1793 251 1816 ICV_20 $T=639860 274720 1 0 $X=639670 $Y=271760
X1669 1 2 1789 358 1818 ICV_20 $T=640780 285600 0 0 $X=640590 $Y=285360
X1670 1 2 1886 356 1903 ICV_20 $T=685400 291040 1 0 $X=685210 $Y=288080
X1671 1 2 1893 359 1906 ICV_20 $T=686320 269280 0 0 $X=686130 $Y=269040
X1672 1 2 1893 357 1921 ICV_20 $T=695520 269280 0 0 $X=695330 $Y=269040
X1673 1 2 1886 363 1923 ICV_20 $T=697820 285600 1 0 $X=697630 $Y=282640
X1674 1 2 1886 364 1925 ICV_20 $T=697820 291040 0 0 $X=697630 $Y=290800
X1675 1 2 456 388 1938 ICV_20 $T=701960 301920 1 0 $X=701770 $Y=298960
X1676 1 2 1943 367 1952 ICV_20 $T=711620 280160 0 0 $X=711430 $Y=279920
X1677 1 2 456 418 1958 ICV_20 $T=713460 307360 1 0 $X=713270 $Y=304400
X1678 1 2 1944 356 1981 ICV_20 $T=727260 291040 0 0 $X=727070 $Y=290800
X1679 1 2 522 11 550 ICV_21 $T=6900 263840 1 0 $X=6710 $Y=260880
X1680 1 2 581 24 613 ICV_21 $T=41400 285600 0 0 $X=41210 $Y=285360
X1681 1 2 707 10 723 ICV_21 $T=93380 274720 1 0 $X=93190 $Y=271760
X1682 1 2 744 14 762 ICV_21 $T=111780 274720 1 0 $X=111590 $Y=271760
X1683 1 2 761 4 778 ICV_21 $T=118220 274720 0 0 $X=118030 $Y=274480
X1684 1 2 744 10 780 ICV_21 $T=120980 269280 1 0 $X=120790 $Y=266320
X1685 1 2 813 11 834 ICV_21 $T=146280 247520 1 0 $X=146090 $Y=244560
X1686 1 2 115 112 124 ICV_21 $T=168820 247520 1 0 $X=168630 $Y=244560
X1687 1 2 906 125 908 ICV_21 $T=190440 296480 0 0 $X=190250 $Y=296240
X1688 1 2 157 110 1034 ICV_21 $T=244720 307360 1 0 $X=244530 $Y=304400
X1689 1 2 1022 125 1031 ICV_21 $T=247480 291040 0 0 $X=247290 $Y=290800
X1690 1 2 166 125 167 ICV_21 $T=261740 312800 1 0 $X=261550 $Y=309840
X1691 1 2 170 111 173 ICV_21 $T=280140 247520 1 0 $X=279950 $Y=244560
X1692 1 2 171 126 175 ICV_21 $T=293940 307360 0 0 $X=293750 $Y=307120
X1693 1 2 1231 217 1238 ICV_21 $T=354200 296480 0 0 $X=354010 $Y=296240
X1694 1 2 1418 227 1432 ICV_21 $T=448500 285600 1 0 $X=448310 $Y=282640
X1695 1 2 1459 250 1475 ICV_21 $T=468280 252960 0 0 $X=468090 $Y=252720
X1696 1 2 177 375 381 ICV_21 $T=511060 301920 0 0 $X=510870 $Y=301680
X1697 1 2 1515 363 1565 ICV_21 $T=514280 269280 1 0 $X=514090 $Y=266320
X1698 1 2 1572 359 1577 ICV_21 $T=522100 285600 0 0 $X=521910 $Y=285360
X1699 1 2 1630 357 1652 ICV_21 $T=560740 296480 1 0 $X=560550 $Y=293520
X1700 1 2 1873 390 1899 ICV_21 $T=682640 312800 1 0 $X=682450 $Y=309840
X1701 1 2 450 358 1922 ICV_21 $T=693680 247520 1 0 $X=693490 $Y=244560
X1702 1 2 1944 359 1957 ICV_21 $T=710700 291040 1 0 $X=710510 $Y=288080
X1703 1 2 525 11 546 546 545 18 ICV_22 $T=6900 280160 0 0 $X=6710 $Y=279920
X1704 1 2 530 10 547 549 555 17 ICV_22 $T=6900 296480 0 0 $X=6710 $Y=296240
X1705 1 2 32 14 609 52 45 16 ICV_22 $T=41400 252960 0 0 $X=41210 $Y=252720
X1706 1 2 62 5 675 682 66 33 ICV_22 $T=74060 307360 0 0 $X=73870 $Y=307120
X1707 1 2 738 5 753 753 757 16 ICV_22 $T=108560 301920 1 0 $X=108370 $Y=298960
X1708 1 2 764 24 798 798 771 33 ICV_22 $T=132480 258400 1 0 $X=132290 $Y=255440
X1709 1 2 809 24 846 847 822 16 ICV_22 $T=153640 274720 0 0 $X=153450 $Y=274480
X1710 1 2 137 112 916 887 119 135 ICV_22 $T=188600 307360 1 0 $X=188410 $Y=304400
X1711 1 2 906 127 944 934 923 117 ICV_22 $T=201940 296480 1 0 $X=201750 $Y=293520
X1712 1 2 899 112 945 945 923 123 ICV_22 $T=202400 285600 0 0 $X=202210 $Y=285360
X1713 1 2 153 127 971 971 154 134 ICV_22 $T=216660 307360 1 0 $X=216470 $Y=304400
X1714 1 2 950 110 988 988 954 122 ICV_22 $T=224020 285600 1 0 $X=223830 $Y=282640
X1715 1 2 1045 111 1080 1080 1059 117 ICV_22 $T=269560 280160 0 0 $X=269370 $Y=279920
X1716 1 2 176 112 1154 1154 184 123 ICV_22 $T=305440 247520 1 0 $X=305250 $Y=244560
X1717 1 2 1230 251 1244 1244 1240 263 ICV_22 $T=356040 263840 0 0 $X=355850 $Y=263600
X1718 1 2 1290 227 1328 1328 1312 252 ICV_22 $T=398820 280160 0 0 $X=398630 $Y=279920
X1719 1 2 1515 367 1571 1562 1534 348 ICV_22 $T=516120 258400 0 0 $X=515930 $Y=258160
X1720 1 2 1641 390 1658 1667 1656 375 ICV_22 $T=563960 312800 1 0 $X=563770 $Y=309840
X1721 1 2 1735 251 1743 1743 435 263 ICV_22 $T=606740 247520 0 0 $X=606550 $Y=247280
X1722 1 2 1820 404 1827 1827 1824 389 ICV_22 $T=648600 301920 1 0 $X=648410 $Y=298960
X1723 1 2 1841 359 1881 1881 1844 341 ICV_22 $T=672980 280160 1 0 $X=672790 $Y=277200
X1724 1 2 1873 404 1882 1882 1875 389 ICV_22 $T=672980 301920 1 0 $X=672790 $Y=298960
X1725 1 2 1900 368 1939 1940 1916 348 ICV_22 $T=701040 263840 1 0 $X=700850 $Y=260880
X1726 1 2 456 404 1963 1961 1926 375 ICV_22 $T=712540 301920 0 0 $X=712350 $Y=301680
X1727 1 2 1946 367 1964 1964 1955 306 ICV_22 $T=713000 269280 0 0 $X=712810 $Y=269040
X1728 1 2 ICV_23 $T=18400 269280 1 0 $X=18210 $Y=266320
X1729 1 2 ICV_23 $T=32200 247520 0 0 $X=32010 $Y=247280
X1730 1 2 ICV_23 $T=46460 301920 1 0 $X=46270 $Y=298960
X1731 1 2 ICV_23 $T=74520 296480 1 0 $X=74330 $Y=293520
X1732 1 2 ICV_23 $T=74520 312800 1 0 $X=74330 $Y=309840
X1733 1 2 ICV_23 $T=88320 252960 0 0 $X=88130 $Y=252720
X1734 1 2 ICV_23 $T=88320 258400 0 0 $X=88130 $Y=258160
X1735 1 2 ICV_23 $T=102580 280160 1 0 $X=102390 $Y=277200
X1736 1 2 ICV_23 $T=144440 280160 0 0 $X=144250 $Y=279920
X1737 1 2 ICV_23 $T=144440 291040 0 0 $X=144250 $Y=290800
X1738 1 2 ICV_23 $T=214820 291040 1 0 $X=214630 $Y=288080
X1739 1 2 ICV_23 $T=270940 291040 1 0 $X=270750 $Y=288080
X1740 1 2 ICV_23 $T=299000 263840 1 0 $X=298810 $Y=260880
X1741 1 2 ICV_23 $T=312800 269280 0 0 $X=312610 $Y=269040
X1742 1 2 ICV_23 $T=340860 247520 0 0 $X=340670 $Y=247280
X1743 1 2 ICV_23 $T=340860 258400 0 0 $X=340670 $Y=258160
X1744 1 2 ICV_23 $T=340860 291040 0 0 $X=340670 $Y=290800
X1745 1 2 ICV_23 $T=355120 296480 1 0 $X=354930 $Y=293520
X1746 1 2 ICV_23 $T=355120 307360 1 0 $X=354930 $Y=304400
X1747 1 2 ICV_23 $T=368920 280160 0 0 $X=368730 $Y=279920
X1748 1 2 ICV_23 $T=368920 291040 0 0 $X=368730 $Y=290800
X1749 1 2 ICV_23 $T=453100 280160 0 0 $X=452910 $Y=279920
X1750 1 2 ICV_23 $T=453100 291040 0 0 $X=452910 $Y=290800
X1751 1 2 ICV_23 $T=467360 258400 1 0 $X=467170 $Y=255440
X1752 1 2 ICV_23 $T=467360 280160 1 0 $X=467170 $Y=277200
X1753 1 2 ICV_23 $T=509220 258400 0 0 $X=509030 $Y=258160
X1754 1 2 ICV_23 $T=509220 285600 0 0 $X=509030 $Y=285360
X1755 1 2 ICV_23 $T=509220 301920 0 0 $X=509030 $Y=301680
X1756 1 2 ICV_23 $T=537280 252960 0 0 $X=537090 $Y=252720
X1757 1 2 ICV_23 $T=537280 285600 0 0 $X=537090 $Y=285360
X1758 1 2 ICV_23 $T=551540 252960 1 0 $X=551350 $Y=250000
X1759 1 2 ICV_23 $T=565340 258400 0 0 $X=565150 $Y=258160
X1760 1 2 ICV_23 $T=579600 247520 1 0 $X=579410 $Y=244560
X1761 1 2 ICV_23 $T=607660 252960 1 0 $X=607470 $Y=250000
X1762 1 2 ICV_23 $T=607660 274720 1 0 $X=607470 $Y=271760
X1763 1 2 ICV_23 $T=635720 296480 1 0 $X=635530 $Y=293520
X1764 1 2 ICV_23 $T=649520 301920 0 0 $X=649330 $Y=301680
X1765 1 2 ICV_23 $T=691840 269280 1 0 $X=691650 $Y=266320
X1766 1 2 ICV_23 $T=691840 296480 1 0 $X=691650 $Y=293520
X1767 1 2 ICV_23 $T=705640 274720 0 0 $X=705450 $Y=274480
X1768 1 2 ICV_23 $T=705640 291040 0 0 $X=705450 $Y=290800
X1769 1 2 ICV_23 $T=733700 307360 0 0 $X=733510 $Y=307120
X1770 1 2 ICV_24 $T=17940 274720 1 0 $X=17750 $Y=271760
X1771 1 2 ICV_24 $T=87860 291040 0 0 $X=87670 $Y=290800
X1772 1 2 ICV_24 $T=87860 307360 0 0 $X=87670 $Y=307120
X1773 1 2 ICV_24 $T=115920 263840 0 0 $X=115730 $Y=263600
X1774 1 2 ICV_24 $T=115920 280160 0 0 $X=115730 $Y=279920
X1775 1 2 ICV_24 $T=130180 274720 1 0 $X=129990 $Y=271760
X1776 1 2 ICV_24 $T=158240 285600 1 0 $X=158050 $Y=282640
X1777 1 2 ICV_24 $T=158240 291040 1 0 $X=158050 $Y=288080
X1778 1 2 ICV_24 $T=158240 301920 1 0 $X=158050 $Y=298960
X1779 1 2 ICV_24 $T=214360 258400 1 0 $X=214170 $Y=255440
X1780 1 2 ICV_24 $T=214360 307360 1 0 $X=214170 $Y=304400
X1781 1 2 ICV_24 $T=228160 285600 0 0 $X=227970 $Y=285360
X1782 1 2 ICV_24 $T=242420 247520 1 0 $X=242230 $Y=244560
X1783 1 2 ICV_24 $T=242420 307360 1 0 $X=242230 $Y=304400
X1784 1 2 ICV_24 $T=284280 252960 0 0 $X=284090 $Y=252720
X1785 1 2 ICV_24 $T=298540 301920 1 0 $X=298350 $Y=298960
X1786 1 2 ICV_24 $T=312340 285600 0 0 $X=312150 $Y=285360
X1787 1 2 ICV_24 $T=368460 307360 0 0 $X=368270 $Y=307120
X1788 1 2 ICV_24 $T=396520 285600 0 0 $X=396330 $Y=285360
X1789 1 2 ICV_24 $T=438840 301920 1 0 $X=438650 $Y=298960
X1790 1 2 ICV_24 $T=494960 247520 1 0 $X=494770 $Y=244560
X1791 1 2 ICV_24 $T=508760 296480 0 0 $X=508570 $Y=296240
X1792 1 2 ICV_24 $T=551080 258400 1 0 $X=550890 $Y=255440
X1793 1 2 ICV_24 $T=551080 263840 1 0 $X=550890 $Y=260880
X1794 1 2 ICV_24 $T=635260 247520 1 0 $X=635070 $Y=244560
X1795 1 2 ICV_24 $T=649060 263840 0 0 $X=648870 $Y=263600
X1796 1 2 ICV_24 $T=663320 258400 1 0 $X=663130 $Y=255440
X1797 1 2 ICV_24 $T=663320 291040 1 0 $X=663130 $Y=288080
X1798 1 2 ICV_24 $T=691380 247520 1 0 $X=691190 $Y=244560
X1799 1 2 ICV_24 $T=691380 252960 1 0 $X=691190 $Y=250000
X1800 1 2 15 2 527 1 sky130_fd_sc_hd__inv_1 $T=25300 252960 1 0 $X=25110 $Y=250000
X1801 1 2 6 2 23 1 sky130_fd_sc_hd__inv_1 $T=25760 247520 1 0 $X=25570 $Y=244560
X1802 1 2 20 2 542 1 sky130_fd_sc_hd__inv_1 $T=25760 274720 1 0 $X=25570 $Y=271760
X1803 1 2 3 2 545 1 sky130_fd_sc_hd__inv_1 $T=29900 285600 0 0 $X=29710 $Y=285360
X1804 1 2 36 2 543 1 sky130_fd_sc_hd__inv_1 $T=31740 307360 1 0 $X=31550 $Y=304400
X1805 1 2 8 2 555 1 sky130_fd_sc_hd__inv_1 $T=33120 296480 1 0 $X=32930 $Y=293520
X1806 1 2 44 2 29 1 sky130_fd_sc_hd__inv_1 $T=40940 312800 1 0 $X=40750 $Y=309840
X1807 1 2 49 2 578 1 sky130_fd_sc_hd__inv_1 $T=49220 274720 1 0 $X=49030 $Y=271760
X1808 1 2 40 2 602 1 sky130_fd_sc_hd__inv_1 $T=50600 285600 1 0 $X=50410 $Y=282640
X1809 1 2 35 2 585 1 sky130_fd_sc_hd__inv_1 $T=50600 291040 0 0 $X=50410 $Y=290800
X1810 1 2 53 2 45 1 sky130_fd_sc_hd__inv_1 $T=52440 252960 1 0 $X=52250 $Y=250000
X1811 1 2 54 2 47 1 sky130_fd_sc_hd__inv_1 $T=60260 307360 0 0 $X=60070 $Y=307120
X1812 1 2 57 2 641 1 sky130_fd_sc_hd__inv_1 $T=67620 280160 1 0 $X=67430 $Y=277200
X1813 1 2 63 2 642 1 sky130_fd_sc_hd__inv_1 $T=73140 296480 1 0 $X=72950 $Y=293520
X1814 1 2 60 2 56 1 sky130_fd_sc_hd__inv_1 $T=74520 252960 1 0 $X=74330 $Y=250000
X1815 1 2 48 2 627 1 sky130_fd_sc_hd__inv_1 $T=80960 263840 0 0 $X=80770 $Y=263600
X1816 1 2 58 2 66 1 sky130_fd_sc_hd__inv_1 $T=83720 307360 1 0 $X=83530 $Y=304400
X1817 1 2 64 2 676 1 sky130_fd_sc_hd__inv_1 $T=87400 274720 0 0 $X=87210 $Y=274480
X1818 1 2 73 2 693 1 sky130_fd_sc_hd__inv_1 $T=90620 301920 0 0 $X=90430 $Y=301680
X1819 1 2 72 2 690 1 sky130_fd_sc_hd__inv_1 $T=97520 263840 0 0 $X=97330 $Y=263600
X1820 1 2 67 2 684 1 sky130_fd_sc_hd__inv_1 $T=101660 285600 0 0 $X=101470 $Y=285360
X1821 1 2 76 2 730 1 sky130_fd_sc_hd__inv_1 $T=111780 269280 1 0 $X=111590 $Y=266320
X1822 1 2 80 2 740 1 sky130_fd_sc_hd__inv_1 $T=115920 285600 0 0 $X=115730 $Y=285360
X1823 1 2 83 2 74 1 sky130_fd_sc_hd__inv_1 $T=120520 258400 1 0 $X=120330 $Y=255440
X1824 1 2 90 2 718 1 sky130_fd_sc_hd__inv_1 $T=128800 274720 1 0 $X=128610 $Y=271760
X1825 1 2 86 2 757 1 sky130_fd_sc_hd__inv_1 $T=139380 301920 1 0 $X=139190 $Y=298960
X1826 1 2 88 2 772 1 sky130_fd_sc_hd__inv_1 $T=143060 291040 0 0 $X=142870 $Y=290800
X1827 1 2 99 2 779 1 sky130_fd_sc_hd__inv_1 $T=143980 285600 1 0 $X=143790 $Y=282640
X1828 1 2 94 2 771 1 sky130_fd_sc_hd__inv_1 $T=146280 252960 0 0 $X=146090 $Y=252720
X1829 1 2 102 2 824 1 sky130_fd_sc_hd__inv_1 $T=156860 301920 1 0 $X=156670 $Y=298960
X1830 1 2 104 2 822 1 sky130_fd_sc_hd__inv_1 $T=161460 274720 1 0 $X=161270 $Y=271760
X1831 1 2 98 2 811 1 sky130_fd_sc_hd__inv_1 $T=163300 263840 0 0 $X=163110 $Y=263600
X1832 1 2 103 2 835 1 sky130_fd_sc_hd__inv_1 $T=166060 252960 0 0 $X=165870 $Y=252720
X1833 1 2 106 2 89 1 sky130_fd_sc_hd__inv_1 $T=166520 312800 1 0 $X=166330 $Y=309840
X1834 1 2 20 2 862 1 sky130_fd_sc_hd__inv_1 $T=172040 269280 0 0 $X=171850 $Y=269040
X1835 1 2 48 2 863 1 sky130_fd_sc_hd__inv_1 $T=172500 263840 0 0 $X=172310 $Y=263600
X1836 1 2 15 2 116 1 sky130_fd_sc_hd__inv_1 $T=174340 252960 0 0 $X=174150 $Y=252720
X1837 1 2 36 2 873 1 sky130_fd_sc_hd__inv_1 $T=175720 301920 1 0 $X=175530 $Y=298960
X1838 1 2 3 2 874 1 sky130_fd_sc_hd__inv_1 $T=186300 285600 1 0 $X=186110 $Y=282640
X1839 1 2 8 2 923 1 sky130_fd_sc_hd__inv_1 $T=198720 291040 1 0 $X=198530 $Y=288080
X1840 1 2 44 2 139 1 sky130_fd_sc_hd__inv_1 $T=200100 301920 0 0 $X=199910 $Y=301680
X1841 1 2 57 2 921 1 sky130_fd_sc_hd__inv_1 $T=200560 280160 0 0 $X=200370 $Y=279920
X1842 1 2 28 2 146 1 sky130_fd_sc_hd__inv_1 $T=206540 252960 1 0 $X=206350 $Y=250000
X1843 1 2 49 2 933 1 sky130_fd_sc_hd__inv_1 $T=208380 269280 1 0 $X=208190 $Y=266320
X1844 1 2 35 2 954 1 sky130_fd_sc_hd__inv_1 $T=219880 291040 0 0 $X=219690 $Y=290800
X1845 1 2 64 2 973 1 sky130_fd_sc_hd__inv_1 $T=225400 274720 1 0 $X=225210 $Y=271760
X1846 1 2 60 2 155 1 sky130_fd_sc_hd__inv_1 $T=229080 252960 1 0 $X=228890 $Y=250000
X1847 1 2 58 2 975 1 sky130_fd_sc_hd__inv_1 $T=230460 307360 0 0 $X=230270 $Y=307120
X1848 1 2 76 2 986 1 sky130_fd_sc_hd__inv_1 $T=231840 258400 0 0 $X=231650 $Y=258160
X1849 1 2 40 2 1012 1 sky130_fd_sc_hd__inv_1 $T=242420 285600 0 0 $X=242230 $Y=285360
X1850 1 2 90 2 1027 1 sky130_fd_sc_hd__inv_1 $T=251160 269280 1 0 $X=250970 $Y=266320
X1851 1 2 160 2 161 1 sky130_fd_sc_hd__inv_1 $T=256220 252960 1 0 $X=256030 $Y=250000
X1852 1 2 72 2 1053 1 sky130_fd_sc_hd__inv_1 $T=264960 258400 1 0 $X=264770 $Y=255440
X1853 1 2 63 2 1059 1 sky130_fd_sc_hd__inv_1 $T=269100 285600 0 0 $X=268910 $Y=285360
X1854 1 2 86 2 1032 1 sky130_fd_sc_hd__inv_1 $T=270480 301920 1 0 $X=270290 $Y=298960
X1855 1 2 73 2 1086 1 sky130_fd_sc_hd__inv_1 $T=287040 301920 0 0 $X=286850 $Y=301680
X1856 1 2 83 2 159 1 sky130_fd_sc_hd__inv_1 $T=288880 252960 0 0 $X=288690 $Y=252720
X1857 1 2 67 2 1104 1 sky130_fd_sc_hd__inv_1 $T=289800 280160 1 0 $X=289610 $Y=277200
X1858 1 2 88 2 1105 1 sky130_fd_sc_hd__inv_1 $T=290720 291040 0 0 $X=290530 $Y=290800
X1859 1 2 102 2 1124 1 sky130_fd_sc_hd__inv_1 $T=297160 301920 1 0 $X=296970 $Y=298960
X1860 1 2 98 2 1146 1 sky130_fd_sc_hd__inv_1 $T=312800 263840 0 0 $X=312610 $Y=263600
X1861 1 2 80 2 1123 1 sky130_fd_sc_hd__inv_1 $T=312800 280160 0 0 $X=312610 $Y=279920
X1862 1 2 94 2 184 1 sky130_fd_sc_hd__inv_1 $T=316940 252960 1 0 $X=316750 $Y=250000
X1863 1 2 106 2 1166 1 sky130_fd_sc_hd__inv_1 $T=322920 307360 0 0 $X=322730 $Y=307120
X1864 1 2 104 2 1183 1 sky130_fd_sc_hd__inv_1 $T=329820 274720 0 0 $X=329630 $Y=274480
X1865 1 2 103 2 1184 1 sky130_fd_sc_hd__inv_1 $T=330280 258400 0 0 $X=330090 $Y=258160
X1866 1 2 99 2 1199 1 sky130_fd_sc_hd__inv_1 $T=338100 285600 1 0 $X=337910 $Y=282640
X1867 1 2 212 2 1203 1 sky130_fd_sc_hd__inv_1 $T=353740 307360 1 0 $X=353550 $Y=304400
X1868 1 2 244 2 247 1 sky130_fd_sc_hd__inv_1 $T=362940 247520 0 0 $X=362750 $Y=247280
X1869 1 2 246 2 1245 1 sky130_fd_sc_hd__inv_1 $T=367080 307360 0 0 $X=366890 $Y=307120
X1870 1 2 242 2 1240 1 sky130_fd_sc_hd__inv_1 $T=379040 269280 1 0 $X=378850 $Y=266320
X1871 1 2 264 2 1253 1 sky130_fd_sc_hd__inv_1 $T=382260 307360 1 0 $X=382070 $Y=304400
X1872 1 2 269 2 1252 1 sky130_fd_sc_hd__inv_1 $T=386860 274720 0 0 $X=386670 $Y=274480
X1873 1 2 278 2 1273 1 sky130_fd_sc_hd__inv_1 $T=398820 247520 0 0 $X=398630 $Y=247280
X1874 1 2 273 2 1299 1 sky130_fd_sc_hd__inv_1 $T=401120 312800 1 0 $X=400930 $Y=309840
X1875 1 2 281 2 1277 1 sky130_fd_sc_hd__inv_1 $T=405260 269280 1 0 $X=405070 $Y=266320
X1876 1 2 294 2 293 1 sky130_fd_sc_hd__inv_1 $T=413540 247520 0 0 $X=413350 $Y=247280
X1877 1 2 297 2 1348 1 sky130_fd_sc_hd__inv_1 $T=416760 269280 0 0 $X=416570 $Y=269040
X1878 1 2 286 2 1312 1 sky130_fd_sc_hd__inv_1 $T=417220 274720 1 0 $X=417030 $Y=271760
X1879 1 2 289 2 1333 1 sky130_fd_sc_hd__inv_1 $T=418600 301920 0 0 $X=418410 $Y=301680
X1880 1 2 300 2 1343 1 sky130_fd_sc_hd__inv_1 $T=426420 258400 1 0 $X=426230 $Y=255440
X1881 1 2 309 2 1370 1 sky130_fd_sc_hd__inv_1 $T=441140 252960 1 0 $X=440950 $Y=250000
X1882 1 2 301 2 1387 1 sky130_fd_sc_hd__inv_1 $T=446660 301920 0 0 $X=446470 $Y=301680
X1883 1 2 313 2 1406 1 sky130_fd_sc_hd__inv_1 $T=451720 269280 1 0 $X=451530 $Y=266320
X1884 1 2 315 2 1420 1 sky130_fd_sc_hd__inv_1 $T=453100 301920 0 0 $X=452910 $Y=301680
X1885 1 2 317 2 1437 1 sky130_fd_sc_hd__inv_1 $T=462300 274720 0 0 $X=462110 $Y=274480
X1886 1 2 322 2 1375 1 sky130_fd_sc_hd__inv_1 $T=466900 263840 1 0 $X=466710 $Y=260880
X1887 1 2 331 2 319 1 sky130_fd_sc_hd__inv_1 $T=469200 247520 1 0 $X=469010 $Y=244560
X1888 1 2 327 2 1467 1 sky130_fd_sc_hd__inv_1 $T=479320 280160 0 0 $X=479130 $Y=279920
X1889 1 2 340 2 1470 1 sky130_fd_sc_hd__inv_1 $T=483000 252960 0 0 $X=482810 $Y=252720
X1890 1 2 329 2 1449 1 sky130_fd_sc_hd__inv_1 $T=483460 296480 1 0 $X=483270 $Y=293520
X1891 1 2 350 2 1484 1 sky130_fd_sc_hd__inv_1 $T=497260 269280 1 0 $X=497070 $Y=266320
X1892 1 2 360 2 1504 1 sky130_fd_sc_hd__inv_1 $T=503700 307360 1 0 $X=503510 $Y=304400
X1893 1 2 242 2 1532 1 sky130_fd_sc_hd__inv_1 $T=505540 285600 1 0 $X=505350 $Y=282640
X1894 1 2 300 2 1534 1 sky130_fd_sc_hd__inv_1 $T=507840 258400 0 0 $X=507650 $Y=258160
X1895 1 2 294 2 1519 1 sky130_fd_sc_hd__inv_1 $T=516580 247520 0 0 $X=516390 $Y=247280
X1896 1 2 297 2 1547 1 sky130_fd_sc_hd__inv_1 $T=524860 269280 0 0 $X=524670 $Y=269040
X1897 1 2 309 2 1576 1 sky130_fd_sc_hd__inv_1 $T=529920 252960 1 0 $X=529730 $Y=250000
X1898 1 2 286 2 1583 1 sky130_fd_sc_hd__inv_1 $T=533140 280160 0 0 $X=532950 $Y=279920
X1899 1 2 212 2 394 1 sky130_fd_sc_hd__inv_1 $T=534980 307360 0 0 $X=534790 $Y=307120
X1900 1 2 281 2 1589 1 sky130_fd_sc_hd__inv_1 $T=539120 269280 1 0 $X=538930 $Y=266320
X1901 1 2 246 2 411 1 sky130_fd_sc_hd__inv_1 $T=553380 312800 1 0 $X=553190 $Y=309840
X1902 1 2 269 2 1620 1 sky130_fd_sc_hd__inv_1 $T=556140 274720 0 0 $X=555950 $Y=274480
X1903 1 2 340 2 1635 1 sky130_fd_sc_hd__inv_1 $T=559820 252960 1 0 $X=559630 $Y=250000
X1904 1 2 322 2 1615 1 sky130_fd_sc_hd__inv_1 $T=567640 263840 1 0 $X=567450 $Y=260880
X1905 1 2 317 2 1650 1 sky130_fd_sc_hd__inv_1 $T=571320 285600 1 0 $X=571130 $Y=282640
X1906 1 2 273 2 1656 1 sky130_fd_sc_hd__inv_1 $T=574540 307360 0 0 $X=574350 $Y=307120
X1907 1 2 414 2 1681 1 sky130_fd_sc_hd__inv_1 $T=582820 274720 0 0 $X=582630 $Y=274480
X1908 1 2 414 2 1685 1 sky130_fd_sc_hd__inv_1 $T=583740 280160 0 0 $X=583550 $Y=279920
X1909 1 2 420 2 1688 1 sky130_fd_sc_hd__inv_1 $T=594780 263840 1 0 $X=594590 $Y=260880
X1910 1 2 254 2 1701 1 sky130_fd_sc_hd__inv_1 $T=595240 301920 0 0 $X=595050 $Y=301680
X1911 1 2 342 2 1739 1 sky130_fd_sc_hd__inv_1 $T=610420 291040 1 0 $X=610230 $Y=288080
X1912 1 2 431 2 1723 1 sky130_fd_sc_hd__inv_1 $T=615480 274720 0 0 $X=615290 $Y=274480
X1913 1 2 301 2 1747 1 sky130_fd_sc_hd__inv_1 $T=615940 307360 1 0 $X=615750 $Y=304400
X1914 1 2 436 2 435 1 sky130_fd_sc_hd__inv_1 $T=627440 252960 1 0 $X=627250 $Y=250000
X1915 1 2 428 2 1730 1 sky130_fd_sc_hd__inv_1 $T=628820 263840 1 0 $X=628630 $Y=260880
X1916 1 2 433 2 1761 1 sky130_fd_sc_hd__inv_1 $T=635260 274720 1 0 $X=635070 $Y=271760
X1917 1 2 442 2 1802 1 sky130_fd_sc_hd__inv_1 $T=647680 263840 0 0 $X=647490 $Y=263600
X1918 1 2 315 2 1824 1 sky130_fd_sc_hd__inv_1 $T=656420 307360 1 0 $X=656230 $Y=304400
X1919 1 2 447 2 444 1 sky130_fd_sc_hd__inv_1 $T=657340 247520 1 0 $X=657150 $Y=244560
X1920 1 2 443 2 1813 1 sky130_fd_sc_hd__inv_1 $T=658720 280160 0 0 $X=658530 $Y=279920
X1921 1 2 439 2 1812 1 sky130_fd_sc_hd__inv_1 $T=662860 252960 1 0 $X=662670 $Y=250000
X1922 1 2 327 2 1804 1 sky130_fd_sc_hd__inv_1 $T=663780 285600 0 0 $X=663590 $Y=285360
X1923 1 2 350 2 1844 1 sky130_fd_sc_hd__inv_1 $T=665620 274720 1 0 $X=665430 $Y=271760
X1924 1 2 433 2 1866 1 sky130_fd_sc_hd__inv_1 $T=672980 285600 1 0 $X=672790 $Y=282640
X1925 1 2 313 2 1853 1 sky130_fd_sc_hd__inv_1 $T=675280 258400 0 0 $X=675090 $Y=258160
X1926 1 2 360 2 1875 1 sky130_fd_sc_hd__inv_1 $T=676660 307360 1 0 $X=676470 $Y=304400
X1927 1 2 449 2 1859 1 sky130_fd_sc_hd__inv_1 $T=678500 247520 1 0 $X=678310 $Y=244560
X1928 1 2 420 2 1910 1 sky130_fd_sc_hd__inv_1 $T=694140 269280 0 0 $X=693950 $Y=269040
X1929 1 2 431 2 1904 1 sky130_fd_sc_hd__inv_1 $T=694140 280160 0 0 $X=693950 $Y=279920
X1930 1 2 436 2 1916 1 sky130_fd_sc_hd__inv_1 $T=700120 247520 0 0 $X=699930 $Y=247280
X1931 1 2 329 2 1926 1 sky130_fd_sc_hd__inv_1 $T=704720 301920 0 0 $X=704530 $Y=301680
X1932 1 2 443 2 1950 1 sky130_fd_sc_hd__inv_1 $T=717140 285600 1 0 $X=716950 $Y=282640
X1933 1 2 428 2 1955 1 sky130_fd_sc_hd__inv_1 $T=719900 263840 1 0 $X=719710 $Y=260880
X1934 1 2 442 2 1965 1 sky130_fd_sc_hd__inv_1 $T=723580 274720 0 0 $X=723390 $Y=274480
X1935 1 2 439 2 462 1 sky130_fd_sc_hd__inv_1 $T=726340 252960 0 0 $X=726150 $Y=252720
X1936 1 2 ICV_25 $T=44620 252960 1 0 $X=44430 $Y=250000
X1937 1 2 ICV_25 $T=72680 291040 1 0 $X=72490 $Y=288080
X1938 1 2 ICV_25 $T=100740 301920 1 0 $X=100550 $Y=298960
X1939 1 2 ICV_25 $T=114540 258400 0 0 $X=114350 $Y=258160
X1940 1 2 ICV_25 $T=156860 247520 1 0 $X=156670 $Y=244560
X1941 1 2 ICV_25 $T=282900 258400 0 0 $X=282710 $Y=258160
X1942 1 2 ICV_25 $T=451260 263840 0 0 $X=451070 $Y=263600
X1943 1 2 ICV_25 $T=465520 269280 1 0 $X=465330 $Y=266320
X1944 1 2 ICV_25 $T=507380 269280 0 0 $X=507190 $Y=269040
X1945 1 2 ICV_25 $T=535440 296480 0 0 $X=535250 $Y=296240
X1946 1 2 ICV_25 $T=563500 263840 0 0 $X=563310 $Y=263600
X1947 1 2 ICV_25 $T=577760 312800 1 0 $X=577570 $Y=309840
X1948 1 2 ICV_25 $T=591560 247520 0 0 $X=591370 $Y=247280
X1949 1 2 ICV_25 $T=619620 307360 0 0 $X=619430 $Y=307120
X1950 1 2 ICV_25 $T=633880 307360 1 0 $X=633690 $Y=304400
X1951 1 2 ICV_25 $T=661940 274720 1 0 $X=661750 $Y=271760
X1952 1 2 ICV_25 $T=675740 269280 0 0 $X=675550 $Y=269040
X1953 1 2 ICV_25 $T=731860 301920 0 0 $X=731670 $Y=301680
X1954 1 2 577 578 13 ICV_26 $T=29900 274720 1 0 $X=29710 $Y=271760
X1955 1 2 587 578 18 ICV_26 $T=40480 258400 1 0 $X=40290 $Y=255440
X1956 1 2 589 578 34 ICV_26 $T=40940 263840 1 0 $X=40750 $Y=260880
X1957 1 2 607 45 17 ICV_26 $T=49220 247520 0 0 $X=49030 $Y=247280
X1958 1 2 625 627 13 ICV_26 $T=57040 263840 0 0 $X=56850 $Y=263600
X1959 1 2 649 642 30 ICV_26 $T=67160 296480 1 0 $X=66970 $Y=293520
X1960 1 2 687 690 19 ICV_26 $T=86940 258400 1 0 $X=86750 $Y=255440
X1961 1 2 85 77 16 ICV_26 $T=106720 307360 0 0 $X=106530 $Y=307120
X1962 1 2 799 771 30 ICV_26 $T=141220 247520 0 0 $X=141030 $Y=247280
X1963 1 2 832 835 30 ICV_26 $T=155020 258400 1 0 $X=154830 $Y=255440
X1964 1 2 868 863 122 ICV_26 $T=174340 258400 0 0 $X=174150 $Y=258160
X1965 1 2 869 873 123 ICV_26 $T=174340 296480 0 0 $X=174150 $Y=296240
X1966 1 2 870 119 121 ICV_26 $T=174340 301920 0 0 $X=174150 $Y=301680
X1967 1 2 865 873 121 ICV_26 $T=174800 296480 1 0 $X=174610 $Y=293520
X1968 1 2 884 863 123 ICV_26 $T=183540 263840 1 0 $X=183350 $Y=260880
X1969 1 2 1011 973 135 ICV_26 $T=241960 274720 0 0 $X=241770 $Y=274480
X1970 1 2 158 159 131 ICV_26 $T=253460 247520 0 0 $X=253270 $Y=247280
X1971 1 2 1057 1027 134 ICV_26 $T=265880 269280 0 0 $X=265690 $Y=269040
X1972 1 2 1071 168 122 ICV_26 $T=272780 307360 1 0 $X=272590 $Y=304400
X1973 1 2 1073 1053 134 ICV_26 $T=275540 258400 1 0 $X=275350 $Y=255440
X1974 1 2 1074 1027 123 ICV_26 $T=277840 269280 0 0 $X=277650 $Y=269040
X1975 1 2 1103 172 134 ICV_26 $T=288420 312800 1 0 $X=288230 $Y=309840
X1976 1 2 1114 1104 131 ICV_26 $T=293020 274720 0 0 $X=292830 $Y=274480
X1977 1 2 1132 159 134 ICV_26 $T=300840 247520 1 0 $X=300650 $Y=244560
X1978 1 2 1197 1199 135 ICV_26 $T=336260 296480 1 0 $X=336070 $Y=293520
X1979 1 2 1213 1203 180 ICV_26 $T=349140 307360 1 0 $X=348950 $Y=304400
X1980 1 2 1285 1252 262 ICV_26 $T=385020 274720 1 0 $X=384830 $Y=271760
X1981 1 2 1327 293 260 ICV_26 $T=407560 247520 0 0 $X=407370 $Y=247280
X1982 1 2 1354 1348 233 ICV_26 $T=421360 285600 1 0 $X=421170 $Y=282640
X1983 1 2 1423 1420 186 ICV_26 $T=454940 291040 0 0 $X=454750 $Y=290800
X1984 1 2 1460 334 185 ICV_26 $T=470120 301920 0 0 $X=469930 $Y=301680
X1985 1 2 1487 343 260 ICV_26 $T=483000 247520 0 0 $X=482810 $Y=247280
X1986 1 2 1563 369 306 ICV_26 $T=525320 247520 0 0 $X=525130 $Y=247280
X1987 1 2 1582 1583 306 ICV_26 $T=532680 285600 0 0 $X=532490 $Y=285360
X1988 1 2 1621 1620 328 ICV_26 $T=553840 285600 0 0 $X=553650 $Y=285360
X1989 1 2 1727 1730 229 ICV_26 $T=604440 269280 1 0 $X=604250 $Y=266320
X1990 1 2 1786 440 400 ICV_26 $T=632500 312800 1 0 $X=632310 $Y=309840
X1991 1 2 1836 1824 376 ICV_26 $T=657800 307360 1 0 $X=657610 $Y=304400
X1992 1 2 1842 1824 400 ICV_26 $T=659640 296480 0 0 $X=659450 $Y=296240
X1993 1 2 1872 1853 341 ICV_26 $T=674360 263840 0 0 $X=674170 $Y=263600
X1994 1 2 1911 1875 361 ICV_26 $T=693680 301920 1 0 $X=693490 $Y=298960
X1995 1 2 1956 463 341 ICV_26 $T=721740 247520 1 0 $X=721550 $Y=244560
X1996 1 2 523 11 556 ICV_28 $T=10580 247520 1 0 $X=10390 $Y=244560
X1997 1 2 21 5 43 ICV_28 $T=31740 312800 1 0 $X=31550 $Y=309840
X1998 1 2 619 24 637 ICV_28 $T=53820 252960 1 0 $X=53630 $Y=250000
X1999 1 2 618 24 668 ICV_28 $T=69460 291040 0 0 $X=69270 $Y=290800
X2000 1 2 665 10 700 ICV_28 $T=84180 291040 1 0 $X=83990 $Y=288080
X2001 1 2 810 14 842 ICV_28 $T=153640 296480 0 0 $X=153450 $Y=296240
X2002 1 2 899 126 924 ICV_28 $T=191360 280160 0 0 $X=191170 $Y=279920
X2003 1 2 1070 128 1087 ICV_28 $T=272780 291040 1 0 $X=272590 $Y=288080
X2004 1 2 176 125 1177 ICV_28 $T=318320 252960 1 0 $X=318130 $Y=250000
X2005 1 2 1180 112 1198 ICV_28 $T=328900 285600 1 0 $X=328710 $Y=282640
X2006 1 2 1247 227 1289 ICV_28 $T=379500 280160 0 0 $X=379310 $Y=279920
X2007 1 2 326 218 1489 ICV_28 $T=476560 312800 1 0 $X=476370 $Y=309840
X2008 1 2 1483 224 1494 ICV_28 $T=480700 280160 1 0 $X=480510 $Y=277200
X2009 1 2 1491 213 1502 ICV_28 $T=484840 296480 1 0 $X=484650 $Y=293520
X2010 1 2 1515 364 1545 ICV_28 $T=505080 269280 1 0 $X=504890 $Y=266320
X2011 1 2 409 401 1643 ICV_28 $T=554760 312800 1 0 $X=554570 $Y=309840
X2012 1 2 1617 358 1646 ICV_28 $T=560740 269280 1 0 $X=560550 $Y=266320
X2013 1 2 1659 253 1673 ICV_28 $T=571780 274720 1 0 $X=571590 $Y=271760
X2014 1 2 618 14 633 ICV_29 $T=51980 291040 0 0 $X=51790 $Y=290800
X2015 1 2 619 26 657 ICV_29 $T=63940 247520 1 0 $X=63750 $Y=244560
X2016 1 2 664 14 691 ICV_29 $T=79120 269280 0 0 $X=78930 $Y=269040
X2017 1 2 664 24 699 ICV_29 $T=83720 274720 1 0 $X=83530 $Y=271760
X2018 1 2 761 26 774 ICV_29 $T=118220 280160 0 0 $X=118030 $Y=279920
X2019 1 2 861 108 876 ICV_29 $T=168820 269280 1 0 $X=168630 $Y=266320
X2020 1 2 919 108 918 ICV_29 $T=195960 274720 1 0 $X=195770 $Y=271760
X2021 1 2 170 108 1126 ICV_29 $T=290720 247520 1 0 $X=290530 $Y=244560
X2022 1 2 1116 108 1131 ICV_29 $T=292100 291040 0 0 $X=291910 $Y=290800
X2023 1 2 1129 108 1148 ICV_29 $T=300840 258400 1 0 $X=300650 $Y=255440
X2024 1 2 1176 127 1186 ICV_29 $T=323840 252960 0 0 $X=323650 $Y=252720
X2025 1 2 1258 213 1250 ICV_29 $T=370760 296480 0 0 $X=370570 $Y=296240
X2026 1 2 1290 224 1307 ICV_29 $T=388240 274720 0 0 $X=388050 $Y=274480
X2027 1 2 1459 251 1476 ICV_29 $T=469200 263840 1 0 $X=469010 $Y=260880
X2028 1 2 1574 368 1585 ICV_29 $T=526240 269280 0 0 $X=526050 $Y=269040
X2029 1 2 379 401 406 ICV_29 $T=532680 312800 1 0 $X=532490 $Y=309840
X2030 1 2 1601 368 1619 ICV_29 $T=543260 296480 1 0 $X=543070 $Y=293520
X2031 1 2 1617 368 1653 ICV_29 $T=562120 274720 1 0 $X=561930 $Y=271760
X2032 1 2 1618 359 1661 ICV_29 $T=564880 258400 1 0 $X=564690 $Y=255440
X2033 1 2 412 223 1684 ICV_29 $T=574540 247520 0 0 $X=574350 $Y=247280
X2034 1 2 1820 401 1842 ICV_29 $T=651360 301920 0 0 $X=651170 $Y=301680
X2035 1 2 1820 407 1855 ICV_29 $T=659640 307360 0 0 $X=659450 $Y=307120
X2036 1 2 1893 367 1936 ICV_29 $T=700120 269280 1 0 $X=699930 $Y=266320
X2037 1 2 550 542 18 541 542 13 ICV_30 $T=17020 258400 0 0 $X=16830 $Y=258160
X2038 1 2 552 555 16 554 555 18 ICV_30 $T=21620 285600 0 0 $X=21430 $Y=285360
X2039 1 2 39 29 13 588 29 34 ICV_30 $T=35880 301920 0 0 $X=35690 $Y=301680
X2040 1 2 584 585 13 601 585 18 ICV_30 $T=38180 301920 1 0 $X=37990 $Y=298960
X2041 1 2 616 602 13 623 585 19 ICV_30 $T=52440 285600 0 0 $X=52250 $Y=285360
X2042 1 2 636 641 33 646 641 19 ICV_30 $T=62100 269280 0 0 $X=61910 $Y=269040
X2043 1 2 634 642 16 633 642 19 ICV_30 $T=62100 296480 0 0 $X=61910 $Y=296240
X2044 1 2 630 641 34 656 641 18 ICV_30 $T=67160 285600 1 0 $X=66970 $Y=282640
X2045 1 2 648 627 34 647 627 18 ICV_30 $T=67620 258400 1 0 $X=67430 $Y=255440
X2046 1 2 659 66 17 660 66 19 ICV_30 $T=74060 301920 0 0 $X=73870 $Y=301680
X2047 1 2 657 56 34 666 56 16 ICV_30 $T=76360 247520 1 0 $X=76170 $Y=244560
X2048 1 2 68 69 19 689 690 18 ICV_30 $T=84640 247520 1 0 $X=84450 $Y=244560
X2049 1 2 678 684 19 696 684 17 ICV_30 $T=87860 280160 1 0 $X=87670 $Y=277200
X2050 1 2 697 693 30 713 693 17 ICV_30 $T=92460 301920 1 0 $X=92270 $Y=298960
X2051 1 2 699 676 33 691 676 19 ICV_30 $T=92920 269280 0 0 $X=92730 $Y=269040
X2052 1 2 706 74 13 717 718 18 ICV_30 $T=95680 263840 1 0 $X=95490 $Y=260880
X2053 1 2 705 77 19 722 693 13 ICV_30 $T=98440 307360 0 0 $X=98250 $Y=307120
X2054 1 2 81 78 13 720 690 34 ICV_30 $T=101660 247520 0 0 $X=101470 $Y=247280
X2055 1 2 723 730 13 731 740 34 ICV_30 $T=105800 280160 1 0 $X=105610 $Y=277200
X2056 1 2 733 730 16 734 730 18 ICV_30 $T=107640 263840 0 0 $X=107450 $Y=263600
X2057 1 2 735 730 33 724 740 13 ICV_30 $T=109020 269280 0 0 $X=108830 $Y=269040
X2058 1 2 91 74 33 762 718 19 ICV_30 $T=117760 247520 1 0 $X=117570 $Y=244560
X2059 1 2 736 730 17 759 718 33 ICV_30 $T=118220 258400 0 0 $X=118030 $Y=258160
X2060 1 2 777 779 33 776 779 30 ICV_30 $T=128340 280160 0 0 $X=128150 $Y=279920
X2061 1 2 794 96 17 782 96 13 ICV_30 $T=146280 307360 0 0 $X=146090 $Y=307120
X2062 1 2 814 89 30 826 824 34 ICV_30 $T=148580 301920 1 0 $X=148390 $Y=298960
X2063 1 2 831 835 34 834 835 18 ICV_30 $T=160540 247520 1 0 $X=160350 $Y=244560
X2064 1 2 838 811 19 780 718 13 ICV_30 $T=160540 269280 1 0 $X=160350 $Y=266320
X2065 1 2 846 822 33 845 822 19 ICV_30 $T=162840 274720 1 0 $X=162650 $Y=271760
X2066 1 2 864 874 121 877 862 117 ICV_30 $T=175260 274720 0 0 $X=175070 $Y=274480
X2067 1 2 904 862 135 903 862 131 ICV_30 $T=192280 280160 1 0 $X=192090 $Y=277200
X2068 1 2 892 874 134 929 921 117 ICV_30 $T=200560 280160 1 0 $X=200370 $Y=277200
X2069 1 2 893 874 135 897 874 131 ICV_30 $T=202400 280160 0 0 $X=202210 $Y=279920
X2070 1 2 941 144 117 843 89 19 ICV_30 $T=214360 301920 0 0 $X=214170 $Y=301680
X2071 1 2 948 146 135 946 933 131 ICV_30 $T=214820 252960 0 0 $X=214630 $Y=252720
X2072 1 2 949 921 131 922 923 121 ICV_30 $T=217580 280160 0 0 $X=217390 $Y=279920
X2073 1 2 1009 986 117 1016 986 136 ICV_30 $T=241500 263840 0 0 $X=241310 $Y=263600
X2074 1 2 1014 975 122 1018 975 123 ICV_30 $T=244260 296480 0 0 $X=244070 $Y=296240
X2075 1 2 1044 1027 135 1040 1027 131 ICV_30 $T=263580 263840 1 0 $X=263390 $Y=260880
X2076 1 2 1051 1032 131 955 139 117 ICV_30 $T=264040 307360 1 0 $X=263850 $Y=304400
X2077 1 2 1065 1032 123 1066 1032 117 ICV_30 $T=270020 296480 0 0 $X=269830 $Y=296240
X2078 1 2 1092 1053 117 1100 1053 135 ICV_30 $T=283360 258400 1 0 $X=283170 $Y=255440
X2079 1 2 1102 1086 134 1113 1086 122 ICV_30 $T=288880 307360 1 0 $X=288690 $Y=304400
X2080 1 2 1138 1104 136 1139 1104 135 ICV_30 $T=304520 269280 0 0 $X=304330 $Y=269040
X2081 1 2 1153 1124 117 1158 189 123 ICV_30 $T=314640 307360 0 0 $X=314450 $Y=307120
X2082 1 2 1156 184 117 1162 1146 117 ICV_30 $T=315560 252960 0 0 $X=315370 $Y=252720
X2083 1 2 1170 1123 121 1181 1183 135 ICV_30 $T=323840 269280 0 0 $X=323650 $Y=269040
X2084 1 2 1186 1184 134 1193 1184 117 ICV_30 $T=332580 258400 0 0 $X=332390 $Y=258160
X2085 1 2 1187 1166 134 1194 1166 135 ICV_30 $T=333500 301920 0 0 $X=333310 $Y=301680
X2086 1 2 1208 1184 136 1209 1184 131 ICV_30 $T=343160 258400 0 0 $X=342970 $Y=258160
X2087 1 2 1205 1184 121 230 231 233 ICV_30 $T=344540 252960 1 0 $X=344350 $Y=250000
X2088 1 2 1223 247 252 1228 247 257 ICV_30 $T=356960 252960 1 0 $X=356770 $Y=250000
X2089 1 2 1255 1240 262 1265 1240 233 ICV_30 $T=370760 263840 0 0 $X=370570 $Y=263600
X2090 1 2 1271 1253 202 1278 1253 192 ICV_30 $T=380880 296480 0 0 $X=380690 $Y=296240
X2091 1 2 1275 1253 186 1288 1253 199 ICV_30 $T=385020 296480 1 0 $X=384830 $Y=293520
X2092 1 2 1286 1277 262 1297 1277 252 ICV_30 $T=387320 263840 0 0 $X=387130 $Y=263600
X2093 1 2 1289 1252 252 1298 1252 257 ICV_30 $T=387320 291040 1 0 $X=387130 $Y=288080
X2094 1 2 1313 1277 260 1320 1277 263 ICV_30 $T=400200 263840 1 0 $X=400010 $Y=260880
X2095 1 2 1301 1312 263 1329 1312 201 ICV_30 $T=407560 269280 0 0 $X=407370 $Y=269040
X2096 1 2 1314 1299 199 1346 1333 192 ICV_30 $T=413080 296480 1 0 $X=412890 $Y=293520
X2097 1 2 1366 1370 260 1368 1370 229 ICV_30 $T=426880 252960 0 0 $X=426690 $Y=252720
X2098 1 2 1364 1348 263 1377 1348 229 ICV_30 $T=426880 274720 0 0 $X=426690 $Y=274480
X2099 1 2 1362 1333 180 1352 1333 188 ICV_30 $T=426880 296480 0 0 $X=426690 $Y=296240
X2100 1 2 1397 1375 229 1411 1375 257 ICV_30 $T=441140 247520 1 0 $X=440950 $Y=244560
X2101 1 2 1386 1387 178 1347 1333 185 ICV_30 $T=441140 301920 1 0 $X=440950 $Y=298960
X2102 1 2 1404 1370 262 1393 1370 263 ICV_30 $T=442520 252960 1 0 $X=442330 $Y=250000
X2103 1 2 1405 1406 262 1395 1406 229 ICV_30 $T=443440 274720 1 0 $X=443250 $Y=271760
X2104 1 2 1416 1375 252 1426 1375 233 ICV_30 $T=451260 263840 1 0 $X=451070 $Y=260880
X2105 1 2 1425 1420 180 1439 1420 188 ICV_30 $T=456320 307360 1 0 $X=456130 $Y=304400
X2106 1 2 1430 1420 185 324 318 199 ICV_30 $T=457240 307360 0 0 $X=457050 $Y=307120
X2107 1 2 1436 1437 233 1434 1437 257 ICV_30 $T=459540 285600 1 0 $X=459350 $Y=282640
X2108 1 2 1451 1437 229 1447 1375 263 ICV_30 $T=469200 274720 1 0 $X=469010 $Y=271760
X2109 1 2 1479 1484 201 1490 1484 263 ICV_30 $T=481160 274720 1 0 $X=480970 $Y=271760
X2110 1 2 1548 1532 303 1555 1532 306 ICV_30 $T=513820 285600 0 0 $X=513630 $Y=285360
X2111 1 2 1565 1534 303 1571 1534 306 ICV_30 $T=525320 263840 1 0 $X=525130 $Y=260880
X2112 1 2 1567 1547 348 1559 1547 382 ICV_30 $T=525320 280160 1 0 $X=525130 $Y=277200
X2113 1 2 1578 1583 337 1590 1583 348 ICV_30 $T=534980 296480 1 0 $X=534790 $Y=293520
X2114 1 2 1595 1583 303 1600 1583 372 ICV_30 $T=540500 291040 1 0 $X=540310 $Y=288080
X2115 1 2 1619 1620 382 1626 1620 372 ICV_30 $T=552000 296480 0 0 $X=551810 $Y=296240
X2116 1 2 1625 1620 306 1622 1620 337 ICV_30 $T=554760 291040 1 0 $X=554570 $Y=288080
X2117 1 2 1642 411 361 1643 411 400 ICV_30 $T=562580 307360 1 0 $X=562390 $Y=304400
X2118 1 2 1644 1635 348 1631 403 372 ICV_30 $T=563500 252960 1 0 $X=563310 $Y=250000
X2119 1 2 1648 1650 303 1649 1650 341 ICV_30 $T=569940 280160 1 0 $X=569750 $Y=277200
X2120 1 2 1654 1656 361 1658 1656 376 ICV_30 $T=571780 307360 1 0 $X=571590 $Y=304400
X2121 1 2 1651 1650 306 1645 1650 337 ICV_30 $T=572240 291040 1 0 $X=572050 $Y=288080
X2122 1 2 1652 1650 348 1665 1650 372 ICV_30 $T=572240 296480 1 0 $X=572050 $Y=293520
X2123 1 2 1657 1615 303 1662 1615 341 ICV_30 $T=572700 269280 1 0 $X=572510 $Y=266320
X2124 1 2 1676 1681 252 1674 1681 257 ICV_30 $T=581440 280160 1 0 $X=581250 $Y=277200
X2125 1 2 1678 415 229 1686 1688 257 ICV_30 $T=581900 263840 1 0 $X=581710 $Y=260880
X2126 1 2 421 415 262 1684 415 260 ICV_30 $T=584200 247520 1 0 $X=584010 $Y=244560
X2127 1 2 1687 423 201 1698 1688 229 ICV_30 $T=586500 252960 0 0 $X=586310 $Y=252720
X2128 1 2 1704 423 257 425 423 252 ICV_30 $T=592480 247520 1 0 $X=592290 $Y=244560
X2129 1 2 1702 1681 233 1705 1681 260 ICV_30 $T=595240 280160 0 0 $X=595050 $Y=279920
X2130 1 2 1776 1761 252 1772 1761 233 ICV_30 $T=631120 280160 0 0 $X=630930 $Y=279920
X2131 1 2 1794 444 229 1808 1812 229 ICV_30 $T=642620 247520 0 0 $X=642430 $Y=247280
X2132 1 2 1817 1813 233 1821 1813 260 ICV_30 $T=651820 285600 1 0 $X=651630 $Y=282640
X2133 1 2 1855 1824 375 1865 1824 373 ICV_30 $T=668380 307360 1 0 $X=668190 $Y=304400
X2134 1 2 1856 1859 382 1870 1853 303 ICV_30 $T=670680 258400 1 0 $X=670490 $Y=255440
X2135 1 2 1860 1866 306 1863 1866 382 ICV_30 $T=672060 291040 1 0 $X=671870 $Y=288080
X2136 1 2 1877 1875 373 1885 1875 375 ICV_30 $T=678040 307360 1 0 $X=677850 $Y=304400
X2137 1 2 1907 1910 303 1906 1910 341 ICV_30 $T=693680 274720 1 0 $X=693490 $Y=271760
X2138 1 2 451 454 382 1918 1916 306 ICV_30 $T=695980 252960 1 0 $X=695790 $Y=250000
X2139 1 2 1923 1904 303 1930 1910 337 ICV_30 $T=703340 280160 1 0 $X=703150 $Y=277200
X2140 1 2 1929 453 306 1935 1916 328 ICV_30 $T=707480 252960 1 0 $X=707290 $Y=250000
X2141 1 2 1954 1965 348 1969 1955 348 ICV_30 $T=721740 274720 1 0 $X=721550 $Y=271760
X2142 1 2 1952 1965 306 1970 1965 372 ICV_30 $T=721740 285600 1 0 $X=721550 $Y=282640
X2143 1 2 1963 1926 389 1962 1926 400 ICV_30 $T=721740 301920 1 0 $X=721550 $Y=298960
X2144 1 2 3 7 2 529 1 sky130_fd_sc_hd__and2_1 $T=7360 285600 1 0 $X=7170 $Y=282640
X2145 1 2 6 7 2 12 1 sky130_fd_sc_hd__and2_1 $T=8280 247520 1 0 $X=8090 $Y=244560
X2146 1 2 8 7 2 531 1 sky130_fd_sc_hd__and2_1 $T=8280 291040 1 0 $X=8090 $Y=288080
X2147 1 2 15 7 2 528 1 sky130_fd_sc_hd__and2_1 $T=13800 258400 0 0 $X=13610 $Y=258160
X2148 1 2 20 7 2 551 1 sky130_fd_sc_hd__and2_1 $T=20240 274720 1 0 $X=20050 $Y=271760
X2149 1 2 28 7 2 31 1 sky130_fd_sc_hd__and2_1 $T=28520 247520 1 0 $X=28330 $Y=244560
X2150 1 2 35 7 2 580 1 sky130_fd_sc_hd__and2_1 $T=31280 285600 0 0 $X=31090 $Y=285360
X2151 1 2 49 7 2 604 1 sky130_fd_sc_hd__and2_1 $T=45540 263840 1 0 $X=45350 $Y=260880
X2152 1 2 48 7 2 605 1 sky130_fd_sc_hd__and2_1 $T=45540 269280 1 0 $X=45350 $Y=266320
X2153 1 2 57 7 2 639 1 sky130_fd_sc_hd__and2_1 $T=62100 291040 1 0 $X=61910 $Y=288080
X2154 1 2 60 7 2 643 1 sky130_fd_sc_hd__and2_1 $T=63020 252960 1 0 $X=62830 $Y=250000
X2155 1 2 63 7 2 653 1 sky130_fd_sc_hd__and2_1 $T=70380 296480 0 0 $X=70190 $Y=296240
X2156 1 2 64 7 2 661 1 sky130_fd_sc_hd__and2_1 $T=73600 274720 1 0 $X=73410 $Y=271760
X2157 1 2 67 7 2 680 1 sky130_fd_sc_hd__and2_1 $T=81880 291040 1 0 $X=81690 $Y=288080
X2158 1 2 73 7 2 702 1 sky130_fd_sc_hd__and2_1 $T=93380 307360 1 0 $X=93190 $Y=304400
X2159 1 2 76 7 2 714 1 sky130_fd_sc_hd__and2_1 $T=97520 280160 0 0 $X=97330 $Y=279920
X2160 1 2 80 7 2 709 1 sky130_fd_sc_hd__and2_1 $T=101200 291040 1 0 $X=101010 $Y=288080
X2161 1 2 83 7 2 732 1 sky130_fd_sc_hd__and2_1 $T=106260 252960 0 0 $X=106070 $Y=252720
X2162 1 2 86 7 2 728 1 sky130_fd_sc_hd__and2_1 $T=107640 301920 0 0 $X=107450 $Y=301680
X2163 1 2 88 7 2 750 1 sky130_fd_sc_hd__and2_1 $T=114540 296480 0 0 $X=114350 $Y=296240
X2164 1 2 90 7 2 751 1 sky130_fd_sc_hd__and2_1 $T=115000 274720 0 0 $X=114810 $Y=274480
X2165 1 2 94 7 2 763 1 sky130_fd_sc_hd__and2_1 $T=124200 252960 0 0 $X=124010 $Y=252720
X2166 1 2 98 7 2 785 1 sky130_fd_sc_hd__and2_1 $T=132480 269280 0 0 $X=132290 $Y=269040
X2167 1 2 99 7 2 788 1 sky130_fd_sc_hd__and2_1 $T=136160 285600 0 0 $X=135970 $Y=285360
X2168 1 2 102 7 2 807 1 sky130_fd_sc_hd__and2_1 $T=143520 296480 0 0 $X=143330 $Y=296240
X2169 1 2 103 7 2 816 1 sky130_fd_sc_hd__and2_1 $T=150420 258400 0 0 $X=150230 $Y=258160
X2170 1 2 104 7 2 817 1 sky130_fd_sc_hd__and2_1 $T=154100 280160 0 0 $X=153910 $Y=279920
X2171 1 2 106 7 2 821 1 sky130_fd_sc_hd__and2_1 $T=156860 307360 1 0 $X=156670 $Y=304400
X2172 1 2 3 107 2 849 1 sky130_fd_sc_hd__and2_1 $T=164220 280160 0 0 $X=164030 $Y=279920
X2173 1 2 48 107 2 858 1 sky130_fd_sc_hd__and2_1 $T=166060 263840 1 0 $X=165870 $Y=260880
X2174 1 2 36 107 2 855 1 sky130_fd_sc_hd__and2_1 $T=166060 301920 1 0 $X=165870 $Y=298960
X2175 1 2 15 107 2 860 1 sky130_fd_sc_hd__and2_1 $T=172040 258400 1 0 $X=171850 $Y=255440
X2176 1 2 53 107 2 900 1 sky130_fd_sc_hd__and2_1 $T=192740 252960 1 0 $X=192550 $Y=250000
X2177 1 2 8 107 2 905 1 sky130_fd_sc_hd__and2_1 $T=198260 291040 0 0 $X=198070 $Y=290800
X2178 1 2 49 107 2 914 1 sky130_fd_sc_hd__and2_1 $T=202400 263840 0 0 $X=202210 $Y=263600
X2179 1 2 35 107 2 947 1 sky130_fd_sc_hd__and2_1 $T=212520 291040 1 0 $X=212330 $Y=288080
X2180 1 2 149 107 2 152 1 sky130_fd_sc_hd__and2_1 $T=213900 312800 1 0 $X=213710 $Y=309840
X2181 1 2 64 107 2 953 1 sky130_fd_sc_hd__and2_1 $T=218500 269280 0 0 $X=218310 $Y=269040
X2182 1 2 58 107 2 980 1 sky130_fd_sc_hd__and2_1 $T=226780 301920 0 0 $X=226590 $Y=301680
X2183 1 2 60 107 2 976 1 sky130_fd_sc_hd__and2_1 $T=230460 252960 0 0 $X=230270 $Y=252720
X2184 1 2 76 107 2 984 1 sky130_fd_sc_hd__and2_1 $T=230460 263840 0 0 $X=230270 $Y=263600
X2185 1 2 40 107 2 985 1 sky130_fd_sc_hd__and2_1 $T=241960 285600 1 0 $X=241770 $Y=282640
X2186 1 2 90 107 2 1017 1 sky130_fd_sc_hd__and2_1 $T=248860 269280 1 0 $X=248670 $Y=266320
X2187 1 2 86 107 2 1028 1 sky130_fd_sc_hd__and2_1 $T=255300 301920 0 0 $X=255110 $Y=301680
X2188 1 2 63 107 2 1041 1 sky130_fd_sc_hd__and2_1 $T=258520 285600 0 0 $X=258330 $Y=285360
X2189 1 2 88 107 2 1095 1 sky130_fd_sc_hd__and2_1 $T=282440 291040 1 0 $X=282250 $Y=288080
X2190 1 2 67 107 2 1098 1 sky130_fd_sc_hd__and2_1 $T=284740 280160 1 0 $X=284550 $Y=277200
X2191 1 2 83 107 2 1094 1 sky130_fd_sc_hd__and2_1 $T=286580 252960 0 0 $X=286390 $Y=252720
X2192 1 2 102 107 2 1101 1 sky130_fd_sc_hd__and2_1 $T=286580 307360 1 0 $X=286390 $Y=304400
X2193 1 2 80 107 2 1136 1 sky130_fd_sc_hd__and2_1 $T=304980 280160 1 0 $X=304790 $Y=277200
X2194 1 2 94 107 2 1135 1 sky130_fd_sc_hd__and2_1 $T=305900 252960 0 0 $X=305710 $Y=252720
X2195 1 2 106 107 2 1160 1 sky130_fd_sc_hd__and2_1 $T=316020 301920 0 0 $X=315830 $Y=301680
X2196 1 2 103 107 2 1167 1 sky130_fd_sc_hd__and2_1 $T=324760 258400 1 0 $X=324570 $Y=255440
X2197 1 2 104 107 2 1178 1 sky130_fd_sc_hd__and2_1 $T=325680 280160 1 0 $X=325490 $Y=277200
X2198 1 2 99 107 2 1168 1 sky130_fd_sc_hd__and2_1 $T=325680 291040 1 0 $X=325490 $Y=288080
X2199 1 2 212 207 2 1200 1 sky130_fd_sc_hd__and2_1 $T=342700 301920 0 0 $X=342510 $Y=301680
X2200 1 2 242 215 2 1226 1 sky130_fd_sc_hd__and2_1 $T=356960 263840 1 0 $X=356770 $Y=260880
X2201 1 2 246 207 2 1227 1 sky130_fd_sc_hd__and2_1 $T=356960 307360 1 0 $X=356770 $Y=304400
X2202 1 2 244 215 2 1232 1 sky130_fd_sc_hd__and2_1 $T=357420 247520 1 0 $X=357230 $Y=244560
X2203 1 2 254 207 2 255 1 sky130_fd_sc_hd__and2_1 $T=362020 312800 1 0 $X=361830 $Y=309840
X2204 1 2 264 207 2 1260 1 sky130_fd_sc_hd__and2_1 $T=372600 307360 1 0 $X=372410 $Y=304400
X2205 1 2 269 215 2 1283 1 sky130_fd_sc_hd__and2_1 $T=382260 280160 1 0 $X=382070 $Y=277200
X2206 1 2 273 207 2 1291 1 sky130_fd_sc_hd__and2_1 $T=387320 301920 0 0 $X=387130 $Y=301680
X2207 1 2 278 215 2 1293 1 sky130_fd_sc_hd__and2_1 $T=395600 247520 0 0 $X=395410 $Y=247280
X2208 1 2 281 215 2 1311 1 sky130_fd_sc_hd__and2_1 $T=397900 263840 1 0 $X=397710 $Y=260880
X2209 1 2 286 215 2 1319 1 sky130_fd_sc_hd__and2_1 $T=402960 274720 1 0 $X=402770 $Y=271760
X2210 1 2 289 207 2 1323 1 sky130_fd_sc_hd__and2_1 $T=406180 307360 1 0 $X=405990 $Y=304400
X2211 1 2 294 215 2 295 1 sky130_fd_sc_hd__and2_1 $T=410320 247520 1 0 $X=410130 $Y=244560
X2212 1 2 300 215 2 1359 1 sky130_fd_sc_hd__and2_1 $T=424120 258400 0 0 $X=423930 $Y=258160
X2213 1 2 301 207 2 1358 1 sky130_fd_sc_hd__and2_1 $T=424580 301920 1 0 $X=424390 $Y=298960
X2214 1 2 309 215 2 1376 1 sky130_fd_sc_hd__and2_1 $T=433320 247520 1 0 $X=433130 $Y=244560
X2215 1 2 313 215 2 1379 1 sky130_fd_sc_hd__and2_1 $T=441140 269280 1 0 $X=440950 $Y=266320
X2216 1 2 315 207 2 1409 1 sky130_fd_sc_hd__and2_1 $T=446200 307360 0 0 $X=446010 $Y=307120
X2217 1 2 317 215 2 1414 1 sky130_fd_sc_hd__and2_1 $T=450800 274720 0 0 $X=450610 $Y=274480
X2218 1 2 322 215 2 1433 1 sky130_fd_sc_hd__and2_1 $T=457700 258400 1 0 $X=457510 $Y=255440
X2219 1 2 327 215 2 1448 1 sky130_fd_sc_hd__and2_1 $T=466440 274720 1 0 $X=466250 $Y=271760
X2220 1 2 329 207 2 1456 1 sky130_fd_sc_hd__and2_1 $T=466440 301920 1 0 $X=466250 $Y=298960
X2221 1 2 342 215 2 1461 1 sky130_fd_sc_hd__and2_1 $T=484380 247520 1 0 $X=484190 $Y=244560
X2222 1 2 344 207 2 345 1 sky130_fd_sc_hd__and2_1 $T=485760 312800 1 0 $X=485570 $Y=309840
X2223 1 2 340 215 2 1482 1 sky130_fd_sc_hd__and2_1 $T=486680 252960 1 0 $X=486490 $Y=250000
X2224 1 2 350 215 2 1499 1 sky130_fd_sc_hd__and2_1 $T=490360 269280 0 0 $X=490170 $Y=269040
X2225 1 2 242 351 2 1501 1 sky130_fd_sc_hd__and2_1 $T=491740 274720 0 0 $X=491550 $Y=274480
X2226 1 2 300 351 2 1505 1 sky130_fd_sc_hd__and2_1 $T=493580 263840 1 0 $X=493390 $Y=260880
X2227 1 2 294 351 2 1500 1 sky130_fd_sc_hd__and2_1 $T=495420 247520 0 0 $X=495230 $Y=247280
X2228 1 2 360 207 2 1517 1 sky130_fd_sc_hd__and2_1 $T=498640 301920 0 0 $X=498450 $Y=301680
X2229 1 2 297 351 2 1522 1 sky130_fd_sc_hd__and2_1 $T=502780 269280 1 0 $X=502590 $Y=266320
X2230 1 2 212 366 2 1543 1 sky130_fd_sc_hd__and2_1 $T=508300 307360 0 0 $X=508110 $Y=307120
X2231 1 2 309 351 2 1560 1 sky130_fd_sc_hd__and2_1 $T=522560 252960 1 0 $X=522370 $Y=250000
X2232 1 2 286 351 2 1568 1 sky130_fd_sc_hd__and2_1 $T=522560 285600 1 0 $X=522370 $Y=282640
X2233 1 2 246 366 2 408 1 sky130_fd_sc_hd__and2_1 $T=542340 312800 1 0 $X=542150 $Y=309840
X2234 1 2 340 351 2 1616 1 sky130_fd_sc_hd__and2_1 $T=549240 252960 1 0 $X=549050 $Y=250000
X2235 1 2 322 351 2 1608 1 sky130_fd_sc_hd__and2_1 $T=551080 258400 0 0 $X=550890 $Y=258160
X2236 1 2 273 366 2 1627 1 sky130_fd_sc_hd__and2_1 $T=557520 307360 1 0 $X=557330 $Y=304400
X2237 1 2 317 351 2 1640 1 sky130_fd_sc_hd__and2_1 $T=563960 280160 0 0 $X=563770 $Y=279920
X2238 1 2 414 215 2 1647 1 sky130_fd_sc_hd__and2_1 $T=567640 280160 1 0 $X=567450 $Y=277200
X2239 1 2 414 351 2 1671 1 sky130_fd_sc_hd__and2_1 $T=578220 280160 1 0 $X=578030 $Y=277200
X2240 1 2 420 215 2 1679 1 sky130_fd_sc_hd__and2_1 $T=581900 274720 1 0 $X=581710 $Y=271760
X2241 1 2 428 215 2 1722 1 sky130_fd_sc_hd__and2_1 $T=605360 252960 1 0 $X=605170 $Y=250000
X2242 1 2 342 351 2 1726 1 sky130_fd_sc_hd__and2_1 $T=606740 285600 1 0 $X=606550 $Y=282640
X2243 1 2 431 215 2 1731 1 sky130_fd_sc_hd__and2_1 $T=607660 274720 0 0 $X=607470 $Y=274480
X2244 1 2 301 366 2 1740 1 sky130_fd_sc_hd__and2_1 $T=609500 312800 1 0 $X=609310 $Y=309840
X2245 1 2 436 215 2 1759 1 sky130_fd_sc_hd__and2_1 $T=620540 247520 0 0 $X=620350 $Y=247280
X2246 1 2 439 215 2 1787 1 sky130_fd_sc_hd__and2_1 $T=633880 258400 1 0 $X=633690 $Y=255440
X2247 1 2 442 215 2 1785 1 sky130_fd_sc_hd__and2_1 $T=634800 258400 0 0 $X=634610 $Y=258160
X2248 1 2 327 351 2 1790 1 sky130_fd_sc_hd__and2_1 $T=634800 285600 1 0 $X=634610 $Y=282640
X2249 1 2 443 215 2 1792 1 sky130_fd_sc_hd__and2_1 $T=637560 274720 1 0 $X=637370 $Y=271760
X2250 1 2 313 351 2 1840 1 sky130_fd_sc_hd__and2_1 $T=665620 263840 1 0 $X=665430 $Y=260880
X2251 1 2 350 351 2 1850 1 sky130_fd_sc_hd__and2_1 $T=665620 269280 1 0 $X=665430 $Y=266320
X2252 1 2 360 366 2 1864 1 sky130_fd_sc_hd__and2_1 $T=672980 312800 1 0 $X=672790 $Y=309840
X2253 1 2 431 351 2 1902 1 sky130_fd_sc_hd__and2_1 $T=690920 280160 1 0 $X=690730 $Y=277200
X2254 1 2 420 351 2 1905 1 sky130_fd_sc_hd__and2_1 $T=691840 263840 0 0 $X=691650 $Y=263600
X2255 1 2 436 351 2 1897 1 sky130_fd_sc_hd__and2_1 $T=693680 252960 1 0 $X=693490 $Y=250000
X2256 1 2 329 366 2 457 1 sky130_fd_sc_hd__and2_1 $T=698740 307360 1 0 $X=698550 $Y=304400
X2257 1 2 447 351 2 460 1 sky130_fd_sc_hd__and2_1 $T=711620 247520 1 0 $X=711430 $Y=244560
X2258 1 2 428 351 2 1941 1 sky130_fd_sc_hd__and2_1 $T=714840 258400 0 0 $X=714650 $Y=258160
X2259 1 2 105 9 2 524 1 sky130_fd_sc_hd__dlclkp_1 $T=6900 312800 1 0 $X=6710 $Y=309840
X2260 1 2 105 528 2 523 1 sky130_fd_sc_hd__dlclkp_1 $T=7360 258400 0 0 $X=7170 $Y=258160
X2261 1 2 105 529 2 525 1 sky130_fd_sc_hd__dlclkp_1 $T=7820 291040 0 0 $X=7630 $Y=290800
X2262 1 2 105 531 2 530 1 sky130_fd_sc_hd__dlclkp_1 $T=14260 291040 0 0 $X=14070 $Y=290800
X2263 1 2 105 551 2 522 1 sky130_fd_sc_hd__dlclkp_1 $T=15180 269280 0 0 $X=14990 $Y=269040
X2264 1 2 105 38 2 32 1 sky130_fd_sc_hd__dlclkp_1 $T=34040 247520 0 0 $X=33850 $Y=247280
X2265 1 2 105 580 2 581 1 sky130_fd_sc_hd__dlclkp_1 $T=40940 291040 1 0 $X=40750 $Y=288080
X2266 1 2 105 604 2 579 1 sky130_fd_sc_hd__dlclkp_1 $T=50600 263840 0 0 $X=50410 $Y=263600
X2267 1 2 105 605 2 628 1 sky130_fd_sc_hd__dlclkp_1 $T=52900 269280 1 0 $X=52710 $Y=266320
X2268 1 2 105 639 2 617 1 sky130_fd_sc_hd__dlclkp_1 $T=60720 285600 1 0 $X=60530 $Y=282640
X2269 1 2 105 643 2 619 1 sky130_fd_sc_hd__dlclkp_1 $T=62100 252960 0 0 $X=61910 $Y=252720
X2270 1 2 105 653 2 618 1 sky130_fd_sc_hd__dlclkp_1 $T=68080 301920 1 0 $X=67890 $Y=298960
X2271 1 2 105 661 2 664 1 sky130_fd_sc_hd__dlclkp_1 $T=72680 269280 0 0 $X=72490 $Y=269040
X2272 1 2 105 680 2 665 1 sky130_fd_sc_hd__dlclkp_1 $T=81420 291040 0 0 $X=81230 $Y=290800
X2273 1 2 105 702 2 685 1 sky130_fd_sc_hd__dlclkp_1 $T=92000 307360 0 0 $X=91810 $Y=307120
X2274 1 2 105 709 2 708 1 sky130_fd_sc_hd__dlclkp_1 $T=94760 291040 1 0 $X=94570 $Y=288080
X2275 1 2 105 714 2 707 1 sky130_fd_sc_hd__dlclkp_1 $T=96140 280160 1 0 $X=95950 $Y=277200
X2276 1 2 105 728 2 738 1 sky130_fd_sc_hd__dlclkp_1 $T=104420 307360 1 0 $X=104230 $Y=304400
X2277 1 2 105 732 2 84 1 sky130_fd_sc_hd__dlclkp_1 $T=105340 252960 1 0 $X=105150 $Y=250000
X2278 1 2 105 750 2 755 1 sky130_fd_sc_hd__dlclkp_1 $T=118220 296480 0 0 $X=118030 $Y=296240
X2279 1 2 105 763 2 764 1 sky130_fd_sc_hd__dlclkp_1 $T=121900 258400 1 0 $X=121710 $Y=255440
X2280 1 2 105 751 2 744 1 sky130_fd_sc_hd__dlclkp_1 $T=122360 274720 1 0 $X=122170 $Y=271760
X2281 1 2 105 785 2 789 1 sky130_fd_sc_hd__dlclkp_1 $T=132480 269280 1 0 $X=132290 $Y=266320
X2282 1 2 105 788 2 761 1 sky130_fd_sc_hd__dlclkp_1 $T=133400 285600 1 0 $X=133210 $Y=282640
X2283 1 2 105 807 2 810 1 sky130_fd_sc_hd__dlclkp_1 $T=141680 301920 1 0 $X=141490 $Y=298960
X2284 1 2 105 816 2 813 1 sky130_fd_sc_hd__dlclkp_1 $T=148580 258400 1 0 $X=148390 $Y=255440
X2285 1 2 105 817 2 809 1 sky130_fd_sc_hd__dlclkp_1 $T=148580 280160 1 0 $X=148390 $Y=277200
X2286 1 2 105 821 2 101 1 sky130_fd_sc_hd__dlclkp_1 $T=150420 307360 1 0 $X=150230 $Y=304400
X2287 1 2 105 849 2 853 1 sky130_fd_sc_hd__dlclkp_1 $T=162380 285600 1 0 $X=162190 $Y=282640
X2288 1 2 105 855 2 854 1 sky130_fd_sc_hd__dlclkp_1 $T=165140 296480 0 0 $X=164950 $Y=296240
X2289 1 2 105 858 2 859 1 sky130_fd_sc_hd__dlclkp_1 $T=166060 263840 0 0 $X=165870 $Y=263600
X2290 1 2 105 860 2 115 1 sky130_fd_sc_hd__dlclkp_1 $T=167440 252960 0 0 $X=167250 $Y=252720
X2291 1 2 105 898 2 906 1 sky130_fd_sc_hd__dlclkp_1 $T=188600 301920 1 0 $X=188410 $Y=298960
X2292 1 2 105 900 2 140 1 sky130_fd_sc_hd__dlclkp_1 $T=189520 247520 1 0 $X=189330 $Y=244560
X2293 1 2 105 905 2 899 1 sky130_fd_sc_hd__dlclkp_1 $T=191820 291040 0 0 $X=191630 $Y=290800
X2294 1 2 105 914 2 927 1 sky130_fd_sc_hd__dlclkp_1 $T=195500 263840 0 0 $X=195310 $Y=263600
X2295 1 2 105 147 2 141 1 sky130_fd_sc_hd__dlclkp_1 $T=207920 247520 0 0 $X=207730 $Y=247280
X2296 1 2 105 947 2 950 1 sky130_fd_sc_hd__dlclkp_1 $T=212060 291040 0 0 $X=211870 $Y=290800
X2297 1 2 105 953 2 956 1 sky130_fd_sc_hd__dlclkp_1 $T=218500 274720 1 0 $X=218310 $Y=271760
X2298 1 2 105 976 2 983 1 sky130_fd_sc_hd__dlclkp_1 $T=226320 258400 1 0 $X=226130 $Y=255440
X2299 1 2 105 984 2 987 1 sky130_fd_sc_hd__dlclkp_1 $T=229540 263840 1 0 $X=229350 $Y=260880
X2300 1 2 105 985 2 990 1 sky130_fd_sc_hd__dlclkp_1 $T=230460 280160 1 0 $X=230270 $Y=277200
X2301 1 2 105 980 2 979 1 sky130_fd_sc_hd__dlclkp_1 $T=230460 301920 0 0 $X=230270 $Y=301680
X2302 1 2 105 1017 2 1020 1 sky130_fd_sc_hd__dlclkp_1 $T=244260 269280 0 0 $X=244070 $Y=269040
X2303 1 2 105 1028 2 1022 1 sky130_fd_sc_hd__dlclkp_1 $T=252080 301920 1 0 $X=251890 $Y=298960
X2304 1 2 105 1041 2 1045 1 sky130_fd_sc_hd__dlclkp_1 $T=256220 291040 1 0 $X=256030 $Y=288080
X2305 1 2 105 1094 2 170 1 sky130_fd_sc_hd__dlclkp_1 $T=282440 252960 1 0 $X=282250 $Y=250000
X2306 1 2 105 1098 2 1097 1 sky130_fd_sc_hd__dlclkp_1 $T=286580 274720 0 0 $X=286390 $Y=274480
X2307 1 2 105 1095 2 1096 1 sky130_fd_sc_hd__dlclkp_1 $T=286580 285600 0 0 $X=286390 $Y=285360
X2308 1 2 105 1101 2 1116 1 sky130_fd_sc_hd__dlclkp_1 $T=288420 301920 0 0 $X=288230 $Y=301680
X2309 1 2 105 1135 2 176 1 sky130_fd_sc_hd__dlclkp_1 $T=302220 252960 1 0 $X=302030 $Y=250000
X2310 1 2 105 1136 2 1142 1 sky130_fd_sc_hd__dlclkp_1 $T=302220 285600 1 0 $X=302030 $Y=282640
X2311 1 2 105 1160 2 1159 1 sky130_fd_sc_hd__dlclkp_1 $T=316940 307360 1 0 $X=316750 $Y=304400
X2312 1 2 105 1167 2 1176 1 sky130_fd_sc_hd__dlclkp_1 $T=322000 258400 0 0 $X=321810 $Y=258160
X2313 1 2 105 1168 2 1180 1 sky130_fd_sc_hd__dlclkp_1 $T=322000 285600 1 0 $X=321810 $Y=282640
X2314 1 2 105 1178 2 1182 1 sky130_fd_sc_hd__dlclkp_1 $T=328900 280160 1 0 $X=328710 $Y=277200
X2315 1 2 479 1200 2 1206 1 sky130_fd_sc_hd__dlclkp_1 $T=335800 307360 0 0 $X=335610 $Y=307120
X2316 1 2 239 1226 2 1230 1 sky130_fd_sc_hd__dlclkp_1 $T=353280 258400 0 0 $X=353090 $Y=258160
X2317 1 2 479 1227 2 1231 1 sky130_fd_sc_hd__dlclkp_1 $T=353280 307360 0 0 $X=353090 $Y=307120
X2318 1 2 239 1232 2 220 1 sky130_fd_sc_hd__dlclkp_1 $T=356500 247520 0 0 $X=356310 $Y=247280
X2319 1 2 479 1260 2 1258 1 sky130_fd_sc_hd__dlclkp_1 $T=371220 307360 0 0 $X=371030 $Y=307120
X2320 1 2 239 1283 2 1247 1 sky130_fd_sc_hd__dlclkp_1 $T=385020 280160 1 0 $X=384830 $Y=277200
X2321 1 2 479 1291 2 1292 1 sky130_fd_sc_hd__dlclkp_1 $T=386860 307360 1 0 $X=386670 $Y=304400
X2322 1 2 239 1293 2 1256 1 sky130_fd_sc_hd__dlclkp_1 $T=389160 247520 0 0 $X=388970 $Y=247280
X2323 1 2 239 1311 2 1274 1 sky130_fd_sc_hd__dlclkp_1 $T=398820 258400 1 0 $X=398630 $Y=255440
X2324 1 2 239 1319 2 1290 1 sky130_fd_sc_hd__dlclkp_1 $T=401120 269280 0 0 $X=400930 $Y=269040
X2325 1 2 479 1323 2 1322 1 sky130_fd_sc_hd__dlclkp_1 $T=403420 301920 0 0 $X=403230 $Y=301680
X2326 1 2 479 1358 2 1369 1 sky130_fd_sc_hd__dlclkp_1 $T=419980 301920 0 0 $X=419790 $Y=301680
X2327 1 2 239 1359 2 1321 1 sky130_fd_sc_hd__dlclkp_1 $T=420440 263840 1 0 $X=420250 $Y=260880
X2328 1 2 239 1376 2 1349 1 sky130_fd_sc_hd__dlclkp_1 $T=429640 247520 0 0 $X=429450 $Y=247280
X2329 1 2 239 1379 2 1380 1 sky130_fd_sc_hd__dlclkp_1 $T=431020 269280 0 0 $X=430830 $Y=269040
X2330 1 2 479 1409 2 1412 1 sky130_fd_sc_hd__dlclkp_1 $T=442060 307360 1 0 $X=441870 $Y=304400
X2331 1 2 239 1414 2 1418 1 sky130_fd_sc_hd__dlclkp_1 $T=446200 280160 1 0 $X=446010 $Y=277200
X2332 1 2 239 1433 2 1396 1 sky130_fd_sc_hd__dlclkp_1 $T=457240 252960 1 0 $X=457050 $Y=250000
X2333 1 2 239 1448 2 1454 1 sky130_fd_sc_hd__dlclkp_1 $T=463680 274720 0 0 $X=463490 $Y=274480
X2334 1 2 479 1456 2 1441 1 sky130_fd_sc_hd__dlclkp_1 $T=469200 301920 1 0 $X=469010 $Y=298960
X2335 1 2 239 1461 2 336 1 sky130_fd_sc_hd__dlclkp_1 $T=470580 247520 1 0 $X=470390 $Y=244560
X2336 1 2 239 1482 2 1459 1 sky130_fd_sc_hd__dlclkp_1 $T=480240 252960 1 0 $X=480050 $Y=250000
X2337 1 2 239 1499 2 1483 1 sky130_fd_sc_hd__dlclkp_1 $T=489900 269280 1 0 $X=489710 $Y=266320
X2338 1 2 239 1500 2 1513 1 sky130_fd_sc_hd__dlclkp_1 $T=490360 252960 1 0 $X=490170 $Y=250000
X2339 1 2 239 1501 2 1514 1 sky130_fd_sc_hd__dlclkp_1 $T=491280 280160 0 0 $X=491090 $Y=279920
X2340 1 2 239 1505 2 1515 1 sky130_fd_sc_hd__dlclkp_1 $T=492200 263840 0 0 $X=492010 $Y=263600
X2341 1 2 479 1517 2 1491 1 sky130_fd_sc_hd__dlclkp_1 $T=497260 307360 1 0 $X=497070 $Y=304400
X2342 1 2 239 1522 2 1521 1 sky130_fd_sc_hd__dlclkp_1 $T=500940 269280 0 0 $X=500750 $Y=269040
X2343 1 2 479 1543 2 379 1 sky130_fd_sc_hd__dlclkp_1 $T=512900 312800 1 0 $X=512710 $Y=309840
X2344 1 2 239 1560 2 1570 1 sky130_fd_sc_hd__dlclkp_1 $T=519340 252960 0 0 $X=519150 $Y=252720
X2345 1 2 239 1568 2 1572 1 sky130_fd_sc_hd__dlclkp_1 $T=526240 285600 1 0 $X=526050 $Y=282640
X2346 1 2 239 1581 2 1574 1 sky130_fd_sc_hd__dlclkp_1 $T=530840 263840 0 0 $X=530650 $Y=263600
X2347 1 2 239 1616 2 1618 1 sky130_fd_sc_hd__dlclkp_1 $T=553380 252960 1 0 $X=553190 $Y=250000
X2348 1 2 479 1627 2 1641 1 sky130_fd_sc_hd__dlclkp_1 $T=557060 301920 0 0 $X=556870 $Y=301680
X2349 1 2 239 1640 2 1630 1 sky130_fd_sc_hd__dlclkp_1 $T=560740 280160 1 0 $X=560550 $Y=277200
X2350 1 2 239 1647 2 1659 1 sky130_fd_sc_hd__dlclkp_1 $T=568100 274720 0 0 $X=567910 $Y=274480
X2351 1 2 239 1679 2 1672 1 sky130_fd_sc_hd__dlclkp_1 $T=580520 269280 0 0 $X=580330 $Y=269040
X2352 1 2 239 1671 2 1677 1 sky130_fd_sc_hd__dlclkp_1 $T=581440 285600 1 0 $X=581250 $Y=282640
X2353 1 2 479 422 2 1690 1 sky130_fd_sc_hd__dlclkp_1 $T=583280 312800 1 0 $X=583090 $Y=309840
X2354 1 2 239 1722 2 1714 1 sky130_fd_sc_hd__dlclkp_1 $T=602600 258400 1 0 $X=602410 $Y=255440
X2355 1 2 239 1726 2 1734 1 sky130_fd_sc_hd__dlclkp_1 $T=603060 285600 0 0 $X=602870 $Y=285360
X2356 1 2 239 1731 2 1708 1 sky130_fd_sc_hd__dlclkp_1 $T=604440 280160 0 0 $X=604250 $Y=279920
X2357 1 2 479 1740 2 1738 1 sky130_fd_sc_hd__dlclkp_1 $T=609500 307360 1 0 $X=609310 $Y=304400
X2358 1 2 239 1759 2 1735 1 sky130_fd_sc_hd__dlclkp_1 $T=617320 247520 1 0 $X=617130 $Y=244560
X2359 1 2 239 1785 2 1788 1 sky130_fd_sc_hd__dlclkp_1 $T=630660 263840 1 0 $X=630470 $Y=260880
X2360 1 2 239 1787 2 1791 1 sky130_fd_sc_hd__dlclkp_1 $T=632040 252960 0 0 $X=631850 $Y=252720
X2361 1 2 239 1790 2 1789 1 sky130_fd_sc_hd__dlclkp_1 $T=634340 285600 0 0 $X=634150 $Y=285360
X2362 1 2 239 1792 2 1793 1 sky130_fd_sc_hd__dlclkp_1 $T=637560 280160 1 0 $X=637370 $Y=277200
X2363 1 2 239 448 2 1846 1 sky130_fd_sc_hd__dlclkp_1 $T=658720 247520 1 0 $X=658530 $Y=244560
X2364 1 2 239 1840 2 1847 1 sky130_fd_sc_hd__dlclkp_1 $T=658720 263840 1 0 $X=658530 $Y=260880
X2365 1 2 239 1850 2 1841 1 sky130_fd_sc_hd__dlclkp_1 $T=669300 269280 0 0 $X=669110 $Y=269040
X2366 1 2 479 1864 2 1873 1 sky130_fd_sc_hd__dlclkp_1 $T=670680 307360 0 0 $X=670490 $Y=307120
X2367 1 2 239 1897 2 1900 1 sky130_fd_sc_hd__dlclkp_1 $T=686780 252960 0 0 $X=686590 $Y=252720
X2368 1 2 239 1905 2 1893 1 sky130_fd_sc_hd__dlclkp_1 $T=693680 269280 1 0 $X=693490 $Y=266320
X2369 1 2 239 1902 2 1886 1 sky130_fd_sc_hd__dlclkp_1 $T=693680 280160 1 0 $X=693490 $Y=277200
X2370 1 2 239 1941 2 1946 1 sky130_fd_sc_hd__dlclkp_1 $T=709780 263840 0 0 $X=709590 $Y=263600
X2371 1 2 523 25 561 ICV_35 $T=20240 258400 1 0 $X=20050 $Y=255440
X2372 1 2 579 10 577 ICV_35 $T=31740 269280 1 0 $X=31550 $Y=266320
X2373 1 2 579 11 587 ICV_35 $T=32200 258400 1 0 $X=32010 $Y=255440
X2374 1 2 579 26 589 ICV_35 $T=32660 263840 1 0 $X=32470 $Y=260880
X2375 1 2 581 5 590 ICV_35 $T=32660 291040 1 0 $X=32470 $Y=288080
X2376 1 2 579 5 598 ICV_35 $T=34040 263840 0 0 $X=33850 $Y=263600
X2377 1 2 582 5 599 ICV_35 $T=34040 274720 0 0 $X=33850 $Y=274480
X2378 1 2 579 14 608 ICV_35 $T=42320 263840 0 0 $X=42130 $Y=263600
X2379 1 2 617 10 632 ICV_35 $T=53360 280160 0 0 $X=53170 $Y=279920
X2380 1 2 617 11 656 ICV_35 $T=64400 291040 1 0 $X=64210 $Y=288080
X2381 1 2 62 4 659 ICV_35 $T=65780 307360 1 0 $X=65590 $Y=304400
X2382 1 2 628 24 663 ICV_35 $T=67620 263840 1 0 $X=67430 $Y=260880
X2383 1 2 670 5 686 ICV_35 $T=80040 252960 0 0 $X=79850 $Y=252720
X2384 1 2 685 24 694 ICV_35 $T=83720 301920 1 0 $X=83530 $Y=298960
X2385 1 2 685 14 698 ICV_35 $T=85100 307360 1 0 $X=84910 $Y=304400
X2386 1 2 71 25 79 ICV_35 $T=92920 247520 1 0 $X=92730 $Y=244560
X2387 1 2 708 10 724 ICV_35 $T=95680 285600 1 0 $X=95490 $Y=282640
X2388 1 2 708 4 727 ICV_35 $T=97980 291040 0 0 $X=97790 $Y=290800
X2389 1 2 707 26 729 ICV_35 $T=98900 263840 0 0 $X=98710 $Y=263600
X2390 1 2 84 10 706 ICV_35 $T=108560 252960 0 0 $X=108370 $Y=252720
X2391 1 2 744 5 768 ICV_35 $T=118220 263840 0 0 $X=118030 $Y=263600
X2392 1 2 764 14 784 ICV_35 $T=126500 252960 0 0 $X=126310 $Y=252720
X2393 1 2 738 24 786 ICV_35 $T=126960 301920 0 0 $X=126770 $Y=301680
X2394 1 2 813 4 833 ICV_35 $T=147660 252960 0 0 $X=147470 $Y=252720
X2395 1 2 789 14 838 ICV_35 $T=151800 269280 1 0 $X=151610 $Y=266320
X2396 1 2 101 24 844 ICV_35 $T=154560 307360 0 0 $X=154370 $Y=307120
X2397 1 2 853 110 871 ICV_35 $T=167900 280160 1 0 $X=167710 $Y=277200
X2398 1 2 109 110 120 ICV_35 $T=167900 312800 1 0 $X=167710 $Y=309840
X2399 1 2 854 128 885 ICV_35 $T=179400 296480 1 0 $X=179210 $Y=293520
X2400 1 2 137 108 917 ICV_35 $T=189980 307360 0 0 $X=189790 $Y=307120
X2401 1 2 140 125 926 ICV_35 $T=193660 247520 0 0 $X=193470 $Y=247280
X2402 1 2 919 110 931 ICV_35 $T=200100 269280 1 0 $X=199910 $Y=266320
X2403 1 2 141 127 150 ICV_35 $T=207460 247520 1 0 $X=207270 $Y=244560
X2404 1 2 141 125 948 ICV_35 $T=207920 252960 1 0 $X=207730 $Y=250000
X2405 1 2 919 127 952 ICV_35 $T=210220 269280 0 0 $X=210030 $Y=269040
X2406 1 2 927 126 965 ICV_35 $T=216660 258400 1 0 $X=216470 $Y=255440
X2407 1 2 956 112 977 ICV_35 $T=220800 269280 0 0 $X=220610 $Y=269040
X2408 1 2 956 110 981 ICV_35 $T=221720 280160 1 0 $X=221530 $Y=277200
X2409 1 2 979 110 1014 ICV_35 $T=236900 301920 0 0 $X=236710 $Y=301680
X2410 1 2 987 128 1038 ICV_35 $T=248860 258400 0 0 $X=248670 $Y=258160
X2411 1 2 1045 127 1062 ICV_35 $T=260820 285600 0 0 $X=260630 $Y=285360
X2412 1 2 1022 111 1066 ICV_35 $T=262660 291040 1 0 $X=262470 $Y=288080
X2413 1 2 1070 112 1085 ICV_35 $T=272780 301920 1 0 $X=272590 $Y=298960
X2414 1 2 1070 127 1102 ICV_35 $T=281060 301920 1 0 $X=280870 $Y=298960
X2415 1 2 1116 110 1141 ICV_35 $T=298080 296480 0 0 $X=297890 $Y=296240
X2416 1 2 1142 128 1119 ICV_35 $T=307280 280160 1 0 $X=307090 $Y=277200
X2417 1 2 176 111 1156 ICV_35 $T=308660 252960 1 0 $X=308470 $Y=250000
X2418 1 2 1159 111 1174 ICV_35 $T=317400 296480 1 0 $X=317210 $Y=293520
X2419 1 2 177 201 1191 ICV_35 $T=332580 247520 0 0 $X=332390 $Y=247280
X2420 1 2 1176 126 1208 ICV_35 $T=336260 263840 1 0 $X=336070 $Y=260880
X2421 1 2 1231 214 1241 ICV_35 $T=356960 301920 1 0 $X=356770 $Y=298960
X2422 1 2 1230 238 1254 ICV_35 $T=359720 258400 0 0 $X=359530 $Y=258160
X2423 1 2 1290 232 1306 ICV_35 $T=389620 274720 1 0 $X=389430 $Y=271760
X2424 1 2 1292 214 1308 ICV_35 $T=389620 301920 0 0 $X=389430 $Y=301680
X2425 1 2 1292 210 1314 ICV_35 $T=393300 296480 1 0 $X=393110 $Y=293520
X2426 1 2 1321 250 1339 ICV_35 $T=406180 263840 0 0 $X=405990 $Y=263600
X2427 1 2 1338 224 1354 ICV_35 $T=413080 285600 1 0 $X=412890 $Y=282640
X2428 1 2 1322 216 1355 ICV_35 $T=413080 291040 1 0 $X=412890 $Y=288080
X2429 1 2 298 222 1360 ICV_35 $T=414460 307360 0 0 $X=414270 $Y=307120
X2430 1 2 1349 253 1368 ICV_35 $T=418140 258400 1 0 $X=417950 $Y=255440
X2431 1 2 177 306 1378 ICV_35 $T=425960 285600 1 0 $X=425770 $Y=282640
X2432 1 2 1369 213 1386 ICV_35 $T=426880 301920 0 0 $X=426690 $Y=301680
X2433 1 2 1380 250 1405 ICV_35 $T=435160 274720 0 0 $X=434970 $Y=274480
X2434 1 2 1396 238 1374 ICV_35 $T=443440 269280 1 0 $X=443250 $Y=266320
X2435 1 2 316 250 1453 ICV_35 $T=460000 252960 0 0 $X=459810 $Y=252720
X2436 1 2 1441 210 1480 ICV_35 $T=473800 296480 0 0 $X=473610 $Y=296240
X2437 1 2 1483 227 1497 ICV_35 $T=483000 274720 0 0 $X=482810 $Y=274480
X2438 1 2 336 250 1508 ICV_35 $T=486680 247520 1 0 $X=486490 $Y=244560
X2439 1 2 1491 210 1538 ICV_35 $T=500480 296480 0 0 $X=500290 $Y=296240
X2440 1 2 1491 218 1540 ICV_35 $T=500940 301920 0 0 $X=500750 $Y=301680
X2441 1 2 177 373 380 ICV_35 $T=511520 307360 1 0 $X=511330 $Y=304400
X2442 1 2 177 376 384 ICV_35 $T=515200 307360 0 0 $X=515010 $Y=307120
X2443 1 2 1521 364 1566 ICV_35 $T=516580 269280 0 0 $X=516390 $Y=269040
X2444 1 2 177 382 1573 ICV_35 $T=519800 296480 0 0 $X=519610 $Y=296240
X2445 1 2 1572 357 1590 ICV_35 $T=529000 291040 0 0 $X=528810 $Y=290800
X2446 1 2 409 404 1614 ICV_35 $T=544640 312800 1 0 $X=544450 $Y=309840
X2447 1 2 1630 356 1645 ICV_35 $T=558440 285600 0 0 $X=558250 $Y=285360
X2448 1 2 1630 367 1651 ICV_35 $T=563040 291040 1 0 $X=562850 $Y=288080
X2449 1 2 1659 232 1674 ICV_35 $T=572700 285600 1 0 $X=572510 $Y=282640
X2450 1 2 1641 404 1675 ICV_35 $T=572700 301920 1 0 $X=572510 $Y=298960
X2451 1 2 1659 238 1680 ICV_35 $T=574540 274720 0 0 $X=574350 $Y=274480
X2452 1 2 1708 227 1733 ICV_35 $T=599380 269280 0 0 $X=599190 $Y=269040
X2453 1 2 1714 223 1762 ICV_35 $T=614560 258400 0 0 $X=614370 $Y=258160
X2454 1 2 1734 364 1764 ICV_35 $T=614560 291040 0 0 $X=614370 $Y=290800
X2455 1 2 437 399 1797 ICV_35 $T=634800 307360 0 0 $X=634610 $Y=307120
X2456 1 2 1793 253 1815 ICV_35 $T=639400 274720 0 0 $X=639210 $Y=274480
X2457 1 2 441 223 446 ICV_35 $T=649060 247520 1 0 $X=648870 $Y=244560
X2458 1 2 1788 250 1822 ICV_35 $T=649060 263840 1 0 $X=648870 $Y=260880
X2459 1 2 1791 232 1837 ICV_35 $T=651360 252960 0 0 $X=651170 $Y=252720
X2460 1 2 1820 385 1839 ICV_35 $T=651360 307360 0 0 $X=651170 $Y=307120
X2461 1 2 1847 358 1869 ICV_35 $T=667000 258400 0 0 $X=666810 $Y=258160
X2462 1 2 1886 368 1901 ICV_35 $T=684940 285600 0 0 $X=684750 $Y=285360
X2463 1 2 1873 399 1912 ICV_35 $T=686780 301920 0 0 $X=686590 $Y=301680
X2464 1 2 459 390 1948 ICV_35 $T=709320 312800 1 0 $X=709130 $Y=309840
X2465 1 2 1944 358 1975 ICV_35 $T=725880 285600 0 0 $X=725690 $Y=285360
X2466 1 2 1946 356 1979 ICV_35 $T=726800 269280 0 0 $X=726610 $Y=269040
X2467 1 2 1943 368 1980 ICV_35 $T=726800 280160 0 0 $X=726610 $Y=279920
X2468 1 2 530 4 549 ICV_36 $T=6900 296480 1 0 $X=6710 $Y=293520
X2469 1 2 617 4 654 ICV_36 $T=62100 274720 0 0 $X=61910 $Y=274480
X2470 1 2 84 26 87 ICV_36 $T=104420 247520 1 0 $X=104230 $Y=244560
X2471 1 2 813 14 851 ICV_36 $T=155940 252960 0 0 $X=155750 $Y=252720
X2472 1 2 115 110 875 ICV_36 $T=167900 252960 1 0 $X=167710 $Y=250000
X2473 1 2 853 126 888 ICV_36 $T=176180 285600 1 0 $X=175990 $Y=282640
X2474 1 2 115 127 895 ICV_36 $T=178020 252960 1 0 $X=177830 $Y=250000
X2475 1 2 899 125 920 ICV_36 $T=188600 291040 1 0 $X=188410 $Y=288080
X2476 1 2 983 111 156 ICV_36 $T=230460 247520 0 0 $X=230270 $Y=247280
X2477 1 2 157 108 1033 ICV_36 $T=245180 301920 0 0 $X=244990 $Y=301680
X2478 1 2 990 127 1036 ICV_36 $T=246560 274720 0 0 $X=246370 $Y=274480
X2479 1 2 166 126 1068 ICV_36 $T=262660 307360 0 0 $X=262470 $Y=307120
X2480 1 2 1070 108 1090 ICV_36 $T=272780 296480 1 0 $X=272590 $Y=293520
X2481 1 2 1142 112 1171 ICV_36 $T=314640 280160 0 0 $X=314450 $Y=279920
X2482 1 2 1159 126 1169 ICV_36 $T=314640 296480 0 0 $X=314450 $Y=296240
X2483 1 2 1142 127 1173 ICV_36 $T=315560 280160 1 0 $X=315370 $Y=277200
X2484 1 2 220 223 236 ICV_36 $T=342700 247520 0 0 $X=342510 $Y=247280
X2485 1 2 1231 218 1248 ICV_36 $T=356500 301920 0 0 $X=356310 $Y=301680
X2486 1 2 1274 232 1276 ICV_36 $T=378120 269280 0 0 $X=377930 $Y=269040
X2487 1 2 1256 232 1300 ICV_36 $T=385020 252960 1 0 $X=384830 $Y=250000
X2488 1 2 1292 219 1304 ICV_36 $T=386860 291040 0 0 $X=386670 $Y=290800
X2489 1 2 1322 217 1346 ICV_36 $T=406180 296480 0 0 $X=405990 $Y=296240
X2490 1 2 314 216 1417 ICV_36 $T=441140 312800 1 0 $X=440950 $Y=309840
X2491 1 2 177 370 378 ICV_36 $T=508760 301920 1 0 $X=508570 $Y=298960
X2492 1 2 362 367 1563 ICV_36 $T=514740 247520 1 0 $X=514550 $Y=244560
X2493 1 2 393 363 402 ICV_36 $T=529460 247520 1 0 $X=529270 $Y=244560
X2494 1 2 393 367 410 ICV_36 $T=539120 247520 0 0 $X=538930 $Y=247280
X2495 1 2 1630 359 1649 ICV_36 $T=560740 285600 1 0 $X=560550 $Y=282640
X2496 1 2 1846 368 1856 ICV_36 $T=659640 252960 0 0 $X=659450 $Y=252720
X2497 1 2 461 357 1959 ICV_36 $T=711620 247520 0 0 $X=711430 $Y=247280
X2498 1 2 32 25 591 ICV_37 $T=33580 252960 0 0 $X=33390 $Y=252720
X2499 1 2 581 4 595 ICV_37 $T=33580 285600 0 0 $X=33390 $Y=285360
X2500 1 2 628 26 648 ICV_37 $T=61640 258400 0 0 $X=61450 $Y=258160
X2501 1 2 628 25 650 ICV_37 $T=61640 263840 0 0 $X=61450 $Y=263600
X2502 1 2 618 25 649 ICV_37 $T=61640 291040 0 0 $X=61450 $Y=290800
X2503 1 2 664 4 677 ICV_37 $T=75900 274720 1 0 $X=75710 $Y=271760
X2504 1 2 62 24 682 ICV_37 $T=75900 307360 1 0 $X=75710 $Y=304400
X2505 1 2 664 25 704 ICV_37 $T=89700 263840 0 0 $X=89510 $Y=263600
X2506 1 2 665 24 712 ICV_37 $T=89700 280160 0 0 $X=89510 $Y=279920
X2507 1 2 707 25 739 ICV_37 $T=103960 258400 1 0 $X=103770 $Y=255440
X2508 1 2 707 5 733 ICV_37 $T=103960 269280 1 0 $X=103770 $Y=266320
X2509 1 2 707 24 735 ICV_37 $T=103960 274720 1 0 $X=103770 $Y=271760
X2510 1 2 764 11 787 ICV_37 $T=132020 252960 1 0 $X=131830 $Y=250000
X2511 1 2 92 5 100 ICV_37 $T=132020 312800 1 0 $X=131830 $Y=309840
X2512 1 2 809 11 819 ICV_37 $T=145820 274720 0 0 $X=145630 $Y=274480
X2513 1 2 810 26 826 ICV_37 $T=145820 296480 0 0 $X=145630 $Y=296240
X2514 1 2 101 25 814 ICV_37 $T=145820 301920 0 0 $X=145630 $Y=301680
X2515 1 2 813 10 856 ICV_37 $T=160080 252960 1 0 $X=159890 $Y=250000
X2516 1 2 809 5 847 ICV_37 $T=160080 280160 1 0 $X=159890 $Y=277200
X2517 1 2 115 108 129 ICV_37 $T=173880 247520 0 0 $X=173690 $Y=247280
X2518 1 2 861 110 879 ICV_37 $T=173880 269280 0 0 $X=173690 $Y=269040
X2519 1 2 853 111 881 ICV_37 $T=173880 285600 0 0 $X=173690 $Y=285360
X2520 1 2 861 125 904 ICV_37 $T=188140 274720 1 0 $X=187950 $Y=271760
X2521 1 2 919 111 929 ICV_37 $T=201940 274720 0 0 $X=201750 $Y=274480
X2522 1 2 950 112 961 ICV_37 $T=216200 285600 1 0 $X=216010 $Y=282640
X2523 1 2 906 110 959 ICV_37 $T=216200 301920 1 0 $X=216010 $Y=298960
X2524 1 2 950 111 995 ICV_37 $T=230000 280160 0 0 $X=229810 $Y=279920
X2525 1 2 987 126 1016 ICV_37 $T=244260 263840 1 0 $X=244070 $Y=260880
X2526 1 2 990 111 1026 ICV_37 $T=244260 285600 1 0 $X=244070 $Y=282640
X2527 1 2 979 111 1006 ICV_37 $T=244260 296480 1 0 $X=244070 $Y=293520
X2528 1 2 979 128 974 ICV_37 $T=244260 301920 1 0 $X=244070 $Y=298960
X2529 1 2 1020 110 1049 ICV_37 $T=258060 269280 0 0 $X=257870 $Y=269040
X2530 1 2 163 112 1077 ICV_37 $T=272320 247520 1 0 $X=272130 $Y=244560
X2531 1 2 163 108 1081 ICV_37 $T=272320 252960 1 0 $X=272130 $Y=250000
X2532 1 2 170 125 1089 ICV_37 $T=286120 247520 0 0 $X=285930 $Y=247280
X2533 1 2 1096 126 1109 ICV_37 $T=286120 280160 0 0 $X=285930 $Y=279920
X2534 1 2 171 127 1103 ICV_37 $T=286120 307360 0 0 $X=285930 $Y=307120
X2535 1 2 1097 126 1138 ICV_37 $T=300380 274720 1 0 $X=300190 $Y=271760
X2536 1 2 1096 128 1121 ICV_37 $T=300380 291040 1 0 $X=300190 $Y=288080
X2537 1 2 1116 125 1137 ICV_37 $T=300380 307360 1 0 $X=300190 $Y=304400
X2538 1 2 1129 111 1162 ICV_37 $T=314180 258400 0 0 $X=313990 $Y=258160
X2539 1 2 1176 111 1193 ICV_37 $T=328440 263840 1 0 $X=328250 $Y=260880
X2540 1 2 1182 125 1181 ICV_37 $T=328440 269280 1 0 $X=328250 $Y=266320
X2541 1 2 1159 125 1194 ICV_37 $T=328440 296480 1 0 $X=328250 $Y=293520
X2542 1 2 1159 127 1187 ICV_37 $T=328440 307360 1 0 $X=328250 $Y=304400
X2543 1 2 1206 218 1218 ICV_37 $T=342240 307360 0 0 $X=342050 $Y=307120
X2544 1 2 1256 253 1268 ICV_37 $T=370300 258400 0 0 $X=370110 $Y=258160
X2545 1 2 1247 238 1249 ICV_37 $T=370300 274720 0 0 $X=370110 $Y=274480
X2546 1 2 1274 227 1297 ICV_37 $T=384560 269280 1 0 $X=384370 $Y=266320
X2547 1 2 1274 251 1320 ICV_37 $T=398360 258400 0 0 $X=398170 $Y=258160
X2548 1 2 1274 224 1316 ICV_37 $T=398360 263840 0 0 $X=398170 $Y=263600
X2549 1 2 284 251 1344 ICV_37 $T=412620 247520 1 0 $X=412430 $Y=244560
X2550 1 2 284 238 1342 ICV_37 $T=412620 252960 1 0 $X=412430 $Y=250000
X2551 1 2 1321 227 1350 ICV_37 $T=412620 263840 1 0 $X=412430 $Y=260880
X2552 1 2 1338 232 1351 ICV_37 $T=412620 280160 1 0 $X=412430 $Y=277200
X2553 1 2 1338 253 1377 ICV_37 $T=426420 280160 0 0 $X=426230 $Y=279920
X2554 1 2 1396 223 1413 ICV_37 $T=440680 263840 1 0 $X=440490 $Y=260880
X2555 1 2 1380 232 1415 ICV_37 $T=440680 285600 1 0 $X=440490 $Y=282640
X2556 1 2 1412 213 1444 ICV_37 $T=454480 296480 0 0 $X=454290 $Y=296240
X2557 1 2 1412 218 1439 ICV_37 $T=454480 301920 0 0 $X=454290 $Y=301680
X2558 1 2 326 222 1460 ICV_37 $T=468740 307360 1 0 $X=468550 $Y=304400
X2559 1 2 326 217 1468 ICV_37 $T=468740 312800 1 0 $X=468550 $Y=309840
X2560 1 2 1459 232 1493 ICV_37 $T=482540 263840 0 0 $X=482350 $Y=263600
X2561 1 2 1483 238 1479 ICV_37 $T=482540 269280 0 0 $X=482350 $Y=269040
X2562 1 2 1483 253 1495 ICV_37 $T=482540 280160 0 0 $X=482350 $Y=279920
X2563 1 2 1483 232 1526 ICV_37 $T=496800 274720 1 0 $X=496610 $Y=271760
X2564 1 2 1514 358 1527 ICV_37 $T=496800 285600 1 0 $X=496610 $Y=282640
X2565 1 2 1513 367 1553 ICV_37 $T=510600 252960 0 0 $X=510410 $Y=252720
X2566 1 2 177 389 395 ICV_37 $T=524860 301920 1 0 $X=524670 $Y=298960
X2567 1 2 379 390 396 ICV_37 $T=524860 312800 1 0 $X=524670 $Y=309840
X2568 1 2 379 404 1602 ICV_37 $T=538660 307360 0 0 $X=538470 $Y=307120
X2569 1 2 1617 356 1633 ICV_37 $T=552920 269280 1 0 $X=552730 $Y=266320
X2570 1 2 1601 359 1634 ICV_37 $T=552920 280160 1 0 $X=552730 $Y=277200
X2571 1 2 1601 367 1625 ICV_37 $T=552920 285600 1 0 $X=552730 $Y=282640
X2572 1 2 1601 364 1626 ICV_37 $T=552920 296480 1 0 $X=552730 $Y=293520
X2573 1 2 412 227 1655 ICV_37 $T=566720 247520 0 0 $X=566530 $Y=247280
X2574 1 2 1630 363 1648 ICV_37 $T=566720 280160 0 0 $X=566530 $Y=279920
X2575 1 2 1641 401 1666 ICV_37 $T=566720 301920 0 0 $X=566530 $Y=301680
X2576 1 2 1641 407 1667 ICV_37 $T=566720 307360 0 0 $X=566530 $Y=307120
X2577 1 2 412 251 1670 ICV_37 $T=580980 252960 1 0 $X=580790 $Y=250000
X2578 1 2 1672 250 1691 ICV_37 $T=580980 258400 1 0 $X=580790 $Y=255440
X2579 1 2 1672 232 1686 ICV_37 $T=580980 269280 1 0 $X=580790 $Y=266320
X2580 1 2 424 253 1715 ICV_37 $T=594780 252960 0 0 $X=594590 $Y=252720
X2581 1 2 1672 251 1711 ICV_37 $T=594780 258400 0 0 $X=594590 $Y=258160
X2582 1 2 1677 358 1713 ICV_37 $T=594780 285600 0 0 $X=594590 $Y=285360
X2583 1 2 1735 232 434 ICV_37 $T=609040 247520 1 0 $X=608850 $Y=244560
X2584 1 2 1734 368 1742 ICV_37 $T=609040 296480 1 0 $X=608850 $Y=293520
X2585 1 2 1735 250 1774 ICV_37 $T=622840 252960 0 0 $X=622650 $Y=252720
X2586 1 2 1763 227 1776 ICV_37 $T=622840 280160 0 0 $X=622650 $Y=279920
X2587 1 2 1734 358 1768 ICV_37 $T=622840 285600 0 0 $X=622650 $Y=285360
X2588 1 2 1788 227 1799 ICV_37 $T=637100 269280 1 0 $X=636910 $Y=266320
X2589 1 2 1789 367 1803 ICV_37 $T=637100 291040 1 0 $X=636910 $Y=288080
X2590 1 2 441 232 1828 ICV_37 $T=650900 247520 0 0 $X=650710 $Y=247280
X2591 1 2 1793 238 1823 ICV_37 $T=650900 274720 0 0 $X=650710 $Y=274480
X2592 1 2 1793 232 1832 ICV_37 $T=650900 280160 0 0 $X=650710 $Y=279920
X2593 1 2 1841 368 1843 ICV_37 $T=665160 280160 1 0 $X=664970 $Y=277200
X2594 1 2 1848 358 1862 ICV_37 $T=665160 285600 1 0 $X=664970 $Y=282640
X2595 1 2 1848 368 1863 ICV_37 $T=665160 296480 1 0 $X=664970 $Y=293520
X2596 1 2 1820 399 1858 ICV_37 $T=665160 301920 1 0 $X=664970 $Y=298960
X2597 1 2 1820 418 1865 ICV_37 $T=665160 312800 1 0 $X=664970 $Y=309840
X2598 1 2 1846 364 1887 ICV_37 $T=678960 252960 0 0 $X=678770 $Y=252720
X2599 1 2 1841 357 1888 ICV_37 $T=678960 280160 0 0 $X=678770 $Y=279920
X2600 1 2 1848 356 1884 ICV_37 $T=678960 291040 0 0 $X=678770 $Y=290800
X2601 1 2 1873 407 1885 ICV_37 $T=678960 307360 0 0 $X=678770 $Y=307120
X2602 1 2 1900 367 1918 ICV_37 $T=693220 258400 1 0 $X=693030 $Y=255440
X2603 1 2 1900 357 1940 ICV_37 $T=707020 258400 0 0 $X=706830 $Y=258160
X2604 1 2 1951 357 466 ICV_37 $T=721280 258400 1 0 $X=721090 $Y=255440
X2605 1 2 1951 364 467 ICV_37 $T=721280 263840 1 0 $X=721090 $Y=260880
X2606 1 2 1946 357 1969 ICV_37 $T=721280 269280 1 0 $X=721090 $Y=266320
X2607 1 2 1943 359 1971 ICV_37 $T=721280 280160 1 0 $X=721090 $Y=277200
X2608 1 2 461 368 1988 ICV_37 $T=735080 247520 0 0 $X=734890 $Y=247280
X2609 1 2 1951 358 1987 ICV_37 $T=735080 252960 0 0 $X=734890 $Y=252720
X2610 1 2 1946 368 1989 ICV_37 $T=735080 269280 0 0 $X=734890 $Y=269040
X2611 1 2 21 26 588 42 14 606 ICV_38 $T=33120 307360 1 0 $X=32930 $Y=304400
X2612 1 2 685 25 697 685 4 713 ICV_38 $T=85560 296480 1 0 $X=85370 $Y=293520
X2613 1 2 738 25 790 755 10 795 ICV_38 $T=128800 296480 0 0 $X=128610 $Y=296240
X2614 1 2 101 14 843 101 10 746 ICV_38 $T=155480 301920 0 0 $X=155290 $Y=301680
X2615 1 2 810 24 839 810 5 841 ICV_38 $T=155940 285600 0 0 $X=155750 $Y=285360
X2616 1 2 163 126 1048 163 110 1060 ICV_38 $T=257600 252960 1 0 $X=257410 $Y=250000
X2617 1 2 1097 127 1117 1097 112 1127 ICV_38 $T=288420 263840 0 0 $X=288230 $Y=263600
X2618 1 2 177 180 187 177 188 193 ICV_38 $T=310960 291040 1 0 $X=310770 $Y=288080
X2619 1 2 208 210 221 208 216 237 ICV_38 $T=339020 312800 1 0 $X=338830 $Y=309840
X2620 1 2 1182 108 1212 177 229 1222 ICV_38 $T=340400 274720 1 0 $X=340210 $Y=271760
X2621 1 2 1247 223 1259 1247 253 1261 ICV_38 $T=366160 280160 1 0 $X=365970 $Y=277200
X2622 1 2 1369 216 1398 1369 219 1400 ICV_38 $T=434700 291040 0 0 $X=434510 $Y=290800
X2623 1 2 1412 216 1423 1412 219 1431 ICV_38 $T=447580 291040 1 0 $X=447390 $Y=288080
X2624 1 2 1418 232 1434 1418 253 1451 ICV_38 $T=452640 280160 1 0 $X=452450 $Y=277200
X2625 1 2 1514 363 1548 1514 367 1555 ICV_38 $T=506920 285600 1 0 $X=506730 $Y=282640
X2626 1 2 1572 358 1598 1572 363 1595 ICV_38 $T=534520 285600 1 0 $X=534330 $Y=282640
X2627 1 2 1841 364 1851 1841 356 1871 ICV_38 $T=660560 274720 0 0 $X=660370 $Y=274480
X2628 1 2 556 527 18 ICV_39 $T=20240 252960 1 0 $X=20050 $Y=250000
X2629 1 2 50 51 18 ICV_39 $T=50140 312800 1 0 $X=49950 $Y=309840
X2630 1 2 658 56 30 ICV_39 $T=76360 252960 1 0 $X=76170 $Y=250000
X2631 1 2 828 822 17 ICV_39 $T=155020 280160 1 0 $X=154830 $Y=277200
X2632 1 2 815 89 34 ICV_39 $T=155020 312800 1 0 $X=154830 $Y=309840
X2633 1 2 851 835 19 ICV_39 $T=164680 258400 0 0 $X=164490 $Y=258160
X2634 1 2 866 873 122 ICV_39 $T=174800 291040 0 0 $X=174610 $Y=290800
X2635 1 2 1106 1105 134 ICV_39 $T=291180 280160 1 0 $X=290990 $Y=277200
X2636 1 2 1147 1146 135 ICV_39 $T=309120 252960 0 0 $X=308930 $Y=252720
X2637 1 2 1155 1124 131 ICV_39 $T=318320 301920 1 0 $X=318130 $Y=298960
X2638 1 2 1169 1166 136 ICV_39 $T=323380 301920 1 0 $X=323190 $Y=298960
X2639 1 2 1149 172 135 ICV_39 $T=323380 307360 1 0 $X=323190 $Y=304400
X2640 1 2 1173 1123 134 ICV_39 $T=325220 280160 0 0 $X=325030 $Y=279920
X2641 1 2 1221 1203 185 ICV_39 $T=356960 312800 1 0 $X=356770 $Y=309840
X2642 1 2 1246 247 229 ICV_39 $T=365240 247520 0 0 $X=365050 $Y=247280
X2643 1 2 1264 1252 263 ICV_39 $T=379500 274720 1 0 $X=379310 $Y=271760
X2644 1 2 1304 1299 202 ICV_39 $T=398820 285600 0 0 $X=398630 $Y=285360
X2645 1 2 1341 1333 199 ICV_39 $T=415380 285600 0 0 $X=415190 $Y=285360
X2646 1 2 1350 1343 252 ICV_39 $T=419060 258400 0 0 $X=418870 $Y=258160
X2647 1 2 1443 1437 260 ICV_39 $T=461380 274720 1 0 $X=461190 $Y=271760
X2648 1 2 1421 319 229 ICV_39 $T=463680 252960 1 0 $X=463490 $Y=250000
X2649 1 2 1468 334 192 ICV_39 $T=477480 307360 0 0 $X=477290 $Y=307120
X2650 1 2 1477 1467 257 ICV_39 $T=483000 285600 0 0 $X=482810 $Y=285360
X2651 1 2 1526 1484 257 ICV_39 $T=505540 274720 0 0 $X=505350 $Y=274480
X2652 1 2 1545 1534 372 ICV_39 $T=512440 263840 0 0 $X=512250 $Y=263600
X2653 1 2 1639 1615 306 ICV_39 $T=561660 274720 0 0 $X=561470 $Y=274480
X2654 1 2 1733 1723 252 ICV_39 $T=609500 269280 1 0 $X=609310 $Y=266320
X2655 1 2 1784 1761 257 ICV_39 $T=632040 291040 1 0 $X=631850 $Y=288080
X2656 1 2 1806 1802 229 ICV_39 $T=651360 269280 0 0 $X=651170 $Y=269040
X2657 1 2 1832 1813 257 ICV_39 $T=660100 285600 1 0 $X=659910 $Y=282640
X2658 1 2 1837 1812 257 ICV_39 $T=665620 258400 1 0 $X=665430 $Y=255440
X2659 1 2 1939 1916 382 ICV_39 $T=714840 263840 1 0 $X=714650 $Y=260880
X2660 1 2 1957 1950 341 ICV_39 $T=721740 291040 1 0 $X=721550 $Y=288080
X2661 1 2 1953 1950 348 ICV_39 $T=721740 296480 1 0 $X=721550 $Y=293520
X2662 1 2 1987 462 328 ICV_39 $T=737840 258400 0 0 $X=737650 $Y=258160
X2663 1 2 1984 1965 337 ICV_39 $T=737840 274720 0 0 $X=737650 $Y=274480
X2664 1 2 1980 1965 382 ICV_39 $T=737840 280160 0 0 $X=737650 $Y=279920
X2665 1 2 561 527 30 ICV_40 $T=27140 252960 1 0 $X=26950 $Y=250000
X2666 1 2 609 45 19 ICV_40 $T=55200 252960 0 0 $X=55010 $Y=252720
X2667 1 2 637 56 33 ICV_40 $T=61640 258400 1 0 $X=61450 $Y=255440
X2668 1 2 631 642 13 ICV_40 $T=62100 301920 1 0 $X=61910 $Y=298960
X2669 1 2 729 730 34 ICV_40 $T=107180 263840 1 0 $X=106990 $Y=260880
X2670 1 2 747 740 19 ICV_40 $T=115000 280160 1 0 $X=114810 $Y=277200
X2671 1 2 768 718 16 ICV_40 $T=126040 247520 1 0 $X=125850 $Y=244560
X2672 1 2 795 772 13 ICV_40 $T=139380 285600 0 0 $X=139190 $Y=285360
X2673 1 2 839 824 33 ICV_40 $T=161920 291040 1 0 $X=161730 $Y=288080
X2674 1 2 840 824 13 ICV_40 $T=161920 307360 1 0 $X=161730 $Y=304400
X2675 1 2 848 822 13 ICV_40 $T=167440 274720 0 0 $X=167250 $Y=274480
X2676 1 2 886 873 135 ICV_40 $T=188600 296480 1 0 $X=188410 $Y=293520
X2677 1 2 938 921 123 ICV_40 $T=209760 269280 1 0 $X=209570 $Y=266320
X2678 1 2 939 144 131 ICV_40 $T=210220 301920 1 0 $X=210030 $Y=298960
X2679 1 2 952 921 134 ICV_40 $T=217120 269280 1 0 $X=216930 $Y=266320
X2680 1 2 1008 154 122 ICV_40 $T=240580 307360 0 0 $X=240390 $Y=307120
X2681 1 2 1085 1086 123 ICV_40 $T=280140 301920 0 0 $X=279950 $Y=301680
X2682 1 2 1131 1124 121 ICV_40 $T=300840 301920 1 0 $X=300650 $Y=298960
X2683 1 2 1137 1124 135 ICV_40 $T=303600 312800 1 0 $X=303410 $Y=309840
X2684 1 2 183 184 121 ICV_40 $T=315100 247520 0 0 $X=314910 $Y=247280
X2685 1 2 1177 184 135 ICV_40 $T=328900 252960 1 0 $X=328710 $Y=250000
X2686 1 2 1219 1203 199 ICV_40 $T=350060 301920 1 0 $X=349870 $Y=298960
X2687 1 2 1238 1245 192 ICV_40 $T=368920 296480 1 0 $X=368730 $Y=293520
X2688 1 2 1251 1245 178 ICV_40 $T=377660 307360 0 0 $X=377470 $Y=307120
X2689 1 2 1269 1252 233 ICV_40 $T=378120 285600 1 0 $X=377930 $Y=282640
X2690 1 2 1267 1273 252 ICV_40 $T=378580 258400 1 0 $X=378390 $Y=255440
X2691 1 2 1268 1273 229 ICV_40 $T=385020 258400 1 0 $X=384830 $Y=255440
X2692 1 2 1280 1253 188 ICV_40 $T=385020 301920 1 0 $X=384830 $Y=298960
X2693 1 2 1317 1299 185 ICV_40 $T=406640 301920 1 0 $X=406450 $Y=298960
X2694 1 2 1351 1348 257 ICV_40 $T=420440 285600 0 0 $X=420250 $Y=285360
X2695 1 2 1383 1387 199 ICV_40 $T=434700 291040 1 0 $X=434510 $Y=288080
X2696 1 2 1400 1387 202 ICV_40 $T=441600 291040 1 0 $X=441410 $Y=288080
X2697 1 2 1415 1406 257 ICV_40 $T=448040 285600 0 0 $X=447850 $Y=285360
X2698 1 2 1458 1449 202 ICV_40 $T=470120 296480 1 0 $X=469930 $Y=293520
X2699 1 2 1476 1470 263 ICV_40 $T=483000 258400 0 0 $X=482810 $Y=258160
X2700 1 2 1457 1449 180 ICV_40 $T=483000 296480 0 0 $X=482810 $Y=296240
X2701 1 2 1497 1484 252 ICV_40 $T=490820 280160 1 0 $X=490630 $Y=277200
X2702 1 2 1508 343 262 ICV_40 $T=497260 247520 1 0 $X=497070 $Y=244560
X2703 1 2 1531 1532 341 ICV_40 $T=504160 280160 0 0 $X=503970 $Y=279920
X2704 1 2 1566 1547 372 ICV_40 $T=525320 269280 1 0 $X=525130 $Y=266320
X2705 1 2 1550 1534 382 ICV_40 $T=533600 263840 1 0 $X=533410 $Y=260880
X2706 1 2 1610 1589 303 ICV_40 $T=546940 274720 1 0 $X=546750 $Y=271760
X2707 1 2 1675 1656 389 ICV_40 $T=581900 301920 1 0 $X=581710 $Y=298960
X2708 1 2 1682 1656 373 ICV_40 $T=582360 307360 1 0 $X=582170 $Y=304400
X2709 1 2 1741 1739 348 ICV_40 $T=613640 291040 1 0 $X=613450 $Y=288080
X2710 1 2 1750 1747 400 ICV_40 $T=616400 301920 0 0 $X=616210 $Y=301680
X2711 1 2 1851 1844 372 ICV_40 $T=668840 280160 0 0 $X=668650 $Y=279920
X2712 1 2 1878 1844 303 ICV_40 $T=680800 274720 0 0 $X=680610 $Y=274480
X2713 1 2 1889 1875 400 ICV_40 $T=686780 301920 1 0 $X=686590 $Y=298960
X2714 1 2 1901 1904 382 ICV_40 $T=691840 291040 0 0 $X=691650 $Y=290800
X2715 1 2 452 455 400 ICV_40 $T=695980 312800 1 0 $X=695790 $Y=309840
X2716 1 2 1934 1926 391 ICV_40 $T=708400 307360 0 0 $X=708210 $Y=307120
X2717 1 2 1978 1955 303 ICV_40 $T=736920 263840 0 0 $X=736730 $Y=263600
X2718 1 2 744 4 758 ICV_43 $T=120980 263840 1 0 $X=120790 $Y=260880
X2719 1 2 761 25 776 ICV_43 $T=120980 280160 1 0 $X=120790 $Y=277200
X2720 1 2 789 25 804 ICV_43 $T=136160 263840 1 0 $X=135970 $Y=260880
X2721 1 2 789 10 837 ICV_43 $T=152720 258400 0 0 $X=152530 $Y=258160
X2722 1 2 101 5 113 ICV_43 $T=162840 307360 0 0 $X=162650 $Y=307120
X2723 1 2 899 128 915 ICV_43 $T=190900 285600 0 0 $X=190710 $Y=285360
X2724 1 2 177 192 197 ICV_43 $T=322460 291040 0 0 $X=322270 $Y=290800
X2725 1 2 1182 128 1201 ICV_43 $T=331200 274720 0 0 $X=331010 $Y=274480
X2726 1 2 220 224 235 ICV_43 $T=345460 247520 1 0 $X=345270 $Y=244560
X2727 1 2 220 227 1223 ICV_43 $T=346840 252960 0 0 $X=346650 $Y=252720
X2728 1 2 1258 216 1275 ICV_43 $T=373520 291040 1 0 $X=373330 $Y=288080
X2729 1 2 1349 250 1404 ICV_43 $T=436080 247520 0 0 $X=435890 $Y=247280
X2730 1 2 316 227 1427 ICV_43 $T=449420 247520 1 0 $X=449230 $Y=244560
X2731 1 2 1441 219 1458 ICV_43 $T=463220 291040 0 0 $X=463030 $Y=290800
X2732 1 2 1789 368 1814 ICV_43 $T=639860 296480 0 0 $X=639670 $Y=296240
X2733 1 2 1841 367 1883 ICV_43 $T=681260 274720 1 0 $X=681070 $Y=271760
X2734 1 2 522 5 533 ICV_47 $T=5520 269280 0 0 $X=5330 $Y=269040
X2735 1 2 523 10 526 ICV_47 $T=6900 252960 0 0 $X=6710 $Y=252720
X2736 1 2 32 4 607 ICV_47 $T=40480 247520 0 0 $X=40290 $Y=247280
X2737 1 2 617 26 630 ICV_47 $T=51980 285600 1 0 $X=51790 $Y=282640
X2738 1 2 619 25 658 ICV_47 $T=65320 252960 1 0 $X=65130 $Y=250000
X2739 1 2 685 26 725 ICV_47 $T=95680 296480 0 0 $X=95490 $Y=296240
X2740 1 2 708 11 748 ICV_47 $T=107180 280160 0 0 $X=106990 $Y=279920
X2741 1 2 84 5 716 ICV_47 $T=111780 258400 1 0 $X=111590 $Y=255440
X2742 1 2 738 11 766 ICV_47 $T=118220 301920 0 0 $X=118030 $Y=301680
X2743 1 2 761 5 792 ICV_47 $T=128800 274720 0 0 $X=128610 $Y=274480
X2744 1 2 789 5 805 ICV_47 $T=134780 269280 0 0 $X=134590 $Y=269040
X2745 1 2 813 26 831 ICV_47 $T=146280 247520 0 0 $X=146090 $Y=247280
X2746 1 2 810 10 840 ICV_47 $T=154100 291040 0 0 $X=153910 $Y=290800
X2747 1 2 854 110 866 ICV_47 $T=166060 296480 1 0 $X=165870 $Y=293520
X2748 1 2 854 125 886 ICV_47 $T=177100 301920 1 0 $X=176910 $Y=298960
X2749 1 2 859 112 884 ICV_47 $T=178940 258400 0 0 $X=178750 $Y=258160
X2750 1 2 115 128 132 ICV_47 $T=179400 247520 1 0 $X=179210 $Y=244560
X2751 1 2 861 128 903 ICV_47 $T=183540 274720 0 0 $X=183350 $Y=274480
X2752 1 2 137 127 925 ICV_47 $T=192740 312800 1 0 $X=192550 $Y=309840
X2753 1 2 956 126 1007 ICV_47 $T=232760 274720 1 0 $X=232570 $Y=271760
X2754 1 2 1022 127 1046 ICV_47 $T=252080 296480 1 0 $X=251890 $Y=293520
X2755 1 2 1054 127 1073 ICV_47 $T=267720 252960 0 0 $X=267530 $Y=252720
X2756 1 2 1054 126 1099 ICV_47 $T=278760 263840 1 0 $X=278570 $Y=260880
X2757 1 2 1097 111 1108 ICV_47 $T=284280 269280 1 0 $X=284090 $Y=266320
X2758 1 2 1142 111 1150 ICV_47 $T=305440 274720 0 0 $X=305250 $Y=274480
X2759 1 2 1142 110 1157 ICV_47 $T=308200 274720 1 0 $X=308010 $Y=271760
X2760 1 2 1142 126 1172 ICV_47 $T=316940 274720 1 0 $X=316750 $Y=271760
X2761 1 2 179 108 194 ICV_47 $T=316940 312800 1 0 $X=316750 $Y=309840
X2762 1 2 176 127 195 ICV_47 $T=319240 247520 1 0 $X=319050 $Y=244560
X2763 1 2 1182 111 1196 ICV_47 $T=328900 274720 1 0 $X=328710 $Y=271760
X2764 1 2 1176 108 1205 ICV_47 $T=333500 252960 0 0 $X=333310 $Y=252720
X2765 1 2 1206 213 1202 ICV_47 $T=340400 301920 1 0 $X=340210 $Y=298960
X2766 1 2 220 238 1243 ICV_47 $T=356960 258400 1 0 $X=356770 $Y=255440
X2767 1 2 1230 250 1255 ICV_47 $T=359260 263840 1 0 $X=359070 $Y=260880
X2768 1 2 1256 227 1267 ICV_47 $T=369380 258400 1 0 $X=369190 $Y=255440
X2769 1 2 1247 224 1269 ICV_47 $T=370760 280160 0 0 $X=370570 $Y=279920
X2770 1 2 1258 219 1271 ICV_47 $T=370760 291040 0 0 $X=370570 $Y=290800
X2771 1 2 261 217 1284 ICV_47 $T=375820 312800 1 0 $X=375630 $Y=309840
X2772 1 2 1274 250 1286 ICV_47 $T=378120 258400 0 0 $X=377930 $Y=258160
X2773 1 2 1247 250 1285 ICV_47 $T=378120 274720 0 0 $X=377930 $Y=274480
X2774 1 2 1322 210 1341 ICV_47 $T=406180 291040 0 0 $X=405990 $Y=290800
X2775 1 2 1418 251 1435 ICV_47 $T=451720 274720 1 0 $X=451530 $Y=271760
X2776 1 2 1521 358 1546 ICV_47 $T=504620 274720 1 0 $X=504430 $Y=271760
X2777 1 2 177 372 1554 ICV_47 $T=511060 296480 0 0 $X=510870 $Y=296240
X2778 1 2 393 359 1592 ICV_47 $T=529920 247520 0 0 $X=529730 $Y=247280
X2779 1 2 379 399 1596 ICV_47 $T=532680 307360 1 0 $X=532490 $Y=304400
X2780 1 2 1601 358 1621 ICV_47 $T=545100 285600 0 0 $X=544910 $Y=285360
X2781 1 2 1617 367 1639 ICV_47 $T=553380 274720 1 0 $X=553190 $Y=271760
X2782 1 2 1641 388 1654 ICV_47 $T=563960 301920 1 0 $X=563770 $Y=298960
X2783 1 2 1659 251 1703 ICV_47 $T=584200 274720 0 0 $X=584010 $Y=274480
X2784 1 2 424 238 1687 ICV_47 $T=588800 252960 1 0 $X=588610 $Y=250000
X2785 1 2 1714 253 1727 ICV_47 $T=600300 263840 1 0 $X=600110 $Y=260880
X2786 1 2 1714 232 1737 ICV_47 $T=602600 263840 0 0 $X=602410 $Y=263600
X2787 1 2 1738 401 1750 ICV_47 $T=609500 301920 1 0 $X=609310 $Y=298960
X2788 1 2 1738 385 1757 ICV_47 $T=610880 307360 0 0 $X=610690 $Y=307120
X2789 1 2 1763 223 1783 ICV_47 $T=623300 274720 0 0 $X=623110 $Y=274480
X2790 1 2 1788 251 1795 ICV_47 $T=633420 263840 0 0 $X=633230 $Y=263600
X2791 1 2 1789 356 1796 ICV_47 $T=633420 291040 0 0 $X=633230 $Y=290800
X2792 1 2 1793 227 1811 ICV_47 $T=639400 280160 0 0 $X=639210 $Y=279920
X2793 1 2 1841 358 1854 ICV_47 $T=660560 269280 0 0 $X=660370 $Y=269040
X2794 1 2 1846 359 1876 ICV_47 $T=670220 247520 0 0 $X=670030 $Y=247280
X2795 1 2 1841 363 1878 ICV_47 $T=672520 274720 1 0 $X=672330 $Y=271760
X2796 1 2 456 390 1928 ICV_47 $T=698280 307360 0 0 $X=698090 $Y=307120
X2797 1 2 1900 358 1935 ICV_47 $T=701040 258400 1 0 $X=700850 $Y=255440
X2798 1 2 1944 357 1953 ICV_47 $T=711160 291040 0 0 $X=710970 $Y=290800
X2799 1 2 1943 357 1954 ICV_47 $T=711620 280160 1 0 $X=711430 $Y=277200
X2800 1 2 456 401 1962 ICV_47 $T=713460 296480 0 0 $X=713270 $Y=296240
X2801 1 2 46 47 18 ICV_48 $T=43700 312800 1 0 $X=43510 $Y=309840
X2802 1 2 626 627 19 ICV_48 $T=57500 269280 0 0 $X=57310 $Y=269040
X2803 1 2 745 74 30 ICV_48 $T=113620 247520 0 0 $X=113430 $Y=247280
X2804 1 2 746 89 13 ICV_48 $T=113620 307360 0 0 $X=113430 $Y=307120
X2805 1 2 97 89 18 ICV_48 $T=127880 301920 1 0 $X=127690 $Y=298960
X2806 1 2 114 116 117 ICV_48 $T=169740 258400 0 0 $X=169550 $Y=258160
X2807 1 2 885 873 131 ICV_48 $T=184000 291040 1 0 $X=183810 $Y=288080
X2808 1 2 918 921 121 ICV_48 $T=197800 269280 0 0 $X=197610 $Y=269040
X2809 1 2 944 139 134 ICV_48 $T=225860 296480 0 0 $X=225670 $Y=296240
X2810 1 2 1030 1012 123 ICV_48 $T=253920 280160 0 0 $X=253730 $Y=279920
X2811 1 2 1031 1032 135 ICV_48 $T=253920 296480 0 0 $X=253730 $Y=296240
X2812 1 2 1061 1059 135 ICV_48 $T=268180 274720 1 0 $X=267990 $Y=271760
X2813 1 2 1089 159 135 ICV_48 $T=281980 263840 0 0 $X=281790 $Y=263600
X2814 1 2 1075 1027 117 ICV_48 $T=281980 274720 0 0 $X=281790 $Y=274480
X2815 1 2 1076 1059 131 ICV_48 $T=281980 285600 0 0 $X=281790 $Y=285360
X2816 1 2 1087 1086 131 ICV_48 $T=281980 296480 0 0 $X=281790 $Y=296240
X2817 1 2 1120 1123 135 ICV_48 $T=296240 285600 1 0 $X=296050 $Y=282640
X2818 1 2 1198 1199 123 ICV_48 $T=338100 285600 0 0 $X=337910 $Y=285360
X2819 1 2 1250 1253 178 ICV_48 $T=366160 285600 0 0 $X=365970 $Y=285360
X2820 1 2 1266 1240 229 ICV_48 $T=380420 263840 1 0 $X=380230 $Y=260880
X2821 1 2 1330 1333 178 ICV_48 $T=408480 285600 1 0 $X=408290 $Y=282640
X2822 1 2 1331 280 199 ICV_48 $T=408480 307360 1 0 $X=408290 $Y=304400
X2823 1 2 311 312 233 ICV_48 $T=436540 247520 1 0 $X=436350 $Y=244560
X2824 1 2 1417 318 186 ICV_48 $T=450340 307360 0 0 $X=450150 $Y=307120
X2825 1 2 1502 1504 178 ICV_48 $T=492660 291040 1 0 $X=492470 $Y=288080
X2826 1 2 1585 1589 382 ICV_48 $T=534520 280160 0 0 $X=534330 $Y=279920
X2827 1 2 1699 1701 400 ICV_48 $T=590640 301920 0 0 $X=590450 $Y=301680
X2828 1 2 429 430 389 ICV_48 $T=604900 307360 1 0 $X=604710 $Y=304400
X2829 1 2 1760 1761 229 ICV_48 $T=618700 274720 0 0 $X=618510 $Y=274480
X2830 1 2 1777 1747 389 ICV_48 $T=632960 301920 1 0 $X=632770 $Y=298960
X2831 1 2 1816 1813 263 ICV_48 $T=646760 269280 0 0 $X=646570 $Y=269040
X2832 1 2 1899 1875 376 ICV_48 $T=689080 307360 1 0 $X=688890 $Y=304400
X2833 1 2 1921 1910 348 ICV_48 $T=702880 263840 0 0 $X=702690 $Y=263600
X2834 1 2 1973 462 303 ICV_48 $T=730940 258400 0 0 $X=730750 $Y=258160
X2835 1 2 526 527 13 523 14 553 ICV_51 $T=8280 258400 1 0 $X=8090 $Y=255440
X2836 1 2 606 47 19 618 10 631 ICV_51 $T=49680 301920 1 0 $X=49490 $Y=298960
X2837 1 2 610 585 30 618 5 634 ICV_51 $T=50140 296480 0 0 $X=49950 $Y=296240
X2838 1 2 612 602 34 617 24 636 ICV_51 $T=50600 274720 1 0 $X=50410 $Y=271760
X2839 1 2 760 718 34 764 10 767 ICV_51 $T=120520 252960 1 0 $X=120330 $Y=250000
X2840 1 2 787 771 18 764 25 799 ICV_51 $T=134780 247520 1 0 $X=134590 $Y=244560
X2841 1 2 808 771 16 813 25 832 ICV_51 $T=143520 252960 1 0 $X=143330 $Y=250000
X2842 1 2 819 822 18 809 14 845 ICV_51 $T=151800 269280 0 0 $X=151610 $Y=269040
X2843 1 2 875 116 122 115 126 896 ICV_51 $T=177100 252960 0 0 $X=176910 $Y=252720
X2844 1 2 908 139 135 141 111 930 ICV_51 $T=195040 252960 1 0 $X=194850 $Y=250000
X2845 1 2 151 144 135 153 108 972 ICV_51 $T=214820 307360 0 0 $X=214630 $Y=307120
X2846 1 2 991 975 135 979 112 1018 ICV_51 $T=235980 291040 0 0 $X=235790 $Y=290800
X2847 1 2 1046 1032 134 1022 110 1063 ICV_51 $T=259440 291040 0 0 $X=259250 $Y=290800
X2848 1 2 1134 1105 135 177 178 182 ICV_51 $T=302680 291040 0 0 $X=302490 $Y=290800
X2849 1 2 1202 1203 178 1206 214 1213 ICV_51 $T=337640 307360 1 0 $X=337450 $Y=304400
X2850 1 2 1242 1245 185 261 210 266 ICV_51 $T=364320 312800 1 0 $X=364130 $Y=309840
X2851 1 2 1303 1273 263 284 227 1326 ICV_51 $T=396060 252960 1 0 $X=395870 $Y=250000
X2852 1 2 1342 293 201 1349 223 1366 ICV_51 $T=414460 252960 0 0 $X=414270 $Y=252720
X2853 1 2 1344 293 263 1349 238 1367 ICV_51 $T=414920 247520 0 0 $X=414730 $Y=247280
X2854 1 2 1374 1375 201 1380 238 1394 ICV_51 $T=429180 269280 1 0 $X=428990 $Y=266320
X2855 1 2 1506 1504 186 1491 214 1536 ICV_51 $T=497260 301920 1 0 $X=497070 $Y=298960
X2856 1 2 1518 1519 348 362 357 1542 ICV_51 $T=499100 247520 0 0 $X=498910 $Y=247280
X2857 1 2 1758 1747 376 437 401 1786 ICV_51 $T=623300 307360 0 0 $X=623110 $Y=307120
X2858 1 2 1811 1813 252 1793 223 1821 ICV_51 $T=645840 280160 1 0 $X=645650 $Y=277200
X2859 1 2 1831 1802 257 1847 364 1852 ICV_51 $T=662860 263840 0 0 $X=662670 $Y=263600
X2860 1 2 1852 1853 372 1847 359 1872 ICV_51 $T=667920 269280 1 0 $X=667730 $Y=266320
X2861 1 2 654 641 17 ICV_52 $T=70380 280160 1 0 $X=70190 $Y=277200
X2862 1 2 701 676 34 ICV_52 $T=98440 269280 1 0 $X=98250 $Y=266320
X2863 1 2 752 757 19 ICV_52 $T=122360 301920 1 0 $X=122170 $Y=298960
X2864 1 2 805 811 16 ICV_52 $T=146280 269280 0 0 $X=146090 $Y=269040
X2865 1 2 803 779 13 ICV_52 $T=146280 285600 0 0 $X=146090 $Y=285360
X2866 1 2 837 811 13 ICV_52 $T=160540 263840 1 0 $X=160350 $Y=260880
X2867 1 2 883 863 117 ICV_52 $T=185840 263840 0 0 $X=185650 $Y=263600
X2868 1 2 966 933 117 ICV_52 $T=224480 252960 0 0 $X=224290 $Y=252720
X2869 1 2 1117 1104 134 ICV_52 $T=294860 269280 1 0 $X=294670 $Y=266320
X2870 1 2 1196 1183 117 ICV_52 $T=336720 263840 0 0 $X=336530 $Y=263600
X2871 1 2 1262 267 260 ICV_52 $T=379040 247520 1 0 $X=378850 $Y=244560
X2872 1 2 1357 1333 202 ICV_52 $T=421360 296480 1 0 $X=421170 $Y=293520
X2873 1 2 1394 1406 201 ICV_52 $T=448960 269280 0 0 $X=448770 $Y=269040
X2874 1 2 1429 1420 199 ICV_52 $T=460920 301920 1 0 $X=460730 $Y=298960
X2875 1 2 1539 355 185 ICV_52 $T=519340 312800 1 0 $X=519150 $Y=309840
X2876 1 2 1588 1589 306 ICV_52 $T=535440 280160 1 0 $X=535250 $Y=277200
X2877 1 2 1737 1730 257 ICV_52 $T=611800 263840 1 0 $X=611610 $Y=260880
X2878 1 2 1754 435 260 ICV_52 $T=621920 252960 1 0 $X=621730 $Y=250000
X2879 1 2 553 527 19 ICV_53 $T=15640 252960 0 0 $X=15450 $Y=252720
X2880 1 2 599 602 16 ICV_53 $T=40020 269280 1 0 $X=39830 $Y=266320
X2881 1 2 668 642 33 ICV_53 $T=76360 296480 1 0 $X=76170 $Y=293520
X2882 1 2 694 693 33 ICV_53 $T=90160 296480 0 0 $X=89970 $Y=296240
X2883 1 2 841 824 16 ICV_53 $T=160540 296480 1 0 $X=160350 $Y=293520
X2884 1 2 842 824 19 ICV_53 $T=160540 301920 1 0 $X=160350 $Y=298960
X2885 1 2 928 146 131 ICV_53 $T=202400 247520 0 0 $X=202210 $Y=247280
X2886 1 2 1048 161 136 ICV_53 $T=262200 252960 0 0 $X=262010 $Y=252720
X2887 1 2 1060 161 122 ICV_53 $T=266340 258400 1 0 $X=266150 $Y=255440
X2888 1 2 1157 1123 122 ICV_53 $T=314640 269280 0 0 $X=314450 $Y=269040
X2889 1 2 1546 1547 328 ICV_53 $T=511060 269280 0 0 $X=510870 $Y=269040
X2890 1 2 1535 1547 341 ICV_53 $T=511060 274720 0 0 $X=510870 $Y=274480
X2891 1 2 1713 1685 328 ICV_53 $T=599380 291040 1 0 $X=599190 $Y=288080
X2892 1 2 1721 423 263 ICV_53 $T=602600 252960 0 0 $X=602410 $Y=252720
X2893 1 2 1799 1802 252 ICV_53 $T=642160 263840 0 0 $X=641970 $Y=263600
X2894 1 2 1854 1844 328 ICV_53 $T=667000 274720 1 0 $X=666810 $Y=271760
X2895 1 2 1879 1866 303 ICV_53 $T=679420 285600 0 0 $X=679230 $Y=285360
X2896 1 2 458 454 372 ICV_53 $T=701500 247520 0 0 $X=701310 $Y=247280
X2897 1 2 1931 1910 328 ICV_53 $T=707480 269280 0 0 $X=707290 $Y=269040
X2898 1 2 1949 462 306 ICV_53 $T=715760 252960 1 0 $X=715570 $Y=250000
X2899 1 2 37 2 7 1 sky130_fd_sc_hd__clkbuf_16 $T=34040 269280 0 0 $X=33850 $Y=269040
X2900 1 2 37 2 207 1 sky130_fd_sc_hd__clkbuf_16 $T=329820 312800 1 0 $X=329630 $Y=309840
X2901 1 2 204 2 215 1 sky130_fd_sc_hd__clkbuf_16 $T=334880 252960 1 0 $X=334690 $Y=250000
X2902 1 2 225 2 238 1 sky130_fd_sc_hd__clkbuf_16 $T=346840 263840 0 0 $X=346650 $Y=263600
X2903 1 2 177 2 239 1 sky130_fd_sc_hd__clkbuf_16 $T=347300 263840 1 0 $X=347110 $Y=260880
X2904 1 2 240 2 128 1 sky130_fd_sc_hd__clkbuf_16 $T=356040 274720 0 0 $X=355850 $Y=274480
X2905 1 2 243 2 253 1 sky130_fd_sc_hd__clkbuf_16 $T=356960 280160 1 0 $X=356770 $Y=277200
X2906 1 2 249 2 110 1 sky130_fd_sc_hd__clkbuf_16 $T=358800 285600 1 0 $X=358610 $Y=282640
X2907 1 2 256 2 125 1 sky130_fd_sc_hd__clkbuf_16 $T=364320 291040 1 0 $X=364130 $Y=288080
X2908 1 2 259 2 108 1 sky130_fd_sc_hd__clkbuf_16 $T=368000 285600 1 0 $X=367810 $Y=282640
X2909 1 2 268 2 112 1 sky130_fd_sc_hd__clkbuf_16 $T=378120 285600 0 0 $X=377930 $Y=285360
X2910 1 2 272 2 126 1 sky130_fd_sc_hd__clkbuf_16 $T=387320 285600 0 0 $X=387130 $Y=285360
X2911 1 2 274 2 127 1 sky130_fd_sc_hd__clkbuf_16 $T=388240 285600 1 0 $X=388050 $Y=282640
X2912 1 2 283 2 111 1 sky130_fd_sc_hd__clkbuf_16 $T=398820 291040 1 0 $X=398630 $Y=288080
X2913 1 2 272 2 399 1 sky130_fd_sc_hd__clkbuf_16 $T=545100 301920 0 0 $X=544910 $Y=301680
X2914 1 2 274 2 388 1 sky130_fd_sc_hd__clkbuf_16 $T=554760 301920 1 0 $X=554570 $Y=298960
X2915 1 2 256 2 404 1 sky130_fd_sc_hd__clkbuf_16 $T=712080 301920 1 0 $X=711890 $Y=298960
X2916 1 2 240 2 401 1 sky130_fd_sc_hd__clkbuf_16 $T=724040 307360 1 0 $X=723850 $Y=304400
X2917 1 2 603 45 34 ICV_56 $T=49220 247520 1 0 $X=49030 $Y=244560
X2918 1 2 675 66 16 ICV_56 $T=82340 301920 0 0 $X=82150 $Y=301680
X2919 1 2 75 77 30 ICV_56 $T=96600 312800 1 0 $X=96410 $Y=309840
X2920 1 2 743 740 16 ICV_56 $T=117760 291040 1 0 $X=117570 $Y=288080
X2921 1 2 766 757 18 ICV_56 $T=125120 307360 1 0 $X=124930 $Y=304400
X2922 1 2 790 757 30 ICV_56 $T=136160 307360 1 0 $X=135970 $Y=304400
X2923 1 2 784 771 19 ICV_56 $T=138460 258400 0 0 $X=138270 $Y=258160
X2924 1 2 924 923 136 ICV_56 $T=210680 280160 0 0 $X=210490 $Y=279920
X2925 1 2 1033 164 121 ICV_56 $T=257140 307360 1 0 $X=256950 $Y=304400
X2926 1 2 1207 1183 136 ICV_56 $T=342700 280160 0 0 $X=342510 $Y=279920
X2927 1 2 1233 1199 121 ICV_56 $T=359260 285600 0 0 $X=359070 $Y=285360
X2928 1 2 1243 247 201 ICV_56 $T=365240 252960 1 0 $X=365050 $Y=250000
X2929 1 2 1284 270 192 ICV_56 $T=383640 307360 0 0 $X=383450 $Y=307120
X2930 1 2 1356 1343 260 ICV_56 $T=422280 269280 1 0 $X=422090 $Y=266320
X2931 1 2 1427 319 252 ICV_56 $T=455860 247520 0 0 $X=455670 $Y=247280
X2932 1 2 1481 1449 185 ICV_56 $T=489900 307360 1 0 $X=489710 $Y=304400
X2933 1 2 1594 1589 372 ICV_56 $T=540040 274720 1 0 $X=539850 $Y=271760
X2934 1 2 1602 394 389 ICV_56 $T=546020 301920 1 0 $X=545830 $Y=298960
X2935 1 2 1796 1804 337 ICV_56 $T=643540 291040 0 0 $X=643350 $Y=290800
X2936 1 2 1874 1859 348 ICV_56 $T=678960 258400 1 0 $X=678770 $Y=255440
X2937 1 2 1927 1904 348 ICV_56 $T=707480 285600 0 0 $X=707290 $Y=285360
X2938 1 2 530 5 552 548 545 13 ICV_58 $T=6900 285600 0 0 $X=6710 $Y=285360
X2939 1 2 664 26 701 704 676 30 ICV_58 $T=83720 269280 1 0 $X=83530 $Y=266320
X2940 1 2 761 10 803 806 779 18 ICV_58 $T=132480 280160 1 0 $X=132290 $Y=277200
X2941 1 2 861 127 902 902 862 134 ICV_58 $T=181700 269280 0 0 $X=181510 $Y=269040
X2942 1 2 899 108 922 881 874 117 ICV_58 $T=188600 285600 1 0 $X=188410 $Y=282640
X2943 1 2 141 126 964 964 146 136 ICV_58 $T=214360 247520 0 0 $X=214170 $Y=247280
X2944 1 2 927 111 966 965 933 136 ICV_58 $T=214360 258400 0 0 $X=214170 $Y=258160
X2945 1 2 983 125 1021 1021 155 135 ICV_58 $T=240580 252960 0 0 $X=240390 $Y=252720
X2946 1 2 1054 112 1069 1069 1053 123 ICV_58 $T=262660 263840 0 0 $X=262470 $Y=263600
X2947 1 2 1159 128 1189 1174 1166 117 ICV_58 $T=324760 296480 0 0 $X=324570 $Y=296240
X2948 1 2 1231 216 1236 1236 1245 186 ICV_58 $T=354200 291040 0 0 $X=354010 $Y=290800
X2949 1 2 298 217 1361 1361 302 192 ICV_58 $T=413080 312800 1 0 $X=412890 $Y=309840
X2950 1 2 1396 232 1411 1413 1375 260 ICV_58 $T=439300 258400 0 0 $X=439110 $Y=258160
X2951 1 2 1459 223 1492 1492 1470 260 ICV_58 $T=478860 263840 1 0 $X=478670 $Y=260880
X2952 1 2 1513 356 1523 1525 1519 341 ICV_58 $T=493120 258400 0 0 $X=492930 $Y=258160
X2953 1 2 1574 359 1587 1587 1589 341 ICV_58 $T=525320 274720 1 0 $X=525130 $Y=271760
X2954 1 2 1672 227 1694 1694 1688 252 ICV_58 $T=578680 263840 0 0 $X=578490 $Y=263600
X2955 1 2 1690 404 1728 1728 1701 389 ICV_58 $T=595240 296480 0 0 $X=595050 $Y=296240
X2956 1 2 1735 223 1754 1751 435 233 ICV_58 $T=608120 252960 0 0 $X=607930 $Y=252720
X2957 1 2 1738 399 1770 1770 1747 370 ICV_58 $T=618240 301920 1 0 $X=618050 $Y=298960
X2958 1 2 1763 232 1784 1783 1761 260 ICV_58 $T=621460 280160 1 0 $X=621270 $Y=277200
X2959 1 2 459 407 1974 1974 464 375 ICV_58 $T=721740 312800 1 0 $X=721550 $Y=309840
X2960 1 2 576 543 34 ICV_62 $T=33580 301920 1 0 $X=33390 $Y=298960
X2961 1 2 598 578 16 ICV_62 $T=48300 269280 1 0 $X=48110 $Y=266320
X2962 1 2 686 690 16 ICV_62 $T=90160 252960 0 0 $X=89970 $Y=252720
X2963 1 2 700 684 13 ICV_62 $T=104420 285600 1 0 $X=104230 $Y=282640
X2964 1 2 778 779 17 ICV_62 $T=132480 274720 1 0 $X=132290 $Y=271760
X2965 1 2 792 779 16 ICV_62 $T=137080 274720 1 0 $X=136890 $Y=271760
X2966 1 2 856 835 13 ICV_62 $T=169280 247520 0 0 $X=169090 $Y=247280
X2967 1 2 871 874 122 ICV_62 $T=175260 280160 0 0 $X=175070 $Y=279920
X2968 1 2 872 874 123 ICV_62 $T=179400 291040 1 0 $X=179210 $Y=288080
X2969 1 2 1007 973 136 ICV_62 $T=244720 274720 1 0 $X=244530 $Y=271760
X2970 1 2 1013 1012 136 ICV_62 $T=244720 280160 1 0 $X=244530 $Y=277200
X2971 1 2 1049 1027 122 ICV_62 $T=263580 274720 1 0 $X=263390 $Y=271760
X2972 1 2 1078 1053 121 ICV_62 $T=277380 263840 0 0 $X=277190 $Y=263600
X2973 1 2 1081 161 121 ICV_62 $T=281520 247520 0 0 $X=281330 $Y=247280
X2974 1 2 1118 159 123 ICV_62 $T=298080 258400 0 0 $X=297890 $Y=258160
X2975 1 2 1127 1104 123 ICV_62 $T=299920 269280 0 0 $X=299730 $Y=269040
X2976 1 2 1204 1183 134 ICV_62 $T=342700 269280 0 0 $X=342510 $Y=269040
X2977 1 2 1257 1245 199 ICV_62 $T=370760 301920 0 0 $X=370570 $Y=301680
X2978 1 2 1261 1252 229 ICV_62 $T=373520 285600 0 0 $X=373330 $Y=285360
X2979 1 2 1308 1299 180 ICV_62 $T=398820 301920 0 0 $X=398630 $Y=301680
X2980 1 2 1326 293 252 ICV_62 $T=408020 252960 1 0 $X=407830 $Y=250000
X2981 1 2 1363 302 199 ICV_62 $T=426880 307360 0 0 $X=426690 $Y=307120
X2982 1 2 1438 1437 201 ICV_62 $T=466440 269280 0 0 $X=466250 $Y=269040
X2983 1 2 1557 1519 382 ICV_62 $T=525320 252960 1 0 $X=525130 $Y=250000
X2984 1 2 1655 415 252 ICV_62 $T=572240 252960 1 0 $X=572050 $Y=250000
X2985 1 2 1689 1688 201 ICV_62 $T=590180 263840 1 0 $X=589990 $Y=260880
X2986 1 2 1711 1688 263 ICV_62 $T=598000 258400 1 0 $X=597810 $Y=255440
X2987 1 2 427 423 233 ICV_62 $T=604440 247520 1 0 $X=604250 $Y=244560
X2988 1 2 1818 1804 328 ICV_62 $T=647220 291040 1 0 $X=647030 $Y=288080
X2989 1 2 1912 1875 370 ICV_62 $T=694140 307360 1 0 $X=693950 $Y=304400
X2990 1 2 1914 1916 372 ICV_62 $T=698280 263840 0 0 $X=698090 $Y=263600
X2991 1 2 667 627 16 ICV_63 $T=76360 258400 1 0 $X=76170 $Y=255440
X2992 1 2 663 627 33 ICV_63 $T=76360 263840 1 0 $X=76170 $Y=260880
X2993 1 2 830 811 18 ICV_63 $T=154560 263840 1 0 $X=154370 $Y=260880
X2994 1 2 833 835 17 ICV_63 $T=155020 252960 1 0 $X=154830 $Y=250000
X2995 1 2 951 921 136 ICV_63 $T=216660 280160 1 0 $X=216470 $Y=277200
X2996 1 2 1141 1124 122 ICV_63 $T=304520 296480 1 0 $X=304330 $Y=293520
X2997 1 2 1210 1199 122 ICV_63 $T=342700 285600 0 0 $X=342510 $Y=285360
X2998 1 2 1241 1245 180 ICV_63 $T=364780 296480 0 0 $X=364590 $Y=296240
X2999 1 2 1249 1252 201 ICV_63 $T=365240 274720 0 0 $X=365050 $Y=274480
X3000 1 2 1287 1277 201 ICV_63 $T=386860 258400 0 0 $X=386670 $Y=258160
X3001 1 2 1310 1312 260 ICV_63 $T=397900 274720 1 0 $X=397710 $Y=271760
X3002 1 2 1335 1343 257 ICV_63 $T=413080 258400 1 0 $X=412890 $Y=255440
X3003 1 2 1403 1406 260 ICV_63 $T=441140 280160 1 0 $X=440950 $Y=277200
X3004 1 2 1428 319 263 ICV_63 $T=454940 252960 0 0 $X=454750 $Y=252720
X3005 1 2 1455 1449 192 ICV_63 $T=469200 285600 1 0 $X=469010 $Y=282640
X3006 1 2 1544 1519 303 ICV_63 $T=511060 258400 0 0 $X=510870 $Y=258160
X3007 1 2 1613 1615 372 ICV_63 $T=547860 269280 1 0 $X=547670 $Y=266320
X3008 1 2 1757 1747 391 ICV_63 $T=617320 307360 1 0 $X=617130 $Y=304400
X3009 1 2 1857 1824 361 ICV_63 $T=667920 296480 0 0 $X=667730 $Y=296240
X3010 1 2 1880 1866 372 ICV_63 $T=680340 291040 1 0 $X=680150 $Y=288080
X3011 1 2 1933 1926 370 ICV_63 $T=707480 301920 0 0 $X=707290 $Y=301680
X3012 1 2 755 4 781 ICV_66 $T=124660 291040 1 0 $X=124470 $Y=288080
X3013 1 2 764 5 808 ICV_66 $T=138460 252960 0 0 $X=138270 $Y=252720
X3014 1 2 853 108 864 ICV_66 $T=166520 280160 0 0 $X=166330 $Y=279920
X3015 1 2 854 108 865 ICV_66 $T=166520 291040 0 0 $X=166330 $Y=290800
X3016 1 2 919 128 949 ICV_66 $T=208840 280160 1 0 $X=208650 $Y=277200
X3017 1 2 990 126 1013 ICV_66 $T=236900 280160 1 0 $X=236710 $Y=277200
X3018 1 2 171 111 174 ICV_66 $T=293020 312800 1 0 $X=292830 $Y=309840
X3019 1 2 176 128 181 ICV_66 $T=306820 247520 0 0 $X=306630 $Y=247280
X3020 1 2 220 232 1228 ICV_66 $T=349140 258400 1 0 $X=348950 $Y=255440
X3021 1 2 1321 232 1335 ICV_66 $T=405260 258400 1 0 $X=405070 $Y=255440
X3022 1 2 1322 213 1330 ICV_66 $T=405260 296480 1 0 $X=405070 $Y=293520
X3023 1 2 1380 253 1395 ICV_66 $T=433320 280160 1 0 $X=433130 $Y=277200
X3024 1 2 316 253 1421 ICV_66 $T=447120 247520 0 0 $X=446930 $Y=247280
X3025 1 2 1521 357 1567 ICV_66 $T=517500 280160 1 0 $X=517310 $Y=277200
X3026 1 2 461 359 1956 ICV_66 $T=713920 247520 1 0 $X=713730 $Y=244560
X3027 1 2 1946 363 1978 ICV_66 $T=727720 263840 0 0 $X=727530 $Y=263600
X3028 1 2 523 4 534 534 527 17 ICV_68 $T=7360 247520 0 0 $X=7170 $Y=247280
X3029 1 2 525 4 538 538 545 17 ICV_68 $T=7820 274720 0 0 $X=7630 $Y=274480
X3030 1 2 582 24 597 597 602 33 ICV_68 $T=34500 274720 1 0 $X=34310 $Y=271760
X3031 1 2 32 10 620 620 45 13 ICV_68 $T=48300 258400 1 0 $X=48110 $Y=255440
X3032 1 2 665 25 674 674 684 30 ICV_68 $T=75900 285600 0 0 $X=75710 $Y=285360
X3033 1 2 670 11 689 692 690 30 ICV_68 $T=81420 252960 1 0 $X=81230 $Y=250000
X3034 1 2 664 10 711 711 676 13 ICV_68 $T=90160 274720 0 0 $X=89970 $Y=274480
X3035 1 2 92 4 794 796 757 17 ICV_68 $T=132020 307360 0 0 $X=131830 $Y=307120
X3036 1 2 810 4 825 825 824 17 ICV_68 $T=146280 296480 1 0 $X=146090 $Y=293520
X3037 1 2 859 108 880 880 863 121 ICV_68 $T=174340 258400 1 0 $X=174150 $Y=255440
X3038 1 2 927 108 958 958 933 121 ICV_68 $T=216200 263840 0 0 $X=216010 $Y=263600
X3039 1 2 153 112 970 970 154 123 ICV_68 $T=218500 312800 1 0 $X=218310 $Y=309840
X3040 1 2 983 112 993 993 155 123 ICV_68 $T=230460 252960 1 0 $X=230270 $Y=250000
X3041 1 2 979 126 999 999 975 136 ICV_68 $T=230920 301920 1 0 $X=230730 $Y=298960
X3042 1 2 990 125 1023 1026 1012 117 ICV_68 $T=244260 285600 0 0 $X=244070 $Y=285360
X3043 1 2 990 110 1037 1036 1012 134 ICV_68 $T=249320 280160 1 0 $X=249130 $Y=277200
X3044 1 2 1097 128 1114 1108 1104 117 ICV_68 $T=287040 274720 1 0 $X=286850 $Y=271760
X3045 1 2 1129 126 1143 1143 1146 136 ICV_68 $T=300840 263840 1 0 $X=300650 $Y=260880
X3046 1 2 1142 125 1120 1150 1123 117 ICV_68 $T=308660 285600 1 0 $X=308470 $Y=282640
X3047 1 2 1129 127 1165 1165 1146 134 ICV_68 $T=314640 263840 0 0 $X=314450 $Y=263600
X3048 1 2 1182 110 1214 1214 1183 122 ICV_68 $T=342700 274720 0 0 $X=342510 $Y=274480
X3049 1 2 1182 112 1215 1215 1183 123 ICV_68 $T=342700 280160 1 0 $X=342510 $Y=277200
X3050 1 2 1206 210 1219 1220 1203 202 ICV_68 $T=343160 291040 1 0 $X=342970 $Y=288080
X3051 1 2 258 251 276 277 267 201 ICV_68 $T=387780 247520 1 0 $X=387590 $Y=244560
X3052 1 2 1290 223 1310 1307 1312 233 ICV_68 $T=391460 280160 1 0 $X=391270 $Y=277200
X3053 1 2 1369 217 1382 1382 1387 192 ICV_68 $T=426880 296480 1 0 $X=426690 $Y=293520
X3054 1 2 1454 238 1465 1465 1467 201 ICV_68 $T=469200 263840 0 0 $X=469010 $Y=263600
X3055 1 2 1454 224 1478 1478 1467 233 ICV_68 $T=474260 285600 1 0 $X=474070 $Y=282640
X3056 1 2 1513 358 1524 1524 1519 328 ICV_68 $T=497260 252960 1 0 $X=497070 $Y=250000
X3057 1 2 1515 358 1564 1564 1534 328 ICV_68 $T=517500 263840 0 0 $X=517310 $Y=263600
X3058 1 2 1617 363 1657 1653 1615 382 ICV_68 $T=567180 269280 0 0 $X=566990 $Y=269040
X3059 1 2 1677 367 1692 1692 1685 306 ICV_68 $T=581440 285600 0 0 $X=581250 $Y=285360
X3060 1 2 1708 223 1753 1753 1723 260 ICV_68 $T=610420 274720 1 0 $X=610230 $Y=271760
X3061 1 2 1763 250 1781 1781 1761 262 ICV_68 $T=624220 269280 0 0 $X=624030 $Y=269040
X3062 1 2 1820 390 1836 1839 1824 391 ICV_68 $T=651820 312800 1 0 $X=651630 $Y=309840
X3063 1 2 1848 367 1860 1862 1866 328 ICV_68 $T=665160 285600 0 0 $X=664970 $Y=285360
X3064 1 2 1900 363 1917 1917 1916 303 ICV_68 $T=693220 252960 0 0 $X=693030 $Y=252720
X3065 1 2 461 364 1972 1972 463 372 ICV_68 $T=721740 247520 0 0 $X=721550 $Y=247280
X3066 1 2 461 358 469 470 463 303 ICV_68 $T=729560 247520 1 0 $X=729370 $Y=244560
X3067 1 2 461 356 1982 1982 463 337 ICV_68 $T=729560 252960 1 0 $X=729370 $Y=250000
X3068 1 2 530 11 554 ICV_69 $T=10580 291040 1 0 $X=10390 $Y=288080
X3069 1 2 32 11 41 ICV_69 $T=30820 247520 1 0 $X=30630 $Y=244560
X3070 1 2 42 25 629 ICV_69 $T=51980 301920 0 0 $X=51790 $Y=301680
X3071 1 2 628 5 667 ICV_69 $T=71300 258400 0 0 $X=71110 $Y=258160
X3072 1 2 670 4 719 ICV_69 $T=94760 252960 1 0 $X=94570 $Y=250000
X3073 1 2 744 11 717 ICV_69 $T=126500 263840 0 0 $X=126310 $Y=263600
X3074 1 2 109 126 891 ICV_69 $T=178940 312800 1 0 $X=178750 $Y=309840
X3075 1 2 853 128 897 ICV_69 $T=181700 285600 0 0 $X=181510 $Y=285360
X3076 1 2 1020 125 1044 ICV_69 $T=252540 269280 1 0 $X=252350 $Y=266320
X3077 1 2 1045 112 1064 ICV_69 $T=262660 280160 1 0 $X=262470 $Y=277200
X3078 1 2 166 110 1071 ICV_69 $T=272780 307360 0 0 $X=272590 $Y=307120
X3079 1 2 171 125 1149 ICV_69 $T=304520 307360 0 0 $X=304330 $Y=307120
X3080 1 2 1180 128 1224 ICV_69 $T=347300 285600 1 0 $X=347110 $Y=282640
X3081 1 2 1231 210 1257 ICV_69 $T=365240 301920 1 0 $X=365050 $Y=298960
X3082 1 2 1258 217 1278 ICV_69 $T=374900 296480 1 0 $X=374710 $Y=293520
X3083 1 2 1247 232 1298 ICV_69 $T=388700 280160 0 0 $X=388510 $Y=279920
X3084 1 2 1338 251 1364 ICV_69 $T=417220 274720 0 0 $X=417030 $Y=274480
X3085 1 2 1454 232 1477 ICV_69 $T=472880 285600 0 0 $X=472690 $Y=285360
X3086 1 2 1491 216 1506 ICV_69 $T=487140 301920 1 0 $X=486950 $Y=298960
X3087 1 2 177 348 1503 ICV_69 $T=487600 285600 1 0 $X=487410 $Y=282640
X3088 1 2 1521 367 1549 ICV_69 $T=508300 280160 1 0 $X=508110 $Y=277200
X3089 1 2 409 399 1623 ICV_69 $T=546480 307360 0 0 $X=546290 $Y=307120
X3090 1 2 1659 227 1676 ICV_69 $T=574540 280160 0 0 $X=574350 $Y=279920
X3091 1 2 1659 224 1702 ICV_69 $T=585120 280160 0 0 $X=584930 $Y=279920
X3092 1 2 1690 401 1699 ICV_69 $T=587880 301920 1 0 $X=587690 $Y=298960
X3093 1 2 1672 253 1698 ICV_69 $T=588800 258400 1 0 $X=588610 $Y=255440
X3094 1 2 1738 390 1758 ICV_69 $T=611800 312800 1 0 $X=611610 $Y=309840
X3095 1 2 1846 357 1874 ICV_69 $T=669760 252960 0 0 $X=669570 $Y=252720
X3096 1 2 1886 358 1924 ICV_69 $T=697360 280160 0 0 $X=697170 $Y=279920
X3097 1 2 40 7 583 583 582 105 ICV_74 $T=36340 285600 1 0 $X=36150 $Y=282640
X3098 1 2 58 7 644 644 62 105 ICV_74 $T=62560 301920 0 0 $X=62370 $Y=301680
X3099 1 2 72 7 695 695 670 105 ICV_74 $T=90160 258400 0 0 $X=89970 $Y=258160
X3100 1 2 20 107 852 852 861 105 ICV_74 $T=163300 269280 0 0 $X=163110 $Y=269040
X3101 1 2 44 107 898 138 137 105 ICV_74 $T=187220 301920 0 0 $X=187030 $Y=301680
X3102 1 2 57 107 907 907 919 105 ICV_74 $T=192740 274720 0 0 $X=192550 $Y=274480
X3103 1 2 72 107 1047 1047 1054 105 ICV_74 $T=258980 258400 0 0 $X=258790 $Y=258160
X3104 1 2 73 107 1067 1067 1070 105 ICV_74 $T=270480 301920 0 0 $X=270290 $Y=301680
X3105 1 2 98 107 1140 1140 1129 105 ICV_74 $T=304060 263840 0 0 $X=303870 $Y=263600
X3106 1 2 297 215 1345 1345 1338 239 ICV_74 $T=413540 269280 1 0 $X=413350 $Y=266320
X3107 1 2 269 351 1597 1597 1601 239 ICV_74 $T=539580 280160 0 0 $X=539390 $Y=279920
X3108 1 2 281 351 1581 1608 1617 239 ICV_74 $T=543260 263840 0 0 $X=543070 $Y=263600
X3109 1 2 433 215 1744 1744 1763 239 ICV_74 $T=614560 269280 1 0 $X=614370 $Y=266320
X3110 1 2 315 366 1819 1819 1820 479 ICV_74 $T=647220 307360 1 0 $X=647030 $Y=304400
X3111 1 2 433 351 1845 1845 1848 239 ICV_74 $T=660100 280160 0 0 $X=659910 $Y=279920
X3112 1 2 443 351 1932 1932 1944 239 ICV_74 $T=707020 285600 1 0 $X=706830 $Y=282640
X3113 1 2 442 351 1937 1937 1943 239 ICV_74 $T=707480 274720 0 0 $X=707290 $Y=274480
X3114 1 2 439 351 1942 1942 1951 239 ICV_74 $T=710240 258400 1 0 $X=710050 $Y=255440
X3115 1 2 581 25 610 ICV_76 $T=46460 296480 1 0 $X=46270 $Y=293520
X3116 1 2 664 11 671 ICV_76 $T=74520 269280 1 0 $X=74330 $Y=266320
X3117 1 2 618 11 681 ICV_76 $T=74520 301920 1 0 $X=74330 $Y=298960
X3118 1 2 899 111 934 ICV_76 $T=200560 291040 0 0 $X=200370 $Y=290800
X3119 1 2 1176 112 1192 ICV_76 $T=327060 258400 1 0 $X=326870 $Y=255440
X3120 1 2 1230 224 1265 ICV_76 $T=368920 269280 0 0 $X=368730 $Y=269040
X3121 1 2 1292 216 1324 ICV_76 $T=396980 291040 0 0 $X=396790 $Y=290800
X3122 1 2 1292 213 1295 ICV_76 $T=396980 296480 0 0 $X=396790 $Y=296240
X3123 1 2 1418 223 1443 ICV_76 $T=453100 274720 0 0 $X=452910 $Y=274480
X3124 1 2 1513 359 1525 ICV_76 $T=495420 258400 1 0 $X=495230 $Y=255440
X3125 1 2 379 388 1579 ICV_76 $T=523480 307360 1 0 $X=523290 $Y=304400
X3126 1 2 1572 364 1600 ICV_76 $T=537280 291040 0 0 $X=537090 $Y=290800
X3127 1 2 393 357 1632 ICV_76 $T=551540 247520 1 0 $X=551350 $Y=244560
X3128 1 2 1630 368 1664 ICV_76 $T=565340 291040 0 0 $X=565150 $Y=290800
X3129 1 2 1672 224 1710 ICV_76 $T=593400 263840 0 0 $X=593210 $Y=263600
X3130 1 2 1738 404 1777 ICV_76 $T=621460 296480 0 0 $X=621270 $Y=296240
X3131 1 2 1873 401 1889 ICV_76 $T=677580 301920 0 0 $X=677390 $Y=301680
X3132 1 2 1900 364 1914 ICV_76 $T=691840 263840 1 0 $X=691650 $Y=260880
X3133 1 2 524 5 537 537 543 16 4 536 536 543 17 ICV_77 $T=7360 301920 1 0 $X=7170 $Y=298960
X3134 1 2 522 26 564 564 542 34 25 563 563 542 30 ICV_77 $T=21160 263840 1 0 $X=20970 $Y=260880
X3135 1 2 530 14 568 568 555 19 25 567 567 555 30 ICV_77 $T=21160 291040 1 0 $X=20970 $Y=288080
X3136 1 2 530 26 574 574 555 34 24 573 573 555 33 ICV_77 $T=21620 296480 1 0 $X=21430 $Y=293520
X3137 1 2 524 26 576 558 543 19 24 575 575 543 33 ICV_77 $T=22080 301920 1 0 $X=21890 $Y=298960
X3138 1 2 582 14 594 594 602 19 25 593 593 602 30 ICV_77 $T=34040 280160 1 0 $X=33850 $Y=277200
X3139 1 2 581 11 601 600 585 34 26 600 547 555 13 ICV_77 $T=34960 296480 1 0 $X=34770 $Y=293520
X3140 1 2 708 5 743 727 740 17 24 742 742 740 33 ICV_77 $T=106260 291040 1 0 $X=106070 $Y=288080
X3141 1 2 859 125 913 913 863 135 128 912 911 863 134 ICV_77 $T=189980 258400 1 0 $X=189790 $Y=255440
X3142 1 2 927 112 937 937 933 123 110 936 936 933 122 ICV_77 $T=202860 258400 1 0 $X=202670 $Y=255440
X3143 1 2 1070 125 1112 1112 1086 135 126 1111 1111 1086 136 ICV_77 $T=286580 296480 1 0 $X=286390 $Y=293520
X3144 1 2 1459 224 1473 1473 1470 233 238 1469 1475 1470 262 ICV_77 $T=471040 258400 1 0 $X=470850 $Y=255440
X3145 1 2 1514 357 1529 1529 1532 348 356 1528 1528 1532 337 ICV_77 $T=497260 291040 1 0 $X=497070 $Y=288080
X3146 1 2 1570 363 1605 1605 1576 303 357 1604 1604 1576 348 ICV_77 $T=539580 258400 1 0 $X=539390 $Y=255440
X3147 1 2 1677 357 1696 1696 1685 348 359 1695 1695 1685 341 ICV_77 $T=582360 291040 1 0 $X=582170 $Y=288080
X3148 1 2 1708 238 1719 1719 1723 201 251 1718 1718 1723 263 ICV_77 $T=596160 274720 1 0 $X=595970 $Y=271760
X3149 1 2 1734 359 1746 1746 1739 341 367 1745 1745 1739 306 ICV_77 $T=609500 285600 1 0 $X=609310 $Y=282640
X3150 1 2 1791 251 1810 1795 1802 263 227 1809 1809 1812 252 ICV_77 $T=638940 258400 1 0 $X=638750 $Y=255440
X3151 1 2 1789 357 1835 1835 1804 348 359 1834 1834 1804 341 ICV_77 $T=651820 291040 1 0 $X=651630 $Y=288080
X3152 1 2 1847 356 1895 1895 1853 337 357 1894 1894 1853 348 ICV_77 $T=680340 263840 1 0 $X=680150 $Y=260880
X3153 1 2 198 200 61 203 1191 205 2 209 1 sky130_fd_sc_hd__mux4_1 $T=330280 247520 1 0 $X=330090 $Y=244560
X3154 1 2 226 228 61 234 1222 205 2 241 1 sky130_fd_sc_hd__mux4_1 $T=347300 269280 0 0 $X=347110 $Y=269040
X3155 1 2 279 282 61 285 1318 205 2 290 1 sky130_fd_sc_hd__mux4_1 $T=397440 285600 1 0 $X=397250 $Y=282640
X3156 1 2 287 288 61 292 1332 205 2 296 1 sky130_fd_sc_hd__mux4_1 $T=403880 285600 0 0 $X=403690 $Y=285360
X3157 1 2 304 305 61 308 1378 205 2 310 1 sky130_fd_sc_hd__mux4_1 $T=426880 285600 0 0 $X=426690 $Y=285360
X3158 1 2 320 321 61 323 1440 205 2 325 1 sky130_fd_sc_hd__mux4_1 $T=455860 285600 0 0 $X=455670 $Y=285360
X3159 1 2 330 333 61 335 1463 205 2 338 1 sky130_fd_sc_hd__mux4_1 $T=469200 291040 1 0 $X=469010 $Y=288080
X3160 1 2 346 349 61 352 1503 205 2 354 1 sky130_fd_sc_hd__mux4_1 $T=488060 285600 0 0 $X=487870 $Y=285360
X3161 1 2 371 374 61 377 1554 205 2 383 1 sky130_fd_sc_hd__mux4_1 $T=512900 296480 1 0 $X=512710 $Y=293520
X3162 1 2 386 387 61 392 1573 205 2 398 1 sky130_fd_sc_hd__mux4_1 $T=525320 296480 1 0 $X=525130 $Y=293520
.ENDS
***************************************
.SUBCKT ICV_79 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380
+ 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400
+ 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420
+ 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440
+ 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460
+ 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480
+ 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500
+ 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520
+ 521 522 523 524 525 526 527
** N=1980 EP=527 IP=15906 FDC=47715
*.SEEDPROM
X0 1 2 Dpar a=2091.2 p=1484.64 m=1 $[nwdiode] $X=5330 $Y=183545 $D=191
X1 1 2 Dpar a=2090.63 p=1485.34 m=1 $[nwdiode] $X=5330 $Y=188985 $D=191
X2 1 2 Dpar a=2091.2 p=1484.64 m=1 $[nwdiode] $X=5330 $Y=194425 $D=191
X3 1 2 Dpar a=2090.3 p=1485.74 m=1 $[nwdiode] $X=5330 $Y=199865 $D=191
X4 1 2 Dpar a=2091.12 p=1484.74 m=1 $[nwdiode] $X=5330 $Y=205305 $D=191
X5 1 2 Dpar a=2090.95 p=1484.94 m=1 $[nwdiode] $X=5330 $Y=210745 $D=191
X6 1 2 Dpar a=2091.44 p=1484.34 m=1 $[nwdiode] $X=5330 $Y=216185 $D=191
X7 1 2 Dpar a=2090.95 p=1484.94 m=1 $[nwdiode] $X=5330 $Y=221625 $D=191
X8 1 2 Dpar a=2090.71 p=1485.24 m=1 $[nwdiode] $X=5330 $Y=227065 $D=191
X9 1 2 Dpar a=2091.6 p=1484.14 m=1 $[nwdiode] $X=5330 $Y=232505 $D=191
X10 1 2 Dpar a=2090.71 p=1485.24 m=1 $[nwdiode] $X=5330 $Y=237945 $D=191
X11 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=17940 198560 0 0 $X=17750 $Y=198320
X12 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=18400 198560 1 0 $X=18210 $Y=195600
X13 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=27600 198560 0 0 $X=27410 $Y=198320
X14 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=48300 242080 0 0 $X=48110 $Y=241840
X15 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=81880 242080 0 0 $X=81690 $Y=241840
X16 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=82340 187680 0 0 $X=82150 $Y=187440
X17 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=84180 204000 1 0 $X=83990 $Y=201040
X18 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=87860 236640 1 0 $X=87670 $Y=233680
X19 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=98440 214880 1 0 $X=98250 $Y=211920
X20 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=121900 242080 1 0 $X=121710 $Y=239120
X21 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=141680 214880 1 0 $X=141490 $Y=211920
X22 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=153640 231200 0 0 $X=153450 $Y=230960
X23 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=154560 220320 0 0 $X=154370 $Y=220080
X24 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=158700 193120 1 0 $X=158510 $Y=190160
X25 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=160540 220320 1 0 $X=160350 $Y=217360
X26 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=168360 204000 0 0 $X=168170 $Y=203760
X27 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=183540 204000 0 0 $X=183350 $Y=203760
X28 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=202400 220320 0 0 $X=202210 $Y=220080
X29 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=228620 214880 0 0 $X=228430 $Y=214640
X30 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=244720 242080 1 0 $X=244530 $Y=239120
X31 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=252540 214880 1 0 $X=252350 $Y=211920
X32 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=258520 236640 0 0 $X=258330 $Y=236400
X33 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=268180 214880 0 0 $X=267990 $Y=214640
X34 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=271400 236640 0 0 $X=271210 $Y=236400
X35 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=272780 182240 1 0 $X=272590 $Y=179280
X36 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=295780 187680 0 0 $X=295590 $Y=187440
X37 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=311420 193120 0 0 $X=311230 $Y=192880
X38 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=312800 198560 0 0 $X=312610 $Y=198320
X39 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=314180 242080 1 0 $X=313990 $Y=239120
X40 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=314640 187680 0 0 $X=314450 $Y=187440
X41 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=327520 225760 0 0 $X=327330 $Y=225520
X42 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=331200 209440 0 0 $X=331010 $Y=209200
X43 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=340860 209440 0 0 $X=340670 $Y=209200
X44 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=340860 214880 0 0 $X=340670 $Y=214640
X45 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=370760 182240 0 0 $X=370570 $Y=182000
X46 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=388240 193120 0 0 $X=388050 $Y=192880
X47 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=413080 220320 1 0 $X=412890 $Y=217360
X48 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=419520 204000 1 0 $X=419330 $Y=201040
X49 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=453100 182240 0 0 $X=452910 $Y=182000
X50 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=453100 193120 0 0 $X=452910 $Y=192880
X51 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=457240 242080 0 0 $X=457050 $Y=241840
X52 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=463220 236640 1 0 $X=463030 $Y=233680
X53 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=469200 187680 1 0 $X=469010 $Y=184720
X54 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=480700 220320 1 0 $X=480510 $Y=217360
X55 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=481160 193120 0 0 $X=480970 $Y=192880
X56 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=483920 236640 1 0 $X=483730 $Y=233680
X57 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=509220 225760 0 0 $X=509030 $Y=225520
X58 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=509220 236640 0 0 $X=509030 $Y=236400
X59 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=510140 204000 1 0 $X=509950 $Y=201040
X60 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=511980 209440 1 0 $X=511790 $Y=206480
X61 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=551540 193120 1 0 $X=551350 $Y=190160
X62 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=565340 220320 0 0 $X=565150 $Y=220080
X63 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=576380 225760 1 0 $X=576190 $Y=222800
X64 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=593400 236640 0 0 $X=593210 $Y=236400
X65 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=609500 236640 1 0 $X=609310 $Y=233680
X66 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=613640 214880 0 0 $X=613450 $Y=214640
X67 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=621460 214880 0 0 $X=621270 $Y=214640
X68 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=649980 231200 1 0 $X=649790 $Y=228240
X69 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=654120 198560 1 0 $X=653930 $Y=195600
X70 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=662860 187680 0 0 $X=662670 $Y=187440
X71 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=663780 204000 1 0 $X=663590 $Y=201040
X72 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=663780 209440 1 0 $X=663590 $Y=206480
X73 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=673900 193120 1 0 $X=673710 $Y=190160
X74 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=679420 209440 0 0 $X=679230 $Y=209200
X75 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=693680 214880 1 0 $X=693490 $Y=211920
X76 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=696440 236640 0 0 $X=696250 $Y=236400
X77 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=707480 220320 0 0 $X=707290 $Y=220080
X78 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=707480 236640 0 0 $X=707290 $Y=236400
X79 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=719900 187680 1 0 $X=719710 $Y=184720
X80 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=721740 225760 1 0 $X=721550 $Y=222800
X81 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=735540 225760 0 0 $X=735350 $Y=225520
X82 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=735540 242080 0 0 $X=735350 $Y=241840
X83 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=741520 225760 1 0 $X=741330 $Y=222800
X84 1 2 ICV_1 $T=744280 214880 0 180 $X=742710 $Y=211920
X85 1 2 ICV_1 $T=744280 242080 0 180 $X=742710 $Y=239120
X86 1 2 ICV_2 $T=5520 182240 1 0 $X=5330 $Y=179280
X87 1 2 ICV_2 $T=5520 193120 1 0 $X=5330 $Y=190160
X88 1 2 ICV_2 $T=5520 204000 1 0 $X=5330 $Y=201040
X89 1 2 ICV_2 $T=5520 214880 1 0 $X=5330 $Y=211920
X90 1 2 ICV_2 $T=5520 225760 1 0 $X=5330 $Y=222800
X91 1 2 ICV_2 $T=5520 236640 1 0 $X=5330 $Y=233680
X92 1 2 ICV_2 $T=744280 182240 0 180 $X=742710 $Y=179280
X93 1 2 ICV_2 $T=744280 193120 0 180 $X=742710 $Y=190160
X94 1 2 ICV_2 $T=744280 204000 0 180 $X=742710 $Y=201040
X95 1 2 ICV_2 $T=744280 220320 0 180 $X=742710 $Y=217360
X96 1 2 ICV_2 $T=744280 231200 0 180 $X=742710 $Y=228240
X229 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 209440 1 0 $X=17750 $Y=206480
X230 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=20240 225760 1 0 $X=20050 $Y=222800
X231 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=34040 225760 0 0 $X=33850 $Y=225520
X232 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=38180 209440 0 0 $X=37990 $Y=209200
X233 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=62100 204000 0 0 $X=61910 $Y=203760
X234 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=69920 182240 1 0 $X=69730 $Y=179280
X235 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=74060 187680 0 0 $X=73870 $Y=187440
X236 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=76360 193120 1 0 $X=76170 $Y=190160
X237 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=79120 209440 0 0 $X=78930 $Y=209200
X238 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=80040 236640 0 0 $X=79850 $Y=236400
X239 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=87860 198560 0 0 $X=87670 $Y=198320
X240 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=122360 220320 0 0 $X=122170 $Y=220080
X241 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=135240 242080 0 0 $X=135050 $Y=241840
X242 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=139840 204000 1 0 $X=139650 $Y=201040
X243 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=150420 204000 0 0 $X=150230 $Y=203760
X244 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=154100 209440 0 0 $X=153910 $Y=209200
X245 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=158240 231200 1 0 $X=158050 $Y=228240
X246 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=181700 193120 0 0 $X=181510 $Y=192880
X247 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=210680 231200 0 0 $X=210490 $Y=230960
X248 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=216660 231200 1 0 $X=216470 $Y=228240
X249 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=228160 204000 1 0 $X=227970 $Y=201040
X250 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=248860 242080 0 0 $X=248670 $Y=241840
X251 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=256220 182240 0 0 $X=256030 $Y=182000
X252 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=258520 193120 0 0 $X=258330 $Y=192880
X253 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=260820 209440 1 0 $X=260630 $Y=206480
X254 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=262660 182240 0 0 $X=262470 $Y=182000
X255 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=293940 209440 0 0 $X=293750 $Y=209200
X256 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=298540 220320 1 0 $X=298350 $Y=217360
X257 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=298540 231200 1 0 $X=298350 $Y=228240
X258 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=326600 220320 1 0 $X=326410 $Y=217360
X259 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=328900 182240 1 0 $X=328710 $Y=179280
X260 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=354660 225760 1 0 $X=354470 $Y=222800
X261 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=361100 198560 1 0 $X=360910 $Y=195600
X262 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=361100 214880 1 0 $X=360910 $Y=211920
X263 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=389160 204000 1 0 $X=388970 $Y=201040
X264 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=398820 220320 0 0 $X=398630 $Y=220080
X265 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=406180 225760 0 0 $X=405990 $Y=225520
X266 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=408020 193120 0 0 $X=407830 $Y=192880
X267 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=409400 182240 0 0 $X=409210 $Y=182000
X268 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=420440 182240 0 0 $X=420250 $Y=182000
X269 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=426880 236640 0 0 $X=426690 $Y=236400
X270 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=435160 242080 0 0 $X=434970 $Y=241840
X271 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=446200 198560 0 0 $X=446010 $Y=198320
X272 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=446200 231200 0 0 $X=446010 $Y=230960
X273 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=448500 242080 1 0 $X=448310 $Y=239120
X274 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=454940 236640 0 0 $X=454750 $Y=236400
X275 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=470580 182240 0 0 $X=470390 $Y=182000
X276 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=490360 198560 0 0 $X=490170 $Y=198320
X277 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=491740 214880 0 0 $X=491550 $Y=214640
X278 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=523020 242080 1 0 $X=522830 $Y=239120
X279 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=525320 187680 1 0 $X=525130 $Y=184720
X280 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=546480 193120 0 0 $X=546290 $Y=192880
X281 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=553380 214880 1 0 $X=553190 $Y=211920
X282 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=587880 214880 0 0 $X=587690 $Y=214640
X283 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=658720 198560 0 0 $X=658530 $Y=198320
X284 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=665620 182240 1 0 $X=665430 $Y=179280
X285 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=681260 242080 1 0 $X=681070 $Y=239120
X286 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=693680 242080 1 0 $X=693490 $Y=239120
X287 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=711620 182240 0 0 $X=711430 $Y=182000
X288 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=735540 231200 0 0 $X=735350 $Y=230960
X289 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 231200 1 0 $X=740870 $Y=228240
X290 1 2 ICV_3 $T=13340 236640 0 0 $X=13150 $Y=236400
X291 1 2 ICV_3 $T=31280 193120 0 0 $X=31090 $Y=192880
X292 1 2 ICV_3 $T=62100 198560 0 0 $X=61910 $Y=198320
X293 1 2 ICV_3 $T=63020 225760 1 0 $X=62830 $Y=222800
X294 1 2 ICV_3 $T=69460 225760 1 0 $X=69270 $Y=222800
X295 1 2 ICV_3 $T=83720 231200 1 0 $X=83530 $Y=228240
X296 1 2 ICV_3 $T=125580 236640 1 0 $X=125390 $Y=233680
X297 1 2 ICV_3 $T=143520 236640 0 0 $X=143330 $Y=236400
X298 1 2 ICV_3 $T=161920 242080 0 0 $X=161730 $Y=241840
X299 1 2 ICV_3 $T=185840 242080 0 0 $X=185650 $Y=241840
X300 1 2 ICV_3 $T=188600 193120 1 0 $X=188410 $Y=190160
X301 1 2 ICV_3 $T=236440 236640 1 0 $X=236250 $Y=233680
X302 1 2 ICV_3 $T=241960 220320 1 0 $X=241770 $Y=217360
X303 1 2 ICV_3 $T=304980 231200 1 0 $X=304790 $Y=228240
X304 1 2 ICV_3 $T=311880 209440 0 0 $X=311690 $Y=209200
X305 1 2 ICV_3 $T=318780 236640 0 0 $X=318590 $Y=236400
X306 1 2 ICV_3 $T=338100 204000 1 0 $X=337910 $Y=201040
X307 1 2 ICV_3 $T=356960 193120 1 0 $X=356770 $Y=190160
X308 1 2 ICV_3 $T=363860 209440 0 0 $X=363670 $Y=209200
X309 1 2 ICV_3 $T=392380 209440 1 0 $X=392190 $Y=206480
X310 1 2 ICV_3 $T=397440 187680 1 0 $X=397250 $Y=184720
X311 1 2 ICV_3 $T=406180 198560 1 0 $X=405990 $Y=195600
X312 1 2 ICV_3 $T=424120 198560 0 0 $X=423930 $Y=198320
X313 1 2 ICV_3 $T=431940 231200 1 0 $X=431750 $Y=228240
X314 1 2 ICV_3 $T=438380 242080 1 0 $X=438190 $Y=239120
X315 1 2 ICV_3 $T=448040 220320 0 0 $X=447850 $Y=220080
X316 1 2 ICV_3 $T=452180 231200 0 0 $X=451990 $Y=230960
X317 1 2 ICV_3 $T=504160 182240 0 0 $X=503970 $Y=182000
X318 1 2 ICV_3 $T=511060 214880 0 0 $X=510870 $Y=214640
X319 1 2 ICV_3 $T=518420 182240 0 0 $X=518230 $Y=182000
X320 1 2 ICV_3 $T=531760 231200 0 0 $X=531570 $Y=230960
X321 1 2 ICV_3 $T=536360 182240 0 0 $X=536170 $Y=182000
X322 1 2 ICV_3 $T=567180 187680 0 0 $X=566990 $Y=187440
X323 1 2 ICV_3 $T=585580 187680 1 0 $X=585390 $Y=184720
X324 1 2 ICV_3 $T=587420 182240 0 0 $X=587230 $Y=182000
X325 1 2 ICV_3 $T=587880 225760 1 0 $X=587690 $Y=222800
X326 1 2 ICV_3 $T=592480 242080 0 0 $X=592290 $Y=241840
X327 1 2 ICV_3 $T=623300 187680 0 0 $X=623110 $Y=187440
X328 1 2 ICV_3 $T=644000 236640 0 0 $X=643810 $Y=236400
X329 1 2 ICV_3 $T=651360 182240 0 0 $X=651170 $Y=182000
X330 1 2 ICV_3 $T=665620 231200 1 0 $X=665430 $Y=228240
X331 1 2 ICV_3 $T=679420 187680 0 0 $X=679230 $Y=187440
X332 1 2 ICV_3 $T=700580 242080 0 0 $X=700390 $Y=241840
X333 1 2 ICV_3 $T=719900 182240 0 0 $X=719710 $Y=182000
X334 1 2 ICV_3 $T=735540 182240 0 0 $X=735350 $Y=182000
X335 1 2 ICV_3 $T=735540 214880 0 0 $X=735350 $Y=214640
X336 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=12420 193120 1 0 $X=12230 $Y=190160
X337 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=16100 231200 0 0 $X=15910 $Y=230960
X338 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=20240 204000 0 0 $X=20050 $Y=203760
X339 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=28060 209440 1 0 $X=27870 $Y=206480
X340 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=58880 209440 0 0 $X=58690 $Y=209200
X341 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=97520 242080 0 0 $X=97330 $Y=241840
X342 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=98900 214880 0 0 $X=98710 $Y=214640
X343 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=124660 204000 1 0 $X=124470 $Y=201040
X344 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=139840 209440 1 0 $X=139650 $Y=206480
X345 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=140300 236640 1 0 $X=140110 $Y=233680
X346 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=146280 193120 0 0 $X=146090 $Y=192880
X347 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=146280 242080 0 0 $X=146090 $Y=241840
X348 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=160540 187680 0 0 $X=160350 $Y=187440
X349 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=169740 225760 1 0 $X=169550 $Y=222800
X350 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=184920 209440 0 0 $X=184730 $Y=209200
X351 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=188600 182240 1 0 $X=188410 $Y=179280
X352 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=269560 204000 1 0 $X=269370 $Y=201040
X353 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=286580 193120 0 0 $X=286390 $Y=192880
X354 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=300840 214880 1 0 $X=300650 $Y=211920
X355 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=300840 236640 1 0 $X=300650 $Y=233680
X356 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=311420 182240 0 0 $X=311230 $Y=182000
X357 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=311420 225760 0 0 $X=311230 $Y=225520
X358 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=328900 242080 1 0 $X=328710 $Y=239120
X359 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=339480 236640 0 0 $X=339290 $Y=236400
X360 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=353740 209440 1 0 $X=353550 $Y=206480
X361 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=353740 231200 1 0 $X=353550 $Y=228240
X362 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=361100 204000 1 0 $X=360910 $Y=201040
X363 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=367540 214880 0 0 $X=367350 $Y=214640
X364 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=370760 214880 0 0 $X=370570 $Y=214640
X365 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=395600 209440 0 0 $X=395410 $Y=209200
X366 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=395600 220320 0 0 $X=395410 $Y=220080
X367 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=437920 204000 1 0 $X=437730 $Y=201040
X368 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=437920 209440 1 0 $X=437730 $Y=206480
X369 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=441140 187680 1 0 $X=440950 $Y=184720
X370 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=451720 242080 0 0 $X=451530 $Y=241840
X371 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=476560 209440 1 0 $X=476370 $Y=206480
X372 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=494040 209440 1 0 $X=493850 $Y=206480
X373 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=525320 214880 1 0 $X=525130 $Y=211920
X374 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=573620 231200 1 0 $X=573430 $Y=228240
X375 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=634340 242080 1 0 $X=634150 $Y=239120
X376 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=642620 182240 0 0 $X=642430 $Y=182000
X377 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=657800 231200 1 0 $X=657610 $Y=228240
X378 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=676660 214880 1 0 $X=676470 $Y=211920
X379 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=714380 220320 1 0 $X=714190 $Y=217360
X380 1 2 ICV_4 $T=118220 204000 0 0 $X=118030 $Y=203760
X381 1 2 ICV_4 $T=226320 220320 1 0 $X=226130 $Y=217360
X382 1 2 ICV_4 $T=269560 204000 0 0 $X=269370 $Y=203760
X383 1 2 ICV_4 $T=316020 236640 1 0 $X=315830 $Y=233680
X384 1 2 ICV_4 $T=367080 204000 0 0 $X=366890 $Y=203760
X385 1 2 ICV_4 $T=367080 231200 0 0 $X=366890 $Y=230960
X386 1 2 ICV_4 $T=518420 225760 0 0 $X=518230 $Y=225520
X387 1 2 ICV_4 $T=535440 236640 0 0 $X=535250 $Y=236400
X388 1 2 ICV_4 $T=536820 220320 1 0 $X=536630 $Y=217360
X389 1 2 ICV_4 $T=563500 242080 0 0 $X=563310 $Y=241840
X390 1 2 ICV_4 $T=567180 193120 0 0 $X=566990 $Y=192880
X391 1 2 ICV_4 $T=581440 204000 1 0 $X=581250 $Y=201040
X392 1 2 ICV_4 $T=595240 198560 0 0 $X=595050 $Y=198320
X393 1 2 ICV_4 $T=605820 220320 1 0 $X=605630 $Y=217360
X394 1 2 ICV_4 $T=708860 209440 1 0 $X=708670 $Y=206480
X395 1 2 ICV_4 $T=739680 220320 0 0 $X=739490 $Y=220080
X396 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 182240 1 0 $X=6710 $Y=179280
X397 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 182240 0 0 $X=6710 $Y=182000
X398 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 193120 0 0 $X=6710 $Y=192880
X399 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 198560 1 0 $X=6710 $Y=195600
X400 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 209440 0 0 $X=6710 $Y=209200
X401 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 214880 1 0 $X=6710 $Y=211920
X402 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 214880 0 0 $X=6710 $Y=214640
X403 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 220320 1 0 $X=6710 $Y=217360
X404 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=16100 236640 1 0 $X=15910 $Y=233680
X405 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=34040 231200 0 0 $X=33850 $Y=230960
X406 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=68080 204000 1 0 $X=67890 $Y=201040
X407 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=70380 225760 0 0 $X=70190 $Y=225520
X408 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=94300 198560 0 0 $X=94110 $Y=198320
X409 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=95220 231200 1 0 $X=95030 $Y=228240
X410 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=104420 242080 1 0 $X=104230 $Y=239120
X411 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=114080 220320 0 0 $X=113890 $Y=220080
X412 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=129720 187680 0 0 $X=129530 $Y=187440
X413 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=129720 225760 0 0 $X=129530 $Y=225520
X414 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=132480 187680 1 0 $X=132290 $Y=184720
X415 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=142140 204000 0 0 $X=141950 $Y=203760
X416 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=164680 231200 1 0 $X=164490 $Y=228240
X417 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=168360 204000 1 0 $X=168170 $Y=201040
X418 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=170200 182240 0 0 $X=170010 $Y=182000
X419 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=173880 214880 1 0 $X=173690 $Y=211920
X420 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=174340 198560 0 0 $X=174150 $Y=198320
X421 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=174340 220320 0 0 $X=174150 $Y=220080
X422 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=177100 236640 1 0 $X=176910 $Y=233680
X423 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=178480 214880 0 0 $X=178290 $Y=214640
X424 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=183080 220320 1 0 $X=182890 $Y=217360
X425 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=184460 187680 1 0 $X=184270 $Y=184720
X426 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=188600 198560 1 0 $X=188410 $Y=195600
X427 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=189060 231200 0 0 $X=188870 $Y=230960
X428 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=197800 220320 0 0 $X=197610 $Y=220080
X429 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=198260 187680 0 0 $X=198070 $Y=187440
X430 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=200100 214880 1 0 $X=199910 $Y=211920
X431 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=207920 225760 0 0 $X=207730 $Y=225520
X432 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=210220 209440 0 0 $X=210030 $Y=209200
X433 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=211140 204000 1 0 $X=210950 $Y=201040
X434 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=226320 182240 0 0 $X=226130 $Y=182000
X435 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=234600 225760 0 0 $X=234410 $Y=225520
X436 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=240120 225760 1 0 $X=239930 $Y=222800
X437 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=244720 182240 1 0 $X=244530 $Y=179280
X438 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=258060 214880 1 0 $X=257870 $Y=211920
X439 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=268640 225760 1 0 $X=268450 $Y=222800
X440 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=271400 225760 0 0 $X=271210 $Y=225520
X441 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=272780 198560 1 0 $X=272590 $Y=195600
X442 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=278300 193120 0 0 $X=278110 $Y=192880
X443 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=282440 236640 0 0 $X=282250 $Y=236400
X444 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=303140 242080 0 0 $X=302950 $Y=241840
X445 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=310960 225760 1 0 $X=310770 $Y=222800
X446 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=318780 193120 0 0 $X=318590 $Y=192880
X447 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=324300 225760 1 0 $X=324110 $Y=222800
X448 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=328900 214880 1 0 $X=328710 $Y=211920
X449 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=336260 220320 1 0 $X=336070 $Y=217360
X450 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=337640 231200 0 0 $X=337450 $Y=230960
X451 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=342700 204000 0 0 $X=342510 $Y=203760
X452 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=375360 193120 0 0 $X=375170 $Y=192880
X453 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=378120 242080 0 0 $X=377930 $Y=241840
X454 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=385020 214880 1 0 $X=384830 $Y=211920
X455 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=385020 220320 1 0 $X=384830 $Y=217360
X456 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=390540 214880 0 0 $X=390350 $Y=214640
X457 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=414000 193120 0 0 $X=413810 $Y=192880
X458 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=415380 220320 0 0 $X=415190 $Y=220080
X459 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=434240 198560 0 0 $X=434050 $Y=198320
X460 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=459080 198560 1 0 $X=458890 $Y=195600
X461 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=476560 193120 1 0 $X=476370 $Y=190160
X462 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=505540 225760 0 0 $X=505350 $Y=225520
X463 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=511060 182240 1 0 $X=510870 $Y=179280
X464 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=520260 214880 0 0 $X=520070 $Y=214640
X465 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=520720 204000 1 0 $X=520530 $Y=201040
X466 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=525320 204000 1 0 $X=525130 $Y=201040
X467 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=525320 209440 1 0 $X=525130 $Y=206480
X468 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=531760 242080 1 0 $X=531570 $Y=239120
X469 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=536820 236640 1 0 $X=536630 $Y=233680
X470 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=543260 242080 0 0 $X=543070 $Y=241840
X471 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=552920 204000 0 0 $X=552730 $Y=203760
X472 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=554300 214880 0 0 $X=554110 $Y=214640
X473 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=557520 193120 1 0 $X=557330 $Y=190160
X474 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=568560 198560 1 0 $X=568370 $Y=195600
X475 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=570860 182240 1 0 $X=570670 $Y=179280
X476 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=572700 225760 1 0 $X=572510 $Y=222800
X477 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=595240 204000 0 0 $X=595050 $Y=203760
X478 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=606740 225760 0 0 $X=606550 $Y=225520
X479 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=609960 214880 0 0 $X=609770 $Y=214640
X480 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=616860 220320 1 0 $X=616670 $Y=217360
X481 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=628820 220320 0 0 $X=628630 $Y=220080
X482 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=650440 198560 1 0 $X=650250 $Y=195600
X483 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=651820 236640 1 0 $X=651630 $Y=233680
X484 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=661020 198560 1 0 $X=660830 $Y=195600
X485 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=665620 193120 1 0 $X=665430 $Y=190160
X486 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=674360 209440 0 0 $X=674170 $Y=209200
X487 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=674820 187680 0 0 $X=674630 $Y=187440
X488 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=674820 236640 1 0 $X=674630 $Y=233680
X489 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=679420 242080 0 0 $X=679230 $Y=241840
X490 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=701040 198560 1 0 $X=700850 $Y=195600
X491 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=703340 193120 0 0 $X=703150 $Y=192880
X492 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=714840 193120 0 0 $X=714650 $Y=192880
X493 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 187680 1 0 $X=6710 $Y=184720
X494 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 187680 0 0 $X=6710 $Y=187440
X495 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 193120 1 0 $X=6710 $Y=190160
X496 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 198560 0 0 $X=6710 $Y=198320
X497 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 204000 1 0 $X=6710 $Y=201040
X498 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 204000 0 0 $X=6710 $Y=203760
X499 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 209440 1 0 $X=6710 $Y=206480
X500 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 220320 0 0 $X=6710 $Y=220080
X501 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 225760 1 0 $X=6710 $Y=222800
X502 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 225760 0 0 $X=6710 $Y=225520
X503 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 231200 1 0 $X=6710 $Y=228240
X504 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=12420 198560 0 0 $X=12230 $Y=198320
X505 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=12420 209440 1 0 $X=12230 $Y=206480
X506 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=12420 220320 0 0 $X=12230 $Y=220080
X507 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=12420 225760 1 0 $X=12230 $Y=222800
X508 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=12420 225760 0 0 $X=12230 $Y=225520
X509 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=12420 231200 1 0 $X=12230 $Y=228240
X510 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=17940 225760 0 0 $X=17750 $Y=225520
X511 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=20240 231200 1 0 $X=20050 $Y=228240
X512 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=22540 220320 0 0 $X=22350 $Y=220080
X513 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=23460 225760 0 0 $X=23270 $Y=225520
X514 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=28060 220320 0 0 $X=27870 $Y=220080
X515 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=48760 209440 0 0 $X=48570 $Y=209200
X516 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=49680 225760 0 0 $X=49490 $Y=225520
X517 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=55200 225760 0 0 $X=55010 $Y=225520
X518 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=57500 225760 1 0 $X=57310 $Y=222800
X519 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=62100 209440 0 0 $X=61910 $Y=209200
X520 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=69000 242080 0 0 $X=68810 $Y=241840
X521 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=118220 182240 0 0 $X=118030 $Y=182000
X522 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=182160 225760 1 0 $X=181970 $Y=222800
X523 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=202400 225760 0 0 $X=202210 $Y=225520
X524 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=213900 214880 0 0 $X=213710 $Y=214640
X525 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=223100 214880 0 0 $X=222910 $Y=214640
X526 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=242880 225760 0 0 $X=242690 $Y=225520
X527 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=243340 242080 0 0 $X=243150 $Y=241840
X528 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=322000 225760 0 0 $X=321810 $Y=225520
X529 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=332120 231200 0 0 $X=331930 $Y=230960
X530 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=336260 242080 0 0 $X=336070 $Y=241840
X531 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=492200 231200 0 0 $X=492010 $Y=230960
X532 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=500020 225760 0 0 $X=499830 $Y=225520
X533 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=504620 242080 0 0 $X=504430 $Y=241840
X534 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=511060 193120 0 0 $X=510870 $Y=192880
X535 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=514740 214880 0 0 $X=514550 $Y=214640
X536 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=517960 220320 1 0 $X=517770 $Y=217360
X537 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=600300 220320 1 0 $X=600110 $Y=217360
X538 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=623300 220320 0 0 $X=623110 $Y=220080
X539 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=665620 214880 1 0 $X=665430 $Y=211920
X540 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=671140 214880 1 0 $X=670950 $Y=211920
X541 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=671600 182240 1 0 $X=671410 $Y=179280
X542 1 2 613 601 2 45 1 sky130_fd_sc_hd__ebufn_2 $T=28980 198560 0 0 $X=28790 $Y=198320
X543 1 2 632 640 2 50 1 sky130_fd_sc_hd__ebufn_2 $T=41860 198560 1 0 $X=41670 $Y=195600
X544 1 2 629 619 2 41 1 sky130_fd_sc_hd__ebufn_2 $T=43240 242080 1 0 $X=43050 $Y=239120
X545 1 2 678 681 2 31 1 sky130_fd_sc_hd__ebufn_2 $T=63940 204000 0 0 $X=63750 $Y=203760
X546 1 2 680 681 2 27 1 sky130_fd_sc_hd__ebufn_2 $T=64400 198560 0 0 $X=64210 $Y=198320
X547 1 2 682 672 2 46 1 sky130_fd_sc_hd__ebufn_2 $T=65320 225760 1 0 $X=65130 $Y=222800
X548 1 2 701 691 2 45 1 sky130_fd_sc_hd__ebufn_2 $T=71760 225760 1 0 $X=71570 $Y=222800
X549 1 2 699 681 2 44 1 sky130_fd_sc_hd__ebufn_2 $T=76360 198560 1 0 $X=76170 $Y=195600
X550 1 2 709 710 2 31 1 sky130_fd_sc_hd__ebufn_2 $T=78200 193120 1 0 $X=78010 $Y=190160
X551 1 2 715 73 2 40 1 sky130_fd_sc_hd__ebufn_2 $T=81880 236640 0 0 $X=81690 $Y=236400
X552 1 2 721 76 2 45 1 sky130_fd_sc_hd__ebufn_2 $T=83720 187680 0 0 $X=83530 $Y=187440
X553 1 2 730 76 2 31 1 sky130_fd_sc_hd__ebufn_2 $T=88320 187680 1 0 $X=88130 $Y=184720
X554 1 2 94 87 2 40 1 sky130_fd_sc_hd__ebufn_2 $T=100280 242080 0 0 $X=100090 $Y=241840
X555 1 2 759 757 2 19 1 sky130_fd_sc_hd__ebufn_2 $T=101660 214880 0 0 $X=101470 $Y=214640
X556 1 2 812 110 2 48 1 sky130_fd_sc_hd__ebufn_2 $T=138000 182240 0 0 $X=137810 $Y=182000
X557 1 2 825 808 2 41 1 sky130_fd_sc_hd__ebufn_2 $T=139380 236640 0 0 $X=139190 $Y=236400
X558 1 2 837 110 2 31 1 sky130_fd_sc_hd__ebufn_2 $T=143980 193120 1 0 $X=143790 $Y=190160
X559 1 2 843 807 2 50 1 sky130_fd_sc_hd__ebufn_2 $T=149040 193120 0 0 $X=148850 $Y=192880
X560 1 2 874 881 2 19 1 sky130_fd_sc_hd__ebufn_2 $T=169740 204000 0 0 $X=169550 $Y=203760
X561 1 2 880 882 2 135 1 sky130_fd_sc_hd__ebufn_2 $T=169740 236640 0 0 $X=169550 $Y=236400
X562 1 2 879 129 2 48 1 sky130_fd_sc_hd__ebufn_2 $T=173880 193120 1 0 $X=173690 $Y=190160
X563 1 2 166 164 2 151 1 sky130_fd_sc_hd__ebufn_2 $T=196420 242080 0 0 $X=196230 $Y=241840
X564 1 2 920 177 2 44 1 sky130_fd_sc_hd__ebufn_2 $T=208840 182240 0 0 $X=208650 $Y=182000
X565 1 2 937 177 2 31 1 sky130_fd_sc_hd__ebufn_2 $T=209300 182240 1 0 $X=209110 $Y=179280
X566 1 2 952 170 2 152 1 sky130_fd_sc_hd__ebufn_2 $T=210680 242080 0 0 $X=210490 $Y=241840
X567 1 2 995 966 2 196 1 sky130_fd_sc_hd__ebufn_2 $T=225400 193120 0 0 $X=225210 $Y=192880
X568 1 2 999 974 2 156 1 sky130_fd_sc_hd__ebufn_2 $T=230460 225760 0 0 $X=230270 $Y=225520
X569 1 2 1007 985 2 211 1 sky130_fd_sc_hd__ebufn_2 $T=235980 225760 1 0 $X=235790 $Y=222800
X570 1 2 1012 193 2 219 1 sky130_fd_sc_hd__ebufn_2 $T=240120 187680 1 0 $X=239930 $Y=184720
X571 1 2 1013 983 2 219 1 sky130_fd_sc_hd__ebufn_2 $T=240120 193120 1 0 $X=239930 $Y=190160
X572 1 2 1034 1020 2 157 1 sky130_fd_sc_hd__ebufn_2 $T=248400 242080 1 0 $X=248210 $Y=239120
X573 1 2 1049 1046 2 198 1 sky130_fd_sc_hd__ebufn_2 $T=253920 214880 1 0 $X=253730 $Y=211920
X574 1 2 1061 224 2 198 1 sky130_fd_sc_hd__ebufn_2 $T=260360 193120 0 0 $X=260170 $Y=192880
X575 1 2 1074 1078 2 195 1 sky130_fd_sc_hd__ebufn_2 $T=272780 209440 1 0 $X=272590 $Y=206480
X576 1 2 1107 1100 2 155 1 sky130_fd_sc_hd__ebufn_2 $T=286580 225760 0 0 $X=286390 $Y=225520
X577 1 2 1101 1100 2 152 1 sky130_fd_sc_hd__ebufn_2 $T=294860 242080 1 0 $X=294670 $Y=239120
X578 1 2 1119 258 2 196 1 sky130_fd_sc_hd__ebufn_2 $T=299460 182240 0 0 $X=299270 $Y=182000
X579 1 2 1150 268 2 219 1 sky130_fd_sc_hd__ebufn_2 $T=314640 182240 1 0 $X=314450 $Y=179280
X580 1 2 1163 268 2 211 1 sky130_fd_sc_hd__ebufn_2 $T=316020 187680 0 0 $X=315830 $Y=187440
X581 1 2 1175 1155 2 185 1 sky130_fd_sc_hd__ebufn_2 $T=331660 187680 0 0 $X=331470 $Y=187440
X582 1 2 294 274 2 155 1 sky130_fd_sc_hd__ebufn_2 $T=332120 242080 0 0 $X=331930 $Y=241840
X583 1 2 1190 1184 2 194 1 sky130_fd_sc_hd__ebufn_2 $T=337640 220320 0 0 $X=337450 $Y=220080
X584 1 2 1263 1248 2 271 1 sky130_fd_sc_hd__ebufn_2 $T=376740 236640 1 0 $X=376550 $Y=233680
X585 1 2 1298 1280 2 261 1 sky130_fd_sc_hd__ebufn_2 $T=394680 209440 1 0 $X=394490 $Y=206480
X586 1 2 1302 351 2 211 1 sky130_fd_sc_hd__ebufn_2 $T=397440 193120 1 0 $X=397250 $Y=190160
X587 1 2 1326 1327 2 261 1 sky130_fd_sc_hd__ebufn_2 $T=408480 198560 1 0 $X=408290 $Y=195600
X588 1 2 1329 1327 2 252 1 sky130_fd_sc_hd__ebufn_2 $T=409860 193120 0 0 $X=409670 $Y=192880
X589 1 2 1324 351 2 216 1 sky130_fd_sc_hd__ebufn_2 $T=413080 193120 1 0 $X=412890 $Y=190160
X590 1 2 1290 1248 2 329 1 sky130_fd_sc_hd__ebufn_2 $T=414460 225760 0 0 $X=414270 $Y=225520
X591 1 2 1335 1297 2 232 1 sky130_fd_sc_hd__ebufn_2 $T=419980 231200 0 0 $X=419790 $Y=230960
X592 1 2 1344 1327 2 263 1 sky130_fd_sc_hd__ebufn_2 $T=421820 204000 0 0 $X=421630 $Y=203760
X593 1 2 1348 1351 2 263 1 sky130_fd_sc_hd__ebufn_2 $T=422280 182240 0 0 $X=422090 $Y=182000
X594 1 2 1361 1366 2 255 1 sky130_fd_sc_hd__ebufn_2 $T=428720 236640 0 0 $X=428530 $Y=236400
X595 1 2 1353 1351 2 254 1 sky130_fd_sc_hd__ebufn_2 $T=430100 187680 1 0 $X=429910 $Y=184720
X596 1 2 1380 1368 2 263 1 sky130_fd_sc_hd__ebufn_2 $T=434700 225760 0 0 $X=434510 $Y=225520
X597 1 2 1402 370 2 238 1 sky130_fd_sc_hd__ebufn_2 $T=448040 231200 0 0 $X=447850 $Y=230960
X598 1 2 1408 1347 2 231 1 sky130_fd_sc_hd__ebufn_2 $T=454940 198560 1 0 $X=454750 $Y=195600
X599 1 2 1450 1449 2 255 1 sky130_fd_sc_hd__ebufn_2 $T=470580 187680 1 0 $X=470390 $Y=184720
X600 1 2 1406 1347 2 194 1 sky130_fd_sc_hd__ebufn_2 $T=476100 198560 0 0 $X=475910 $Y=198320
X601 1 2 1459 392 2 232 1 sky130_fd_sc_hd__ebufn_2 $T=477020 182240 0 0 $X=476830 $Y=182000
X602 1 2 1464 393 2 329 1 sky130_fd_sc_hd__ebufn_2 $T=478400 236640 0 0 $X=478210 $Y=236400
X603 1 2 401 393 2 249 1 sky130_fd_sc_hd__ebufn_2 $T=494040 242080 0 0 $X=493850 $Y=241840
X604 1 2 1498 1477 2 285 1 sky130_fd_sc_hd__ebufn_2 $T=494500 225760 0 0 $X=494310 $Y=225520
X605 1 2 1521 1499 2 330 1 sky130_fd_sc_hd__ebufn_2 $T=506000 187680 0 0 $X=505810 $Y=187440
X606 1 2 410 411 2 415 1 sky130_fd_sc_hd__ebufn_2 $T=506460 182240 0 0 $X=506270 $Y=182000
X607 1 2 1524 1465 2 232 1 sky130_fd_sc_hd__ebufn_2 $T=509680 214880 1 0 $X=509490 $Y=211920
X608 1 2 1536 1534 2 330 1 sky130_fd_sc_hd__ebufn_2 $T=518420 187680 1 0 $X=518230 $Y=184720
X609 1 2 1544 426 2 414 1 sky130_fd_sc_hd__ebufn_2 $T=520720 182240 0 0 $X=520530 $Y=182000
X610 1 2 1556 1534 2 251 1 sky130_fd_sc_hd__ebufn_2 $T=527160 193120 1 0 $X=526970 $Y=190160
X611 1 2 1607 1580 2 415 1 sky130_fd_sc_hd__ebufn_2 $T=552460 225760 0 0 $X=552270 $Y=225520
X612 1 2 1621 1605 2 329 1 sky130_fd_sc_hd__ebufn_2 $T=561200 193120 1 0 $X=561010 $Y=190160
X613 1 2 458 460 2 285 1 sky130_fd_sc_hd__ebufn_2 $T=575460 236640 0 0 $X=575270 $Y=236400
X614 1 2 1669 1652 2 285 1 sky130_fd_sc_hd__ebufn_2 $T=596160 220320 1 0 $X=595970 $Y=217360
X615 1 2 1705 1704 2 255 1 sky130_fd_sc_hd__ebufn_2 $T=609500 204000 1 0 $X=609310 $Y=201040
X616 1 2 1712 1713 2 249 1 sky130_fd_sc_hd__ebufn_2 $T=610880 236640 1 0 $X=610690 $Y=233680
X617 1 2 1785 1739 2 255 1 sky130_fd_sc_hd__ebufn_2 $T=646300 236640 0 0 $X=646110 $Y=236400
X618 1 2 1791 1739 2 329 1 sky130_fd_sc_hd__ebufn_2 $T=651360 236640 0 0 $X=651170 $Y=236400
X619 1 2 1797 1759 2 330 1 sky130_fd_sc_hd__ebufn_2 $T=655960 214880 0 0 $X=655770 $Y=214640
X620 1 2 1798 1783 2 238 1 sky130_fd_sc_hd__ebufn_2 $T=656880 198560 1 0 $X=656690 $Y=195600
X621 1 2 1810 500 2 330 1 sky130_fd_sc_hd__ebufn_2 $T=660560 242080 1 0 $X=660370 $Y=239120
X622 1 2 1817 1812 2 414 1 sky130_fd_sc_hd__ebufn_2 $T=665620 242080 1 0 $X=665430 $Y=239120
X623 1 2 1823 501 2 414 1 sky130_fd_sc_hd__ebufn_2 $T=667460 182240 1 0 $X=667270 $Y=179280
X624 1 2 1834 1831 2 427 1 sky130_fd_sc_hd__ebufn_2 $T=670680 187680 0 0 $X=670490 $Y=187440
X625 1 2 1887 509 2 427 1 sky130_fd_sc_hd__ebufn_2 $T=695520 242080 1 0 $X=695330 $Y=239120
X626 1 2 1893 1856 2 430 1 sky130_fd_sc_hd__ebufn_2 $T=702420 231200 0 0 $X=702230 $Y=230960
X627 1 2 1919 510 2 415 1 sky130_fd_sc_hd__ebufn_2 $T=712080 225760 0 0 $X=711890 $Y=225520
X628 1 2 1930 1901 2 415 1 sky130_fd_sc_hd__ebufn_2 $T=717140 193120 1 0 $X=716950 $Y=190160
X629 1 2 1931 1932 2 427 1 sky130_fd_sc_hd__ebufn_2 $T=717140 220320 1 0 $X=716950 $Y=217360
X630 1 2 1956 1901 2 412 1 sky130_fd_sc_hd__ebufn_2 $T=730480 182240 0 0 $X=730290 $Y=182000
X631 1 2 1951 1954 2 412 1 sky130_fd_sc_hd__ebufn_2 $T=730940 204000 0 0 $X=730750 $Y=203760
X632 1 2 1952 1932 2 412 1 sky130_fd_sc_hd__ebufn_2 $T=730940 209440 0 0 $X=730750 $Y=209200
X765 1 2 595 601 19 ICV_6 $T=19780 198560 1 0 $X=19590 $Y=195600
X766 1 2 597 603 19 ICV_6 $T=19780 209440 1 0 $X=19590 $Y=206480
X767 1 2 596 603 27 ICV_6 $T=19780 214880 1 0 $X=19590 $Y=211920
X768 1 2 624 603 44 ICV_6 $T=33580 209440 0 0 $X=33390 $Y=209200
X769 1 2 610 3 46 ICV_6 $T=33580 236640 0 0 $X=33390 $Y=236400
X770 1 2 728 710 27 ICV_6 $T=89700 198560 0 0 $X=89510 $Y=198320
X771 1 2 772 757 44 ICV_6 $T=117760 209440 0 0 $X=117570 $Y=209200
X772 1 2 103 98 39 ICV_6 $T=117760 220320 0 0 $X=117570 $Y=220080
X773 1 2 817 780 44 ICV_6 $T=145820 204000 0 0 $X=145630 $Y=203760
X774 1 2 855 119 45 ICV_6 $T=160080 193120 1 0 $X=159890 $Y=190160
X775 1 2 864 834 31 ICV_6 $T=160080 214880 1 0 $X=159890 $Y=211920
X776 1 2 861 824 32 ICV_6 $T=160080 231200 1 0 $X=159890 $Y=228240
X777 1 2 863 824 41 ICV_6 $T=160080 242080 1 0 $X=159890 $Y=239120
X778 1 2 885 881 28 ICV_6 $T=173880 214880 0 0 $X=173690 $Y=214640
X779 1 2 917 882 157 ICV_6 $T=188140 242080 1 0 $X=187950 $Y=239120
X780 1 2 940 929 27 ICV_6 $T=201940 209440 0 0 $X=201750 $Y=209200
X781 1 2 186 187 155 ICV_6 $T=216200 242080 1 0 $X=216010 $Y=239120
X782 1 2 1030 224 185 ICV_6 $T=244260 187680 1 0 $X=244070 $Y=184720
X783 1 2 1051 234 216 ICV_6 $T=258060 182240 0 0 $X=257870 $Y=182000
X784 1 2 1085 1078 211 ICV_6 $T=272320 214880 1 0 $X=272130 $Y=211920
X785 1 2 1112 1091 195 ICV_6 $T=286120 204000 0 0 $X=285930 $Y=203760
X786 1 2 1135 1138 135 ICV_6 $T=300380 231200 1 0 $X=300190 $Y=228240
X787 1 2 1161 1155 212 ICV_6 $T=314180 193120 0 0 $X=313990 $Y=192880
X788 1 2 1160 1138 157 ICV_6 $T=314180 236640 0 0 $X=313990 $Y=236400
X789 1 2 1194 1184 254 ICV_6 $T=342240 214880 0 0 $X=342050 $Y=214640
X790 1 2 1214 1201 219 ICV_6 $T=356500 198560 1 0 $X=356310 $Y=195600
X791 1 2 1222 1201 198 ICV_6 $T=356500 204000 1 0 $X=356310 $Y=201040
X792 1 2 1227 1212 261 ICV_6 $T=356500 214880 1 0 $X=356310 $Y=211920
X793 1 2 1220 309 238 ICV_6 $T=356500 231200 1 0 $X=356310 $Y=228240
X794 1 2 1229 1193 185 ICV_6 $T=370300 187680 0 0 $X=370110 $Y=187440
X795 1 2 1274 1255 185 ICV_6 $T=384560 187680 1 0 $X=384370 $Y=184720
X796 1 2 1279 1268 211 ICV_6 $T=384560 204000 1 0 $X=384370 $Y=201040
X797 1 2 1325 351 212 ICV_6 $T=412620 187680 1 0 $X=412430 $Y=184720
X798 1 2 1319 1297 254 ICV_6 $T=412620 214880 1 0 $X=412430 $Y=211920
X799 1 2 358 355 285 ICV_6 $T=412620 242080 1 0 $X=412430 $Y=239120
X800 1 2 1362 364 244 ICV_6 $T=426420 182240 0 0 $X=426230 $Y=182000
X801 1 2 379 375 232 ICV_6 $T=454480 182240 0 0 $X=454290 $Y=182000
X802 1 2 1445 1423 238 ICV_6 $T=468740 225760 1 0 $X=468550 $Y=222800
X803 1 2 1469 1449 330 ICV_6 $T=482540 187680 0 0 $X=482350 $Y=187440
X804 1 2 1467 1449 249 ICV_6 $T=482540 193120 0 0 $X=482350 $Y=192880
X805 1 2 395 393 330 ICV_6 $T=482540 242080 0 0 $X=482350 $Y=241840
X806 1 2 1501 1477 255 ICV_6 $T=496800 225760 1 0 $X=496610 $Y=222800
X807 1 2 1500 393 285 ICV_6 $T=496800 242080 1 0 $X=496610 $Y=239120
X808 1 2 1529 420 413 ICV_6 $T=510600 236640 0 0 $X=510410 $Y=236400
X809 1 2 1548 420 427 ICV_6 $T=524860 242080 1 0 $X=524670 $Y=239120
X810 1 2 438 437 424 ICV_6 $T=538660 242080 0 0 $X=538470 $Y=241840
X811 1 2 1596 1581 285 ICV_6 $T=552920 193120 1 0 $X=552730 $Y=190160
X812 1 2 1611 1580 414 ICV_6 $T=552920 220320 1 0 $X=552730 $Y=217360
X813 1 2 1608 1612 415 ICV_6 $T=552920 236640 1 0 $X=552730 $Y=233680
X814 1 2 1610 1612 414 ICV_6 $T=552920 242080 1 0 $X=552730 $Y=239120
X815 1 2 1622 443 271 ICV_6 $T=566720 182240 0 0 $X=566530 $Y=182000
X816 1 2 1631 1636 255 ICV_6 $T=566720 220320 0 0 $X=566530 $Y=220080
X817 1 2 1633 1612 424 ICV_6 $T=566720 231200 0 0 $X=566530 $Y=230960
X818 1 2 1620 443 238 ICV_6 $T=580980 187680 1 0 $X=580790 $Y=184720
X819 1 2 1656 1649 238 ICV_6 $T=580980 209440 1 0 $X=580790 $Y=206480
X820 1 2 1677 1653 330 ICV_6 $T=594780 225760 0 0 $X=594590 $Y=225520
X821 1 2 1711 1713 285 ICV_6 $T=609040 242080 1 0 $X=608850 $Y=239120
X822 1 2 1729 1736 271 ICV_6 $T=622840 214880 0 0 $X=622650 $Y=214640
X823 1 2 1734 1713 330 ICV_6 $T=622840 236640 0 0 $X=622650 $Y=236400
X824 1 2 1847 1818 414 ICV_6 $T=678960 214880 0 0 $X=678770 $Y=214640
X825 1 2 1848 1818 412 ICV_6 $T=678960 220320 0 0 $X=678770 $Y=220080
X826 1 2 1840 1812 427 ICV_6 $T=678960 231200 0 0 $X=678770 $Y=230960
X827 1 2 1877 1865 427 ICV_6 $T=693220 204000 1 0 $X=693030 $Y=201040
X828 1 2 1875 1844 412 ICV_6 $T=693220 225760 1 0 $X=693030 $Y=222800
X829 1 2 1904 506 429 ICV_6 $T=707020 182240 0 0 $X=706830 $Y=182000
X830 1 2 1936 1938 415 ICV_6 $T=721280 231200 1 0 $X=721090 $Y=228240
X831 1 2 1946 1938 427 ICV_6 $T=735080 220320 0 0 $X=734890 $Y=220080
X970 1 2 9 11 2 592 1 sky130_fd_sc_hd__dfxtp_1 $T=12420 187680 0 0 $X=12230 $Y=187440
X971 1 2 589 33 2 624 1 sky130_fd_sc_hd__dfxtp_1 $T=25300 209440 0 0 $X=25110 $Y=209200
X972 1 2 608 6 2 638 1 sky130_fd_sc_hd__dfxtp_1 $T=37720 231200 0 0 $X=37530 $Y=230960
X973 1 2 608 21 2 651 1 sky130_fd_sc_hd__dfxtp_1 $T=39560 236640 0 0 $X=39370 $Y=236400
X974 1 2 49 11 2 654 1 sky130_fd_sc_hd__dfxtp_1 $T=45540 187680 0 0 $X=45350 $Y=187440
X975 1 2 660 33 2 699 1 sky130_fd_sc_hd__dfxtp_1 $T=64860 198560 1 0 $X=64670 $Y=195600
X976 1 2 660 36 2 705 1 sky130_fd_sc_hd__dfxtp_1 $T=68080 209440 1 0 $X=67890 $Y=206480
X977 1 2 702 14 2 79 1 sky130_fd_sc_hd__dfxtp_1 $T=73600 231200 0 0 $X=73410 $Y=230960
X978 1 2 702 7 2 713 1 sky130_fd_sc_hd__dfxtp_1 $T=74060 225760 0 0 $X=73870 $Y=225520
X979 1 2 702 21 2 715 1 sky130_fd_sc_hd__dfxtp_1 $T=74520 242080 0 0 $X=74330 $Y=241840
X980 1 2 89 11 2 749 1 sky130_fd_sc_hd__dfxtp_1 $T=92460 187680 0 0 $X=92270 $Y=187440
X981 1 2 86 24 2 733 1 sky130_fd_sc_hd__dfxtp_1 $T=98440 236640 0 0 $X=98250 $Y=236400
X982 1 2 751 10 2 755 1 sky130_fd_sc_hd__dfxtp_1 $T=106720 220320 0 0 $X=106530 $Y=220080
X983 1 2 97 24 2 782 1 sky130_fd_sc_hd__dfxtp_1 $T=108100 242080 1 0 $X=107910 $Y=239120
X984 1 2 793 7 2 830 1 sky130_fd_sc_hd__dfxtp_1 $T=133400 225760 0 0 $X=133210 $Y=225520
X985 1 2 104 10 2 837 1 sky130_fd_sc_hd__dfxtp_1 $T=136160 187680 1 0 $X=135970 $Y=184720
X986 1 2 813 36 2 841 1 sky130_fd_sc_hd__dfxtp_1 $T=141220 225760 1 0 $X=141030 $Y=222800
X987 1 2 116 12 2 851 1 sky130_fd_sc_hd__dfxtp_1 $T=146740 182240 1 0 $X=146550 $Y=179280
X988 1 2 813 10 2 864 1 sky130_fd_sc_hd__dfxtp_1 $T=153640 214880 0 0 $X=153450 $Y=214640
X989 1 2 127 46 2 884 1 sky130_fd_sc_hd__dfxtp_1 $T=165600 225760 0 0 $X=165410 $Y=225520
X990 1 2 875 132 2 891 1 sky130_fd_sc_hd__dfxtp_1 $T=169740 236640 1 0 $X=169550 $Y=233680
X991 1 2 875 148 2 916 1 sky130_fd_sc_hd__dfxtp_1 $T=181700 231200 0 0 $X=181510 $Y=230960
X992 1 2 911 10 2 935 1 sky130_fd_sc_hd__dfxtp_1 $T=193200 204000 0 0 $X=193010 $Y=203760
X993 1 2 905 13 2 950 1 sky130_fd_sc_hd__dfxtp_1 $T=199180 198560 1 0 $X=198990 $Y=195600
X994 1 2 905 10 2 951 1 sky130_fd_sc_hd__dfxtp_1 $T=203780 204000 1 0 $X=203590 $Y=201040
X995 1 2 127 28 2 961 1 sky130_fd_sc_hd__dfxtp_1 $T=206540 220320 0 0 $X=206350 $Y=220080
X996 1 2 127 32 2 969 1 sky130_fd_sc_hd__dfxtp_1 $T=207920 225760 1 0 $X=207730 $Y=222800
X997 1 2 127 8 2 971 1 sky130_fd_sc_hd__dfxtp_1 $T=211600 225760 0 0 $X=211410 $Y=225520
X998 1 2 955 138 2 972 1 sky130_fd_sc_hd__dfxtp_1 $T=211600 236640 0 0 $X=211410 $Y=236400
X999 1 2 180 183 2 978 1 sky130_fd_sc_hd__dfxtp_1 $T=214360 182240 0 0 $X=214170 $Y=182000
X1000 1 2 955 132 2 998 1 sky130_fd_sc_hd__dfxtp_1 $T=221720 231200 0 0 $X=221530 $Y=230960
X1001 1 2 228 183 2 1050 1 sky130_fd_sc_hd__dfxtp_1 $T=248400 182240 1 0 $X=248210 $Y=179280
X1002 1 2 127 230 2 1054 1 sky130_fd_sc_hd__dfxtp_1 $T=250240 220320 0 0 $X=250050 $Y=220080
X1003 1 2 1048 146 2 1057 1 sky130_fd_sc_hd__dfxtp_1 $T=260360 231200 1 0 $X=260170 $Y=228240
X1004 1 2 228 200 2 1082 1 sky130_fd_sc_hd__dfxtp_1 $T=264500 182240 1 0 $X=264310 $Y=179280
X1005 1 2 1062 199 2 1085 1 sky130_fd_sc_hd__dfxtp_1 $T=266340 220320 0 0 $X=266150 $Y=220080
X1006 1 2 1092 147 2 1101 1 sky130_fd_sc_hd__dfxtp_1 $T=275080 236640 0 0 $X=274890 $Y=236400
X1007 1 2 1096 199 2 1110 1 sky130_fd_sc_hd__dfxtp_1 $T=278300 220320 0 0 $X=278110 $Y=220080
X1008 1 2 127 249 2 1019 1 sky130_fd_sc_hd__dfxtp_1 $T=285200 214880 1 0 $X=285010 $Y=211920
X1009 1 2 1108 183 2 1119 1 sky130_fd_sc_hd__dfxtp_1 $T=285660 182240 1 0 $X=285470 $Y=179280
X1010 1 2 1108 182 2 1120 1 sky130_fd_sc_hd__dfxtp_1 $T=286120 187680 1 0 $X=285930 $Y=184720
X1011 1 2 1116 138 2 1139 1 sky130_fd_sc_hd__dfxtp_1 $T=295320 236640 0 0 $X=295130 $Y=236400
X1012 1 2 1156 181 2 1165 1 sky130_fd_sc_hd__dfxtp_1 $T=312340 209440 1 0 $X=312150 $Y=206480
X1013 1 2 1197 181 2 1224 1 sky130_fd_sc_hd__dfxtp_1 $T=348220 193120 1 0 $X=348030 $Y=190160
X1014 1 2 1202 300 2 314 1 sky130_fd_sc_hd__dfxtp_1 $T=348680 242080 1 0 $X=348490 $Y=239120
X1015 1 2 1183 183 2 1226 1 sky130_fd_sc_hd__dfxtp_1 $T=350060 198560 0 0 $X=349870 $Y=198320
X1016 1 2 1203 278 2 1227 1 sky130_fd_sc_hd__dfxtp_1 $T=350060 209440 0 0 $X=349870 $Y=209200
X1017 1 2 1197 182 2 1229 1 sky130_fd_sc_hd__dfxtp_1 $T=350980 182240 0 0 $X=350790 $Y=182000
X1018 1 2 1234 284 2 1244 1 sky130_fd_sc_hd__dfxtp_1 $T=359720 209440 1 0 $X=359530 $Y=206480
X1019 1 2 127 155 2 328 1 sky130_fd_sc_hd__dfxtp_1 $T=361100 231200 1 0 $X=360910 $Y=228240
X1020 1 2 1237 205 2 1254 1 sky130_fd_sc_hd__dfxtp_1 $T=365240 187680 1 0 $X=365050 $Y=184720
X1021 1 2 1234 282 2 1257 1 sky130_fd_sc_hd__dfxtp_1 $T=367080 220320 1 0 $X=366890 $Y=217360
X1022 1 2 1252 201 2 1272 1 sky130_fd_sc_hd__dfxtp_1 $T=373060 198560 0 0 $X=372870 $Y=198320
X1023 1 2 1237 201 2 1275 1 sky130_fd_sc_hd__dfxtp_1 $T=377200 187680 1 0 $X=377010 $Y=184720
X1024 1 2 1252 199 2 1279 1 sky130_fd_sc_hd__dfxtp_1 $T=378120 204000 0 0 $X=377930 $Y=203760
X1025 1 2 1262 280 2 1281 1 sky130_fd_sc_hd__dfxtp_1 $T=378120 214880 0 0 $X=377930 $Y=214640
X1026 1 2 1262 267 2 1300 1 sky130_fd_sc_hd__dfxtp_1 $T=388700 220320 1 0 $X=388510 $Y=217360
X1027 1 2 1339 284 2 1353 1 sky130_fd_sc_hd__dfxtp_1 $T=418140 187680 0 0 $X=417950 $Y=187440
X1028 1 2 1339 278 2 1355 1 sky130_fd_sc_hd__dfxtp_1 $T=420440 198560 1 0 $X=420250 $Y=195600
X1029 1 2 1342 280 2 1367 1 sky130_fd_sc_hd__dfxtp_1 $T=421360 220320 1 0 $X=421170 $Y=217360
X1030 1 2 1339 279 2 1348 1 sky130_fd_sc_hd__dfxtp_1 $T=425500 193120 1 0 $X=425310 $Y=190160
X1031 1 2 1342 275 2 1385 1 sky130_fd_sc_hd__dfxtp_1 $T=429640 214880 1 0 $X=429450 $Y=211920
X1032 1 2 1412 299 2 1439 1 sky130_fd_sc_hd__dfxtp_1 $T=456780 242080 1 0 $X=456590 $Y=239120
X1033 1 2 1428 317 2 1421 1 sky130_fd_sc_hd__dfxtp_1 $T=467820 225760 0 0 $X=467630 $Y=225520
X1034 1 2 1428 298 2 1441 1 sky130_fd_sc_hd__dfxtp_1 $T=468740 220320 0 0 $X=468550 $Y=220080
X1035 1 2 1440 299 2 1466 1 sky130_fd_sc_hd__dfxtp_1 $T=473800 198560 1 0 $X=473610 $Y=195600
X1036 1 2 389 318 2 1464 1 sky130_fd_sc_hd__dfxtp_1 $T=475180 242080 0 0 $X=474990 $Y=241840
X1037 1 2 1476 280 2 1524 1 sky130_fd_sc_hd__dfxtp_1 $T=504620 209440 1 0 $X=504430 $Y=206480
X1038 1 2 1526 298 2 1537 1 sky130_fd_sc_hd__dfxtp_1 $T=511060 193120 1 0 $X=510870 $Y=190160
X1039 1 2 1594 406 2 1608 1 sky130_fd_sc_hd__dfxtp_1 $T=545560 242080 1 0 $X=545370 $Y=239120
X1040 1 2 1617 286 2 1630 1 sky130_fd_sc_hd__dfxtp_1 $T=557980 214880 0 0 $X=557790 $Y=214640
X1041 1 2 1617 288 2 1631 1 sky130_fd_sc_hd__dfxtp_1 $T=557980 220320 0 0 $X=557790 $Y=220080
X1042 1 2 1598 318 2 454 1 sky130_fd_sc_hd__dfxtp_1 $T=560740 187680 1 0 $X=560550 $Y=184720
X1043 1 2 1637 298 2 1647 1 sky130_fd_sc_hd__dfxtp_1 $T=572240 198560 1 0 $X=572050 $Y=195600
X1044 1 2 1637 299 2 1656 1 sky130_fd_sc_hd__dfxtp_1 $T=573620 209440 1 0 $X=573430 $Y=206480
X1045 1 2 1642 318 2 1651 1 sky130_fd_sc_hd__dfxtp_1 $T=574080 225760 0 0 $X=573890 $Y=225520
X1046 1 2 1643 317 2 1650 1 sky130_fd_sc_hd__dfxtp_1 $T=575000 209440 0 0 $X=574810 $Y=209200
X1047 1 2 1643 286 2 1675 1 sky130_fd_sc_hd__dfxtp_1 $T=584660 209440 0 0 $X=584470 $Y=209200
X1048 1 2 1685 298 2 1707 1 sky130_fd_sc_hd__dfxtp_1 $T=599380 225760 0 0 $X=599190 $Y=225520
X1049 1 2 1688 318 2 1709 1 sky130_fd_sc_hd__dfxtp_1 $T=602600 231200 0 0 $X=602410 $Y=230960
X1050 1 2 473 318 2 1679 1 sky130_fd_sc_hd__dfxtp_1 $T=603520 182240 0 0 $X=603330 $Y=182000
X1051 1 2 1714 318 2 1756 1 sky130_fd_sc_hd__dfxtp_1 $T=625600 209440 1 0 $X=625410 $Y=206480
X1052 1 2 1795 423 2 1811 1 sky130_fd_sc_hd__dfxtp_1 $T=655500 236640 1 0 $X=655310 $Y=233680
X1053 1 2 1795 406 2 1833 1 sky130_fd_sc_hd__dfxtp_1 $T=663780 236640 0 0 $X=663590 $Y=236400
X1054 1 2 1816 406 2 1842 1 sky130_fd_sc_hd__dfxtp_1 $T=670680 193120 0 0 $X=670490 $Y=192880
X1055 1 2 1802 404 2 1847 1 sky130_fd_sc_hd__dfxtp_1 $T=671600 214880 0 0 $X=671410 $Y=214640
X1056 1 2 1802 403 2 1848 1 sky130_fd_sc_hd__dfxtp_1 $T=671600 220320 0 0 $X=671410 $Y=220080
X1057 1 2 1815 421 2 1850 1 sky130_fd_sc_hd__dfxtp_1 $T=672980 209440 1 0 $X=672790 $Y=206480
X1058 1 2 1815 403 2 1853 1 sky130_fd_sc_hd__dfxtp_1 $T=681260 204000 1 0 $X=681070 $Y=201040
X1059 1 2 1816 409 2 1858 1 sky130_fd_sc_hd__dfxtp_1 $T=682180 187680 1 0 $X=681990 $Y=184720
X1060 1 2 1839 422 2 1873 1 sky130_fd_sc_hd__dfxtp_1 $T=683560 231200 0 0 $X=683370 $Y=230960
X1061 1 2 1866 422 2 1877 1 sky130_fd_sc_hd__dfxtp_1 $T=685860 198560 0 0 $X=685670 $Y=198320
X1062 1 2 1867 404 2 1883 1 sky130_fd_sc_hd__dfxtp_1 $T=687240 209440 0 0 $X=687050 $Y=209200
X1063 1 2 505 423 2 1904 1 sky130_fd_sc_hd__dfxtp_1 $T=698740 182240 0 0 $X=698550 $Y=182000
X1064 1 2 1866 406 2 1916 1 sky130_fd_sc_hd__dfxtp_1 $T=707480 204000 1 0 $X=707290 $Y=201040
X1065 1 2 1876 422 2 1924 1 sky130_fd_sc_hd__dfxtp_1 $T=710240 187680 1 0 $X=710050 $Y=184720
X1066 1 2 1917 403 2 1937 1 sky130_fd_sc_hd__dfxtp_1 $T=713000 231200 1 0 $X=712810 $Y=228240
X1067 1 2 1935 421 2 1948 1 sky130_fd_sc_hd__dfxtp_1 $T=718980 214880 0 0 $X=718790 $Y=214640
X1068 1 2 1917 423 2 1963 1 sky130_fd_sc_hd__dfxtp_1 $T=727720 220320 0 0 $X=727530 $Y=220080
X1069 1 2 1923 405 2 1898 1 sky130_fd_sc_hd__dfxtp_1 $T=730020 242080 1 0 $X=729830 $Y=239120
X1070 1 2 611 3 41 587 25 611 ICV_13 $T=20240 242080 1 0 $X=20050 $Y=239120
X1071 1 2 620 601 44 588 35 621 ICV_13 $T=24380 198560 1 0 $X=24190 $Y=195600
X1072 1 2 53 55 46 608 25 629 ICV_13 $T=31740 242080 1 0 $X=31550 $Y=239120
X1073 1 2 635 640 44 626 35 632 ICV_13 $T=34500 204000 1 0 $X=34310 $Y=201040
X1074 1 2 633 641 28 627 34 637 ICV_13 $T=34960 220320 1 0 $X=34770 $Y=217360
X1075 1 2 639 640 31 626 10 639 ICV_13 $T=35420 209440 1 0 $X=35230 $Y=206480
X1076 1 2 662 641 27 627 13 662 ICV_13 $T=48300 214880 1 0 $X=48110 $Y=211920
X1077 1 2 663 641 31 627 10 663 ICV_13 $T=48300 220320 1 0 $X=48110 $Y=217360
X1078 1 2 665 640 27 626 11 661 ICV_13 $T=49220 198560 0 0 $X=49030 $Y=198320
X1079 1 2 666 672 32 653 6 666 ICV_13 $T=50140 231200 0 0 $X=49950 $Y=230960
X1080 1 2 677 681 45 660 34 677 ICV_13 $T=56580 204000 1 0 $X=56390 $Y=201040
X1081 1 2 671 672 18 653 24 682 ICV_13 $T=58880 231200 1 0 $X=58690 $Y=228240
X1082 1 2 688 672 8 653 5 688 ICV_13 $T=62100 231200 0 0 $X=61910 $Y=230960
X1083 1 2 692 694 28 676 12 692 ICV_13 $T=62560 220320 1 0 $X=62370 $Y=217360
X1084 1 2 716 73 46 676 34 712 ICV_13 $T=74060 220320 0 0 $X=73870 $Y=220080
X1085 1 2 706 681 19 703 10 709 ICV_13 $T=76360 198560 0 0 $X=76170 $Y=198320
X1086 1 2 718 694 19 676 11 718 ICV_13 $T=76360 220320 1 0 $X=76170 $Y=217360
X1087 1 2 719 73 32 702 6 719 ICV_13 $T=76360 236640 1 0 $X=76170 $Y=233680
X1088 1 2 720 73 41 702 25 720 ICV_13 $T=76360 242080 1 0 $X=76170 $Y=239120
X1089 1 2 731 710 44 703 33 731 ICV_13 $T=82340 193120 1 0 $X=82150 $Y=190160
X1090 1 2 746 750 48 735 36 746 ICV_13 $T=92000 204000 1 0 $X=91810 $Y=201040
X1091 1 2 748 93 31 89 10 748 ICV_13 $T=92460 187680 1 0 $X=92270 $Y=184720
X1092 1 2 739 691 27 734 11 687 ICV_13 $T=97520 209440 0 0 $X=97330 $Y=209200
X1093 1 2 761 750 44 735 33 761 ICV_13 $T=97980 198560 0 0 $X=97790 $Y=198320
X1094 1 2 765 773 18 760 7 765 ICV_13 $T=104420 225760 0 0 $X=104230 $Y=225520
X1095 1 2 767 773 41 760 25 767 ICV_13 $T=104420 236640 1 0 $X=104230 $Y=233680
X1096 1 2 771 757 48 751 33 772 ICV_13 $T=105800 214880 0 0 $X=105610 $Y=214640
X1097 1 2 774 773 66 760 14 774 ICV_13 $T=105800 236640 0 0 $X=105610 $Y=236400
X1098 1 2 790 792 50 784 35 790 ICV_13 $T=115920 193120 1 0 $X=115730 $Y=190160
X1099 1 2 794 792 48 784 36 794 ICV_13 $T=118220 187680 0 0 $X=118030 $Y=187440
X1100 1 2 795 773 32 760 6 795 ICV_13 $T=118220 225760 0 0 $X=118030 $Y=225520
X1101 1 2 801 757 28 751 12 801 ICV_13 $T=120060 214880 1 0 $X=119870 $Y=211920
X1102 1 2 823 792 19 784 11 823 ICV_13 $T=132480 193120 1 0 $X=132290 $Y=190160
X1103 1 2 826 792 44 784 33 826 ICV_13 $T=133400 187680 0 0 $X=133210 $Y=187440
X1104 1 2 829 834 28 813 12 829 ICV_13 $T=133400 220320 0 0 $X=133210 $Y=220080
X1105 1 2 835 110 44 104 33 835 ICV_13 $T=135240 182240 1 0 $X=135050 $Y=179280
X1106 1 2 842 807 27 819 33 849 ICV_13 $T=146280 198560 0 0 $X=146090 $Y=198320
X1107 1 2 862 824 66 836 5 865 ICV_13 $T=153640 236640 0 0 $X=153450 $Y=236400
X1108 1 2 877 881 50 866 35 877 ICV_13 $T=162380 209440 0 0 $X=162190 $Y=209200
X1109 1 2 887 868 27 860 13 887 ICV_13 $T=167900 198560 1 0 $X=167710 $Y=195600
X1110 1 2 889 881 31 860 33 893 ICV_13 $T=172040 204000 1 0 $X=171850 $Y=201040
X1111 1 2 899 129 31 125 10 899 ICV_13 $T=174340 187680 0 0 $X=174150 $Y=187440
X1112 1 2 888 882 151 136 138 145 ICV_13 $T=174340 242080 0 0 $X=174150 $Y=241840
X1113 1 2 902 882 153 875 149 917 ICV_13 $T=181700 236640 0 0 $X=181510 $Y=236400
X1114 1 2 928 929 45 911 34 928 ICV_13 $T=188600 214880 1 0 $X=188410 $Y=211920
X1115 1 2 958 929 19 911 36 956 ICV_13 $T=202400 214880 0 0 $X=202210 $Y=214640
X1116 1 2 956 929 48 911 11 958 ICV_13 $T=203780 214880 1 0 $X=203590 $Y=211920
X1117 1 2 979 983 185 962 181 976 ICV_13 $T=213900 193120 0 0 $X=213710 $Y=192880
X1118 1 2 986 193 195 180 188 986 ICV_13 $T=216660 182240 1 0 $X=216470 $Y=179280
X1119 1 2 987 983 195 962 188 987 ICV_13 $T=216660 187680 1 0 $X=216470 $Y=184720
X1120 1 2 976 983 198 962 182 979 ICV_13 $T=216660 193120 1 0 $X=216470 $Y=190160
X1121 1 2 989 966 198 963 181 989 ICV_13 $T=216660 198560 1 0 $X=216470 $Y=195600
X1122 1 2 990 966 195 963 188 990 ICV_13 $T=216660 204000 1 0 $X=216470 $Y=201040
X1123 1 2 991 985 195 967 188 991 ICV_13 $T=216660 209440 1 0 $X=216470 $Y=206480
X1124 1 2 992 985 198 967 181 992 ICV_13 $T=216660 214880 1 0 $X=216470 $Y=211920
X1125 1 2 972 974 153 955 137 975 ICV_13 $T=216660 236640 1 0 $X=216470 $Y=233680
X1126 1 2 993 985 196 967 183 993 ICV_13 $T=217580 204000 0 0 $X=217390 $Y=203760
X1127 1 2 997 974 151 955 149 996 ICV_13 $T=220800 242080 1 0 $X=220610 $Y=239120
X1128 1 2 1014 983 216 962 205 1014 ICV_13 $T=230460 193120 0 0 $X=230270 $Y=192880
X1129 1 2 1017 966 212 963 201 1016 ICV_13 $T=230460 198560 0 0 $X=230270 $Y=198320
X1130 1 2 1006 985 219 963 200 1017 ICV_13 $T=230460 204000 0 0 $X=230270 $Y=203760
X1131 1 2 1018 985 212 967 200 1018 ICV_13 $T=230460 209440 0 0 $X=230270 $Y=209200
X1132 1 2 1039 224 211 1028 201 1047 ICV_13 $T=246100 187680 0 0 $X=245910 $Y=187440
X1133 1 2 1044 1046 216 1022 181 1049 ICV_13 $T=246560 214880 0 0 $X=246370 $Y=214640
X1134 1 2 1052 234 211 228 199 1052 ICV_13 $T=248860 187680 1 0 $X=248670 $Y=184720
X1135 1 2 246 247 153 240 147 1094 ICV_13 $T=270020 242080 0 0 $X=269830 $Y=241840
X1136 1 2 1104 1091 198 127 244 982 ICV_13 $T=274620 214880 0 0 $X=274430 $Y=214640
X1137 1 2 1095 1087 195 1066 201 1097 ICV_13 $T=276460 193120 1 0 $X=276270 $Y=190160
X1138 1 2 1106 1087 212 1066 200 1106 ICV_13 $T=276460 198560 1 0 $X=276270 $Y=195600
X1139 1 2 1109 1091 216 1096 205 1109 ICV_13 $T=278300 220320 1 0 $X=278110 $Y=217360
X1140 1 2 1110 1091 211 127 251 1008 ICV_13 $T=286580 214880 0 0 $X=286390 $Y=214640
X1141 1 2 1124 1100 142 1092 132 1124 ICV_13 $T=287040 231200 1 0 $X=286850 $Y=228240
X1142 1 2 1129 258 212 1108 200 1129 ICV_13 $T=288880 198560 0 0 $X=288690 $Y=198320
X1143 1 2 1147 1136 211 1121 182 1146 ICV_13 $T=300840 209440 1 0 $X=300650 $Y=206480
X1144 1 2 1149 1138 151 1116 130 1149 ICV_13 $T=302680 236640 0 0 $X=302490 $Y=236400
X1145 1 2 1151 268 212 262 201 1150 ICV_13 $T=303140 182240 1 0 $X=302950 $Y=179280
X1146 1 2 1158 1155 195 1141 188 1158 ICV_13 $T=305900 193120 1 0 $X=305710 $Y=190160
X1147 1 2 1174 1155 216 1141 182 1175 ICV_13 $T=320160 187680 0 0 $X=319970 $Y=187440
X1148 1 2 1177 274 156 264 148 1177 ICV_13 $T=320620 242080 0 0 $X=320430 $Y=241840
X1149 1 2 1169 1172 219 1156 183 1170 ICV_13 $T=322000 198560 0 0 $X=321810 $Y=198320
X1150 1 2 1185 1155 198 1141 181 1185 ICV_13 $T=327060 193120 0 0 $X=326870 $Y=192880
X1151 1 2 1186 292 211 283 199 1186 ICV_13 $T=328900 187680 1 0 $X=328710 $Y=184720
X1152 1 2 1187 1155 211 1141 199 1187 ICV_13 $T=328900 193120 1 0 $X=328710 $Y=190160
X1153 1 2 1195 1201 216 1183 199 1198 ICV_13 $T=333960 209440 1 0 $X=333770 $Y=206480
X1154 1 2 1204 1184 231 1173 296 1204 ICV_13 $T=336260 225760 1 0 $X=336070 $Y=222800
X1155 1 2 303 292 185 283 183 1205 ICV_13 $T=336720 182240 1 0 $X=336530 $Y=179280
X1156 1 2 1210 309 251 1202 297 1216 ICV_13 $T=342700 236640 0 0 $X=342510 $Y=236400
X1157 1 2 1219 1212 231 1203 296 1219 ICV_13 $T=344540 220320 1 0 $X=344350 $Y=217360
X1158 1 2 1223 1201 212 1183 200 1223 ICV_13 $T=346380 204000 0 0 $X=346190 $Y=203760
X1159 1 2 1216 309 249 1202 318 1241 ICV_13 $T=356960 242080 1 0 $X=356770 $Y=239120
X1160 1 2 1253 1255 212 1237 200 1253 ICV_13 $T=364780 193120 1 0 $X=364590 $Y=190160
X1161 1 2 1265 1248 251 1249 286 1265 ICV_13 $T=370760 225760 0 0 $X=370570 $Y=225520
X1162 1 2 1266 336 249 331 297 1266 ICV_13 $T=370760 236640 0 0 $X=370570 $Y=236400
X1163 1 2 1269 1268 195 1252 188 1269 ICV_13 $T=372140 198560 1 0 $X=371950 $Y=195600
X1164 1 2 1275 1255 219 1237 182 1274 ICV_13 $T=377200 182240 0 0 $X=377010 $Y=182000
X1165 1 2 1284 336 251 331 286 1284 ICV_13 $T=381800 242080 0 0 $X=381610 $Y=241840
X1166 1 2 1289 1268 185 1252 182 1289 ICV_13 $T=385020 198560 1 0 $X=384830 $Y=195600
X1167 1 2 1291 1248 249 1249 297 1291 ICV_13 $T=385020 236640 1 0 $X=384830 $Y=233680
X1168 1 2 1292 336 285 331 298 1292 ICV_13 $T=385020 242080 1 0 $X=384830 $Y=239120
X1169 1 2 1293 1268 216 1252 205 1293 ICV_13 $T=385480 204000 0 0 $X=385290 $Y=203760
X1170 1 2 1299 1280 254 1262 278 1298 ICV_13 $T=388700 214880 1 0 $X=388510 $Y=211920
X1171 1 2 1315 1311 330 1301 317 1315 ICV_13 $T=398820 236640 0 0 $X=398630 $Y=236400
X1172 1 2 1318 1327 232 1308 267 1321 ICV_13 $T=401120 209440 1 0 $X=400930 $Y=206480
X1173 1 2 1343 1327 244 1308 282 1343 ICV_13 $T=412620 198560 0 0 $X=412430 $Y=198320
X1174 1 2 1345 1311 249 1301 297 1345 ICV_13 $T=413080 236640 1 0 $X=412890 $Y=233680
X1175 1 2 1358 1368 244 1342 267 1363 ICV_13 $T=419980 225760 1 0 $X=419790 $Y=222800
X1176 1 2 1373 364 231 360 296 1373 ICV_13 $T=426880 182240 1 0 $X=426690 $Y=179280
X1177 1 2 1359 1366 285 361 317 1371 ICV_13 $T=426880 231200 0 0 $X=426690 $Y=230960
X1178 1 2 1374 1351 252 1339 282 1378 ICV_13 $T=427800 198560 1 0 $X=427610 $Y=195600
X1179 1 2 1381 1368 231 1342 296 1381 ICV_13 $T=428720 220320 1 0 $X=428530 $Y=217360
X1180 1 2 1388 1389 254 1369 280 1390 ICV_13 $T=431940 204000 0 0 $X=431750 $Y=203760
X1181 1 2 1400 370 255 1375 288 1400 ICV_13 $T=441140 231200 1 0 $X=440950 $Y=228240
X1182 1 2 1401 370 251 1375 286 1401 ICV_13 $T=441140 236640 0 0 $X=440950 $Y=236400
X1183 1 2 1393 364 252 360 279 1386 ICV_13 $T=441600 182240 0 0 $X=441410 $Y=182000
X1184 1 2 374 375 194 1395 279 1346 ICV_13 $T=442980 187680 0 0 $X=442790 $Y=187440
X1185 1 2 1397 1337 254 1391 278 1417 ICV_13 $T=448040 214880 1 0 $X=447850 $Y=211920
X1186 1 2 1433 1438 249 1415 297 1433 ICV_13 $T=455400 204000 1 0 $X=455210 $Y=201040
X1187 1 2 1446 1422 330 1412 317 1446 ICV_13 $T=462300 231200 0 0 $X=462110 $Y=230960
X1188 1 2 1471 1449 251 1440 286 1471 ICV_13 $T=474720 187680 1 0 $X=474530 $Y=184720
X1189 1 2 1487 1477 330 1456 317 1487 ICV_13 $T=483000 225760 0 0 $X=482810 $Y=225520
X1190 1 2 1488 1491 271 1474 300 1488 ICV_13 $T=483460 204000 1 0 $X=483270 $Y=201040
X1191 1 2 1489 1465 261 1476 278 1489 ICV_13 $T=483460 214880 1 0 $X=483270 $Y=211920
X1192 1 2 1494 1499 249 1481 298 1495 ICV_13 $T=487140 193120 0 0 $X=486950 $Y=192880
X1193 1 2 1505 1499 251 1481 286 1505 ICV_13 $T=492660 182240 0 0 $X=492470 $Y=182000
X1194 1 2 1509 1491 249 1474 297 1509 ICV_13 $T=497260 204000 0 0 $X=497070 $Y=203760
X1195 1 2 1514 1520 413 1504 405 1514 ICV_13 $T=497720 236640 0 0 $X=497530 $Y=236400
X1196 1 2 1517 1491 330 1474 317 1517 ICV_13 $T=498640 198560 0 0 $X=498450 $Y=198320
X1197 1 2 1537 1534 285 1526 317 1536 ICV_13 $T=511060 187680 0 0 $X=510870 $Y=187440
X1198 1 2 1538 1534 271 1526 300 1538 ICV_13 $T=511060 198560 1 0 $X=510870 $Y=195600
X1199 1 2 1541 1520 424 1504 409 1541 ICV_13 $T=511060 231200 0 0 $X=510870 $Y=230960
X1200 1 2 1540 1520 429 408 405 1529 ICV_13 $T=511520 242080 1 0 $X=511330 $Y=239120
X1201 1 2 1547 420 429 408 422 1548 ICV_13 $T=516120 242080 0 0 $X=515930 $Y=241840
X1202 1 2 1565 426 415 416 406 1565 ICV_13 $T=524860 182240 0 0 $X=524670 $Y=182000
X1203 1 2 1566 1534 249 1526 297 1566 ICV_13 $T=525320 198560 1 0 $X=525130 $Y=195600
X1204 1 2 1555 1530 429 1508 421 1558 ICV_13 $T=525320 220320 1 0 $X=525130 $Y=217360
X1205 1 2 1567 1568 424 1551 409 1567 ICV_13 $T=525320 236640 1 0 $X=525130 $Y=233680
X1206 1 2 1574 1546 413 1535 405 1574 ICV_13 $T=529000 204000 1 0 $X=528810 $Y=201040
X1207 1 2 1575 1546 412 1535 403 1575 ICV_13 $T=529000 209440 1 0 $X=528810 $Y=206480
X1208 1 2 1586 1581 330 1563 317 1586 ICV_13 $T=535440 187680 1 0 $X=535250 $Y=184720
X1209 1 2 1591 1580 424 1576 409 1591 ICV_13 $T=537280 214880 1 0 $X=537090 $Y=211920
X1210 1 2 1577 1581 255 1563 300 1593 ICV_13 $T=540040 193120 1 0 $X=539850 $Y=190160
X1211 1 2 1609 1580 413 1576 405 1609 ICV_13 $T=546480 220320 0 0 $X=546290 $Y=220080
X1212 1 2 1619 437 413 436 405 1619 ICV_13 $T=552000 242080 0 0 $X=551810 $Y=241840
X1213 1 2 1650 1652 330 1617 318 1638 ICV_13 $T=569480 214880 1 0 $X=569290 $Y=211920
X1214 1 2 1655 1653 238 1642 298 1661 ICV_13 $T=580980 231200 0 0 $X=580790 $Y=230960
X1215 1 2 1668 1667 271 463 300 1668 ICV_13 $T=581900 193120 0 0 $X=581710 $Y=192880
X1216 1 2 1657 1652 238 1643 298 1669 ICV_13 $T=581900 220320 0 0 $X=581710 $Y=220080
X1217 1 2 1680 1653 271 1642 300 1680 ICV_13 $T=586040 236640 1 0 $X=585850 $Y=233680
X1218 1 2 1693 1699 255 1685 288 1693 ICV_13 $T=596620 225760 1 0 $X=596430 $Y=222800
X1219 1 2 1718 1699 329 1685 318 1718 ICV_13 $T=609500 231200 1 0 $X=609310 $Y=228240
X1220 1 2 1720 1699 271 1685 300 1720 ICV_13 $T=610420 225760 0 0 $X=610230 $Y=225520
X1221 1 2 1733 1713 255 1688 317 1734 ICV_13 $T=615020 236640 1 0 $X=614830 $Y=233680
X1222 1 2 1740 1745 249 1727 297 1740 ICV_13 $T=620080 225760 1 0 $X=619890 $Y=222800
X1223 1 2 1742 1745 251 1727 286 1742 ICV_13 $T=620540 220320 1 0 $X=620350 $Y=217360
X1224 1 2 1751 493 271 488 299 1752 ICV_13 $T=625140 198560 1 0 $X=624950 $Y=195600
X1225 1 2 1761 1739 238 1743 298 1762 ICV_13 $T=628360 231200 0 0 $X=628170 $Y=230960
X1226 1 2 1769 1745 271 1727 288 1772 ICV_13 $T=637560 225760 1 0 $X=637370 $Y=222800
X1227 1 2 1773 500 249 495 297 1773 ICV_13 $T=637560 242080 1 0 $X=637370 $Y=239120
X1228 1 2 1782 1783 271 1768 300 1782 ICV_13 $T=639400 198560 0 0 $X=639210 $Y=198320
X1229 1 2 1786 1787 329 1770 297 1784 ICV_13 $T=639860 187680 1 0 $X=639670 $Y=184720
X1230 1 2 1796 500 251 495 286 1796 ICV_13 $T=649060 242080 1 0 $X=648870 $Y=239120
X1231 1 2 1803 1787 251 1770 286 1803 ICV_13 $T=651360 187680 1 0 $X=651170 $Y=184720
X1232 1 2 1804 1787 330 1770 317 1804 ICV_13 $T=651360 187680 0 0 $X=651170 $Y=187440
X1233 1 2 1805 1787 285 1770 298 1805 ICV_13 $T=651360 193120 0 0 $X=651170 $Y=192880
X1234 1 2 1806 1783 285 1768 298 1806 ICV_13 $T=651360 204000 0 0 $X=651170 $Y=203760
X1235 1 2 1807 1759 251 1765 286 1807 ICV_13 $T=651360 209440 0 0 $X=651170 $Y=209200
X1236 1 2 502 500 238 495 317 1810 ICV_13 $T=651360 242080 0 0 $X=651170 $Y=241840
X1237 1 2 1821 1818 424 1802 409 1821 ICV_13 $T=660100 214880 0 0 $X=659910 $Y=214640
X1238 1 2 1832 1826 414 1815 406 1827 ICV_13 $T=662860 209440 0 0 $X=662670 $Y=209200
X1239 1 2 1836 1831 429 1816 423 1836 ICV_13 $T=665620 198560 1 0 $X=665430 $Y=195600
X1240 1 2 1838 1812 424 1795 409 1838 ICV_13 $T=666540 231200 0 0 $X=666350 $Y=230960
X1241 1 2 1843 1812 430 1795 421 1843 ICV_13 $T=669760 242080 1 0 $X=669570 $Y=239120
X1242 1 2 1845 1818 430 1802 421 1845 ICV_13 $T=671140 220320 1 0 $X=670950 $Y=217360
X1243 1 2 1868 1831 412 1816 403 1868 ICV_13 $T=679420 193120 0 0 $X=679230 $Y=192880
X1244 1 2 1850 1826 430 1815 405 1852 ICV_13 $T=680340 209440 1 0 $X=680150 $Y=206480
X1245 1 2 1878 1865 413 1866 405 1878 ICV_13 $T=685860 204000 0 0 $X=685670 $Y=203760
X1246 1 2 1889 1856 414 1839 404 1889 ICV_13 $T=690920 231200 0 0 $X=690730 $Y=230960
X1247 1 2 1894 1886 427 1867 422 1894 ICV_13 $T=694600 209440 0 0 $X=694410 $Y=209200
X1248 1 2 1902 1844 430 1861 421 1902 ICV_13 $T=697820 225760 1 0 $X=697630 $Y=222800
X1249 1 2 1906 1844 424 1861 409 1906 ICV_13 $T=699200 231200 1 0 $X=699010 $Y=228240
X1250 1 2 1925 1886 424 1867 409 1925 ICV_13 $T=707480 209440 0 0 $X=707290 $Y=209200
X1251 1 2 1926 1886 430 1867 421 1926 ICV_13 $T=707480 214880 0 0 $X=707290 $Y=214640
X1252 1 2 1928 509 429 508 423 1928 ICV_13 $T=709320 242080 1 0 $X=709130 $Y=239120
X1253 1 2 1940 519 430 514 421 1940 ICV_13 $T=714840 242080 0 0 $X=714650 $Y=241840
X1254 1 2 1937 1938 412 1917 421 1943 ICV_13 $T=716220 225760 0 0 $X=716030 $Y=225520
X1255 1 2 1949 1901 430 1933 406 1930 ICV_13 $T=718520 193120 0 0 $X=718330 $Y=192880
X1256 1 2 1944 510 430 1923 406 1919 ICV_13 $T=723580 236640 0 0 $X=723390 $Y=236400
X1257 1 2 1966 1938 413 1917 405 1966 ICV_13 $T=730020 225760 1 0 $X=729830 $Y=222800
X1258 1 2 1970 1901 414 513 405 1967 ICV_13 $T=730480 187680 1 0 $X=730290 $Y=184720
X1259 1 2 1971 1954 414 1934 404 1971 ICV_13 $T=731400 198560 1 0 $X=731210 $Y=195600
X1260 1 2 627 33 656 656 641 44 ICV_14 $T=45080 214880 0 0 $X=44890 $Y=214640
X1261 1 2 652 33 664 664 659 44 ICV_14 $T=48300 182240 0 0 $X=48110 $Y=182000
X1262 1 2 660 10 678 674 681 50 ICV_14 $T=55660 209440 1 0 $X=55470 $Y=206480
X1263 1 2 653 21 696 696 672 40 ICV_14 $T=62100 236640 1 0 $X=61910 $Y=233680
X1264 1 2 74 12 707 707 76 28 ICV_14 $T=69460 182240 0 0 $X=69270 $Y=182000
X1265 1 2 676 13 722 723 694 44 ICV_14 $T=76360 214880 1 0 $X=76170 $Y=211920
X1266 1 2 735 11 737 737 750 19 ICV_14 $T=90160 193120 0 0 $X=89970 $Y=192880
X1267 1 2 734 35 744 743 750 45 ICV_14 $T=90620 209440 1 0 $X=90430 $Y=206480
X1268 1 2 764 10 788 788 780 31 ICV_14 $T=112240 204000 1 0 $X=112050 $Y=201040
X1269 1 2 784 13 797 797 792 27 ICV_14 $T=118220 193120 0 0 $X=118030 $Y=192880
X1270 1 2 104 13 800 800 110 27 ICV_14 $T=118680 182240 1 0 $X=118490 $Y=179280
X1271 1 2 793 5 806 815 808 66 ICV_14 $T=126960 236640 0 0 $X=126770 $Y=236400
X1272 1 2 764 33 817 818 780 48 ICV_14 $T=129720 204000 0 0 $X=129530 $Y=203760
X1273 1 2 784 34 827 827 792 45 ICV_14 $T=132480 198560 1 0 $X=132290 $Y=195600
X1274 1 2 813 11 828 828 834 19 ICV_14 $T=132480 220320 1 0 $X=132290 $Y=217360
X1275 1 2 897 12 924 900 868 19 ICV_14 $T=185840 187680 0 0 $X=185650 $Y=187440
X1276 1 2 967 182 980 980 985 185 ICV_14 $T=213900 209440 0 0 $X=213710 $Y=209200
X1277 1 2 189 130 994 994 187 151 ICV_14 $T=217120 242080 0 0 $X=216930 $Y=241840
X1278 1 2 963 199 1015 1015 966 211 ICV_14 $T=229540 198560 1 0 $X=229350 $Y=195600
X1279 1 2 1002 149 1034 1036 1020 151 ICV_14 $T=241040 236640 0 0 $X=240850 $Y=236400
X1280 1 2 1048 132 1079 1079 1055 142 ICV_14 $T=263120 231200 0 0 $X=262930 $Y=230960
X1281 1 2 1121 205 1144 1144 1136 216 ICV_14 $T=298080 214880 0 0 $X=297890 $Y=214640
X1282 1 2 127 152 332 1240 309 330 ICV_14 $T=364320 236640 1 0 $X=364130 $Y=233680
X1283 1 2 1234 279 1258 1243 1239 252 ICV_14 $T=367080 209440 1 0 $X=366890 $Y=206480
X1284 1 2 361 300 1376 1376 1366 271 ICV_14 $T=425960 242080 1 0 $X=425770 $Y=239120
X1285 1 2 1339 267 1377 1378 1351 244 ICV_14 $T=426880 193120 0 0 $X=426690 $Y=192880
X1286 1 2 1375 317 1403 1396 370 285 ICV_14 $T=441140 225760 0 0 $X=440950 $Y=225520
X1287 1 2 373 267 1434 383 382 252 ICV_14 $T=454940 182240 1 0 $X=454750 $Y=179280
X1288 1 2 1415 317 1435 1435 1438 330 ICV_14 $T=454940 209440 0 0 $X=454750 $Y=209200
X1289 1 2 1440 298 1451 1451 1449 285 ICV_14 $T=463680 198560 0 0 $X=463490 $Y=198320
X1290 1 2 1476 282 1515 1515 1465 244 ICV_14 $T=497260 214880 1 0 $X=497070 $Y=211920
X1291 1 2 1582 299 1599 1578 1581 238 ICV_14 $T=540500 204000 1 0 $X=540310 $Y=201040
X1292 1 2 1582 297 1601 1601 1605 249 ICV_14 $T=540500 209440 1 0 $X=540310 $Y=206480
X1293 1 2 1594 421 1613 1613 1612 430 ICV_14 $T=546480 231200 0 0 $X=546290 $Y=230960
X1294 1 2 1582 286 1625 1625 1605 251 ICV_14 $T=555680 204000 1 0 $X=555490 $Y=201040
X1295 1 2 1643 318 1662 1660 1652 249 ICV_14 $T=575460 214880 0 0 $X=575270 $Y=214640
X1296 1 2 1637 318 1682 1683 1649 330 ICV_14 $T=585580 209440 1 0 $X=585390 $Y=206480
X1297 1 2 1685 317 1696 1696 1699 330 ICV_14 $T=596160 231200 1 0 $X=595970 $Y=228240
X1298 1 2 1768 318 1776 1776 1783 329 ICV_14 $T=637560 209440 1 0 $X=637370 $Y=206480
X1299 1 2 1768 317 1801 1801 1783 330 ICV_14 $T=649980 209440 1 0 $X=649790 $Y=206480
X1300 1 2 1765 299 1808 1808 1759 238 ICV_14 $T=650440 214880 1 0 $X=650250 $Y=211920
X1301 1 2 1795 405 1813 1813 1812 413 ICV_14 $T=654120 231200 0 0 $X=653930 $Y=230960
X1302 1 2 1876 421 1891 1891 1885 430 ICV_14 $T=690920 193120 0 0 $X=690730 $Y=192880
X1303 1 2 1935 405 1973 1974 1932 414 ICV_14 $T=730480 214880 1 0 $X=730290 $Y=211920
X1304 1 2 9 10 16 593 15 28 ICV_16 $T=10580 182240 0 0 $X=10390 $Y=182000
X1305 1 2 588 13 594 594 601 27 ICV_16 $T=10580 193120 0 0 $X=10390 $Y=192880
X1306 1 2 9 36 617 617 15 48 ICV_16 $T=23000 182240 1 0 $X=22810 $Y=179280
X1307 1 2 627 12 633 634 641 48 ICV_16 $T=34040 220320 0 0 $X=33850 $Y=220080
X1308 1 2 627 11 657 637 641 45 ICV_16 $T=46000 220320 0 0 $X=45810 $Y=220080
X1309 1 2 652 12 670 670 659 28 ICV_16 $T=50600 193120 1 0 $X=50410 $Y=190160
X1310 1 2 652 13 690 690 659 27 ICV_16 $T=62100 187680 0 0 $X=61910 $Y=187440
X1311 1 2 676 36 693 693 694 48 ICV_16 $T=62100 220320 0 0 $X=61910 $Y=220080
X1312 1 2 74 34 721 80 76 48 ICV_16 $T=76360 187680 1 0 $X=76170 $Y=184720
X1313 1 2 89 36 747 747 93 48 ICV_16 $T=92000 182240 1 0 $X=91810 $Y=179280
X1314 1 2 89 13 768 768 93 27 ICV_16 $T=104420 187680 1 0 $X=104230 $Y=184720
X1315 1 2 751 34 799 109 98 66 ICV_16 $T=119140 220320 1 0 $X=118950 $Y=217360
X1316 1 2 159 132 946 936 170 135 ICV_16 $T=196880 236640 1 0 $X=196690 $Y=233680
X1317 1 2 962 183 988 988 983 196 ICV_16 $T=216200 187680 0 0 $X=216010 $Y=187440
X1318 1 2 962 199 1004 1004 983 211 ICV_16 $T=228160 187680 1 0 $X=227970 $Y=184720
X1319 1 2 962 200 1005 1005 983 212 ICV_16 $T=228160 193120 1 0 $X=227970 $Y=190160
X1320 1 2 1002 147 1025 1026 1020 153 ICV_16 $T=232300 242080 1 0 $X=232110 $Y=239120
X1321 1 2 1022 183 1042 1041 1046 195 ICV_16 $T=244260 204000 0 0 $X=244070 $Y=203760
X1322 1 2 1092 130 1115 1115 1100 151 ICV_16 $T=281060 236640 1 0 $X=280870 $Y=233680
X1323 1 2 1108 201 1127 1126 258 198 ICV_16 $T=287960 193120 1 0 $X=287770 $Y=190160
X1324 1 2 1203 279 1228 1235 1212 244 ICV_16 $T=352820 220320 0 0 $X=352630 $Y=220080
X1325 1 2 1202 288 1236 1236 309 255 ICV_16 $T=354200 236640 0 0 $X=354010 $Y=236400
X1326 1 2 127 142 324 1226 1201 196 ICV_16 $T=357420 198560 0 0 $X=357230 $Y=198320
X1327 1 2 319 199 325 326 311 216 ICV_16 $T=358800 182240 1 0 $X=358610 $Y=179280
X1328 1 2 1301 298 1340 1340 1311 285 ICV_16 $T=410320 236640 0 0 $X=410130 $Y=236400
X1329 1 2 361 318 1370 1371 1366 330 ICV_16 $T=424580 236640 1 0 $X=424390 $Y=233680
X1330 1 2 1415 318 1455 1457 1438 271 ICV_16 $T=467360 209440 0 0 $X=467170 $Y=209200
X1331 1 2 388 280 1459 391 392 252 ICV_16 $T=469200 182240 1 0 $X=469010 $Y=179280
X1332 1 2 1456 318 1490 1490 1477 329 ICV_16 $T=483000 220320 0 0 $X=482810 $Y=220080
X1333 1 2 1504 403 1512 1512 1520 412 ICV_16 $T=497260 231200 1 0 $X=497070 $Y=228240
X1334 1 2 1504 404 1513 1513 1520 414 ICV_16 $T=497260 236640 1 0 $X=497070 $Y=233680
X1335 1 2 1504 406 1516 1516 1520 415 ICV_16 $T=497720 231200 0 0 $X=497530 $Y=230960
X1336 1 2 1481 299 1519 1519 1499 238 ICV_16 $T=498640 193120 0 0 $X=498450 $Y=192880
X1337 1 2 1508 423 1555 1558 1530 430 ICV_16 $T=519800 220320 0 0 $X=519610 $Y=220080
X1338 1 2 1526 288 1560 1560 1534 255 ICV_16 $T=522560 187680 0 0 $X=522370 $Y=187440
X1339 1 2 1551 421 1561 1561 1568 430 ICV_16 $T=523480 236640 0 0 $X=523290 $Y=236400
X1340 1 2 1551 422 1584 1584 1568 427 ICV_16 $T=534520 231200 1 0 $X=534330 $Y=228240
X1341 1 2 1563 297 1590 1557 1534 329 ICV_16 $T=536820 198560 1 0 $X=536630 $Y=195600
X1342 1 2 1637 288 1645 1646 1649 249 ICV_16 $T=568100 204000 1 0 $X=567910 $Y=201040
X1343 1 2 467 300 479 1689 477 251 ICV_16 $T=597080 242080 1 0 $X=596890 $Y=239120
X1344 1 2 1685 299 1716 1717 1699 251 ICV_16 $T=608580 220320 0 0 $X=608390 $Y=220080
X1345 1 2 1714 286 1753 1753 1736 251 ICV_16 $T=624680 204000 1 0 $X=624490 $Y=201040
X1346 1 2 1768 288 1774 1774 1783 255 ICV_16 $T=637560 204000 1 0 $X=637370 $Y=201040
X1347 1 2 1770 300 1781 1781 1787 271 ICV_16 $T=638940 193120 0 0 $X=638750 $Y=192880
X1348 1 2 1768 299 1798 1800 1783 251 ICV_16 $T=649520 204000 1 0 $X=649330 $Y=201040
X1349 1 2 1795 403 1837 1837 1812 412 ICV_16 $T=665620 242080 0 0 $X=665430 $Y=241840
X1350 1 2 1867 403 1914 1914 1886 412 ICV_16 $T=703340 214880 1 0 $X=703150 $Y=211920
X1351 1 2 1935 403 1952 1948 1932 430 ICV_16 $T=718980 209440 0 0 $X=718790 $Y=209200
X1352 1 2 1923 404 1968 525 517 429 ICV_16 $T=730020 236640 1 0 $X=729830 $Y=233680
X1353 1 2 589 10 598 598 603 31 ICV_17 $T=10580 214880 0 0 $X=10390 $Y=214640
X1354 1 2 784 10 798 798 792 31 ICV_17 $T=117760 198560 1 0 $X=117570 $Y=195600
X1355 1 2 875 130 888 891 882 142 ICV_17 $T=166980 242080 1 0 $X=166790 $Y=239120
X1356 1 2 127 27 930 923 929 50 ICV_17 $T=188600 220320 1 0 $X=188410 $Y=217360
X1357 1 2 897 11 953 954 177 27 ICV_17 $T=199180 193120 1 0 $X=198990 $Y=190160
X1358 1 2 180 199 1009 1009 193 211 ICV_17 $T=228160 182240 1 0 $X=227970 $Y=179280
X1359 1 2 1002 146 1033 1035 1020 156 ICV_17 $T=240120 231200 0 0 $X=239930 $Y=230960
X1360 1 2 1028 205 1058 1058 224 216 ICV_17 $T=252080 198560 1 0 $X=251890 $Y=195600
X1361 1 2 1108 188 1125 1125 258 195 ICV_17 $T=286580 182240 0 0 $X=286390 $Y=182000
X1362 1 2 1116 132 1145 1145 1138 142 ICV_17 $T=298540 225760 0 0 $X=298350 $Y=225520
X1363 1 2 1237 199 1273 1273 1255 211 ICV_17 $T=374900 187680 0 0 $X=374710 $Y=187440
X1364 1 2 1249 298 1287 1283 1248 238 ICV_17 $T=382260 225760 0 0 $X=382070 $Y=225520
X1365 1 2 1301 300 1312 1312 1311 271 ICV_17 $T=396520 236640 1 0 $X=396330 $Y=233680
X1366 1 2 1306 296 1313 1300 1280 194 ICV_17 $T=397440 220320 1 0 $X=397250 $Y=217360
X1367 1 2 360 267 1354 1354 364 194 ICV_17 $T=417220 187680 1 0 $X=417030 $Y=184720
X1368 1 2 1342 279 1380 1363 1368 194 ICV_17 $T=426880 220320 0 0 $X=426690 $Y=220080
X1369 1 2 1369 296 1404 1404 1389 231 ICV_17 $T=441140 209440 0 0 $X=440950 $Y=209200
X1370 1 2 1415 298 1437 1437 1438 285 ICV_17 $T=454940 209440 1 0 $X=454750 $Y=206480
X1371 1 2 1428 288 1460 1462 1465 263 ICV_17 $T=469660 214880 0 0 $X=469470 $Y=214640
X1372 1 2 1474 286 1483 1483 1491 251 ICV_17 $T=481160 198560 1 0 $X=480970 $Y=195600
X1373 1 2 1476 284 1492 1492 1465 254 ICV_17 $T=483000 209440 0 0 $X=482810 $Y=209200
X1374 1 2 1476 275 1511 1511 1465 252 ICV_17 $T=495880 209440 0 0 $X=495690 $Y=209200
X1375 1 2 1474 318 1518 1510 1491 255 ICV_17 $T=497260 204000 1 0 $X=497070 $Y=201040
X1376 1 2 1617 299 1640 1640 1636 238 ICV_17 $T=560740 231200 1 0 $X=560550 $Y=228240
X1377 1 2 463 286 1670 1670 1667 251 ICV_17 $T=581440 182240 1 0 $X=581250 $Y=179280
X1378 1 2 463 298 1671 1671 1667 285 ICV_17 $T=581440 198560 0 0 $X=581250 $Y=198320
X1379 1 2 473 317 478 480 471 251 ICV_17 $T=595700 182240 1 0 $X=595510 $Y=179280
X1380 1 2 481 286 1721 1721 486 251 ICV_17 $T=609500 182240 1 0 $X=609310 $Y=179280
X1381 1 2 481 298 1722 1697 471 285 ICV_17 $T=609500 193120 1 0 $X=609310 $Y=190160
X1382 1 2 488 288 1748 1748 493 255 ICV_17 $T=623300 182240 0 0 $X=623110 $Y=182000
X1383 1 2 488 318 1749 1750 493 285 ICV_17 $T=623300 187680 1 0 $X=623110 $Y=184720
X1384 1 2 1765 297 1777 1777 1759 249 ICV_17 $T=637560 209440 0 0 $X=637370 $Y=209200
X1385 1 2 1765 300 1778 1778 1759 271 ICV_17 $T=637560 214880 1 0 $X=637370 $Y=211920
X1386 1 2 1802 406 1822 1820 1818 429 ICV_17 $T=658720 220320 0 0 $X=658530 $Y=220080
X1387 1 2 1815 423 1824 1827 1826 415 ICV_17 $T=662860 204000 0 0 $X=662670 $Y=203760
X1388 1 2 508 406 1911 1911 509 415 ICV_17 $T=701040 236640 1 0 $X=700850 $Y=233680
X1389 1 2 1876 406 1918 1920 1885 412 ICV_17 $T=704720 198560 1 0 $X=704530 $Y=195600
X1390 1 2 1934 403 1951 1955 1932 415 ICV_17 $T=718060 204000 0 0 $X=717870 $Y=203760
X1391 1 2 676 10 685 685 694 31 ICV_19 $T=59800 214880 1 0 $X=59610 $Y=211920
X1392 1 2 676 35 697 697 694 50 ICV_19 $T=62100 214880 0 0 $X=61910 $Y=214640
X1393 1 2 652 10 698 698 659 31 ICV_19 $T=62560 193120 1 0 $X=62370 $Y=190160
X1394 1 2 676 33 723 722 694 27 ICV_19 $T=75440 214880 0 0 $X=75250 $Y=214640
X1395 1 2 703 12 724 705 681 48 ICV_19 $T=75900 204000 0 0 $X=75710 $Y=203760
X1396 1 2 735 35 770 776 750 27 ICV_19 $T=104420 198560 1 0 $X=104230 $Y=195600
X1397 1 2 813 35 831 831 834 50 ICV_19 $T=132020 214880 0 0 $X=131830 $Y=214640
X1398 1 2 167 13 947 947 158 27 ICV_19 $T=195960 182240 1 0 $X=195770 $Y=179280
X1399 1 2 333 181 1271 1271 337 198 ICV_19 $T=370760 182240 1 0 $X=370570 $Y=179280
X1400 1 2 1456 286 1472 1472 1477 251 ICV_19 $T=473340 225760 1 0 $X=473150 $Y=222800
X1401 1 2 388 267 1484 396 392 261 ICV_19 $T=481160 182240 1 0 $X=480970 $Y=179280
X1402 1 2 1504 423 1540 1539 1520 427 ICV_19 $T=509220 231200 1 0 $X=509030 $Y=228240
X1403 1 2 473 299 1694 1694 471 238 ICV_19 $T=595240 193120 0 0 $X=595050 $Y=192880
X1404 1 2 1685 297 1695 1695 1699 249 ICV_19 $T=595240 220320 0 0 $X=595050 $Y=220080
X1405 1 2 1727 317 1741 1744 1736 238 ICV_19 $T=618700 214880 1 0 $X=618510 $Y=211920
X1406 1 2 488 300 1751 1722 486 285 ICV_19 $T=623300 193120 0 0 $X=623110 $Y=192880
X1407 1 2 1714 298 1754 1754 1736 285 ICV_19 $T=623300 204000 0 0 $X=623110 $Y=203760
X1408 1 2 1768 297 1775 1775 1783 249 ICV_19 $T=636640 204000 0 0 $X=636450 $Y=203760
X1409 1 2 1770 288 1780 1784 1787 249 ICV_19 $T=637560 193120 1 0 $X=637370 $Y=190160
X1410 1 2 1935 409 1969 1963 1938 429 ICV_19 $T=729100 220320 1 0 $X=728910 $Y=217360
X1411 1 2 9 12 593 ICV_20 $T=10580 182240 1 0 $X=10390 $Y=179280
X1412 1 2 588 11 595 ICV_20 $T=10580 198560 1 0 $X=10390 $Y=195600
X1413 1 2 588 12 604 ICV_20 $T=12420 204000 0 0 $X=12230 $Y=203760
X1414 1 2 9 34 38 ICV_20 $T=22540 182240 0 0 $X=22350 $Y=182000
X1415 1 2 56 6 60 ICV_20 $T=40480 242080 0 0 $X=40290 $Y=241840
X1416 1 2 660 35 674 ICV_20 $T=53820 204000 0 0 $X=53630 $Y=203760
X1417 1 2 660 12 700 ICV_20 $T=68080 204000 0 0 $X=67890 $Y=203760
X1418 1 2 660 11 706 ICV_20 $T=68540 198560 0 0 $X=68350 $Y=198320
X1419 1 2 703 34 714 ICV_20 $T=76360 204000 1 0 $X=76170 $Y=201040
X1420 1 2 74 10 730 ICV_20 $T=81880 182240 0 0 $X=81690 $Y=182000
X1421 1 2 735 12 769 ICV_20 $T=104420 204000 1 0 $X=104230 $Y=201040
X1422 1 2 793 25 825 ICV_20 $T=132480 236640 1 0 $X=132290 $Y=233680
X1423 1 2 819 10 839 ICV_20 $T=138000 209440 0 0 $X=137810 $Y=209200
X1424 1 2 819 34 840 ICV_20 $T=146280 209440 0 0 $X=146090 $Y=209200
X1425 1 2 836 6 861 ICV_20 $T=152260 236640 1 0 $X=152070 $Y=233680
X1426 1 2 860 36 873 ICV_20 $T=160540 204000 1 0 $X=160350 $Y=201040
X1427 1 2 860 10 867 ICV_20 $T=160540 204000 0 0 $X=160350 $Y=203760
X1428 1 2 866 33 910 ICV_20 $T=178020 209440 1 0 $X=177830 $Y=206480
X1429 1 2 911 13 940 ICV_20 $T=194580 209440 1 0 $X=194390 $Y=206480
X1430 1 2 905 12 942 ICV_20 $T=195960 204000 1 0 $X=195770 $Y=201040
X1431 1 2 127 31 968 ICV_20 $T=207460 220320 1 0 $X=207270 $Y=217360
X1432 1 2 967 201 1006 ICV_20 $T=228160 209440 1 0 $X=227970 $Y=206480
X1433 1 2 967 199 1007 ICV_20 $T=228160 214880 1 0 $X=227970 $Y=211920
X1434 1 2 1022 201 1045 ICV_20 $T=244720 214880 1 0 $X=244530 $Y=211920
X1435 1 2 228 205 1051 ICV_20 $T=248400 182240 0 0 $X=248210 $Y=182000
X1436 1 2 127 237 1067 ICV_20 $T=258520 220320 0 0 $X=258330 $Y=220080
X1437 1 2 1062 205 1077 ICV_20 $T=262200 220320 1 0 $X=262010 $Y=217360
X1438 1 2 1048 137 1073 ICV_20 $T=263580 225760 0 0 $X=263390 $Y=225520
X1439 1 2 1092 137 1099 ICV_20 $T=275080 225760 0 0 $X=274890 $Y=225520
X1440 1 2 1066 181 1103 ICV_20 $T=276000 198560 0 0 $X=275810 $Y=198320
X1441 1 2 127 255 1118 ICV_20 $T=290720 225760 0 0 $X=290530 $Y=225520
X1442 1 2 1121 201 1134 ICV_20 $T=292560 214880 1 0 $X=292370 $Y=211920
X1443 1 2 1121 188 1143 ICV_20 $T=297160 204000 0 0 $X=296970 $Y=203760
X1444 1 2 262 205 1154 ICV_20 $T=303600 182240 0 0 $X=303410 $Y=182000
X1445 1 2 1141 201 1153 ICV_20 $T=303600 193120 0 0 $X=303410 $Y=192880
X1446 1 2 1116 146 1159 ICV_20 $T=306360 231200 0 0 $X=306170 $Y=230960
X1447 1 2 1141 200 1161 ICV_20 $T=306820 198560 1 0 $X=306630 $Y=195600
X1448 1 2 1116 147 1162 ICV_20 $T=308200 236640 1 0 $X=308010 $Y=233680
X1449 1 2 1156 201 1169 ICV_20 $T=314640 198560 1 0 $X=314450 $Y=195600
X1450 1 2 1141 205 1174 ICV_20 $T=317400 193120 1 0 $X=317210 $Y=190160
X1451 1 2 1173 278 1196 ICV_20 $T=333040 214880 0 0 $X=332850 $Y=214640
X1452 1 2 1197 183 1209 ICV_20 $T=340400 193120 1 0 $X=340210 $Y=190160
X1453 1 2 1202 286 1210 ICV_20 $T=340860 242080 1 0 $X=340670 $Y=239120
X1454 1 2 1203 275 1211 ICV_20 $T=341780 214880 1 0 $X=341590 $Y=211920
X1455 1 2 1203 267 1217 ICV_20 $T=342700 220320 0 0 $X=342510 $Y=220080
X1456 1 2 1234 280 1238 ICV_20 $T=359720 214880 0 0 $X=359530 $Y=214640
X1457 1 2 127 151 348 ICV_20 $T=389620 231200 0 0 $X=389430 $Y=230960
X1458 1 2 127 343 350 ICV_20 $T=390540 198560 0 0 $X=390350 $Y=198320
X1459 1 2 1306 284 1319 ICV_20 $T=400200 214880 1 0 $X=400010 $Y=211920
X1460 1 2 339 200 1325 ICV_20 $T=401580 193120 1 0 $X=401390 $Y=190160
X1461 1 2 1308 275 1329 ICV_20 $T=402500 204000 1 0 $X=402310 $Y=201040
X1462 1 2 1306 279 1295 ICV_20 $T=404800 225760 1 0 $X=404610 $Y=222800
X1463 1 2 361 298 1359 ICV_20 $T=418600 225760 0 0 $X=418410 $Y=225520
X1464 1 2 360 282 1362 ICV_20 $T=419060 182240 1 0 $X=418870 $Y=179280
X1465 1 2 1369 284 1388 ICV_20 $T=430100 209440 1 0 $X=429910 $Y=206480
X1466 1 2 1375 298 1396 ICV_20 $T=438380 231200 0 0 $X=438190 $Y=230960
X1467 1 2 1391 275 1416 ICV_20 $T=446660 214880 0 0 $X=446470 $Y=214640
X1468 1 2 1412 286 1425 ICV_20 $T=452640 231200 1 0 $X=452450 $Y=228240
X1469 1 2 1395 275 1429 ICV_20 $T=454020 187680 1 0 $X=453830 $Y=184720
X1470 1 2 1440 300 1447 ICV_20 $T=463680 193120 0 0 $X=463490 $Y=192880
X1471 1 2 389 298 1500 ICV_20 $T=488060 242080 1 0 $X=487870 $Y=239120
X1472 1 2 1508 405 1525 ICV_20 $T=502780 214880 0 0 $X=502590 $Y=214640
X1473 1 2 408 404 1527 ICV_20 $T=503700 242080 1 0 $X=503510 $Y=239120
X1474 1 2 1551 406 1564 ICV_20 $T=523940 231200 0 0 $X=523750 $Y=230960
X1475 1 2 1576 404 1611 ICV_20 $T=546480 214880 0 0 $X=546290 $Y=214640
X1476 1 2 1598 286 1614 ICV_20 $T=549700 182240 0 0 $X=549510 $Y=182000
X1477 1 2 1582 298 1623 ICV_20 $T=555680 209440 0 0 $X=555490 $Y=209200
X1478 1 2 1617 300 1627 ICV_20 $T=556600 225760 0 0 $X=556410 $Y=225520
X1479 1 2 1594 403 1628 ICV_20 $T=556600 236640 0 0 $X=556410 $Y=236400
X1480 1 2 1594 423 1632 ICV_20 $T=558900 231200 0 0 $X=558710 $Y=230960
X1481 1 2 1617 297 1639 ICV_20 $T=561660 214880 1 0 $X=561470 $Y=211920
X1482 1 2 447 406 455 ICV_20 $T=563040 182240 1 0 $X=562850 $Y=179280
X1483 1 2 1642 288 1681 ICV_20 $T=585580 236640 0 0 $X=585390 $Y=236400
X1484 1 2 473 300 1691 ICV_20 $T=595700 193120 1 0 $X=595510 $Y=190160
X1485 1 2 1686 300 1702 ICV_20 $T=598000 214880 1 0 $X=597810 $Y=211920
X1486 1 2 1686 317 1700 ICV_20 $T=598920 204000 1 0 $X=598730 $Y=201040
X1487 1 2 1688 298 1711 ICV_20 $T=605820 242080 0 0 $X=605630 $Y=241840
X1488 1 2 1688 288 1733 ICV_20 $T=614560 231200 0 0 $X=614370 $Y=230960
X1489 1 2 1743 317 1738 ICV_20 $T=627440 236640 0 0 $X=627250 $Y=236400
X1490 1 2 1770 318 1786 ICV_20 $T=639860 187680 0 0 $X=639670 $Y=187440
X1491 1 2 1743 297 1788 ICV_20 $T=639860 231200 0 0 $X=639670 $Y=230960
X1492 1 2 1802 423 1820 ICV_20 $T=657340 225760 1 0 $X=657150 $Y=222800
X1493 1 2 1816 421 1830 ICV_20 $T=662860 193120 0 0 $X=662670 $Y=192880
X1494 1 2 1816 404 1857 ICV_20 $T=674360 187680 1 0 $X=674170 $Y=184720
X1495 1 2 1866 423 1870 ICV_20 $T=685400 198560 1 0 $X=685210 $Y=195600
X1496 1 2 508 422 1887 ICV_20 $T=688620 236640 0 0 $X=688430 $Y=236400
X1497 1 2 1861 422 1895 ICV_20 $T=694140 220320 0 0 $X=693950 $Y=220080
X1498 1 2 1923 421 1944 ICV_20 $T=715760 236640 0 0 $X=715570 $Y=236400
X1499 1 2 608 7 628 ICV_21 $T=25760 231200 1 0 $X=25570 $Y=228240
X1500 1 2 626 36 645 ICV_21 $T=34040 204000 0 0 $X=33850 $Y=203760
X1501 1 2 608 20 650 ICV_21 $T=36340 231200 1 0 $X=36150 $Y=228240
X1502 1 2 653 7 671 ICV_21 $T=48300 231200 1 0 $X=48110 $Y=228240
X1503 1 2 703 11 711 ICV_21 $T=70840 193120 0 0 $X=70650 $Y=192880
X1504 1 2 760 24 779 ICV_21 $T=111780 231200 1 0 $X=111590 $Y=228240
X1505 1 2 764 12 810 ICV_21 $T=120980 209440 1 0 $X=120790 $Y=206480
X1506 1 2 116 34 855 ICV_21 $T=146280 182240 0 0 $X=146090 $Y=182000
X1507 1 2 866 13 908 ICV_21 $T=174340 209440 0 0 $X=174150 $Y=209200
X1508 1 2 127 221 227 ICV_21 $T=237820 182240 0 0 $X=237630 $Y=182000
X1509 1 2 1116 137 1135 ICV_21 $T=286580 231200 0 0 $X=286390 $Y=230960
X1510 1 2 1237 188 1251 ICV_21 $T=359720 193120 0 0 $X=359530 $Y=192880
X1511 1 2 339 181 1303 ICV_21 $T=387780 187680 0 0 $X=387590 $Y=187440
X1512 1 2 339 205 1324 ICV_21 $T=398820 187680 0 0 $X=398630 $Y=187440
X1513 1 2 360 275 1393 ICV_21 $T=431020 182240 0 0 $X=430830 $Y=182000
X1514 1 2 1391 284 1397 ICV_21 $T=436080 214880 0 0 $X=435890 $Y=214640
X1515 1 2 1440 288 1450 ICV_21 $T=462300 187680 0 0 $X=462110 $Y=187440
X1516 1 2 1456 298 1498 ICV_21 $T=485300 231200 1 0 $X=485110 $Y=228240
X1517 1 2 1563 288 1577 ICV_21 $T=528080 193120 0 0 $X=527890 $Y=192880
X1518 1 2 1563 299 1578 ICV_21 $T=528080 198560 0 0 $X=527890 $Y=198320
X1519 1 2 1598 297 1618 ICV_21 $T=548320 187680 0 0 $X=548130 $Y=187440
X1520 1 2 1643 297 1660 ICV_21 $T=571320 220320 0 0 $X=571130 $Y=220080
X1521 1 2 1802 422 1841 ICV_21 $T=665620 225760 1 0 $X=665430 $Y=222800
X1522 1 2 1867 423 1881 ICV_21 $T=683560 214880 0 0 $X=683370 $Y=214640
X1523 1 2 9 33 612 600 15 27 ICV_22 $T=20240 187680 1 0 $X=20050 $Y=184720
X1524 1 2 627 35 636 636 641 50 ICV_22 $T=32660 214880 1 0 $X=32470 $Y=211920
X1525 1 2 653 14 668 649 619 66 ICV_22 $T=48300 236640 1 0 $X=48110 $Y=233680
X1526 1 2 652 11 683 684 659 45 ICV_22 $T=57040 187680 1 0 $X=56850 $Y=184720
X1527 1 2 735 10 738 738 750 31 ICV_22 $T=88780 198560 1 0 $X=88590 $Y=195600
X1528 1 2 751 35 804 804 757 50 ICV_22 $T=118220 214880 0 0 $X=118030 $Y=214640
X1529 1 2 125 11 895 895 129 19 ICV_22 $T=170660 187680 1 0 $X=170470 $Y=184720
X1530 1 2 1002 132 1024 1024 1020 142 ICV_22 $T=230000 231200 1 0 $X=229810 $Y=228240
X1531 1 2 1066 183 1086 1084 1087 216 ICV_22 $T=264500 193120 0 0 $X=264310 $Y=192880
X1532 1 2 1173 282 1182 1182 1184 244 ICV_22 $T=323840 220320 0 0 $X=323650 $Y=220080
X1533 1 2 331 318 1267 1267 336 329 ICV_22 $T=368460 242080 1 0 $X=368270 $Y=239120
X1534 1 2 1306 278 1322 1313 1297 231 ICV_22 $T=398820 214880 0 0 $X=398630 $Y=214640
X1535 1 2 1301 299 1334 1314 1311 329 ICV_22 $T=406180 231200 0 0 $X=405990 $Y=230960
X1536 1 2 1395 267 1406 376 375 263 ICV_22 $T=441140 193120 1 0 $X=440950 $Y=190160
X1537 1 2 1395 296 1408 1407 1347 244 ICV_22 $T=441140 198560 1 0 $X=440950 $Y=195600
X1538 1 2 1369 282 1409 1409 1389 244 ICV_22 $T=441140 209440 1 0 $X=440950 $Y=206480
X1539 1 2 1412 298 1419 1398 1337 194 ICV_22 $T=449420 236640 1 0 $X=449230 $Y=233680
X1540 1 2 1481 300 1522 1522 1499 271 ICV_22 $T=497260 193120 1 0 $X=497070 $Y=190160
X1541 1 2 1508 404 1531 1531 1530 414 ICV_22 $T=504160 220320 1 0 $X=503970 $Y=217360
X1542 1 2 1582 300 1600 1600 1605 271 ICV_22 $T=539120 204000 0 0 $X=538930 $Y=203760
X1543 1 2 473 298 1697 1690 471 255 ICV_22 $T=595240 187680 0 0 $X=595050 $Y=187440
X1544 1 2 481 300 1723 1723 486 271 ICV_22 $T=608580 193120 0 0 $X=608390 $Y=192880
X1545 1 2 481 318 1725 1726 486 249 ICV_22 $T=609500 187680 1 0 $X=609310 $Y=184720
X1546 1 2 1802 405 1825 1825 1818 413 ICV_22 $T=658260 225760 0 0 $X=658070 $Y=225520
X1547 1 2 1934 421 1947 1947 1954 430 ICV_22 $T=716220 198560 0 0 $X=716030 $Y=198320
X1548 1 2 1917 404 1965 1964 1938 424 ICV_22 $T=727260 231200 1 0 $X=727070 $Y=228240
X1549 1 2 1933 404 1970 1972 1954 429 ICV_22 $T=729100 193120 1 0 $X=728910 $Y=190160
X1550 1 2 1934 423 1972 1973 1932 413 ICV_22 $T=729100 209440 1 0 $X=728910 $Y=206480
X1551 1 2 ICV_23 $T=18400 182240 1 0 $X=18210 $Y=179280
X1552 1 2 ICV_23 $T=18400 242080 1 0 $X=18210 $Y=239120
X1553 1 2 ICV_23 $T=46460 214880 1 0 $X=46270 $Y=211920
X1554 1 2 ICV_23 $T=46460 220320 1 0 $X=46270 $Y=217360
X1555 1 2 ICV_23 $T=74520 236640 1 0 $X=74330 $Y=233680
X1556 1 2 ICV_23 $T=74520 242080 1 0 $X=74330 $Y=239120
X1557 1 2 ICV_23 $T=102580 198560 1 0 $X=102390 $Y=195600
X1558 1 2 ICV_23 $T=116380 182240 0 0 $X=116190 $Y=182000
X1559 1 2 ICV_23 $T=130640 198560 1 0 $X=130450 $Y=195600
X1560 1 2 ICV_23 $T=144440 198560 0 0 $X=144250 $Y=198320
X1561 1 2 ICV_23 $T=158700 182240 1 0 $X=158510 $Y=179280
X1562 1 2 ICV_23 $T=172500 242080 0 0 $X=172310 $Y=241840
X1563 1 2 ICV_23 $T=186760 220320 1 0 $X=186570 $Y=217360
X1564 1 2 ICV_23 $T=186760 231200 1 0 $X=186570 $Y=228240
X1565 1 2 ICV_23 $T=200560 193120 0 0 $X=200370 $Y=192880
X1566 1 2 ICV_23 $T=200560 204000 0 0 $X=200370 $Y=203760
X1567 1 2 ICV_23 $T=214820 198560 1 0 $X=214630 $Y=195600
X1568 1 2 ICV_23 $T=214820 204000 1 0 $X=214630 $Y=201040
X1569 1 2 ICV_23 $T=228620 198560 0 0 $X=228430 $Y=198320
X1570 1 2 ICV_23 $T=228620 236640 0 0 $X=228430 $Y=236400
X1571 1 2 ICV_23 $T=256680 193120 0 0 $X=256490 $Y=192880
X1572 1 2 ICV_23 $T=270940 187680 1 0 $X=270750 $Y=184720
X1573 1 2 ICV_23 $T=340860 204000 0 0 $X=340670 $Y=203760
X1574 1 2 ICV_23 $T=396980 204000 0 0 $X=396790 $Y=203760
X1575 1 2 ICV_23 $T=439300 198560 1 0 $X=439110 $Y=195600
X1576 1 2 ICV_23 $T=467360 182240 1 0 $X=467170 $Y=179280
X1577 1 2 ICV_23 $T=523480 220320 1 0 $X=523290 $Y=217360
X1578 1 2 ICV_23 $T=523480 236640 1 0 $X=523290 $Y=233680
X1579 1 2 ICV_23 $T=551540 182240 1 0 $X=551350 $Y=179280
X1580 1 2 ICV_23 $T=565340 193120 0 0 $X=565150 $Y=192880
X1581 1 2 ICV_23 $T=565340 214880 0 0 $X=565150 $Y=214640
X1582 1 2 ICV_23 $T=579600 198560 1 0 $X=579410 $Y=195600
X1583 1 2 ICV_23 $T=593400 209440 0 0 $X=593210 $Y=209200
X1584 1 2 ICV_23 $T=593400 220320 0 0 $X=593210 $Y=220080
X1585 1 2 ICV_23 $T=635720 236640 1 0 $X=635530 $Y=233680
X1586 1 2 ICV_23 $T=677580 242080 0 0 $X=677390 $Y=241840
X1587 1 2 ICV_23 $T=691840 209440 1 0 $X=691650 $Y=206480
X1588 1 2 ICV_23 $T=705640 204000 0 0 $X=705450 $Y=203760
X1589 1 2 ICV_24 $T=17940 225760 1 0 $X=17750 $Y=222800
X1590 1 2 ICV_24 $T=17940 231200 1 0 $X=17750 $Y=228240
X1591 1 2 ICV_24 $T=31740 214880 0 0 $X=31550 $Y=214640
X1592 1 2 ICV_24 $T=46000 204000 1 0 $X=45810 $Y=201040
X1593 1 2 ICV_24 $T=46000 225760 1 0 $X=45810 $Y=222800
X1594 1 2 ICV_24 $T=74060 220320 1 0 $X=73870 $Y=217360
X1595 1 2 ICV_24 $T=115920 225760 0 0 $X=115730 $Y=225520
X1596 1 2 ICV_24 $T=143980 193120 0 0 $X=143790 $Y=192880
X1597 1 2 ICV_24 $T=256220 204000 0 0 $X=256030 $Y=203760
X1598 1 2 ICV_24 $T=326600 214880 1 0 $X=326410 $Y=211920
X1599 1 2 ICV_24 $T=326600 231200 1 0 $X=326410 $Y=228240
X1600 1 2 ICV_24 $T=368460 225760 0 0 $X=368270 $Y=225520
X1601 1 2 ICV_24 $T=452640 236640 0 0 $X=452450 $Y=236400
X1602 1 2 ICV_24 $T=466900 204000 1 0 $X=466710 $Y=201040
X1603 1 2 ICV_24 $T=494960 187680 1 0 $X=494770 $Y=184720
X1604 1 2 ICV_24 $T=494960 204000 1 0 $X=494770 $Y=201040
X1605 1 2 ICV_24 $T=494960 214880 1 0 $X=494770 $Y=211920
X1606 1 2 ICV_24 $T=508760 204000 0 0 $X=508570 $Y=203760
X1607 1 2 ICV_24 $T=635260 209440 1 0 $X=635070 $Y=206480
X1608 1 2 ICV_24 $T=677120 182240 0 0 $X=676930 $Y=182000
X1609 1 2 23 2 601 1 sky130_fd_sc_hd__inv_1 $T=26680 193120 1 0 $X=26490 $Y=190160
X1610 1 2 37 2 603 1 sky130_fd_sc_hd__inv_1 $T=26680 209440 1 0 $X=26490 $Y=206480
X1611 1 2 52 2 619 1 sky130_fd_sc_hd__inv_1 $T=38180 236640 0 0 $X=37990 $Y=236400
X1612 1 2 54 2 641 1 sky130_fd_sc_hd__inv_1 $T=42320 209440 0 0 $X=42130 $Y=209200
X1613 1 2 59 2 640 1 sky130_fd_sc_hd__inv_1 $T=46000 198560 1 0 $X=45810 $Y=195600
X1614 1 2 71 2 659 1 sky130_fd_sc_hd__inv_1 $T=63940 182240 1 0 $X=63750 $Y=179280
X1615 1 2 64 2 672 1 sky130_fd_sc_hd__inv_1 $T=73140 242080 1 0 $X=72950 $Y=239120
X1616 1 2 84 2 710 1 sky130_fd_sc_hd__inv_1 $T=87860 187680 0 0 $X=87670 $Y=187440
X1617 1 2 77 2 694 1 sky130_fd_sc_hd__inv_1 $T=88780 214880 1 0 $X=88590 $Y=211920
X1618 1 2 91 2 691 1 sky130_fd_sc_hd__inv_1 $T=101200 204000 0 0 $X=101010 $Y=203760
X1619 1 2 83 2 87 1 sky130_fd_sc_hd__inv_1 $T=104420 242080 0 0 $X=104230 $Y=241840
X1620 1 2 102 2 773 1 sky130_fd_sc_hd__inv_1 $T=124200 236640 1 0 $X=124010 $Y=233680
X1621 1 2 106 2 757 1 sky130_fd_sc_hd__inv_1 $T=129720 209440 0 0 $X=129530 $Y=209200
X1622 1 2 107 2 808 1 sky130_fd_sc_hd__inv_1 $T=132480 242080 1 0 $X=132290 $Y=239120
X1623 1 2 111 2 780 1 sky130_fd_sc_hd__inv_1 $T=134320 198560 0 0 $X=134130 $Y=198320
X1624 1 2 101 2 792 1 sky130_fd_sc_hd__inv_1 $T=143520 187680 1 0 $X=143330 $Y=184720
X1625 1 2 114 2 807 1 sky130_fd_sc_hd__inv_1 $T=153640 198560 1 0 $X=153450 $Y=195600
X1626 1 2 115 2 824 1 sky130_fd_sc_hd__inv_1 $T=160540 242080 0 0 $X=160350 $Y=241840
X1627 1 2 126 2 882 1 sky130_fd_sc_hd__inv_1 $T=171120 242080 0 0 $X=170930 $Y=241840
X1628 1 2 121 2 868 1 sky130_fd_sc_hd__inv_1 $T=178020 193120 1 0 $X=177830 $Y=190160
X1629 1 2 123 2 881 1 sky130_fd_sc_hd__inv_1 $T=182160 204000 0 0 $X=181970 $Y=203760
X1630 1 2 42 2 170 1 sky130_fd_sc_hd__inv_1 $T=200560 242080 0 0 $X=200370 $Y=241840
X1631 1 2 169 2 909 1 sky130_fd_sc_hd__inv_1 $T=206540 198560 1 0 $X=206350 $Y=195600
X1632 1 2 175 2 929 1 sky130_fd_sc_hd__inv_1 $T=208840 209440 0 0 $X=208650 $Y=209200
X1633 1 2 179 2 177 1 sky130_fd_sc_hd__inv_1 $T=212980 182240 0 0 $X=212790 $Y=182000
X1634 1 2 64 2 974 1 sky130_fd_sc_hd__inv_1 $T=218960 236640 0 0 $X=218770 $Y=236400
X1635 1 2 59 2 966 1 sky130_fd_sc_hd__inv_1 $T=228160 198560 1 0 $X=227970 $Y=195600
X1636 1 2 23 2 983 1 sky130_fd_sc_hd__inv_1 $T=228620 187680 0 0 $X=228430 $Y=187440
X1637 1 2 37 2 985 1 sky130_fd_sc_hd__inv_1 $T=235980 209440 1 0 $X=235790 $Y=206480
X1638 1 2 83 2 1020 1 sky130_fd_sc_hd__inv_1 $T=236900 242080 0 0 $X=236710 $Y=241840
X1639 1 2 77 2 1046 1 sky130_fd_sc_hd__inv_1 $T=255760 209440 0 0 $X=255570 $Y=209200
X1640 1 2 72 2 1055 1 sky130_fd_sc_hd__inv_1 $T=256680 236640 0 0 $X=256490 $Y=236400
X1641 1 2 84 2 224 1 sky130_fd_sc_hd__inv_1 $T=260360 187680 1 0 $X=260170 $Y=184720
X1642 1 2 54 2 1078 1 sky130_fd_sc_hd__inv_1 $T=270940 214880 1 0 $X=270750 $Y=211920
X1643 1 2 67 2 1087 1 sky130_fd_sc_hd__inv_1 $T=275080 193120 1 0 $X=274890 $Y=190160
X1644 1 2 102 2 1100 1 sky130_fd_sc_hd__inv_1 $T=293940 236640 0 0 $X=293750 $Y=236400
X1645 1 2 91 2 1091 1 sky130_fd_sc_hd__inv_1 $T=294400 204000 1 0 $X=294210 $Y=201040
X1646 1 2 115 2 1138 1 sky130_fd_sc_hd__inv_1 $T=299000 242080 1 0 $X=298810 $Y=239120
X1647 1 2 106 2 1136 1 sky130_fd_sc_hd__inv_1 $T=310500 209440 0 0 $X=310310 $Y=209200
X1648 1 2 121 2 1155 1 sky130_fd_sc_hd__inv_1 $T=312800 193120 0 0 $X=312610 $Y=192880
X1649 1 2 111 2 1172 1 sky130_fd_sc_hd__inv_1 $T=322920 204000 0 0 $X=322730 $Y=203760
X1650 1 2 114 2 1201 1 sky130_fd_sc_hd__inv_1 $T=345920 198560 1 0 $X=345730 $Y=195600
X1651 1 2 301 2 1184 1 sky130_fd_sc_hd__inv_1 $T=346840 214880 0 0 $X=346650 $Y=214640
X1652 1 2 307 2 1212 1 sky130_fd_sc_hd__inv_1 $T=356960 220320 1 0 $X=356770 $Y=217360
X1653 1 2 295 2 1193 1 sky130_fd_sc_hd__inv_1 $T=357420 182240 1 0 $X=357230 $Y=179280
X1654 1 2 315 2 1239 1 sky130_fd_sc_hd__inv_1 $T=374440 214880 1 0 $X=374250 $Y=211920
X1655 1 2 118 2 1268 1 sky130_fd_sc_hd__inv_1 $T=380420 198560 0 0 $X=380230 $Y=198320
X1656 1 2 334 2 1248 1 sky130_fd_sc_hd__inv_1 $T=383180 225760 1 0 $X=382990 $Y=222800
X1657 1 2 334 2 1280 1 sky130_fd_sc_hd__inv_1 $T=396060 220320 1 0 $X=395870 $Y=217360
X1658 1 2 340 2 336 1 sky130_fd_sc_hd__inv_1 $T=396520 242080 1 0 $X=396330 $Y=239120
X1659 1 2 112 2 351 1 sky130_fd_sc_hd__inv_1 $T=399740 182240 0 0 $X=399550 $Y=182000
X1660 1 2 356 2 1311 1 sky130_fd_sc_hd__inv_1 $T=413080 231200 1 0 $X=412890 $Y=228240
X1661 1 2 353 2 1327 1 sky130_fd_sc_hd__inv_1 $T=418140 204000 1 0 $X=417950 $Y=201040
X1662 1 2 363 2 1366 1 sky130_fd_sc_hd__inv_1 $T=433320 225760 0 0 $X=433130 $Y=225520
X1663 1 2 356 2 1351 1 sky130_fd_sc_hd__inv_1 $T=434240 187680 1 0 $X=434050 $Y=184720
X1664 1 2 368 2 364 1 sky130_fd_sc_hd__inv_1 $T=438380 182240 1 0 $X=438190 $Y=179280
X1665 1 2 369 2 370 1 sky130_fd_sc_hd__inv_1 $T=448500 225760 1 0 $X=448310 $Y=222800
X1666 1 2 363 2 1389 1 sky130_fd_sc_hd__inv_1 $T=452640 204000 0 0 $X=452450 $Y=203760
X1667 1 2 365 2 1337 1 sky130_fd_sc_hd__inv_1 $T=455860 220320 0 0 $X=455670 $Y=220080
X1668 1 2 367 2 1347 1 sky130_fd_sc_hd__inv_1 $T=462300 193120 0 0 $X=462110 $Y=192880
X1669 1 2 378 2 1422 1 sky130_fd_sc_hd__inv_1 $T=473800 231200 0 0 $X=473610 $Y=230960
X1670 1 2 380 2 1423 1 sky130_fd_sc_hd__inv_1 $T=477020 220320 0 0 $X=476830 $Y=220080
X1671 1 2 368 2 1438 1 sky130_fd_sc_hd__inv_1 $T=480240 198560 0 0 $X=480050 $Y=198320
X1672 1 2 381 2 1449 1 sky130_fd_sc_hd__inv_1 $T=481160 182240 0 0 $X=480970 $Y=182000
X1673 1 2 399 2 393 1 sky130_fd_sc_hd__inv_1 $T=492660 242080 0 0 $X=492470 $Y=241840
X1674 1 2 402 2 392 1 sky130_fd_sc_hd__inv_1 $T=494500 182240 1 0 $X=494310 $Y=179280
X1675 1 2 390 2 1477 1 sky130_fd_sc_hd__inv_1 $T=498640 225760 0 0 $X=498450 $Y=225520
X1676 1 2 400 2 1491 1 sky130_fd_sc_hd__inv_1 $T=504160 198560 1 0 $X=503970 $Y=195600
X1677 1 2 397 2 1499 1 sky130_fd_sc_hd__inv_1 $T=507380 187680 1 0 $X=507190 $Y=184720
X1678 1 2 394 2 1465 1 sky130_fd_sc_hd__inv_1 $T=508760 209440 0 0 $X=508570 $Y=209200
X1679 1 2 353 2 1530 1 sky130_fd_sc_hd__inv_1 $T=513360 214880 0 0 $X=513170 $Y=214640
X1680 1 2 340 2 1520 1 sky130_fd_sc_hd__inv_1 $T=522560 231200 0 0 $X=522370 $Y=230960
X1681 1 2 428 2 1534 1 sky130_fd_sc_hd__inv_1 $T=525780 193120 1 0 $X=525590 $Y=190160
X1682 1 2 315 2 420 1 sky130_fd_sc_hd__inv_1 $T=527620 242080 0 0 $X=527430 $Y=241840
X1683 1 2 356 2 1568 1 sky130_fd_sc_hd__inv_1 $T=536360 225760 0 0 $X=536170 $Y=225520
X1684 1 2 369 2 1580 1 sky130_fd_sc_hd__inv_1 $T=540040 220320 1 0 $X=539850 $Y=217360
X1685 1 2 442 2 1605 1 sky130_fd_sc_hd__inv_1 $T=561200 198560 0 0 $X=561010 $Y=198320
X1686 1 2 448 2 1636 1 sky130_fd_sc_hd__inv_1 $T=567180 209440 0 0 $X=566990 $Y=209200
X1687 1 2 457 2 460 1 sky130_fd_sc_hd__inv_1 $T=579600 236640 0 0 $X=579410 $Y=236400
X1688 1 2 461 2 1653 1 sky130_fd_sc_hd__inv_1 $T=581900 225760 0 0 $X=581710 $Y=225520
X1689 1 2 464 2 1652 1 sky130_fd_sc_hd__inv_1 $T=592020 209440 0 0 $X=591830 $Y=209200
X1690 1 2 446 2 1649 1 sky130_fd_sc_hd__inv_1 $T=593400 193120 0 0 $X=593210 $Y=192880
X1691 1 2 472 2 1667 1 sky130_fd_sc_hd__inv_1 $T=594320 182240 1 0 $X=594130 $Y=179280
X1692 1 2 476 2 1704 1 sky130_fd_sc_hd__inv_1 $T=609500 198560 1 0 $X=609310 $Y=195600
X1693 1 2 469 2 1699 1 sky130_fd_sc_hd__inv_1 $T=614100 225760 1 0 $X=613910 $Y=222800
X1694 1 2 470 2 1713 1 sky130_fd_sc_hd__inv_1 $T=620540 236640 0 0 $X=620350 $Y=236400
X1695 1 2 487 2 1736 1 sky130_fd_sc_hd__inv_1 $T=631580 198560 0 0 $X=631390 $Y=198320
X1696 1 2 482 2 1745 1 sky130_fd_sc_hd__inv_1 $T=638020 220320 1 0 $X=637830 $Y=217360
X1697 1 2 498 2 1739 1 sky130_fd_sc_hd__inv_1 $T=648600 231200 1 0 $X=648410 $Y=228240
X1698 1 2 496 2 1783 1 sky130_fd_sc_hd__inv_1 $T=655500 198560 1 0 $X=655310 $Y=195600
X1699 1 2 497 2 1787 1 sky130_fd_sc_hd__inv_1 $T=658260 182240 0 0 $X=658070 $Y=182000
X1700 1 2 494 2 1759 1 sky130_fd_sc_hd__inv_1 $T=662400 209440 1 0 $X=662210 $Y=206480
X1701 1 2 385 2 1812 1 sky130_fd_sc_hd__inv_1 $T=662860 236640 1 0 $X=662670 $Y=233680
X1702 1 2 457 2 1818 1 sky130_fd_sc_hd__inv_1 $T=663780 220320 1 0 $X=663590 $Y=217360
X1703 1 2 428 2 1831 1 sky130_fd_sc_hd__inv_1 $T=672980 187680 1 0 $X=672790 $Y=184720
X1704 1 2 400 2 1826 1 sky130_fd_sc_hd__inv_1 $T=675280 198560 0 0 $X=675090 $Y=198320
X1705 1 2 470 2 1844 1 sky130_fd_sc_hd__inv_1 $T=676200 225760 1 0 $X=676010 $Y=222800
X1706 1 2 494 2 1865 1 sky130_fd_sc_hd__inv_1 $T=684480 198560 0 0 $X=684290 $Y=198320
X1707 1 2 446 2 506 1 sky130_fd_sc_hd__inv_1 $T=691840 182240 1 0 $X=691650 $Y=179280
X1708 1 2 464 2 1886 1 sky130_fd_sc_hd__inv_1 $T=698740 214880 0 0 $X=698550 $Y=214640
X1709 1 2 462 2 509 1 sky130_fd_sc_hd__inv_1 $T=699660 242080 1 0 $X=699470 $Y=239120
X1710 1 2 496 2 1885 1 sky130_fd_sc_hd__inv_1 $T=707480 187680 0 0 $X=707290 $Y=187440
X1711 1 2 461 2 1938 1 sky130_fd_sc_hd__inv_1 $T=719440 225760 1 0 $X=719250 $Y=222800
X1712 1 2 498 2 510 1 sky130_fd_sc_hd__inv_1 $T=725880 231200 1 0 $X=725690 $Y=228240
X1713 1 2 489 2 519 1 sky130_fd_sc_hd__inv_1 $T=726340 242080 0 0 $X=726150 $Y=241840
X1714 1 2 497 2 1901 1 sky130_fd_sc_hd__inv_1 $T=729100 187680 1 0 $X=728910 $Y=184720
X1715 1 2 448 2 1932 1 sky130_fd_sc_hd__inv_1 $T=729100 214880 1 0 $X=728910 $Y=211920
X1716 1 2 482 2 1954 1 sky130_fd_sc_hd__inv_1 $T=730020 198560 1 0 $X=729830 $Y=195600
X1717 1 2 ICV_25 $T=30360 182240 0 0 $X=30170 $Y=182000
X1718 1 2 ICV_25 $T=44620 182240 1 0 $X=44430 $Y=179280
X1719 1 2 ICV_25 $T=100740 236640 1 0 $X=100550 $Y=233680
X1720 1 2 ICV_25 $T=156860 225760 1 0 $X=156670 $Y=222800
X1721 1 2 ICV_25 $T=282900 225760 0 0 $X=282710 $Y=225520
X1722 1 2 ICV_25 $T=297160 198560 1 0 $X=296970 $Y=195600
X1723 1 2 ICV_25 $T=325220 187680 1 0 $X=325030 $Y=184720
X1724 1 2 ICV_25 $T=325220 193120 1 0 $X=325030 $Y=190160
X1725 1 2 ICV_25 $T=409400 193120 1 0 $X=409210 $Y=190160
X1726 1 2 ICV_25 $T=409400 236640 1 0 $X=409210 $Y=233680
X1727 1 2 ICV_25 $T=465520 220320 1 0 $X=465330 $Y=217360
X1728 1 2 ICV_25 $T=493580 220320 1 0 $X=493390 $Y=217360
X1729 1 2 ICV_25 $T=493580 236640 1 0 $X=493390 $Y=233680
X1730 1 2 ICV_25 $T=563500 187680 0 0 $X=563310 $Y=187440
X1731 1 2 ICV_25 $T=605820 214880 1 0 $X=605630 $Y=211920
X1732 1 2 ICV_25 $T=647680 187680 0 0 $X=647490 $Y=187440
X1733 1 2 ICV_25 $T=647680 231200 0 0 $X=647490 $Y=230960
X1734 1 2 ICV_25 $T=675740 204000 0 0 $X=675550 $Y=203760
X1735 1 2 ICV_25 $T=675740 236640 0 0 $X=675550 $Y=236400
X1736 1 2 592 15 19 ICV_26 $T=15180 193120 1 0 $X=14990 $Y=190160
X1737 1 2 599 603 28 ICV_26 $T=17940 220320 0 0 $X=17750 $Y=220080
X1738 1 2 616 619 46 ICV_26 $T=28980 225760 0 0 $X=28790 $Y=225520
X1739 1 2 623 603 50 ICV_26 $T=30820 209440 1 0 $X=30630 $Y=206480
X1740 1 2 661 640 19 ICV_26 $T=54280 209440 0 0 $X=54090 $Y=209200
X1741 1 2 70 69 18 ICV_26 $T=62100 242080 0 0 $X=61910 $Y=241840
X1742 1 2 683 659 19 ICV_26 $T=65320 182240 1 0 $X=65130 $Y=179280
X1743 1 2 713 73 18 ICV_26 $T=81420 225760 0 0 $X=81230 $Y=225520
X1744 1 2 805 807 19 ICV_26 $T=127420 193120 1 0 $X=127230 $Y=190160
X1745 1 2 803 780 50 ICV_26 $T=127420 204000 1 0 $X=127230 $Y=201040
X1746 1 2 820 792 28 ICV_26 $T=139380 193120 0 0 $X=139190 $Y=192880
X1747 1 2 830 808 18 ICV_26 $T=140760 225760 0 0 $X=140570 $Y=225520
X1748 1 2 840 807 45 ICV_26 $T=144900 220320 1 0 $X=144710 $Y=217360
X1749 1 2 851 119 28 ICV_26 $T=154100 182240 1 0 $X=153910 $Y=179280
X1750 1 2 853 119 27 ICV_26 $T=155940 187680 0 0 $X=155750 $Y=187440
X1751 1 2 122 119 48 ICV_26 $T=156860 182240 0 0 $X=156670 $Y=182000
X1752 1 2 876 881 48 ICV_26 $T=169280 214880 0 0 $X=169090 $Y=214640
X1753 1 2 907 909 19 ICV_26 $T=183540 204000 1 0 $X=183350 $Y=201040
X1754 1 2 154 158 28 ICV_26 $T=191360 182240 1 0 $X=191170 $Y=179280
X1755 1 2 964 966 185 ICV_26 $T=212980 204000 0 0 $X=212790 $Y=203760
X1756 1 2 978 193 196 ICV_26 $T=221720 182240 0 0 $X=221530 $Y=182000
X1757 1 2 1011 985 216 ICV_26 $T=235980 214880 1 0 $X=235790 $Y=211920
X1758 1 2 1023 1020 135 ICV_26 $T=238280 225760 0 0 $X=238090 $Y=225520
X1759 1 2 1056 1055 156 ICV_26 $T=258520 231200 0 0 $X=258330 $Y=230960
X1760 1 2 1063 224 195 ICV_26 $T=260360 193120 1 0 $X=260170 $Y=190160
X1761 1 2 1068 234 219 ICV_26 $T=265880 187680 0 0 $X=265690 $Y=187440
X1762 1 2 1073 1055 135 ICV_26 $T=267720 231200 1 0 $X=267530 $Y=228240
X1763 1 2 1088 1091 219 ICV_26 $T=273700 220320 0 0 $X=273510 $Y=220080
X1764 1 2 1120 258 185 ICV_26 $T=293480 187680 1 0 $X=293290 $Y=184720
X1765 1 2 1133 1136 196 ICV_26 $T=295780 204000 1 0 $X=295590 $Y=201040
X1766 1 2 1142 1138 156 ICV_26 $T=303600 236640 1 0 $X=303410 $Y=233680
X1767 1 2 1165 1172 198 ICV_26 $T=322000 214880 1 0 $X=321810 $Y=211920
X1768 1 2 1170 1172 196 ICV_26 $T=322460 193120 0 0 $X=322270 $Y=192880
X1769 1 2 1171 1172 195 ICV_26 $T=323840 204000 1 0 $X=323650 $Y=201040
X1770 1 2 320 311 196 ICV_26 $T=358340 182240 0 0 $X=358150 $Y=182000
X1771 1 2 1225 1193 212 ICV_26 $T=358340 187680 0 0 $X=358150 $Y=187440
X1772 1 2 1251 1255 195 ICV_26 $T=370760 193120 0 0 $X=370570 $Y=192880
X1773 1 2 1250 1255 196 ICV_26 $T=372600 187680 1 0 $X=372410 $Y=184720
X1774 1 2 1257 1239 244 ICV_26 $T=373520 214880 0 0 $X=373330 $Y=214640
X1775 1 2 1307 1297 252 ICV_26 $T=398820 198560 0 0 $X=398630 $Y=198320
X1776 1 2 1316 355 329 ICV_26 $T=407100 242080 1 0 $X=406910 $Y=239120
X1777 1 2 1317 355 251 ICV_26 $T=407100 242080 0 0 $X=406910 $Y=241840
X1778 1 2 1323 351 196 ICV_26 $T=408020 187680 1 0 $X=407830 $Y=184720
X1779 1 2 1322 1297 261 ICV_26 $T=408020 214880 1 0 $X=407830 $Y=211920
X1780 1 2 1334 1311 238 ICV_26 $T=414460 231200 1 0 $X=414270 $Y=228240
X1781 1 2 1336 1337 263 ICV_26 $T=415380 225760 1 0 $X=415190 $Y=222800
X1782 1 2 1350 1337 232 ICV_26 $T=421820 214880 0 0 $X=421630 $Y=214640
X1783 1 2 1364 1366 251 ICV_26 $T=427340 231200 1 0 $X=427150 $Y=228240
X1784 1 2 1441 1423 285 ICV_26 $T=464140 225760 1 0 $X=463950 $Y=222800
X1785 1 2 1439 1422 238 ICV_26 $T=464140 242080 1 0 $X=463950 $Y=239120
X1786 1 2 1447 1449 271 ICV_26 $T=469200 198560 1 0 $X=469010 $Y=195600
X1787 1 2 1448 1422 255 ICV_26 $T=469200 236640 1 0 $X=469010 $Y=233680
X1788 1 2 1507 1465 231 ICV_26 $T=499560 220320 1 0 $X=499370 $Y=217360
X1789 1 2 1552 1546 430 ICV_26 $T=523940 214880 0 0 $X=523750 $Y=214640
X1790 1 2 1618 443 249 ICV_26 $T=558900 187680 0 0 $X=558710 $Y=187440
X1791 1 2 1635 1636 285 ICV_26 $T=568100 225760 1 0 $X=567910 $Y=222800
X1792 1 2 1651 1653 329 ICV_26 $T=576380 231200 1 0 $X=576190 $Y=228240
X1793 1 2 1661 1653 285 ICV_26 $T=580980 236640 0 0 $X=580790 $Y=236400
X1794 1 2 1665 1667 329 ICV_26 $T=587880 187680 0 0 $X=587690 $Y=187440
X1795 1 2 1691 471 271 ICV_26 $T=603520 193120 1 0 $X=603330 $Y=190160
X1796 1 2 1692 471 249 ICV_26 $T=603980 187680 1 0 $X=603790 $Y=184720
X1797 1 2 1709 1713 329 ICV_26 $T=609960 231200 0 0 $X=609770 $Y=230960
X1798 1 2 1708 1713 271 ICV_26 $T=610880 236640 0 0 $X=610690 $Y=236400
X1799 1 2 1730 1736 249 ICV_26 $T=621000 209440 1 0 $X=620810 $Y=206480
X1800 1 2 1779 501 430 ICV_26 $T=645380 182240 0 0 $X=645190 $Y=182000
X1801 1 2 1780 1787 255 ICV_26 $T=645840 198560 1 0 $X=645650 $Y=195600
X1802 1 2 1811 1812 429 ICV_26 $T=660560 231200 1 0 $X=660370 $Y=228240
X1803 1 2 1830 1831 430 ICV_26 $T=669300 193120 1 0 $X=669110 $Y=190160
X1804 1 2 1833 1812 415 ICV_26 $T=671140 236640 0 0 $X=670950 $Y=236400
X1805 1 2 1841 1818 427 ICV_26 $T=674360 225760 0 0 $X=674170 $Y=225520
X1806 1 2 1851 506 427 ICV_26 $T=679420 182240 0 0 $X=679230 $Y=182000
X1807 1 2 1852 1826 413 ICV_26 $T=679420 214880 1 0 $X=679230 $Y=211920
X1808 1 2 1870 1865 429 ICV_26 $T=688620 204000 1 0 $X=688430 $Y=201040
X1809 1 2 1879 1886 413 ICV_26 $T=694140 214880 0 0 $X=693950 $Y=214640
X1810 1 2 1899 1865 412 ICV_26 $T=704260 209440 1 0 $X=704070 $Y=206480
X1811 1 2 1945 510 424 ICV_26 $T=723120 231200 0 0 $X=722930 $Y=230960
X1812 1 2 1967 518 413 ICV_26 $T=737380 182240 1 0 $X=737190 $Y=179280
X1813 1 2 526 517 413 ICV_26 $T=737380 242080 1 0 $X=737190 $Y=239120
X1814 1 2 587 7 590 ICV_28 $T=6900 231200 0 0 $X=6710 $Y=230960
X1815 1 2 587 6 591 ICV_28 $T=6900 236640 1 0 $X=6710 $Y=233680
X1816 1 2 587 5 586 ICV_28 $T=6900 242080 0 0 $X=6710 $Y=241840
X1817 1 2 608 24 616 ICV_28 $T=27600 236640 1 0 $X=27410 $Y=233680
X1818 1 2 866 12 885 ICV_28 $T=164680 214880 1 0 $X=164490 $Y=211920
X1819 1 2 127 44 894 ICV_28 $T=171120 220320 1 0 $X=170930 $Y=217360
X1820 1 2 127 45 931 ICV_28 $T=188600 220320 0 0 $X=188410 $Y=220080
X1821 1 2 159 137 936 ICV_28 $T=191820 225760 0 0 $X=191630 $Y=225520
X1822 1 2 1028 199 1039 ICV_28 $T=241960 198560 0 0 $X=241770 $Y=198320
X1823 1 2 127 231 925 ICV_28 $T=248400 225760 0 0 $X=248210 $Y=225520
X1824 1 2 1028 181 1061 ICV_28 $T=252080 204000 1 0 $X=251890 $Y=201040
X1825 1 2 228 201 1068 ICV_28 $T=261740 187680 1 0 $X=261550 $Y=184720
X1826 1 2 1108 181 1126 ICV_28 $T=286580 187680 0 0 $X=286390 $Y=187440
X1827 1 2 127 252 981 ICV_28 $T=286580 220320 0 0 $X=286390 $Y=220080
X1828 1 2 1108 205 1132 ICV_28 $T=287960 198560 1 0 $X=287770 $Y=195600
X1829 1 2 1156 188 1171 ICV_28 $T=314640 204000 1 0 $X=314450 $Y=201040
X1830 1 2 1173 280 1178 ICV_28 $T=322000 209440 0 0 $X=321810 $Y=209200
X1831 1 2 127 285 1157 ICV_28 $T=322920 231200 0 0 $X=322730 $Y=230960
X1832 1 2 1173 275 1181 ICV_28 $T=323840 214880 0 0 $X=323650 $Y=214640
X1833 1 2 1197 200 1225 ICV_28 $T=347300 198560 1 0 $X=347110 $Y=195600
X1834 1 2 1197 199 1230 ICV_28 $T=349140 187680 0 0 $X=348950 $Y=187440
X1835 1 2 1234 275 1243 ICV_28 $T=357880 204000 0 0 $X=357690 $Y=203760
X1836 1 2 1249 299 1283 ICV_28 $T=378120 231200 0 0 $X=377930 $Y=230960
X1837 1 2 339 188 349 ICV_28 $T=388700 182240 0 0 $X=388510 $Y=182000
X1838 1 2 354 318 1316 ICV_28 $T=397900 242080 1 0 $X=397710 $Y=239120
X1839 1 2 1306 275 1307 ICV_28 $T=398820 209440 0 0 $X=398630 $Y=209200
X1840 1 2 1369 279 1413 ICV_28 $T=443440 204000 0 0 $X=443250 $Y=203760
X1841 1 2 1551 405 1570 ICV_28 $T=525320 231200 1 0 $X=525130 $Y=228240
X1842 1 2 1576 406 1607 ICV_28 $T=543720 225760 1 0 $X=543530 $Y=222800
X1843 1 2 1637 297 1646 ICV_28 $T=567180 204000 0 0 $X=566990 $Y=203760
X1844 1 2 463 288 1664 ICV_28 $T=578220 182240 0 0 $X=578030 $Y=182000
X1845 1 2 1637 317 1683 ICV_28 $T=585120 204000 0 0 $X=584930 $Y=203760
X1846 1 2 1743 286 1763 ICV_28 $T=626520 236640 1 0 $X=626330 $Y=233680
X1847 1 2 1727 298 1764 ICV_28 $T=627440 214880 0 0 $X=627250 $Y=214640
X1848 1 2 499 421 1779 ICV_28 $T=637560 182240 1 0 $X=637370 $Y=179280
X1849 1 2 1795 422 1840 ICV_28 $T=665620 236640 1 0 $X=665430 $Y=233680
X1850 1 2 1867 405 1879 ICV_28 $T=684020 214880 1 0 $X=683830 $Y=211920
X1851 1 2 513 403 1939 ICV_28 $T=712080 182240 1 0 $X=711890 $Y=179280
X1852 1 2 608 5 625 ICV_29 $T=23920 236640 0 0 $X=23730 $Y=236400
X1853 1 2 49 35 58 ICV_29 $T=34960 182240 1 0 $X=34770 $Y=179280
X1854 1 2 89 34 100 ICV_29 $T=104420 182240 0 0 $X=104230 $Y=182000
X1855 1 2 793 24 811 ICV_29 $T=122360 231200 1 0 $X=122170 $Y=228240
X1856 1 2 793 21 814 ICV_29 $T=125580 242080 0 0 $X=125390 $Y=241840
X1857 1 2 116 13 853 ICV_29 $T=146280 187680 0 0 $X=146090 $Y=187440
X1858 1 2 127 66 886 ICV_29 $T=164220 231200 0 0 $X=164030 $Y=230960
X1859 1 2 897 33 920 ICV_29 $T=181700 182240 0 0 $X=181510 $Y=182000
X1860 1 2 1002 137 1023 ICV_29 $T=230460 231200 0 0 $X=230270 $Y=230960
X1861 1 2 1048 147 1064 ICV_29 $T=252080 236640 1 0 $X=251890 $Y=233680
X1862 1 2 1062 181 1070 ICV_29 $T=258520 214880 0 0 $X=258330 $Y=214640
X1863 1 2 262 200 1151 ICV_29 $T=300840 187680 1 0 $X=300650 $Y=184720
X1864 1 2 1183 182 1208 ICV_29 $T=336260 198560 1 0 $X=336070 $Y=195600
X1865 1 2 1342 278 1357 ICV_29 $T=416760 209440 0 0 $X=416570 $Y=209200
X1866 1 2 1339 296 1382 ICV_29 $T=426880 187680 0 0 $X=426690 $Y=187440
X1867 1 2 1391 296 1411 ICV_29 $T=448500 220320 1 0 $X=448310 $Y=217360
X1868 1 2 1440 297 1467 ICV_29 $T=471500 193120 0 0 $X=471310 $Y=192880
X1869 1 2 1526 318 1557 ICV_29 $T=518420 198560 0 0 $X=518230 $Y=198320
X1870 1 2 1642 297 1658 ICV_29 $T=571320 231200 0 0 $X=571130 $Y=230960
X1871 1 2 1686 298 1698 ICV_29 $T=595240 209440 0 0 $X=595050 $Y=209200
X1872 1 2 1743 300 1790 ICV_29 $T=638940 225760 0 0 $X=638750 $Y=225520
X1873 1 2 499 422 503 ICV_29 $T=655040 182240 1 0 $X=654850 $Y=179280
X1874 1 2 505 409 1896 ICV_29 $T=693680 182240 1 0 $X=693490 $Y=179280
X1875 1 2 1866 409 1909 ICV_29 $T=697820 204000 1 0 $X=697630 $Y=201040
X1876 1 2 590 3 18 591 3 32 ICV_30 $T=15640 236640 0 0 $X=15450 $Y=236400
X1877 1 2 604 601 28 602 601 31 ICV_30 $T=19320 198560 0 0 $X=19130 $Y=198320
X1878 1 2 638 619 32 650 619 39 ICV_30 $T=41400 225760 0 0 $X=41210 $Y=225520
X1879 1 2 631 57 27 647 57 31 ICV_30 $T=42320 193120 0 0 $X=42130 $Y=192880
X1880 1 2 62 57 44 644 57 45 ICV_30 $T=48300 182240 1 0 $X=48110 $Y=179280
X1881 1 2 645 640 48 655 640 28 ICV_30 $T=48300 204000 1 0 $X=48110 $Y=201040
X1882 1 2 714 710 45 726 710 48 ICV_30 $T=80960 209440 0 0 $X=80770 $Y=209200
X1883 1 2 745 691 44 736 691 31 ICV_30 $T=104420 209440 1 0 $X=104230 $Y=206480
X1884 1 2 744 691 50 778 780 19 ICV_30 $T=109480 198560 0 0 $X=109290 $Y=198320
X1885 1 2 763 98 18 779 773 46 ICV_30 $T=109480 231200 0 0 $X=109290 $Y=230960
X1886 1 2 789 780 27 786 780 45 ICV_30 $T=121440 204000 0 0 $X=121250 $Y=203760
X1887 1 2 841 834 48 839 807 31 ICV_30 $T=146280 220320 0 0 $X=146090 $Y=220080
X1888 1 2 847 824 18 846 824 39 ICV_30 $T=149960 231200 1 0 $X=149770 $Y=228240
X1889 1 2 844 807 28 858 807 48 ICV_30 $T=152260 204000 0 0 $X=152070 $Y=203760
X1890 1 2 856 834 27 857 834 45 ICV_30 $T=155940 220320 0 0 $X=155750 $Y=220080
X1891 1 2 867 868 31 873 868 48 ICV_30 $T=163300 198560 0 0 $X=163110 $Y=198320
X1892 1 2 869 129 45 878 129 28 ICV_30 $T=165600 193120 1 0 $X=165410 $Y=190160
X1893 1 2 872 868 50 901 868 45 ICV_30 $T=179400 198560 1 0 $X=179210 $Y=195600
X1894 1 2 910 881 44 918 909 45 ICV_30 $T=184920 204000 0 0 $X=184730 $Y=203760
X1895 1 2 915 882 152 160 164 135 ICV_30 $T=188140 242080 0 0 $X=187950 $Y=241840
X1896 1 2 914 882 155 162 164 152 ICV_30 $T=188600 231200 1 0 $X=188410 $Y=228240
X1897 1 2 916 882 156 163 164 157 ICV_30 $T=188600 236640 1 0 $X=188410 $Y=233680
X1898 1 2 919 909 44 927 909 50 ICV_30 $T=190900 193120 1 0 $X=190710 $Y=190160
X1899 1 2 935 929 31 951 909 31 ICV_30 $T=202400 204000 0 0 $X=202210 $Y=203760
X1900 1 2 932 170 156 946 170 142 ICV_30 $T=202400 231200 0 0 $X=202210 $Y=230960
X1901 1 2 933 170 155 176 170 151 ICV_30 $T=202400 242080 0 0 $X=202210 $Y=241840
X1902 1 2 942 909 28 950 909 27 ICV_30 $T=203320 198560 0 0 $X=203130 $Y=198320
X1903 1 2 998 974 142 996 974 157 ICV_30 $T=228160 236640 1 0 $X=227970 $Y=233680
X1904 1 2 1016 966 219 1040 224 212 ICV_30 $T=248400 193120 0 0 $X=248210 $Y=192880
X1905 1 2 1083 1087 211 1076 1078 219 ICV_30 $T=272780 204000 0 0 $X=272590 $Y=203760
X1906 1 2 1080 1055 151 1081 1055 153 ICV_30 $T=272780 236640 1 0 $X=272590 $Y=233680
X1907 1 2 1097 1087 219 1102 1087 185 ICV_30 $T=277840 187680 1 0 $X=277650 $Y=184720
X1908 1 2 1140 1136 212 1148 1136 198 ICV_30 $T=303600 214880 1 0 $X=303410 $Y=211920
X1909 1 2 1123 1091 196 1153 1155 219 ICV_30 $T=305900 187680 0 0 $X=305710 $Y=187440
X1910 1 2 1154 268 216 1164 268 198 ICV_30 $T=314640 182240 0 0 $X=314450 $Y=182000
X1911 1 2 1159 1138 155 1162 1138 152 ICV_30 $T=314640 231200 0 0 $X=314450 $Y=230960
X1912 1 2 1168 1172 212 1167 1172 211 ICV_30 $T=324300 204000 0 0 $X=324110 $Y=203760
X1913 1 2 1181 1184 252 1178 1184 232 ICV_30 $T=332580 209440 0 0 $X=332390 $Y=209200
X1914 1 2 1188 1155 196 1208 1201 185 ICV_30 $T=342700 193120 0 0 $X=342510 $Y=192880
X1915 1 2 1200 1201 195 1209 1193 196 ICV_30 $T=345460 209440 1 0 $X=345270 $Y=206480
X1916 1 2 1205 292 196 310 311 219 ICV_30 $T=348220 182240 1 0 $X=348030 $Y=179280
X1917 1 2 1224 1193 198 1230 1193 211 ICV_30 $T=356960 187680 1 0 $X=356770 $Y=184720
X1918 1 2 316 313 238 1221 313 255 ICV_30 $T=357420 242080 0 0 $X=357230 $Y=241840
X1919 1 2 1244 1239 254 1256 1239 261 ICV_30 $T=370760 209440 0 0 $X=370570 $Y=209200
X1920 1 2 1272 1268 219 1276 1255 198 ICV_30 $T=379960 193120 0 0 $X=379770 $Y=192880
X1921 1 2 1303 351 198 1294 351 185 ICV_30 $T=399740 187680 1 0 $X=399550 $Y=184720
X1922 1 2 1346 1347 263 1355 1351 261 ICV_30 $T=420900 204000 1 0 $X=420710 $Y=201040
X1923 1 2 1356 1366 249 366 1366 238 ICV_30 $T=426880 242080 0 0 $X=426690 $Y=241840
X1924 1 2 1365 1368 254 1367 1368 232 ICV_30 $T=427800 214880 0 0 $X=427610 $Y=214640
X1925 1 2 1387 1389 261 1390 1389 232 ICV_30 $T=437920 198560 0 0 $X=437730 $Y=198320
X1926 1 2 1394 370 329 1392 370 249 ICV_30 $T=441140 236640 1 0 $X=440950 $Y=233680
X1927 1 2 1413 1389 263 1417 1337 261 ICV_30 $T=454940 204000 0 0 $X=454750 $Y=203760
X1928 1 2 1425 1422 251 1432 1422 249 ICV_30 $T=459540 225760 0 0 $X=459350 $Y=225520
X1929 1 2 1427 1347 261 1431 1347 232 ICV_30 $T=460460 193120 1 0 $X=460270 $Y=190160
X1930 1 2 1434 382 194 1429 1347 252 ICV_30 $T=462300 182240 0 0 $X=462110 $Y=182000
X1931 1 2 1478 1477 249 1479 1477 271 ICV_30 $T=483920 231200 0 0 $X=483730 $Y=230960
X1932 1 2 1455 1438 329 1485 1491 285 ICV_30 $T=485760 209440 1 0 $X=485570 $Y=206480
X1933 1 2 431 432 413 433 432 412 ICV_30 $T=527160 187680 1 0 $X=526970 $Y=184720
X1934 1 2 1559 1530 415 1550 1530 427 ICV_30 $T=528080 225760 0 0 $X=527890 $Y=225520
X1935 1 2 1573 1546 427 1554 1546 429 ICV_30 $T=539120 209440 0 0 $X=538930 $Y=209200
X1936 1 2 1564 1568 415 1589 1568 429 ICV_30 $T=539120 225760 0 0 $X=538930 $Y=225520
X1937 1 2 1579 1581 251 1593 1581 271 ICV_30 $T=540040 187680 0 0 $X=539850 $Y=187440
X1938 1 2 1585 1568 414 1587 1568 412 ICV_30 $T=541420 236640 1 0 $X=541230 $Y=233680
X1939 1 2 1597 1580 429 1599 1605 238 ICV_30 $T=547400 209440 0 0 $X=547210 $Y=209200
X1940 1 2 1630 1636 251 1639 1636 249 ICV_30 $T=567180 214880 0 0 $X=566990 $Y=214640
X1941 1 2 1628 1612 412 1632 1612 429 ICV_30 $T=567180 236640 0 0 $X=566990 $Y=236400
X1942 1 2 1663 1649 271 1662 1652 329 ICV_30 $T=584660 204000 1 0 $X=584470 $Y=201040
X1943 1 2 1732 1736 255 1728 1736 330 ICV_30 $T=623300 198560 0 0 $X=623110 $Y=198320
X1944 1 2 1758 1759 329 1766 1745 329 ICV_30 $T=632500 220320 0 0 $X=632310 $Y=220080
X1945 1 2 1752 493 238 1749 493 329 ICV_30 $T=637560 198560 1 0 $X=637370 $Y=195600
X1946 1 2 1772 1745 255 1790 1739 271 ICV_30 $T=649060 225760 1 0 $X=648870 $Y=222800
X1947 1 2 1824 1826 429 1835 1826 427 ICV_30 $T=667000 198560 0 0 $X=666810 $Y=198320
X1948 1 2 1855 1856 429 1863 1856 424 ICV_30 $T=680340 236640 0 0 $X=680150 $Y=236400
X1949 1 2 1857 1831 414 1862 1831 413 ICV_30 $T=681720 187680 0 0 $X=681530 $Y=187440
X1950 1 2 1872 1844 429 1859 1856 415 ICV_30 $T=690000 225760 0 0 $X=689810 $Y=225520
X1951 1 2 1874 506 413 1890 506 415 ICV_30 $T=693680 187680 1 0 $X=693490 $Y=184720
X1952 1 2 1884 1885 429 1892 1885 413 ICV_30 $T=694600 193120 1 0 $X=694410 $Y=190160
X1953 1 2 1883 1886 414 1881 1886 429 ICV_30 $T=695060 214880 1 0 $X=694870 $Y=211920
X1954 1 2 1880 1856 412 1873 1856 427 ICV_30 $T=697820 236640 0 0 $X=697630 $Y=236400
X1955 1 2 1900 1901 429 1907 1885 424 ICV_30 $T=703800 193120 1 0 $X=703610 $Y=190160
X1956 1 2 1903 1865 430 1916 1865 415 ICV_30 $T=707480 204000 0 0 $X=707290 $Y=203760
X1957 1 2 1912 1885 414 1924 1885 427 ICV_30 $T=709780 187680 0 0 $X=709590 $Y=187440
X1958 1 2 1941 1901 427 1950 1954 427 ICV_30 $T=721740 198560 1 0 $X=721550 $Y=195600
X1959 1 2 1942 510 412 521 517 427 ICV_30 $T=721740 236640 1 0 $X=721550 $Y=233680
X1960 1 2 516 517 415 520 517 412 ICV_30 $T=721740 242080 1 0 $X=721550 $Y=239120
X1961 1 2 1939 518 412 1953 518 415 ICV_30 $T=722200 182240 0 0 $X=722010 $Y=182000
X1962 1 2 23 26 2 606 1 sky130_fd_sc_hd__and2_1 $T=20700 187680 0 0 $X=20510 $Y=187440
X1963 1 2 37 26 2 605 1 sky130_fd_sc_hd__and2_1 $T=24380 209440 1 0 $X=24190 $Y=206480
X1964 1 2 54 26 2 630 1 sky130_fd_sc_hd__and2_1 $T=40020 209440 0 0 $X=39830 $Y=209200
X1965 1 2 59 26 2 646 1 sky130_fd_sc_hd__and2_1 $T=48300 193120 1 0 $X=48110 $Y=190160
X1966 1 2 67 26 2 679 1 sky130_fd_sc_hd__and2_1 $T=62100 193120 0 0 $X=61910 $Y=192880
X1967 1 2 72 43 2 686 1 sky130_fd_sc_hd__and2_1 $T=66700 242080 0 0 $X=66510 $Y=241840
X1968 1 2 83 43 2 725 1 sky130_fd_sc_hd__and2_1 $T=87860 242080 1 0 $X=87670 $Y=239120
X1969 1 2 84 26 2 708 1 sky130_fd_sc_hd__and2_1 $T=90160 187680 0 0 $X=89970 $Y=187440
X1970 1 2 91 26 2 727 1 sky130_fd_sc_hd__and2_1 $T=98900 204000 0 0 $X=98710 $Y=203760
X1971 1 2 92 26 2 758 1 sky130_fd_sc_hd__and2_1 $T=99820 187680 0 0 $X=99630 $Y=187440
X1972 1 2 101 26 2 775 1 sky130_fd_sc_hd__and2_1 $T=114080 182240 0 0 $X=113890 $Y=182000
X1973 1 2 102 43 2 785 1 sky130_fd_sc_hd__and2_1 $T=114540 242080 0 0 $X=114350 $Y=241840
X1974 1 2 106 26 2 783 1 sky130_fd_sc_hd__and2_1 $T=122360 209440 0 0 $X=122170 $Y=209200
X1975 1 2 107 43 2 796 1 sky130_fd_sc_hd__and2_1 $T=123280 242080 1 0 $X=123090 $Y=239120
X1976 1 2 111 26 2 802 1 sky130_fd_sc_hd__and2_1 $T=132020 198560 0 0 $X=131830 $Y=198320
X1977 1 2 114 26 2 816 1 sky130_fd_sc_hd__and2_1 $T=142140 198560 0 0 $X=141950 $Y=198320
X1978 1 2 115 43 2 822 1 sky130_fd_sc_hd__and2_1 $T=143520 242080 0 0 $X=143330 $Y=241840
X1979 1 2 118 26 2 838 1 sky130_fd_sc_hd__and2_1 $T=149500 214880 1 0 $X=149310 $Y=211920
X1980 1 2 121 26 2 852 1 sky130_fd_sc_hd__and2_1 $T=156400 193120 1 0 $X=156210 $Y=190160
X1981 1 2 126 128 2 870 1 sky130_fd_sc_hd__and2_1 $T=164680 242080 1 0 $X=164490 $Y=239120
X1982 1 2 169 26 2 934 1 sky130_fd_sc_hd__and2_1 $T=198260 193120 0 0 $X=198070 $Y=192880
X1983 1 2 175 26 2 944 1 sky130_fd_sc_hd__and2_1 $T=206540 209440 0 0 $X=206350 $Y=209200
X1984 1 2 37 178 2 959 1 sky130_fd_sc_hd__and2_1 $T=210680 204000 0 0 $X=210490 $Y=203760
X1985 1 2 59 178 2 957 1 sky130_fd_sc_hd__and2_1 $T=211600 198560 0 0 $X=211410 $Y=198320
X1986 1 2 23 178 2 960 1 sky130_fd_sc_hd__and2_1 $T=213440 182240 1 0 $X=213250 $Y=179280
X1987 1 2 52 128 2 184 1 sky130_fd_sc_hd__and2_1 $T=214820 242080 0 0 $X=214630 $Y=241840
X1988 1 2 83 128 2 1003 1 sky130_fd_sc_hd__and2_1 $T=230460 236640 0 0 $X=230270 $Y=236400
X1989 1 2 222 178 2 223 1 sky130_fd_sc_hd__and2_1 $T=241960 182240 1 0 $X=241770 $Y=179280
X1990 1 2 84 178 2 1027 1 sky130_fd_sc_hd__and2_1 $T=241960 198560 1 0 $X=241770 $Y=195600
X1991 1 2 77 178 2 1021 1 sky130_fd_sc_hd__and2_1 $T=241960 204000 0 0 $X=241770 $Y=203760
X1992 1 2 72 128 2 1032 1 sky130_fd_sc_hd__and2_1 $T=246100 242080 1 0 $X=245910 $Y=239120
X1993 1 2 107 128 2 1053 1 sky130_fd_sc_hd__and2_1 $T=254380 236640 0 0 $X=254190 $Y=236400
X1994 1 2 54 178 2 1059 1 sky130_fd_sc_hd__and2_1 $T=258520 204000 0 0 $X=258330 $Y=203760
X1995 1 2 67 178 2 1069 1 sky130_fd_sc_hd__and2_1 $T=272780 193120 1 0 $X=272590 $Y=190160
X1996 1 2 102 128 2 1089 1 sky130_fd_sc_hd__and2_1 $T=272780 236640 0 0 $X=272590 $Y=236400
X1997 1 2 71 178 2 1093 1 sky130_fd_sc_hd__and2_1 $T=274160 182240 1 0 $X=273970 $Y=179280
X1998 1 2 106 178 2 1114 1 sky130_fd_sc_hd__and2_1 $T=286580 198560 0 0 $X=286390 $Y=198320
X1999 1 2 121 178 2 1137 1 sky130_fd_sc_hd__and2_1 $T=297160 187680 0 0 $X=296970 $Y=187440
X2000 1 2 101 178 2 1128 1 sky130_fd_sc_hd__and2_1 $T=300840 182240 1 0 $X=300650 $Y=179280
X2001 1 2 111 178 2 1152 1 sky130_fd_sc_hd__and2_1 $T=310500 198560 0 0 $X=310310 $Y=198320
X2002 1 2 295 178 2 1191 1 sky130_fd_sc_hd__and2_1 $T=335800 187680 0 0 $X=335610 $Y=187440
X2003 1 2 301 302 2 1206 1 sky130_fd_sc_hd__and2_1 $T=342700 225760 0 0 $X=342510 $Y=225520
X2004 1 2 301 308 2 1213 1 sky130_fd_sc_hd__and2_1 $T=350060 231200 0 0 $X=349870 $Y=230960
X2005 1 2 307 302 2 1218 1 sky130_fd_sc_hd__and2_1 $T=350520 220320 0 0 $X=350330 $Y=220080
X2006 1 2 118 178 2 1242 1 sky130_fd_sc_hd__and2_1 $T=370760 198560 0 0 $X=370570 $Y=198320
X2007 1 2 334 308 2 1270 1 sky130_fd_sc_hd__and2_1 $T=380880 225760 1 0 $X=380690 $Y=222800
X2008 1 2 340 308 2 1285 1 sky130_fd_sc_hd__and2_1 $T=387320 231200 0 0 $X=387130 $Y=230960
X2009 1 2 346 302 2 1305 1 sky130_fd_sc_hd__and2_1 $T=396060 225760 0 0 $X=395870 $Y=225520
X2010 1 2 353 302 2 1304 1 sky130_fd_sc_hd__and2_1 $T=398820 209440 1 0 $X=398630 $Y=206480
X2011 1 2 356 302 2 1331 1 sky130_fd_sc_hd__and2_1 $T=409400 187680 0 0 $X=409210 $Y=187440
X2012 1 2 356 308 2 1330 1 sky130_fd_sc_hd__and2_1 $T=413080 225760 1 0 $X=412890 $Y=222800
X2013 1 2 363 302 2 1352 1 sky130_fd_sc_hd__and2_1 $T=421360 209440 1 0 $X=421170 $Y=206480
X2014 1 2 363 308 2 1360 1 sky130_fd_sc_hd__and2_1 $T=424120 231200 0 0 $X=423930 $Y=230960
X2015 1 2 365 302 2 1372 1 sky130_fd_sc_hd__and2_1 $T=431480 225760 1 0 $X=431290 $Y=222800
X2016 1 2 369 308 2 1383 1 sky130_fd_sc_hd__and2_1 $T=438840 225760 0 0 $X=438650 $Y=225520
X2017 1 2 368 308 2 1405 1 sky130_fd_sc_hd__and2_1 $T=450800 193120 0 0 $X=450610 $Y=192880
X2018 1 2 378 308 2 1414 1 sky130_fd_sc_hd__and2_1 $T=454940 242080 0 0 $X=454750 $Y=241840
X2019 1 2 380 308 2 1420 1 sky130_fd_sc_hd__and2_1 $T=455860 214880 0 0 $X=455670 $Y=214640
X2020 1 2 381 308 2 1430 1 sky130_fd_sc_hd__and2_1 $T=460000 182240 0 0 $X=459810 $Y=182000
X2021 1 2 385 308 2 1426 1 sky130_fd_sc_hd__and2_1 $T=465060 242080 0 0 $X=464870 $Y=241840
X2022 1 2 390 308 2 1452 1 sky130_fd_sc_hd__and2_1 $T=475180 225760 0 0 $X=474990 $Y=225520
X2023 1 2 394 302 2 1470 1 sky130_fd_sc_hd__and2_1 $T=479320 209440 0 0 $X=479130 $Y=209200
X2024 1 2 397 308 2 1480 1 sky130_fd_sc_hd__and2_1 $T=490360 182240 0 0 $X=490170 $Y=182000
X2025 1 2 340 398 2 1493 1 sky130_fd_sc_hd__and2_1 $T=491280 236640 1 0 $X=491090 $Y=233680
X2026 1 2 400 308 2 1496 1 sky130_fd_sc_hd__and2_1 $T=494040 198560 1 0 $X=493850 $Y=195600
X2027 1 2 353 398 2 1503 1 sky130_fd_sc_hd__and2_1 $T=497260 220320 1 0 $X=497070 $Y=217360
X2028 1 2 315 398 2 1506 1 sky130_fd_sc_hd__and2_1 $T=501400 242080 1 0 $X=501210 $Y=239120
X2029 1 2 301 398 2 1532 1 sky130_fd_sc_hd__and2_1 $T=513820 214880 1 0 $X=513630 $Y=211920
X2030 1 2 428 308 2 1543 1 sky130_fd_sc_hd__and2_1 $T=522560 187680 1 0 $X=522370 $Y=184720
X2031 1 2 356 398 2 1549 1 sky130_fd_sc_hd__and2_1 $T=522560 231200 1 0 $X=522370 $Y=228240
X2032 1 2 378 398 2 1562 1 sky130_fd_sc_hd__and2_1 $T=529460 242080 1 0 $X=529270 $Y=239120
X2033 1 2 369 398 2 1569 1 sky130_fd_sc_hd__and2_1 $T=532680 225760 1 0 $X=532490 $Y=222800
X2034 1 2 441 308 2 1592 1 sky130_fd_sc_hd__and2_1 $T=549240 182240 1 0 $X=549050 $Y=179280
X2035 1 2 390 398 2 1602 1 sky130_fd_sc_hd__and2_1 $T=549700 236640 1 0 $X=549510 $Y=233680
X2036 1 2 442 308 2 1606 1 sky130_fd_sc_hd__and2_1 $T=553380 204000 1 0 $X=553190 $Y=201040
X2037 1 2 446 308 2 1626 1 sky130_fd_sc_hd__and2_1 $T=563040 193120 0 0 $X=562850 $Y=192880
X2038 1 2 448 308 2 1615 1 sky130_fd_sc_hd__and2_1 $T=563500 209440 0 0 $X=563310 $Y=209200
X2039 1 2 457 308 2 1644 1 sky130_fd_sc_hd__and2_1 $T=574540 242080 0 0 $X=574350 $Y=241840
X2040 1 2 461 308 2 1654 1 sky130_fd_sc_hd__and2_1 $T=577760 225760 1 0 $X=577570 $Y=222800
X2041 1 2 464 308 2 1641 1 sky130_fd_sc_hd__and2_1 $T=582360 209440 0 0 $X=582170 $Y=209200
X2042 1 2 469 308 2 1678 1 sky130_fd_sc_hd__and2_1 $T=592480 225760 0 0 $X=592290 $Y=225520
X2043 1 2 470 308 2 1684 1 sky130_fd_sc_hd__and2_1 $T=592480 231200 0 0 $X=592290 $Y=230960
X2044 1 2 476 308 2 1687 1 sky130_fd_sc_hd__and2_1 $T=602600 198560 1 0 $X=602410 $Y=195600
X2045 1 2 482 308 2 1719 1 sky130_fd_sc_hd__and2_1 $T=616400 214880 1 0 $X=616210 $Y=211920
X2046 1 2 487 308 2 1715 1 sky130_fd_sc_hd__and2_1 $T=622380 204000 1 0 $X=622190 $Y=201040
X2047 1 2 489 308 2 1746 1 sky130_fd_sc_hd__and2_1 $T=627900 242080 0 0 $X=627710 $Y=241840
X2048 1 2 494 308 2 1757 1 sky130_fd_sc_hd__and2_1 $T=632960 209440 1 0 $X=632770 $Y=206480
X2049 1 2 496 308 2 1760 1 sky130_fd_sc_hd__and2_1 $T=636640 193120 0 0 $X=636450 $Y=192880
X2050 1 2 497 308 2 1767 1 sky130_fd_sc_hd__and2_1 $T=637560 187680 1 0 $X=637370 $Y=184720
X2051 1 2 498 308 2 1737 1 sky130_fd_sc_hd__and2_1 $T=637560 231200 1 0 $X=637370 $Y=228240
X2052 1 2 457 398 2 1792 1 sky130_fd_sc_hd__and2_1 $T=648600 225760 0 0 $X=648410 $Y=225520
X2053 1 2 400 398 2 1814 1 sky130_fd_sc_hd__and2_1 $T=661480 204000 1 0 $X=661290 $Y=201040
X2054 1 2 428 398 2 1819 1 sky130_fd_sc_hd__and2_1 $T=662860 187680 1 0 $X=662670 $Y=184720
X2055 1 2 380 398 2 1828 1 sky130_fd_sc_hd__and2_1 $T=672060 225760 0 0 $X=671870 $Y=225520
X2056 1 2 494 398 2 1846 1 sky130_fd_sc_hd__and2_1 $T=676660 198560 0 0 $X=676470 $Y=198320
X2057 1 2 470 398 2 1849 1 sky130_fd_sc_hd__and2_1 $T=683560 220320 0 0 $X=683370 $Y=220080
X2058 1 2 496 398 2 1869 1 sky130_fd_sc_hd__and2_1 $T=690000 187680 0 0 $X=689810 $Y=187440
X2059 1 2 464 398 2 1860 1 sky130_fd_sc_hd__and2_1 $T=693680 209440 1 0 $X=693490 $Y=206480
X2060 1 2 461 398 2 1915 1 sky130_fd_sc_hd__and2_1 $T=708860 220320 0 0 $X=708670 $Y=220080
X2061 1 2 498 398 2 1913 1 sky130_fd_sc_hd__and2_1 $T=710700 231200 1 0 $X=710510 $Y=228240
X2062 1 2 448 398 2 1921 1 sky130_fd_sc_hd__and2_1 $T=712080 209440 1 0 $X=711890 $Y=206480
X2063 1 2 482 398 2 1929 1 sky130_fd_sc_hd__and2_1 $T=715760 204000 0 0 $X=715570 $Y=203760
X2064 1 2 497 398 2 1927 1 sky130_fd_sc_hd__and2_1 $T=717600 187680 1 0 $X=717410 $Y=184720
X2065 1 2 ICV_31 $T=45540 236640 1 0 $X=45350 $Y=233680
X2066 1 2 ICV_31 $T=59340 193120 0 0 $X=59150 $Y=192880
X2067 1 2 ICV_31 $T=129720 225760 1 0 $X=129530 $Y=222800
X2068 1 2 ICV_31 $T=171580 198560 0 0 $X=171390 $Y=198320
X2069 1 2 ICV_31 $T=185840 209440 1 0 $X=185650 $Y=206480
X2070 1 2 ICV_31 $T=199640 198560 0 0 $X=199450 $Y=198320
X2071 1 2 ICV_31 $T=227700 225760 0 0 $X=227510 $Y=225520
X2072 1 2 ICV_31 $T=270020 220320 1 0 $X=269830 $Y=217360
X2073 1 2 ICV_31 $T=283820 198560 0 0 $X=283630 $Y=198320
X2074 1 2 ICV_31 $T=283820 231200 0 0 $X=283630 $Y=230960
X2075 1 2 ICV_31 $T=298080 187680 1 0 $X=297890 $Y=184720
X2076 1 2 ICV_31 $T=382260 242080 1 0 $X=382070 $Y=239120
X2077 1 2 ICV_31 $T=410320 204000 1 0 $X=410130 $Y=201040
X2078 1 2 ICV_31 $T=410320 220320 1 0 $X=410130 $Y=217360
X2079 1 2 ICV_31 $T=522560 198560 1 0 $X=522370 $Y=195600
X2080 1 2 ICV_31 $T=564420 225760 0 0 $X=564230 $Y=225520
X2081 1 2 ICV_31 $T=564420 236640 0 0 $X=564230 $Y=236400
X2082 1 2 ICV_31 $T=592480 187680 0 0 $X=592290 $Y=187440
X2083 1 2 ICV_31 $T=606740 204000 1 0 $X=606550 $Y=201040
X2084 1 2 ICV_31 $T=606740 209440 1 0 $X=606550 $Y=206480
X2085 1 2 ICV_31 $T=620540 220320 0 0 $X=620350 $Y=220080
X2086 1 2 ICV_31 $T=662860 214880 1 0 $X=662670 $Y=211920
X2087 1 2 ICV_31 $T=690920 220320 1 0 $X=690730 $Y=217360
X2088 1 2 287 4 2 587 1 sky130_fd_sc_hd__dlclkp_1 $T=6900 236640 0 0 $X=6710 $Y=236400
X2089 1 2 266 605 2 589 1 sky130_fd_sc_hd__dlclkp_1 $T=18860 209440 0 0 $X=18670 $Y=209200
X2090 1 2 266 606 2 588 1 sky130_fd_sc_hd__dlclkp_1 $T=20240 193120 1 0 $X=20050 $Y=190160
X2091 1 2 287 51 2 608 1 sky130_fd_sc_hd__dlclkp_1 $T=34040 242080 0 0 $X=33850 $Y=241840
X2092 1 2 266 630 2 627 1 sky130_fd_sc_hd__dlclkp_1 $T=38640 214880 0 0 $X=38450 $Y=214640
X2093 1 2 266 646 2 626 1 sky130_fd_sc_hd__dlclkp_1 $T=42780 198560 0 0 $X=42590 $Y=198320
X2094 1 2 266 63 2 652 1 sky130_fd_sc_hd__dlclkp_1 $T=57500 182240 1 0 $X=57310 $Y=179280
X2095 1 2 287 675 2 653 1 sky130_fd_sc_hd__dlclkp_1 $T=62100 236640 0 0 $X=61910 $Y=236400
X2096 1 2 266 679 2 660 1 sky130_fd_sc_hd__dlclkp_1 $T=64400 193120 0 0 $X=64210 $Y=192880
X2097 1 2 287 686 2 702 1 sky130_fd_sc_hd__dlclkp_1 $T=66700 242080 1 0 $X=66510 $Y=239120
X2098 1 2 266 704 2 676 1 sky130_fd_sc_hd__dlclkp_1 $T=72680 209440 0 0 $X=72490 $Y=209200
X2099 1 2 266 708 2 703 1 sky130_fd_sc_hd__dlclkp_1 $T=75900 187680 0 0 $X=75710 $Y=187440
X2100 1 2 266 78 2 74 1 sky130_fd_sc_hd__dlclkp_1 $T=76820 182240 1 0 $X=76630 $Y=179280
X2101 1 2 287 725 2 86 1 sky130_fd_sc_hd__dlclkp_1 $T=83260 242080 0 0 $X=83070 $Y=241840
X2102 1 2 266 727 2 734 1 sky130_fd_sc_hd__dlclkp_1 $T=85560 204000 1 0 $X=85370 $Y=201040
X2103 1 2 266 758 2 735 1 sky130_fd_sc_hd__dlclkp_1 $T=104420 193120 1 0 $X=104230 $Y=190160
X2104 1 2 266 775 2 784 1 sky130_fd_sc_hd__dlclkp_1 $T=111320 187680 0 0 $X=111130 $Y=187440
X2105 1 2 266 783 2 751 1 sky130_fd_sc_hd__dlclkp_1 $T=113620 214880 1 0 $X=113430 $Y=211920
X2106 1 2 287 785 2 760 1 sky130_fd_sc_hd__dlclkp_1 $T=115460 242080 1 0 $X=115270 $Y=239120
X2107 1 2 266 802 2 764 1 sky130_fd_sc_hd__dlclkp_1 $T=125580 198560 0 0 $X=125390 $Y=198320
X2108 1 2 287 796 2 793 1 sky130_fd_sc_hd__dlclkp_1 $T=125580 242080 1 0 $X=125390 $Y=239120
X2109 1 2 266 816 2 819 1 sky130_fd_sc_hd__dlclkp_1 $T=135700 198560 0 0 $X=135510 $Y=198320
X2110 1 2 287 822 2 836 1 sky130_fd_sc_hd__dlclkp_1 $T=137080 242080 0 0 $X=136890 $Y=241840
X2111 1 2 266 838 2 813 1 sky130_fd_sc_hd__dlclkp_1 $T=143060 214880 1 0 $X=142870 $Y=211920
X2112 1 2 266 852 2 860 1 sky130_fd_sc_hd__dlclkp_1 $T=153180 193120 0 0 $X=152990 $Y=192880
X2113 1 2 266 859 2 866 1 sky130_fd_sc_hd__dlclkp_1 $T=155940 209440 0 0 $X=155750 $Y=209200
X2114 1 2 287 870 2 875 1 sky130_fd_sc_hd__dlclkp_1 $T=164220 242080 0 0 $X=164030 $Y=241840
X2115 1 2 266 173 2 897 1 sky130_fd_sc_hd__dlclkp_1 $T=202400 182240 0 0 $X=202210 $Y=182000
X2116 1 2 266 934 2 905 1 sky130_fd_sc_hd__dlclkp_1 $T=202400 193120 0 0 $X=202210 $Y=192880
X2117 1 2 266 944 2 911 1 sky130_fd_sc_hd__dlclkp_1 $T=202400 209440 1 0 $X=202210 $Y=206480
X2118 1 2 287 948 2 955 1 sky130_fd_sc_hd__dlclkp_1 $T=205160 236640 0 0 $X=204970 $Y=236400
X2119 1 2 266 957 2 963 1 sky130_fd_sc_hd__dlclkp_1 $T=208380 198560 1 0 $X=208190 $Y=195600
X2120 1 2 266 959 2 967 1 sky130_fd_sc_hd__dlclkp_1 $T=208840 209440 1 0 $X=208650 $Y=206480
X2121 1 2 266 960 2 962 1 sky130_fd_sc_hd__dlclkp_1 $T=209760 187680 0 0 $X=209570 $Y=187440
X2122 1 2 287 1003 2 1002 1 sky130_fd_sc_hd__dlclkp_1 $T=230460 242080 0 0 $X=230270 $Y=241840
X2123 1 2 266 1021 2 1022 1 sky130_fd_sc_hd__dlclkp_1 $T=237360 209440 1 0 $X=237170 $Y=206480
X2124 1 2 266 1027 2 1028 1 sky130_fd_sc_hd__dlclkp_1 $T=241960 193120 0 0 $X=241770 $Y=192880
X2125 1 2 287 1032 2 1048 1 sky130_fd_sc_hd__dlclkp_1 $T=250700 242080 0 0 $X=250510 $Y=241840
X2126 1 2 266 1059 2 1062 1 sky130_fd_sc_hd__dlclkp_1 $T=258520 198560 0 0 $X=258330 $Y=198320
X2127 1 2 287 1053 2 240 1 sky130_fd_sc_hd__dlclkp_1 $T=258520 242080 0 0 $X=258330 $Y=241840
X2128 1 2 266 1069 2 1066 1 sky130_fd_sc_hd__dlclkp_1 $T=264960 193120 1 0 $X=264770 $Y=190160
X2129 1 2 266 1090 2 1096 1 sky130_fd_sc_hd__dlclkp_1 $T=273240 204000 1 0 $X=273050 $Y=201040
X2130 1 2 287 1089 2 1092 1 sky130_fd_sc_hd__dlclkp_1 $T=273700 242080 1 0 $X=273510 $Y=239120
X2131 1 2 266 1093 2 1108 1 sky130_fd_sc_hd__dlclkp_1 $T=278760 182240 0 0 $X=278570 $Y=182000
X2132 1 2 266 1114 2 1121 1 sky130_fd_sc_hd__dlclkp_1 $T=290720 204000 0 0 $X=290530 $Y=203760
X2133 1 2 266 1128 2 262 1 sky130_fd_sc_hd__dlclkp_1 $T=293940 182240 1 0 $X=293750 $Y=179280
X2134 1 2 287 1131 2 1116 1 sky130_fd_sc_hd__dlclkp_1 $T=296700 242080 0 0 $X=296510 $Y=241840
X2135 1 2 266 1137 2 1141 1 sky130_fd_sc_hd__dlclkp_1 $T=299460 187680 0 0 $X=299270 $Y=187440
X2136 1 2 266 1152 2 1156 1 sky130_fd_sc_hd__dlclkp_1 $T=308200 204000 1 0 $X=308010 $Y=201040
X2137 1 2 266 281 2 283 1 sky130_fd_sc_hd__dlclkp_1 $T=322000 182240 1 0 $X=321810 $Y=179280
X2138 1 2 266 1180 2 1183 1 sky130_fd_sc_hd__dlclkp_1 $T=331660 204000 1 0 $X=331470 $Y=201040
X2139 1 2 266 1191 2 1197 1 sky130_fd_sc_hd__dlclkp_1 $T=342700 187680 0 0 $X=342510 $Y=187440
X2140 1 2 338 1206 2 1173 1 sky130_fd_sc_hd__dlclkp_1 $T=345000 225760 0 0 $X=344810 $Y=225520
X2141 1 2 338 1213 2 1202 1 sky130_fd_sc_hd__dlclkp_1 $T=347300 231200 1 0 $X=347110 $Y=228240
X2142 1 2 338 1218 2 1203 1 sky130_fd_sc_hd__dlclkp_1 $T=348220 225760 1 0 $X=348030 $Y=222800
X2143 1 2 338 1232 2 1234 1 sky130_fd_sc_hd__dlclkp_1 $T=357420 209440 0 0 $X=357230 $Y=209200
X2144 1 2 266 323 2 1237 1 sky130_fd_sc_hd__dlclkp_1 $T=362940 187680 0 0 $X=362750 $Y=187440
X2145 1 2 266 1242 2 1252 1 sky130_fd_sc_hd__dlclkp_1 $T=363860 204000 1 0 $X=363670 $Y=201040
X2146 1 2 338 1260 2 1262 1 sky130_fd_sc_hd__dlclkp_1 $T=374440 225760 1 0 $X=374250 $Y=222800
X2147 1 2 338 1270 2 1249 1 sky130_fd_sc_hd__dlclkp_1 $T=377200 231200 1 0 $X=377010 $Y=228240
X2148 1 2 338 1285 2 331 1 sky130_fd_sc_hd__dlclkp_1 $T=391000 236640 0 0 $X=390810 $Y=236400
X2149 1 2 338 1304 2 1308 1 sky130_fd_sc_hd__dlclkp_1 $T=396060 204000 1 0 $X=395870 $Y=201040
X2150 1 2 338 1305 2 1306 1 sky130_fd_sc_hd__dlclkp_1 $T=398360 225760 1 0 $X=398170 $Y=222800
X2151 1 2 338 1330 2 1301 1 sky130_fd_sc_hd__dlclkp_1 $T=408020 225760 0 0 $X=407830 $Y=225520
X2152 1 2 338 1331 2 1339 1 sky130_fd_sc_hd__dlclkp_1 $T=411700 187680 0 0 $X=411510 $Y=187440
X2153 1 2 338 359 2 354 1 sky130_fd_sc_hd__dlclkp_1 $T=412620 242080 0 0 $X=412430 $Y=241840
X2154 1 2 338 1332 2 1342 1 sky130_fd_sc_hd__dlclkp_1 $T=415380 214880 0 0 $X=415190 $Y=214640
X2155 1 2 338 1352 2 1369 1 sky130_fd_sc_hd__dlclkp_1 $T=423660 209440 1 0 $X=423470 $Y=206480
X2156 1 2 338 1360 2 361 1 sky130_fd_sc_hd__dlclkp_1 $T=426880 225760 0 0 $X=426690 $Y=225520
X2157 1 2 338 1372 2 1391 1 sky130_fd_sc_hd__dlclkp_1 $T=433780 225760 1 0 $X=433590 $Y=222800
X2158 1 2 338 1383 2 1375 1 sky130_fd_sc_hd__dlclkp_1 $T=434240 231200 1 0 $X=434050 $Y=228240
X2159 1 2 338 1379 2 1395 1 sky130_fd_sc_hd__dlclkp_1 $T=436540 187680 0 0 $X=436350 $Y=187440
X2160 1 2 338 1405 2 1415 1 sky130_fd_sc_hd__dlclkp_1 $T=448040 198560 0 0 $X=447850 $Y=198320
X2161 1 2 338 1414 2 1412 1 sky130_fd_sc_hd__dlclkp_1 $T=450340 242080 1 0 $X=450150 $Y=239120
X2162 1 2 338 1426 2 384 1 sky130_fd_sc_hd__dlclkp_1 $T=458620 242080 0 0 $X=458430 $Y=241840
X2163 1 2 338 1420 2 1428 1 sky130_fd_sc_hd__dlclkp_1 $T=459080 220320 1 0 $X=458890 $Y=217360
X2164 1 2 338 1430 2 1440 1 sky130_fd_sc_hd__dlclkp_1 $T=462300 187680 1 0 $X=462110 $Y=184720
X2165 1 2 338 1452 2 1456 1 sky130_fd_sc_hd__dlclkp_1 $T=470120 231200 1 0 $X=469930 $Y=228240
X2166 1 2 338 1470 2 1476 1 sky130_fd_sc_hd__dlclkp_1 $T=479320 209440 1 0 $X=479130 $Y=206480
X2167 1 2 338 1480 2 1481 1 sky130_fd_sc_hd__dlclkp_1 $T=483920 182240 0 0 $X=483730 $Y=182000
X2168 1 2 338 1493 2 1504 1 sky130_fd_sc_hd__dlclkp_1 $T=491280 236640 0 0 $X=491090 $Y=236400
X2169 1 2 338 1496 2 1474 1 sky130_fd_sc_hd__dlclkp_1 $T=492200 198560 0 0 $X=492010 $Y=198320
X2170 1 2 338 1503 2 1508 1 sky130_fd_sc_hd__dlclkp_1 $T=494960 220320 0 0 $X=494770 $Y=220080
X2171 1 2 338 1506 2 408 1 sky130_fd_sc_hd__dlclkp_1 $T=498180 242080 0 0 $X=497990 $Y=241840
X2172 1 2 338 1532 2 1535 1 sky130_fd_sc_hd__dlclkp_1 $T=513360 209440 1 0 $X=513170 $Y=206480
X2173 1 2 338 1543 2 1526 1 sky130_fd_sc_hd__dlclkp_1 $T=518420 193120 1 0 $X=518230 $Y=190160
X2174 1 2 338 1549 2 1551 1 sky130_fd_sc_hd__dlclkp_1 $T=521640 225760 0 0 $X=521450 $Y=225520
X2175 1 2 338 1562 2 436 1 sky130_fd_sc_hd__dlclkp_1 $T=529000 242080 0 0 $X=528810 $Y=241840
X2176 1 2 338 1569 2 1576 1 sky130_fd_sc_hd__dlclkp_1 $T=532220 220320 0 0 $X=532030 $Y=220080
X2177 1 2 338 1572 2 1563 1 sky130_fd_sc_hd__dlclkp_1 $T=533600 182240 1 0 $X=533410 $Y=179280
X2178 1 2 338 1592 2 1598 1 sky130_fd_sc_hd__dlclkp_1 $T=542800 182240 1 0 $X=542610 $Y=179280
X2179 1 2 338 1602 2 1594 1 sky130_fd_sc_hd__dlclkp_1 $T=546480 231200 1 0 $X=546290 $Y=228240
X2180 1 2 338 1606 2 1582 1 sky130_fd_sc_hd__dlclkp_1 $T=550160 198560 0 0 $X=549970 $Y=198320
X2181 1 2 338 1615 2 1617 1 sky130_fd_sc_hd__dlclkp_1 $T=555220 214880 1 0 $X=555030 $Y=211920
X2182 1 2 338 1626 2 1637 1 sky130_fd_sc_hd__dlclkp_1 $T=562120 198560 1 0 $X=561930 $Y=195600
X2183 1 2 338 1641 2 1643 1 sky130_fd_sc_hd__dlclkp_1 $T=568560 209440 0 0 $X=568370 $Y=209200
X2184 1 2 338 1644 2 453 1 sky130_fd_sc_hd__dlclkp_1 $T=571780 242080 1 0 $X=571590 $Y=239120
X2185 1 2 338 459 2 463 1 sky130_fd_sc_hd__dlclkp_1 $T=574540 182240 1 0 $X=574350 $Y=179280
X2186 1 2 338 1654 2 1642 1 sky130_fd_sc_hd__dlclkp_1 $T=581440 225760 1 0 $X=581250 $Y=222800
X2187 1 2 338 1659 2 467 1 sky130_fd_sc_hd__dlclkp_1 $T=586040 242080 0 0 $X=585850 $Y=241840
X2188 1 2 338 1678 2 1685 1 sky130_fd_sc_hd__dlclkp_1 $T=590180 225760 1 0 $X=589990 $Y=222800
X2189 1 2 338 1687 2 1686 1 sky130_fd_sc_hd__dlclkp_1 $T=596160 198560 1 0 $X=595970 $Y=195600
X2190 1 2 338 1684 2 1688 1 sky130_fd_sc_hd__dlclkp_1 $T=596160 231200 0 0 $X=595970 $Y=230960
X2191 1 2 338 1715 2 1714 1 sky130_fd_sc_hd__dlclkp_1 $T=612720 198560 0 0 $X=612530 $Y=198320
X2192 1 2 338 1719 2 1727 1 sky130_fd_sc_hd__dlclkp_1 $T=615020 214880 0 0 $X=614830 $Y=214640
X2193 1 2 338 1737 2 1743 1 sky130_fd_sc_hd__dlclkp_1 $T=621460 231200 1 0 $X=621270 $Y=228240
X2194 1 2 338 1746 2 495 1 sky130_fd_sc_hd__dlclkp_1 $T=627900 242080 1 0 $X=627710 $Y=239120
X2195 1 2 338 1757 2 1765 1 sky130_fd_sc_hd__dlclkp_1 $T=631120 209440 0 0 $X=630930 $Y=209200
X2196 1 2 338 1760 2 1768 1 sky130_fd_sc_hd__dlclkp_1 $T=632960 198560 0 0 $X=632770 $Y=198320
X2197 1 2 338 1767 2 1770 1 sky130_fd_sc_hd__dlclkp_1 $T=636180 182240 0 0 $X=635990 $Y=182000
X2198 1 2 338 1793 2 1795 1 sky130_fd_sc_hd__dlclkp_1 $T=651360 231200 1 0 $X=651170 $Y=228240
X2199 1 2 338 1792 2 1802 1 sky130_fd_sc_hd__dlclkp_1 $T=651820 225760 0 0 $X=651630 $Y=225520
X2200 1 2 338 1814 2 1815 1 sky130_fd_sc_hd__dlclkp_1 $T=660560 198560 0 0 $X=660370 $Y=198320
X2201 1 2 338 1819 2 1816 1 sky130_fd_sc_hd__dlclkp_1 $T=664240 187680 0 0 $X=664050 $Y=187440
X2202 1 2 338 1828 2 1839 1 sky130_fd_sc_hd__dlclkp_1 $T=667920 231200 1 0 $X=667730 $Y=228240
X2203 1 2 338 1829 2 505 1 sky130_fd_sc_hd__dlclkp_1 $T=670680 182240 0 0 $X=670490 $Y=182000
X2204 1 2 338 1849 2 1861 1 sky130_fd_sc_hd__dlclkp_1 $T=677580 225760 1 0 $X=677390 $Y=222800
X2205 1 2 338 1860 2 1867 1 sky130_fd_sc_hd__dlclkp_1 $T=680800 209440 0 0 $X=680610 $Y=209200
X2206 1 2 338 1864 2 508 1 sky130_fd_sc_hd__dlclkp_1 $T=683100 242080 1 0 $X=682910 $Y=239120
X2207 1 2 338 1869 2 1876 1 sky130_fd_sc_hd__dlclkp_1 $T=686780 193120 1 0 $X=686590 $Y=190160
X2208 1 2 338 1846 2 1866 1 sky130_fd_sc_hd__dlclkp_1 $T=693220 198560 0 0 $X=693030 $Y=198320
X2209 1 2 338 1913 2 1923 1 sky130_fd_sc_hd__dlclkp_1 $T=707940 231200 0 0 $X=707750 $Y=230960
X2210 1 2 338 512 2 514 1 sky130_fd_sc_hd__dlclkp_1 $T=708400 242080 0 0 $X=708210 $Y=241840
X2211 1 2 338 1915 2 1917 1 sky130_fd_sc_hd__dlclkp_1 $T=711160 220320 0 0 $X=710970 $Y=220080
X2212 1 2 338 1927 2 1933 1 sky130_fd_sc_hd__dlclkp_1 $T=713460 182240 0 0 $X=713270 $Y=182000
X2213 1 2 338 1921 2 1935 1 sky130_fd_sc_hd__dlclkp_1 $T=714380 209440 1 0 $X=714190 $Y=206480
X2214 1 2 338 1929 2 1934 1 sky130_fd_sc_hd__dlclkp_1 $T=714840 204000 1 0 $X=714650 $Y=201040
X2215 1 2 ICV_32 $T=44160 187680 1 0 $X=43970 $Y=184720
X2216 1 2 ICV_32 $T=57960 220320 0 0 $X=57770 $Y=220080
X2217 1 2 ICV_32 $T=86020 225760 0 0 $X=85830 $Y=225520
X2218 1 2 ICV_32 $T=86020 231200 0 0 $X=85830 $Y=230960
X2219 1 2 ICV_32 $T=142140 182240 0 0 $X=141950 $Y=182000
X2220 1 2 ICV_32 $T=156400 204000 1 0 $X=156210 $Y=201040
X2221 1 2 ICV_32 $T=226320 209440 0 0 $X=226130 $Y=209200
X2222 1 2 ICV_32 $T=240580 214880 1 0 $X=240390 $Y=211920
X2223 1 2 ICV_32 $T=310500 214880 0 0 $X=310310 $Y=214640
X2224 1 2 ICV_32 $T=324760 242080 1 0 $X=324570 $Y=239120
X2225 1 2 ICV_32 $T=338560 193120 0 0 $X=338370 $Y=192880
X2226 1 2 ICV_32 $T=380880 236640 1 0 $X=380690 $Y=233680
X2227 1 2 ICV_32 $T=577300 193120 1 0 $X=577110 $Y=190160
X2228 1 2 ICV_32 $T=619160 182240 0 0 $X=618970 $Y=182000
X2229 1 2 ICV_32 $T=619160 187680 0 0 $X=618970 $Y=187440
X2230 1 2 ICV_32 $T=619160 198560 0 0 $X=618970 $Y=198320
X2231 1 2 ICV_32 $T=689540 187680 1 0 $X=689350 $Y=184720
X2232 1 2 ICV_32 $T=689540 242080 1 0 $X=689350 $Y=239120
X2233 1 2 ICV_32 $T=717600 198560 1 0 $X=717410 $Y=195600
X2234 1 2 589 13 596 ICV_35 $T=10580 209440 0 0 $X=10390 $Y=209200
X2235 1 2 589 11 597 ICV_35 $T=10580 214880 1 0 $X=10390 $Y=211920
X2236 1 2 589 36 622 ICV_35 $T=23460 214880 0 0 $X=23270 $Y=214640
X2237 1 2 589 35 623 ICV_35 $T=24380 214880 1 0 $X=24190 $Y=211920
X2238 1 2 626 33 635 ICV_35 $T=34040 198560 0 0 $X=33850 $Y=198320
X2239 1 2 626 13 665 ICV_35 $T=48300 198560 1 0 $X=48110 $Y=195600
X2240 1 2 660 13 680 ICV_35 $T=56580 198560 1 0 $X=56390 $Y=195600
X2241 1 2 653 20 695 ICV_35 $T=62100 225760 0 0 $X=61910 $Y=225520
X2242 1 2 703 13 728 ICV_35 $T=80500 198560 1 0 $X=80310 $Y=195600
X2243 1 2 703 35 732 ICV_35 $T=81420 193120 0 0 $X=81230 $Y=192880
X2244 1 2 734 13 739 ICV_35 $T=90160 214880 1 0 $X=89970 $Y=211920
X2245 1 2 734 12 740 ICV_35 $T=90160 220320 0 0 $X=89970 $Y=220080
X2246 1 2 86 25 741 ICV_35 $T=90160 236640 0 0 $X=89970 $Y=236400
X2247 1 2 86 6 742 ICV_35 $T=90160 242080 1 0 $X=89970 $Y=239120
X2248 1 2 751 11 759 ICV_35 $T=98440 220320 0 0 $X=98250 $Y=220080
X2249 1 2 751 36 771 ICV_35 $T=104420 214880 1 0 $X=104230 $Y=211920
X2250 1 2 764 13 789 ICV_35 $T=112700 209440 1 0 $X=112510 $Y=206480
X2251 1 2 760 21 791 ICV_35 $T=115920 236640 1 0 $X=115730 $Y=233680
X2252 1 2 116 33 848 ICV_35 $T=144900 187680 1 0 $X=144710 $Y=184720
X2253 1 2 116 11 854 ICV_35 $T=148120 193120 1 0 $X=147930 $Y=190160
X2254 1 2 813 34 857 ICV_35 $T=148580 225760 1 0 $X=148390 $Y=222800
X2255 1 2 866 11 874 ICV_35 $T=160540 209440 1 0 $X=160350 $Y=206480
X2256 1 2 866 36 876 ICV_35 $T=161000 214880 0 0 $X=160810 $Y=214640
X2257 1 2 127 39 890 ICV_35 $T=168360 231200 1 0 $X=168170 $Y=228240
X2258 1 2 875 147 915 ICV_35 $T=179860 242080 1 0 $X=179670 $Y=239120
X2259 1 2 911 12 938 ICV_35 $T=193660 214880 0 0 $X=193470 $Y=214640
X2260 1 2 955 130 997 ICV_35 $T=220340 236640 0 0 $X=220150 $Y=236400
X2261 1 2 1002 138 1026 ICV_35 $T=232760 236640 0 0 $X=232570 $Y=236400
X2262 1 2 127 215 225 ICV_35 $T=237820 187680 0 0 $X=237630 $Y=187440
X2263 1 2 1028 183 235 ICV_35 $T=252080 193120 1 0 $X=251890 $Y=190160
X2264 1 2 1048 148 1056 ICV_35 $T=252080 231200 1 0 $X=251890 $Y=228240
X2265 1 2 1062 188 1074 ICV_35 $T=261280 204000 1 0 $X=261090 $Y=201040
X2266 1 2 1066 205 1084 ICV_35 $T=264960 198560 0 0 $X=264770 $Y=198320
X2267 1 2 1092 146 1107 ICV_35 $T=275540 231200 0 0 $X=275350 $Y=230960
X2268 1 2 1096 181 1104 ICV_35 $T=276920 214880 1 0 $X=276730 $Y=211920
X2269 1 2 127 261 906 ICV_35 $T=295780 220320 0 0 $X=295590 $Y=220080
X2270 1 2 1116 149 1160 ICV_35 $T=305900 242080 1 0 $X=305710 $Y=239120
X2271 1 2 1156 205 1176 ICV_35 $T=319700 209440 1 0 $X=319510 $Y=206480
X2272 1 2 1183 205 1195 ICV_35 $T=332580 204000 0 0 $X=332390 $Y=203760
X2273 1 2 1183 188 1200 ICV_35 $T=333500 198560 0 0 $X=333310 $Y=198320
X2274 1 2 1197 188 1207 ICV_35 $T=342700 182240 0 0 $X=342510 $Y=182000
X2275 1 2 1237 181 1276 ICV_35 $T=376280 193120 1 0 $X=376090 $Y=190160
X2276 1 2 339 199 1302 ICV_35 $T=389160 187680 1 0 $X=388970 $Y=184720
X2277 1 2 354 286 1317 ICV_35 $T=398820 242080 0 0 $X=398630 $Y=241840
X2278 1 2 339 183 1323 ICV_35 $T=401120 182240 0 0 $X=400930 $Y=182000
X2279 1 2 1339 280 1349 ICV_35 $T=417220 193120 1 0 $X=417030 $Y=190160
X2280 1 2 361 286 1364 ICV_35 $T=419060 231200 1 0 $X=418870 $Y=228240
X2281 1 2 1375 297 1392 ICV_35 $T=432860 236640 0 0 $X=432670 $Y=236400
X2282 1 2 1391 267 1398 ICV_35 $T=439760 220320 0 0 $X=439570 $Y=220080
X2283 1 2 1412 318 1442 ICV_35 $T=460460 231200 1 0 $X=460270 $Y=228240
X2284 1 2 408 423 1547 ICV_35 $T=515200 236640 0 0 $X=515010 $Y=236400
X2285 1 2 1508 422 1550 ICV_35 $T=516120 225760 1 0 $X=515930 $Y=222800
X2286 1 2 1598 299 1620 ICV_35 $T=553380 198560 1 0 $X=553190 $Y=195600
X2287 1 2 453 317 465 ICV_35 $T=576840 242080 0 0 $X=576650 $Y=241840
X2288 1 2 1642 286 1673 ICV_35 $T=583280 225760 0 0 $X=583090 $Y=225520
X2289 1 2 467 297 474 ICV_35 $T=588800 242080 1 0 $X=588610 $Y=239120
X2290 1 2 473 288 1690 ICV_35 $T=595240 182240 0 0 $X=595050 $Y=182000
X2291 1 2 1688 297 1712 ICV_35 $T=602600 236640 0 0 $X=602410 $Y=236400
X2292 1 2 481 288 485 ICV_35 $T=610880 182240 0 0 $X=610690 $Y=182000
X2293 1 2 1727 300 1769 ICV_35 $T=630660 225760 0 0 $X=630470 $Y=225520
X2294 1 2 499 409 1794 ICV_35 $T=646760 182240 1 0 $X=646570 $Y=179280
X2295 1 2 1795 404 1817 ICV_35 $T=655500 236640 0 0 $X=655310 $Y=236400
X2296 1 2 499 404 1823 ICV_35 $T=659640 182240 0 0 $X=659450 $Y=182000
X2297 1 2 1815 409 1854 ICV_35 $T=672980 204000 1 0 $X=672790 $Y=201040
X2298 1 2 1839 406 1859 ICV_35 $T=674360 231200 1 0 $X=674170 $Y=228240
X2299 1 2 1816 405 1862 ICV_35 $T=677120 198560 1 0 $X=676930 $Y=195600
X2300 1 2 1861 423 1872 ICV_35 $T=682640 220320 1 0 $X=682450 $Y=217360
X2301 1 2 1861 405 1882 ICV_35 $T=685860 220320 0 0 $X=685670 $Y=220080
X2302 1 2 1866 403 1899 ICV_35 $T=695980 209440 1 0 $X=695790 $Y=206480
X2303 1 2 1866 421 1903 ICV_35 $T=697360 204000 0 0 $X=697170 $Y=203760
X2304 1 2 1861 404 1905 ICV_35 $T=698280 225760 0 0 $X=698090 $Y=225520
X2305 1 2 508 403 1910 ICV_35 $T=701040 242080 1 0 $X=700850 $Y=239120
X2306 1 2 1876 404 1912 ICV_35 $T=701960 187680 1 0 $X=701770 $Y=184720
X2307 1 2 1933 422 1941 ICV_35 $T=718060 187680 0 0 $X=717870 $Y=187440
X2308 1 2 513 409 523 ICV_35 $T=729100 182240 1 0 $X=728910 $Y=179280
X2309 1 2 49 34 644 ICV_36 $T=34040 187680 1 0 $X=33850 $Y=184720
X2310 1 2 836 14 862 ICV_36 $T=149960 242080 1 0 $X=149770 $Y=239120
X2311 1 2 125 35 131 ICV_36 $T=160540 182240 1 0 $X=160350 $Y=179280
X2312 1 2 125 34 869 ICV_36 $T=160540 187680 1 0 $X=160350 $Y=184720
X2313 1 2 127 48 912 ICV_36 $T=176640 231200 1 0 $X=176450 $Y=228240
X2314 1 2 897 10 937 ICV_36 $T=191360 182240 0 0 $X=191170 $Y=182000
X2315 1 2 1062 200 1071 ICV_36 $T=258520 209440 0 0 $X=258330 $Y=209200
X2316 1 2 1048 138 1081 ICV_36 $T=261280 242080 1 0 $X=261090 $Y=239120
X2317 1 2 283 200 1199 ICV_36 $T=331660 182240 0 0 $X=331470 $Y=182000
X2318 1 2 1249 317 1245 ICV_36 $T=364320 225760 1 0 $X=364130 $Y=222800
X2319 1 2 1456 297 1478 ICV_36 $T=473800 236640 1 0 $X=473610 $Y=233680
X2320 1 2 1456 288 1501 ICV_36 $T=486680 225760 1 0 $X=486490 $Y=222800
X2321 1 2 1481 317 1521 ICV_36 $T=497260 187680 1 0 $X=497070 $Y=184720
X2322 1 2 1582 317 1603 ICV_36 $T=539120 198560 0 0 $X=538930 $Y=198320
X2323 1 2 481 297 1726 ICV_36 $T=609040 187680 0 0 $X=608850 $Y=187440
X2324 1 2 1917 406 1936 ICV_36 $T=709320 225760 1 0 $X=709130 $Y=222800
X2325 1 2 587 24 610 ICV_37 $T=19780 236640 1 0 $X=19590 $Y=233680
X2326 1 2 49 13 631 ICV_37 $T=33580 193120 0 0 $X=33390 $Y=192880
X2327 1 2 626 12 655 ICV_37 $T=47840 209440 1 0 $X=47650 $Y=206480
X2328 1 2 652 34 684 ICV_37 $T=61640 182240 0 0 $X=61450 $Y=182000
X2329 1 2 702 24 716 ICV_37 $T=75900 225760 1 0 $X=75710 $Y=222800
X2330 1 2 702 20 717 ICV_37 $T=75900 231200 1 0 $X=75710 $Y=228240
X2331 1 2 734 10 736 ICV_37 $T=89700 209440 0 0 $X=89510 $Y=209200
X2332 1 2 86 5 90 ICV_37 $T=89700 242080 0 0 $X=89510 $Y=241840
X2333 1 2 760 20 766 ICV_37 $T=103960 231200 1 0 $X=103770 $Y=228240
X2334 1 2 764 11 778 ICV_37 $T=117760 198560 0 0 $X=117570 $Y=198320
X2335 1 2 760 5 787 ICV_37 $T=117760 231200 0 0 $X=117570 $Y=230960
X2336 1 2 97 25 108 ICV_37 $T=117760 242080 0 0 $X=117570 $Y=241840
X2337 1 2 764 35 803 ICV_37 $T=132020 204000 1 0 $X=131830 $Y=201040
X2338 1 2 764 36 818 ICV_37 $T=132020 209440 1 0 $X=131830 $Y=206480
X2339 1 2 813 33 850 ICV_37 $T=145820 214880 0 0 $X=145630 $Y=214640
X2340 1 2 836 7 847 ICV_37 $T=145820 231200 0 0 $X=145630 $Y=230960
X2341 1 2 836 24 821 ICV_37 $T=145820 236640 0 0 $X=145630 $Y=236400
X2342 1 2 860 35 872 ICV_37 $T=160080 198560 1 0 $X=159890 $Y=195600
X2343 1 2 125 33 143 ICV_37 $T=173880 182240 0 0 $X=173690 $Y=182000
X2344 1 2 860 11 900 ICV_37 $T=173880 193120 0 0 $X=173690 $Y=192880
X2345 1 2 860 34 901 ICV_37 $T=173880 204000 0 0 $X=173690 $Y=203760
X2346 1 2 875 137 880 ICV_37 $T=173880 231200 0 0 $X=173690 $Y=230960
X2347 1 2 875 138 902 ICV_37 $T=173880 236640 0 0 $X=173690 $Y=236400
X2348 1 2 897 34 165 ICV_37 $T=188140 187680 1 0 $X=187950 $Y=184720
X2349 1 2 905 11 907 ICV_37 $T=188140 204000 1 0 $X=187950 $Y=201040
X2350 1 2 897 13 954 ICV_37 $T=201940 187680 0 0 $X=201750 $Y=187440
X2351 1 2 180 201 1012 ICV_37 $T=230000 182240 0 0 $X=229810 $Y=182000
X2352 1 2 962 201 1013 ICV_37 $T=230000 187680 0 0 $X=229810 $Y=187440
X2353 1 2 967 205 1011 ICV_37 $T=230000 214880 0 0 $X=229810 $Y=214640
X2354 1 2 1028 182 1030 ICV_37 $T=244260 193120 1 0 $X=244070 $Y=190160
X2355 1 2 1028 200 1040 ICV_37 $T=244260 198560 1 0 $X=244070 $Y=195600
X2356 1 2 1022 188 1041 ICV_37 $T=244260 204000 1 0 $X=244070 $Y=201040
X2357 1 2 1022 182 1043 ICV_37 $T=244260 209440 1 0 $X=244070 $Y=206480
X2358 1 2 1022 205 1044 ICV_37 $T=244260 220320 1 0 $X=244070 $Y=217360
X2359 1 2 1002 148 1035 ICV_37 $T=244260 231200 1 0 $X=244070 $Y=228240
X2360 1 2 1002 130 1036 ICV_37 $T=244260 236640 1 0 $X=244070 $Y=233680
X2361 1 2 1028 188 1063 ICV_37 $T=258060 187680 0 0 $X=257870 $Y=187440
X2362 1 2 127 243 1098 ICV_37 $T=272320 225760 1 0 $X=272130 $Y=222800
X2363 1 2 1096 201 1088 ICV_37 $T=286120 209440 0 0 $X=285930 $Y=209200
X2364 1 2 1092 149 1122 ICV_37 $T=286120 236640 0 0 $X=285930 $Y=236400
X2365 1 2 250 147 256 ICV_37 $T=286120 242080 0 0 $X=285930 $Y=241840
X2366 1 2 1121 183 1133 ICV_37 $T=300380 204000 1 0 $X=300190 $Y=201040
X2367 1 2 1121 199 1147 ICV_37 $T=300380 220320 1 0 $X=300190 $Y=217360
X2368 1 2 1156 182 1166 ICV_37 $T=314180 198560 0 0 $X=313990 $Y=198320
X2369 1 2 1156 199 1167 ICV_37 $T=314180 204000 0 0 $X=313990 $Y=203760
X2370 1 2 1156 200 1168 ICV_37 $T=314180 209440 0 0 $X=313990 $Y=209200
X2371 1 2 127 271 1037 ICV_37 $T=314180 225760 0 0 $X=313990 $Y=225520
X2372 1 2 1141 183 1188 ICV_37 $T=328440 198560 1 0 $X=328250 $Y=195600
X2373 1 2 1173 279 1189 ICV_37 $T=328440 220320 1 0 $X=328250 $Y=217360
X2374 1 2 1173 267 1190 ICV_37 $T=328440 225760 1 0 $X=328250 $Y=222800
X2375 1 2 1183 201 1214 ICV_37 $T=342240 198560 0 0 $X=342050 $Y=198320
X2376 1 2 1203 284 1215 ICV_37 $T=342240 209440 0 0 $X=342050 $Y=209200
X2377 1 2 127 157 306 ICV_37 $T=342240 231200 0 0 $X=342050 $Y=230960
X2378 1 2 1203 282 1235 ICV_37 $T=356500 225760 1 0 $X=356310 $Y=222800
X2379 1 2 1202 317 1240 ICV_37 $T=356500 236640 1 0 $X=356310 $Y=233680
X2380 1 2 1234 267 1264 ICV_37 $T=370300 204000 0 0 $X=370110 $Y=203760
X2381 1 2 1249 300 1263 ICV_37 $T=370300 231200 0 0 $X=370110 $Y=230960
X2382 1 2 331 300 335 ICV_37 $T=370300 242080 0 0 $X=370110 $Y=241840
X2383 1 2 1252 200 1288 ICV_37 $T=384560 209440 1 0 $X=384370 $Y=206480
X2384 1 2 1249 318 1290 ICV_37 $T=384560 231200 1 0 $X=384370 $Y=228240
X2385 1 2 1301 286 1310 ICV_37 $T=398360 225760 0 0 $X=398170 $Y=225520
X2386 1 2 1301 318 1314 ICV_37 $T=398360 231200 0 0 $X=398170 $Y=230960
X2387 1 2 1308 296 1341 ICV_37 $T=412620 198560 1 0 $X=412430 $Y=195600
X2388 1 2 1308 279 1344 ICV_37 $T=412620 209440 1 0 $X=412430 $Y=206480
X2389 1 2 1339 275 1374 ICV_37 $T=426420 198560 0 0 $X=426230 $Y=198320
X2390 1 2 1391 280 1350 ICV_37 $T=440680 220320 1 0 $X=440490 $Y=217360
X2391 1 2 1391 279 1336 ICV_37 $T=440680 225760 1 0 $X=440490 $Y=222800
X2392 1 2 1375 318 1394 ICV_37 $T=440680 242080 1 0 $X=440490 $Y=239120
X2393 1 2 1395 280 1431 ICV_37 $T=454480 187680 0 0 $X=454290 $Y=187440
X2394 1 2 1395 278 1427 ICV_37 $T=454480 193120 0 0 $X=454290 $Y=192880
X2395 1 2 1412 297 1432 ICV_37 $T=454480 231200 0 0 $X=454290 $Y=230960
X2396 1 2 1440 318 1453 ICV_37 $T=468740 193120 1 0 $X=468550 $Y=190160
X2397 1 2 1415 300 1457 ICV_37 $T=468740 209440 1 0 $X=468550 $Y=206480
X2398 1 2 1474 298 1485 ICV_37 $T=482540 198560 0 0 $X=482350 $Y=198320
X2399 1 2 389 288 1482 ICV_37 $T=482540 236640 0 0 $X=482350 $Y=236400
X2400 1 2 1474 288 1510 ICV_37 $T=496800 209440 1 0 $X=496610 $Y=206480
X2401 1 2 416 421 425 ICV_37 $T=510600 182240 0 0 $X=510410 $Y=182000
X2402 1 2 1526 299 1533 ICV_37 $T=510600 198560 0 0 $X=510410 $Y=198320
X2403 1 2 1504 422 1539 ICV_37 $T=510600 225760 0 0 $X=510410 $Y=225520
X2404 1 2 416 405 434 ICV_37 $T=524860 182240 1 0 $X=524670 $Y=179280
X2405 1 2 1508 406 1559 ICV_37 $T=524860 225760 1 0 $X=524670 $Y=222800
X2406 1 2 1563 318 1595 ICV_37 $T=538660 182240 0 0 $X=538470 $Y=182000
X2407 1 2 1563 298 1596 ICV_37 $T=538660 193120 0 0 $X=538470 $Y=192880
X2408 1 2 1576 423 1597 ICV_37 $T=538660 214880 0 0 $X=538470 $Y=214640
X2409 1 2 1576 421 1583 ICV_37 $T=538660 220320 0 0 $X=538470 $Y=220080
X2410 1 2 1551 423 1589 ICV_37 $T=538660 231200 0 0 $X=538470 $Y=230960
X2411 1 2 1551 404 1585 ICV_37 $T=538660 236640 0 0 $X=538470 $Y=236400
X2412 1 2 1598 288 445 ICV_37 $T=552920 187680 1 0 $X=552730 $Y=184720
X2413 1 2 1594 422 1616 ICV_37 $T=552920 231200 1 0 $X=552730 $Y=228240
X2414 1 2 453 300 456 ICV_37 $T=566720 242080 0 0 $X=566530 $Y=241840
X2415 1 2 453 286 466 ICV_37 $T=580980 242080 1 0 $X=580790 $Y=239120
X2416 1 2 467 286 1689 ICV_37 $T=594780 236640 0 0 $X=594590 $Y=236400
X2417 1 2 467 299 475 ICV_37 $T=594780 242080 0 0 $X=594590 $Y=241840
X2418 1 2 1685 286 1717 ICV_37 $T=609040 220320 1 0 $X=608850 $Y=217360
X2419 1 2 1714 299 1744 ICV_37 $T=622840 209440 0 0 $X=622650 $Y=209200
X2420 1 2 1727 299 1747 ICV_37 $T=622840 225760 0 0 $X=622650 $Y=225520
X2421 1 2 1768 286 1800 ICV_37 $T=650900 198560 0 0 $X=650710 $Y=198320
X2422 1 2 1765 317 1797 ICV_37 $T=650900 220320 0 0 $X=650710 $Y=220080
X2423 1 2 1816 422 1834 ICV_37 $T=665160 187680 1 0 $X=664970 $Y=184720
X2424 1 2 1815 422 1835 ICV_37 $T=665160 204000 1 0 $X=664970 $Y=201040
X2425 1 2 1815 404 1832 ICV_37 $T=665160 209440 1 0 $X=664970 $Y=206480
X2426 1 2 1839 423 1855 ICV_37 $T=678960 225760 0 0 $X=678770 $Y=225520
X2427 1 2 1876 405 1892 ICV_37 $T=693220 198560 1 0 $X=693030 $Y=195600
X2428 1 2 1839 421 1893 ICV_37 $T=693220 236640 1 0 $X=693030 $Y=233680
X2429 1 2 1876 403 1920 ICV_37 $T=707020 193120 0 0 $X=706830 $Y=192880
X2430 1 2 513 406 1953 ICV_37 $T=721280 182240 1 0 $X=721090 $Y=179280
X2431 1 2 1933 403 1956 ICV_37 $T=721280 187680 1 0 $X=721090 $Y=184720
X2432 1 2 1933 421 1949 ICV_37 $T=721280 193120 1 0 $X=721090 $Y=190160
X2433 1 2 1934 406 1957 ICV_37 $T=721280 204000 1 0 $X=721090 $Y=201040
X2434 1 2 1934 422 1950 ICV_37 $T=721280 209440 1 0 $X=721090 $Y=206480
X2435 1 2 1935 406 1955 ICV_37 $T=721280 214880 1 0 $X=721090 $Y=211920
X2436 1 2 1935 422 1931 ICV_37 $T=721280 220320 1 0 $X=721090 $Y=217360
X2437 1 2 1933 405 1959 ICV_37 $T=735080 187680 0 0 $X=734890 $Y=187440
X2438 1 2 1933 423 1900 ICV_37 $T=735080 193120 0 0 $X=734890 $Y=192880
X2439 1 2 1934 409 1960 ICV_37 $T=735080 198560 0 0 $X=734890 $Y=198320
X2440 1 2 1934 405 1958 ICV_37 $T=735080 204000 0 0 $X=734890 $Y=203760
X2441 1 2 1935 404 1974 ICV_37 $T=735080 209440 0 0 $X=734890 $Y=209200
X2442 1 2 1923 423 527 ICV_37 $T=735080 236640 0 0 $X=734890 $Y=236400
X2443 1 2 819 13 842 819 11 805 ICV_38 $T=141680 204000 1 0 $X=141490 $Y=201040
X2444 1 2 819 12 844 819 36 858 ICV_38 $T=142600 209440 1 0 $X=142410 $Y=206480
X2445 1 2 905 33 919 905 35 927 ICV_38 $T=183540 193120 0 0 $X=183350 $Y=192880
X2446 1 2 905 36 922 905 34 918 ICV_38 $T=184920 198560 0 0 $X=184730 $Y=198320
X2447 1 2 159 146 933 159 147 952 ICV_38 $T=192740 242080 1 0 $X=192550 $Y=239120
X2448 1 2 963 182 964 963 183 995 ICV_38 $T=213900 198560 0 0 $X=213710 $Y=198320
X2449 1 2 1066 188 1095 1066 182 1102 ICV_38 $T=270480 187680 0 0 $X=270290 $Y=187440
X2450 1 2 1096 188 1112 1096 183 1123 ICV_38 $T=279680 204000 1 0 $X=279490 $Y=201040
X2451 1 2 1121 200 1140 1121 181 1148 ICV_38 $T=295780 209440 0 0 $X=295590 $Y=209200
X2452 1 2 262 181 1164 262 199 1163 ICV_38 $T=310500 187680 1 0 $X=310310 $Y=184720
X2453 1 2 127 153 304 1202 299 1220 ICV_38 $T=338100 236640 1 0 $X=337910 $Y=233680
X2454 1 2 127 135 321 1202 298 1247 ICV_38 $T=352360 231200 0 0 $X=352170 $Y=230960
X2455 1 2 1306 267 1320 1306 282 1333 ICV_38 $T=400660 220320 0 0 $X=400470 $Y=220080
X2456 1 2 1375 300 372 1375 299 1402 ICV_38 $T=437000 242080 0 0 $X=436810 $Y=241840
X2457 1 2 1535 404 1553 1535 409 1545 ICV_38 $T=520260 204000 0 0 $X=520070 $Y=203760
X2458 1 2 1598 298 444 1598 300 1622 ICV_38 $T=548320 193120 0 0 $X=548130 $Y=192880
X2459 1 2 1686 288 1705 1686 318 1710 ICV_38 $T=598920 204000 0 0 $X=598730 $Y=203760
X2460 1 2 505 421 507 505 422 1851 ICV_38 $T=677120 182240 1 0 $X=676930 $Y=179280
X2461 1 2 1839 409 1863 1839 403 1880 ICV_38 $T=678500 236640 1 0 $X=678310 $Y=233680
X2462 1 2 505 405 1874 505 406 1890 ICV_38 $T=684020 182240 0 0 $X=683830 $Y=182000
X2463 1 2 1876 423 1884 1876 409 1907 ICV_38 $T=692300 187680 0 0 $X=692110 $Y=187440
X2464 1 2 1861 406 1897 1867 406 1922 ICV_38 $T=699660 220320 1 0 $X=699470 $Y=217360
X2465 1 2 654 57 19 ICV_39 $T=70840 187680 1 0 $X=70650 $Y=184720
X2466 1 2 732 710 50 ICV_39 $T=93840 193120 1 0 $X=93650 $Y=190160
X2467 1 2 749 93 19 ICV_39 $T=98900 193120 1 0 $X=98710 $Y=190160
X2468 1 2 742 87 32 ICV_39 $T=98900 231200 1 0 $X=98710 $Y=228240
X2469 1 2 740 691 28 ICV_39 $T=99360 225760 0 0 $X=99170 $Y=225520
X2470 1 2 756 87 39 ICV_39 $T=104420 231200 0 0 $X=104230 $Y=230960
X2471 1 2 953 177 19 ICV_39 $T=208840 193120 0 0 $X=208650 $Y=192880
X2472 1 2 1033 1020 155 ICV_39 $T=253000 231200 0 0 $X=252810 $Y=230960
X2473 1 2 1064 1055 152 ICV_39 $T=264960 242080 0 0 $X=264770 $Y=241840
X2474 1 2 1077 1078 216 ICV_39 $T=269560 214880 0 0 $X=269370 $Y=214640
X2475 1 2 1075 1078 196 ICV_39 $T=281060 204000 0 0 $X=280870 $Y=203760
X2476 1 2 1127 258 219 ICV_39 $T=300840 193120 1 0 $X=300650 $Y=190160
X2477 1 2 272 274 152 ICV_39 $T=315560 242080 0 0 $X=315370 $Y=241840
X2478 1 2 1166 1172 185 ICV_39 $T=323380 198560 1 0 $X=323190 $Y=195600
X2479 1 2 1176 1172 216 ICV_39 $T=328900 209440 1 0 $X=328710 $Y=206480
X2480 1 2 1254 1255 216 ICV_39 $T=372140 182240 0 0 $X=371950 $Y=182000
X2481 1 2 1258 1239 263 ICV_39 $T=379040 209440 0 0 $X=378850 $Y=209200
X2482 1 2 1264 1239 194 ICV_39 $T=379500 209440 1 0 $X=379310 $Y=206480
X2483 1 2 1288 1268 212 ICV_39 $T=391000 204000 1 0 $X=390810 $Y=201040
X2484 1 2 345 336 255 ICV_39 $T=393300 242080 0 0 $X=393110 $Y=241840
X2485 1 2 1321 1327 194 ICV_39 $T=413080 204000 1 0 $X=412890 $Y=201040
X2486 1 2 1382 1351 231 ICV_39 $T=435620 193120 1 0 $X=435430 $Y=190160
X2487 1 2 1527 420 414 ICV_39 $T=511060 242080 0 0 $X=510870 $Y=241840
X2488 1 2 1588 1580 412 ICV_39 $T=547400 225760 0 0 $X=547210 $Y=225520
X2489 1 2 468 1667 330 ICV_39 $T=589720 182240 0 0 $X=589530 $Y=182000
X2490 1 2 1672 1652 271 ICV_39 $T=589720 214880 0 0 $X=589530 $Y=214640
X2491 1 2 1756 1736 329 ICV_39 $T=632040 214880 1 0 $X=631850 $Y=211920
X2492 1 2 1741 1745 330 ICV_39 $T=632040 220320 1 0 $X=631850 $Y=217360
X2493 1 2 1918 1885 415 ICV_39 $T=712080 193120 1 0 $X=711890 $Y=190160
X2494 1 2 1957 1954 415 ICV_39 $T=730020 198560 0 0 $X=729830 $Y=198320
X2495 1 2 1961 1901 424 ICV_39 $T=737840 182240 0 0 $X=737650 $Y=182000
X2496 1 2 1962 1932 429 ICV_39 $T=737840 204000 1 0 $X=737650 $Y=201040
X2497 1 2 1969 1932 424 ICV_39 $T=737840 214880 0 0 $X=737650 $Y=214640
X2498 1 2 621 601 50 ICV_40 $T=35880 198560 1 0 $X=35690 $Y=195600
X2499 1 2 769 750 28 ICV_40 $T=111780 204000 0 0 $X=111590 $Y=203760
X2500 1 2 762 93 44 ICV_40 $T=116380 187680 1 0 $X=116190 $Y=184720
X2501 1 2 782 98 46 ICV_40 $T=139840 231200 0 0 $X=139650 $Y=230960
X2502 1 2 848 119 44 ICV_40 $T=154100 187680 1 0 $X=153910 $Y=184720
X2503 1 2 908 881 27 ICV_40 $T=188600 209440 1 0 $X=188410 $Y=206480
X2504 1 2 938 929 28 ICV_40 $T=201480 220320 1 0 $X=201290 $Y=217360
X2505 1 2 1042 1046 196 ICV_40 $T=252080 198560 0 0 $X=251890 $Y=198320
X2506 1 2 1132 258 216 ICV_40 $T=300840 198560 1 0 $X=300650 $Y=195600
X2507 1 2 1179 292 216 ICV_40 $T=330740 182240 1 0 $X=330550 $Y=179280
X2508 1 2 1198 1201 211 ICV_40 $T=340400 204000 1 0 $X=340210 $Y=201040
X2509 1 2 1215 1212 254 ICV_40 $T=350520 214880 1 0 $X=350330 $Y=211920
X2510 1 2 1328 351 219 ICV_40 $T=413080 182240 1 0 $X=412890 $Y=179280
X2511 1 2 1436 1438 255 ICV_40 $T=462760 198560 1 0 $X=462570 $Y=195600
X2512 1 2 1473 1477 238 ICV_40 $T=485300 236640 1 0 $X=485110 $Y=233680
X2513 1 2 1595 1581 329 ICV_40 $T=546940 187680 1 0 $X=546750 $Y=184720
X2514 1 2 1614 443 251 ICV_40 $T=557060 182240 1 0 $X=556870 $Y=179280
X2515 1 2 1638 1636 329 ICV_40 $T=567640 209440 1 0 $X=567450 $Y=206480
X2516 1 2 1682 1649 329 ICV_40 $T=592940 204000 1 0 $X=592750 $Y=201040
X2517 1 2 490 484 329 ICV_40 $T=630200 242080 0 0 $X=630010 $Y=241840
X2518 1 2 1842 1831 415 ICV_40 $T=675280 193120 1 0 $X=675090 $Y=190160
X2519 1 2 1882 1844 413 ICV_40 $T=693680 220320 1 0 $X=693490 $Y=217360
X2520 1 2 1895 1844 427 ICV_40 $T=701040 214880 0 0 $X=700850 $Y=214640
X2521 1 2 1922 1886 415 ICV_40 $T=715300 214880 1 0 $X=715110 $Y=211920
X2522 1 2 1965 1938 414 ICV_40 $T=736920 225760 0 0 $X=736730 $Y=225520
X2523 1 2 524 519 414 ICV_40 $T=736920 242080 0 0 $X=736730 $Y=241840
X2524 1 2 9 35 614 ICV_41 $T=23000 187680 0 0 $X=22810 $Y=187440
X2525 1 2 588 34 613 ICV_41 $T=23000 204000 0 0 $X=22810 $Y=203760
X2526 1 2 734 36 754 ICV_41 $T=93840 225760 1 0 $X=93650 $Y=222800
X2527 1 2 813 13 856 ICV_41 $T=149500 220320 1 0 $X=149310 $Y=217360
X2528 1 2 125 36 879 ICV_41 $T=163300 187680 0 0 $X=163110 $Y=187440
X2529 1 2 866 34 903 ICV_41 $T=177560 214880 1 0 $X=177370 $Y=211920
X2530 1 2 127 218 1029 ICV_41 $T=240120 220320 0 0 $X=239930 $Y=220080
X2531 1 2 127 232 892 ICV_41 $T=252080 220320 1 0 $X=251890 $Y=217360
X2532 1 2 127 238 1065 ICV_41 $T=261740 236640 1 0 $X=261550 $Y=233680
X2533 1 2 127 263 1001 ICV_41 $T=304060 220320 0 0 $X=303870 $Y=220080
X2534 1 2 1183 181 1222 ICV_41 $T=346380 204000 1 0 $X=346190 $Y=201040
X2535 1 2 1395 284 1410 ICV_41 $T=443900 187680 1 0 $X=443710 $Y=184720
X2536 1 2 1412 288 1448 ICV_41 $T=468280 236640 0 0 $X=468090 $Y=236400
X2537 1 2 416 404 1544 ICV_41 $T=514740 182240 1 0 $X=514550 $Y=179280
X2538 1 2 1535 422 1573 ICV_41 $T=528540 214880 0 0 $X=528350 $Y=214640
X2539 1 2 1551 403 1587 ICV_41 $T=535440 242080 1 0 $X=535250 $Y=239120
X2540 1 2 1594 404 1610 ICV_41 $T=546480 236640 0 0 $X=546290 $Y=236400
X2541 1 2 1582 318 1621 ICV_41 $T=556600 204000 0 0 $X=556410 $Y=203760
X2542 1 2 1765 318 1758 ICV_41 $T=640780 220320 0 0 $X=640590 $Y=220080
X2543 1 2 1839 405 1871 ICV_41 $T=682640 231200 1 0 $X=682450 $Y=228240
X2544 1 2 1917 422 1946 ICV_41 $T=717600 220320 0 0 $X=717410 $Y=220080
X2545 1 2 658 659 50 669 659 48 ICV_44 $T=52900 187680 0 0 $X=52710 $Y=187440
X2546 1 2 787 773 8 791 773 40 ICV_44 $T=118220 236640 0 0 $X=118030 $Y=236400
X2547 1 2 833 808 39 832 808 32 ICV_44 $T=141220 231200 1 0 $X=141030 $Y=228240
X2548 1 2 975 974 135 970 974 152 ICV_44 $T=218960 225760 0 0 $X=218770 $Y=225520
X2549 1 2 1043 1046 185 1045 1046 219 ICV_44 $T=252080 209440 1 0 $X=251890 $Y=206480
X2550 1 2 1050 234 196 1047 224 219 ICV_44 $T=255760 182240 1 0 $X=255570 $Y=179280
X2551 1 2 1071 1078 212 1072 1078 185 ICV_44 $T=268640 209440 0 0 $X=268450 $Y=209200
X2552 1 2 1143 1136 195 1146 1136 185 ICV_44 $T=304980 204000 0 0 $X=304790 $Y=203760
X2553 1 2 1199 292 212 1207 1193 195 ICV_44 $T=340400 187680 1 0 $X=340210 $Y=184720
X2554 1 2 1281 1280 232 1278 1280 263 ICV_44 $T=385020 225760 1 0 $X=384830 $Y=222800
X2555 1 2 1528 1530 424 1525 1530 413 ICV_44 $T=511060 220320 0 0 $X=510870 $Y=220080
X2556 1 2 1698 1704 285 1710 1704 329 ICV_44 $T=604900 209440 0 0 $X=604710 $Y=209200
X2557 1 2 1763 1739 251 1762 1739 285 ICV_44 $T=635260 236640 0 0 $X=635070 $Y=236400
X2558 1 2 511 506 414 1896 506 424 ICV_44 $T=703340 182240 1 0 $X=703150 $Y=179280
X2559 1 2 1908 1865 414 1909 1865 424 ICV_44 $T=707480 198560 0 0 $X=707290 $Y=198320
X2560 1 2 1958 1954 413 1960 1954 424 ICV_44 $T=729100 204000 1 0 $X=728910 $Y=201040
X2561 1 2 589 12 599 ICV_47 $T=10580 220320 1 0 $X=10390 $Y=217360
X2562 1 2 588 33 620 ICV_47 $T=22540 193120 0 0 $X=22350 $Y=192880
X2563 1 2 608 14 649 ICV_47 $T=36800 236640 1 0 $X=36610 $Y=233680
X2564 1 2 652 35 658 ICV_47 $T=48300 187680 1 0 $X=48110 $Y=184720
X2565 1 2 652 36 669 ICV_47 $T=50600 193120 0 0 $X=50410 $Y=192880
X2566 1 2 74 11 88 ICV_47 $T=83260 182240 1 0 $X=83070 $Y=179280
X2567 1 2 735 34 743 ICV_47 $T=90160 204000 0 0 $X=89970 $Y=203760
X2568 1 2 734 33 745 ICV_47 $T=90160 214880 0 0 $X=89970 $Y=214640
X2569 1 2 97 7 763 ICV_47 $T=105800 242080 0 0 $X=105610 $Y=241840
X2570 1 2 764 34 786 ICV_47 $T=109020 209440 0 0 $X=108830 $Y=209200
X2571 1 2 784 12 820 ICV_47 $T=130640 193120 0 0 $X=130450 $Y=192880
X2572 1 2 793 6 832 ICV_47 $T=132480 225760 1 0 $X=132290 $Y=222800
X2573 1 2 793 20 833 ICV_47 $T=132480 231200 1 0 $X=132290 $Y=228240
X2574 1 2 819 35 843 ICV_47 $T=144900 198560 1 0 $X=144710 $Y=195600
X2575 1 2 125 12 878 ICV_47 $T=161460 182240 0 0 $X=161270 $Y=182000
X2576 1 2 127 50 883 ICV_47 $T=164220 220320 0 0 $X=164030 $Y=220080
X2577 1 2 127 40 904 ICV_47 $T=174340 225760 0 0 $X=174150 $Y=225520
X2578 1 2 897 35 913 ICV_47 $T=179400 193120 1 0 $X=179210 $Y=190160
X2579 1 2 127 18 921 ICV_47 $T=183080 225760 0 0 $X=182890 $Y=225520
X2580 1 2 159 138 939 ICV_47 $T=193200 236640 0 0 $X=193010 $Y=236400
X2581 1 2 955 147 970 ICV_47 $T=207460 242080 1 0 $X=207270 $Y=239120
X2582 1 2 127 19 984 ICV_47 $T=213900 220320 0 0 $X=213710 $Y=220080
X2583 1 2 1022 199 1031 ICV_47 $T=237820 214880 0 0 $X=237630 $Y=214640
X2584 1 2 1022 200 1038 ICV_47 $T=241960 209440 0 0 $X=241770 $Y=209200
X2585 1 2 1048 149 1060 ICV_47 $T=252540 242080 1 0 $X=252350 $Y=239120
X2586 1 2 1062 183 1075 ICV_47 $T=260820 204000 0 0 $X=260630 $Y=203760
X2587 1 2 1096 200 1111 ICV_47 $T=277380 209440 0 0 $X=277190 $Y=209200
X2588 1 2 127 254 943 ICV_47 $T=289800 220320 1 0 $X=289610 $Y=217360
X2589 1 2 283 205 1179 ICV_47 $T=322920 182240 0 0 $X=322730 $Y=182000
X2590 1 2 1197 205 1231 ICV_47 $T=350980 193120 0 0 $X=350790 $Y=192880
X2591 1 2 1234 296 1246 ICV_47 $T=358340 220320 1 0 $X=358150 $Y=217360
X2592 1 2 1249 288 1259 ICV_47 $T=368460 231200 1 0 $X=368270 $Y=228240
X2593 1 2 1262 275 1277 ICV_47 $T=375820 214880 1 0 $X=375630 $Y=211920
X2594 1 2 1252 183 1286 ICV_47 $T=381800 198560 0 0 $X=381610 $Y=198320
X2595 1 2 331 317 342 ICV_47 $T=382260 236640 0 0 $X=382070 $Y=236400
X2596 1 2 339 182 1294 ICV_47 $T=385020 182240 1 0 $X=384830 $Y=179280
X2597 1 2 1262 296 1296 ICV_47 $T=386860 220320 0 0 $X=386670 $Y=220080
X2598 1 2 1308 280 1318 ICV_47 $T=398820 204000 0 0 $X=398630 $Y=203760
X2599 1 2 1306 280 1335 ICV_47 $T=408020 209440 0 0 $X=407830 $Y=209200
X2600 1 2 361 297 1356 ICV_47 $T=417220 242080 1 0 $X=417030 $Y=239120
X2601 1 2 1369 278 1387 ICV_47 $T=429180 204000 1 0 $X=428990 $Y=201040
X2602 1 2 373 282 377 ICV_47 $T=446200 182240 1 0 $X=446010 $Y=179280
X2603 1 2 1415 288 1436 ICV_47 $T=454940 198560 0 0 $X=454750 $Y=198320
X2604 1 2 1428 297 1443 ICV_47 $T=459540 214880 1 0 $X=459350 $Y=211920
X2605 1 2 1440 317 1469 ICV_47 $T=472880 187680 0 0 $X=472690 $Y=187440
X2606 1 2 1456 300 1479 ICV_47 $T=476560 231200 1 0 $X=476370 $Y=228240
X2607 1 2 1476 267 1475 ICV_47 $T=483000 214880 0 0 $X=482810 $Y=214640
X2608 1 2 1481 288 1497 ICV_47 $T=486220 187680 1 0 $X=486030 $Y=184720
X2609 1 2 1535 421 1552 ICV_47 $T=516120 214880 1 0 $X=515930 $Y=211920
X2610 1 2 1563 286 1579 ICV_47 $T=531300 193120 1 0 $X=531110 $Y=190160
X2611 1 2 1576 403 1588 ICV_47 $T=534980 225760 1 0 $X=534790 $Y=222800
X2612 1 2 1642 299 1655 ICV_47 $T=571780 236640 1 0 $X=571590 $Y=233680
X2613 1 2 1643 299 1657 ICV_47 $T=572240 220320 1 0 $X=572050 $Y=217360
X2614 1 2 1637 300 1663 ICV_47 $T=576380 204000 0 0 $X=576190 $Y=203760
X2615 1 2 1643 300 1672 ICV_47 $T=581440 214880 1 0 $X=581250 $Y=211920
X2616 1 2 1686 286 1706 ICV_47 $T=598000 209440 1 0 $X=597810 $Y=206480
X2617 1 2 1714 288 1732 ICV_47 $T=613640 204000 1 0 $X=613450 $Y=201040
X2618 1 2 1688 299 1735 ICV_47 $T=613640 242080 0 0 $X=613450 $Y=241840
X2619 1 2 1765 288 1789 ICV_47 $T=639400 220320 1 0 $X=639210 $Y=217360
X2620 1 2 1743 318 1791 ICV_47 $T=639860 231200 1 0 $X=639670 $Y=228240
X2621 1 2 1923 403 1942 ICV_47 $T=714380 231200 0 0 $X=714190 $Y=230960
X2622 1 2 1933 409 1961 ICV_47 $T=726340 187680 0 0 $X=726150 $Y=187440
X2623 1 2 1935 423 1962 ICV_47 $T=726340 214880 0 0 $X=726150 $Y=214640
X2624 1 2 657 641 19 ICV_48 $T=57500 214880 0 0 $X=57310 $Y=214640
X2625 1 2 75 76 50 ICV_48 $T=71760 182240 1 0 $X=71570 $Y=179280
X2626 1 2 700 681 28 ICV_48 $T=71760 204000 1 0 $X=71570 $Y=201040
X2627 1 2 712 694 45 ICV_48 $T=85560 220320 0 0 $X=85370 $Y=220080
X2628 1 2 754 691 48 ICV_48 $T=99820 214880 1 0 $X=99630 $Y=211920
X2629 1 2 755 757 31 ICV_48 $T=99820 220320 1 0 $X=99630 $Y=217360
X2630 1 2 806 808 8 ICV_48 $T=127880 236640 1 0 $X=127690 $Y=233680
X2631 1 2 913 177 50 ICV_48 $T=212060 193120 1 0 $X=211870 $Y=190160
X2632 1 2 1103 1087 198 ICV_48 $T=281980 193120 0 0 $X=281790 $Y=192880
X2633 1 2 1134 1136 219 ICV_48 $T=296240 209440 1 0 $X=296050 $Y=206480
X2634 1 2 1192 1193 219 ICV_48 $T=338100 187680 0 0 $X=337910 $Y=187440
X2635 1 2 1189 1184 263 ICV_48 $T=338100 225760 0 0 $X=337910 $Y=225520
X2636 1 2 1245 1248 330 ICV_48 $T=366160 209440 0 0 $X=365970 $Y=209200
X2637 1 2 1247 309 285 ICV_48 $T=366160 236640 0 0 $X=365970 $Y=236400
X2638 1 2 1295 1297 263 ICV_48 $T=394220 193120 0 0 $X=394030 $Y=192880
X2639 1 2 1296 1280 231 ICV_48 $T=394220 214880 0 0 $X=394030 $Y=214640
X2640 1 2 1349 1351 232 ICV_48 $T=422280 193120 0 0 $X=422090 $Y=192880
X2641 1 2 1320 1297 194 ICV_48 $T=422280 236640 0 0 $X=422090 $Y=236400
X2642 1 2 1386 364 263 ICV_48 $T=436540 187680 1 0 $X=436350 $Y=184720
X2643 1 2 1370 1366 329 ICV_48 $T=436540 236640 1 0 $X=436350 $Y=233680
X2644 1 2 1411 1337 231 ICV_48 $T=450340 220320 0 0 $X=450150 $Y=220080
X2645 1 2 1442 1422 329 ICV_48 $T=464600 236640 1 0 $X=464410 $Y=233680
X2646 1 2 1463 1423 251 ICV_48 $T=478400 220320 0 0 $X=478210 $Y=220080
X2647 1 2 1460 1423 255 ICV_48 $T=478400 225760 0 0 $X=478210 $Y=225520
X2648 1 2 1545 1546 424 ICV_48 $T=520720 209440 1 0 $X=520530 $Y=206480
X2649 1 2 435 432 414 ICV_48 $T=534520 187680 0 0 $X=534330 $Y=187440
X2650 1 2 1571 1546 415 ICV_48 $T=534520 209440 0 0 $X=534330 $Y=209200
X2651 1 2 1590 1581 249 ICV_48 $T=548780 198560 1 0 $X=548590 $Y=195600
X2652 1 2 1604 1580 427 ICV_48 $T=548780 214880 1 0 $X=548590 $Y=211920
X2653 1 2 1623 1605 285 ICV_48 $T=562580 198560 0 0 $X=562390 $Y=198320
X2654 1 2 1700 1704 330 ICV_48 $T=604900 198560 1 0 $X=604710 $Y=195600
X2655 1 2 1897 1844 415 ICV_48 $T=702880 220320 0 0 $X=702690 $Y=220080
X2656 1 2 1898 510 413 ICV_48 $T=702880 242080 0 0 $X=702690 $Y=241840
X2657 1 2 588 36 615 615 601 48 ICV_49 $T=20240 204000 1 0 $X=20050 $Y=201040
X2658 1 2 49 36 643 643 57 48 ICV_49 $T=34040 182240 0 0 $X=33850 $Y=182000
X2659 1 2 703 36 726 724 710 28 ICV_49 $T=76360 209440 1 0 $X=76170 $Y=206480
X2660 1 2 89 35 752 752 93 50 ICV_49 $T=90160 182240 0 0 $X=89970 $Y=182000
X2661 1 2 86 7 753 753 87 18 ICV_49 $T=90160 231200 0 0 $X=89970 $Y=230960
X2662 1 2 89 12 777 777 93 28 ICV_49 $T=104420 182240 1 0 $X=104230 $Y=179280
X2663 1 2 104 36 812 809 110 28 ICV_49 $T=123740 182240 0 0 $X=123550 $Y=182000
X2664 1 2 793 14 815 811 808 46 ICV_49 $T=125580 231200 0 0 $X=125390 $Y=230960
X2665 1 2 1092 148 1105 1105 1100 156 ICV_49 $T=272780 231200 1 0 $X=272590 $Y=228240
X2666 1 2 1308 284 1338 1338 1327 254 ICV_49 $T=407560 204000 0 0 $X=407370 $Y=203760
X2667 1 2 1369 275 1384 1385 1368 252 ICV_49 $T=426880 209440 0 0 $X=426690 $Y=209200
X2668 1 2 1428 300 1461 1461 1423 271 ICV_49 $T=469200 214880 1 0 $X=469010 $Y=211920
X2669 1 2 1481 318 1502 1497 1499 255 ICV_49 $T=487140 187680 0 0 $X=486950 $Y=187440
X2670 1 2 1504 421 1542 1542 1520 430 ICV_49 $T=509220 236640 1 0 $X=509030 $Y=233680
X2671 1 2 1582 288 1624 1624 1605 255 ICV_49 $T=553380 209440 1 0 $X=553190 $Y=206480
X2672 1 2 1594 409 1633 1629 1612 413 ICV_49 $T=557520 236640 1 0 $X=557330 $Y=233680
X2673 1 2 1637 286 1648 1648 1649 251 ICV_49 $T=567180 198560 0 0 $X=566990 $Y=198320
X2674 1 2 488 317 491 492 493 251 ICV_49 $T=622380 182240 1 0 $X=622190 $Y=179280
X2675 1 2 488 298 1750 1755 493 249 ICV_49 $T=622380 193120 1 0 $X=622190 $Y=190160
X2676 1 2 1743 288 1785 1788 1739 249 ICV_49 $T=637560 236640 1 0 $X=637370 $Y=233680
X2677 1 2 586 3 8 587 14 17 ICV_51 $T=6900 242080 1 0 $X=6710 $Y=239120
X2678 1 2 614 15 50 49 10 647 ICV_51 $T=34040 187680 0 0 $X=33850 $Y=187440
X2679 1 2 689 73 8 702 5 689 ICV_51 $T=68540 236640 0 0 $X=68350 $Y=236400
X2680 1 2 733 87 46 86 20 756 ICV_51 $T=89240 236640 1 0 $X=89050 $Y=233680
X2681 1 2 711 710 19 735 13 776 ICV_51 $T=102580 193120 0 0 $X=102390 $Y=192880
X2682 1 2 821 824 46 836 21 845 ICV_51 $T=138460 242080 1 0 $X=138270 $Y=239120
X2683 1 2 845 824 40 836 25 863 ICV_51 $T=149040 242080 0 0 $X=148850 $Y=241840
X2684 1 2 903 881 45 911 35 923 ICV_51 $T=182160 214880 0 0 $X=181970 $Y=214640
X2685 1 2 973 974 155 955 148 999 ICV_51 $T=218500 231200 1 0 $X=218310 $Y=228240
X2686 1 2 1060 1055 157 1048 130 1080 ICV_51 $T=259900 236640 0 0 $X=259710 $Y=236400
X2687 1 2 1211 1212 252 1203 280 1233 ICV_51 $T=348220 214880 0 0 $X=348030 $Y=214640
X2688 1 2 1228 1212 263 127 156 327 ICV_51 $T=356960 225760 0 0 $X=356770 $Y=225520
X2689 1 2 1238 1239 232 1234 278 1256 ICV_51 $T=362940 214880 1 0 $X=362750 $Y=211920
X2690 1 2 1259 1248 255 1262 282 1282 ICV_51 $T=375360 220320 0 0 $X=375170 $Y=220080
X2691 1 2 1277 1280 252 1262 284 1299 ICV_51 $T=384100 209440 0 0 $X=383910 $Y=209200
X2692 1 2 1377 1351 194 1395 282 1407 ICV_51 $T=439300 193120 0 0 $X=439110 $Y=192880
X2693 1 2 1419 1422 285 1412 300 1444 ICV_51 $T=456780 236640 0 0 $X=456590 $Y=236400
X2694 1 2 1421 1423 330 1428 299 1445 ICV_51 $T=457240 220320 0 0 $X=457050 $Y=220080
X2695 1 2 1424 1423 329 1428 318 1424 ICV_51 $T=458160 214880 0 0 $X=457970 $Y=214640
X2696 1 2 1443 1423 249 1428 286 1463 ICV_51 $T=469200 220320 1 0 $X=469010 $Y=217360
X2697 1 2 1475 1465 194 1476 279 1462 ICV_51 $T=482080 220320 1 0 $X=481890 $Y=217360
X2698 1 2 1533 1534 238 1526 286 1556 ICV_51 $T=516580 193120 0 0 $X=516390 $Y=192880
X2699 1 2 1583 1580 430 1576 422 1604 ICV_51 $T=541420 220320 1 0 $X=541230 $Y=217360
X2700 1 2 1616 1612 427 1617 298 1635 ICV_51 $T=556600 225760 1 0 $X=556410 $Y=222800
X2701 1 2 1647 1649 285 463 318 1665 ICV_51 $T=576380 187680 0 0 $X=576190 $Y=187440
X2702 1 2 1679 471 329 473 297 1692 ICV_51 $T=592480 187680 1 0 $X=592290 $Y=184720
X2703 1 2 1681 1653 255 1688 300 1708 ICV_51 $T=597540 236640 1 0 $X=597350 $Y=233680
X2704 1 2 1706 1704 251 1714 300 1729 ICV_51 $T=609500 209440 1 0 $X=609310 $Y=206480
X2705 1 2 628 619 18 ICV_52 $T=35880 225760 0 0 $X=35690 $Y=225520
X2706 1 2 695 672 39 ICV_52 $T=70380 231200 1 0 $X=70190 $Y=228240
X2707 1 2 849 807 44 ICV_52 $T=157780 198560 0 0 $X=157590 $Y=198320
X2708 1 2 949 177 48 ICV_52 $T=210680 187680 1 0 $X=210490 $Y=184720
X2709 1 2 1025 1020 152 ICV_52 $T=238740 236640 1 0 $X=238550 $Y=233680
X2710 1 2 1070 1078 198 ICV_52 $T=272780 220320 1 0 $X=272590 $Y=217360
X2711 1 2 259 260 153 ICV_52 $T=294860 225760 1 0 $X=294670 $Y=222800
X2712 1 2 1217 1212 194 ICV_52 $T=351440 225760 0 0 $X=351250 $Y=225520
X2713 1 2 1231 1193 216 ICV_52 $T=359260 193120 1 0 $X=359070 $Y=190160
X2714 1 2 1233 1212 232 ICV_52 $T=364780 220320 0 0 $X=364590 $Y=220080
X2715 1 2 1309 1311 255 ICV_52 $T=407100 231200 1 0 $X=406910 $Y=228240
X2716 1 2 1410 1347 254 ICV_52 $T=454940 193120 1 0 $X=454750 $Y=190160
X2717 1 2 1518 1491 329 ICV_52 $T=505540 198560 1 0 $X=505350 $Y=195600
X2718 1 2 1645 1649 255 ICV_52 $T=576380 193120 0 0 $X=576190 $Y=192880
X2719 1 2 1747 1745 238 ICV_52 $T=631580 225760 1 0 $X=631390 $Y=222800
X2720 1 2 1854 1826 424 ICV_52 $T=680340 204000 0 0 $X=680150 $Y=203760
X2721 1 2 1858 1831 424 ICV_52 $T=681260 193120 1 0 $X=681070 $Y=190160
X2722 1 2 1871 1856 413 ICV_52 $T=693680 231200 1 0 $X=693490 $Y=228240
X2723 1 2 1968 510 414 ICV_52 $T=737380 231200 0 0 $X=737190 $Y=230960
X2724 1 2 29 2 12 1 sky130_fd_sc_hd__clkbuf_16 $T=22080 225760 1 0 $X=21890 $Y=222800
X2725 1 2 61 2 36 1 sky130_fd_sc_hd__clkbuf_16 $T=48300 225760 1 0 $X=48110 $Y=222800
X2726 1 2 29 2 25 1 sky130_fd_sc_hd__clkbuf_16 $T=48300 242080 1 0 $X=48110 $Y=239120
X2727 1 2 61 2 21 1 sky130_fd_sc_hd__clkbuf_16 $T=49680 242080 0 0 $X=49490 $Y=241840
X2728 1 2 81 2 13 1 sky130_fd_sc_hd__clkbuf_16 $T=84640 225760 1 0 $X=84450 $Y=222800
X2729 1 2 82 2 20 1 sky130_fd_sc_hd__clkbuf_16 $T=86020 231200 1 0 $X=85830 $Y=228240
X2730 1 2 81 2 7 1 sky130_fd_sc_hd__clkbuf_16 $T=90160 225760 0 0 $X=89970 $Y=225520
X2731 1 2 95 2 99 1 sky130_fd_sc_hd__clkbuf_16 $T=102580 204000 0 0 $X=102390 $Y=203760
X2732 1 2 96 2 26 1 sky130_fd_sc_hd__clkbuf_16 $T=104420 225760 1 0 $X=104230 $Y=222800
X2733 1 2 105 2 6 1 sky130_fd_sc_hd__clkbuf_16 $T=120520 225760 1 0 $X=120330 $Y=222800
X2734 1 2 105 2 10 1 sky130_fd_sc_hd__clkbuf_16 $T=124200 220320 0 0 $X=124010 $Y=220080
X2735 1 2 82 2 33 1 sky130_fd_sc_hd__clkbuf_16 $T=132480 214880 1 0 $X=132290 $Y=211920
X2736 1 2 117 2 24 1 sky130_fd_sc_hd__clkbuf_16 $T=147200 225760 0 0 $X=147010 $Y=225520
X2737 1 2 120 2 14 1 sky130_fd_sc_hd__clkbuf_16 $T=155020 231200 0 0 $X=154830 $Y=230960
X2738 1 2 120 2 34 1 sky130_fd_sc_hd__clkbuf_16 $T=156400 225760 0 0 $X=156210 $Y=225520
X2739 1 2 124 2 11 1 sky130_fd_sc_hd__clkbuf_16 $T=160540 225760 1 0 $X=160350 $Y=222800
X2740 1 2 124 2 5 1 sky130_fd_sc_hd__clkbuf_16 $T=160540 236640 1 0 $X=160350 $Y=233680
X2741 1 2 117 2 35 1 sky130_fd_sc_hd__clkbuf_16 $T=161920 220320 1 0 $X=161730 $Y=217360
X2742 1 2 245 2 178 1 sky130_fd_sc_hd__clkbuf_16 $T=276460 182240 1 0 $X=276270 $Y=179280
X2743 1 2 127 2 266 1 sky130_fd_sc_hd__clkbuf_16 $T=301300 198560 0 0 $X=301110 $Y=198320
X2744 1 2 120 2 267 1 sky130_fd_sc_hd__clkbuf_16 $T=301760 225760 1 0 $X=301570 $Y=222800
X2745 1 2 105 2 275 1 sky130_fd_sc_hd__clkbuf_16 $T=308200 220320 1 0 $X=308010 $Y=217360
X2746 1 2 82 2 278 1 sky130_fd_sc_hd__clkbuf_16 $T=312800 214880 1 0 $X=312610 $Y=211920
X2747 1 2 117 2 280 1 sky130_fd_sc_hd__clkbuf_16 $T=314640 214880 0 0 $X=314450 $Y=214640
X2748 1 2 124 2 279 1 sky130_fd_sc_hd__clkbuf_16 $T=314640 220320 0 0 $X=314450 $Y=220080
X2749 1 2 29 2 282 1 sky130_fd_sc_hd__clkbuf_16 $T=315100 225760 1 0 $X=314910 $Y=222800
X2750 1 2 245 2 128 1 sky130_fd_sc_hd__clkbuf_16 $T=315560 242080 1 0 $X=315370 $Y=239120
X2751 1 2 81 2 284 1 sky130_fd_sc_hd__clkbuf_16 $T=317400 220320 1 0 $X=317210 $Y=217360
X2752 1 2 276 2 286 1 sky130_fd_sc_hd__clkbuf_16 $T=317400 231200 1 0 $X=317210 $Y=228240
X2753 1 2 277 2 288 1 sky130_fd_sc_hd__clkbuf_16 $T=319240 236640 1 0 $X=319050 $Y=233680
X2754 1 2 127 2 287 1 sky130_fd_sc_hd__clkbuf_16 $T=321080 236640 0 0 $X=320890 $Y=236400
X2755 1 2 61 2 296 1 sky130_fd_sc_hd__clkbuf_16 $T=328900 225760 0 0 $X=328710 $Y=225520
X2756 1 2 289 2 297 1 sky130_fd_sc_hd__clkbuf_16 $T=328900 231200 1 0 $X=328710 $Y=228240
X2757 1 2 290 2 298 1 sky130_fd_sc_hd__clkbuf_16 $T=328900 236640 1 0 $X=328710 $Y=233680
X2758 1 2 291 2 299 1 sky130_fd_sc_hd__clkbuf_16 $T=330280 236640 0 0 $X=330090 $Y=236400
X2759 1 2 293 2 300 1 sky130_fd_sc_hd__clkbuf_16 $T=331660 242080 1 0 $X=331470 $Y=239120
X2760 1 2 96 2 302 1 sky130_fd_sc_hd__clkbuf_16 $T=338100 231200 1 0 $X=337910 $Y=228240
X2761 1 2 322 2 201 1 sky130_fd_sc_hd__clkbuf_16 $T=362940 198560 1 0 $X=362750 $Y=195600
X2762 1 2 341 2 183 1 sky130_fd_sc_hd__clkbuf_16 $T=388240 193120 1 0 $X=388050 $Y=190160
X2763 1 2 344 2 205 1 sky130_fd_sc_hd__clkbuf_16 $T=393760 182240 1 0 $X=393570 $Y=179280
X2764 1 2 347 2 182 1 sky130_fd_sc_hd__clkbuf_16 $T=396980 198560 1 0 $X=396790 $Y=195600
X2765 1 2 352 2 181 1 sky130_fd_sc_hd__clkbuf_16 $T=398820 193120 0 0 $X=398630 $Y=192880
X2766 1 2 357 2 362 1 sky130_fd_sc_hd__clkbuf_16 $T=411240 182240 0 0 $X=411050 $Y=182000
X2767 1 2 407 2 405 1 sky130_fd_sc_hd__clkbuf_16 $T=501860 182240 1 0 $X=501670 $Y=179280
X2768 1 2 357 2 404 1 sky130_fd_sc_hd__clkbuf_16 $T=509220 187680 1 0 $X=509030 $Y=184720
X2769 1 2 417 2 421 1 sky130_fd_sc_hd__clkbuf_16 $T=511060 204000 0 0 $X=510870 $Y=203760
X2770 1 2 418 2 422 1 sky130_fd_sc_hd__clkbuf_16 $T=511060 209440 0 0 $X=510870 $Y=209200
X2771 1 2 419 2 409 1 sky130_fd_sc_hd__clkbuf_16 $T=511520 204000 1 0 $X=511330 $Y=201040
X2772 1 2 766 773 39 ICV_56 $T=113620 225760 1 0 $X=113430 $Y=222800
X2773 1 2 810 780 28 ICV_56 $T=131100 209440 0 0 $X=130910 $Y=209200
X2774 1 2 893 868 44 ICV_56 $T=178020 198560 0 0 $X=177830 $Y=198320
X2775 1 2 922 909 48 ICV_56 $T=192280 198560 1 0 $X=192090 $Y=195600
X2776 1 2 939 170 153 ICV_56 $T=208840 236640 1 0 $X=208650 $Y=233680
X2777 1 2 1122 1100 157 ICV_56 $T=293020 236640 1 0 $X=292830 $Y=233680
X2778 1 2 1333 1297 244 ICV_56 $T=414460 220320 1 0 $X=414270 $Y=217360
X2779 1 2 1384 1389 252 ICV_56 $T=441140 214880 1 0 $X=440950 $Y=211920
X2780 1 2 386 387 238 ICV_56 $T=468280 242080 0 0 $X=468090 $Y=241840
X2781 1 2 1466 1449 238 ICV_56 $T=480240 193120 1 0 $X=480050 $Y=190160
X2782 1 2 1495 1499 285 ICV_56 $T=497260 198560 1 0 $X=497070 $Y=195600
X2783 1 2 1627 1636 271 ICV_56 $T=567180 225760 0 0 $X=566990 $Y=225520
X2784 1 2 1675 1652 251 ICV_56 $T=591100 214880 1 0 $X=590910 $Y=211920
X2785 1 2 1702 1704 271 ICV_56 $T=609500 214880 1 0 $X=609310 $Y=211920
X2786 1 2 1910 509 412 ICV_56 $T=708860 236640 0 0 $X=708670 $Y=236400
X2787 1 2 1943 1938 430 ICV_56 $T=723120 225760 1 0 $X=722930 $Y=222800
X2788 1 2 587 21 609 609 3 40 ICV_58 $T=16100 242080 0 0 $X=15910 $Y=241840
X2789 1 2 589 34 618 618 603 45 ICV_58 $T=20240 220320 1 0 $X=20050 $Y=217360
X2790 1 2 627 36 634 625 619 8 ICV_58 $T=31280 225760 1 0 $X=31090 $Y=222800
X2791 1 2 49 12 642 642 57 28 ICV_58 $T=33120 193120 1 0 $X=32930 $Y=190160
X2792 1 2 653 25 667 667 672 41 ICV_58 $T=46920 236640 0 0 $X=46730 $Y=236400
X2793 1 2 751 13 781 781 757 27 ICV_58 $T=104420 220320 1 0 $X=104230 $Y=217360
X2794 1 2 897 36 949 924 177 28 ICV_58 $T=195960 187680 1 0 $X=195770 $Y=184720
X2795 1 2 1096 182 1113 1111 1091 212 ICV_58 $T=276920 209440 1 0 $X=276730 $Y=206480
X2796 1 2 1092 138 1117 1117 1100 153 ICV_58 $T=280140 242080 1 0 $X=279950 $Y=239120
X2797 1 2 305 288 1221 312 313 271 ICV_58 $T=342700 242080 0 0 $X=342510 $Y=241840
X2798 1 2 1301 288 1309 1310 1311 251 ICV_58 $T=392380 231200 1 0 $X=392190 $Y=228240
X2799 1 2 1508 409 1528 1523 1530 412 ICV_58 $T=501400 225760 1 0 $X=501210 $Y=222800
X2800 1 2 1617 317 1634 1634 1636 330 ICV_58 $T=557520 220320 1 0 $X=557330 $Y=217360
X2801 1 2 463 299 1674 1674 1667 238 ICV_58 $T=581440 198560 1 0 $X=581250 $Y=195600
X2802 1 2 1643 288 1676 1676 1652 255 ICV_58 $T=581440 220320 1 0 $X=581250 $Y=217360
X2803 1 2 1642 317 1677 1673 1653 251 ICV_58 $T=581440 231200 1 0 $X=581250 $Y=228240
X2804 1 2 1686 299 1703 1703 1704 238 ICV_58 $T=595240 214880 0 0 $X=595050 $Y=214640
X2805 1 2 1765 298 1809 1809 1759 285 ICV_58 $T=648140 220320 1 0 $X=647950 $Y=217360
X2806 1 2 508 405 1888 1888 509 413 ICV_58 $T=685860 242080 0 0 $X=685670 $Y=241840
X2807 1 2 587 20 607 607 3 39 ICV_60 $T=18860 231200 0 0 $X=18670 $Y=230960
X2808 1 2 860 12 871 871 868 28 ICV_60 $T=159620 193120 0 0 $X=159430 $Y=192880
X2809 1 2 125 13 896 896 129 27 ICV_60 $T=173420 182240 1 0 $X=173230 $Y=179280
X2810 1 2 911 33 926 926 929 44 ICV_60 $T=187680 209440 0 0 $X=187490 $Y=209200
X2811 1 2 963 205 1010 1010 966 216 ICV_60 $T=230000 204000 1 0 $X=229810 $Y=201040
X2812 1 2 228 181 242 1082 234 212 ICV_60 $T=264500 182240 0 0 $X=264310 $Y=182000
X2813 1 2 1108 199 1130 1130 258 211 ICV_60 $T=289340 193120 0 0 $X=289150 $Y=192880
X2814 1 2 1252 181 1261 1261 1268 198 ICV_60 $T=370300 204000 1 0 $X=370110 $Y=201040
X2815 1 2 1369 267 1399 1399 1389 194 ICV_60 $T=441140 204000 1 0 $X=440950 $Y=201040
X2816 1 2 1391 282 1418 1418 1337 244 ICV_60 $T=449880 225760 1 0 $X=449690 $Y=222800
X2817 1 2 1415 299 1454 1454 1438 238 ICV_60 $T=467820 204000 0 0 $X=467630 $Y=203760
X2818 1 2 1415 286 1458 1458 1438 251 ICV_60 $T=469200 204000 1 0 $X=469010 $Y=201040
X2819 1 2 389 300 1468 1468 393 271 ICV_60 $T=473800 242080 1 0 $X=473610 $Y=239120
X2820 1 2 1474 299 1486 1486 1491 238 ICV_60 $T=483000 204000 0 0 $X=482810 $Y=203760
X2821 1 2 1535 423 1554 1553 1546 414 ICV_60 $T=520260 209440 0 0 $X=520070 $Y=209200
X2822 1 2 1594 405 1629 450 437 429 ICV_60 $T=557520 242080 1 0 $X=557330 $Y=239120
X2823 1 2 463 297 1666 1666 1667 249 ICV_60 $T=581440 193120 1 0 $X=581250 $Y=190160
X2824 1 2 1686 297 1701 1701 1704 249 ICV_60 $T=598460 198560 0 0 $X=598270 $Y=198320
X2825 1 2 481 299 1724 1724 486 238 ICV_60 $T=610880 198560 1 0 $X=610690 $Y=195600
X2826 1 2 1688 286 1731 1731 1713 251 ICV_60 $T=613640 242080 1 0 $X=613450 $Y=239120
X2827 1 2 488 297 1755 1725 486 329 ICV_60 $T=625600 187680 0 0 $X=625410 $Y=187440
X2828 1 2 495 288 1771 1771 500 255 ICV_60 $T=636180 242080 0 0 $X=635990 $Y=241840
X2829 1 2 1727 318 1766 1764 1745 285 ICV_60 $T=636640 214880 0 0 $X=636450 $Y=214640
X2830 1 2 1770 299 1799 1799 1787 238 ICV_60 $T=650900 193120 1 0 $X=650710 $Y=190160
X2831 1 2 67 681 ICV_61 $T=72220 198560 1 0 $X=72030 $Y=195600
X2832 1 2 72 73 ICV_61 $T=86020 236640 0 0 $X=85830 $Y=236400
X2833 1 2 92 750 ICV_61 $T=114080 193120 0 0 $X=113890 $Y=192880
X2834 1 2 118 834 ICV_61 $T=156860 214880 1 0 $X=156670 $Y=211920
X2835 1 2 101 268 ICV_61 $T=318780 182240 1 0 $X=318590 $Y=179280
X2836 1 2 301 309 ICV_61 $T=353280 236640 1 0 $X=353090 $Y=233680
X2837 1 2 169 1255 ICV_61 $T=385020 193120 1 0 $X=384830 $Y=190160
X2838 1 2 346 1297 ICV_61 $T=417220 214880 1 0 $X=417030 $Y=211920
X2839 1 2 340 1368 ICV_61 $T=437000 214880 1 0 $X=436810 $Y=211920
X2840 1 2 301 1546 ICV_61 $T=534980 204000 0 0 $X=534790 $Y=203760
X2841 1 2 378 437 ICV_61 $T=535440 242080 0 0 $X=535250 $Y=241840
X2842 1 2 439 1581 ICV_61 $T=546480 182240 0 0 $X=546290 $Y=182000
X2843 1 2 390 1612 ICV_61 $T=553380 225760 1 0 $X=553190 $Y=222800
X2844 1 2 441 443 ICV_61 $T=553840 182240 1 0 $X=553650 $Y=179280
X2845 1 2 462 477 ICV_61 $T=602600 242080 0 0 $X=602410 $Y=241840
X2846 1 2 380 1856 ICV_61 $T=686780 225760 0 0 $X=686590 $Y=225520
X2847 1 2 622 603 48 ICV_62 $T=34040 214880 0 0 $X=33850 $Y=214640
X2848 1 2 651 619 40 ICV_62 $T=45540 231200 0 0 $X=45350 $Y=230960
X2849 1 2 668 672 66 ICV_62 $T=57500 242080 1 0 $X=57310 $Y=239120
X2850 1 2 68 69 46 ICV_62 $T=62100 242080 1 0 $X=61910 $Y=239120
X2851 1 2 814 808 40 ICV_62 $T=133860 242080 1 0 $X=133670 $Y=239120
X2852 1 2 865 824 8 ICV_62 $T=165140 236640 0 0 $X=164950 $Y=236400
X2853 1 2 1031 1046 211 ICV_62 $T=254380 225760 1 0 $X=254190 $Y=222800
X2854 1 2 1086 1087 196 ICV_62 $T=273240 187680 1 0 $X=273050 $Y=184720
X2855 1 2 1094 247 152 ICV_62 $T=281520 242080 0 0 $X=281330 $Y=241840
X2856 1 2 1113 1091 185 ICV_62 $T=291640 209440 1 0 $X=291450 $Y=206480
X2857 1 2 1196 1184 261 ICV_62 $T=339940 220320 1 0 $X=339750 $Y=217360
X2858 1 2 1241 309 329 ICV_62 $T=365700 242080 0 0 $X=365510 $Y=241840
X2859 1 2 1246 1239 231 ICV_62 $T=370760 220320 0 0 $X=370570 $Y=220080
X2860 1 2 1286 1268 196 ICV_62 $T=389620 193120 0 0 $X=389430 $Y=192880
X2861 1 2 1287 1248 285 ICV_62 $T=393760 225760 1 0 $X=393570 $Y=222800
X2862 1 2 1341 1327 231 ICV_62 $T=417680 193120 0 0 $X=417490 $Y=192880
X2863 1 2 1403 370 330 ICV_62 $T=454940 225760 0 0 $X=454750 $Y=225520
X2864 1 2 1416 1337 252 ICV_62 $T=463220 204000 0 0 $X=463030 $Y=203760
X2865 1 2 1444 1422 271 ICV_62 $T=469200 242080 1 0 $X=469010 $Y=239120
X2866 1 2 1453 1449 329 ICV_62 $T=472420 182240 0 0 $X=472230 $Y=182000
X2867 1 2 1482 393 255 ICV_62 $T=488060 242080 0 0 $X=487870 $Y=241840
X2868 1 2 1484 392 194 ICV_62 $T=497260 182240 1 0 $X=497070 $Y=179280
X2869 1 2 1502 1499 329 ICV_62 $T=501400 187680 0 0 $X=501210 $Y=187440
X2870 1 2 1570 1568 413 ICV_62 $T=534060 231200 0 0 $X=533870 $Y=230960
X2871 1 2 440 437 430 ICV_62 $T=547400 242080 0 0 $X=547210 $Y=241840
X2872 1 2 1603 1605 330 ICV_62 $T=556600 198560 0 0 $X=556410 $Y=198320
X2873 1 2 1658 1653 249 ICV_62 $T=581440 236640 1 0 $X=581250 $Y=233680
X2874 1 2 1664 1667 255 ICV_62 $T=587880 187680 1 0 $X=587690 $Y=184720
X2875 1 2 1707 1699 285 ICV_62 $T=609500 225760 1 0 $X=609310 $Y=222800
X2876 1 2 1716 1699 238 ICV_62 $T=615480 225760 1 0 $X=615290 $Y=222800
X2877 1 2 1735 1713 238 ICV_62 $T=623300 242080 0 0 $X=623110 $Y=241840
X2878 1 2 1789 1759 255 ICV_62 $T=651360 214880 0 0 $X=651170 $Y=214640
X2879 1 2 1794 501 424 ICV_62 $T=653660 182240 0 0 $X=653470 $Y=182000
X2880 1 2 1822 1818 415 ICV_62 $T=666540 220320 1 0 $X=666350 $Y=217360
X2881 1 2 1905 1844 414 ICV_62 $T=707480 225760 0 0 $X=707290 $Y=225520
X2882 1 2 612 15 44 ICV_63 $T=28060 193120 1 0 $X=27870 $Y=190160
X2883 1 2 648 640 45 ICV_63 $T=43700 209440 0 0 $X=43510 $Y=209200
X2884 1 2 687 691 19 ICV_63 $T=67620 209440 0 0 $X=67430 $Y=209200
X2885 1 2 717 73 39 ICV_63 $T=80960 231200 0 0 $X=80770 $Y=230960
X2886 1 2 741 87 41 ICV_63 $T=98440 242080 1 0 $X=98250 $Y=239120
X2887 1 2 770 750 50 ICV_63 $T=110860 193120 1 0 $X=110670 $Y=190160
X2888 1 2 799 757 45 ICV_63 $T=124660 209440 0 0 $X=124470 $Y=209200
X2889 1 2 850 834 44 ICV_63 $T=151800 214880 1 0 $X=151610 $Y=211920
X2890 1 2 854 119 19 ICV_63 $T=155020 198560 1 0 $X=154830 $Y=195600
X2891 1 2 214 217 153 ICV_63 $T=238280 242080 0 0 $X=238090 $Y=241840
X2892 1 2 1038 1046 212 ICV_63 $T=250700 209440 0 0 $X=250510 $Y=209200
X2893 1 2 1057 1055 155 ICV_63 $T=258520 225760 0 0 $X=258330 $Y=225520
X2894 1 2 1099 1100 135 ICV_63 $T=280140 225760 1 0 $X=279950 $Y=222800
X2895 1 2 1139 1138 153 ICV_63 $T=300840 242080 1 0 $X=300650 $Y=239120
X2896 1 2 1282 1280 244 ICV_63 $T=385480 214880 0 0 $X=385290 $Y=214640
X2897 1 2 1357 1368 261 ICV_63 $T=426880 204000 0 0 $X=426690 $Y=203760
X2898 1 2 371 364 254 ICV_63 $T=441140 182240 1 0 $X=440950 $Y=179280
X2899 1 2 483 484 285 ICV_63 $T=615480 236640 0 0 $X=615290 $Y=236400
X2900 1 2 1738 1739 330 ICV_63 $T=623300 231200 0 0 $X=623110 $Y=230960
X2901 1 2 1853 1826 412 ICV_63 $T=679420 198560 0 0 $X=679230 $Y=198320
X2902 1 2 1959 1901 413 ICV_63 $T=730020 193120 0 0 $X=729830 $Y=192880
X2903 1 2 22 26 30 ICV_65 $T=20240 182240 1 0 $X=20050 $Y=179280
X2904 1 2 42 43 47 ICV_65 $T=30820 242080 0 0 $X=30630 $Y=241840
X2905 1 2 64 43 675 ICV_65 $T=58880 242080 0 0 $X=58690 $Y=241840
X2906 1 2 77 26 704 ICV_65 $T=73140 214880 1 0 $X=72950 $Y=211920
X2907 1 2 112 26 113 ICV_65 $T=132480 182240 1 0 $X=132290 $Y=179280
X2908 1 2 123 26 859 ICV_65 $T=157320 209440 1 0 $X=157130 $Y=206480
X2909 1 2 133 26 134 ICV_65 $T=170660 182240 1 0 $X=170470 $Y=179280
X2910 1 2 64 128 948 ICV_65 $T=202400 236640 0 0 $X=202210 $Y=236400
X2911 1 2 91 178 1090 ICV_65 $T=273240 198560 0 0 $X=273050 $Y=198320
X2912 1 2 115 128 1131 ICV_65 $T=293940 242080 0 0 $X=293750 $Y=241840
X2913 1 2 114 178 1180 ICV_65 $T=328900 204000 1 0 $X=328710 $Y=201040
X2914 1 2 315 302 1232 ICV_65 $T=356960 209440 1 0 $X=356770 $Y=206480
X2915 1 2 334 302 1260 ICV_65 $T=374440 220320 1 0 $X=374250 $Y=217360
X2916 1 2 340 302 1332 ICV_65 $T=412620 214880 0 0 $X=412430 $Y=214640
X2917 1 2 367 302 1379 ICV_65 $T=432860 193120 1 0 $X=432670 $Y=190160
X2918 1 2 439 308 1572 ICV_65 $T=540040 182240 1 0 $X=539850 $Y=179280
X2919 1 2 462 308 1659 ICV_65 $T=578220 242080 1 0 $X=578030 $Y=239120
X2920 1 2 385 398 1793 ICV_65 $T=651360 231200 0 0 $X=651170 $Y=230960
X2921 1 2 469 398 504 ICV_65 $T=662860 242080 0 0 $X=662670 $Y=241840
X2922 1 2 446 398 1829 ICV_65 $T=667920 182240 0 0 $X=667730 $Y=182000
X2923 1 2 462 398 1864 ICV_65 $T=683100 242080 0 0 $X=682910 $Y=241840
X2924 1 2 9 13 600 ICV_66 $T=12420 187680 1 0 $X=12230 $Y=184720
X2925 1 2 588 10 602 ICV_66 $T=12420 204000 1 0 $X=12230 $Y=201040
X2926 1 2 875 146 914 ICV_66 $T=180780 236640 1 0 $X=180590 $Y=233680
X2927 1 2 127 194 941 ICV_66 $T=222640 220320 0 0 $X=222450 $Y=220080
X2928 1 2 1066 199 1083 ICV_66 $T=264960 198560 1 0 $X=264770 $Y=195600
X2929 1 2 264 130 270 ICV_66 $T=306820 242080 0 0 $X=306630 $Y=241840
X2930 1 2 1197 201 1192 ICV_66 $T=349140 187680 1 0 $X=348950 $Y=184720
X2931 1 2 1237 183 1250 ICV_66 $T=362940 182240 0 0 $X=362750 $Y=182000
X2932 1 2 1262 279 1278 ICV_66 $T=377200 220320 1 0 $X=377010 $Y=217360
X2933 1 2 1342 282 1358 ICV_66 $T=419060 220320 0 0 $X=418870 $Y=220080
X2934 1 2 361 288 1361 ICV_66 $T=419060 242080 0 0 $X=418870 $Y=241840
X2935 1 2 1456 299 1473 ICV_66 $T=475180 231200 0 0 $X=474990 $Y=230960
X2936 1 2 1866 404 1908 ICV_66 $T=699660 198560 0 0 $X=699470 $Y=198320
X2937 1 2 1923 422 515 ICV_66 $T=713920 236640 1 0 $X=713730 $Y=233680
X2938 1 2 1917 409 1964 ICV_66 $T=727720 225760 0 0 $X=727530 $Y=225520
X2939 1 2 1923 409 1945 ICV_66 $T=727720 231200 0 0 $X=727530 $Y=230960
X2940 1 2 514 409 522 ICV_66 $T=727720 242080 0 0 $X=727530 $Y=241840
X2941 1 2 451 452 2 249 1 sky130_fd_sc_hd__ebufn_4 $T=565340 193120 1 0 $X=565150 $Y=190160
X2942 1 2 451 452 2 255 1 sky130_fd_sc_hd__ebufn_4 $T=569020 187680 1 0 $X=568830 $Y=184720
X2943 1 2 451 452 2 285 1 sky130_fd_sc_hd__ebufn_4 $T=569480 187680 0 0 $X=569290 $Y=187440
X2944 1 2 451 452 2 238 1 sky130_fd_sc_hd__ebufn_4 $T=570400 193120 0 0 $X=570210 $Y=192880
X2945 1 2 451 452 2 271 1 sky130_fd_sc_hd__ebufn_4 $T=571320 193120 1 0 $X=571130 $Y=190160
X2946 1 2 451 452 2 330 1 sky130_fd_sc_hd__ebufn_4 $T=572240 182240 0 0 $X=572050 $Y=182000
X2947 1 2 451 452 2 329 1 sky130_fd_sc_hd__ebufn_4 $T=575000 187680 1 0 $X=574810 $Y=184720
X2948 1 2 673 2 65 1 sky130_fd_sc_hd__clkbuf_4 $T=59800 220320 1 0 $X=59610 $Y=217360
X2949 1 2 729 2 85 1 sky130_fd_sc_hd__clkbuf_4 $T=87860 220320 1 0 $X=87670 $Y=217360
X2950 1 2 898 2 144 1 sky130_fd_sc_hd__clkbuf_4 $T=180320 220320 1 0 $X=180130 $Y=217360
X2951 1 2 945 2 174 1 sky130_fd_sc_hd__clkbuf_4 $T=203780 220320 0 0 $X=203590 $Y=220080
X2952 1 2 977 2 190 1 sky130_fd_sc_hd__clkbuf_4 $T=220340 214880 0 0 $X=220150 $Y=214640
X2953 1 2 1000 2 203 1 sky130_fd_sc_hd__clkbuf_4 $T=229540 220320 1 0 $X=229350 $Y=217360
X2954 1 2 626 34 648 ICV_69 $T=44620 204000 0 0 $X=44430 $Y=203760
X2955 1 2 734 34 701 ICV_69 $T=90620 220320 1 0 $X=90430 $Y=217360
X2956 1 2 89 33 762 ICV_69 $T=102120 187680 0 0 $X=101930 $Y=187440
X2957 1 2 104 12 809 ICV_69 $T=122360 187680 1 0 $X=122170 $Y=184720
X2958 1 2 836 20 846 ICV_69 $T=143060 236640 1 0 $X=142870 $Y=233680
X2959 1 2 866 10 889 ICV_69 $T=168820 209440 1 0 $X=168630 $Y=206480
X2960 1 2 159 148 932 ICV_69 $T=192740 231200 0 0 $X=192550 $Y=230960
X2961 1 2 127 41 965 ICV_69 $T=207000 231200 1 0 $X=206810 $Y=228240
X2962 1 2 955 146 973 ICV_69 $T=212520 231200 0 0 $X=212330 $Y=230960
X2963 1 2 1062 182 1072 ICV_69 $T=261740 214880 1 0 $X=261550 $Y=211920
X2964 1 2 1062 201 1076 ICV_69 $T=262660 209440 1 0 $X=262470 $Y=206480
X2965 1 2 1116 148 1142 ICV_69 $T=297160 231200 0 0 $X=296970 $Y=230960
X2966 1 2 1173 284 1194 ICV_69 $T=332580 214880 1 0 $X=332390 $Y=211920
X2967 1 2 339 201 1328 ICV_69 $T=402960 182240 1 0 $X=402770 $Y=179280
X2968 1 2 1308 278 1326 ICV_69 $T=403420 198560 0 0 $X=403230 $Y=198320
X2969 1 2 1342 284 1365 ICV_69 $T=420440 214880 1 0 $X=420250 $Y=211920
X2970 1 2 1481 297 1494 ICV_69 $T=487140 193120 1 0 $X=486950 $Y=190160
X2971 1 2 1476 296 1507 ICV_69 $T=493580 214880 0 0 $X=493390 $Y=214640
X2972 1 2 1508 403 1523 ICV_69 $T=501400 220320 0 0 $X=501210 $Y=220080
X2973 1 2 1535 406 1571 ICV_69 $T=528080 214880 1 0 $X=527890 $Y=211920
X2974 1 2 1598 317 449 ICV_69 $T=557520 182240 0 0 $X=557330 $Y=182000
X2975 1 2 1714 317 1728 ICV_69 $T=613640 204000 0 0 $X=613450 $Y=203760
X2976 1 2 1714 297 1730 ICV_69 $T=613640 209440 0 0 $X=613450 $Y=209200
X2977 1 2 1743 299 1761 ICV_69 $T=627900 231200 1 0 $X=627710 $Y=228240
X2978 1 2 1861 403 1875 ICV_69 $T=684020 225760 1 0 $X=683830 $Y=222800
X2979 1 2 883 884 139 140 892 141 2 898 1 sky130_fd_sc_hd__mux4_1 $T=172500 225760 1 0 $X=172310 $Y=222800
X2980 1 2 894 890 139 150 906 141 2 729 1 sky130_fd_sc_hd__mux4_1 $T=178940 220320 0 0 $X=178750 $Y=220080
X2981 1 2 912 904 139 161 925 141 2 168 1 sky130_fd_sc_hd__mux4_1 $T=188600 225760 1 0 $X=188410 $Y=222800
X2982 1 2 931 886 139 171 941 141 2 945 1 sky130_fd_sc_hd__mux4_1 $T=197340 231200 1 0 $X=197150 $Y=228240
X2983 1 2 930 921 139 172 943 141 2 673 1 sky130_fd_sc_hd__mux4_1 $T=198260 225760 1 0 $X=198070 $Y=222800
X2984 1 2 968 969 139 191 981 141 2 977 1 sky130_fd_sc_hd__mux4_1 $T=216660 220320 1 0 $X=216470 $Y=217360
X2985 1 2 961 965 139 192 982 141 2 197 1 sky130_fd_sc_hd__mux4_1 $T=216660 225760 1 0 $X=216470 $Y=222800
X2986 1 2 984 971 139 204 1001 141 2 1000 1 sky130_fd_sc_hd__mux4_1 $T=226320 225760 1 0 $X=226130 $Y=222800
X2987 1 2 202 206 139 209 1008 141 2 213 1 sky130_fd_sc_hd__mux4_1 $T=230460 220320 0 0 $X=230270 $Y=220080
X2988 1 2 207 208 139 210 1019 141 2 220 1 sky130_fd_sc_hd__mux4_1 $T=232300 220320 1 0 $X=232110 $Y=217360
X2989 1 2 1029 226 139 229 1037 141 2 233 1 sky130_fd_sc_hd__mux4_1 $T=244720 225760 1 0 $X=244530 $Y=222800
X2990 1 2 1054 236 139 239 1065 141 2 241 1 sky130_fd_sc_hd__mux4_1 $T=258980 225760 1 0 $X=258790 $Y=222800
X2991 1 2 1067 248 139 253 1118 141 2 257 1 sky130_fd_sc_hd__mux4_1 $T=285200 225760 1 0 $X=285010 $Y=222800
X2992 1 2 1098 265 139 269 1157 141 2 273 1 sky130_fd_sc_hd__mux4_1 $T=307280 231200 1 0 $X=307090 $Y=228240
.ENDS
***************************************
.SUBCKT ICV_80 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=26
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=7360 0 0 0 $X=7170 $Y=-240
X1 1 2 3 4 2 5 1 sky130_fd_sc_hd__dfxtp_1 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_81 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=460 0 0 0 $X=270 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_82
** N=2 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_sc_hd__and3b_4 VNB VPB B C A_N VPWR X VGND
** N=81 EP=8 IP=0 FDC=16
*.SEEDPROM
M0 11 9 10 VNB nshort L=0.15 W=0.65 AD=0.121875 AS=0.19825 PD=1.025 PS=1.91 NRD=24.456 NRS=0 m=1 r=4.33333 sa=75000.2 sb=75003.4 a=0.0975 p=1.6 mult=1 $X=610 $Y=235 $D=9
M1 12 B 11 VNB nshort L=0.15 W=0.65 AD=0.07475 AS=0.121875 PD=0.88 PS=1.025 NRD=11.076 NRS=24.456 m=1 r=4.33333 sa=75000.8 sb=75002.8 a=0.0975 p=1.6 mult=1 $X=1135 $Y=235 $D=8
M2 VGND C 12 VNB nshort L=0.15 W=0.65 AD=0.138125 AS=0.07475 PD=1.075 PS=0.88 NRD=25.836 NRS=11.076 m=1 r=4.33333 sa=75001.1 sb=75002.4 a=0.0975 p=1.6 mult=1 $X=1515 $Y=235 $D=9
M3 X 10 VGND VNB nshort L=0.15 W=0.65 AD=0.091 AS=0.138125 PD=0.93 PS=1.075 NRD=0 NRS=0.912 m=1 r=4.33333 sa=75001.7 sb=75001.9 a=0.0975 p=1.6 mult=1 $X=2090 $Y=235 $D=9
M4 VGND 10 X VNB nshort L=0.15 W=0.65 AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 m=1 r=4.33333 sa=75002.1 sb=75001.4 a=0.0975 p=1.6 mult=1 $X=2520 $Y=235 $D=9
M5 X 10 VGND VNB nshort L=0.15 W=0.65 AD=0.091 AS=0.091 PD=0.93 PS=0.93 NRD=0 NRS=0 m=1 r=4.33333 sa=75002.6 sb=75001 a=0.0975 p=1.6 mult=1 $X=2950 $Y=235 $D=9
M6 VGND 10 X VNB nshort L=0.15 W=0.65 AD=0.131671 AS=0.091 PD=1.2271 PS=0.93 NRD=0 NRS=0 m=1 r=4.33333 sa=75003 sb=75000.6 a=0.0975 p=1.6 mult=1 $X=3380 $Y=235 $D=9
M7 9 A_N VGND VNB nshort L=0.15 W=0.42 AD=0.1491 AS=0.0850794 PD=1.55 PS=0.792897 NRD=19.992 NRS=42.156 m=1 r=2.8 sa=75003.5 sb=75000.3 a=0.063 p=1.14 mult=1 $X=3890 $Y=465 $D=9
M8 VPWR 9 10 VPB phighvt L=0.15 W=1 AD=0.1875 AS=0.33 PD=1.375 PS=2.66 NRD=12.7853 NRS=8.8453 m=1 r=6.66667 sa=75000.3 sb=75003.2 a=0.15 p=2.3 mult=1 $X=610 $Y=1485 $D=89
M9 10 B VPWR VPB phighvt L=0.15 W=1 AD=0.15 AS=0.1875 PD=1.3 PS=1.375 NRD=3.9203 NRS=5.8903 m=1 r=6.66667 sa=75000.8 sb=75002.7 a=0.15 p=2.3 mult=1 $X=1135 $Y=1485 $D=89
M10 VPWR C 10 VPB phighvt L=0.15 W=1 AD=0.1775 AS=0.15 PD=1.355 PS=1.3 NRD=6.8753 NRS=0 m=1 r=6.66667 sa=75001.2 sb=75002.2 a=0.15 p=2.3 mult=1 $X=1585 $Y=1485 $D=89
M11 X 10 VPWR VPB phighvt L=0.15 W=1 AD=0.145 AS=0.1775 PD=1.29 PS=1.355 NRD=1.9503 NRS=7.8603 m=1 r=6.66667 sa=75001.7 sb=75001.7 a=0.15 p=2.3 mult=1 $X=2090 $Y=1485 $D=89
M12 VPWR 10 X VPB phighvt L=0.15 W=1 AD=0.135 AS=0.145 PD=1.27 PS=1.29 NRD=0 NRS=0 m=1 r=6.66667 sa=75002.2 sb=75001.3 a=0.15 p=2.3 mult=1 $X=2530 $Y=1485 $D=89
M13 X 10 VPWR VPB phighvt L=0.15 W=1 AD=0.14 AS=0.135 PD=1.28 PS=1.27 NRD=0 NRS=0 m=1 r=6.66667 sa=75002.6 sb=75000.9 a=0.15 p=2.3 mult=1 $X=2950 $Y=1485 $D=89
M14 VPWR 10 X VPB phighvt L=0.15 W=1 AD=0.222887 AS=0.14 PD=1.91549 PS=1.28 NRD=0 NRS=0 m=1 r=6.66667 sa=75003 sb=75000.4 a=0.15 p=2.3 mult=1 $X=3380 $Y=1485 $D=89
M15 9 A_N VPWR VPB phighvt L=0.15 W=0.42 AD=0.1197 AS=0.0936127 PD=1.41 PS=0.804507 NRD=0 NRS=78.7409 m=1 r=2.8 sa=75003.5 sb=75000.2 a=0.063 p=1.14 mult=1 $X=3890 $Y=1725 $D=89
.ENDS
***************************************
.SUBCKT ICV_83 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380
+ 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400
+ 401 402 403 404 405 406 407 408 409 410 411 412 413 414 415 416 417 418 419 420
+ 421 422 423 424 425 426 427 428 429 430 431 432 433 434 435 436 437 438 439 440
+ 441 442 443 444 445 446 447 448 449 450 451 452 453 454 455 456 457 458 459 460
+ 461 462 463 464 465 466 467 468 469 470 471 472 473 474 475 476 477 478 479 480
+ 481 482 483 484 485 486 487 488 489 490 491 492 493 494 495 496 497 498 499 500
+ 501 502 503 504 505 506 507 508 509 510 511 512 513 514 515 516 517 518 519 520
+ 521 522 523 524 525 526 527 528 529 530 531 532 533 534 535 536 537 538 539 540
+ 541 542 543 544 545 546 547 548 549 550 551 552
** N=1978 EP=552 IP=16760 FDC=48295
*.SEEDPROM
X0 1 2 Dpar a=2090.95 p=1484.94 m=1 $[nwdiode] $X=5330 $Y=118265 $D=191
X1 1 2 Dpar a=2091.28 p=1484.54 m=1 $[nwdiode] $X=5330 $Y=123705 $D=191
X2 1 2 Dpar a=2090.63 p=1485.34 m=1 $[nwdiode] $X=5330 $Y=129145 $D=191
X3 1 2 Dpar a=2090.63 p=1485.34 m=1 $[nwdiode] $X=5330 $Y=134585 $D=191
X4 1 2 Dpar a=2090.95 p=1484.94 m=1 $[nwdiode] $X=5330 $Y=140025 $D=191
X5 1 2 Dpar a=2091.12 p=1484.74 m=1 $[nwdiode] $X=5330 $Y=145465 $D=191
X6 1 2 Dpar a=2090.55 p=1485.44 m=1 $[nwdiode] $X=5330 $Y=150905 $D=191
X7 1 2 Dpar a=2091.28 p=1484.54 m=1 $[nwdiode] $X=5330 $Y=156345 $D=191
X8 1 2 Dpar a=2090.63 p=1485.34 m=1 $[nwdiode] $X=5330 $Y=161785 $D=191
X9 1 2 Dpar a=2090.71 p=1485.24 m=1 $[nwdiode] $X=5330 $Y=167225 $D=191
X10 1 2 Dpar a=2090.95 p=1484.94 m=1 $[nwdiode] $X=5330 $Y=172665 $D=191
X11 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=16100 138720 0 0 $X=15910 $Y=138480
X12 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=18400 176800 1 0 $X=18210 $Y=173840
X13 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=38180 122400 1 0 $X=37990 $Y=119440
X14 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=42320 133280 1 0 $X=42130 $Y=130320
X15 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=84180 122400 0 0 $X=83990 $Y=122160
X16 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=102580 122400 1 0 $X=102390 $Y=119440
X17 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=116380 116960 0 0 $X=116190 $Y=116720
X18 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=116380 122400 0 0 $X=116190 $Y=122160
X19 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=118220 138720 0 0 $X=118030 $Y=138480
X20 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=130640 171360 1 0 $X=130450 $Y=168400
X21 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=131100 127840 0 0 $X=130910 $Y=127600
X22 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=145820 176800 1 0 $X=145630 $Y=173840
X23 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=146280 116960 0 0 $X=146090 $Y=116720
X24 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=160540 116960 1 0 $X=160350 $Y=114000
X25 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=160540 133280 1 0 $X=160350 $Y=130320
X26 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=172500 116960 0 0 $X=172310 $Y=116720
X27 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=175720 133280 0 0 $X=175530 $Y=133040
X28 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=198260 116960 1 0 $X=198070 $Y=114000
X29 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=202400 149600 0 0 $X=202210 $Y=149360
X30 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=202400 155040 0 0 $X=202210 $Y=154800
X31 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=208840 160480 1 0 $X=208650 $Y=157520
X32 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=216660 116960 1 0 $X=216470 $Y=114000
X33 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=224020 149600 0 0 $X=223830 $Y=149360
X34 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=242880 127840 1 0 $X=242690 $Y=124880
X35 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=244720 160480 1 0 $X=244530 $Y=157520
X36 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=252540 155040 0 0 $X=252350 $Y=154800
X37 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=253920 116960 1 0 $X=253730 $Y=114000
X38 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=257600 165920 1 0 $X=257410 $Y=162960
X39 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=262660 122400 0 0 $X=262470 $Y=122160
X40 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=272780 171360 1 0 $X=272590 $Y=168400
X41 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=284740 176800 1 0 $X=284550 $Y=173840
X42 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=290260 155040 0 0 $X=290070 $Y=154800
X43 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=291180 138720 0 0 $X=290990 $Y=138480
X44 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=308660 165920 1 0 $X=308470 $Y=162960
X45 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=312340 133280 1 0 $X=312150 $Y=130320
X46 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=314640 133280 0 0 $X=314450 $Y=133040
X47 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=318320 149600 0 0 $X=318130 $Y=149360
X48 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=327060 176800 1 0 $X=326870 $Y=173840
X49 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=342700 155040 0 0 $X=342510 $Y=154800
X50 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=344540 144160 1 0 $X=344350 $Y=141200
X51 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=350980 133280 1 0 $X=350790 $Y=130320
X52 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=361100 176800 1 0 $X=360910 $Y=173840
X53 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=365700 160480 1 0 $X=365510 $Y=157520
X54 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=368920 133280 0 0 $X=368730 $Y=133040
X55 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=383180 138720 1 0 $X=382990 $Y=135760
X56 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=385020 133280 1 0 $X=384830 $Y=130320
X57 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=397440 116960 1 0 $X=397250 $Y=114000
X58 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=402960 176800 0 0 $X=402770 $Y=176560
X59 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=417220 155040 0 0 $X=417030 $Y=154800
X60 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=425040 165920 0 0 $X=424850 $Y=165680
X61 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=439300 149600 1 0 $X=439110 $Y=146640
X62 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=448960 127840 1 0 $X=448770 $Y=124880
X63 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=456780 138720 1 0 $X=456590 $Y=135760
X64 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=477020 171360 0 0 $X=476830 $Y=171120
X65 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=481160 122400 1 0 $X=480970 $Y=119440
X66 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=485760 127840 1 0 $X=485570 $Y=124880
X67 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=493120 149600 1 0 $X=492930 $Y=146640
X68 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=495420 127840 1 0 $X=495230 $Y=124880
X69 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=498180 160480 0 0 $X=497990 $Y=160240
X70 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=509220 160480 0 0 $X=509030 $Y=160240
X71 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=535900 144160 1 0 $X=535710 $Y=141200
X72 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=544640 138720 0 0 $X=544450 $Y=138480
X73 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=553380 165920 1 0 $X=553190 $Y=162960
X74 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=558900 138720 0 0 $X=558710 $Y=138480
X75 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=561200 171360 0 0 $X=561010 $Y=171120
X76 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=565340 155040 0 0 $X=565150 $Y=154800
X77 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=581440 165920 1 0 $X=581250 $Y=162960
X78 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=581440 176800 1 0 $X=581250 $Y=173840
X79 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=595240 144160 0 0 $X=595050 $Y=143920
X80 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=614100 138720 1 0 $X=613910 $Y=135760
X81 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=615940 138720 0 0 $X=615750 $Y=138480
X82 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=620080 138720 1 0 $X=619890 $Y=135760
X83 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=621000 149600 1 0 $X=620810 $Y=146640
X84 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=627440 133280 0 0 $X=627250 $Y=133040
X85 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=627440 160480 0 0 $X=627250 $Y=160240
X86 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=628820 116960 0 0 $X=628630 $Y=116720
X87 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=657340 127840 1 0 $X=657150 $Y=124880
X88 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=658720 165920 0 0 $X=658530 $Y=165680
X89 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=659640 176800 1 0 $X=659450 $Y=173840
X90 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=680340 171360 1 0 $X=680150 $Y=168400
X91 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=690920 138720 0 0 $X=690730 $Y=138480
X92 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=693680 116960 1 0 $X=693490 $Y=114000
X93 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=693680 127840 1 0 $X=693490 $Y=124880
X94 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=695060 133280 0 0 $X=694870 $Y=133040
X95 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=703340 176800 0 0 $X=703150 $Y=176560
X96 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=712080 116960 1 0 $X=711890 $Y=114000
X97 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=719900 116960 1 0 $X=719710 $Y=114000
X98 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=721740 122400 1 0 $X=721550 $Y=119440
X99 1 2 ICV_1 $T=744280 116960 0 180 $X=742710 $Y=114000
X100 1 2 ICV_1 $T=744280 122400 0 180 $X=742710 $Y=119440
X101 1 2 ICV_1 $T=744280 127840 0 180 $X=742710 $Y=124880
X102 1 2 ICV_1 $T=744280 176800 0 180 $X=742710 $Y=173840
X103 1 2 ICV_2 $T=5520 116960 1 0 $X=5330 $Y=114000
X104 1 2 ICV_2 $T=5520 127840 1 0 $X=5330 $Y=124880
X105 1 2 ICV_2 $T=5520 138720 1 0 $X=5330 $Y=135760
X106 1 2 ICV_2 $T=5520 149600 1 0 $X=5330 $Y=146640
X107 1 2 ICV_2 $T=5520 160480 1 0 $X=5330 $Y=157520
X108 1 2 ICV_2 $T=5520 171360 1 0 $X=5330 $Y=168400
X109 1 2 ICV_2 $T=744280 133280 0 180 $X=742710 $Y=130320
X110 1 2 ICV_2 $T=744280 144160 0 180 $X=742710 $Y=141200
X111 1 2 ICV_2 $T=744280 155040 0 180 $X=742710 $Y=152080
X112 1 2 ICV_2 $T=744280 165920 0 180 $X=742710 $Y=162960
X284 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=15640 116960 1 0 $X=15450 $Y=114000
X285 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=25300 176800 0 0 $X=25110 $Y=176560
X286 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=59800 155040 0 0 $X=59610 $Y=154800
X287 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=79580 155040 0 0 $X=79390 $Y=154800
X288 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=102120 127840 1 0 $X=101930 $Y=124880
X289 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=104420 155040 1 0 $X=104230 $Y=152080
X290 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=111780 144160 0 0 $X=111590 $Y=143920
X291 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=115920 127840 0 0 $X=115730 $Y=127600
X292 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=115920 133280 0 0 $X=115730 $Y=133040
X293 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=118220 160480 0 0 $X=118030 $Y=160240
X294 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=137540 155040 0 0 $X=137350 $Y=154800
X295 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=143980 149600 0 0 $X=143790 $Y=149360
X296 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=150420 165920 0 0 $X=150230 $Y=165680
X297 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=172040 144160 0 0 $X=171850 $Y=143920
X298 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=172040 149600 0 0 $X=171850 $Y=149360
X299 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=202400 116960 0 0 $X=202210 $Y=116720
X300 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=213900 133280 0 0 $X=213710 $Y=133040
X301 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=222180 155040 0 0 $X=221990 $Y=154800
X302 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=242420 149600 0 0 $X=242230 $Y=149360
X303 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=298540 138720 1 0 $X=298350 $Y=135760
X304 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=312340 127840 0 0 $X=312150 $Y=127600
X305 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=318320 149600 1 0 $X=318130 $Y=146640
X306 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=320160 171360 1 0 $X=319970 $Y=168400
X307 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=322460 122400 1 0 $X=322270 $Y=119440
X308 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=326600 149600 1 0 $X=326410 $Y=146640
X309 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=354660 160480 1 0 $X=354470 $Y=157520
X310 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=367540 155040 1 0 $X=367350 $Y=152080
X311 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=378580 165920 0 0 $X=378390 $Y=165680
X312 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=410780 160480 1 0 $X=410590 $Y=157520
X313 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=413080 133280 1 0 $X=412890 $Y=130320
X314 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=424580 127840 0 0 $X=424390 $Y=127600
X315 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=434700 155040 1 0 $X=434510 $Y=152080
X316 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=452640 122400 0 0 $X=452450 $Y=122160
X317 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=466900 127840 0 0 $X=466710 $Y=127600
X318 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=479320 171360 1 0 $X=479130 $Y=168400
X319 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=480700 127840 0 0 $X=480510 $Y=127600
X320 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=507840 171360 1 0 $X=507650 $Y=168400
X321 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=512900 116960 1 0 $X=512710 $Y=114000
X322 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=525320 165920 1 0 $X=525130 $Y=162960
X323 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=539120 122400 1 0 $X=538930 $Y=119440
X324 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=564880 176800 0 0 $X=564690 $Y=176560
X325 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=574540 176800 0 0 $X=574350 $Y=176560
X326 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=575000 138720 0 0 $X=574810 $Y=138480
X327 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=577760 133280 0 0 $X=577570 $Y=133040
X328 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=577760 155040 0 0 $X=577570 $Y=154800
X329 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=592940 127840 0 0 $X=592750 $Y=127600
X330 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=614560 160480 0 0 $X=614370 $Y=160240
X331 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=623300 165920 0 0 $X=623110 $Y=165680
X332 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=644920 165920 1 0 $X=644730 $Y=162960
X333 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=649060 160480 0 0 $X=648870 $Y=160240
X334 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=662400 138720 0 0 $X=662210 $Y=138480
X335 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=690920 127840 0 0 $X=690730 $Y=127600
X336 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=697820 176800 1 0 $X=697630 $Y=173840
X337 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=707480 122400 0 0 $X=707290 $Y=122160
X338 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=713000 165920 1 0 $X=712810 $Y=162960
X339 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=735540 176800 0 0 $X=735350 $Y=176560
X340 1 2 ICV_3 $T=12420 176800 0 0 $X=12230 $Y=176560
X341 1 2 ICV_3 $T=17480 171360 1 0 $X=17290 $Y=168400
X342 1 2 ICV_3 $T=26220 138720 0 0 $X=26030 $Y=138480
X343 1 2 ICV_3 $T=59340 160480 0 0 $X=59150 $Y=160240
X344 1 2 ICV_3 $T=61180 116960 1 0 $X=60990 $Y=114000
X345 1 2 ICV_3 $T=62100 149600 0 0 $X=61910 $Y=149360
X346 1 2 ICV_3 $T=69460 138720 0 0 $X=69270 $Y=138480
X347 1 2 ICV_3 $T=73600 138720 1 0 $X=73410 $Y=135760
X348 1 2 ICV_3 $T=73600 144160 1 0 $X=73410 $Y=141200
X349 1 2 ICV_3 $T=101660 133280 1 0 $X=101470 $Y=130320
X350 1 2 ICV_3 $T=121900 155040 1 0 $X=121710 $Y=152080
X351 1 2 ICV_3 $T=129720 149600 1 0 $X=129530 $Y=146640
X352 1 2 ICV_3 $T=136620 122400 1 0 $X=136430 $Y=119440
X353 1 2 ICV_3 $T=143520 122400 0 0 $X=143330 $Y=122160
X354 1 2 ICV_3 $T=143520 155040 0 0 $X=143330 $Y=154800
X355 1 2 ICV_3 $T=157780 144160 1 0 $X=157590 $Y=141200
X356 1 2 ICV_3 $T=160540 155040 1 0 $X=160350 $Y=152080
X357 1 2 ICV_3 $T=163760 116960 0 0 $X=163570 $Y=116720
X358 1 2 ICV_3 $T=174340 127840 0 0 $X=174150 $Y=127600
X359 1 2 ICV_3 $T=178020 176800 1 0 $X=177830 $Y=173840
X360 1 2 ICV_3 $T=185840 171360 1 0 $X=185650 $Y=168400
X361 1 2 ICV_3 $T=187680 149600 0 0 $X=187490 $Y=149360
X362 1 2 ICV_3 $T=199640 144160 0 0 $X=199450 $Y=143920
X363 1 2 ICV_3 $T=199640 165920 0 0 $X=199450 $Y=165680
X364 1 2 ICV_3 $T=205160 176800 1 0 $X=204970 $Y=173840
X365 1 2 ICV_3 $T=213900 155040 1 0 $X=213710 $Y=152080
X366 1 2 ICV_3 $T=227700 171360 0 0 $X=227510 $Y=171120
X367 1 2 ICV_3 $T=230000 160480 1 0 $X=229810 $Y=157520
X368 1 2 ICV_3 $T=239200 176800 0 0 $X=239010 $Y=176560
X369 1 2 ICV_3 $T=251160 138720 1 0 $X=250970 $Y=135760
X370 1 2 ICV_3 $T=272780 149600 1 0 $X=272590 $Y=146640
X371 1 2 ICV_3 $T=280140 116960 1 0 $X=279950 $Y=114000
X372 1 2 ICV_3 $T=293020 155040 0 0 $X=292830 $Y=154800
X373 1 2 ICV_3 $T=298080 116960 1 0 $X=297890 $Y=114000
X374 1 2 ICV_3 $T=298080 155040 1 0 $X=297890 $Y=152080
X375 1 2 ICV_3 $T=311880 138720 0 0 $X=311690 $Y=138480
X376 1 2 ICV_3 $T=311880 144160 0 0 $X=311690 $Y=143920
X377 1 2 ICV_3 $T=311880 165920 0 0 $X=311690 $Y=165680
X378 1 2 ICV_3 $T=326140 155040 1 0 $X=325950 $Y=152080
X379 1 2 ICV_3 $T=363860 144160 0 0 $X=363670 $Y=143920
X380 1 2 ICV_3 $T=368000 155040 0 0 $X=367810 $Y=154800
X381 1 2 ICV_3 $T=382260 149600 1 0 $X=382070 $Y=146640
X382 1 2 ICV_3 $T=405260 155040 0 0 $X=405070 $Y=154800
X383 1 2 ICV_3 $T=406180 171360 0 0 $X=405990 $Y=171120
X384 1 2 ICV_3 $T=409860 160480 0 0 $X=409670 $Y=160240
X385 1 2 ICV_3 $T=410320 165920 1 0 $X=410130 $Y=162960
X386 1 2 ICV_3 $T=410320 176800 1 0 $X=410130 $Y=173840
X387 1 2 ICV_3 $T=413080 138720 1 0 $X=412890 $Y=135760
X388 1 2 ICV_3 $T=417680 171360 0 0 $X=417490 $Y=171120
X389 1 2 ICV_3 $T=424120 133280 0 0 $X=423930 $Y=133040
X390 1 2 ICV_3 $T=424120 171360 0 0 $X=423930 $Y=171120
X391 1 2 ICV_3 $T=426880 116960 0 0 $X=426690 $Y=116720
X392 1 2 ICV_3 $T=429640 176800 1 0 $X=429450 $Y=173840
X393 1 2 ICV_3 $T=432400 127840 0 0 $X=432210 $Y=127600
X394 1 2 ICV_3 $T=435160 171360 0 0 $X=434970 $Y=171120
X395 1 2 ICV_3 $T=438380 133280 1 0 $X=438190 $Y=130320
X396 1 2 ICV_3 $T=442060 165920 0 0 $X=441870 $Y=165680
X397 1 2 ICV_3 $T=454940 165920 0 0 $X=454750 $Y=165680
X398 1 2 ICV_3 $T=476100 138720 0 0 $X=475910 $Y=138480
X399 1 2 ICV_3 $T=477480 165920 1 0 $X=477290 $Y=162960
X400 1 2 ICV_3 $T=480240 160480 0 0 $X=480050 $Y=160240
X401 1 2 ICV_3 $T=491740 138720 0 0 $X=491550 $Y=138480
X402 1 2 ICV_3 $T=508300 155040 0 0 $X=508110 $Y=154800
X403 1 2 ICV_3 $T=522560 144160 1 0 $X=522370 $Y=141200
X404 1 2 ICV_3 $T=525320 160480 1 0 $X=525130 $Y=157520
X405 1 2 ICV_3 $T=533600 155040 1 0 $X=533410 $Y=152080
X406 1 2 ICV_3 $T=536360 144160 0 0 $X=536170 $Y=143920
X407 1 2 ICV_3 $T=550160 116960 0 0 $X=549970 $Y=116720
X408 1 2 ICV_3 $T=564420 133280 0 0 $X=564230 $Y=133040
X409 1 2 ICV_3 $T=567180 149600 0 0 $X=566990 $Y=149360
X410 1 2 ICV_3 $T=569480 160480 1 0 $X=569290 $Y=157520
X411 1 2 ICV_3 $T=578680 122400 1 0 $X=578490 $Y=119440
X412 1 2 ICV_3 $T=578680 138720 1 0 $X=578490 $Y=135760
X413 1 2 ICV_3 $T=606280 171360 0 0 $X=606090 $Y=171120
X414 1 2 ICV_3 $T=634800 116960 1 0 $X=634610 $Y=114000
X415 1 2 ICV_3 $T=634800 155040 1 0 $X=634610 $Y=152080
X416 1 2 ICV_3 $T=653660 155040 1 0 $X=653470 $Y=152080
X417 1 2 ICV_3 $T=662860 138720 1 0 $X=662670 $Y=135760
X418 1 2 ICV_3 $T=662860 160480 1 0 $X=662670 $Y=157520
X419 1 2 ICV_3 $T=677120 144160 1 0 $X=676930 $Y=141200
X420 1 2 ICV_3 $T=690920 144160 1 0 $X=690730 $Y=141200
X421 1 2 ICV_3 $T=704720 133280 0 0 $X=704530 $Y=133040
X422 1 2 ICV_3 $T=718980 155040 1 0 $X=718790 $Y=152080
X423 1 2 ICV_3 $T=735540 122400 0 0 $X=735350 $Y=122160
X424 1 2 ICV_3 $T=735540 144160 0 0 $X=735350 $Y=143920
X425 1 2 ICV_3 $T=735540 160480 0 0 $X=735350 $Y=160240
X426 1 2 ICV_3 $T=735540 165920 0 0 $X=735350 $Y=165680
X427 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=16560 160480 1 0 $X=16370 $Y=157520
X428 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=17480 165920 0 0 $X=17290 $Y=165680
X429 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=20240 122400 1 0 $X=20050 $Y=119440
X430 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=34040 165920 0 0 $X=33850 $Y=165680
X431 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=40480 144160 1 0 $X=40290 $Y=141200
X432 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=44620 171360 1 0 $X=44430 $Y=168400
X433 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=45080 127840 1 0 $X=44890 $Y=124880
X434 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=48300 155040 1 0 $X=48110 $Y=152080
X435 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=52440 165920 1 0 $X=52250 $Y=162960
X436 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=58880 116960 0 0 $X=58690 $Y=116720
X437 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=72680 127840 1 0 $X=72490 $Y=124880
X438 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=73140 122400 1 0 $X=72950 $Y=119440
X439 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=74980 127840 0 0 $X=74790 $Y=127600
X440 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=86480 176800 0 0 $X=86290 $Y=176560
X441 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=91080 165920 1 0 $X=90890 $Y=162960
X442 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=93840 155040 1 0 $X=93650 $Y=152080
X443 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=115000 165920 0 0 $X=114810 $Y=165680
X444 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=129260 144160 1 0 $X=129070 $Y=141200
X445 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=136620 127840 1 0 $X=136430 $Y=124880
X446 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=170660 171360 0 0 $X=170470 $Y=171120
X447 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=184920 127840 1 0 $X=184730 $Y=124880
X448 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=184920 138720 1 0 $X=184730 $Y=135760
X449 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=195960 133280 1 0 $X=195770 $Y=130320
X450 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=196880 138720 1 0 $X=196690 $Y=135760
X451 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=202400 160480 0 0 $X=202210 $Y=160240
X452 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=216660 122400 1 0 $X=216470 $Y=119440
X453 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=255300 122400 0 0 $X=255110 $Y=122160
X454 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=263120 171360 1 0 $X=262930 $Y=168400
X455 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=280140 144160 1 0 $X=279950 $Y=141200
X456 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=297620 171360 1 0 $X=297430 $Y=168400
X457 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=304980 176800 1 0 $X=304790 $Y=173840
X458 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=307280 155040 0 0 $X=307090 $Y=154800
X459 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=370760 171360 0 0 $X=370570 $Y=171120
X460 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=370760 176800 0 0 $X=370570 $Y=176560
X461 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=374900 138720 0 0 $X=374710 $Y=138480
X462 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=381800 171360 1 0 $X=381610 $Y=168400
X463 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=398820 144160 0 0 $X=398630 $Y=143920
X464 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=405720 171360 1 0 $X=405530 $Y=168400
X465 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=413080 127840 1 0 $X=412890 $Y=124880
X466 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=458160 155040 1 0 $X=457970 $Y=152080
X467 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=465980 165920 1 0 $X=465790 $Y=162960
X468 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=467360 144160 0 0 $X=467170 $Y=143920
X469 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=491280 144160 0 0 $X=491090 $Y=143920
X470 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=507380 171360 0 0 $X=507190 $Y=171120
X471 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=520720 116960 0 0 $X=520530 $Y=116720
X472 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=521640 165920 1 0 $X=521450 $Y=162960
X473 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=526700 133280 0 0 $X=526510 $Y=133040
X474 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=545100 122400 1 0 $X=544910 $Y=119440
X475 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=546020 138720 1 0 $X=545830 $Y=135760
X476 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=549700 155040 1 0 $X=549510 $Y=152080
X477 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=557980 144160 0 0 $X=557790 $Y=143920
X478 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=558440 127840 1 0 $X=558250 $Y=124880
X479 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=567180 165920 0 0 $X=566990 $Y=165680
X480 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=569480 176800 1 0 $X=569290 $Y=173840
X481 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=577760 165920 1 0 $X=577570 $Y=162960
X482 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=592020 155040 0 0 $X=591830 $Y=154800
X483 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=606280 138720 1 0 $X=606090 $Y=135760
X484 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=608580 138720 0 0 $X=608390 $Y=138480
X485 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=612260 116960 0 0 $X=612070 $Y=116720
X486 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=634340 122400 1 0 $X=634150 $Y=119440
X487 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=634340 133280 1 0 $X=634150 $Y=130320
X488 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=640780 165920 0 0 $X=640590 $Y=165680
X489 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=644920 122400 1 0 $X=644730 $Y=119440
X490 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=648140 165920 0 0 $X=647950 $Y=165680
X491 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=662400 149600 1 0 $X=662210 $Y=146640
X492 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=662400 165920 1 0 $X=662210 $Y=162960
X493 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=693680 160480 1 0 $X=693490 $Y=157520
X494 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=703800 116960 0 0 $X=703610 $Y=116720
X495 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=712540 149600 0 0 $X=712350 $Y=149360
X496 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=718520 127840 1 0 $X=718330 $Y=124880
X497 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=729100 149600 1 0 $X=728910 $Y=146640
X498 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=729100 155040 1 0 $X=728910 $Y=152080
X499 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=729100 171360 1 0 $X=728910 $Y=168400
X500 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=731860 144160 0 0 $X=731670 $Y=143920
X501 1 2 ICV_4 $T=6900 133280 0 0 $X=6710 $Y=133040
X502 1 2 ICV_4 $T=16560 144160 1 0 $X=16370 $Y=141200
X503 1 2 ICV_4 $T=44620 149600 1 0 $X=44430 $Y=146640
X504 1 2 ICV_4 $T=44620 165920 1 0 $X=44430 $Y=162960
X505 1 2 ICV_4 $T=48300 122400 1 0 $X=48110 $Y=119440
X506 1 2 ICV_4 $T=55660 176800 1 0 $X=55470 $Y=173840
X507 1 2 ICV_4 $T=76360 127840 1 0 $X=76170 $Y=124880
X508 1 2 ICV_4 $T=128800 122400 1 0 $X=128610 $Y=119440
X509 1 2 ICV_4 $T=166060 133280 1 0 $X=165870 $Y=130320
X510 1 2 ICV_4 $T=184920 138720 0 0 $X=184730 $Y=138480
X511 1 2 ICV_4 $T=203780 116960 1 0 $X=203590 $Y=114000
X512 1 2 ICV_4 $T=226780 165920 0 0 $X=226590 $Y=165680
X513 1 2 ICV_4 $T=230460 138720 0 0 $X=230270 $Y=138480
X514 1 2 ICV_4 $T=230460 160480 0 0 $X=230270 $Y=160240
X515 1 2 ICV_4 $T=232760 144160 1 0 $X=232570 $Y=141200
X516 1 2 ICV_4 $T=241040 171360 1 0 $X=240850 $Y=168400
X517 1 2 ICV_4 $T=241960 127840 0 0 $X=241770 $Y=127600
X518 1 2 ICV_4 $T=282900 116960 0 0 $X=282710 $Y=116720
X519 1 2 ICV_4 $T=300840 133280 1 0 $X=300650 $Y=130320
X520 1 2 ICV_4 $T=310960 122400 0 0 $X=310770 $Y=122160
X521 1 2 ICV_4 $T=310960 160480 0 0 $X=310770 $Y=160240
X522 1 2 ICV_4 $T=310960 171360 0 0 $X=310770 $Y=171120
X523 1 2 ICV_4 $T=342700 144160 0 0 $X=342510 $Y=143920
X524 1 2 ICV_4 $T=371220 160480 1 0 $X=371030 $Y=157520
X525 1 2 ICV_4 $T=382720 116960 0 0 $X=382530 $Y=116720
X526 1 2 ICV_4 $T=393760 149600 1 0 $X=393570 $Y=146640
X527 1 2 ICV_4 $T=438840 127840 0 0 $X=438650 $Y=127600
X528 1 2 ICV_4 $T=445280 138720 1 0 $X=445090 $Y=135760
X529 1 2 ICV_4 $T=454940 144160 0 0 $X=454750 $Y=143920
X530 1 2 ICV_4 $T=497260 138720 1 0 $X=497070 $Y=135760
X531 1 2 ICV_4 $T=507380 138720 0 0 $X=507190 $Y=138480
X532 1 2 ICV_4 $T=511060 165920 0 0 $X=510870 $Y=165680
X533 1 2 ICV_4 $T=511980 138720 1 0 $X=511790 $Y=135760
X534 1 2 ICV_4 $T=530380 138720 0 0 $X=530190 $Y=138480
X535 1 2 ICV_4 $T=538200 116960 1 0 $X=538010 $Y=114000
X536 1 2 ICV_4 $T=539120 155040 0 0 $X=538930 $Y=154800
X537 1 2 ICV_4 $T=577760 160480 1 0 $X=577570 $Y=157520
X538 1 2 ICV_4 $T=586040 122400 1 0 $X=585850 $Y=119440
X539 1 2 ICV_4 $T=602600 116960 0 0 $X=602410 $Y=116720
X540 1 2 ICV_4 $T=621460 165920 1 0 $X=621270 $Y=162960
X541 1 2 ICV_4 $T=623300 155040 1 0 $X=623110 $Y=152080
X542 1 2 ICV_4 $T=641240 144160 0 0 $X=641050 $Y=143920
X543 1 2 ICV_4 $T=665620 171360 1 0 $X=665430 $Y=168400
X544 1 2 ICV_4 $T=675740 171360 0 0 $X=675550 $Y=171120
X545 1 2 ICV_4 $T=731860 138720 0 0 $X=731670 $Y=138480
X546 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 133280 1 0 $X=6710 $Y=130320
X547 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 165920 1 0 $X=6710 $Y=162960
X548 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 171360 0 0 $X=6710 $Y=171120
X549 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 176800 1 0 $X=6710 $Y=173840
X550 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=29900 122400 0 0 $X=29710 $Y=122160
X551 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=29900 155040 0 0 $X=29710 $Y=154800
X552 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=34500 122400 1 0 $X=34310 $Y=119440
X553 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=57960 144160 0 0 $X=57770 $Y=143920
X554 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=83720 160480 1 0 $X=83530 $Y=157520
X555 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=86020 144160 0 0 $X=85830 $Y=143920
X556 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=90160 127840 0 0 $X=89970 $Y=127600
X557 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=91080 127840 1 0 $X=90890 $Y=124880
X558 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=93840 176800 1 0 $X=93650 $Y=173840
X559 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=98440 176800 0 0 $X=98250 $Y=176560
X560 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=118220 144160 1 0 $X=118030 $Y=141200
X561 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=118220 165920 0 0 $X=118030 $Y=165680
X562 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=120980 127840 1 0 $X=120790 $Y=124880
X563 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=128340 155040 1 0 $X=128150 $Y=152080
X564 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=139840 160480 1 0 $X=139650 $Y=157520
X565 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=142140 138720 0 0 $X=141950 $Y=138480
X566 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=150420 127840 0 0 $X=150230 $Y=127600
X567 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=153640 144160 0 0 $X=153450 $Y=143920
X568 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=165600 122400 1 0 $X=165410 $Y=119440
X569 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=165600 127840 1 0 $X=165410 $Y=124880
X570 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=170200 127840 0 0 $X=170010 $Y=127600
X571 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=184460 144160 1 0 $X=184270 $Y=141200
X572 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=184460 176800 1 0 $X=184270 $Y=173840
X573 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=197340 122400 0 0 $X=197150 $Y=122160
X574 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=212520 149600 1 0 $X=212330 $Y=146640
X575 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=226320 176800 0 0 $X=226130 $Y=176560
X576 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=242420 155040 0 0 $X=242230 $Y=154800
X577 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=252080 171360 1 0 $X=251890 $Y=168400
X578 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=264500 149600 0 0 $X=264310 $Y=149360
X579 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=275540 133280 0 0 $X=275350 $Y=133040
X580 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=276920 133280 1 0 $X=276730 $Y=130320
X581 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=281980 155040 1 0 $X=281790 $Y=152080
X582 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=286580 155040 0 0 $X=286390 $Y=154800
X583 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=298080 149600 0 0 $X=297890 $Y=149360
X584 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=299920 171360 0 0 $X=299730 $Y=171120
X585 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=309120 171360 1 0 $X=308930 $Y=168400
X586 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=314640 149600 0 0 $X=314450 $Y=149360
X587 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=322000 160480 0 0 $X=321810 $Y=160240
X588 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=333960 133280 0 0 $X=333770 $Y=133040
X589 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=338560 116960 0 0 $X=338370 $Y=116720
X590 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=345460 155040 1 0 $X=345270 $Y=152080
X591 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=347300 133280 1 0 $X=347110 $Y=130320
X592 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=352820 127840 1 0 $X=352630 $Y=124880
X593 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=380880 122400 1 0 $X=380690 $Y=119440
X594 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=381340 155040 0 0 $X=381150 $Y=154800
X595 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=385020 122400 1 0 $X=384830 $Y=119440
X596 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=387320 127840 0 0 $X=387130 $Y=127600
X597 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=394680 138720 0 0 $X=394490 $Y=138480
X598 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=398820 133280 0 0 $X=398630 $Y=133040
X599 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=398820 160480 0 0 $X=398630 $Y=160240
X600 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=408940 133280 0 0 $X=408750 $Y=133040
X601 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=422740 155040 0 0 $X=422550 $Y=154800
X602 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=435620 127840 1 0 $X=435430 $Y=124880
X603 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=436080 149600 0 0 $X=435890 $Y=149360
X604 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=438380 133280 0 0 $X=438190 $Y=133040
X605 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=439760 122400 0 0 $X=439570 $Y=122160
X606 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=448500 171360 1 0 $X=448310 $Y=168400
X607 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=450800 155040 0 0 $X=450610 $Y=154800
X608 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=483000 160480 0 0 $X=482810 $Y=160240
X609 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=487140 149600 0 0 $X=486950 $Y=149360
X610 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=491280 116960 0 0 $X=491090 $Y=116720
X611 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=493120 138720 1 0 $X=492930 $Y=135760
X612 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=500480 149600 0 0 $X=500290 $Y=149360
X613 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=502780 165920 0 0 $X=502590 $Y=165680
X614 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=506460 133280 1 0 $X=506270 $Y=130320
X615 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=506920 155040 1 0 $X=506730 $Y=152080
X616 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=521180 160480 1 0 $X=520990 $Y=157520
X617 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=521180 171360 1 0 $X=520990 $Y=168400
X618 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=521180 176800 1 0 $X=520990 $Y=173840
X619 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=538200 171360 1 0 $X=538010 $Y=168400
X620 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=565340 144160 1 0 $X=565150 $Y=141200
X621 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=571780 171360 0 0 $X=571590 $Y=171120
X622 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=595240 171360 0 0 $X=595050 $Y=171120
X623 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=615940 155040 0 0 $X=615750 $Y=154800
X624 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=630660 155040 0 0 $X=630470 $Y=154800
X625 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=644920 116960 1 0 $X=644730 $Y=114000
X626 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=644920 127840 1 0 $X=644730 $Y=124880
X627 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=689540 149600 1 0 $X=689350 $Y=146640
X628 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=690920 176800 0 0 $X=690730 $Y=176560
X629 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=693680 149600 1 0 $X=693490 $Y=146640
X630 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=697820 155040 1 0 $X=697630 $Y=152080
X631 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=698740 160480 1 0 $X=698550 $Y=157520
X632 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=699200 127840 1 0 $X=699010 $Y=124880
X633 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=717140 171360 0 0 $X=716950 $Y=171120
X634 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=727260 122400 1 0 $X=727070 $Y=119440
X635 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=731400 122400 0 0 $X=731210 $Y=122160
X636 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 116960 0 0 $X=6710 $Y=116720
X637 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 176800 0 0 $X=6710 $Y=176560
X638 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=85560 165920 1 0 $X=85370 $Y=162960
X639 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=111780 160480 1 0 $X=111590 $Y=157520
X640 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=154560 122400 1 0 $X=154370 $Y=119440
X641 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=210220 122400 1 0 $X=210030 $Y=119440
X642 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=213900 171360 0 0 $X=213710 $Y=171120
X643 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=214820 127840 0 0 $X=214630 $Y=127600
X644 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=346840 138720 0 0 $X=346650 $Y=138480
X645 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=347300 127840 1 0 $X=347110 $Y=124880
X646 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=352360 138720 0 0 $X=352170 $Y=138480
X647 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=363400 127840 0 0 $X=363210 $Y=127600
X648 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=417220 144160 1 0 $X=417030 $Y=141200
X649 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=457700 122400 1 0 $X=457510 $Y=119440
X650 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=475640 127840 1 0 $X=475450 $Y=124880
X651 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=515200 133280 0 0 $X=515010 $Y=133040
X652 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=532680 122400 0 0 $X=532490 $Y=122160
X653 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=657340 160480 1 0 $X=657150 $Y=157520
X654 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=687240 160480 1 0 $X=687050 $Y=157520
X655 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=701040 165920 0 0 $X=700850 $Y=165680
X656 1 2 13 15 2 19 1 sky130_fd_sc_hd__ebufn_2 $T=14720 176800 0 0 $X=14530 $Y=176560
X657 1 2 608 615 2 19 1 sky130_fd_sc_hd__ebufn_2 $T=26680 165920 0 0 $X=26490 $Y=165680
X658 1 2 635 589 2 37 1 sky130_fd_sc_hd__ebufn_2 $T=36340 144160 1 0 $X=36150 $Y=141200
X659 1 2 650 48 2 37 1 sky130_fd_sc_hd__ebufn_2 $T=43700 133280 1 0 $X=43510 $Y=130320
X660 1 2 49 51 2 38 1 sky130_fd_sc_hd__ebufn_2 $T=43700 176800 1 0 $X=43510 $Y=173840
X661 1 2 668 48 2 21 1 sky130_fd_sc_hd__ebufn_2 $T=51060 127840 1 0 $X=50870 $Y=124880
X662 1 2 665 48 2 38 1 sky130_fd_sc_hd__ebufn_2 $T=54740 116960 1 0 $X=54550 $Y=114000
X663 1 2 697 661 2 19 1 sky130_fd_sc_hd__ebufn_2 $T=63940 155040 0 0 $X=63750 $Y=154800
X664 1 2 715 695 2 21 1 sky130_fd_sc_hd__ebufn_2 $T=70840 127840 0 0 $X=70650 $Y=127600
X665 1 2 716 710 2 20 1 sky130_fd_sc_hd__ebufn_2 $T=71760 138720 0 0 $X=71570 $Y=138480
X666 1 2 793 752 2 32 1 sky130_fd_sc_hd__ebufn_2 $T=110860 165920 0 0 $X=110670 $Y=165680
X667 1 2 83 85 2 71 1 sky130_fd_sc_hd__ebufn_2 $T=111320 116960 1 0 $X=111130 $Y=114000
X668 1 2 809 814 2 19 1 sky130_fd_sc_hd__ebufn_2 $T=121900 165920 0 0 $X=121710 $Y=165680
X669 1 2 817 798 2 38 1 sky130_fd_sc_hd__ebufn_2 $T=124200 155040 1 0 $X=124010 $Y=152080
X670 1 2 811 790 2 37 1 sky130_fd_sc_hd__ebufn_2 $T=126500 138720 1 0 $X=126310 $Y=135760
X671 1 2 848 844 2 21 1 sky130_fd_sc_hd__ebufn_2 $T=139380 155040 0 0 $X=139190 $Y=154800
X672 1 2 887 858 2 21 1 sky130_fd_sc_hd__ebufn_2 $T=158700 165920 0 0 $X=158510 $Y=165680
X673 1 2 895 899 2 21 1 sky130_fd_sc_hd__ebufn_2 $T=161920 133280 1 0 $X=161730 $Y=130320
X674 1 2 900 892 2 21 1 sky130_fd_sc_hd__ebufn_2 $T=162840 155040 1 0 $X=162650 $Y=152080
X675 1 2 904 882 2 19 1 sky130_fd_sc_hd__ebufn_2 $T=166060 127840 0 0 $X=165870 $Y=127600
X676 1 2 907 882 2 38 1 sky130_fd_sc_hd__ebufn_2 $T=180320 144160 1 0 $X=180130 $Y=141200
X677 1 2 917 882 2 32 1 sky130_fd_sc_hd__ebufn_2 $T=180320 149600 1 0 $X=180130 $Y=146640
X678 1 2 935 911 2 32 1 sky130_fd_sc_hd__ebufn_2 $T=180320 176800 1 0 $X=180130 $Y=173840
X679 1 2 943 944 2 32 1 sky130_fd_sc_hd__ebufn_2 $T=185380 160480 0 0 $X=185190 $Y=160240
X680 1 2 978 944 2 20 1 sky130_fd_sc_hd__ebufn_2 $T=205160 165920 0 0 $X=204970 $Y=165680
X681 1 2 965 969 2 32 1 sky130_fd_sc_hd__ebufn_2 $T=209760 155040 1 0 $X=209570 $Y=152080
X682 1 2 1003 1004 2 162 1 sky130_fd_sc_hd__ebufn_2 $T=219420 122400 1 0 $X=219230 $Y=119440
X683 1 2 1056 1047 2 207 1 sky130_fd_sc_hd__ebufn_2 $T=251160 122400 0 0 $X=250970 $Y=122160
X684 1 2 1063 1054 2 189 1 sky130_fd_sc_hd__ebufn_2 $T=253920 165920 0 0 $X=253730 $Y=165680
X685 1 2 1085 212 2 162 1 sky130_fd_sc_hd__ebufn_2 $T=268180 176800 1 0 $X=267990 $Y=173840
X686 1 2 1100 1102 2 167 1 sky130_fd_sc_hd__ebufn_2 $T=274160 171360 1 0 $X=273970 $Y=168400
X687 1 2 1144 1117 2 201 1 sky130_fd_sc_hd__ebufn_2 $T=295320 155040 0 0 $X=295130 $Y=154800
X688 1 2 1177 1161 2 185 1 sky130_fd_sc_hd__ebufn_2 $T=310040 165920 1 0 $X=309850 $Y=162960
X689 1 2 1179 1160 2 200 1 sky130_fd_sc_hd__ebufn_2 $T=313720 133280 1 0 $X=313530 $Y=130320
X690 1 2 1204 1205 2 201 1 sky130_fd_sc_hd__ebufn_2 $T=324300 122400 1 0 $X=324110 $Y=119440
X691 1 2 1178 1142 2 201 1 sky130_fd_sc_hd__ebufn_2 $T=324300 133280 1 0 $X=324110 $Y=130320
X692 1 2 1287 1276 2 162 1 sky130_fd_sc_hd__ebufn_2 $T=367080 160480 1 0 $X=366890 $Y=157520
X693 1 2 1300 1272 2 167 1 sky130_fd_sc_hd__ebufn_2 $T=376740 122400 1 0 $X=376550 $Y=119440
X694 1 2 1364 1367 2 162 1 sky130_fd_sc_hd__ebufn_2 $T=408480 171360 1 0 $X=408290 $Y=168400
X695 1 2 1378 1367 2 188 1 sky130_fd_sc_hd__ebufn_2 $T=418600 155040 0 0 $X=418410 $Y=154800
X696 1 2 1384 1367 2 185 1 sky130_fd_sc_hd__ebufn_2 $T=419980 171360 0 0 $X=419790 $Y=171120
X697 1 2 1405 1400 2 216 1 sky130_fd_sc_hd__ebufn_2 $T=434700 127840 0 0 $X=434510 $Y=127600
X698 1 2 1438 319 2 316 1 sky130_fd_sc_hd__ebufn_2 $T=452180 171360 1 0 $X=451990 $Y=168400
X699 1 2 1444 321 2 325 1 sky130_fd_sc_hd__ebufn_2 $T=454480 116960 1 0 $X=454290 $Y=114000
X700 1 2 1451 1452 2 325 1 sky130_fd_sc_hd__ebufn_2 $T=458160 138720 1 0 $X=457970 $Y=135760
X701 1 2 1485 1487 2 342 1 sky130_fd_sc_hd__ebufn_2 $T=477940 138720 1 0 $X=477750 $Y=135760
X702 1 2 1486 1490 2 304 1 sky130_fd_sc_hd__ebufn_2 $T=478400 171360 0 0 $X=478210 $Y=171120
X703 1 2 1559 1538 2 325 1 sky130_fd_sc_hd__ebufn_2 $T=516580 149600 1 0 $X=516390 $Y=146640
X704 1 2 1574 1538 2 305 1 sky130_fd_sc_hd__ebufn_2 $T=527620 160480 1 0 $X=527430 $Y=157520
X705 1 2 1593 1596 2 365 1 sky130_fd_sc_hd__ebufn_2 $T=537280 144160 1 0 $X=537090 $Y=141200
X706 1 2 1603 1604 2 354 1 sky130_fd_sc_hd__ebufn_2 $T=540960 122400 1 0 $X=540770 $Y=119440
X707 1 2 1610 1596 2 351 1 sky130_fd_sc_hd__ebufn_2 $T=546020 138720 0 0 $X=545830 $Y=138480
X708 1 2 1662 1638 2 409 1 sky130_fd_sc_hd__ebufn_2 $T=590180 171360 0 0 $X=589990 $Y=171120
X709 1 2 1663 1638 2 405 1 sky130_fd_sc_hd__ebufn_2 $T=590640 165920 0 0 $X=590450 $Y=165680
X710 1 2 1632 440 2 423 1 sky130_fd_sc_hd__ebufn_2 $T=601680 155040 1 0 $X=601490 $Y=152080
X711 1 2 1692 1672 2 320 1 sky130_fd_sc_hd__ebufn_2 $T=604440 138720 0 0 $X=604250 $Y=138480
X712 1 2 1721 1722 2 397 1 sky130_fd_sc_hd__ebufn_2 $T=618700 160480 1 0 $X=618510 $Y=157520
X713 1 2 1742 517 2 320 1 sky130_fd_sc_hd__ebufn_2 $T=630200 116960 0 0 $X=630010 $Y=116720
X714 1 2 1813 531 2 365 1 sky130_fd_sc_hd__ebufn_2 $T=668380 127840 1 0 $X=668190 $Y=124880
X715 1 2 1807 1804 2 409 1 sky130_fd_sc_hd__ebufn_2 $T=674820 176800 1 0 $X=674630 $Y=173840
X716 1 2 1829 1837 2 356 1 sky130_fd_sc_hd__ebufn_2 $T=683100 160480 1 0 $X=682910 $Y=157520
X717 1 2 1864 1866 2 344 1 sky130_fd_sc_hd__ebufn_2 $T=695060 127840 1 0 $X=694870 $Y=124880
X718 1 2 1884 1892 2 342 1 sky130_fd_sc_hd__ebufn_2 $T=713460 155040 1 0 $X=713270 $Y=152080
X719 1 2 1906 1868 2 351 1 sky130_fd_sc_hd__ebufn_2 $T=717140 138720 1 0 $X=716950 $Y=135760
X720 1 2 1922 1920 2 371 1 sky130_fd_sc_hd__ebufn_2 $T=723120 122400 1 0 $X=722930 $Y=119440
X721 1 2 1932 549 2 354 1 sky130_fd_sc_hd__ebufn_2 $T=730940 116960 0 0 $X=730750 $Y=116720
X834 1 2 598 605 19 ICV_6 $T=19780 144160 1 0 $X=19590 $Y=141200
X835 1 2 596 589 21 ICV_6 $T=19780 149600 1 0 $X=19590 $Y=146640
X836 1 2 607 615 20 ICV_6 $T=19780 171360 1 0 $X=19590 $Y=168400
X837 1 2 612 615 11 ICV_6 $T=19780 176800 1 0 $X=19590 $Y=173840
X838 1 2 629 599 38 ICV_6 $T=33580 116960 0 0 $X=33390 $Y=116720
X839 1 2 628 605 40 ICV_6 $T=33580 133280 0 0 $X=33390 $Y=133040
X840 1 2 662 649 40 ICV_6 $T=47840 149600 1 0 $X=47650 $Y=146640
X841 1 2 657 649 38 ICV_6 $T=47840 165920 1 0 $X=47650 $Y=162960
X842 1 2 722 710 11 ICV_6 $T=75900 116960 1 0 $X=75710 $Y=114000
X843 1 2 689 695 11 ICV_6 $T=75900 133280 1 0 $X=75710 $Y=130320
X844 1 2 709 683 11 ICV_6 $T=75900 171360 1 0 $X=75710 $Y=168400
X845 1 2 704 710 32 ICV_6 $T=89700 133280 0 0 $X=89510 $Y=133040
X846 1 2 738 744 37 ICV_6 $T=89700 149600 0 0 $X=89510 $Y=149360
X847 1 2 771 754 38 ICV_6 $T=103960 122400 1 0 $X=103770 $Y=119440
X848 1 2 774 754 19 ICV_6 $T=103960 127840 1 0 $X=103770 $Y=124880
X849 1 2 781 783 11 ICV_6 $T=103960 133280 1 0 $X=103770 $Y=130320
X850 1 2 764 744 32 ICV_6 $T=103960 144160 1 0 $X=103770 $Y=141200
X851 1 2 778 752 40 ICV_6 $T=103960 171360 1 0 $X=103770 $Y=168400
X852 1 2 803 783 20 ICV_6 $T=117760 116960 0 0 $X=117570 $Y=116720
X853 1 2 805 783 40 ICV_6 $T=117760 122400 0 0 $X=117570 $Y=122160
X854 1 2 802 783 37 ICV_6 $T=117760 127840 0 0 $X=117570 $Y=127600
X855 1 2 801 783 21 ICV_6 $T=117760 133280 0 0 $X=117570 $Y=133040
X856 1 2 836 824 20 ICV_6 $T=132020 122400 1 0 $X=131830 $Y=119440
X857 1 2 833 824 40 ICV_6 $T=132020 127840 1 0 $X=131830 $Y=124880
X858 1 2 831 824 21 ICV_6 $T=132020 133280 1 0 $X=131830 $Y=130320
X859 1 2 821 93 11 ICV_6 $T=132020 176800 1 0 $X=131830 $Y=173840
X860 1 2 861 103 37 ICV_6 $T=145820 127840 0 0 $X=145630 $Y=127600
X861 1 2 863 858 40 ICV_6 $T=145820 165920 0 0 $X=145630 $Y=165680
X862 1 2 919 892 37 ICV_6 $T=173880 149600 0 0 $X=173690 $Y=149360
X863 1 2 886 112 38 ICV_6 $T=173880 176800 0 0 $X=173690 $Y=176560
X864 1 2 942 892 32 ICV_6 $T=188140 155040 1 0 $X=187950 $Y=152080
X865 1 2 1020 1004 150 ICV_6 $T=230000 116960 0 0 $X=229810 $Y=116720
X866 1 2 1043 195 189 ICV_6 $T=244260 122400 1 0 $X=244070 $Y=119440
X867 1 2 1065 195 166 ICV_6 $T=258060 116960 0 0 $X=257870 $Y=116720
X868 1 2 1066 195 150 ICV_6 $T=258060 122400 0 0 $X=257870 $Y=122160
X869 1 2 1064 212 166 ICV_6 $T=258060 176800 0 0 $X=257870 $Y=176560
X870 1 2 1089 1097 207 ICV_6 $T=272320 133280 1 0 $X=272130 $Y=130320
X871 1 2 222 212 167 ICV_6 $T=272320 176800 1 0 $X=272130 $Y=173840
X872 1 2 1121 1102 162 ICV_6 $T=286120 165920 0 0 $X=285930 $Y=165680
X873 1 2 1120 1102 188 ICV_6 $T=286120 171360 0 0 $X=285930 $Y=171120
X874 1 2 1119 1102 186 ICV_6 $T=286120 176800 0 0 $X=285930 $Y=176560
X875 1 2 1154 1118 167 ICV_6 $T=300380 160480 1 0 $X=300190 $Y=157520
X876 1 2 1151 1118 185 ICV_6 $T=300380 176800 1 0 $X=300190 $Y=173840
X877 1 2 1174 1142 214 ICV_6 $T=314180 122400 0 0 $X=313990 $Y=122160
X878 1 2 1165 1142 207 ICV_6 $T=314180 127840 0 0 $X=313990 $Y=127600
X879 1 2 1207 1205 200 ICV_6 $T=328440 133280 1 0 $X=328250 $Y=130320
X880 1 2 1212 1191 150 ICV_6 $T=328440 144160 1 0 $X=328250 $Y=141200
X881 1 2 1235 1191 167 ICV_6 $T=342240 138720 0 0 $X=342050 $Y=138480
X882 1 2 1242 1214 167 ICV_6 $T=342240 165920 0 0 $X=342050 $Y=165680
X883 1 2 1243 1214 188 ICV_6 $T=342240 171360 0 0 $X=342050 $Y=171120
X884 1 2 1271 1272 188 ICV_6 $T=356500 127840 1 0 $X=356310 $Y=124880
X885 1 2 1263 1261 186 ICV_6 $T=356500 138720 1 0 $X=356310 $Y=135760
X886 1 2 1269 1274 162 ICV_6 $T=356500 149600 1 0 $X=356310 $Y=146640
X887 1 2 1267 1276 185 ICV_6 $T=356500 165920 1 0 $X=356310 $Y=162960
X888 1 2 1268 244 188 ICV_6 $T=356500 176800 1 0 $X=356310 $Y=173840
X889 1 2 1288 1272 150 ICV_6 $T=370300 116960 0 0 $X=370110 $Y=116720
X890 1 2 1292 1261 188 ICV_6 $T=370300 133280 0 0 $X=370110 $Y=133040
X891 1 2 1293 1261 166 ICV_6 $T=370300 138720 0 0 $X=370110 $Y=138480
X892 1 2 1295 1274 189 ICV_6 $T=370300 149600 0 0 $X=370110 $Y=149360
X893 1 2 1319 1326 167 ICV_6 $T=384560 138720 1 0 $X=384370 $Y=135760
X894 1 2 1317 1324 162 ICV_6 $T=384560 144160 1 0 $X=384370 $Y=141200
X895 1 2 1346 259 186 ICV_6 $T=398360 127840 0 0 $X=398170 $Y=127600
X896 1 2 1344 1326 188 ICV_6 $T=398360 138720 0 0 $X=398170 $Y=138480
X897 1 2 1339 1324 150 ICV_6 $T=398360 165920 0 0 $X=398170 $Y=165680
X898 1 2 268 270 166 ICV_6 $T=398360 176800 0 0 $X=398170 $Y=176560
X899 1 2 1373 1372 188 ICV_6 $T=412620 144160 1 0 $X=412430 $Y=141200
X900 1 2 1368 1367 166 ICV_6 $T=412620 171360 1 0 $X=412430 $Y=168400
X901 1 2 1390 1372 166 ICV_6 $T=426420 127840 0 0 $X=426230 $Y=127600
X902 1 2 1389 1372 185 ICV_6 $T=426420 138720 0 0 $X=426230 $Y=138480
X903 1 2 1414 293 185 ICV_6 $T=440680 122400 1 0 $X=440490 $Y=119440
X904 1 2 1412 1410 214 ICV_6 $T=440680 138720 1 0 $X=440490 $Y=135760
X905 1 2 1404 1410 216 ICV_6 $T=440680 149600 1 0 $X=440490 $Y=146640
X906 1 2 1439 321 300 ICV_6 $T=454480 116960 0 0 $X=454290 $Y=116720
X907 1 2 1465 321 309 ICV_6 $T=468740 122400 1 0 $X=468550 $Y=119440
X908 1 2 1496 1501 345 ICV_6 $T=482540 122400 0 0 $X=482350 $Y=122160
X909 1 2 1493 1487 354 ICV_6 $T=482540 127840 0 0 $X=482350 $Y=127600
X910 1 2 1491 1490 320 ICV_6 $T=482540 149600 0 0 $X=482350 $Y=149360
X911 1 2 374 361 356 ICV_6 $T=496800 116960 1 0 $X=496610 $Y=114000
X912 1 2 1520 1501 371 ICV_6 $T=496800 122400 1 0 $X=496610 $Y=119440
X913 1 2 1542 1534 342 ICV_6 $T=510600 133280 0 0 $X=510410 $Y=133040
X914 1 2 1540 1534 356 ICV_6 $T=510600 138720 0 0 $X=510410 $Y=138480
X915 1 2 1566 386 405 ICV_6 $T=524860 171360 1 0 $X=524670 $Y=168400
X916 1 2 1591 1600 405 ICV_6 $T=538660 165920 0 0 $X=538470 $Y=165680
X917 1 2 1595 1600 407 ICV_6 $T=538660 171360 0 0 $X=538470 $Y=171120
X918 1 2 1581 393 423 ICV_6 $T=538660 176800 0 0 $X=538470 $Y=176560
X919 1 2 1619 1600 423 ICV_6 $T=552920 160480 1 0 $X=552730 $Y=157520
X920 1 2 1617 1600 444 ICV_6 $T=552920 171360 1 0 $X=552730 $Y=168400
X921 1 2 1641 1596 344 ICV_6 $T=566720 155040 0 0 $X=566530 $Y=154800
X922 1 2 1660 1639 304 ICV_6 $T=580980 127840 1 0 $X=580790 $Y=124880
X923 1 2 1655 1596 345 ICV_6 $T=580980 133280 1 0 $X=580790 $Y=130320
X924 1 2 1658 1638 397 ICV_6 $T=580980 160480 1 0 $X=580790 $Y=157520
X925 1 2 1674 1679 294 ICV_6 $T=594780 138720 0 0 $X=594590 $Y=138480
X926 1 2 1675 1679 300 ICV_6 $T=594780 149600 0 0 $X=594590 $Y=149360
X927 1 2 1680 1682 396 ICV_6 $T=594780 165920 0 0 $X=594590 $Y=165680
X928 1 2 1699 1682 391 ICV_6 $T=609040 165920 1 0 $X=608850 $Y=162960
X929 1 2 1696 1682 409 ICV_6 $T=609040 171360 1 0 $X=608850 $Y=168400
X930 1 2 1703 1682 423 ICV_6 $T=609040 176800 1 0 $X=608850 $Y=173840
X931 1 2 1726 488 300 ICV_6 $T=622840 116960 0 0 $X=622650 $Y=116720
X932 1 2 1717 1719 305 ICV_6 $T=622840 127840 0 0 $X=622650 $Y=127600
X933 1 2 1725 1722 391 ICV_6 $T=622840 160480 0 0 $X=622650 $Y=160240
X934 1 2 1752 1756 316 ICV_6 $T=637100 138720 1 0 $X=636910 $Y=135760
X935 1 2 1754 1756 300 ICV_6 $T=637100 144160 1 0 $X=636910 $Y=141200
X936 1 2 1775 1756 309 ICV_6 $T=650900 144160 0 0 $X=650710 $Y=143920
X937 1 2 1764 1771 407 ICV_6 $T=650900 171360 0 0 $X=650710 $Y=171120
X938 1 2 1782 523 444 ICV_6 $T=650900 176800 0 0 $X=650710 $Y=176560
X939 1 2 1802 1794 351 ICV_6 $T=665160 138720 1 0 $X=664970 $Y=135760
X940 1 2 1803 1794 371 ICV_6 $T=665160 149600 1 0 $X=664970 $Y=146640
X941 1 2 1836 531 354 ICV_6 $T=678960 122400 0 0 $X=678770 $Y=122160
X942 1 2 1831 1837 351 ICV_6 $T=678960 144160 0 0 $X=678770 $Y=143920
X943 1 2 1828 1837 371 ICV_6 $T=678960 160480 0 0 $X=678770 $Y=160240
X944 1 2 1857 1837 345 ICV_6 $T=693220 155040 1 0 $X=693030 $Y=152080
X945 1 2 1860 1841 397 ICV_6 $T=693220 165920 1 0 $X=693030 $Y=162960
X946 1 2 1865 1841 409 ICV_6 $T=693220 171360 1 0 $X=693030 $Y=168400
X947 1 2 1850 1841 405 ICV_6 $T=693220 176800 1 0 $X=693030 $Y=173840
X948 1 2 1917 1892 354 ICV_6 $T=721280 160480 1 0 $X=721090 $Y=157520
X1036 1 2 583 9 2 609 1 sky130_fd_sc_hd__dfxtp_1 $T=10580 133280 1 0 $X=10390 $Y=130320
X1037 1 2 587 26 2 632 1 sky130_fd_sc_hd__dfxtp_1 $T=24380 171360 1 0 $X=24190 $Y=168400
X1038 1 2 44 27 2 650 1 sky130_fd_sc_hd__dfxtp_1 $T=36800 127840 0 0 $X=36610 $Y=127600
X1039 1 2 639 28 2 662 1 sky130_fd_sc_hd__dfxtp_1 $T=38640 155040 1 0 $X=38450 $Y=152080
X1040 1 2 702 9 2 719 1 sky130_fd_sc_hd__dfxtp_1 $T=68540 133280 1 0 $X=68350 $Y=130320
X1041 1 2 685 9 2 722 1 sky130_fd_sc_hd__dfxtp_1 $T=69460 133280 0 0 $X=69270 $Y=133040
X1042 1 2 62 27 2 725 1 sky130_fd_sc_hd__dfxtp_1 $T=79120 176800 0 0 $X=78930 $Y=176560
X1043 1 2 73 6 2 774 1 sky130_fd_sc_hd__dfxtp_1 $T=94760 127840 1 0 $X=94570 $Y=124880
X1044 1 2 745 6 2 779 1 sky130_fd_sc_hd__dfxtp_1 $T=97520 160480 0 0 $X=97330 $Y=160240
X1045 1 2 761 6 2 786 1 sky130_fd_sc_hd__dfxtp_1 $T=99820 138720 0 0 $X=99630 $Y=138480
X1046 1 2 761 27 2 811 1 sky130_fd_sc_hd__dfxtp_1 $T=111780 138720 1 0 $X=111590 $Y=135760
X1047 1 2 761 5 2 826 1 sky130_fd_sc_hd__dfxtp_1 $T=121900 144160 1 0 $X=121710 $Y=141200
X1048 1 2 816 6 2 834 1 sky130_fd_sc_hd__dfxtp_1 $T=124660 127840 1 0 $X=124470 $Y=124880
X1049 1 2 829 26 2 854 1 sky130_fd_sc_hd__dfxtp_1 $T=139840 149600 1 0 $X=139650 $Y=146640
X1050 1 2 100 9 2 874 1 sky130_fd_sc_hd__dfxtp_1 $T=144900 133280 1 0 $X=144710 $Y=130320
X1051 1 2 884 6 2 904 1 sky130_fd_sc_hd__dfxtp_1 $T=157780 138720 0 0 $X=157590 $Y=138480
X1052 1 2 906 27 2 925 1 sky130_fd_sc_hd__dfxtp_1 $T=169740 138720 1 0 $X=169550 $Y=135760
X1053 1 2 928 26 2 946 1 sky130_fd_sc_hd__dfxtp_1 $T=180780 133280 1 0 $X=180590 $Y=130320
X1054 1 2 941 29 2 973 1 sky130_fd_sc_hd__dfxtp_1 $T=192280 144160 0 0 $X=192090 $Y=143920
X1055 1 2 933 9 2 994 1 sky130_fd_sc_hd__dfxtp_1 $T=205620 165920 1 0 $X=205430 $Y=162960
X1056 1 2 998 156 2 1003 1 sky130_fd_sc_hd__dfxtp_1 $T=222180 122400 0 0 $X=221990 $Y=122160
X1057 1 2 998 155 2 1020 1 sky130_fd_sc_hd__dfxtp_1 $T=222640 116960 0 0 $X=222450 $Y=116720
X1058 1 2 1000 178 2 1038 1 sky130_fd_sc_hd__dfxtp_1 $T=235980 138720 1 0 $X=235790 $Y=135760
X1059 1 2 183 153 2 1065 1 sky130_fd_sc_hd__dfxtp_1 $T=248400 116960 0 0 $X=248210 $Y=116720
X1060 1 2 1041 206 2 1070 1 sky130_fd_sc_hd__dfxtp_1 $T=252080 127840 1 0 $X=251890 $Y=124880
X1061 1 2 1040 178 2 1063 1 sky130_fd_sc_hd__dfxtp_1 $T=255760 171360 1 0 $X=255570 $Y=168400
X1062 1 2 1076 194 2 1101 1 sky130_fd_sc_hd__dfxtp_1 $T=268180 149600 0 0 $X=267990 $Y=149360
X1063 1 2 225 153 2 1147 1 sky130_fd_sc_hd__dfxtp_1 $T=290720 116960 1 0 $X=290530 $Y=114000
X1064 1 2 1133 206 2 1149 1 sky130_fd_sc_hd__dfxtp_1 $T=292100 127840 1 0 $X=291910 $Y=124880
X1065 1 2 1124 154 2 1154 1 sky130_fd_sc_hd__dfxtp_1 $T=293020 160480 1 0 $X=292830 $Y=157520
X1066 1 2 1133 204 2 1139 1 sky130_fd_sc_hd__dfxtp_1 $T=293480 122400 0 0 $X=293290 $Y=122160
X1067 1 2 1156 155 2 1176 1 sky130_fd_sc_hd__dfxtp_1 $T=303600 160480 0 0 $X=303410 $Y=160240
X1068 1 2 1156 175 2 1177 1 sky130_fd_sc_hd__dfxtp_1 $T=303600 171360 0 0 $X=303410 $Y=171120
X1069 1 2 1133 193 2 1178 1 sky130_fd_sc_hd__dfxtp_1 $T=304980 127840 0 0 $X=304790 $Y=127600
X1070 1 2 1156 176 2 1188 1 sky130_fd_sc_hd__dfxtp_1 $T=312800 171360 1 0 $X=312610 $Y=168400
X1071 1 2 1187 206 2 1219 1 sky130_fd_sc_hd__dfxtp_1 $T=326600 127840 0 0 $X=326410 $Y=127600
X1072 1 2 243 179 2 1268 1 sky130_fd_sc_hd__dfxtp_1 $T=349140 176800 0 0 $X=348950 $Y=176560
X1073 1 2 1253 176 2 1275 1 sky130_fd_sc_hd__dfxtp_1 $T=350980 160480 0 0 $X=350790 $Y=160240
X1074 1 2 243 178 2 248 1 sky130_fd_sc_hd__dfxtp_1 $T=356500 171360 0 0 $X=356310 $Y=171120
X1075 1 2 1257 155 2 1288 1 sky130_fd_sc_hd__dfxtp_1 $T=361100 127840 1 0 $X=360910 $Y=124880
X1076 1 2 1257 154 2 1300 1 sky130_fd_sc_hd__dfxtp_1 $T=366620 116960 1 0 $X=366430 $Y=114000
X1077 1 2 255 156 2 1306 1 sky130_fd_sc_hd__dfxtp_1 $T=370760 176800 1 0 $X=370570 $Y=173840
X1078 1 2 1301 176 2 1320 1 sky130_fd_sc_hd__dfxtp_1 $T=375820 155040 1 0 $X=375630 $Y=152080
X1079 1 2 1301 175 2 1331 1 sky130_fd_sc_hd__dfxtp_1 $T=385020 155040 0 0 $X=384830 $Y=154800
X1080 1 2 1327 153 2 1334 1 sky130_fd_sc_hd__dfxtp_1 $T=386400 165920 0 0 $X=386210 $Y=165680
X1081 1 2 1312 154 2 1343 1 sky130_fd_sc_hd__dfxtp_1 $T=391000 127840 0 0 $X=390810 $Y=127600
X1082 1 2 1350 155 2 1366 1 sky130_fd_sc_hd__dfxtp_1 $T=402500 160480 0 0 $X=402310 $Y=160240
X1083 1 2 1350 178 2 1365 1 sky130_fd_sc_hd__dfxtp_1 $T=403420 160480 1 0 $X=403230 $Y=157520
X1084 1 2 269 154 2 277 1 sky130_fd_sc_hd__dfxtp_1 $T=405260 116960 1 0 $X=405070 $Y=114000
X1085 1 2 1354 153 2 1390 1 sky130_fd_sc_hd__dfxtp_1 $T=416300 133280 1 0 $X=416110 $Y=130320
X1086 1 2 279 283 2 1397 1 sky130_fd_sc_hd__dfxtp_1 $T=422280 176800 1 0 $X=422090 $Y=173840
X1087 1 2 1377 154 2 1418 1 sky130_fd_sc_hd__dfxtp_1 $T=434240 116960 0 0 $X=434050 $Y=116720
X1088 1 2 1466 338 2 1480 1 sky130_fd_sc_hd__dfxtp_1 $T=468740 138720 0 0 $X=468550 $Y=138480
X1089 1 2 1467 340 2 1502 1 sky130_fd_sc_hd__dfxtp_1 $T=477020 133280 1 0 $X=476830 $Y=130320
X1090 1 2 1466 343 2 1488 1 sky130_fd_sc_hd__dfxtp_1 $T=477940 144160 1 0 $X=477750 $Y=141200
X1091 1 2 1475 283 2 1519 1 sky130_fd_sc_hd__dfxtp_1 $T=488060 165920 1 0 $X=487870 $Y=162960
X1092 1 2 1523 357 2 1540 1 sky130_fd_sc_hd__dfxtp_1 $T=500020 138720 0 0 $X=499830 $Y=138480
X1093 1 2 1524 379 2 385 1 sky130_fd_sc_hd__dfxtp_1 $T=500020 171360 0 0 $X=499830 $Y=171120
X1094 1 2 1523 341 2 1542 1 sky130_fd_sc_hd__dfxtp_1 $T=500480 127840 0 0 $X=500290 $Y=127600
X1095 1 2 1580 378 2 1597 1 sky130_fd_sc_hd__dfxtp_1 $T=531300 160480 0 0 $X=531110 $Y=160240
X1096 1 2 1606 343 2 1615 1 sky130_fd_sc_hd__dfxtp_1 $T=542340 155040 1 0 $X=542150 $Y=152080
X1097 1 2 428 382 2 435 1 sky130_fd_sc_hd__dfxtp_1 $T=544180 176800 1 0 $X=543990 $Y=173840
X1098 1 2 1588 358 2 1624 1 sky130_fd_sc_hd__dfxtp_1 $T=547860 127840 0 0 $X=547670 $Y=127600
X1099 1 2 1626 357 2 1620 1 sky130_fd_sc_hd__dfxtp_1 $T=557060 133280 0 0 $X=556870 $Y=133040
X1100 1 2 1628 281 2 1637 1 sky130_fd_sc_hd__dfxtp_1 $T=559820 122400 1 0 $X=559630 $Y=119440
X1101 1 2 1625 395 2 1658 1 sky130_fd_sc_hd__dfxtp_1 $T=570400 165920 1 0 $X=570210 $Y=162960
X1102 1 2 452 303 2 1656 1 sky130_fd_sc_hd__dfxtp_1 $T=578680 116960 0 0 $X=578490 $Y=116720
X1103 1 2 1666 281 2 1675 1 sky130_fd_sc_hd__dfxtp_1 $T=586500 138720 0 0 $X=586310 $Y=138480
X1104 1 2 1668 380 2 1696 1 sky130_fd_sc_hd__dfxtp_1 $T=598920 171360 0 0 $X=598730 $Y=171120
X1105 1 2 500 475 2 1712 1 sky130_fd_sc_hd__dfxtp_1 $T=610880 176800 0 0 $X=610690 $Y=176560
X1106 1 2 477 283 2 1723 1 sky130_fd_sc_hd__dfxtp_1 $T=614100 116960 1 0 $X=613910 $Y=114000
X1107 1 2 1710 379 2 1728 1 sky130_fd_sc_hd__dfxtp_1 $T=615020 171360 0 0 $X=614830 $Y=171120
X1108 1 2 1710 399 2 1746 1 sky130_fd_sc_hd__dfxtp_1 $T=625600 171360 0 0 $X=625410 $Y=171120
X1109 1 2 1748 298 2 1760 1 sky130_fd_sc_hd__dfxtp_1 $T=634340 155040 0 0 $X=634150 $Y=154800
X1110 1 2 522 379 2 1782 1 sky130_fd_sc_hd__dfxtp_1 $T=643540 176800 0 0 $X=643350 $Y=176560
X1111 1 2 1749 307 2 1772 1 sky130_fd_sc_hd__dfxtp_1 $T=649060 133280 1 0 $X=648870 $Y=130320
X1112 1 2 1779 338 2 1805 1 sky130_fd_sc_hd__dfxtp_1 $T=657340 144160 0 0 $X=657150 $Y=143920
X1113 1 2 529 358 2 1815 1 sky130_fd_sc_hd__dfxtp_1 $T=662860 122400 0 0 $X=662670 $Y=122160
X1114 1 2 529 357 2 535 1 sky130_fd_sc_hd__dfxtp_1 $T=670220 116960 1 0 $X=670030 $Y=114000
X1115 1 2 1806 340 2 1847 1 sky130_fd_sc_hd__dfxtp_1 $T=679420 133280 1 0 $X=679230 $Y=130320
X1116 1 2 1844 339 2 1864 1 sky130_fd_sc_hd__dfxtp_1 $T=687240 122400 0 0 $X=687050 $Y=122160
X1117 1 2 1835 400 2 1870 1 sky130_fd_sc_hd__dfxtp_1 $T=691840 160480 0 0 $X=691650 $Y=160240
X1118 1 2 1871 378 2 1882 1 sky130_fd_sc_hd__dfxtp_1 $T=697820 165920 1 0 $X=697630 $Y=162960
X1119 1 2 1869 341 2 1884 1 sky130_fd_sc_hd__dfxtp_1 $T=698740 144160 0 0 $X=698550 $Y=143920
X1120 1 2 1869 357 2 1886 1 sky130_fd_sc_hd__dfxtp_1 $T=699200 155040 0 0 $X=699010 $Y=154800
X1121 1 2 1869 338 2 1893 1 sky130_fd_sc_hd__dfxtp_1 $T=702420 160480 1 0 $X=702230 $Y=157520
X1122 1 2 1869 343 2 1917 1 sky130_fd_sc_hd__dfxtp_1 $T=712080 155040 0 0 $X=711890 $Y=154800
X1123 1 2 606 605 21 586 8 606 ICV_13 $T=10120 133280 0 0 $X=9930 $Y=133040
X1124 1 2 619 599 37 583 27 619 ICV_13 $T=22080 127840 1 0 $X=21890 $Y=124880
X1125 1 2 624 602 37 584 26 617 ICV_13 $T=22080 149600 0 0 $X=21890 $Y=149360
X1126 1 2 626 599 40 583 28 626 ICV_13 $T=23000 122400 1 0 $X=22810 $Y=119440
X1127 1 2 640 45 47 4 34 640 ICV_13 $T=28520 116960 1 0 $X=28330 $Y=114000
X1128 1 2 643 605 38 586 29 643 ICV_13 $T=30820 133280 1 0 $X=30630 $Y=130320
X1129 1 2 645 649 19 639 6 645 ICV_13 $T=34960 160480 0 0 $X=34770 $Y=160240
X1130 1 2 647 654 37 641 27 647 ICV_13 $T=35880 138720 0 0 $X=35690 $Y=138480
X1131 1 2 659 661 38 639 27 652 ICV_13 $T=36800 155040 0 0 $X=36610 $Y=154800
X1132 1 2 653 649 21 639 8 653 ICV_13 $T=36800 165920 0 0 $X=36610 $Y=165680
X1133 1 2 660 48 20 44 5 660 ICV_13 $T=38180 116960 0 0 $X=37990 $Y=116720
X1134 1 2 681 661 37 666 29 659 ICV_13 $T=48300 155040 0 0 $X=48110 $Y=154800
X1135 1 2 682 683 37 664 27 682 ICV_13 $T=48300 171360 1 0 $X=48110 $Y=168400
X1136 1 2 690 661 40 666 28 690 ICV_13 $T=55200 165920 1 0 $X=55010 $Y=162960
X1137 1 2 692 695 19 675 27 694 ICV_13 $T=57040 133280 1 0 $X=56850 $Y=130320
X1138 1 2 700 683 21 664 8 700 ICV_13 $T=58880 176800 1 0 $X=58690 $Y=173840
X1139 1 2 706 710 19 685 28 711 ICV_13 $T=63480 149600 1 0 $X=63290 $Y=146640
X1140 1 2 713 695 32 675 26 713 ICV_13 $T=63940 122400 0 0 $X=63750 $Y=122160
X1141 1 2 717 723 19 701 26 718 ICV_13 $T=68080 155040 0 0 $X=67890 $Y=154800
X1142 1 2 719 741 11 702 29 731 ICV_13 $T=77740 127840 0 0 $X=77550 $Y=127600
X1143 1 2 733 741 20 702 5 733 ICV_13 $T=78200 116960 0 0 $X=78010 $Y=116720
X1144 1 2 718 723 32 701 5 736 ICV_13 $T=78200 149600 0 0 $X=78010 $Y=149360
X1145 1 2 742 744 20 726 5 742 ICV_13 $T=79120 138720 1 0 $X=78930 $Y=135760
X1146 1 2 730 741 21 702 6 740 ICV_13 $T=79580 127840 1 0 $X=79390 $Y=124880
X1147 1 2 746 70 71 63 7 746 ICV_13 $T=80500 116960 1 0 $X=80310 $Y=114000
X1148 1 2 747 741 40 702 28 747 ICV_13 $T=80500 133280 1 0 $X=80310 $Y=130320
X1149 1 2 758 760 21 745 8 758 ICV_13 $T=87400 160480 1 0 $X=87210 $Y=157520
X1150 1 2 772 754 21 73 27 773 ICV_13 $T=94300 133280 0 0 $X=94110 $Y=133040
X1151 1 2 775 754 40 73 28 775 ICV_13 $T=95220 122400 0 0 $X=95030 $Y=122160
X1152 1 2 795 760 32 745 26 795 ICV_13 $T=104880 160480 0 0 $X=104690 $Y=160240
X1153 1 2 820 814 20 791 26 822 ICV_13 $T=119140 171360 1 0 $X=118950 $Y=168400
X1154 1 2 828 790 11 761 9 828 ICV_13 $T=121900 138720 0 0 $X=121710 $Y=138480
X1155 1 2 834 824 19 816 26 838 ICV_13 $T=132020 122400 0 0 $X=131830 $Y=122160
X1156 1 2 845 824 38 816 29 845 ICV_13 $T=132480 116960 0 0 $X=132290 $Y=116720
X1157 1 2 853 93 32 89 26 853 ICV_13 $T=133860 176800 0 0 $X=133670 $Y=176560
X1158 1 2 855 851 40 837 28 855 ICV_13 $T=134320 138720 1 0 $X=134130 $Y=135760
X1159 1 2 865 103 40 100 28 865 ICV_13 $T=139380 127840 1 0 $X=139190 $Y=124880
X1160 1 2 850 844 37 829 9 872 ICV_13 $T=143520 160480 1 0 $X=143330 $Y=157520
X1161 1 2 890 899 37 108 8 895 ICV_13 $T=154560 133280 0 0 $X=154370 $Y=133040
X1162 1 2 889 899 32 108 6 897 ICV_13 $T=161460 122400 0 0 $X=161270 $Y=122160
X1163 1 2 909 911 20 898 5 909 ICV_13 $T=161920 165920 1 0 $X=161730 $Y=162960
X1164 1 2 923 927 21 906 8 923 ICV_13 $T=169280 133280 1 0 $X=169090 $Y=130320
X1165 1 2 936 927 32 906 26 936 ICV_13 $T=174340 122400 0 0 $X=174150 $Y=122160
X1166 1 2 961 951 21 932 8 961 ICV_13 $T=185840 122400 0 0 $X=185650 $Y=122160
X1167 1 2 946 950 32 941 8 963 ICV_13 $T=188140 138720 0 0 $X=187950 $Y=138480
X1168 1 2 964 969 37 941 26 965 ICV_13 $T=188600 149600 1 0 $X=188410 $Y=146640
X1169 1 2 968 944 21 933 8 968 ICV_13 $T=189520 160480 0 0 $X=189330 $Y=160240
X1170 1 2 981 950 40 928 28 981 ICV_13 $T=199640 138720 1 0 $X=199450 $Y=135760
X1171 1 2 979 950 20 928 9 985 ICV_13 $T=202400 133280 0 0 $X=202210 $Y=133040
X1172 1 2 983 969 11 932 9 982 ICV_13 $T=204240 127840 1 0 $X=204050 $Y=124880
X1173 1 2 1008 995 166 1001 153 1008 ICV_13 $T=215280 165920 0 0 $X=215090 $Y=165680
X1174 1 2 1012 1004 167 998 154 1012 ICV_13 $T=216660 127840 1 0 $X=216470 $Y=124880
X1175 1 2 1017 995 167 1001 154 1017 ICV_13 $T=216660 171360 1 0 $X=216470 $Y=168400
X1176 1 2 1027 1004 188 998 179 1027 ICV_13 $T=230460 122400 0 0 $X=230270 $Y=122160
X1177 1 2 1028 1004 189 998 178 1028 ICV_13 $T=230460 127840 0 0 $X=230270 $Y=127600
X1178 1 2 1030 997 188 1002 179 1030 ICV_13 $T=230460 144160 0 0 $X=230270 $Y=143920
X1179 1 2 1035 997 186 1002 176 1035 ICV_13 $T=230920 149600 0 0 $X=230730 $Y=149360
X1180 1 2 1036 995 188 1001 179 1036 ICV_13 $T=230920 165920 1 0 $X=230730 $Y=162960
X1181 1 2 1037 1004 186 998 176 1037 ICV_13 $T=232760 122400 1 0 $X=232570 $Y=119440
X1182 1 2 1057 1047 203 1041 197 1057 ICV_13 $T=244720 133280 1 0 $X=244530 $Y=130320
X1183 1 2 1053 1042 210 1044 193 1055 ICV_13 $T=244720 149600 1 0 $X=244530 $Y=146640
X1184 1 2 1059 1054 185 1040 175 1059 ICV_13 $T=244720 176800 1 0 $X=244530 $Y=173840
X1185 1 2 1079 1042 214 1044 205 1079 ICV_13 $T=258520 138720 0 0 $X=258330 $Y=138480
X1186 1 2 1081 1047 211 1041 213 1081 ICV_13 $T=259440 127840 1 0 $X=259250 $Y=124880
X1187 1 2 1099 1096 214 1076 196 1105 ICV_13 $T=272780 160480 1 0 $X=272590 $Y=157520
X1188 1 2 1104 1102 166 1084 155 1115 ICV_13 $T=275540 165920 1 0 $X=275350 $Y=162960
X1189 1 2 1122 1102 189 1084 178 1122 ICV_13 $T=278300 171360 1 0 $X=278110 $Y=168400
X1190 1 2 1112 1094 214 1075 204 1126 ICV_13 $T=280140 122400 1 0 $X=279950 $Y=119440
X1191 1 2 1140 1097 200 1077 204 1140 ICV_13 $T=287040 138720 1 0 $X=286850 $Y=135760
X1192 1 2 1126 1094 200 1077 193 1128 ICV_13 $T=288420 133280 1 0 $X=288230 $Y=130320
X1193 1 2 1147 227 166 225 156 1155 ICV_13 $T=293940 116960 0 0 $X=293750 $Y=116720
X1194 1 2 1181 1142 203 1133 213 1173 ICV_13 $T=308200 127840 1 0 $X=308010 $Y=124880
X1195 1 2 1180 1160 211 1148 213 1180 ICV_13 $T=308200 138720 1 0 $X=308010 $Y=135760
X1196 1 2 1175 1142 210 1133 197 1181 ICV_13 $T=310960 122400 1 0 $X=310770 $Y=119440
X1197 1 2 1193 1161 189 1153 156 1196 ICV_13 $T=314640 155040 0 0 $X=314450 $Y=154800
X1198 1 2 1201 1160 207 1148 196 1201 ICV_13 $T=316480 144160 1 0 $X=316290 $Y=141200
X1199 1 2 1209 1205 210 1187 194 1209 ICV_13 $T=321080 122400 0 0 $X=320890 $Y=122160
X1200 1 2 1211 1191 162 1192 156 1211 ICV_13 $T=321540 138720 0 0 $X=321350 $Y=138480
X1201 1 2 1216 1191 189 1192 178 1216 ICV_13 $T=322460 133280 0 0 $X=322270 $Y=133040
X1202 1 2 1224 233 189 232 178 1224 ICV_13 $T=327060 116960 0 0 $X=326870 $Y=116720
X1203 1 2 1227 1218 167 1208 153 1226 ICV_13 $T=328900 144160 0 0 $X=328710 $Y=143920
X1204 1 2 1231 1191 166 1192 153 1231 ICV_13 $T=333040 144160 1 0 $X=332850 $Y=141200
X1205 1 2 1234 1191 186 1192 176 1234 ICV_13 $T=334880 138720 1 0 $X=334690 $Y=135760
X1206 1 2 1232 1205 207 1187 205 1238 ICV_13 $T=335800 127840 1 0 $X=335610 $Y=124880
X1207 1 2 1240 1205 211 1187 213 1240 ICV_13 $T=336260 122400 1 0 $X=336070 $Y=119440
X1208 1 2 1241 1214 162 1206 156 1241 ICV_13 $T=336260 165920 1 0 $X=336070 $Y=162960
X1209 1 2 1260 244 167 235 156 245 ICV_13 $T=345000 176800 1 0 $X=344810 $Y=173840
X1210 1 2 1262 1261 189 1248 178 1262 ICV_13 $T=347300 127840 0 0 $X=347110 $Y=127600
X1211 1 2 1266 1276 166 1252 153 1277 ICV_13 $T=352360 144160 0 0 $X=352170 $Y=143920
X1212 1 2 1280 244 166 243 155 250 ICV_13 $T=358340 165920 0 0 $X=358150 $Y=165680
X1213 1 2 1291 1276 188 1253 156 1287 ICV_13 $T=361100 165920 1 0 $X=360910 $Y=162960
X1214 1 2 1290 1274 186 1252 154 1298 ICV_13 $T=365240 144160 1 0 $X=365050 $Y=141200
X1215 1 2 1304 1272 162 1257 178 1302 ICV_13 $T=368460 127840 1 0 $X=368270 $Y=124880
X1216 1 2 1307 258 189 255 155 1310 ICV_13 $T=372600 165920 1 0 $X=372410 $Y=162960
X1217 1 2 1286 1276 150 1301 178 1318 ICV_13 $T=374900 149600 0 0 $X=374710 $Y=149360
X1218 1 2 1335 259 189 257 155 264 ICV_13 $T=385940 116960 0 0 $X=385750 $Y=116720
X1219 1 2 1341 259 185 1312 175 1341 ICV_13 $T=388700 122400 1 0 $X=388510 $Y=119440
X1220 1 2 1343 259 167 1312 176 1346 ICV_13 $T=391460 133280 1 0 $X=391270 $Y=130320
X1221 1 2 1356 1284 186 1327 175 1340 ICV_13 $T=398820 176800 1 0 $X=398630 $Y=173840
X1222 1 2 1352 1326 150 1349 153 1361 ICV_13 $T=401580 144160 0 0 $X=401390 $Y=143920
X1223 1 2 1371 1372 167 1354 155 1379 ICV_13 $T=412620 133280 0 0 $X=412430 $Y=133040
X1224 1 2 1382 1360 186 1349 176 1382 ICV_13 $T=413540 149600 0 0 $X=413350 $Y=149360
X1225 1 2 1406 302 304 1396 296 1406 ICV_13 $T=428260 165920 1 0 $X=428070 $Y=162960
X1226 1 2 1408 302 305 1396 298 1408 ICV_13 $T=429180 171360 1 0 $X=428990 $Y=168400
X1227 1 2 1430 1410 210 1398 194 1430 ICV_13 $T=441600 144160 0 0 $X=441410 $Y=143920
X1228 1 2 1431 1400 210 1395 213 1423 ICV_13 $T=442060 127840 0 0 $X=441870 $Y=127600
X1229 1 2 1427 1400 207 1395 194 1431 ICV_13 $T=442060 133280 0 0 $X=441870 $Y=133040
X1230 1 2 1454 1452 294 1440 283 1454 ICV_13 $T=454940 138720 0 0 $X=454750 $Y=138480
X1231 1 2 1448 1449 300 160 200 327 ICV_13 $T=455400 149600 0 0 $X=455210 $Y=149360
X1232 1 2 1443 319 304 314 307 328 ICV_13 $T=455860 176800 0 0 $X=455670 $Y=176560
X1233 1 2 1457 319 300 314 281 1457 ICV_13 $T=456320 171360 1 0 $X=456130 $Y=168400
X1234 1 2 1460 1452 304 1440 296 1460 ICV_13 $T=457240 133280 1 0 $X=457050 $Y=130320
X1235 1 2 1468 1452 320 1440 295 1468 ICV_13 $T=462300 122400 0 0 $X=462110 $Y=122160
X1236 1 2 1469 1449 316 1426 303 1469 ICV_13 $T=462300 155040 0 0 $X=462110 $Y=154800
X1237 1 2 1480 1473 345 1466 340 1483 ICV_13 $T=470120 144160 0 0 $X=469930 $Y=143920
X1238 1 2 1482 349 316 335 295 1484 ICV_13 $T=470120 176800 1 0 $X=469930 $Y=173840
X1239 1 2 1507 349 304 335 296 1507 ICV_13 $T=483000 176800 0 0 $X=482810 $Y=176560
X1240 1 2 1509 1487 344 1467 339 1509 ICV_13 $T=484380 133280 1 0 $X=484190 $Y=130320
X1241 1 2 1513 1487 365 1466 360 1504 ICV_13 $T=485300 144160 1 0 $X=485110 $Y=141200
X1242 1 2 1515 1490 316 1475 303 1515 ICV_13 $T=486680 160480 0 0 $X=486490 $Y=160240
X1243 1 2 1526 1501 351 1476 357 1525 ICV_13 $T=494960 116960 0 0 $X=494770 $Y=116720
X1244 1 2 1543 1534 354 1523 343 1543 ICV_13 $T=500480 138720 1 0 $X=500290 $Y=135760
X1245 1 2 1545 361 371 347 358 1545 ICV_13 $T=501400 116960 1 0 $X=501210 $Y=114000
X1246 1 2 1558 1538 304 1547 296 1558 ICV_13 $T=509680 160480 1 0 $X=509490 $Y=157520
X1247 1 2 1578 1555 304 1548 303 1583 ICV_13 $T=525320 122400 1 0 $X=525130 $Y=119440
X1248 1 2 1573 1555 325 1548 298 1576 ICV_13 $T=525320 127840 1 0 $X=525130 $Y=124880
X1249 1 2 1612 433 351 424 343 1611 ICV_13 $T=541420 116960 1 0 $X=541230 $Y=114000
X1250 1 2 1615 1602 354 1606 338 1616 ICV_13 $T=542340 155040 0 0 $X=542150 $Y=154800
X1251 1 2 1614 1600 409 1580 379 1617 ICV_13 $T=543260 165920 0 0 $X=543070 $Y=165680
X1252 1 2 1621 1600 397 1580 395 1621 ICV_13 $T=546480 160480 0 0 $X=546290 $Y=160240
X1253 1 2 1616 1602 345 1606 357 1631 ICV_13 $T=553840 155040 0 0 $X=553650 $Y=154800
X1254 1 2 1613 1602 351 1606 339 1633 ICV_13 $T=554300 149600 1 0 $X=554110 $Y=146640
X1255 1 2 1637 1639 300 1588 341 1622 ICV_13 $T=555220 122400 0 0 $X=555030 $Y=122160
X1256 1 2 1634 1604 365 1588 360 1634 ICV_13 $T=555220 127840 0 0 $X=555030 $Y=127600
X1257 1 2 1649 1639 325 1628 310 1649 ICV_13 $T=567180 122400 1 0 $X=566990 $Y=119440
X1258 1 2 1653 1638 407 1625 382 1653 ICV_13 $T=568100 171360 1 0 $X=567910 $Y=168400
X1259 1 2 1654 1596 371 1626 358 1654 ICV_13 $T=569020 144160 1 0 $X=568830 $Y=141200
X1260 1 2 1656 463 316 452 283 466 ICV_13 $T=569480 116960 1 0 $X=569290 $Y=114000
X1261 1 2 1669 1639 294 1628 283 1669 ICV_13 $T=583280 122400 0 0 $X=583090 $Y=122160
X1262 1 2 1673 1672 325 1665 307 1681 ICV_13 $T=589260 122400 1 0 $X=589070 $Y=119440
X1263 1 2 1683 1682 405 1668 382 1685 ICV_13 $T=596620 171360 1 0 $X=596430 $Y=168400
X1264 1 2 1689 1672 305 1665 281 1691 ICV_13 $T=597080 133280 1 0 $X=596890 $Y=130320
X1265 1 2 1695 1679 320 1666 295 1695 ICV_13 $T=597540 149600 1 0 $X=597350 $Y=146640
X1266 1 2 1697 1682 444 1668 379 1697 ICV_13 $T=599380 165920 0 0 $X=599190 $Y=165680
X1267 1 2 1690 1682 397 1668 400 1703 ICV_13 $T=603060 160480 0 0 $X=602870 $Y=160240
X1268 1 2 1708 1707 294 1688 283 1708 ICV_13 $T=604440 155040 0 0 $X=604250 $Y=154800
X1269 1 2 1716 1719 320 1704 295 1716 ICV_13 $T=611340 127840 1 0 $X=611150 $Y=124880
X1270 1 2 1720 1719 325 1704 298 1717 ICV_13 $T=611340 127840 0 0 $X=611150 $Y=127600
X1271 1 2 1727 1722 407 1710 380 1734 ICV_13 $T=622380 171360 1 0 $X=622190 $Y=168400
X1272 1 2 1739 1719 294 1704 283 1739 ICV_13 $T=623300 122400 0 0 $X=623110 $Y=122160
X1273 1 2 1745 1722 396 1710 388 1745 ICV_13 $T=624680 165920 1 0 $X=624490 $Y=162960
X1274 1 2 1758 517 305 519 298 1758 ICV_13 $T=634340 116960 0 0 $X=634150 $Y=116720
X1275 1 2 1767 1743 294 1755 388 1768 ICV_13 $T=637560 160480 0 0 $X=637370 $Y=160240
X1276 1 2 1770 1771 405 1755 399 1770 ICV_13 $T=637560 171360 1 0 $X=637370 $Y=168400
X1277 1 2 1791 1763 325 519 310 1788 ICV_13 $T=647680 122400 1 0 $X=647490 $Y=119440
X1278 1 2 1793 517 304 519 307 1790 ICV_13 $T=648600 116960 1 0 $X=648410 $Y=114000
X1279 1 2 1796 1763 294 1749 283 1796 ICV_13 $T=651360 122400 0 0 $X=651170 $Y=122160
X1280 1 2 1805 1794 345 1779 341 1816 ICV_13 $T=665620 144160 1 0 $X=665430 $Y=141200
X1281 1 2 534 523 397 522 380 1819 ICV_13 $T=666080 176800 0 0 $X=665890 $Y=176560
X1282 1 2 1827 1804 405 1795 399 1827 ICV_13 $T=668840 171360 1 0 $X=668650 $Y=168400
X1283 1 2 1830 531 345 529 343 1836 ICV_13 $T=672520 127840 1 0 $X=672330 $Y=124880
X1284 1 2 1843 531 342 529 341 1843 ICV_13 $T=677580 116960 1 0 $X=677390 $Y=114000
X1285 1 2 1846 1824 365 1806 360 1846 ICV_13 $T=679420 127840 0 0 $X=679230 $Y=127600
X1286 1 2 1849 1824 371 1806 358 1849 ICV_13 $T=679420 138720 0 0 $X=679230 $Y=138480
X1287 1 2 540 539 405 536 382 1851 ICV_13 $T=679420 176800 0 0 $X=679230 $Y=176560
X1288 1 2 1878 1866 342 1844 341 1878 ICV_13 $T=694600 122400 0 0 $X=694410 $Y=122160
X1289 1 2 543 537 345 538 357 1890 ICV_13 $T=700580 116960 1 0 $X=700390 $Y=114000
X1290 1 2 1890 537 356 538 341 1905 ICV_13 $T=707480 116960 0 0 $X=707290 $Y=116720
X1291 1 2 1901 1891 397 1871 388 1899 ICV_13 $T=707480 160480 0 0 $X=707290 $Y=160240
X1292 1 2 1894 1892 365 1871 400 1910 ICV_13 $T=709780 160480 1 0 $X=709590 $Y=157520
X1293 1 2 1923 546 397 544 399 1924 ICV_13 $T=714840 176800 0 0 $X=714650 $Y=176560
X1294 1 2 1934 1914 371 1916 340 1931 ICV_13 $T=718980 133280 0 0 $X=718790 $Y=133040
X1295 1 2 1938 1914 354 1916 343 1938 ICV_13 $T=720360 138720 0 0 $X=720170 $Y=138480
X1296 1 2 1948 546 391 544 378 1948 ICV_13 $T=730480 176800 1 0 $X=730290 $Y=173840
X1297 1 2 1949 1920 365 1904 360 1949 ICV_13 $T=730940 122400 1 0 $X=730750 $Y=119440
X1298 1 2 1952 1928 391 1919 378 1952 ICV_13 $T=730940 165920 1 0 $X=730750 $Y=162960
X1299 1 2 585 5 592 592 602 20 ICV_14 $T=6900 155040 1 0 $X=6710 $Y=152080
X1300 1 2 585 6 593 593 602 19 ICV_14 $T=6900 155040 0 0 $X=6710 $Y=154800
X1301 1 2 641 26 676 676 654 32 ICV_14 $T=46460 133280 0 0 $X=46270 $Y=133040
X1302 1 2 664 5 712 712 683 20 ICV_14 $T=62560 171360 1 0 $X=62370 $Y=168400
X1303 1 2 701 28 724 720 723 37 ICV_14 $T=68540 165920 0 0 $X=68350 $Y=165680
X1304 1 2 702 27 732 732 741 37 ICV_14 $T=76820 133280 0 0 $X=76630 $Y=133040
X1305 1 2 788 6 807 807 783 19 ICV_14 $T=108560 127840 1 0 $X=108370 $Y=124880
X1306 1 2 837 29 852 852 851 38 ICV_14 $T=132940 144160 0 0 $X=132750 $Y=143920
X1307 1 2 884 27 921 915 882 20 ICV_14 $T=167900 144160 1 0 $X=167710 $Y=141200
X1308 1 2 884 8 920 902 882 40 ICV_14 $T=167900 149600 1 0 $X=167710 $Y=146640
X1309 1 2 941 9 983 973 969 38 ICV_14 $T=200100 149600 1 0 $X=199910 $Y=146640
X1310 1 2 151 154 1006 1006 163 167 ICV_14 $T=213900 176800 0 0 $X=213710 $Y=176560
X1311 1 2 1108 206 1138 1138 1117 216 ICV_14 $T=285660 155040 1 0 $X=285470 $Y=152080
X1312 1 2 230 153 1190 1194 231 150 ICV_14 $T=312340 176800 1 0 $X=312150 $Y=173840
X1313 1 2 232 176 1199 1199 233 186 ICV_14 $T=314640 116960 1 0 $X=314450 $Y=114000
X1314 1 2 232 175 1200 1200 233 185 ICV_14 $T=314640 116960 0 0 $X=314450 $Y=116720
X1315 1 2 1208 179 1245 1245 1218 188 ICV_14 $T=336260 149600 1 0 $X=336070 $Y=146640
X1316 1 2 1252 175 1294 1294 1274 185 ICV_14 $T=361100 149600 1 0 $X=360910 $Y=146640
X1317 1 2 1257 176 1299 1299 1272 186 ICV_14 $T=364320 122400 1 0 $X=364130 $Y=119440
X1318 1 2 257 153 1332 1332 265 166 ICV_14 $T=385020 116960 1 0 $X=384830 $Y=114000
X1319 1 2 1303 176 1347 1347 1326 186 ICV_14 $T=390540 138720 1 0 $X=390350 $Y=135760
X1320 1 2 1349 156 1363 1361 1360 166 ICV_14 $T=401120 149600 0 0 $X=400930 $Y=149360
X1321 1 2 1350 154 1383 1383 1367 167 ICV_14 $T=412620 165920 0 0 $X=412430 $Y=165680
X1322 1 2 1349 154 1385 1385 1360 167 ICV_14 $T=413080 144160 0 0 $X=412890 $Y=143920
X1323 1 2 1349 175 1386 1386 1360 185 ICV_14 $T=413080 149600 1 0 $X=412890 $Y=146640
X1324 1 2 1395 205 1401 1401 1400 214 ICV_14 $T=425960 133280 1 0 $X=425770 $Y=130320
X1325 1 2 1440 303 1456 1456 1452 316 ICV_14 $T=454940 133280 0 0 $X=454750 $Y=133040
X1326 1 2 1466 341 1471 1483 1473 351 ICV_14 $T=469200 149600 1 0 $X=469010 $Y=146640
X1327 1 2 160 354 1530 1536 1538 294 ICV_14 $T=497260 160480 1 0 $X=497070 $Y=157520
X1328 1 2 1524 382 1565 1567 393 407 ICV_14 $T=512440 171360 0 0 $X=512250 $Y=171120
X1329 1 2 1688 303 1709 1709 1707 316 ICV_14 $T=605820 149600 0 0 $X=605630 $Y=149360
X1330 1 2 1733 298 1753 1753 1756 305 ICV_14 $T=627900 138720 0 0 $X=627710 $Y=138480
X1331 1 2 1755 400 1785 1785 1771 423 ICV_14 $T=644920 160480 1 0 $X=644730 $Y=157520
X1332 1 2 529 340 1811 1811 531 351 ICV_14 $T=660100 116960 0 0 $X=659910 $Y=116720
X1333 1 2 1918 339 1929 1940 1921 371 ICV_14 $T=721740 149600 0 0 $X=721550 $Y=149360
X1334 1 2 1904 357 1951 1951 1920 356 ICV_14 $T=730020 133280 1 0 $X=729830 $Y=130320
X1335 1 2 545 338 551 1953 1914 365 ICV_14 $T=730480 116960 1 0 $X=730290 $Y=114000
X1336 1 2 1916 360 1953 1958 1921 365 ICV_14 $T=730480 138720 1 0 $X=730290 $Y=135760
X1337 1 2 703 695 20 675 29 696 688 695 40 ICV_15 $T=57500 122400 1 0 $X=57310 $Y=119440
X1338 1 2 797 798 32 782 26 797 796 798 20 ICV_15 $T=106260 155040 1 0 $X=106070 $Y=152080
X1339 1 2 873 103 32 100 6 864 864 103 19 ICV_15 $T=138920 122400 1 0 $X=138730 $Y=119440
X1340 1 2 924 927 19 906 28 922 922 927 40 ICV_15 $T=169280 127840 1 0 $X=169090 $Y=124880
X1341 1 2 962 950 37 932 27 949 952 950 21 ICV_15 $T=182620 127840 0 0 $X=182430 $Y=127600
X1342 1 2 1019 997 162 1002 156 1019 1007 1014 150 ICV_15 $T=217120 144160 1 0 $X=216930 $Y=141200
X1343 1 2 1116 1118 150 1084 175 1107 1107 1102 185 ICV_15 $T=270480 176800 0 0 $X=270290 $Y=176560
X1344 1 2 1228 239 189 235 154 1222 1222 239 167 ICV_15 $T=326140 176800 0 0 $X=325950 $Y=176560
X1345 1 2 1541 1534 365 1523 358 1529 1529 1534 371 ICV_15 $T=497720 144160 1 0 $X=497530 $Y=141200
X1346 1 2 1568 386 397 1524 400 1569 1544 386 409 ICV_15 $T=514280 165920 0 0 $X=514090 $Y=165680
X1347 1 2 1605 1604 344 1588 357 1607 1607 1604 356 ICV_15 $T=536820 127840 1 0 $X=536630 $Y=124880
X1348 1 2 1747 1722 423 1710 400 1747 1728 1722 444 ICV_15 $T=625140 165920 0 0 $X=624950 $Y=165680
X1349 1 2 1765 1763 320 1749 303 1762 1762 1763 316 ICV_15 $T=634800 122400 0 0 $X=634610 $Y=122160
X1350 1 2 1769 1771 397 1755 378 1787 1787 1771 391 ICV_15 $T=646760 165920 1 0 $X=646570 $Y=162960
X1351 1 2 1895 1866 351 1844 358 1896 1897 1866 354 ICV_15 $T=702880 127840 1 0 $X=702690 $Y=124880
X1352 1 2 1944 1921 345 1918 343 1933 1933 1921 354 ICV_15 $T=719440 155040 0 0 $X=719250 $Y=154800
X1353 1 2 587 8 611 611 615 21 ICV_16 $T=10580 171360 0 0 $X=10390 $Y=171120
X1354 1 2 586 26 620 620 605 32 ICV_16 $T=21620 133280 0 0 $X=21430 $Y=133040
X1355 1 2 587 29 630 618 602 32 ICV_16 $T=23460 165920 1 0 $X=23270 $Y=162960
X1356 1 2 584 28 634 634 589 40 ICV_16 $T=24380 144160 1 0 $X=24190 $Y=141200
X1357 1 2 584 29 627 597 589 19 ICV_16 $T=24380 149600 1 0 $X=24190 $Y=146640
X1358 1 2 639 9 651 656 654 11 ICV_16 $T=36340 149600 0 0 $X=36150 $Y=149360
X1359 1 2 726 28 743 739 744 21 ICV_16 $T=78660 149600 1 0 $X=78470 $Y=146640
X1360 1 2 729 8 751 751 752 21 ICV_16 $T=81880 171360 1 0 $X=81690 $Y=168400
X1361 1 2 726 26 764 765 744 38 ICV_16 $T=90620 149600 1 0 $X=90430 $Y=146640
X1362 1 2 782 28 794 776 790 32 ICV_16 $T=104420 149600 1 0 $X=104230 $Y=146640
X1363 1 2 782 5 796 794 798 40 ICV_16 $T=104880 149600 0 0 $X=104690 $Y=149360
X1364 1 2 788 29 804 804 783 38 ICV_16 $T=108560 122400 1 0 $X=108370 $Y=119440
X1365 1 2 782 29 817 806 814 38 ICV_16 $T=117300 160480 1 0 $X=117110 $Y=157520
X1366 1 2 829 8 848 847 851 11 ICV_16 $T=132020 149600 0 0 $X=131830 $Y=149360
X1367 1 2 108 9 894 894 899 11 ICV_16 $T=154100 127840 0 0 $X=153910 $Y=127600
X1368 1 2 906 29 926 931 927 20 ICV_16 $T=170200 116960 1 0 $X=170010 $Y=114000
X1369 1 2 898 29 934 934 911 38 ICV_16 $T=173420 165920 1 0 $X=173230 $Y=162960
X1370 1 2 898 6 938 938 911 19 ICV_16 $T=173880 171360 1 0 $X=173690 $Y=168400
X1371 1 2 1002 153 1015 1015 997 166 ICV_16 $T=216200 144160 0 0 $X=216010 $Y=143920
X1372 1 2 151 176 1022 1022 163 186 ICV_16 $T=228160 176800 1 0 $X=227970 $Y=173840
X1373 1 2 1040 153 1074 218 219 150 ICV_16 $T=256220 176800 1 0 $X=256030 $Y=173840
X1374 1 2 1108 204 1141 1130 1117 214 ICV_16 $T=286580 144160 0 0 $X=286390 $Y=143920
X1375 1 2 1206 175 1221 1223 1214 186 ICV_16 $T=325220 171360 0 0 $X=325030 $Y=171120
X1376 1 2 1301 154 1336 1333 1324 188 ICV_16 $T=386400 149600 0 0 $X=386210 $Y=149360
X1377 1 2 269 153 1357 1357 274 166 ICV_16 $T=400200 122400 1 0 $X=400010 $Y=119440
X1378 1 2 1440 307 1455 1455 1452 309 ICV_16 $T=454940 127840 0 0 $X=454750 $Y=127600
X1379 1 2 1440 281 1459 1453 1452 305 ICV_16 $T=456780 127840 1 0 $X=456590 $Y=124880
X1380 1 2 1467 358 1516 1516 1487 371 ICV_16 $T=487140 127840 0 0 $X=486950 $Y=127600
X1381 1 2 392 400 1581 415 393 409 ICV_16 $T=523940 176800 0 0 $X=523750 $Y=176560
X1382 1 2 1606 358 1630 1630 1602 371 ICV_16 $T=553380 155040 1 0 $X=553190 $Y=152080
X1383 1 2 473 475 480 1646 440 396 ICV_16 $T=582360 176800 0 0 $X=582170 $Y=176560
X1384 1 2 1704 303 1736 1736 1719 316 ICV_16 $T=622380 122400 1 0 $X=622190 $Y=119440
X1385 1 2 1806 341 1822 1822 1824 342 ICV_16 $T=665160 127840 0 0 $X=664970 $Y=127600
X1386 1 2 1806 343 1842 1842 1824 354 ICV_16 $T=675740 138720 1 0 $X=675550 $Y=135760
X1387 1 2 1835 388 1852 1852 1841 396 ICV_16 $T=679420 165920 1 0 $X=679230 $Y=162960
X1388 1 2 1869 360 1894 1886 1892 356 ICV_16 $T=701500 155040 1 0 $X=701310 $Y=152080
X1389 1 2 1859 360 1900 1903 1868 345 ICV_16 $T=705180 138720 1 0 $X=704990 $Y=135760
X1390 1 2 545 343 1932 1905 537 342 ICV_16 $T=718980 116960 0 0 $X=718790 $Y=116720
X1391 1 2 583 6 594 594 599 19 ICV_17 $T=6900 127840 1 0 $X=6710 $Y=124880
X1392 1 2 586 5 595 595 605 20 ICV_17 $T=6900 138720 1 0 $X=6710 $Y=135760
X1393 1 2 664 6 678 684 683 40 ICV_17 $T=46000 176800 0 0 $X=45810 $Y=176560
X1394 1 2 666 8 679 679 661 21 ICV_17 $T=46460 160480 0 0 $X=46270 $Y=160240
X1395 1 2 761 29 787 787 790 38 ICV_17 $T=98900 144160 0 0 $X=98710 $Y=143920
X1396 1 2 816 27 832 832 824 37 ICV_17 $T=122360 133280 0 0 $X=122170 $Y=133040
X1397 1 2 829 28 869 869 844 40 ICV_17 $T=139840 155040 1 0 $X=139650 $Y=152080
X1398 1 2 1001 176 1023 1023 995 186 ICV_17 $T=228160 171360 1 0 $X=227970 $Y=168400
X1399 1 2 1040 155 1060 1060 1054 150 ICV_17 $T=244720 165920 1 0 $X=244530 $Y=162960
X1400 1 2 1124 176 1150 1150 1118 186 ICV_17 $T=290720 165920 0 0 $X=290530 $Y=165680
X1401 1 2 1148 205 1164 1164 1160 214 ICV_17 $T=299000 138720 0 0 $X=298810 $Y=138480
X1402 1 2 1303 156 1322 1315 1324 166 ICV_17 $T=375360 144160 0 0 $X=375170 $Y=143920
X1403 1 2 1327 155 1283 1334 1284 166 ICV_17 $T=385020 171360 1 0 $X=384830 $Y=168400
X1404 1 2 1301 155 1339 1320 1324 186 ICV_17 $T=386860 155040 1 0 $X=386670 $Y=152080
X1405 1 2 1349 155 1359 1363 1360 162 ICV_17 $T=399740 155040 1 0 $X=399550 $Y=152080
X1406 1 2 1377 153 292 1375 274 188 ICV_17 $T=420440 116960 1 0 $X=420250 $Y=114000
X1407 1 2 1398 193 1433 1433 1410 201 ICV_17 $T=441140 144160 1 0 $X=440950 $Y=141200
X1408 1 2 314 295 1436 1446 319 294 ICV_17 $T=454940 171360 0 0 $X=454750 $Y=171120
X1409 1 2 1548 310 1573 1576 1555 305 ICV_17 $T=519800 122400 0 0 $X=519610 $Y=122160
X1410 1 2 411 281 418 1583 1555 316 ICV_17 $T=525320 116960 1 0 $X=525130 $Y=114000
X1411 1 2 1665 296 1677 1677 1672 304 ICV_17 $T=585580 127840 1 0 $X=585390 $Y=124880
X1412 1 2 1704 281 1713 1713 1719 300 ICV_17 $T=609040 122400 0 0 $X=608850 $Y=122160
X1413 1 2 1704 307 1715 1715 1719 309 ICV_17 $T=609500 122400 1 0 $X=609310 $Y=119440
X1414 1 2 522 400 1773 1773 523 423 ICV_17 $T=637560 176800 1 0 $X=637370 $Y=173840
X1415 1 2 1779 357 1798 1798 1794 356 ICV_17 $T=651820 144160 1 0 $X=651630 $Y=141200
X1416 1 2 1835 378 1855 1855 1841 391 ICV_17 $T=679420 165920 0 0 $X=679230 $Y=165680
X1417 1 2 1871 379 1908 1908 1891 444 ICV_17 $T=706100 171360 1 0 $X=705910 $Y=168400
X1437 1 2 585 28 622 622 602 40 ICV_19 $T=20240 160480 1 0 $X=20050 $Y=157520
X1438 1 2 641 28 672 672 654 40 ICV_19 $T=44620 144160 0 0 $X=44430 $Y=143920
X1439 1 2 701 29 737 737 723 38 ICV_19 $T=76360 160480 0 0 $X=76170 $Y=160240
X1440 1 2 782 8 818 818 798 21 ICV_19 $T=116380 149600 1 0 $X=116190 $Y=146640
X1441 1 2 898 8 910 910 911 21 ICV_19 $T=160540 171360 1 0 $X=160350 $Y=168400
X1442 1 2 998 175 1024 1024 1004 185 ICV_19 $T=228160 127840 1 0 $X=227970 $Y=124880
X1443 1 2 1000 176 1025 1025 1014 186 ICV_19 $T=228160 133280 1 0 $X=227970 $Y=130320
X1444 1 2 1002 178 1026 1031 997 185 ICV_19 $T=228160 149600 1 0 $X=227970 $Y=146640
X1445 1 2 1044 197 1058 1058 1042 203 ICV_19 $T=242880 138720 0 0 $X=242690 $Y=138480
X1446 1 2 1354 156 1370 1370 1372 162 ICV_19 $T=402960 127840 0 0 $X=402770 $Y=127600
X1447 1 2 1398 196 1429 1429 1410 207 ICV_19 $T=439760 138720 0 0 $X=439570 $Y=138480
X1448 1 2 313 307 1465 1463 321 316 ICV_19 $T=459080 116960 0 0 $X=458890 $Y=116720
X1449 1 2 335 298 1508 1508 349 305 ICV_19 $T=481620 176800 1 0 $X=481430 $Y=173840
X1450 1 2 1748 281 1757 1761 1743 316 ICV_19 $T=632040 149600 0 0 $X=631850 $Y=149360
X1451 1 2 1749 298 1759 1759 1763 305 ICV_19 $T=632500 127840 0 0 $X=632310 $Y=127600
X1452 1 2 1733 310 1778 1776 1756 294 ICV_19 $T=641700 138720 1 0 $X=641510 $Y=135760
X1453 1 2 1818 343 1853 1853 1837 354 ICV_19 $T=678500 155040 1 0 $X=678310 $Y=152080
X1454 1 2 1904 338 1950 1956 1920 342 ICV_19 $T=729100 127840 1 0 $X=728910 $Y=124880
X1455 1 2 583 5 590 ICV_20 $T=6900 122400 1 0 $X=6710 $Y=119440
X1456 1 2 587 9 612 ICV_20 $T=10580 176800 1 0 $X=10390 $Y=173840
X1457 1 2 584 27 635 ICV_20 $T=24380 144160 0 0 $X=24190 $Y=143920
X1458 1 2 44 6 648 ICV_20 $T=35880 122400 0 0 $X=35690 $Y=122160
X1459 1 2 46 27 50 ICV_20 $T=36800 176800 0 0 $X=36610 $Y=176560
X1460 1 2 44 29 665 ICV_20 $T=40020 116960 1 0 $X=39830 $Y=114000
X1461 1 2 675 6 692 ICV_20 $T=55200 127840 1 0 $X=55010 $Y=124880
X1462 1 2 726 27 738 ICV_20 $T=78200 144160 1 0 $X=78010 $Y=141200
X1463 1 2 726 8 739 ICV_20 $T=78200 144160 0 0 $X=78010 $Y=143920
X1464 1 2 73 5 770 ICV_20 $T=93380 116960 1 0 $X=93190 $Y=114000
X1465 1 2 73 26 753 ICV_20 $T=94760 122400 1 0 $X=94570 $Y=119440
X1466 1 2 729 28 778 ICV_20 $T=96600 165920 0 0 $X=96410 $Y=165680
X1467 1 2 788 26 800 ICV_20 $T=108100 127840 0 0 $X=107910 $Y=127600
X1468 1 2 788 5 803 ICV_20 $T=108560 116960 0 0 $X=108370 $Y=116720
X1469 1 2 782 9 808 ICV_20 $T=109940 155040 0 0 $X=109750 $Y=154800
X1470 1 2 816 8 831 ICV_20 $T=123280 133280 1 0 $X=123090 $Y=130320
X1471 1 2 829 5 842 ICV_20 $T=129720 155040 0 0 $X=129530 $Y=154800
X1472 1 2 108 27 890 ICV_20 $T=152260 133280 1 0 $X=152070 $Y=130320
X1473 1 2 108 28 893 ICV_20 $T=153640 122400 0 0 $X=153450 $Y=122160
X1474 1 2 108 5 896 ICV_20 $T=154560 116960 0 0 $X=154370 $Y=116720
X1475 1 2 898 27 912 ICV_20 $T=162840 165920 0 0 $X=162650 $Y=165680
X1476 1 2 906 9 916 ICV_20 $T=166060 133280 0 0 $X=165870 $Y=133040
X1477 1 2 876 27 919 ICV_20 $T=166980 155040 1 0 $X=166790 $Y=152080
X1478 1 2 906 6 924 ICV_20 $T=169280 122400 1 0 $X=169090 $Y=119440
X1479 1 2 898 26 935 ICV_20 $T=174340 171360 0 0 $X=174150 $Y=171120
X1480 1 2 928 29 939 ICV_20 $T=177100 138720 1 0 $X=176910 $Y=135760
X1481 1 2 876 26 942 ICV_20 $T=178480 149600 0 0 $X=178290 $Y=149360
X1482 1 2 933 27 953 ICV_20 $T=182620 165920 0 0 $X=182430 $Y=165680
X1483 1 2 160 152 177 ICV_20 $T=223100 165920 1 0 $X=222910 $Y=162960
X1484 1 2 1000 175 1021 ICV_20 $T=228160 138720 1 0 $X=227970 $Y=135760
X1485 1 2 183 178 1043 ICV_20 $T=236440 116960 1 0 $X=236250 $Y=114000
X1486 1 2 1041 205 1068 ICV_20 $T=250240 133280 0 0 $X=250050 $Y=133040
X1487 1 2 1044 213 1062 ICV_20 $T=256220 149600 1 0 $X=256030 $Y=146640
X1488 1 2 1084 176 1119 ICV_20 $T=276920 176800 1 0 $X=276730 $Y=173840
X1489 1 2 1075 213 1113 ICV_20 $T=278300 122400 0 0 $X=278110 $Y=122160
X1490 1 2 1077 213 1125 ICV_20 $T=279220 138720 1 0 $X=279030 $Y=135760
X1491 1 2 1077 194 1129 ICV_20 $T=280600 133280 1 0 $X=280410 $Y=130320
X1492 1 2 1124 178 1135 ICV_20 $T=289800 171360 1 0 $X=289610 $Y=168400
X1493 1 2 1153 153 1162 ICV_20 $T=299460 155040 0 0 $X=299270 $Y=154800
X1494 1 2 1156 153 1169 ICV_20 $T=300840 165920 1 0 $X=300650 $Y=162960
X1495 1 2 1148 204 1179 ICV_20 $T=306360 133280 0 0 $X=306170 $Y=133040
X1496 1 2 1187 204 1207 ICV_20 $T=318780 127840 0 0 $X=318590 $Y=127600
X1497 1 2 1206 178 1230 ICV_20 $T=334420 160480 0 0 $X=334230 $Y=160240
X1498 1 2 1252 155 1265 ICV_20 $T=348680 149600 1 0 $X=348490 $Y=146640
X1499 1 2 1253 179 1291 ICV_20 $T=360640 160480 0 0 $X=360450 $Y=160240
X1500 1 2 255 178 1307 ICV_20 $T=370760 165920 0 0 $X=370570 $Y=165680
X1501 1 2 257 178 260 ICV_20 $T=374900 116960 0 0 $X=374710 $Y=116720
X1502 1 2 1303 154 1319 ICV_20 $T=375360 138720 1 0 $X=375170 $Y=135760
X1503 1 2 1303 153 1323 ICV_20 $T=376740 144160 1 0 $X=376550 $Y=141200
X1504 1 2 1303 178 1342 ICV_20 $T=389160 144160 1 0 $X=388970 $Y=141200
X1505 1 2 1327 176 1356 ICV_20 $T=397900 171360 1 0 $X=397710 $Y=168400
X1506 1 2 1377 176 1393 ICV_20 $T=418600 122400 0 0 $X=418410 $Y=122160
X1507 1 2 160 186 1407 ICV_20 $T=428720 160480 0 0 $X=428530 $Y=160240
X1508 1 2 1377 175 1414 ICV_20 $T=431940 122400 0 0 $X=431750 $Y=122160
X1509 1 2 1396 283 1419 ICV_20 $T=434240 165920 0 0 $X=434050 $Y=165680
X1510 1 2 1395 193 1428 ICV_20 $T=441140 127840 1 0 $X=440950 $Y=124880
X1511 1 2 160 207 323 ICV_20 $T=448500 165920 1 0 $X=448310 $Y=162960
X1512 1 2 1426 296 1470 ICV_20 $T=462300 160480 0 0 $X=462110 $Y=160240
X1513 1 2 160 162 1479 ICV_20 $T=466900 149600 0 0 $X=466710 $Y=149360
X1514 1 2 1467 338 1481 ICV_20 $T=469200 133280 1 0 $X=469010 $Y=130320
X1515 1 2 335 303 1482 ICV_20 $T=469200 171360 0 0 $X=469010 $Y=171120
X1516 1 2 1475 281 1489 ICV_20 $T=471500 171360 1 0 $X=471310 $Y=168400
X1517 1 2 1476 339 1495 ICV_20 $T=473340 122400 1 0 $X=473150 $Y=119440
X1518 1 2 160 344 1498 ICV_20 $T=474720 149600 0 0 $X=474530 $Y=149360
X1519 1 2 1467 357 1517 ICV_20 $T=487600 133280 0 0 $X=487410 $Y=133040
X1520 1 2 1524 380 1544 ICV_20 $T=500020 171360 1 0 $X=499830 $Y=168400
X1521 1 2 1580 399 1591 ICV_20 $T=529920 165920 0 0 $X=529730 $Y=165680
X1522 1 2 424 340 1612 ICV_20 $T=540960 116960 0 0 $X=540770 $Y=116720
X1523 1 2 1606 340 1613 ICV_20 $T=541420 149600 1 0 $X=541230 $Y=146640
X1524 1 2 1626 360 1593 ICV_20 $T=556140 138720 1 0 $X=555950 $Y=135760
X1525 1 2 1626 339 1641 ICV_20 $T=557520 144160 1 0 $X=557330 $Y=141200
X1526 1 2 428 388 1646 ICV_20 $T=561660 176800 1 0 $X=561470 $Y=173840
X1527 1 2 1626 338 1655 ICV_20 $T=569020 144160 0 0 $X=568830 $Y=143920
X1528 1 2 1626 343 1657 ICV_20 $T=569940 133280 0 0 $X=569750 $Y=133040
X1529 1 2 1665 283 1671 ICV_20 $T=585580 133280 1 0 $X=585390 $Y=130320
X1530 1 2 1666 303 1676 ICV_20 $T=586040 144160 1 0 $X=585850 $Y=141200
X1531 1 2 1668 388 1680 ICV_20 $T=588800 165920 1 0 $X=588610 $Y=162960
X1532 1 2 1668 395 1690 ICV_20 $T=595240 160480 0 0 $X=595050 $Y=160240
X1533 1 2 1710 378 1725 ICV_20 $T=613640 165920 1 0 $X=613450 $Y=162960
X1534 1 2 512 486 518 ICV_20 $T=624680 176800 0 0 $X=624490 $Y=176560
X1535 1 2 1733 307 1775 ICV_20 $T=641700 144160 1 0 $X=641510 $Y=141200
X1536 1 2 1733 296 1777 ICV_20 $T=643080 133280 0 0 $X=642890 $Y=133040
X1537 1 2 1755 379 1781 ICV_20 $T=643080 171360 0 0 $X=642890 $Y=171120
X1538 1 2 1748 310 1784 ICV_20 $T=644920 149600 1 0 $X=644730 $Y=146640
X1539 1 2 1779 360 1800 ICV_20 $T=655040 138720 1 0 $X=654850 $Y=135760
X1540 1 2 1795 395 1825 ICV_20 $T=668840 160480 0 0 $X=668650 $Y=160240
X1541 1 2 1871 395 1901 ICV_20 $T=705180 165920 1 0 $X=704990 $Y=162960
X1542 1 2 1869 358 1915 ICV_20 $T=711620 149600 1 0 $X=711430 $Y=146640
X1543 1 2 1919 400 1945 ICV_20 $T=727260 160480 0 0 $X=727070 $Y=160240
X1544 1 2 1919 388 1946 ICV_20 $T=727260 165920 0 0 $X=727070 $Y=165680
X1545 1 2 587 5 607 ICV_21 $T=6900 165920 0 0 $X=6710 $Y=165680
X1546 1 2 587 6 608 ICV_21 $T=6900 171360 1 0 $X=6710 $Y=168400
X1547 1 2 585 29 625 ICV_21 $T=19320 155040 0 0 $X=19130 $Y=154800
X1548 1 2 586 28 628 ICV_21 $T=20240 133280 1 0 $X=20050 $Y=130320
X1549 1 2 641 5 655 ICV_21 $T=34040 144160 0 0 $X=33850 $Y=143920
X1550 1 2 843 26 883 ICV_21 $T=146280 171360 0 0 $X=146090 $Y=171120
X1551 1 2 876 5 930 ICV_21 $T=167900 160480 1 0 $X=167710 $Y=157520
X1552 1 2 932 28 977 ICV_21 $T=193660 127840 1 0 $X=193470 $Y=124880
X1553 1 2 1076 193 1092 ICV_21 $T=261740 155040 1 0 $X=261550 $Y=152080
X1554 1 2 1108 197 1123 ICV_21 $T=275540 149600 0 0 $X=275350 $Y=149360
X1555 1 2 1253 178 1282 ICV_21 $T=356960 155040 1 0 $X=356770 $Y=152080
X1556 1 2 1252 176 1290 ICV_21 $T=357880 138720 0 0 $X=357690 $Y=138480
X1557 1 2 1354 179 1373 ICV_21 $T=402960 138720 0 0 $X=402770 $Y=138480
X1558 1 2 1523 339 1531 ICV_21 $T=495420 133280 0 0 $X=495230 $Y=133040
X1559 1 2 1547 307 1575 ICV_21 $T=518420 155040 0 0 $X=518230 $Y=154800
X1560 1 2 1547 298 1574 ICV_21 $T=518420 160480 0 0 $X=518230 $Y=160240
X1561 1 2 1625 379 1644 ICV_21 $T=557520 171360 1 0 $X=557330 $Y=168400
X1562 1 2 1666 283 1674 ICV_21 $T=582820 144160 0 0 $X=582630 $Y=143920
X1563 1 2 1666 298 1701 ICV_21 $T=598460 144160 1 0 $X=598270 $Y=141200
X1564 1 2 522 382 1808 ICV_21 $T=655500 176800 0 0 $X=655310 $Y=176560
X1565 1 2 1818 358 1828 ICV_21 $T=667920 155040 1 0 $X=667730 $Y=152080
X1566 1 2 1818 339 1854 ICV_21 $T=678960 149600 1 0 $X=678770 $Y=146640
X1567 1 2 583 8 600 600 599 21 ICV_22 $T=6900 122400 0 0 $X=6710 $Y=122160
X1568 1 2 585 9 604 603 602 21 ICV_22 $T=6900 160480 0 0 $X=6710 $Y=160240
X1569 1 2 685 6 706 705 710 37 ICV_22 $T=59800 144160 1 0 $X=59610 $Y=141200
X1570 1 2 726 9 735 735 744 11 ICV_22 $T=75900 138720 0 0 $X=75710 $Y=138480
X1571 1 2 73 29 771 770 754 20 ICV_22 $T=91540 116960 0 0 $X=91350 $Y=116720
X1572 1 2 782 6 825 825 798 19 ICV_22 $T=118220 149600 0 0 $X=118030 $Y=149360
X1573 1 2 837 5 877 877 851 20 ICV_22 $T=143980 144160 1 0 $X=143790 $Y=141200
X1574 1 2 1124 153 1145 1134 1118 188 ICV_22 $T=286580 160480 0 0 $X=286390 $Y=160240
X1575 1 2 230 156 1171 1171 231 162 ICV_22 $T=300380 176800 0 0 $X=300190 $Y=176560
X1576 1 2 225 178 1172 1172 227 189 ICV_22 $T=300840 116960 1 0 $X=300650 $Y=114000
X1577 1 2 1153 176 1195 1195 1163 186 ICV_22 $T=312340 155040 1 0 $X=312150 $Y=152080
X1578 1 2 1252 156 1269 1265 1274 150 ICV_22 $T=347300 149600 0 0 $X=347110 $Y=149360
X1579 1 2 335 307 346 1484 349 320 ICV_22 $T=467360 176800 0 0 $X=467170 $Y=176560
X1580 1 2 1467 341 1485 1481 1487 345 ICV_22 $T=468740 133280 0 0 $X=468550 $Y=133040
X1581 1 2 1606 341 1635 1631 1602 356 ICV_22 $T=552920 149600 0 0 $X=552730 $Y=149360
X1582 1 2 1628 303 1643 1645 1639 309 ICV_22 $T=558440 133280 1 0 $X=558250 $Y=130320
X1583 1 2 1665 303 1693 1693 1672 316 ICV_22 $T=595240 122400 0 0 $X=595050 $Y=122160
X1584 1 2 1916 341 1911 1957 1921 342 ICV_22 $T=729100 144160 1 0 $X=728910 $Y=141200
X1585 1 2 ICV_23 $T=32200 144160 0 0 $X=32010 $Y=143920
X1586 1 2 ICV_23 $T=32200 165920 0 0 $X=32010 $Y=165680
X1587 1 2 ICV_23 $T=60260 149600 0 0 $X=60070 $Y=149360
X1588 1 2 ICV_23 $T=102580 116960 1 0 $X=102390 $Y=114000
X1589 1 2 ICV_23 $T=102580 149600 1 0 $X=102390 $Y=146640
X1590 1 2 ICV_23 $T=116380 138720 0 0 $X=116190 $Y=138480
X1591 1 2 ICV_23 $T=116380 160480 0 0 $X=116190 $Y=160240
X1592 1 2 ICV_23 $T=186760 149600 1 0 $X=186570 $Y=146640
X1593 1 2 ICV_23 $T=186760 165920 1 0 $X=186570 $Y=162960
X1594 1 2 ICV_23 $T=200560 133280 0 0 $X=200370 $Y=133040
X1595 1 2 ICV_23 $T=242880 133280 1 0 $X=242690 $Y=130320
X1596 1 2 ICV_23 $T=242880 149600 1 0 $X=242690 $Y=146640
X1597 1 2 ICV_23 $T=256680 149600 0 0 $X=256490 $Y=149360
X1598 1 2 ICV_23 $T=270940 127840 1 0 $X=270750 $Y=124880
X1599 1 2 ICV_23 $T=284740 155040 0 0 $X=284550 $Y=154800
X1600 1 2 ICV_23 $T=368920 127840 0 0 $X=368730 $Y=127600
X1601 1 2 ICV_23 $T=368920 176800 0 0 $X=368730 $Y=176560
X1602 1 2 ICV_23 $T=383180 116960 1 0 $X=382990 $Y=114000
X1603 1 2 ICV_23 $T=383180 155040 1 0 $X=382990 $Y=152080
X1604 1 2 ICV_23 $T=396980 122400 0 0 $X=396790 $Y=122160
X1605 1 2 ICV_23 $T=425040 149600 0 0 $X=424850 $Y=149360
X1606 1 2 ICV_23 $T=439300 127840 1 0 $X=439110 $Y=124880
X1607 1 2 ICV_23 $T=453100 138720 0 0 $X=452910 $Y=138480
X1608 1 2 ICV_23 $T=453100 144160 0 0 $X=452910 $Y=143920
X1609 1 2 ICV_23 $T=467360 116960 1 0 $X=467170 $Y=114000
X1610 1 2 ICV_23 $T=467360 149600 1 0 $X=467170 $Y=146640
X1611 1 2 ICV_23 $T=467360 160480 1 0 $X=467170 $Y=157520
X1612 1 2 ICV_23 $T=481160 116960 0 0 $X=480970 $Y=116720
X1613 1 2 ICV_23 $T=481160 176800 0 0 $X=480970 $Y=176560
X1614 1 2 ICV_23 $T=495420 165920 1 0 $X=495230 $Y=162960
X1615 1 2 ICV_23 $T=537280 149600 0 0 $X=537090 $Y=149360
X1616 1 2 ICV_23 $T=551540 176800 1 0 $X=551350 $Y=173840
X1617 1 2 ICV_23 $T=579600 171360 1 0 $X=579410 $Y=168400
X1618 1 2 ICV_23 $T=593400 144160 0 0 $X=593210 $Y=143920
X1619 1 2 ICV_23 $T=621460 138720 0 0 $X=621270 $Y=138480
X1620 1 2 ICV_23 $T=677580 176800 0 0 $X=677390 $Y=176560
X1621 1 2 ICV_23 $T=705640 160480 0 0 $X=705450 $Y=160240
X1622 1 2 ICV_24 $T=17940 133280 1 0 $X=17750 $Y=130320
X1623 1 2 ICV_24 $T=31740 171360 0 0 $X=31550 $Y=171120
X1624 1 2 ICV_24 $T=46000 155040 1 0 $X=45810 $Y=152080
X1625 1 2 ICV_24 $T=143980 116960 0 0 $X=143790 $Y=116720
X1626 1 2 ICV_24 $T=228160 144160 0 0 $X=227970 $Y=143920
X1627 1 2 ICV_24 $T=242420 165920 1 0 $X=242230 $Y=162960
X1628 1 2 ICV_24 $T=256220 138720 0 0 $X=256030 $Y=138480
X1629 1 2 ICV_24 $T=340400 144160 0 0 $X=340210 $Y=143920
X1630 1 2 ICV_24 $T=368460 160480 0 0 $X=368270 $Y=160240
X1631 1 2 ICV_24 $T=382720 133280 1 0 $X=382530 $Y=130320
X1632 1 2 ICV_24 $T=396520 144160 0 0 $X=396330 $Y=143920
X1633 1 2 ICV_24 $T=438840 144160 1 0 $X=438650 $Y=141200
X1634 1 2 ICV_24 $T=494960 176800 1 0 $X=494770 $Y=173840
X1635 1 2 ICV_24 $T=523020 116960 1 0 $X=522830 $Y=114000
X1636 1 2 ICV_24 $T=564880 165920 0 0 $X=564690 $Y=165680
X1637 1 2 ICV_24 $T=635260 171360 1 0 $X=635070 $Y=168400
X1638 1 2 ICV_24 $T=677120 127840 0 0 $X=676930 $Y=127600
X1639 1 2 ICV_24 $T=705180 171360 0 0 $X=704990 $Y=171120
X1640 1 2 16 2 599 1 sky130_fd_sc_hd__inv_1 $T=27140 116960 1 0 $X=26950 $Y=114000
X1641 1 2 31 2 15 1 sky130_fd_sc_hd__inv_1 $T=27140 176800 0 0 $X=26950 $Y=176560
X1642 1 2 24 2 615 1 sky130_fd_sc_hd__inv_1 $T=30820 165920 0 0 $X=30630 $Y=165680
X1643 1 2 33 2 605 1 sky130_fd_sc_hd__inv_1 $T=38180 133280 0 0 $X=37990 $Y=133040
X1644 1 2 43 2 51 1 sky130_fd_sc_hd__inv_1 $T=44620 176800 0 0 $X=44430 $Y=176560
X1645 1 2 41 2 649 1 sky130_fd_sc_hd__inv_1 $T=48300 149600 0 0 $X=48110 $Y=149360
X1646 1 2 42 2 654 1 sky130_fd_sc_hd__inv_1 $T=55660 133280 1 0 $X=55470 $Y=130320
X1647 1 2 53 2 661 1 sky130_fd_sc_hd__inv_1 $T=58880 149600 0 0 $X=58690 $Y=149360
X1648 1 2 58 2 683 1 sky130_fd_sc_hd__inv_1 $T=62100 160480 0 0 $X=61910 $Y=160240
X1649 1 2 55 2 695 1 sky130_fd_sc_hd__inv_1 $T=63480 116960 1 0 $X=63290 $Y=114000
X1650 1 2 56 2 710 1 sky130_fd_sc_hd__inv_1 $T=72220 138720 1 0 $X=72030 $Y=135760
X1651 1 2 68 2 66 1 sky130_fd_sc_hd__inv_1 $T=80500 171360 1 0 $X=80310 $Y=168400
X1652 1 2 64 2 723 1 sky130_fd_sc_hd__inv_1 $T=82800 155040 1 0 $X=82610 $Y=152080
X1653 1 2 60 2 741 1 sky130_fd_sc_hd__inv_1 $T=90160 116960 0 0 $X=89970 $Y=116720
X1654 1 2 72 2 70 1 sky130_fd_sc_hd__inv_1 $T=92000 116960 1 0 $X=91810 $Y=114000
X1655 1 2 76 2 744 1 sky130_fd_sc_hd__inv_1 $T=97980 138720 1 0 $X=97790 $Y=135760
X1656 1 2 77 2 754 1 sky130_fd_sc_hd__inv_1 $T=101200 116960 1 0 $X=101010 $Y=114000
X1657 1 2 75 2 760 1 sky130_fd_sc_hd__inv_1 $T=103500 149600 0 0 $X=103310 $Y=149360
X1658 1 2 78 2 752 1 sky130_fd_sc_hd__inv_1 $T=108560 171360 1 0 $X=108370 $Y=168400
X1659 1 2 81 2 84 1 sky130_fd_sc_hd__inv_1 $T=111320 176800 0 0 $X=111130 $Y=176560
X1660 1 2 79 2 783 1 sky130_fd_sc_hd__inv_1 $T=115460 116960 1 0 $X=115270 $Y=114000
X1661 1 2 87 2 824 1 sky130_fd_sc_hd__inv_1 $T=126500 116960 1 0 $X=126310 $Y=114000
X1662 1 2 90 2 790 1 sky130_fd_sc_hd__inv_1 $T=130640 138720 1 0 $X=130450 $Y=135760
X1663 1 2 91 2 798 1 sky130_fd_sc_hd__inv_1 $T=131560 144160 0 0 $X=131370 $Y=143920
X1664 1 2 98 2 814 1 sky130_fd_sc_hd__inv_1 $T=132480 165920 1 0 $X=132290 $Y=162960
X1665 1 2 101 2 93 1 sky130_fd_sc_hd__inv_1 $T=146280 176800 0 0 $X=146090 $Y=176560
X1666 1 2 104 2 844 1 sky130_fd_sc_hd__inv_1 $T=153640 149600 0 0 $X=153450 $Y=149360
X1667 1 2 105 2 112 1 sky130_fd_sc_hd__inv_1 $T=158700 176800 1 0 $X=158510 $Y=173840
X1668 1 2 113 2 858 1 sky130_fd_sc_hd__inv_1 $T=160540 165920 1 0 $X=160350 $Y=162960
X1669 1 2 107 2 899 1 sky130_fd_sc_hd__inv_1 $T=162380 116960 0 0 $X=162190 $Y=116720
X1670 1 2 120 2 882 1 sky130_fd_sc_hd__inv_1 $T=174340 133280 0 0 $X=174150 $Y=133040
X1671 1 2 121 2 927 1 sky130_fd_sc_hd__inv_1 $T=178020 122400 1 0 $X=177830 $Y=119440
X1672 1 2 122 2 117 1 sky130_fd_sc_hd__inv_1 $T=178480 176800 0 0 $X=178290 $Y=176560
X1673 1 2 118 2 911 1 sky130_fd_sc_hd__inv_1 $T=185380 165920 1 0 $X=185190 $Y=162960
X1674 1 2 126 2 892 1 sky130_fd_sc_hd__inv_1 $T=186300 149600 0 0 $X=186110 $Y=149360
X1675 1 2 129 2 951 1 sky130_fd_sc_hd__inv_1 $T=196420 116960 0 0 $X=196230 $Y=116720
X1676 1 2 134 2 950 1 sky130_fd_sc_hd__inv_1 $T=200560 127840 0 0 $X=200370 $Y=127600
X1677 1 2 143 2 128 1 sky130_fd_sc_hd__inv_1 $T=209300 165920 0 0 $X=209110 $Y=165680
X1678 1 2 135 2 969 1 sky130_fd_sc_hd__inv_1 $T=213900 138720 0 0 $X=213710 $Y=138480
X1679 1 2 24 2 995 1 sky130_fd_sc_hd__inv_1 $T=237820 165920 0 0 $X=237630 $Y=165680
X1680 1 2 31 2 163 1 sky130_fd_sc_hd__inv_1 $T=237820 176800 0 0 $X=237630 $Y=176560
X1681 1 2 42 2 1004 1 sky130_fd_sc_hd__inv_1 $T=241500 127840 1 0 $X=241310 $Y=124880
X1682 1 2 22 2 1014 1 sky130_fd_sc_hd__inv_1 $T=241500 133280 1 0 $X=241310 $Y=130320
X1683 1 2 41 2 997 1 sky130_fd_sc_hd__inv_1 $T=241500 149600 1 0 $X=241310 $Y=146640
X1684 1 2 190 2 1042 1 sky130_fd_sc_hd__inv_1 $T=242420 144160 0 0 $X=242230 $Y=143920
X1685 1 2 31 2 1047 1 sky130_fd_sc_hd__inv_1 $T=245180 127840 0 0 $X=244990 $Y=127600
X1686 1 2 43 2 212 1 sky130_fd_sc_hd__inv_1 $T=256680 176800 0 0 $X=256490 $Y=176560
X1687 1 2 17 2 1054 1 sky130_fd_sc_hd__inv_1 $T=264500 160480 0 0 $X=264310 $Y=160240
X1688 1 2 209 2 1094 1 sky130_fd_sc_hd__inv_1 $T=271860 116960 0 0 $X=271670 $Y=116720
X1689 1 2 217 2 1097 1 sky130_fd_sc_hd__inv_1 $T=274160 133280 0 0 $X=273970 $Y=133040
X1690 1 2 52 2 1117 1 sky130_fd_sc_hd__inv_1 $T=283360 149600 1 0 $X=283170 $Y=146640
X1691 1 2 33 2 1118 1 sky130_fd_sc_hd__inv_1 $T=291640 155040 0 0 $X=291450 $Y=154800
X1692 1 2 57 2 229 1 sky130_fd_sc_hd__inv_1 $T=299000 176800 0 0 $X=298810 $Y=176560
X1693 1 2 124 2 1142 1 sky130_fd_sc_hd__inv_1 $T=300840 122400 1 0 $X=300650 $Y=119440
X1694 1 2 81 2 1161 1 sky130_fd_sc_hd__inv_1 $T=304060 165920 0 0 $X=303870 $Y=165680
X1695 1 2 228 2 1160 1 sky130_fd_sc_hd__inv_1 $T=304980 133280 0 0 $X=304790 $Y=133040
X1696 1 2 53 2 1163 1 sky130_fd_sc_hd__inv_1 $T=308200 149600 1 0 $X=308010 $Y=146640
X1697 1 2 56 2 1191 1 sky130_fd_sc_hd__inv_1 $T=319700 138720 1 0 $X=319510 $Y=135760
X1698 1 2 76 2 233 1 sky130_fd_sc_hd__inv_1 $T=327060 116960 1 0 $X=326870 $Y=114000
X1699 1 2 237 2 1205 1 sky130_fd_sc_hd__inv_1 $T=332580 122400 0 0 $X=332390 $Y=122160
X1700 1 2 64 2 1218 1 sky130_fd_sc_hd__inv_1 $T=333500 149600 0 0 $X=333310 $Y=149360
X1701 1 2 234 2 239 1 sky130_fd_sc_hd__inv_1 $T=342700 176800 0 0 $X=342510 $Y=176560
X1702 1 2 98 2 244 1 sky130_fd_sc_hd__inv_1 $T=350980 171360 1 0 $X=350790 $Y=168400
X1703 1 2 91 2 1261 1 sky130_fd_sc_hd__inv_1 $T=355120 138720 1 0 $X=354930 $Y=135760
X1704 1 2 121 2 1272 1 sky130_fd_sc_hd__inv_1 $T=368920 116960 0 0 $X=368730 $Y=116720
X1705 1 2 113 2 1274 1 sky130_fd_sc_hd__inv_1 $T=368920 138720 0 0 $X=368730 $Y=138480
X1706 1 2 122 2 258 1 sky130_fd_sc_hd__inv_1 $T=379040 176800 1 0 $X=378850 $Y=173840
X1707 1 2 105 2 1324 1 sky130_fd_sc_hd__inv_1 $T=385480 155040 1 0 $X=385290 $Y=152080
X1708 1 2 120 2 1326 1 sky130_fd_sc_hd__inv_1 $T=389160 138720 1 0 $X=388970 $Y=135760
X1709 1 2 137 2 259 1 sky130_fd_sc_hd__inv_1 $T=395600 122400 0 0 $X=395410 $Y=122160
X1710 1 2 75 2 1360 1 sky130_fd_sc_hd__inv_1 $T=407560 155040 0 0 $X=407370 $Y=154800
X1711 1 2 272 2 1372 1 sky130_fd_sc_hd__inv_1 $T=414920 133280 1 0 $X=414730 $Y=130320
X1712 1 2 143 2 274 1 sky130_fd_sc_hd__inv_1 $T=416300 116960 0 0 $X=416110 $Y=116720
X1713 1 2 266 2 1367 1 sky130_fd_sc_hd__inv_1 $T=420440 160480 1 0 $X=420250 $Y=157520
X1714 1 2 136 2 293 1 sky130_fd_sc_hd__inv_1 $T=430100 122400 1 0 $X=429910 $Y=119440
X1715 1 2 266 2 1400 1 sky130_fd_sc_hd__inv_1 $T=431020 127840 0 0 $X=430830 $Y=127600
X1716 1 2 289 2 302 1 sky130_fd_sc_hd__inv_1 $T=444360 165920 0 0 $X=444170 $Y=165680
X1717 1 2 322 2 1452 1 sky130_fd_sc_hd__inv_1 $T=467360 133280 0 0 $X=467170 $Y=133040
X1718 1 2 312 2 319 1 sky130_fd_sc_hd__inv_1 $T=467820 171360 0 0 $X=467630 $Y=171120
X1719 1 2 308 2 1449 1 sky130_fd_sc_hd__inv_1 $T=469200 160480 1 0 $X=469010 $Y=157520
X1720 1 2 330 2 1473 1 sky130_fd_sc_hd__inv_1 $T=476560 144160 1 0 $X=476370 $Y=141200
X1721 1 2 333 2 1487 1 sky130_fd_sc_hd__inv_1 $T=482080 138720 1 0 $X=481890 $Y=135760
X1722 1 2 337 2 361 1 sky130_fd_sc_hd__inv_1 $T=486680 116960 1 0 $X=486490 $Y=114000
X1723 1 2 352 2 1490 1 sky130_fd_sc_hd__inv_1 $T=492660 165920 0 0 $X=492470 $Y=165680
X1724 1 2 336 2 1501 1 sky130_fd_sc_hd__inv_1 $T=499100 127840 0 0 $X=498910 $Y=127600
X1725 1 2 352 2 1534 1 sky130_fd_sc_hd__inv_1 $T=509220 144160 0 0 $X=509030 $Y=143920
X1726 1 2 366 2 386 1 sky130_fd_sc_hd__inv_1 $T=511060 171360 0 0 $X=510870 $Y=171120
X1727 1 2 336 2 1555 1 sky130_fd_sc_hd__inv_1 $T=518420 122400 0 0 $X=518230 $Y=122160
X1728 1 2 306 2 393 1 sky130_fd_sc_hd__inv_1 $T=522560 176800 0 0 $X=522370 $Y=176560
X1729 1 2 384 2 1538 1 sky130_fd_sc_hd__inv_1 $T=529000 155040 0 0 $X=528810 $Y=154800
X1730 1 2 350 2 1600 1 sky130_fd_sc_hd__inv_1 $T=541880 165920 1 0 $X=541690 $Y=162960
X1731 1 2 308 2 1604 1 sky130_fd_sc_hd__inv_1 $T=546480 127840 0 0 $X=546290 $Y=127600
X1732 1 2 312 2 433 1 sky130_fd_sc_hd__inv_1 $T=548780 116960 0 0 $X=548590 $Y=116720
X1733 1 2 410 2 1602 1 sky130_fd_sc_hd__inv_1 $T=551540 149600 0 0 $X=551350 $Y=149360
X1734 1 2 421 2 440 1 sky130_fd_sc_hd__inv_1 $T=552000 176800 0 0 $X=551810 $Y=176560
X1735 1 2 430 2 1596 1 sky130_fd_sc_hd__inv_1 $T=560280 138720 0 0 $X=560090 $Y=138480
X1736 1 2 434 2 1638 1 sky130_fd_sc_hd__inv_1 $T=563500 165920 0 0 $X=563310 $Y=165680
X1737 1 2 447 2 1682 1 sky130_fd_sc_hd__inv_1 $T=598920 165920 1 0 $X=598730 $Y=162960
X1738 1 2 489 2 1679 1 sky130_fd_sc_hd__inv_1 $T=602140 144160 0 0 $X=601950 $Y=143920
X1739 1 2 479 2 491 1 sky130_fd_sc_hd__inv_1 $T=602600 176800 1 0 $X=602410 $Y=173840
X1740 1 2 472 2 1672 1 sky130_fd_sc_hd__inv_1 $T=609500 133280 1 0 $X=609310 $Y=130320
X1741 1 2 501 2 503 1 sky130_fd_sc_hd__inv_1 $T=623300 176800 0 0 $X=623110 $Y=176560
X1742 1 2 495 2 488 1 sky130_fd_sc_hd__inv_1 $T=627440 116960 0 0 $X=627250 $Y=116720
X1743 1 2 508 2 1707 1 sky130_fd_sc_hd__inv_1 $T=630660 149600 0 0 $X=630470 $Y=149360
X1744 1 2 490 2 1719 1 sky130_fd_sc_hd__inv_1 $T=631120 127840 0 0 $X=630930 $Y=127600
X1745 1 2 499 2 1722 1 sky130_fd_sc_hd__inv_1 $T=633880 171360 1 0 $X=633690 $Y=168400
X1746 1 2 510 2 520 1 sky130_fd_sc_hd__inv_1 $T=635260 176800 1 0 $X=635070 $Y=173840
X1747 1 2 429 2 523 1 sky130_fd_sc_hd__inv_1 $T=642160 176800 0 0 $X=641970 $Y=176560
X1748 1 2 504 2 1756 1 sky130_fd_sc_hd__inv_1 $T=651360 138720 0 0 $X=651170 $Y=138480
X1749 1 2 404 2 1794 1 sky130_fd_sc_hd__inv_1 $T=655960 144160 0 0 $X=655770 $Y=143920
X1750 1 2 511 2 517 1 sky130_fd_sc_hd__inv_1 $T=658720 116960 0 0 $X=658530 $Y=116720
X1751 1 2 432 2 1824 1 sky130_fd_sc_hd__inv_1 $T=674360 138720 1 0 $X=674170 $Y=135760
X1752 1 2 406 2 1804 1 sky130_fd_sc_hd__inv_1 $T=676660 160480 0 0 $X=676470 $Y=160240
X1753 1 2 490 2 531 1 sky130_fd_sc_hd__inv_1 $T=685860 122400 0 0 $X=685670 $Y=122160
X1754 1 2 479 2 1841 1 sky130_fd_sc_hd__inv_1 $T=691380 165920 1 0 $X=691190 $Y=162960
X1755 1 2 461 2 1837 1 sky130_fd_sc_hd__inv_1 $T=691840 155040 1 0 $X=691650 $Y=152080
X1756 1 2 472 2 1866 1 sky130_fd_sc_hd__inv_1 $T=693680 133280 0 0 $X=693490 $Y=133040
X1757 1 2 509 2 1868 1 sky130_fd_sc_hd__inv_1 $T=701040 144160 1 0 $X=700850 $Y=141200
X1758 1 2 510 2 1891 1 sky130_fd_sc_hd__inv_1 $T=715760 171360 0 0 $X=715570 $Y=171120
X1759 1 2 508 2 1892 1 sky130_fd_sc_hd__inv_1 $T=717600 155040 1 0 $X=717410 $Y=152080
X1760 1 2 504 2 1920 1 sky130_fd_sc_hd__inv_1 $T=719900 133280 1 0 $X=719710 $Y=130320
X1761 1 2 489 2 1921 1 sky130_fd_sc_hd__inv_1 $T=719900 149600 1 0 $X=719710 $Y=146640
X1762 1 2 502 2 1928 1 sky130_fd_sc_hd__inv_1 $T=725880 160480 1 0 $X=725690 $Y=157520
X1763 1 2 468 2 546 1 sky130_fd_sc_hd__inv_1 $T=726340 176800 0 0 $X=726150 $Y=176560
X1764 1 2 511 2 549 1 sky130_fd_sc_hd__inv_1 $T=729100 116960 1 0 $X=728910 $Y=114000
X1765 1 2 513 2 1914 1 sky130_fd_sc_hd__inv_1 $T=729100 138720 1 0 $X=728910 $Y=135760
X1766 1 2 590 599 20 ICV_26 $T=14720 122400 1 0 $X=14530 $Y=119440
X1767 1 2 591 589 20 ICV_26 $T=15180 149600 1 0 $X=14990 $Y=146640
X1768 1 2 625 602 38 ICV_26 $T=28980 160480 0 0 $X=28790 $Y=160240
X1769 1 2 636 615 37 ICV_26 $T=31740 171360 1 0 $X=31550 $Y=168400
X1770 1 2 655 654 20 ICV_26 $T=43240 144160 1 0 $X=43050 $Y=141200
X1771 1 2 698 661 20 ICV_26 $T=63480 160480 0 0 $X=63290 $Y=160240
X1772 1 2 767 754 11 ICV_26 $T=99360 138720 1 0 $X=99170 $Y=135760
X1773 1 2 784 760 11 ICV_26 $T=104420 165920 1 0 $X=104230 $Y=162960
X1774 1 2 826 790 20 ICV_26 $T=126960 144160 0 0 $X=126770 $Y=143920
X1775 1 2 839 814 21 ICV_26 $T=132480 165920 0 0 $X=132290 $Y=165680
X1776 1 2 948 951 38 ICV_26 $T=188600 122400 1 0 $X=188410 $Y=119440
X1777 1 2 980 944 40 ICV_26 $T=205160 160480 0 0 $X=204970 $Y=160240
X1778 1 2 993 995 150 ICV_26 $T=210680 165920 0 0 $X=210490 $Y=165680
X1779 1 2 1105 1096 207 ICV_26 $T=275080 160480 0 0 $X=274890 $Y=160240
X1780 1 2 1123 1117 203 ICV_26 $T=284740 149600 1 0 $X=284550 $Y=146640
X1781 1 2 1125 1097 211 ICV_26 $T=286580 138720 0 0 $X=286390 $Y=138480
X1782 1 2 1170 1161 188 ICV_26 $T=307740 176800 1 0 $X=307550 $Y=173840
X1783 1 2 1219 1205 216 ICV_26 $T=331200 127840 1 0 $X=331010 $Y=124880
X1784 1 2 1229 1191 188 ICV_26 $T=337640 133280 0 0 $X=337450 $Y=133040
X1785 1 2 1233 1205 203 ICV_26 $T=342700 127840 0 0 $X=342510 $Y=127600
X1786 1 2 1236 1218 185 ICV_26 $T=342700 149600 0 0 $X=342510 $Y=149360
X1787 1 2 1273 1261 167 ICV_26 $T=356960 133280 1 0 $X=356770 $Y=130320
X1788 1 2 1278 1272 185 ICV_26 $T=358800 127840 0 0 $X=358610 $Y=127600
X1789 1 2 1298 1274 167 ICV_26 $T=370760 144160 0 0 $X=370570 $Y=143920
X1790 1 2 1311 259 162 ICV_26 $T=379960 127840 1 0 $X=379770 $Y=124880
X1791 1 2 1329 259 166 ICV_26 $T=386400 133280 0 0 $X=386210 $Y=133040
X1792 1 2 1338 1284 167 ICV_26 $T=393760 165920 0 0 $X=393570 $Y=165680
X1793 1 2 1340 1284 185 ICV_26 $T=394220 176800 1 0 $X=394030 $Y=173840
X1794 1 2 1376 274 150 ICV_26 $T=415840 127840 1 0 $X=415650 $Y=124880
X1795 1 2 1416 293 162 ICV_26 $T=441600 116960 0 0 $X=441410 $Y=116720
X1796 1 2 1494 1501 342 ICV_26 $T=481160 127840 1 0 $X=480970 $Y=124880
X1797 1 2 1502 1487 351 ICV_26 $T=483000 133280 0 0 $X=482810 $Y=133040
X1798 1 2 1533 1534 351 ICV_26 $T=506000 133280 0 0 $X=505810 $Y=133040
X1799 1 2 1611 433 354 ICV_26 $T=547860 122400 1 0 $X=547670 $Y=119440
X1800 1 2 1620 1596 356 ICV_26 $T=552460 133280 0 0 $X=552270 $Y=133040
X1801 1 2 1644 1638 444 ICV_26 $T=567180 171360 0 0 $X=566990 $Y=171120
X1802 1 2 1661 1639 305 ICV_26 $T=581440 122400 1 0 $X=581250 $Y=119440
X1803 1 2 1671 1672 294 ICV_26 $T=590180 133280 0 0 $X=589990 $Y=133040
X1804 1 2 1676 1679 316 ICV_26 $T=593860 144160 1 0 $X=593670 $Y=141200
X1805 1 2 498 488 325 ICV_26 $T=609500 116960 1 0 $X=609310 $Y=114000
X1806 1 2 1712 503 455 ICV_26 $T=615940 176800 1 0 $X=615750 $Y=173840
X1807 1 2 506 503 451 ICV_26 $T=618240 176800 0 0 $X=618050 $Y=176560
X1808 1 2 1760 1743 305 ICV_26 $T=640320 155040 1 0 $X=640130 $Y=152080
X1809 1 2 1768 1771 396 ICV_26 $T=643540 165920 0 0 $X=643350 $Y=165680
X1810 1 2 1789 1771 409 ICV_26 $T=654120 165920 0 0 $X=653930 $Y=165680
X1811 1 2 530 531 344 ICV_26 $T=665620 116960 1 0 $X=665430 $Y=114000
X1812 1 2 1816 1794 342 ICV_26 $T=669760 138720 1 0 $X=669570 $Y=135760
X1813 1 2 1826 1804 407 ICV_26 $T=674360 165920 0 0 $X=674170 $Y=165680
X1814 1 2 1893 1892 345 ICV_26 $T=707480 155040 0 0 $X=707290 $Y=154800
X1815 1 2 1911 1914 342 ICV_26 $T=715760 138720 0 0 $X=715570 $Y=138480
X1816 1 2 1943 1914 345 ICV_26 $T=730480 133280 0 0 $X=730290 $Y=133040
X1817 1 2 584 9 588 17 589 ICV_27 $T=15640 144160 0 0 $X=15450 $Y=143920
X1818 1 2 585 27 624 22 602 ICV_27 $T=22540 155040 1 0 $X=22350 $Y=152080
X1819 1 2 100 5 867 99 103 ICV_27 $T=141680 116960 1 0 $X=141490 $Y=114000
X1820 1 2 837 26 880 102 851 ICV_27 $T=149040 138720 0 0 $X=148850 $Y=138480
X1821 1 2 933 28 980 136 944 ICV_27 $T=200100 160480 1 0 $X=199910 $Y=157520
X1822 1 2 1076 197 1088 72 1096 ICV_27 $T=264500 155040 0 0 $X=264310 $Y=154800
X1823 1 2 1084 153 1104 58 1102 ICV_27 $T=268640 165920 0 0 $X=268450 $Y=165680
X1824 1 2 1206 153 1220 68 1214 ICV_27 $T=325680 160480 0 0 $X=325490 $Y=160240
X1825 1 2 1253 154 1270 78 1276 ICV_27 $T=350060 155040 0 0 $X=349870 $Y=154800
X1826 1 2 1327 154 1338 118 1284 ICV_27 $T=391920 165920 1 0 $X=391730 $Y=162960
X1827 1 2 1398 205 1412 122 1410 ICV_27 $T=431020 138720 0 0 $X=430830 $Y=138480
X1828 1 2 1628 296 1660 461 1639 ICV_27 $T=572240 127840 1 0 $X=572050 $Y=124880
X1829 1 2 1748 296 1783 509 1743 ICV_27 $T=644920 155040 1 0 $X=644730 $Y=152080
X1830 1 2 1749 296 1792 513 1763 ICV_27 $T=648600 127840 1 0 $X=648410 $Y=124880
X1831 1 2 1755 380 1789 501 1771 ICV_27 $T=649060 171360 1 0 $X=648870 $Y=168400
X1832 1 2 538 343 1858 495 537 ICV_27 $T=685860 116960 0 0 $X=685670 $Y=116720
X1833 1 2 586 6 598 ICV_28 $T=6900 138720 0 0 $X=6710 $Y=138480
X1834 1 2 586 27 621 ICV_28 $T=20240 138720 1 0 $X=20050 $Y=135760
X1835 1 2 583 26 623 ICV_28 $T=20700 122400 0 0 $X=20510 $Y=122160
X1836 1 2 587 28 633 ICV_28 $T=22540 171360 0 0 $X=22350 $Y=171120
X1837 1 2 639 26 646 ICV_28 $T=33580 160480 1 0 $X=33390 $Y=157520
X1838 1 2 639 29 657 ICV_28 $T=35420 165920 1 0 $X=35230 $Y=162960
X1839 1 2 641 8 663 ICV_28 $T=38180 138720 1 0 $X=37990 $Y=135760
X1840 1 2 44 28 669 ICV_28 $T=43700 122400 0 0 $X=43510 $Y=122160
X1841 1 2 666 9 686 ICV_28 $T=49680 149600 0 0 $X=49490 $Y=149360
X1842 1 2 675 9 689 ICV_28 $T=52440 127840 0 0 $X=52250 $Y=127600
X1843 1 2 666 5 698 ICV_28 $T=55660 160480 1 0 $X=55470 $Y=157520
X1844 1 2 701 6 717 ICV_28 $T=66240 155040 1 0 $X=66050 $Y=152080
X1845 1 2 701 27 720 ICV_28 $T=66700 165920 1 0 $X=66510 $Y=162960
X1846 1 2 702 26 734 ICV_28 $T=76360 122400 1 0 $X=76170 $Y=119440
X1847 1 2 729 5 792 ICV_28 $T=100280 171360 0 0 $X=100090 $Y=171120
X1848 1 2 843 6 856 ICV_28 $T=136620 176800 1 0 $X=136430 $Y=173840
X1849 1 2 106 29 886 ICV_28 $T=149500 176800 1 0 $X=149310 $Y=173840
X1850 1 2 108 26 889 ICV_28 $T=150880 127840 1 0 $X=150690 $Y=124880
X1851 1 2 876 8 900 ICV_28 $T=153640 155040 0 0 $X=153450 $Y=154800
X1852 1 2 941 6 958 ICV_28 $T=183080 144160 0 0 $X=182890 $Y=143920
X1853 1 2 1002 175 1031 ICV_28 $T=228620 155040 1 0 $X=228430 $Y=152080
X1854 1 2 215 155 221 ICV_28 $T=262660 116960 0 0 $X=262470 $Y=116720
X1855 1 2 1076 205 1099 ICV_28 $T=265880 160480 0 0 $X=265690 $Y=160240
X1856 1 2 1084 154 1100 ICV_28 $T=265880 171360 0 0 $X=265690 $Y=171120
X1857 1 2 1124 175 1151 ICV_28 $T=290720 171360 0 0 $X=290530 $Y=171120
X1858 1 2 1192 154 1235 ICV_28 $T=333040 138720 0 0 $X=332850 $Y=138480
X1859 1 2 1208 176 1246 ICV_28 $T=336260 155040 1 0 $X=336070 $Y=152080
X1860 1 2 243 156 1259 ICV_28 $T=346840 165920 0 0 $X=346650 $Y=165680
X1861 1 2 1253 155 1286 ICV_28 $T=358800 155040 0 0 $X=358610 $Y=154800
X1862 1 2 1248 153 1293 ICV_28 $T=359720 133280 0 0 $X=359530 $Y=133040
X1863 1 2 255 153 1309 ICV_28 $T=370760 160480 0 0 $X=370570 $Y=160240
X1864 1 2 255 176 1316 ICV_28 $T=372600 171360 1 0 $X=372410 $Y=168400
X1865 1 2 257 156 261 ICV_28 $T=373980 116960 1 0 $X=373790 $Y=114000
X1866 1 2 1303 175 1325 ICV_28 $T=377200 133280 0 0 $X=377010 $Y=133040
X1867 1 2 1327 178 1285 ICV_28 $T=385020 176800 1 0 $X=384830 $Y=173840
X1868 1 2 160 203 273 ICV_28 $T=394220 160480 1 0 $X=394030 $Y=157520
X1869 1 2 269 179 1375 ICV_28 $T=407100 116960 0 0 $X=406910 $Y=116720
X1870 1 2 1354 175 1389 ICV_28 $T=413540 138720 0 0 $X=413350 $Y=138480
X1871 1 2 160 216 286 ICV_28 $T=417220 171360 1 0 $X=417030 $Y=168400
X1872 1 2 1377 156 1416 ICV_28 $T=431480 122400 1 0 $X=431290 $Y=119440
X1873 1 2 1396 307 1413 ICV_28 $T=436540 160480 0 0 $X=436350 $Y=160240
X1874 1 2 1475 310 1505 ICV_28 $T=480240 160480 1 0 $X=480050 $Y=157520
X1875 1 2 1475 307 1511 ICV_28 $T=483000 165920 0 0 $X=482810 $Y=165680
X1876 1 2 1476 358 1520 ICV_28 $T=487140 122400 0 0 $X=486950 $Y=122160
X1877 1 2 1523 340 1533 ICV_28 $T=497260 133280 1 0 $X=497070 $Y=130320
X1878 1 2 1548 281 1563 ICV_28 $T=510140 122400 1 0 $X=509950 $Y=119440
X1879 1 2 1547 281 1571 ICV_28 $T=518420 149600 0 0 $X=518230 $Y=149360
X1880 1 2 428 378 439 ICV_28 $T=543260 171360 0 0 $X=543070 $Y=171120
X1881 1 2 1665 295 1692 ICV_28 $T=595240 133280 0 0 $X=595050 $Y=133040
X1882 1 2 484 486 492 ICV_28 $T=595240 176800 0 0 $X=595050 $Y=176560
X1883 1 2 1733 281 1754 ICV_28 $T=626980 144160 1 0 $X=626790 $Y=141200
X1884 1 2 1748 307 1780 ICV_28 $T=641700 155040 0 0 $X=641510 $Y=154800
X1885 1 2 1818 340 1831 ICV_28 $T=669760 149600 1 0 $X=669570 $Y=146640
X1886 1 2 1844 360 1862 ICV_28 $T=684020 127840 1 0 $X=683830 $Y=124880
X1887 1 2 538 360 1879 ICV_28 $T=693680 122400 1 0 $X=693490 $Y=119440
X1888 1 2 538 340 1880 ICV_28 $T=694600 116960 0 0 $X=694410 $Y=116720
X1889 1 2 1859 343 1898 ICV_28 $T=702420 144160 1 0 $X=702230 $Y=141200
X1890 1 2 586 9 601 ICV_29 $T=6900 144160 1 0 $X=6710 $Y=141200
X1891 1 2 585 8 603 ICV_29 $T=6900 160480 1 0 $X=6710 $Y=157520
X1892 1 2 675 8 715 ICV_29 $T=63020 127840 1 0 $X=62830 $Y=124880
X1893 1 2 62 28 67 ICV_29 $T=69460 176800 0 0 $X=69270 $Y=176560
X1894 1 2 745 28 757 ICV_29 $T=84180 155040 1 0 $X=83990 $Y=152080
X1895 1 2 73 8 772 ICV_29 $T=92000 133280 1 0 $X=91810 $Y=130320
X1896 1 2 788 28 805 ICV_29 $T=106720 122400 0 0 $X=106530 $Y=122160
X1897 1 2 761 8 799 ICV_29 $T=108560 144160 1 0 $X=108370 $Y=141200
X1898 1 2 816 28 833 ICV_29 $T=122360 122400 0 0 $X=122170 $Y=122160
X1899 1 2 791 28 840 ICV_29 $T=125580 171360 0 0 $X=125390 $Y=171120
X1900 1 2 100 27 861 ICV_29 $T=135240 133280 0 0 $X=135050 $Y=133040
X1901 1 2 108 29 888 ICV_29 $T=150420 116960 1 0 $X=150230 $Y=114000
X1902 1 2 933 29 947 ICV_29 $T=178480 160480 1 0 $X=178290 $Y=157520
X1903 1 2 1075 205 1112 ICV_29 $T=273240 116960 0 0 $X=273050 $Y=116720
X1904 1 2 1108 194 1114 ICV_29 $T=276000 144160 0 0 $X=275810 $Y=143920
X1905 1 2 243 154 1260 ICV_29 $T=346840 171360 0 0 $X=346650 $Y=171120
X1906 1 2 1312 156 1311 ICV_29 $T=378120 122400 0 0 $X=377930 $Y=122160
X1907 1 2 269 156 1358 ICV_29 $T=398820 122400 0 0 $X=398630 $Y=122160
X1908 1 2 1350 153 1368 ICV_29 $T=400660 165920 1 0 $X=400470 $Y=162960
X1909 1 2 1350 156 1364 ICV_29 $T=402960 165920 0 0 $X=402770 $Y=165680
X1910 1 2 160 150 1417 ICV_29 $T=431020 160480 1 0 $X=430830 $Y=157520
X1911 1 2 1426 283 1447 ICV_29 $T=447580 160480 1 0 $X=447390 $Y=157520
X1912 1 2 160 210 329 ICV_29 $T=455400 149600 1 0 $X=455210 $Y=146640
X1913 1 2 160 211 331 ICV_29 $T=456320 165920 1 0 $X=456130 $Y=162960
X1914 1 2 1475 295 1491 ICV_29 $T=470580 160480 1 0 $X=470390 $Y=157520
X1915 1 2 1467 343 1493 ICV_29 $T=471040 127840 0 0 $X=470850 $Y=127600
X1916 1 2 1467 360 1513 ICV_29 $T=483460 138720 1 0 $X=483270 $Y=135760
X1917 1 2 1524 378 1539 ICV_29 $T=497260 165920 1 0 $X=497070 $Y=162960
X1918 1 2 1548 307 1564 ICV_29 $T=511060 116960 0 0 $X=510870 $Y=116720
X1919 1 2 477 298 485 ICV_29 $T=588800 116960 1 0 $X=588610 $Y=114000
X1920 1 2 1733 283 1776 ICV_29 $T=640320 138720 0 0 $X=640130 $Y=138480
X1921 1 2 1779 340 1802 ICV_29 $T=652740 138720 0 0 $X=652550 $Y=138480
X1922 1 2 1779 358 1803 ICV_29 $T=652740 149600 1 0 $X=652550 $Y=146640
X1923 1 2 1818 341 1856 ICV_29 $T=679420 149600 0 0 $X=679230 $Y=149360
X1924 1 2 1818 338 1857 ICV_29 $T=679420 155040 0 0 $X=679230 $Y=154800
X1925 1 2 588 589 11 604 602 11 ICV_30 $T=11500 165920 1 0 $X=11310 $Y=162960
X1926 1 2 609 599 11 601 605 11 ICV_30 $T=17020 127840 0 0 $X=16830 $Y=127600
X1927 1 2 617 589 32 627 589 38 ICV_30 $T=25300 127840 0 0 $X=25110 $Y=127600
X1928 1 2 633 615 40 630 615 38 ICV_30 $T=34040 171360 0 0 $X=33850 $Y=171120
X1929 1 2 644 48 32 648 48 19 ICV_30 $T=39560 122400 1 0 $X=39370 $Y=119440
X1930 1 2 663 654 21 670 48 11 ICV_30 $T=48300 138720 1 0 $X=48110 $Y=135760
X1931 1 2 658 649 20 651 649 11 ICV_30 $T=48300 165920 0 0 $X=48110 $Y=165680
X1932 1 2 699 661 32 686 661 11 ICV_30 $T=64400 149600 0 0 $X=64210 $Y=149360
X1933 1 2 707 710 21 711 710 40 ICV_30 $T=69920 144160 0 0 $X=69730 $Y=143920
X1934 1 2 724 723 40 721 723 11 ICV_30 $T=77280 165920 1 0 $X=77090 $Y=162960
X1935 1 2 728 723 21 736 723 20 ICV_30 $T=81420 155040 0 0 $X=81230 $Y=154800
X1936 1 2 731 741 38 734 741 32 ICV_30 $T=86480 122400 1 0 $X=86290 $Y=119440
X1937 1 2 748 66 20 74 66 11 ICV_30 $T=90160 176800 0 0 $X=89970 $Y=176560
X1938 1 2 763 760 20 779 760 19 ICV_30 $T=101660 155040 0 0 $X=101470 $Y=154800
X1939 1 2 789 790 40 786 790 19 ICV_30 $T=108100 138720 0 0 $X=107910 $Y=138480
X1940 1 2 808 798 11 815 814 37 ICV_30 $T=120060 160480 0 0 $X=119870 $Y=160240
X1941 1 2 800 783 32 92 85 95 ICV_30 $T=120520 122400 1 0 $X=120330 $Y=119440
X1942 1 2 822 814 32 835 814 11 ICV_30 $T=128340 160480 0 0 $X=128150 $Y=160240
X1943 1 2 838 824 32 830 824 11 ICV_30 $T=132480 127840 0 0 $X=132290 $Y=127600
X1944 1 2 842 844 20 859 858 38 ICV_30 $T=137540 160480 0 0 $X=137350 $Y=160240
X1945 1 2 860 103 21 874 103 11 ICV_30 $T=146280 133280 0 0 $X=146090 $Y=133040
X1946 1 2 862 858 20 875 858 11 ICV_30 $T=146280 160480 0 0 $X=146090 $Y=160240
X1947 1 2 878 844 38 872 844 11 ICV_30 $T=154560 160480 0 0 $X=154370 $Y=160240
X1948 1 2 881 882 11 891 892 11 ICV_30 $T=155480 149600 0 0 $X=155290 $Y=149360
X1949 1 2 883 858 32 901 112 19 ICV_30 $T=160540 176800 1 0 $X=160350 $Y=173840
X1950 1 2 896 899 20 888 899 38 ICV_30 $T=161920 116960 1 0 $X=161730 $Y=114000
X1951 1 2 903 892 19 908 892 38 ICV_30 $T=163760 149600 0 0 $X=163570 $Y=149360
X1952 1 2 116 117 38 913 911 40 ICV_30 $T=169740 176800 1 0 $X=169550 $Y=173840
X1953 1 2 912 911 37 914 911 11 ICV_30 $T=174340 165920 0 0 $X=174150 $Y=165680
X1954 1 2 920 882 21 921 882 37 ICV_30 $T=174800 144160 0 0 $X=174610 $Y=143920
X1955 1 2 940 950 19 939 950 38 ICV_30 $T=188600 138720 1 0 $X=188410 $Y=135760
X1956 1 2 959 128 38 953 944 37 ICV_30 $T=191360 165920 0 0 $X=191170 $Y=165680
X1957 1 2 971 128 19 139 142 32 ICV_30 $T=196880 176800 1 0 $X=196690 $Y=173840
X1958 1 2 976 951 19 982 951 11 ICV_30 $T=203320 122400 0 0 $X=203130 $Y=122160
X1959 1 2 970 944 19 994 944 11 ICV_30 $T=207000 171360 1 0 $X=206810 $Y=168400
X1960 1 2 1021 1014 185 1038 1014 189 ICV_30 $T=235980 144160 1 0 $X=235790 $Y=141200
X1961 1 2 198 195 188 1045 195 162 ICV_30 $T=245640 116960 1 0 $X=245450 $Y=114000
X1962 1 2 1052 1054 186 1050 1054 188 ICV_30 $T=249780 171360 0 0 $X=249590 $Y=171120
X1963 1 2 1071 1054 162 1073 1054 167 ICV_30 $T=258980 165920 1 0 $X=258790 $Y=162960
X1964 1 2 1087 1094 216 1106 1094 207 ICV_30 $T=272780 127840 1 0 $X=272590 $Y=124880
X1965 1 2 1090 1097 216 1080 1042 200 ICV_30 $T=272780 138720 0 0 $X=272590 $Y=138480
X1966 1 2 1088 1096 203 1093 1096 216 ICV_30 $T=273240 155040 0 0 $X=273050 $Y=154800
X1967 1 2 1092 1096 201 1091 1096 211 ICV_30 $T=273700 155040 1 0 $X=273510 $Y=152080
X1968 1 2 1101 1096 210 1103 1096 200 ICV_30 $T=275080 149600 1 0 $X=274890 $Y=146640
X1969 1 2 223 224 188 1109 224 166 ICV_30 $T=282440 116960 1 0 $X=282250 $Y=114000
X1970 1 2 1135 1118 189 1145 1118 166 ICV_30 $T=292100 165920 1 0 $X=291910 $Y=162960
X1971 1 2 1158 1160 203 1141 1117 200 ICV_30 $T=303600 144160 0 0 $X=303410 $Y=143920
X1972 1 2 1159 1160 210 1166 1160 201 ICV_30 $T=304060 133280 1 0 $X=303870 $Y=130320
X1973 1 2 1169 1161 166 1188 1161 186 ICV_30 $T=314640 165920 0 0 $X=314450 $Y=165680
X1974 1 2 1184 1163 185 1196 1163 162 ICV_30 $T=319700 149600 0 0 $X=319510 $Y=149360
X1975 1 2 1213 1214 150 1221 1214 185 ICV_30 $T=327980 165920 0 0 $X=327790 $Y=165680
X1976 1 2 1215 233 150 238 233 166 ICV_30 $T=328900 116960 1 0 $X=328710 $Y=114000
X1977 1 2 1217 1218 162 1226 1218 166 ICV_30 $T=330740 160480 1 0 $X=330550 $Y=157520
X1978 1 2 1225 1218 150 1237 1218 189 ICV_30 $T=339020 160480 1 0 $X=338830 $Y=157520
X1979 1 2 1244 241 162 242 241 166 ICV_30 $T=343160 116960 0 0 $X=342970 $Y=116720
X1980 1 2 1256 241 189 246 241 186 ICV_30 $T=351440 116960 0 0 $X=351250 $Y=116720
X1981 1 2 1264 1274 188 1277 1274 166 ICV_30 $T=356960 144160 1 0 $X=356770 $Y=141200
X1982 1 2 1275 1276 186 1270 1276 167 ICV_30 $T=357420 160480 1 0 $X=357230 $Y=157520
X1983 1 2 1279 1272 166 249 241 188 ICV_30 $T=359720 116960 0 0 $X=359530 $Y=116720
X1984 1 2 247 244 185 1285 1284 189 ICV_30 $T=362480 176800 1 0 $X=362290 $Y=173840
X1985 1 2 1296 1261 162 1302 1272 189 ICV_30 $T=370760 127840 0 0 $X=370570 $Y=127600
X1986 1 2 1309 258 166 1310 258 150 ICV_30 $T=380420 160480 0 0 $X=380230 $Y=160240
X1987 1 2 1325 1326 185 1323 1326 166 ICV_30 $T=386400 138720 0 0 $X=386210 $Y=138480
X1988 1 2 1318 1324 189 1322 1326 162 ICV_30 $T=388240 144160 0 0 $X=388050 $Y=143920
X1989 1 2 1306 258 162 1337 1284 162 ICV_30 $T=390080 176800 0 0 $X=389890 $Y=176560
X1990 1 2 1351 274 189 1358 274 162 ICV_30 $T=403420 127840 1 0 $X=403230 $Y=124880
X1991 1 2 1365 1367 189 1366 1367 150 ICV_30 $T=408940 155040 0 0 $X=408750 $Y=154800
X1992 1 2 1369 1372 189 1379 1372 150 ICV_30 $T=416300 127840 0 0 $X=416110 $Y=127600
X1993 1 2 1397 291 294 1394 291 300 ICV_30 $T=426880 176800 0 0 $X=426690 $Y=176560
X1994 1 2 1413 302 309 1419 302 294 ICV_30 $T=437460 171360 0 0 $X=437270 $Y=171120
X1995 1 2 1418 293 167 1415 293 189 ICV_30 $T=441140 116960 1 0 $X=440950 $Y=114000
X1996 1 2 1423 1400 211 1428 1400 201 ICV_30 $T=444360 122400 0 0 $X=444170 $Y=122160
X1997 1 2 1432 1400 200 1425 1410 200 ICV_30 $T=448500 138720 1 0 $X=448310 $Y=135760
X1998 1 2 1450 1449 305 1442 1449 309 ICV_30 $T=457240 165920 0 0 $X=457050 $Y=165680
X1999 1 2 1470 1449 304 1477 1449 320 ICV_30 $T=469200 165920 1 0 $X=469010 $Y=162960
X2000 1 2 1471 1473 342 1478 1473 344 ICV_30 $T=469660 138720 1 0 $X=469470 $Y=135760
X2001 1 2 1492 1490 305 1489 1490 300 ICV_30 $T=479780 165920 1 0 $X=479590 $Y=162960
X2002 1 2 1495 1501 344 1503 361 354 ICV_30 $T=483000 116960 0 0 $X=482810 $Y=116720
X2003 1 2 1504 1473 365 1510 1473 371 ICV_30 $T=487140 127840 1 0 $X=486950 $Y=124880
X2004 1 2 1519 1490 294 1511 1490 309 ICV_30 $T=494500 165920 0 0 $X=494310 $Y=165680
X2005 1 2 1525 1501 356 1528 1501 365 ICV_30 $T=501860 122400 1 0 $X=501670 $Y=119440
X2006 1 2 1546 1534 345 1551 1538 320 ICV_30 $T=508300 149600 1 0 $X=508110 $Y=146640
X2007 1 2 1554 1555 320 1563 1555 300 ICV_30 $T=514740 116960 1 0 $X=514550 $Y=114000
X2008 1 2 1569 386 423 1597 1600 391 ICV_30 $T=533600 165920 1 0 $X=533410 $Y=162960
X2009 1 2 441 443 446 448 443 451 ICV_30 $T=553380 176800 1 0 $X=553190 $Y=173840
X2010 1 2 1636 1638 391 1642 1638 396 ICV_30 $T=562120 165920 1 0 $X=561930 $Y=162960
X2011 1 2 462 463 300 467 463 325 ICV_30 $T=572700 133280 1 0 $X=572510 $Y=130320
X2012 1 2 1651 440 405 483 440 444 ICV_30 $T=592480 160480 1 0 $X=592290 $Y=157520
X2013 1 2 1659 1596 342 1640 440 397 ICV_30 $T=593400 155040 1 0 $X=593210 $Y=152080
X2014 1 2 1686 488 304 1678 488 309 ICV_30 $T=600760 122400 1 0 $X=600570 $Y=119440
X2015 1 2 1701 1679 305 1705 1679 309 ICV_30 $T=609960 144160 1 0 $X=609770 $Y=141200
X2016 1 2 1731 1707 304 1738 1707 309 ICV_30 $T=626520 155040 1 0 $X=626330 $Y=152080
X2017 1 2 1734 1722 409 1746 1722 405 ICV_30 $T=626980 176800 1 0 $X=626790 $Y=173840
X2018 1 2 1777 1756 304 1778 1756 325 ICV_30 $T=651360 133280 0 0 $X=651170 $Y=133040
X2019 1 2 1781 1771 444 527 520 455 ICV_30 $T=651360 176800 1 0 $X=651170 $Y=173840
X2020 1 2 1783 1743 304 1780 1743 309 ICV_30 $T=652280 149600 0 0 $X=652090 $Y=149360
X2021 1 2 1808 523 407 1819 523 409 ICV_30 $T=666540 176800 1 0 $X=666350 $Y=173840
X2022 1 2 1814 1804 423 1825 1804 397 ICV_30 $T=668380 160480 1 0 $X=668190 $Y=157520
X2023 1 2 1863 1841 444 1870 1841 423 ICV_30 $T=692760 165920 0 0 $X=692570 $Y=165680
X2024 1 2 1867 1868 342 1877 1868 344 ICV_30 $T=696440 133280 0 0 $X=696250 $Y=133040
X2025 1 2 1880 537 351 1879 537 365 ICV_30 $T=705180 133280 1 0 $X=704990 $Y=130320
X2026 1 2 1881 1892 344 1898 1868 354 ICV_30 $T=707480 138720 0 0 $X=707290 $Y=138480
X2027 1 2 1882 1891 391 1899 1891 396 ICV_30 $T=707480 165920 0 0 $X=707290 $Y=165680
X2028 1 2 1885 1891 405 1888 1891 409 ICV_30 $T=707480 171360 0 0 $X=707290 $Y=171120
X2029 1 2 1926 1914 344 1931 1914 351 ICV_30 $T=721740 133280 1 0 $X=721550 $Y=130320
X2030 1 2 1924 546 405 1936 1928 407 ICV_30 $T=722200 176800 1 0 $X=722010 $Y=173840
X2031 1 2 1927 1928 397 1935 1928 444 ICV_30 $T=722660 165920 1 0 $X=722470 $Y=162960
X2032 1 2 1925 1920 354 1930 1920 344 ICV_30 $T=723120 122400 0 0 $X=722930 $Y=122160
X2033 1 2 1929 1921 344 1939 1921 351 ICV_30 $T=723580 144160 0 0 $X=723390 $Y=143920
X2034 1 2 1937 1920 351 1942 1914 356 ICV_30 $T=726800 127840 0 0 $X=726610 $Y=127600
X2035 1 2 16 18 2 613 1 sky130_fd_sc_hd__and2_1 $T=17480 116960 1 0 $X=17290 $Y=114000
X2036 1 2 22 18 2 610 1 sky130_fd_sc_hd__and2_1 $T=20240 155040 1 0 $X=20050 $Y=152080
X2037 1 2 24 18 2 616 1 sky130_fd_sc_hd__and2_1 $T=21160 165920 1 0 $X=20970 $Y=162960
X2038 1 2 36 18 2 39 1 sky130_fd_sc_hd__and2_1 $T=31280 116960 0 0 $X=31090 $Y=116720
X2039 1 2 41 18 2 637 1 sky130_fd_sc_hd__and2_1 $T=34040 149600 0 0 $X=33850 $Y=149360
X2040 1 2 42 18 2 642 1 sky130_fd_sc_hd__and2_1 $T=34500 127840 0 0 $X=34310 $Y=127600
X2041 1 2 43 18 2 638 1 sky130_fd_sc_hd__and2_1 $T=34500 176800 0 0 $X=34310 $Y=176560
X2042 1 2 52 25 2 667 1 sky130_fd_sc_hd__and2_1 $T=49680 116960 0 0 $X=49490 $Y=116720
X2043 1 2 53 18 2 671 1 sky130_fd_sc_hd__and2_1 $T=52440 149600 1 0 $X=52250 $Y=146640
X2044 1 2 55 18 2 674 1 sky130_fd_sc_hd__and2_1 $T=58880 116960 1 0 $X=58690 $Y=114000
X2045 1 2 56 18 2 687 1 sky130_fd_sc_hd__and2_1 $T=58880 133280 0 0 $X=58690 $Y=133040
X2046 1 2 57 18 2 59 1 sky130_fd_sc_hd__and2_1 $T=58880 176800 0 0 $X=58690 $Y=176560
X2047 1 2 58 18 2 691 1 sky130_fd_sc_hd__and2_1 $T=60260 171360 1 0 $X=60070 $Y=168400
X2048 1 2 64 18 2 727 1 sky130_fd_sc_hd__and2_1 $T=76360 149600 1 0 $X=76170 $Y=146640
X2049 1 2 68 18 2 69 1 sky130_fd_sc_hd__and2_1 $T=78660 171360 0 0 $X=78470 $Y=171120
X2050 1 2 76 18 2 756 1 sky130_fd_sc_hd__and2_1 $T=97520 138720 0 0 $X=97330 $Y=138480
X2051 1 2 78 18 2 777 1 sky130_fd_sc_hd__and2_1 $T=101660 171360 1 0 $X=101470 $Y=168400
X2052 1 2 79 18 2 785 1 sky130_fd_sc_hd__and2_1 $T=106260 116960 0 0 $X=106070 $Y=116720
X2053 1 2 81 18 2 780 1 sky130_fd_sc_hd__and2_1 $T=109020 176800 0 0 $X=108830 $Y=176560
X2054 1 2 90 18 2 813 1 sky130_fd_sc_hd__and2_1 $T=119600 138720 0 0 $X=119410 $Y=138480
X2055 1 2 91 18 2 812 1 sky130_fd_sc_hd__and2_1 $T=124660 144160 0 0 $X=124470 $Y=143920
X2056 1 2 98 18 2 827 1 sky130_fd_sc_hd__and2_1 $T=129260 160480 1 0 $X=129070 $Y=157520
X2057 1 2 104 18 2 870 1 sky130_fd_sc_hd__and2_1 $T=147200 149600 1 0 $X=147010 $Y=146640
X2058 1 2 105 18 2 866 1 sky130_fd_sc_hd__and2_1 $T=147200 176800 1 0 $X=147010 $Y=173840
X2059 1 2 107 18 2 109 1 sky130_fd_sc_hd__and2_1 $T=152260 116960 0 0 $X=152070 $Y=116720
X2060 1 2 113 18 2 879 1 sky130_fd_sc_hd__and2_1 $T=170660 165920 0 0 $X=170470 $Y=165680
X2061 1 2 118 18 2 918 1 sky130_fd_sc_hd__and2_1 $T=171580 160480 0 0 $X=171390 $Y=160240
X2062 1 2 120 18 2 905 1 sky130_fd_sc_hd__and2_1 $T=174340 138720 0 0 $X=174150 $Y=138480
X2063 1 2 126 18 2 929 1 sky130_fd_sc_hd__and2_1 $T=184460 149600 1 0 $X=184270 $Y=146640
X2064 1 2 129 18 2 957 1 sky130_fd_sc_hd__and2_1 $T=193200 122400 1 0 $X=193010 $Y=119440
X2065 1 2 134 18 2 967 1 sky130_fd_sc_hd__and2_1 $T=198260 127840 0 0 $X=198070 $Y=127600
X2066 1 2 135 18 2 974 1 sky130_fd_sc_hd__and2_1 $T=199640 138720 0 0 $X=199450 $Y=138480
X2067 1 2 136 18 2 966 1 sky130_fd_sc_hd__and2_1 $T=199640 155040 0 0 $X=199450 $Y=154800
X2068 1 2 137 18 2 140 1 sky130_fd_sc_hd__and2_1 $T=199640 176800 0 0 $X=199450 $Y=176560
X2069 1 2 143 18 2 975 1 sky130_fd_sc_hd__and2_1 $T=202860 165920 0 0 $X=202670 $Y=165680
X2070 1 2 42 146 2 991 1 sky130_fd_sc_hd__and2_1 $T=211600 122400 0 0 $X=211410 $Y=122160
X2071 1 2 24 146 2 999 1 sky130_fd_sc_hd__and2_1 $T=212980 165920 1 0 $X=212790 $Y=162960
X2072 1 2 41 146 2 992 1 sky130_fd_sc_hd__and2_1 $T=213900 144160 0 0 $X=213710 $Y=143920
X2073 1 2 16 146 2 184 1 sky130_fd_sc_hd__and2_1 $T=235060 116960 0 0 $X=234870 $Y=116720
X2074 1 2 190 191 2 1048 1 sky130_fd_sc_hd__and2_1 $T=244720 144160 1 0 $X=244530 $Y=141200
X2075 1 2 209 191 2 1067 1 sky130_fd_sc_hd__and2_1 $T=255760 116960 0 0 $X=255570 $Y=116720
X2076 1 2 72 191 2 1069 1 sky130_fd_sc_hd__and2_1 $T=255760 160480 0 0 $X=255570 $Y=160240
X2077 1 2 58 146 2 1083 1 sky130_fd_sc_hd__and2_1 $T=266340 165920 0 0 $X=266150 $Y=165680
X2078 1 2 52 191 2 1095 1 sky130_fd_sc_hd__and2_1 $T=270480 138720 0 0 $X=270290 $Y=138480
X2079 1 2 33 146 2 1111 1 sky130_fd_sc_hd__and2_1 $T=282440 155040 0 0 $X=282250 $Y=154800
X2080 1 2 124 191 2 1131 1 sky130_fd_sc_hd__and2_1 $T=289800 127840 1 0 $X=289610 $Y=124880
X2081 1 2 228 191 2 1143 1 sky130_fd_sc_hd__and2_1 $T=297620 144160 1 0 $X=297430 $Y=141200
X2082 1 2 53 146 2 1152 1 sky130_fd_sc_hd__and2_1 $T=298080 149600 1 0 $X=297890 $Y=146640
X2083 1 2 81 146 2 1157 1 sky130_fd_sc_hd__and2_1 $T=301300 160480 0 0 $X=301110 $Y=160240
X2084 1 2 64 146 2 1183 1 sky130_fd_sc_hd__and2_1 $T=315100 144160 0 0 $X=314910 $Y=143920
X2085 1 2 56 146 2 1185 1 sky130_fd_sc_hd__and2_1 $T=318780 122400 0 0 $X=318590 $Y=122160
X2086 1 2 68 146 2 1202 1 sky130_fd_sc_hd__and2_1 $T=322920 171360 0 0 $X=322730 $Y=171120
X2087 1 2 234 146 2 236 1 sky130_fd_sc_hd__and2_1 $T=324760 176800 1 0 $X=324570 $Y=173840
X2088 1 2 237 191 2 1189 1 sky130_fd_sc_hd__and2_1 $T=328900 127840 1 0 $X=328710 $Y=124880
X2089 1 2 91 146 2 1239 1 sky130_fd_sc_hd__and2_1 $T=342700 133280 0 0 $X=342510 $Y=133040
X2090 1 2 113 146 2 1250 1 sky130_fd_sc_hd__and2_1 $T=345920 144160 1 0 $X=345730 $Y=141200
X2091 1 2 121 146 2 1254 1 sky130_fd_sc_hd__and2_1 $T=354200 122400 1 0 $X=354010 $Y=119440
X2092 1 2 98 146 2 1255 1 sky130_fd_sc_hd__and2_1 $T=356040 165920 0 0 $X=355850 $Y=165680
X2093 1 2 78 146 2 1249 1 sky130_fd_sc_hd__and2_1 $T=358340 160480 0 0 $X=358150 $Y=160240
X2094 1 2 122 146 2 1281 1 sky130_fd_sc_hd__and2_1 $T=363860 171360 0 0 $X=363670 $Y=171120
X2095 1 2 129 146 2 251 1 sky130_fd_sc_hd__and2_1 $T=364320 116960 1 0 $X=364130 $Y=114000
X2096 1 2 253 146 2 254 1 sky130_fd_sc_hd__and2_1 $T=366620 176800 0 0 $X=366430 $Y=176560
X2097 1 2 105 146 2 1297 1 sky130_fd_sc_hd__and2_1 $T=370760 155040 0 0 $X=370570 $Y=154800
X2098 1 2 137 146 2 1305 1 sky130_fd_sc_hd__and2_1 $T=374900 133280 0 0 $X=374710 $Y=133040
X2099 1 2 118 146 2 1330 1 sky130_fd_sc_hd__and2_1 $T=388700 160480 0 0 $X=388510 $Y=160240
X2100 1 2 266 146 2 1345 1 sky130_fd_sc_hd__and2_1 $T=396060 160480 0 0 $X=395870 $Y=160240
X2101 1 2 75 146 2 1348 1 sky130_fd_sc_hd__and2_1 $T=398820 149600 0 0 $X=398630 $Y=149360
X2102 1 2 272 146 2 1353 1 sky130_fd_sc_hd__and2_1 $T=402960 138720 1 0 $X=402770 $Y=135760
X2103 1 2 266 191 2 1387 1 sky130_fd_sc_hd__and2_1 $T=423660 133280 1 0 $X=423470 $Y=130320
X2104 1 2 122 191 2 1392 1 sky130_fd_sc_hd__and2_1 $T=423660 138720 0 0 $X=423470 $Y=138480
X2105 1 2 289 290 2 1391 1 sky130_fd_sc_hd__and2_1 $T=426880 171360 1 0 $X=426690 $Y=168400
X2106 1 2 306 290 2 1403 1 sky130_fd_sc_hd__and2_1 $T=438380 176800 1 0 $X=438190 $Y=173840
X2107 1 2 308 290 2 1420 1 sky130_fd_sc_hd__and2_1 $T=441140 155040 1 0 $X=440950 $Y=152080
X2108 1 2 312 290 2 1422 1 sky130_fd_sc_hd__and2_1 $T=443440 176800 0 0 $X=443250 $Y=176560
X2109 1 2 322 290 2 1437 1 sky130_fd_sc_hd__and2_1 $T=455400 122400 1 0 $X=455210 $Y=119440
X2110 1 2 330 332 2 1458 1 sky130_fd_sc_hd__and2_1 $T=465060 149600 1 0 $X=464870 $Y=146640
X2111 1 2 333 332 2 1461 1 sky130_fd_sc_hd__and2_1 $T=466440 138720 0 0 $X=466250 $Y=138480
X2112 1 2 336 332 2 1472 1 sky130_fd_sc_hd__and2_1 $T=468740 127840 0 0 $X=468550 $Y=127600
X2113 1 2 337 290 2 1462 1 sky130_fd_sc_hd__and2_1 $T=469200 171360 1 0 $X=469010 $Y=168400
X2114 1 2 352 290 2 1500 1 sky130_fd_sc_hd__and2_1 $T=480240 165920 0 0 $X=480050 $Y=165680
X2115 1 2 352 332 2 1521 1 sky130_fd_sc_hd__and2_1 $T=494500 149600 1 0 $X=494310 $Y=146640
X2116 1 2 384 290 2 1535 1 sky130_fd_sc_hd__and2_1 $T=504620 155040 1 0 $X=504430 $Y=152080
X2117 1 2 306 370 2 1537 1 sky130_fd_sc_hd__and2_1 $T=506460 176800 1 0 $X=506270 $Y=173840
X2118 1 2 336 290 2 1532 1 sky130_fd_sc_hd__and2_1 $T=507840 127840 0 0 $X=507650 $Y=127600
X2119 1 2 350 370 2 1577 1 sky130_fd_sc_hd__and2_1 $T=529000 160480 0 0 $X=528810 $Y=160240
X2120 1 2 308 332 2 1582 1 sky130_fd_sc_hd__and2_1 $T=536360 127840 0 0 $X=536170 $Y=127600
X2121 1 2 421 370 2 1598 1 sky130_fd_sc_hd__and2_1 $T=536360 176800 0 0 $X=536170 $Y=176560
X2122 1 2 312 332 2 1587 1 sky130_fd_sc_hd__and2_1 $T=536820 122400 1 0 $X=536630 $Y=119440
X2123 1 2 410 332 2 1594 1 sky130_fd_sc_hd__and2_1 $T=539120 149600 1 0 $X=538930 $Y=146640
X2124 1 2 434 370 2 1627 1 sky130_fd_sc_hd__and2_1 $T=557520 160480 1 0 $X=557330 $Y=157520
X2125 1 2 468 469 2 471 1 sky130_fd_sc_hd__and2_1 $T=578680 176800 1 0 $X=578490 $Y=173840
X2126 1 2 472 290 2 1664 1 sky130_fd_sc_hd__and2_1 $T=581440 138720 1 0 $X=581250 $Y=135760
X2127 1 2 447 370 2 1667 1 sky130_fd_sc_hd__and2_1 $T=596620 165920 1 0 $X=596430 $Y=162960
X2128 1 2 489 290 2 1687 1 sky130_fd_sc_hd__and2_1 $T=605820 155040 1 0 $X=605630 $Y=152080
X2129 1 2 495 290 2 1700 1 sky130_fd_sc_hd__and2_1 $T=606280 116960 1 0 $X=606090 $Y=114000
X2130 1 2 499 370 2 1706 1 sky130_fd_sc_hd__and2_1 $T=610880 165920 0 0 $X=610690 $Y=165680
X2131 1 2 501 469 2 1698 1 sky130_fd_sc_hd__and2_1 $T=613640 176800 1 0 $X=613450 $Y=173840
X2132 1 2 504 290 2 1724 1 sky130_fd_sc_hd__and2_1 $T=619160 133280 1 0 $X=618970 $Y=130320
X2133 1 2 508 290 2 1718 1 sky130_fd_sc_hd__and2_1 $T=620540 155040 0 0 $X=620350 $Y=154800
X2134 1 2 510 469 2 1729 1 sky130_fd_sc_hd__and2_1 $T=623300 171360 0 0 $X=623110 $Y=171120
X2135 1 2 509 290 2 1735 1 sky130_fd_sc_hd__and2_1 $T=627440 144160 0 0 $X=627250 $Y=143920
X2136 1 2 404 332 2 1774 1 sky130_fd_sc_hd__and2_1 $T=649520 144160 1 0 $X=649330 $Y=141200
X2137 1 2 490 332 2 1799 1 sky130_fd_sc_hd__and2_1 $T=662860 127840 0 0 $X=662670 $Y=127600
X2138 1 2 461 332 2 1809 1 sky130_fd_sc_hd__and2_1 $T=665620 155040 1 0 $X=665430 $Y=152080
X2139 1 2 472 332 2 1834 1 sky130_fd_sc_hd__and2_1 $T=677120 133280 1 0 $X=676930 $Y=130320
X2140 1 2 479 370 2 1833 1 sky130_fd_sc_hd__and2_1 $T=677120 165920 1 0 $X=676930 $Y=162960
X2141 1 2 495 332 2 1838 1 sky130_fd_sc_hd__and2_1 $T=683560 122400 0 0 $X=683370 $Y=122160
X2142 1 2 509 332 2 1845 1 sky130_fd_sc_hd__and2_1 $T=684020 144160 0 0 $X=683830 $Y=143920
X2143 1 2 510 370 2 1873 1 sky130_fd_sc_hd__and2_1 $T=696440 160480 1 0 $X=696250 $Y=157520
X2144 1 2 468 370 2 1889 1 sky130_fd_sc_hd__and2_1 $T=704720 176800 0 0 $X=704530 $Y=176560
X2145 1 2 511 332 2 1902 1 sky130_fd_sc_hd__and2_1 $T=711620 122400 1 0 $X=711430 $Y=119440
X2146 1 2 504 332 2 1909 1 sky130_fd_sc_hd__and2_1 $T=714840 127840 0 0 $X=714650 $Y=127600
X2147 1 2 489 332 2 1912 1 sky130_fd_sc_hd__and2_1 $T=714840 144160 0 0 $X=714650 $Y=143920
X2148 1 2 502 370 2 1913 1 sky130_fd_sc_hd__and2_1 $T=718980 171360 1 0 $X=718790 $Y=168400
X2149 1 2 111 610 2 585 1 sky130_fd_sc_hd__dlclkp_1 $T=15640 149600 0 0 $X=15450 $Y=149360
X2150 1 2 111 23 2 30 1 sky130_fd_sc_hd__dlclkp_1 $T=18860 176800 0 0 $X=18670 $Y=176560
X2151 1 2 111 613 2 583 1 sky130_fd_sc_hd__dlclkp_1 $T=20240 116960 1 0 $X=20050 $Y=114000
X2152 1 2 111 616 2 587 1 sky130_fd_sc_hd__dlclkp_1 $T=20240 165920 0 0 $X=20050 $Y=165680
X2153 1 2 111 637 2 639 1 sky130_fd_sc_hd__dlclkp_1 $T=32200 155040 1 0 $X=32010 $Y=152080
X2154 1 2 111 638 2 46 1 sky130_fd_sc_hd__dlclkp_1 $T=32660 176800 1 0 $X=32470 $Y=173840
X2155 1 2 111 642 2 641 1 sky130_fd_sc_hd__dlclkp_1 $T=40020 133280 0 0 $X=39830 $Y=133040
X2156 1 2 111 667 2 54 1 sky130_fd_sc_hd__dlclkp_1 $T=48300 116960 1 0 $X=48110 $Y=114000
X2157 1 2 111 671 2 666 1 sky130_fd_sc_hd__dlclkp_1 $T=51060 155040 1 0 $X=50870 $Y=152080
X2158 1 2 111 674 2 675 1 sky130_fd_sc_hd__dlclkp_1 $T=52440 116960 0 0 $X=52250 $Y=116720
X2159 1 2 111 687 2 685 1 sky130_fd_sc_hd__dlclkp_1 $T=57040 138720 1 0 $X=56850 $Y=135760
X2160 1 2 111 691 2 664 1 sky130_fd_sc_hd__dlclkp_1 $T=62100 165920 0 0 $X=61910 $Y=165680
X2161 1 2 111 61 2 63 1 sky130_fd_sc_hd__dlclkp_1 $T=69460 116960 1 0 $X=69270 $Y=114000
X2162 1 2 111 727 2 701 1 sky130_fd_sc_hd__dlclkp_1 $T=76360 155040 1 0 $X=76170 $Y=152080
X2163 1 2 111 756 2 726 1 sky130_fd_sc_hd__dlclkp_1 $T=91540 138720 1 0 $X=91350 $Y=135760
X2164 1 2 111 780 2 80 1 sky130_fd_sc_hd__dlclkp_1 $T=102580 176800 0 0 $X=102390 $Y=176560
X2165 1 2 111 777 2 729 1 sky130_fd_sc_hd__dlclkp_1 $T=104420 165920 0 0 $X=104230 $Y=165680
X2166 1 2 111 785 2 788 1 sky130_fd_sc_hd__dlclkp_1 $T=104880 116960 1 0 $X=104690 $Y=114000
X2167 1 2 111 812 2 782 1 sky130_fd_sc_hd__dlclkp_1 $T=118220 144160 0 0 $X=118030 $Y=143920
X2168 1 2 111 813 2 761 1 sky130_fd_sc_hd__dlclkp_1 $T=120060 138720 1 0 $X=119870 $Y=135760
X2169 1 2 111 827 2 791 1 sky130_fd_sc_hd__dlclkp_1 $T=126040 165920 0 0 $X=125850 $Y=165680
X2170 1 2 111 97 2 89 1 sky130_fd_sc_hd__dlclkp_1 $T=127420 176800 0 0 $X=127230 $Y=176560
X2171 1 2 111 866 2 106 1 sky130_fd_sc_hd__dlclkp_1 $T=144900 171360 1 0 $X=144710 $Y=168400
X2172 1 2 111 870 2 829 1 sky130_fd_sc_hd__dlclkp_1 $T=147200 149600 0 0 $X=147010 $Y=149360
X2173 1 2 111 879 2 843 1 sky130_fd_sc_hd__dlclkp_1 $T=152260 165920 0 0 $X=152070 $Y=165680
X2174 1 2 111 905 2 884 1 sky130_fd_sc_hd__dlclkp_1 $T=163300 138720 1 0 $X=163110 $Y=135760
X2175 1 2 111 114 2 906 1 sky130_fd_sc_hd__dlclkp_1 $T=166060 116960 0 0 $X=165870 $Y=116720
X2176 1 2 111 115 2 119 1 sky130_fd_sc_hd__dlclkp_1 $T=167440 176800 0 0 $X=167250 $Y=176560
X2177 1 2 111 918 2 898 1 sky130_fd_sc_hd__dlclkp_1 $T=174340 160480 0 0 $X=174150 $Y=160240
X2178 1 2 111 929 2 876 1 sky130_fd_sc_hd__dlclkp_1 $T=175720 155040 1 0 $X=175530 $Y=152080
X2179 1 2 111 957 2 932 1 sky130_fd_sc_hd__dlclkp_1 $T=189980 116960 0 0 $X=189790 $Y=116720
X2180 1 2 111 966 2 933 1 sky130_fd_sc_hd__dlclkp_1 $T=193660 160480 1 0 $X=193470 $Y=157520
X2181 1 2 111 967 2 928 1 sky130_fd_sc_hd__dlclkp_1 $T=194120 133280 0 0 $X=193930 $Y=133040
X2182 1 2 111 975 2 125 1 sky130_fd_sc_hd__dlclkp_1 $T=200560 171360 1 0 $X=200370 $Y=168400
X2183 1 2 111 974 2 941 1 sky130_fd_sc_hd__dlclkp_1 $T=202860 144160 1 0 $X=202670 $Y=141200
X2184 1 2 111 991 2 998 1 sky130_fd_sc_hd__dlclkp_1 $T=208380 127840 0 0 $X=208190 $Y=127600
X2185 1 2 111 992 2 1002 1 sky130_fd_sc_hd__dlclkp_1 $T=209760 144160 1 0 $X=209570 $Y=141200
X2186 1 2 111 999 2 1001 1 sky130_fd_sc_hd__dlclkp_1 $T=216660 165920 1 0 $X=216470 $Y=162960
X2187 1 2 111 192 2 199 1 sky130_fd_sc_hd__dlclkp_1 $T=241500 176800 0 0 $X=241310 $Y=176560
X2188 1 2 111 1048 2 1044 1 sky130_fd_sc_hd__dlclkp_1 $T=244720 138720 1 0 $X=244530 $Y=135760
X2189 1 2 111 1067 2 1075 1 sky130_fd_sc_hd__dlclkp_1 $T=258060 122400 1 0 $X=257870 $Y=119440
X2190 1 2 111 1069 2 1076 1 sky130_fd_sc_hd__dlclkp_1 $T=258520 160480 1 0 $X=258330 $Y=157520
X2191 1 2 111 1083 2 1084 1 sky130_fd_sc_hd__dlclkp_1 $T=265880 171360 1 0 $X=265690 $Y=168400
X2192 1 2 111 1095 2 1108 1 sky130_fd_sc_hd__dlclkp_1 $T=273700 144160 1 0 $X=273510 $Y=141200
X2193 1 2 111 1111 2 1124 1 sky130_fd_sc_hd__dlclkp_1 $T=279680 160480 0 0 $X=279490 $Y=160240
X2194 1 2 111 1131 2 1133 1 sky130_fd_sc_hd__dlclkp_1 $T=292560 127840 0 0 $X=292370 $Y=127600
X2195 1 2 111 1143 2 1148 1 sky130_fd_sc_hd__dlclkp_1 $T=292560 138720 0 0 $X=292370 $Y=138480
X2196 1 2 111 1152 2 1153 1 sky130_fd_sc_hd__dlclkp_1 $T=301760 149600 0 0 $X=301570 $Y=149360
X2197 1 2 111 1157 2 1156 1 sky130_fd_sc_hd__dlclkp_1 $T=305440 165920 0 0 $X=305250 $Y=165680
X2198 1 2 111 1185 2 1192 1 sky130_fd_sc_hd__dlclkp_1 $T=316020 133280 0 0 $X=315830 $Y=133040
X2199 1 2 111 1189 2 1187 1 sky130_fd_sc_hd__dlclkp_1 $T=317860 133280 1 0 $X=317670 $Y=130320
X2200 1 2 111 1183 2 1208 1 sky130_fd_sc_hd__dlclkp_1 $T=320160 149600 1 0 $X=319970 $Y=146640
X2201 1 2 111 1202 2 1206 1 sky130_fd_sc_hd__dlclkp_1 $T=322000 171360 1 0 $X=321810 $Y=168400
X2202 1 2 111 1239 2 1248 1 sky130_fd_sc_hd__dlclkp_1 $T=340860 133280 1 0 $X=340670 $Y=130320
X2203 1 2 111 1249 2 1253 1 sky130_fd_sc_hd__dlclkp_1 $T=344540 160480 0 0 $X=344350 $Y=160240
X2204 1 2 111 1250 2 1252 1 sky130_fd_sc_hd__dlclkp_1 $T=345920 144160 0 0 $X=345730 $Y=143920
X2205 1 2 111 1254 2 1257 1 sky130_fd_sc_hd__dlclkp_1 $T=347760 122400 1 0 $X=347570 $Y=119440
X2206 1 2 111 1255 2 243 1 sky130_fd_sc_hd__dlclkp_1 $T=348220 160480 1 0 $X=348030 $Y=157520
X2207 1 2 111 1281 2 255 1 sky130_fd_sc_hd__dlclkp_1 $T=366160 171360 1 0 $X=365970 $Y=168400
X2208 1 2 111 1297 2 1301 1 sky130_fd_sc_hd__dlclkp_1 $T=369380 155040 1 0 $X=369190 $Y=152080
X2209 1 2 111 1305 2 1312 1 sky130_fd_sc_hd__dlclkp_1 $T=376280 133280 1 0 $X=376090 $Y=130320
X2210 1 2 111 1330 2 1327 1 sky130_fd_sc_hd__dlclkp_1 $T=385480 165920 1 0 $X=385290 $Y=162960
X2211 1 2 111 1348 2 1349 1 sky130_fd_sc_hd__dlclkp_1 $T=396980 149600 1 0 $X=396790 $Y=146640
X2212 1 2 111 271 2 269 1 sky130_fd_sc_hd__dlclkp_1 $T=398820 116960 1 0 $X=398630 $Y=114000
X2213 1 2 111 1345 2 1350 1 sky130_fd_sc_hd__dlclkp_1 $T=398820 155040 0 0 $X=398630 $Y=154800
X2214 1 2 111 1353 2 1354 1 sky130_fd_sc_hd__dlclkp_1 $T=402500 133280 0 0 $X=402310 $Y=133040
X2215 1 2 111 1387 2 1395 1 sky130_fd_sc_hd__dlclkp_1 $T=420440 127840 1 0 $X=420250 $Y=124880
X2216 1 2 481 1391 2 1396 1 sky130_fd_sc_hd__dlclkp_1 $T=421820 165920 1 0 $X=421630 $Y=162960
X2217 1 2 111 1392 2 1398 1 sky130_fd_sc_hd__dlclkp_1 $T=423660 144160 1 0 $X=423470 $Y=141200
X2218 1 2 481 1403 2 279 1 sky130_fd_sc_hd__dlclkp_1 $T=431940 176800 1 0 $X=431750 $Y=173840
X2219 1 2 481 1420 2 1426 1 sky130_fd_sc_hd__dlclkp_1 $T=441140 160480 1 0 $X=440950 $Y=157520
X2220 1 2 481 1422 2 314 1 sky130_fd_sc_hd__dlclkp_1 $T=441600 176800 1 0 $X=441410 $Y=173840
X2221 1 2 481 1437 2 1440 1 sky130_fd_sc_hd__dlclkp_1 $T=450340 127840 1 0 $X=450150 $Y=124880
X2222 1 2 481 1458 2 1466 1 sky130_fd_sc_hd__dlclkp_1 $T=461840 144160 1 0 $X=461650 $Y=141200
X2223 1 2 481 1461 2 1467 1 sky130_fd_sc_hd__dlclkp_1 $T=462300 138720 1 0 $X=462110 $Y=135760
X2224 1 2 481 1462 2 335 1 sky130_fd_sc_hd__dlclkp_1 $T=462300 176800 1 0 $X=462110 $Y=173840
X2225 1 2 481 1472 2 1476 1 sky130_fd_sc_hd__dlclkp_1 $T=469200 127840 1 0 $X=469010 $Y=124880
X2226 1 2 481 1500 2 1475 1 sky130_fd_sc_hd__dlclkp_1 $T=481160 171360 1 0 $X=480970 $Y=168400
X2227 1 2 481 1521 2 1523 1 sky130_fd_sc_hd__dlclkp_1 $T=494040 144160 0 0 $X=493850 $Y=143920
X2228 1 2 481 1532 2 1548 1 sky130_fd_sc_hd__dlclkp_1 $T=504160 122400 0 0 $X=503970 $Y=122160
X2229 1 2 481 1535 2 1547 1 sky130_fd_sc_hd__dlclkp_1 $T=504160 149600 0 0 $X=503970 $Y=149360
X2230 1 2 481 1537 2 392 1 sky130_fd_sc_hd__dlclkp_1 $T=504160 176800 0 0 $X=503970 $Y=176560
X2231 1 2 481 1577 2 1580 1 sky130_fd_sc_hd__dlclkp_1 $T=527160 165920 1 0 $X=526970 $Y=162960
X2232 1 2 481 1582 2 1588 1 sky130_fd_sc_hd__dlclkp_1 $T=529920 127840 0 0 $X=529730 $Y=127600
X2233 1 2 481 1587 2 424 1 sky130_fd_sc_hd__dlclkp_1 $T=532220 116960 0 0 $X=532030 $Y=116720
X2234 1 2 481 1594 2 1606 1 sky130_fd_sc_hd__dlclkp_1 $T=535900 155040 1 0 $X=535710 $Y=152080
X2235 1 2 481 1598 2 428 1 sky130_fd_sc_hd__dlclkp_1 $T=537740 176800 1 0 $X=537550 $Y=173840
X2236 1 2 481 1627 2 1625 1 sky130_fd_sc_hd__dlclkp_1 $T=554760 165920 1 0 $X=554570 $Y=162960
X2237 1 2 481 1664 2 1665 1 sky130_fd_sc_hd__dlclkp_1 $T=583740 133280 0 0 $X=583550 $Y=133040
X2238 1 2 481 1667 2 1668 1 sky130_fd_sc_hd__dlclkp_1 $T=587420 160480 0 0 $X=587230 $Y=160240
X2239 1 2 481 1687 2 1666 1 sky130_fd_sc_hd__dlclkp_1 $T=599380 149600 0 0 $X=599190 $Y=149360
X2240 1 2 481 1698 2 500 1 sky130_fd_sc_hd__dlclkp_1 $T=604440 176800 0 0 $X=604250 $Y=176560
X2241 1 2 481 1700 2 477 1 sky130_fd_sc_hd__dlclkp_1 $T=605820 116960 0 0 $X=605630 $Y=116720
X2242 1 2 481 1706 2 1710 1 sky130_fd_sc_hd__dlclkp_1 $T=608580 171360 0 0 $X=608390 $Y=171120
X2243 1 2 481 1718 2 1688 1 sky130_fd_sc_hd__dlclkp_1 $T=616400 160480 0 0 $X=616210 $Y=160240
X2244 1 2 481 1729 2 512 1 sky130_fd_sc_hd__dlclkp_1 $T=620540 176800 1 0 $X=620350 $Y=173840
X2245 1 2 481 1724 2 1733 1 sky130_fd_sc_hd__dlclkp_1 $T=621460 138720 1 0 $X=621270 $Y=135760
X2246 1 2 481 1735 2 1748 1 sky130_fd_sc_hd__dlclkp_1 $T=626980 149600 1 0 $X=626790 $Y=146640
X2247 1 2 481 515 2 519 1 sky130_fd_sc_hd__dlclkp_1 $T=628360 116960 1 0 $X=628170 $Y=114000
X2248 1 2 481 1774 2 1779 1 sky130_fd_sc_hd__dlclkp_1 $T=644460 144160 0 0 $X=644270 $Y=143920
X2249 1 2 481 1799 2 529 1 sky130_fd_sc_hd__dlclkp_1 $T=658720 127840 1 0 $X=658530 $Y=124880
X2250 1 2 481 1809 2 1818 1 sky130_fd_sc_hd__dlclkp_1 $T=665160 149600 0 0 $X=664970 $Y=149360
X2251 1 2 481 1833 2 1835 1 sky130_fd_sc_hd__dlclkp_1 $T=676660 160480 1 0 $X=676470 $Y=157520
X2252 1 2 481 1838 2 538 1 sky130_fd_sc_hd__dlclkp_1 $T=679420 116960 0 0 $X=679230 $Y=116720
X2253 1 2 481 1845 2 1859 1 sky130_fd_sc_hd__dlclkp_1 $T=684480 144160 1 0 $X=684290 $Y=141200
X2254 1 2 481 1834 2 1844 1 sky130_fd_sc_hd__dlclkp_1 $T=686780 133280 1 0 $X=686590 $Y=130320
X2255 1 2 481 1873 2 1871 1 sky130_fd_sc_hd__dlclkp_1 $T=699200 160480 0 0 $X=699010 $Y=160240
X2256 1 2 481 1889 2 544 1 sky130_fd_sc_hd__dlclkp_1 $T=708400 176800 0 0 $X=708210 $Y=176560
X2257 1 2 481 1902 2 545 1 sky130_fd_sc_hd__dlclkp_1 $T=713460 116960 1 0 $X=713270 $Y=114000
X2258 1 2 481 1909 2 1904 1 sky130_fd_sc_hd__dlclkp_1 $T=713460 133280 1 0 $X=713270 $Y=130320
X2259 1 2 481 1913 2 1919 1 sky130_fd_sc_hd__dlclkp_1 $T=714840 165920 1 0 $X=714650 $Y=162960
X2260 1 2 481 1912 2 1918 1 sky130_fd_sc_hd__dlclkp_1 $T=715300 149600 0 0 $X=715110 $Y=149360
X2261 1 2 584 5 591 ICV_35 $T=6900 149600 1 0 $X=6710 $Y=146640
X2262 1 2 585 26 618 ICV_35 $T=20700 160480 0 0 $X=20510 $Y=160240
X2263 1 2 587 27 636 ICV_35 $T=24380 176800 1 0 $X=24190 $Y=173840
X2264 1 2 641 9 656 ICV_35 $T=36340 149600 1 0 $X=36150 $Y=146640
X2265 1 2 639 5 658 ICV_35 $T=36340 171360 1 0 $X=36150 $Y=168400
X2266 1 2 44 8 668 ICV_35 $T=44160 127840 0 0 $X=43970 $Y=127600
X2267 1 2 664 9 709 ICV_35 $T=62100 171360 0 0 $X=61910 $Y=171120
X2268 1 2 701 9 721 ICV_35 $T=68080 160480 0 0 $X=67890 $Y=160240
X2269 1 2 62 29 65 ICV_35 $T=70380 171360 0 0 $X=70190 $Y=171120
X2270 1 2 729 9 749 ICV_35 $T=80960 171360 0 0 $X=80770 $Y=171120
X2271 1 2 791 6 809 ICV_35 $T=109480 171360 0 0 $X=109290 $Y=171120
X2272 1 2 791 9 835 ICV_35 $T=123740 165920 1 0 $X=123550 $Y=162960
X2273 1 2 100 8 860 ICV_35 $T=136620 133280 1 0 $X=136430 $Y=130320
X2274 1 2 843 27 885 ICV_35 $T=151340 171360 1 0 $X=151150 $Y=168400
X2275 1 2 898 9 914 ICV_35 $T=162840 160480 0 0 $X=162650 $Y=160240
X2276 1 2 928 6 940 ICV_35 $T=176640 138720 0 0 $X=176450 $Y=138480
X2277 1 2 932 29 948 ICV_35 $T=181700 116960 0 0 $X=181510 $Y=116720
X2278 1 2 933 5 978 ICV_35 $T=197340 165920 1 0 $X=197150 $Y=162960
X2279 1 2 998 153 1005 ICV_35 $T=213900 122400 0 0 $X=213710 $Y=122160
X2280 1 2 160 161 172 ICV_35 $T=219420 171360 0 0 $X=219230 $Y=171120
X2281 1 2 1041 193 1051 ICV_35 $T=241960 133280 0 0 $X=241770 $Y=133040
X2282 1 2 183 155 1066 ICV_35 $T=248860 122400 1 0 $X=248670 $Y=119440
X2283 1 2 1076 213 1091 ICV_35 $T=264040 149600 1 0 $X=263850 $Y=146640
X2284 1 2 1077 205 1098 ICV_35 $T=265880 133280 0 0 $X=265690 $Y=133040
X2285 1 2 1084 156 1121 ICV_35 $T=277380 165920 0 0 $X=277190 $Y=165680
X2286 1 2 1124 155 1116 ICV_35 $T=290720 176800 0 0 $X=290530 $Y=176560
X2287 1 2 1156 179 1170 ICV_35 $T=300840 171360 1 0 $X=300650 $Y=168400
X2288 1 2 1148 206 1182 ICV_35 $T=308200 144160 1 0 $X=308010 $Y=141200
X2289 1 2 1187 196 1232 ICV_35 $T=333960 122400 0 0 $X=333770 $Y=122160
X2290 1 2 1187 197 1233 ICV_35 $T=333960 127840 0 0 $X=333770 $Y=127600
X2291 1 2 240 156 1244 ICV_35 $T=337180 116960 1 0 $X=336990 $Y=114000
X2292 1 2 1252 179 1264 ICV_35 $T=348220 144160 1 0 $X=348030 $Y=141200
X2293 1 2 1252 178 1295 ICV_35 $T=361100 149600 0 0 $X=360910 $Y=149360
X2294 1 2 1301 153 1315 ICV_35 $T=373060 155040 0 0 $X=372870 $Y=154800
X2295 1 2 1312 179 1328 ICV_35 $T=379040 127840 0 0 $X=378850 $Y=127600
X2296 1 2 269 178 1351 ICV_35 $T=398820 116960 0 0 $X=398630 $Y=116720
X2297 1 2 1350 175 1384 ICV_35 $T=413080 165920 1 0 $X=412890 $Y=162960
X2298 1 2 1398 206 1404 ICV_35 $T=426880 144160 0 0 $X=426690 $Y=143920
X2299 1 2 1396 295 301 ICV_35 $T=426880 171360 0 0 $X=426690 $Y=171120
X2300 1 2 279 303 311 ICV_35 $T=435160 176800 0 0 $X=434970 $Y=176560
X2301 1 2 313 281 1439 ICV_35 $T=446200 116960 0 0 $X=446010 $Y=116720
X2302 1 2 1466 357 1497 ICV_35 $T=483000 144160 0 0 $X=482810 $Y=143920
X2303 1 2 160 351 1585 ICV_35 $T=525320 155040 1 0 $X=525130 $Y=152080
X2304 1 2 160 365 1590 ICV_35 $T=530380 155040 0 0 $X=530190 $Y=154800
X2305 1 2 428 380 436 ICV_35 $T=543260 176800 0 0 $X=543070 $Y=176560
X2306 1 2 1668 399 1683 ICV_35 $T=588340 171360 1 0 $X=588150 $Y=168400
X2307 1 2 1688 295 1702 ICV_35 $T=600760 160480 1 0 $X=600570 $Y=157520
X2308 1 2 1704 310 1720 ICV_35 $T=610880 133280 1 0 $X=610690 $Y=130320
X2309 1 2 1733 303 1752 ICV_35 $T=627900 138720 1 0 $X=627710 $Y=135760
X2310 1 2 1795 388 1812 ICV_35 $T=660560 160480 0 0 $X=660370 $Y=160240
X2311 1 2 1835 395 1860 ICV_35 $T=683560 160480 0 0 $X=683370 $Y=160240
X2312 1 2 1835 380 1865 ICV_35 $T=686780 171360 0 0 $X=686590 $Y=171120
X2313 1 2 1871 399 1885 ICV_35 $T=697820 171360 1 0 $X=697630 $Y=168400
X2314 1 2 1869 340 1887 ICV_35 $T=698740 149600 0 0 $X=698550 $Y=149360
X2315 1 2 1919 395 1927 ICV_35 $T=718980 160480 0 0 $X=718790 $Y=160240
X2316 1 2 729 29 766 ICV_36 $T=90160 171360 0 0 $X=89970 $Y=171120
X2317 1 2 788 27 802 ICV_36 $T=105800 133280 0 0 $X=105610 $Y=133040
X2318 1 2 89 9 821 ICV_36 $T=115920 176800 1 0 $X=115730 $Y=173840
X2319 1 2 816 5 836 ICV_36 $T=122360 116960 0 0 $X=122170 $Y=116720
X2320 1 2 843 28 863 ICV_36 $T=135240 171360 0 0 $X=135050 $Y=171120
X2321 1 2 1076 204 1103 ICV_36 $T=265880 144160 0 0 $X=265690 $Y=143920
X2322 1 2 1084 179 1120 ICV_36 $T=275080 171360 0 0 $X=274890 $Y=171120
X2323 1 2 1133 194 1175 ICV_36 $T=300840 122400 0 0 $X=300650 $Y=122160
X2324 1 2 243 176 252 ICV_36 $T=356500 176800 0 0 $X=356310 $Y=176560
X2325 1 2 269 155 1376 ICV_36 $T=408480 122400 0 0 $X=408290 $Y=122160
X2326 1 2 313 310 1444 ICV_36 $T=445280 122400 1 0 $X=445090 $Y=119440
X2327 1 2 160 166 1445 ICV_36 $T=445280 149600 1 0 $X=445090 $Y=146640
X2328 1 2 1426 310 1464 ICV_36 $T=457240 160480 1 0 $X=457050 $Y=157520
X2329 1 2 1475 298 1492 ICV_36 $T=470120 160480 0 0 $X=469930 $Y=160240
X2330 1 2 1523 360 1541 ICV_36 $T=497260 149600 1 0 $X=497070 $Y=146640
X2331 1 2 1666 296 1684 ICV_36 $T=587420 149600 1 0 $X=587230 $Y=146640
X2332 1 2 1755 382 1764 ICV_36 $T=632960 171360 0 0 $X=632770 $Y=171120
X2333 1 2 1795 379 1801 ICV_36 $T=655500 171360 0 0 $X=655310 $Y=171120
X2334 1 2 1795 382 1826 ICV_36 $T=665620 171360 0 0 $X=665430 $Y=171120
X2335 1 2 1871 382 1883 ICV_36 $T=695060 171360 0 0 $X=694870 $Y=171120
X2336 1 2 44 9 670 ICV_37 $T=47840 133280 1 0 $X=47650 $Y=130320
X2337 1 2 666 27 681 ICV_37 $T=47840 160480 1 0 $X=47650 $Y=157520
X2338 1 2 664 28 684 ICV_37 $T=47840 176800 1 0 $X=47650 $Y=173840
X2339 1 2 675 5 703 ICV_37 $T=61640 116960 0 0 $X=61450 $Y=116720
X2340 1 2 685 26 704 ICV_37 $T=61640 133280 0 0 $X=61450 $Y=133040
X2341 1 2 685 27 705 ICV_37 $T=61640 138720 0 0 $X=61450 $Y=138480
X2342 1 2 685 8 707 ICV_37 $T=61640 144160 0 0 $X=61450 $Y=143920
X2343 1 2 664 26 708 ICV_37 $T=61640 176800 0 0 $X=61450 $Y=176560
X2344 1 2 701 8 728 ICV_37 $T=75900 160480 1 0 $X=75710 $Y=157520
X2345 1 2 726 6 755 ICV_37 $T=89700 138720 0 0 $X=89510 $Y=138480
X2346 1 2 745 27 759 ICV_37 $T=89700 160480 0 0 $X=89510 $Y=160240
X2347 1 2 761 28 789 ICV_37 $T=103960 138720 1 0 $X=103770 $Y=135760
X2348 1 2 745 9 784 ICV_37 $T=103960 160480 1 0 $X=103770 $Y=157520
X2349 1 2 791 5 820 ICV_37 $T=117760 171360 0 0 $X=117570 $Y=171120
X2350 1 2 837 9 847 ICV_37 $T=132020 149600 1 0 $X=131830 $Y=146640
X2351 1 2 829 6 849 ICV_37 $T=132020 155040 1 0 $X=131830 $Y=152080
X2352 1 2 829 27 850 ICV_37 $T=132020 160480 1 0 $X=131830 $Y=157520
X2353 1 2 791 8 839 ICV_37 $T=132020 171360 1 0 $X=131830 $Y=168400
X2354 1 2 100 26 873 ICV_37 $T=145820 122400 0 0 $X=145630 $Y=122160
X2355 1 2 837 27 871 ICV_37 $T=145820 144160 0 0 $X=145630 $Y=143920
X2356 1 2 829 29 878 ICV_37 $T=145820 155040 0 0 $X=145630 $Y=154800
X2357 1 2 884 29 907 ICV_37 $T=160080 144160 1 0 $X=159890 $Y=141200
X2358 1 2 884 9 881 ICV_37 $T=160080 149600 1 0 $X=159890 $Y=146640
X2359 1 2 876 6 903 ICV_37 $T=160080 160480 1 0 $X=159890 $Y=157520
X2360 1 2 906 5 931 ICV_37 $T=173880 116960 0 0 $X=173690 $Y=116720
X2361 1 2 876 28 937 ICV_37 $T=173880 155040 0 0 $X=173690 $Y=154800
X2362 1 2 928 27 962 ICV_37 $T=188140 133280 1 0 $X=187950 $Y=130320
X2363 1 2 1001 155 993 ICV_37 $T=216200 160480 1 0 $X=216010 $Y=157520
X2364 1 2 1001 178 1032 ICV_37 $T=230000 165920 0 0 $X=229810 $Y=165680
X2365 1 2 151 179 1034 ICV_37 $T=230000 176800 0 0 $X=229810 $Y=176560
X2366 1 2 1041 196 1056 ICV_37 $T=244260 127840 1 0 $X=244070 $Y=124880
X2367 1 2 1040 176 1052 ICV_37 $T=244260 171360 1 0 $X=244070 $Y=168400
X2368 1 2 1041 194 1072 ICV_37 $T=258060 133280 0 0 $X=257870 $Y=133040
X2369 1 2 1044 204 1080 ICV_37 $T=258060 144160 0 0 $X=257870 $Y=143920
X2370 1 2 1040 156 1071 ICV_37 $T=258060 165920 0 0 $X=257870 $Y=165680
X2371 1 2 1040 154 1073 ICV_37 $T=258060 171360 0 0 $X=257870 $Y=171120
X2372 1 2 215 153 1109 ICV_37 $T=272320 116960 1 0 $X=272130 $Y=114000
X2373 1 2 1075 196 1106 ICV_37 $T=272320 122400 1 0 $X=272130 $Y=119440
X2374 1 2 1075 194 1132 ICV_37 $T=286120 116960 0 0 $X=285930 $Y=116720
X2375 1 2 1133 196 1165 ICV_37 $T=300380 127840 1 0 $X=300190 $Y=124880
X2376 1 2 1148 193 1166 ICV_37 $T=300380 138720 1 0 $X=300190 $Y=135760
X2377 1 2 1148 197 1158 ICV_37 $T=300380 144160 1 0 $X=300190 $Y=141200
X2378 1 2 1153 179 1167 ICV_37 $T=300380 149600 1 0 $X=300190 $Y=146640
X2379 1 2 1156 156 1197 ICV_37 $T=314180 160480 0 0 $X=313990 $Y=160240
X2380 1 2 1156 154 1198 ICV_37 $T=314180 171360 0 0 $X=313990 $Y=171120
X2381 1 2 232 155 1215 ICV_37 $T=328440 122400 1 0 $X=328250 $Y=119440
X2382 1 2 1208 154 1227 ICV_37 $T=328440 149600 1 0 $X=328250 $Y=146640
X2383 1 2 1208 156 1217 ICV_37 $T=328440 155040 1 0 $X=328250 $Y=152080
X2384 1 2 1206 155 1213 ICV_37 $T=328440 165920 1 0 $X=328250 $Y=162960
X2385 1 2 1206 176 1223 ICV_37 $T=328440 171360 1 0 $X=328250 $Y=168400
X2386 1 2 235 178 1228 ICV_37 $T=328440 176800 1 0 $X=328250 $Y=173840
X2387 1 2 240 178 1256 ICV_37 $T=356500 116960 1 0 $X=356310 $Y=114000
X2388 1 2 1257 153 1279 ICV_37 $T=356500 122400 1 0 $X=356310 $Y=119440
X2389 1 2 1257 156 1304 ICV_37 $T=370300 122400 0 0 $X=370110 $Y=122160
X2390 1 2 1312 153 1329 ICV_37 $T=384560 127840 1 0 $X=384370 $Y=124880
X2391 1 2 1327 179 1355 ICV_37 $T=398360 171360 0 0 $X=398170 $Y=171120
X2392 1 2 269 176 280 ICV_37 $T=412620 116960 1 0 $X=412430 $Y=114000
X2393 1 2 1350 176 1381 ICV_37 $T=412620 160480 1 0 $X=412430 $Y=157520
X2394 1 2 1396 281 299 ICV_37 $T=426420 165920 0 0 $X=426230 $Y=165680
X2395 1 2 1395 196 1427 ICV_37 $T=440680 133280 1 0 $X=440490 $Y=130320
X2396 1 2 1396 310 315 ICV_37 $T=440680 165920 1 0 $X=440490 $Y=162960
X2397 1 2 1396 303 1424 ICV_37 $T=440680 171360 1 0 $X=440490 $Y=168400
X2398 1 2 1440 298 1453 ICV_37 $T=454480 122400 0 0 $X=454290 $Y=122160
X2399 1 2 1426 298 1450 ICV_37 $T=454480 160480 0 0 $X=454290 $Y=160240
X2400 1 2 1466 339 1478 ICV_37 $T=468740 144160 1 0 $X=468550 $Y=141200
X2401 1 2 1426 295 1477 ICV_37 $T=468740 155040 1 0 $X=468550 $Y=152080
X2402 1 2 335 283 364 ICV_37 $T=482540 171360 0 0 $X=482350 $Y=171120
X2403 1 2 1476 360 1528 ICV_37 $T=496800 127840 1 0 $X=496610 $Y=124880
X2404 1 2 160 371 1527 ICV_37 $T=496800 155040 1 0 $X=496610 $Y=152080
X2405 1 2 1548 283 1561 ICV_37 $T=510600 122400 0 0 $X=510410 $Y=122160
X2406 1 2 1547 310 1559 ICV_37 $T=510600 149600 0 0 $X=510410 $Y=149360
X2407 1 2 1547 303 1562 ICV_37 $T=510600 155040 0 0 $X=510410 $Y=154800
X2408 1 2 1547 283 1536 ICV_37 $T=510600 160480 0 0 $X=510410 $Y=160240
X2409 1 2 1588 343 1603 ICV_37 $T=538660 122400 0 0 $X=538470 $Y=122160
X2410 1 2 1588 338 1608 ICV_37 $T=538660 127840 0 0 $X=538470 $Y=127600
X2411 1 2 1580 388 1609 ICV_37 $T=538660 160480 0 0 $X=538470 $Y=160240
X2412 1 2 424 358 1629 ICV_37 $T=552920 116960 1 0 $X=552730 $Y=114000
X2413 1 2 1628 295 1650 ICV_37 $T=566720 122400 0 0 $X=566530 $Y=122160
X2414 1 2 1625 400 1647 ICV_37 $T=566720 160480 0 0 $X=566530 $Y=160240
X2415 1 2 428 399 1651 ICV_37 $T=566720 176800 0 0 $X=566530 $Y=176560
X2416 1 2 452 298 478 ICV_37 $T=580980 116960 1 0 $X=580790 $Y=114000
X2417 1 2 477 296 1686 ICV_37 $T=594780 116960 0 0 $X=594590 $Y=116720
X2418 1 2 1665 298 1689 ICV_37 $T=594780 127840 0 0 $X=594590 $Y=127600
X2419 1 2 1688 296 1731 ICV_37 $T=622840 149600 0 0 $X=622650 $Y=149360
X2420 1 2 1688 298 1741 ICV_37 $T=622840 155040 0 0 $X=622650 $Y=154800
X2421 1 2 519 281 524 ICV_37 $T=637100 116960 1 0 $X=636910 $Y=114000
X2422 1 2 519 295 1742 ICV_37 $T=637100 122400 1 0 $X=636910 $Y=119440
X2423 1 2 1749 295 1765 ICV_37 $T=637100 127840 1 0 $X=636910 $Y=124880
X2424 1 2 1748 303 1761 ICV_37 $T=637100 149600 1 0 $X=636910 $Y=146640
X2425 1 2 1748 283 1767 ICV_37 $T=637100 160480 1 0 $X=636910 $Y=157520
X2426 1 2 1755 395 1769 ICV_37 $T=637100 165920 1 0 $X=636910 $Y=162960
X2427 1 2 519 296 1793 ICV_37 $T=650900 116960 0 0 $X=650710 $Y=116720
X2428 1 2 1835 399 1850 ICV_37 $T=678960 171360 0 0 $X=678770 $Y=171120
X2429 1 2 1859 358 1875 ICV_37 $T=693220 144160 1 0 $X=693030 $Y=141200
X2430 1 2 1844 343 1897 ICV_37 $T=707020 127840 0 0 $X=706830 $Y=127600
X2431 1 2 1859 338 1903 ICV_37 $T=707020 144160 0 0 $X=706830 $Y=143920
X2432 1 2 545 358 548 ICV_37 $T=721280 116960 1 0 $X=721090 $Y=114000
X2433 1 2 1904 340 1937 ICV_37 $T=721280 127840 1 0 $X=721090 $Y=124880
X2434 1 2 1916 339 1926 ICV_37 $T=721280 138720 1 0 $X=721090 $Y=135760
X2435 1 2 1916 358 1934 ICV_37 $T=721280 144160 1 0 $X=721090 $Y=141200
X2436 1 2 1918 340 1939 ICV_37 $T=721280 149600 1 0 $X=721090 $Y=146640
X2437 1 2 1918 358 1940 ICV_37 $T=721280 155040 1 0 $X=721090 $Y=152080
X2438 1 2 1919 399 1941 ICV_37 $T=721280 171360 1 0 $X=721090 $Y=168400
X2439 1 2 545 360 552 ICV_37 $T=735080 116960 0 0 $X=734890 $Y=116720
X2440 1 2 1904 341 1956 ICV_37 $T=735080 127840 0 0 $X=734890 $Y=127600
X2441 1 2 1916 357 1942 ICV_37 $T=735080 133280 0 0 $X=734890 $Y=133040
X2442 1 2 1916 338 1943 ICV_37 $T=735080 138720 0 0 $X=734890 $Y=138480
X2443 1 2 1918 360 1958 ICV_37 $T=735080 149600 0 0 $X=734890 $Y=149360
X2444 1 2 1918 338 1944 ICV_37 $T=735080 155040 0 0 $X=734890 $Y=154800
X2445 1 2 788 8 801 788 9 781 ICV_38 $T=108560 133280 1 0 $X=108370 $Y=130320
X2446 1 2 791 29 806 791 27 815 ICV_38 $T=109020 165920 1 0 $X=108830 $Y=162960
X2447 1 2 843 9 875 843 8 887 ICV_38 $T=145360 165920 1 0 $X=145170 $Y=162960
X2448 1 2 884 28 902 884 5 915 ICV_38 $T=157320 144160 0 0 $X=157130 $Y=143920
X2449 1 2 125 8 127 125 27 960 ICV_38 $T=184920 176800 0 0 $X=184730 $Y=176560
X2450 1 2 932 5 972 932 6 976 ICV_38 $T=195500 122400 1 0 $X=195310 $Y=119440
X2451 1 2 1108 205 1130 1108 213 1146 ICV_38 $T=282900 144160 1 0 $X=282710 $Y=141200
X2452 1 2 1206 179 1243 1206 154 1242 ICV_38 $T=336260 171360 1 0 $X=336070 $Y=168400
X2453 1 2 1248 155 1258 1248 154 1273 ICV_38 $T=345000 133280 0 0 $X=344810 $Y=133040
X2454 1 2 1248 179 1292 1248 156 1296 ICV_38 $T=361560 133280 1 0 $X=361370 $Y=130320
X2455 1 2 1303 155 1352 1349 179 1362 ICV_38 $T=396980 144160 1 0 $X=396790 $Y=141200
X2456 1 2 160 188 1421 160 185 1435 ICV_38 $T=436080 155040 0 0 $X=435890 $Y=154800
X2457 1 2 1398 204 1425 160 189 1441 ICV_38 $T=439760 149600 0 0 $X=439570 $Y=149360
X2458 1 2 160 167 1434 1426 281 1448 ICV_38 $T=443440 155040 1 0 $X=443250 $Y=152080
X2459 1 2 1524 388 1549 1524 395 1568 ICV_38 $T=506920 165920 1 0 $X=506730 $Y=162960
X2460 1 2 1626 340 1610 1626 341 1659 ICV_38 $T=563960 138720 1 0 $X=563770 $Y=135760
X2461 1 2 1666 307 1705 1666 310 1714 ICV_38 $T=603520 144160 0 0 $X=603330 $Y=143920
X2462 1 2 621 605 37 ICV_39 $T=28520 138720 0 0 $X=28330 $Y=138480
X2463 1 2 673 683 38 ICV_39 $T=56580 165920 0 0 $X=56390 $Y=165680
X2464 1 2 86 84 32 ICV_39 $T=112700 176800 0 0 $X=112510 $Y=176560
X2465 1 2 823 93 38 ICV_39 $T=126960 176800 1 0 $X=126770 $Y=173840
X2466 1 2 854 844 32 ICV_39 $T=140760 127840 0 0 $X=140570 $Y=127600
X2467 1 2 871 851 37 ICV_39 $T=149500 149600 1 0 $X=149310 $Y=146640
X2468 1 2 857 851 19 ICV_39 $T=155020 138720 1 0 $X=154830 $Y=135760
X2469 1 2 849 844 19 ICV_39 $T=155020 160480 1 0 $X=154830 $Y=157520
X2470 1 2 123 117 37 ICV_39 $T=179860 176800 0 0 $X=179670 $Y=176560
X2471 1 2 958 969 19 ICV_39 $T=198720 155040 1 0 $X=198530 $Y=152080
X2472 1 2 977 951 40 ICV_39 $T=203320 127840 0 0 $X=203130 $Y=127600
X2473 1 2 985 950 11 ICV_39 $T=211140 138720 1 0 $X=210950 $Y=135760
X2474 1 2 1055 1042 201 ICV_39 $T=250700 155040 1 0 $X=250510 $Y=152080
X2475 1 2 1070 1047 216 ICV_39 $T=259440 127840 0 0 $X=259250 $Y=127600
X2476 1 2 1074 1054 166 ICV_39 $T=267260 165920 1 0 $X=267070 $Y=162960
X2477 1 2 1115 1102 150 ICV_39 $T=287040 165920 1 0 $X=286850 $Y=162960
X2478 1 2 1128 1097 201 ICV_39 $T=287500 127840 0 0 $X=287310 $Y=127600
X2479 1 2 1127 1094 201 ICV_39 $T=288420 122400 0 0 $X=288230 $Y=122160
X2480 1 2 1146 1117 211 ICV_39 $T=298540 144160 0 0 $X=298350 $Y=143920
X2481 1 2 1198 1161 167 ICV_39 $T=322920 165920 0 0 $X=322730 $Y=165680
X2482 1 2 1210 1191 185 ICV_39 $T=329820 138720 1 0 $X=329630 $Y=135760
X2483 1 2 1247 239 166 ICV_39 $T=344080 176800 0 0 $X=343890 $Y=176560
X2484 1 2 1328 259 188 ICV_39 $T=386400 133280 1 0 $X=386210 $Y=130320
X2485 1 2 1336 1324 167 ICV_39 $T=393300 155040 0 0 $X=393110 $Y=154800
X2486 1 2 1342 1326 189 ICV_39 $T=403420 149600 1 0 $X=403230 $Y=146640
X2487 1 2 1399 293 188 ICV_39 $T=429180 116960 0 0 $X=428990 $Y=116720
X2488 1 2 317 318 150 ICV_39 $T=449420 116960 1 0 $X=449230 $Y=114000
X2489 1 2 1464 1449 325 ICV_39 $T=466440 165920 0 0 $X=466250 $Y=165680
X2490 1 2 1571 1538 300 ICV_39 $T=529920 149600 1 0 $X=529730 $Y=146640
X2491 1 2 1685 1682 407 ICV_39 $T=597540 176800 1 0 $X=597350 $Y=173840
X2492 1 2 1691 1672 300 ICV_39 $T=603980 127840 1 0 $X=603790 $Y=124880
X2493 1 2 493 491 455 ICV_39 $T=603980 176800 1 0 $X=603790 $Y=173840
X2494 1 2 525 517 316 ICV_39 $T=645840 116960 0 0 $X=645650 $Y=116720
X2495 1 2 1766 1763 300 ICV_39 $T=645840 127840 0 0 $X=645650 $Y=127600
X2496 1 2 528 517 294 ICV_39 $T=660100 116960 1 0 $X=659910 $Y=114000
X2497 1 2 1832 1837 365 ICV_39 $T=679420 144160 1 0 $X=679230 $Y=141200
X2498 1 2 1950 1920 345 ICV_39 $T=737840 122400 0 0 $X=737650 $Y=122160
X2499 1 2 1954 1921 356 ICV_39 $T=737840 144160 0 0 $X=737650 $Y=143920
X2500 1 2 1945 1928 423 ICV_39 $T=737840 160480 1 0 $X=737650 $Y=157520
X2501 1 2 1955 1928 409 ICV_39 $T=737840 160480 0 0 $X=737650 $Y=160240
X2502 1 2 1946 1928 396 ICV_39 $T=737840 165920 0 0 $X=737650 $Y=165680
X2503 1 2 669 48 40 ICV_40 $T=51520 122400 1 0 $X=51330 $Y=119440
X2504 1 2 694 695 37 ICV_40 $T=64860 127840 0 0 $X=64670 $Y=127600
X2505 1 2 743 744 40 ICV_40 $T=86480 144160 1 0 $X=86290 $Y=141200
X2506 1 2 750 752 37 ICV_40 $T=90620 165920 0 0 $X=90430 $Y=165680
X2507 1 2 759 760 37 ICV_40 $T=93840 165920 1 0 $X=93650 $Y=162960
X2508 1 2 916 927 11 ICV_40 $T=176640 127840 0 0 $X=176450 $Y=127600
X2509 1 2 925 927 37 ICV_40 $T=177100 133280 0 0 $X=176910 $Y=133040
X2510 1 2 926 927 38 ICV_40 $T=182160 116960 1 0 $X=181970 $Y=114000
X2511 1 2 937 892 40 ICV_40 $T=182160 155040 1 0 $X=181970 $Y=152080
X2512 1 2 1032 995 189 ICV_40 $T=247940 165920 0 0 $X=247750 $Y=165680
X2513 1 2 208 195 167 ICV_40 $T=255300 116960 1 0 $X=255110 $Y=114000
X2514 1 2 1068 1047 214 ICV_40 $T=258980 138720 1 0 $X=258790 $Y=135760
X2515 1 2 1098 1097 214 ICV_40 $T=273240 138720 1 0 $X=273050 $Y=135760
X2516 1 2 1110 1097 203 ICV_40 $T=280140 133280 0 0 $X=279950 $Y=133040
X2517 1 2 1129 1097 210 ICV_40 $T=287500 133280 0 0 $X=287310 $Y=133040
X2518 1 2 1149 1142 216 ICV_40 $T=299000 127840 0 0 $X=298810 $Y=127600
X2519 1 2 1167 1163 188 ICV_40 $T=308200 149600 0 0 $X=308010 $Y=149360
X2520 1 2 1182 1160 216 ICV_40 $T=315560 138720 0 0 $X=315370 $Y=138480
X2521 1 2 1220 1214 166 ICV_40 $T=336260 165920 0 0 $X=336070 $Y=165680
X2522 1 2 1246 1218 186 ICV_40 $T=344080 155040 0 0 $X=343890 $Y=154800
X2523 1 2 1313 258 185 ICV_40 $T=380420 165920 0 0 $X=380230 $Y=165680
X2524 1 2 1316 258 186 ICV_40 $T=381340 171360 0 0 $X=381150 $Y=171120
X2525 1 2 1505 1490 325 ICV_40 $T=492660 155040 0 0 $X=492470 $Y=154800
X2526 1 2 1517 1487 356 ICV_40 $T=494040 138720 0 0 $X=493850 $Y=138480
X2527 1 2 1608 1604 345 ICV_40 $T=546940 133280 1 0 $X=546750 $Y=130320
X2528 1 2 1609 1600 396 ICV_40 $T=546940 160480 1 0 $X=546750 $Y=157520
X2529 1 2 1622 1604 342 ICV_40 $T=553840 122400 1 0 $X=553650 $Y=119440
X2530 1 2 1633 1602 344 ICV_40 $T=560740 144160 0 0 $X=560550 $Y=143920
X2531 1 2 1647 1638 423 ICV_40 $T=569940 165920 0 0 $X=569750 $Y=165680
X2532 1 2 1723 488 294 ICV_40 $T=622380 116960 1 0 $X=622190 $Y=114000
X2533 1 2 1790 517 309 ICV_40 $T=659180 122400 1 0 $X=658990 $Y=119440
X2534 1 2 532 533 351 ICV_40 $T=672980 116960 0 0 $X=672790 $Y=116720
X2535 1 2 1896 1866 371 ICV_40 $T=709320 122400 0 0 $X=709130 $Y=122160
X2536 1 2 666 6 697 ICV_43 $T=64860 160480 1 0 $X=64670 $Y=157520
X2537 1 2 106 6 901 ICV_43 $T=156400 176800 0 0 $X=156210 $Y=176560
X2538 1 2 876 29 908 ICV_43 $T=162840 155040 0 0 $X=162650 $Y=154800
X2539 1 2 928 8 952 ICV_43 $T=183080 133280 0 0 $X=182890 $Y=133040
X2540 1 2 125 6 971 ICV_43 $T=190900 171360 0 0 $X=190710 $Y=171120
X2541 1 2 183 156 1045 ICV_43 $T=237360 116960 0 0 $X=237170 $Y=116720
X2542 1 2 1044 196 1061 ICV_43 $T=247020 144160 1 0 $X=246830 $Y=141200
X2543 1 2 215 154 220 ICV_43 $T=261280 116960 1 0 $X=261090 $Y=114000
X2544 1 2 1153 178 1203 ICV_43 $T=317400 160480 1 0 $X=317210 $Y=157520
X2545 1 2 240 155 1251 ICV_43 $T=345460 116960 1 0 $X=345270 $Y=114000
X2546 1 2 1257 175 1278 ICV_43 $T=359260 122400 0 0 $X=359070 $Y=122160
X2547 1 2 1327 156 1337 ICV_43 $T=387320 171360 0 0 $X=387130 $Y=171120
X2548 1 2 1312 155 267 ICV_43 $T=392380 127840 1 0 $X=392190 $Y=124880
X2549 1 2 1398 197 1409 ICV_43 $T=429640 138720 1 0 $X=429450 $Y=135760
X2550 1 2 1580 380 1614 ICV_43 $T=541880 171360 1 0 $X=541690 $Y=168400
X2551 1 2 1628 307 1645 ICV_43 $T=561200 127840 1 0 $X=561010 $Y=124880
X2552 1 2 1918 341 1957 ICV_43 $T=731860 149600 1 0 $X=731670 $Y=146640
X2553 1 2 1918 357 1954 ICV_43 $T=731860 155040 1 0 $X=731670 $Y=152080
X2554 1 2 1919 380 1955 ICV_43 $T=731860 171360 1 0 $X=731670 $Y=168400
X2555 1 2 4 7 12 ICV_47 $T=6900 116960 1 0 $X=6710 $Y=114000
X2556 1 2 584 8 596 ICV_47 $T=6900 144160 0 0 $X=6710 $Y=143920
X2557 1 2 584 6 597 ICV_47 $T=6900 149600 0 0 $X=6710 $Y=149360
X2558 1 2 583 29 629 ICV_47 $T=22540 116960 0 0 $X=22350 $Y=116720
X2559 1 2 675 28 688 ICV_47 $T=52900 122400 0 0 $X=52710 $Y=122160
X2560 1 2 685 29 693 ICV_47 $T=54740 149600 1 0 $X=54550 $Y=146640
X2561 1 2 666 26 699 ICV_47 $T=57500 155040 1 0 $X=57310 $Y=152080
X2562 1 2 685 5 716 ICV_47 $T=63480 138720 1 0 $X=63290 $Y=135760
X2563 1 2 702 8 730 ICV_47 $T=75440 122400 0 0 $X=75250 $Y=122160
X2564 1 2 729 27 750 ICV_47 $T=80960 165920 0 0 $X=80770 $Y=165680
X2565 1 2 726 29 765 ICV_47 $T=90160 144160 0 0 $X=89970 $Y=143920
X2566 1 2 89 29 823 ICV_47 $T=118220 176800 0 0 $X=118030 $Y=176560
X2567 1 2 816 9 830 ICV_47 $T=122360 127840 0 0 $X=122170 $Y=127600
X2568 1 2 837 6 857 ICV_47 $T=133400 138720 0 0 $X=133210 $Y=138480
X2569 1 2 106 28 110 ICV_47 $T=147660 176800 0 0 $X=147470 $Y=176560
X2570 1 2 898 28 913 ICV_47 $T=161920 171360 0 0 $X=161730 $Y=171120
X2571 1 2 884 26 917 ICV_47 $T=165140 138720 0 0 $X=164950 $Y=138480
X2572 1 2 932 26 945 ICV_47 $T=179400 122400 1 0 $X=179210 $Y=119440
X2573 1 2 933 26 943 ICV_47 $T=181700 155040 0 0 $X=181510 $Y=154800
X2574 1 2 125 26 955 ICV_47 $T=182160 171360 0 0 $X=181970 $Y=171120
X2575 1 2 933 6 970 ICV_47 $T=188600 165920 1 0 $X=188410 $Y=162960
X2576 1 2 1124 179 1134 ICV_47 $T=284280 160480 1 0 $X=284090 $Y=157520
X2577 1 2 1133 205 1174 ICV_47 $T=302220 122400 1 0 $X=302030 $Y=119440
X2578 1 2 1153 155 1186 ICV_47 $T=309580 149600 1 0 $X=309390 $Y=146640
X2579 1 2 1187 193 1204 ICV_47 $T=319700 127840 1 0 $X=319510 $Y=124880
X2580 1 2 1208 155 1225 ICV_47 $T=326140 155040 0 0 $X=325950 $Y=154800
X2581 1 2 235 153 1247 ICV_47 $T=336260 176800 1 0 $X=336070 $Y=173840
X2582 1 2 1248 176 1263 ICV_47 $T=346380 138720 1 0 $X=346190 $Y=135760
X2583 1 2 1253 175 1267 ICV_47 $T=347760 165920 1 0 $X=347570 $Y=162960
X2584 1 2 243 153 1280 ICV_47 $T=356960 171360 1 0 $X=356770 $Y=168400
X2585 1 2 1301 156 1317 ICV_47 $T=373520 149600 1 0 $X=373330 $Y=146640
X2586 1 2 1301 179 1333 ICV_47 $T=385020 149600 1 0 $X=384830 $Y=146640
X2587 1 2 1354 178 1369 ICV_47 $T=402960 133280 1 0 $X=402770 $Y=130320
X2588 1 2 1377 155 285 ICV_47 $T=417680 116960 0 0 $X=417490 $Y=116720
X2589 1 2 1395 206 1405 ICV_47 $T=426880 127840 1 0 $X=426690 $Y=124880
X2590 1 2 1398 213 1411 ICV_47 $T=430100 144160 1 0 $X=429910 $Y=141200
X2591 1 2 1426 307 1442 ICV_47 $T=445740 160480 0 0 $X=445550 $Y=160240
X2592 1 2 314 303 1438 ICV_47 $T=445740 171360 0 0 $X=445550 $Y=171120
X2593 1 2 314 296 1443 ICV_47 $T=445740 176800 0 0 $X=445550 $Y=176560
X2594 1 2 313 303 1463 ICV_47 $T=458620 116960 1 0 $X=458430 $Y=114000
X2595 1 2 1476 341 1494 ICV_47 $T=472420 116960 0 0 $X=472230 $Y=116720
X2596 1 2 160 345 1499 ICV_47 $T=473800 155040 0 0 $X=473610 $Y=154800
X2597 1 2 1466 358 1510 ICV_47 $T=483000 138720 0 0 $X=482810 $Y=138480
X2598 1 2 1523 338 1546 ICV_47 $T=500480 144160 0 0 $X=500290 $Y=143920
X2599 1 2 1580 382 1595 ICV_47 $T=529460 171360 1 0 $X=529270 $Y=168400
X2600 1 2 1580 400 1619 ICV_47 $T=543260 165920 1 0 $X=543070 $Y=162960
X2601 1 2 1588 340 1623 ICV_47 $T=546480 122400 0 0 $X=546290 $Y=122160
X2602 1 2 428 400 1632 ICV_47 $T=552460 171360 0 0 $X=552270 $Y=171120
X2603 1 2 1625 378 1636 ICV_47 $T=554760 165920 0 0 $X=554570 $Y=165680
X2604 1 2 1625 388 1642 ICV_47 $T=557980 160480 0 0 $X=557790 $Y=160240
X2605 1 2 452 307 458 ICV_47 $T=560740 116960 1 0 $X=560550 $Y=114000
X2606 1 2 1628 298 1661 ICV_47 $T=574540 122400 0 0 $X=574350 $Y=122160
X2607 1 2 477 307 1678 ICV_47 $T=586040 116960 0 0 $X=585850 $Y=116720
X2608 1 2 1710 395 1721 ICV_47 $T=613180 165920 0 0 $X=612990 $Y=165680
X2609 1 2 1710 382 1727 ICV_47 $T=613640 171360 1 0 $X=613450 $Y=168400
X2610 1 2 1688 281 1730 ICV_47 $T=614560 155040 1 0 $X=614370 $Y=152080
X2611 1 2 1818 357 1829 ICV_47 $T=669760 155040 0 0 $X=669570 $Y=154800
X2612 1 2 529 338 1830 ICV_47 $T=670220 122400 0 0 $X=670030 $Y=122160
X2613 1 2 536 378 542 ICV_47 $T=694600 176800 0 0 $X=694410 $Y=176560
X2614 1 2 1904 339 1930 ICV_47 $T=717140 127840 0 0 $X=716950 $Y=127600
X2615 1 2 35 15 32 ICV_48 $T=29440 176800 0 0 $X=29250 $Y=176560
X2616 1 2 740 741 19 ICV_48 $T=85560 122400 0 0 $X=85370 $Y=122160
X2617 1 2 769 752 19 ICV_48 $T=99820 165920 1 0 $X=99630 $Y=162960
X2618 1 2 799 790 21 ICV_48 $T=113620 144160 0 0 $X=113430 $Y=143920
X2619 1 2 94 96 95 ICV_48 $T=127880 116960 1 0 $X=127690 $Y=114000
X2620 1 2 972 951 20 ICV_48 $T=197800 116960 0 0 $X=197610 $Y=116720
X2621 1 2 1034 163 188 ICV_48 $T=240120 176800 1 0 $X=239930 $Y=173840
X2622 1 2 1062 1042 211 ICV_48 $T=253920 155040 0 0 $X=253730 $Y=154800
X2623 1 2 1113 1094 211 ICV_48 $T=281980 127840 0 0 $X=281790 $Y=127600
X2624 1 2 1114 1117 210 ICV_48 $T=281980 138720 0 0 $X=281790 $Y=138480
X2625 1 2 226 227 150 ICV_48 $T=296240 122400 1 0 $X=296050 $Y=119440
X2626 1 2 1173 1142 211 ICV_48 $T=310040 116960 0 0 $X=309850 $Y=116720
X2627 1 2 1176 1161 150 ICV_48 $T=310040 155040 0 0 $X=309850 $Y=154800
X2628 1 2 1258 1261 150 ICV_48 $T=352360 133280 1 0 $X=352170 $Y=130320
X2629 1 2 1259 244 162 ICV_48 $T=352360 171360 1 0 $X=352170 $Y=168400
X2630 1 2 1282 1276 189 ICV_48 $T=366160 144160 0 0 $X=365970 $Y=143920
X2631 1 2 1283 1284 150 ICV_48 $T=366160 171360 0 0 $X=365970 $Y=171120
X2632 1 2 1314 258 188 ICV_48 $T=380420 176800 1 0 $X=380230 $Y=173840
X2633 1 2 1362 1360 188 ICV_48 $T=408480 149600 1 0 $X=408290 $Y=146640
X2634 1 2 1411 1410 211 ICV_48 $T=436540 155040 1 0 $X=436350 $Y=152080
X2635 1 2 1436 319 320 ICV_48 $T=450340 165920 0 0 $X=450150 $Y=165680
X2636 1 2 1488 1473 354 ICV_48 $T=478400 138720 0 0 $X=478210 $Y=138480
X2637 1 2 1518 361 344 ICV_48 $T=506460 116960 0 0 $X=506270 $Y=116720
X2638 1 2 1539 386 391 ICV_48 $T=506460 165920 0 0 $X=506270 $Y=165680
X2639 1 2 454 443 455 ICV_48 $T=562580 171360 0 0 $X=562390 $Y=171120
X2640 1 2 1801 1804 444 ICV_48 $T=661020 176800 1 0 $X=660830 $Y=173840
X2641 1 2 1858 537 354 ICV_48 $T=689080 116960 1 0 $X=688890 $Y=114000
X2642 1 2 623 599 32 44 26 644 ICV_51 $T=33580 127840 1 0 $X=33390 $Y=124880
X2643 1 2 725 66 37 62 5 748 ICV_51 $T=77280 176800 1 0 $X=77090 $Y=173840
X2644 1 2 755 744 19 761 26 776 ICV_51 $T=92460 144160 1 0 $X=92270 $Y=141200
X2645 1 2 840 814 40 843 5 862 ICV_51 $T=133860 165920 1 0 $X=133670 $Y=162960
X2646 1 2 996 997 150 1002 155 996 ICV_51 $T=212520 149600 0 0 $X=212330 $Y=149360
X2647 1 2 1049 1047 200 1041 204 1049 ICV_51 $T=246560 127840 0 0 $X=246370 $Y=127600
X2648 1 2 1072 1047 210 1077 196 1089 ICV_51 $T=260820 133280 1 0 $X=260630 $Y=130320
X2649 1 2 1139 1142 200 1148 194 1159 ICV_51 $T=293480 133280 0 0 $X=293290 $Y=133040
X2650 1 2 1162 1163 166 1153 175 1184 ICV_51 $T=305900 160480 1 0 $X=305710 $Y=157520
X2651 1 2 1186 1163 150 1192 155 1212 ICV_51 $T=317400 144160 0 0 $X=317210 $Y=143920
X2652 1 2 1251 241 150 1257 179 1271 ICV_51 $T=347760 122400 0 0 $X=347570 $Y=122160
X2653 1 2 1497 1473 356 160 342 1512 ICV_51 $T=481620 149600 1 0 $X=481430 $Y=146640
X2654 1 2 1549 386 396 1524 399 1566 ICV_51 $T=509680 171360 1 0 $X=509490 $Y=168400
X2655 1 2 1550 393 397 392 382 1567 ICV_51 $T=509680 176800 1 0 $X=509490 $Y=173840
X2656 1 2 1601 1602 365 1606 360 1601 ICV_51 $T=540040 149600 0 0 $X=539850 $Y=149360
X2657 1 2 442 443 445 428 395 1640 ICV_51 $T=553380 176800 0 0 $X=553190 $Y=176560
X2658 1 2 1648 463 320 1665 310 1673 ICV_51 $T=581440 127840 0 0 $X=581250 $Y=127600
X2659 1 2 1740 1743 320 1748 295 1740 ICV_51 $T=629740 144160 0 0 $X=629550 $Y=143920
X2660 1 2 1839 537 344 538 339 1839 ICV_51 $T=681720 122400 1 0 $X=681530 $Y=119440
X2661 1 2 1840 1841 407 1835 379 1863 ICV_51 $T=681720 171360 1 0 $X=681530 $Y=168400
X2662 1 2 1854 1837 344 1859 357 1872 ICV_51 $T=687240 144160 0 0 $X=687050 $Y=143920
X2663 1 2 1910 1891 423 1919 379 1935 ICV_51 $T=715760 165920 0 0 $X=715570 $Y=165680
X2664 1 2 708 683 32 ICV_52 $T=70380 176800 1 0 $X=70190 $Y=173840
X2665 1 2 693 710 38 ICV_52 $T=72680 149600 0 0 $X=72490 $Y=149360
X2666 1 2 766 752 38 ICV_52 $T=98440 176800 1 0 $X=98250 $Y=173840
X2667 1 2 880 851 32 ICV_52 $T=154560 149600 1 0 $X=154370 $Y=146640
X2668 1 2 960 128 37 ICV_52 $T=191360 176800 1 0 $X=191170 $Y=173840
X2669 1 2 1061 1042 207 ICV_52 $T=253460 138720 1 0 $X=253270 $Y=135760
X2670 1 2 1203 1163 189 ICV_52 $T=327980 149600 0 0 $X=327790 $Y=149360
X2671 1 2 1355 1284 188 ICV_52 $T=404340 176800 0 0 $X=404150 $Y=176560
X2672 1 2 1409 1410 203 ICV_52 $T=436080 144160 0 0 $X=435890 $Y=143920
X2673 1 2 1447 1449 294 ICV_52 $T=456780 155040 0 0 $X=456590 $Y=154800
X2674 1 2 1575 1538 309 ICV_52 $T=541420 160480 1 0 $X=541230 $Y=157520
X2675 1 2 1635 1602 342 ICV_52 $T=575460 149600 1 0 $X=575270 $Y=146640
X2676 1 2 1657 1596 354 ICV_52 $T=576840 138720 0 0 $X=576650 $Y=138480
X2677 1 2 1684 1679 304 ICV_52 $T=596620 144160 0 0 $X=596430 $Y=143920
X2678 1 2 1681 1672 309 ICV_52 $T=598460 127840 1 0 $X=598270 $Y=124880
X2679 1 2 1757 1743 300 ICV_52 $T=645380 149600 0 0 $X=645190 $Y=149360
X2680 1 2 1848 1824 356 ICV_52 $T=687700 138720 1 0 $X=687510 $Y=135760
X2681 1 2 1862 1866 365 ICV_52 $T=695060 116960 1 0 $X=694870 $Y=114000
X2682 1 2 1915 1892 371 ICV_52 $T=718060 144160 0 0 $X=717870 $Y=143920
X2683 1 2 1947 546 423 ICV_52 $T=737380 171360 0 0 $X=737190 $Y=171120
X2684 1 2 550 546 396 ICV_52 $T=737380 176800 0 0 $X=737190 $Y=176560
X2685 1 2 ICV_54 $T=19780 127840 1 0 $X=19590 $Y=124880
X2686 1 2 ICV_54 $T=33580 122400 0 0 $X=33390 $Y=122160
X2687 1 2 ICV_54 $T=33580 138720 0 0 $X=33390 $Y=138480
X2688 1 2 ICV_54 $T=61640 122400 0 0 $X=61450 $Y=122160
X2689 1 2 ICV_54 $T=61640 155040 0 0 $X=61450 $Y=154800
X2690 1 2 ICV_54 $T=75900 144160 1 0 $X=75710 $Y=141200
X2691 1 2 ICV_54 $T=132020 138720 1 0 $X=131830 $Y=135760
X2692 1 2 ICV_54 $T=286120 122400 0 0 $X=285930 $Y=122160
X2693 1 2 ICV_54 $T=328440 160480 1 0 $X=328250 $Y=157520
X2694 1 2 ICV_54 $T=342240 160480 0 0 $X=342050 $Y=160240
X2695 1 2 ICV_54 $T=426420 160480 0 0 $X=426230 $Y=160240
X2696 1 2 ICV_54 $T=454480 155040 0 0 $X=454290 $Y=154800
X2697 1 2 ICV_54 $T=538660 116960 0 0 $X=538470 $Y=116720
X2698 1 2 ICV_54 $T=566720 144160 0 0 $X=566530 $Y=143920
X2699 1 2 ICV_54 $T=609040 127840 1 0 $X=608850 $Y=124880
X2700 1 2 ICV_54 $T=735080 171360 0 0 $X=734890 $Y=171120
X2701 1 2 3 2 14 1 sky130_fd_sc_hd__clkbuf_16 $T=6900 127840 0 0 $X=6710 $Y=127600
X2702 1 2 10 2 25 1 sky130_fd_sc_hd__clkbuf_16 $T=13340 116960 0 0 $X=13150 $Y=116720
X2703 1 2 82 2 88 1 sky130_fd_sc_hd__clkbuf_16 $T=109940 171360 1 0 $X=109750 $Y=168400
X2704 1 2 144 2 147 1 sky130_fd_sc_hd__clkbuf_16 $T=204240 116960 0 0 $X=204050 $Y=116720
X2705 1 2 145 2 148 1 sky130_fd_sc_hd__clkbuf_16 $T=207000 116960 1 0 $X=206810 $Y=114000
X2706 1 2 149 2 158 1 sky130_fd_sc_hd__clkbuf_16 $T=213440 116960 0 0 $X=213250 $Y=116720
X2707 1 2 157 2 165 1 sky130_fd_sc_hd__clkbuf_16 $T=218040 116960 1 0 $X=217850 $Y=114000
X2708 1 2 159 2 169 1 sky130_fd_sc_hd__clkbuf_16 $T=220340 127840 0 0 $X=220150 $Y=127600
X2709 1 2 164 2 180 1 sky130_fd_sc_hd__clkbuf_16 $T=223560 122400 1 0 $X=223370 $Y=119440
X2710 1 2 171 2 7 1 sky130_fd_sc_hd__clkbuf_16 $T=227240 116960 1 0 $X=227050 $Y=114000
X2711 1 2 181 2 34 1 sky130_fd_sc_hd__clkbuf_16 $T=233680 138720 0 0 $X=233490 $Y=138480
X2712 1 2 187 2 191 1 sky130_fd_sc_hd__clkbuf_16 $T=240580 160480 0 0 $X=240390 $Y=160240
X2713 1 2 256 2 197 1 sky130_fd_sc_hd__clkbuf_16 $T=374440 160480 1 0 $X=374250 $Y=157520
X2714 1 2 262 2 206 1 sky130_fd_sc_hd__clkbuf_16 $T=385020 160480 1 0 $X=384830 $Y=157520
X2715 1 2 275 2 179 1 sky130_fd_sc_hd__clkbuf_16 $T=408480 171360 0 0 $X=408290 $Y=171120
X2716 1 2 276 2 175 1 sky130_fd_sc_hd__clkbuf_16 $T=409860 176800 0 0 $X=409670 $Y=176560
X2717 1 2 278 2 153 1 sky130_fd_sc_hd__clkbuf_16 $T=413080 176800 1 0 $X=412890 $Y=173840
X2718 1 2 282 2 196 1 sky130_fd_sc_hd__clkbuf_16 $T=421820 160480 1 0 $X=421630 $Y=157520
X2719 1 2 284 2 193 1 sky130_fd_sc_hd__clkbuf_16 $T=425500 155040 1 0 $X=425310 $Y=152080
X2720 1 2 287 2 204 1 sky130_fd_sc_hd__clkbuf_16 $T=426880 149600 0 0 $X=426690 $Y=149360
X2721 1 2 288 2 213 1 sky130_fd_sc_hd__clkbuf_16 $T=426880 155040 0 0 $X=426690 $Y=154800
X2722 1 2 297 2 194 1 sky130_fd_sc_hd__clkbuf_16 $T=430100 149600 1 0 $X=429910 $Y=146640
X2723 1 2 326 2 332 1 sky130_fd_sc_hd__clkbuf_16 $T=458160 144160 0 0 $X=457970 $Y=143920
X2724 1 2 187 2 370 1 sky130_fd_sc_hd__clkbuf_16 $T=487600 171360 1 0 $X=487410 $Y=168400
X2725 1 2 282 2 382 1 sky130_fd_sc_hd__clkbuf_16 $T=494500 176800 0 0 $X=494310 $Y=176560
X2726 1 2 284 2 379 1 sky130_fd_sc_hd__clkbuf_16 $T=497260 176800 1 0 $X=497070 $Y=173840
X2727 1 2 390 2 1552 1 sky130_fd_sc_hd__clkbuf_16 $T=510140 133280 1 0 $X=509950 $Y=130320
X2728 1 2 394 2 1553 1 sky130_fd_sc_hd__clkbuf_16 $T=511060 127840 0 0 $X=510870 $Y=127600
X2729 1 2 403 2 1556 1 sky130_fd_sc_hd__clkbuf_16 $T=520260 127840 0 0 $X=520070 $Y=127600
X2730 1 2 287 2 400 1 sky130_fd_sc_hd__clkbuf_16 $T=529460 171360 0 0 $X=529270 $Y=171120
X2731 1 2 450 2 343 1 sky130_fd_sc_hd__clkbuf_16 $T=560280 160480 1 0 $X=560090 $Y=157520
X2732 1 2 275 2 358 1 sky130_fd_sc_hd__clkbuf_16 $T=595240 155040 0 0 $X=595050 $Y=154800
X2733 1 2 497 2 338 1 sky130_fd_sc_hd__clkbuf_16 $T=609500 160480 1 0 $X=609310 $Y=157520
X2734 1 2 276 2 357 1 sky130_fd_sc_hd__clkbuf_16 $T=651360 155040 0 0 $X=651170 $Y=154800
X2735 1 2 526 2 339 1 sky130_fd_sc_hd__clkbuf_16 $T=655960 155040 1 0 $X=655770 $Y=152080
X2736 1 2 278 2 340 1 sky130_fd_sc_hd__clkbuf_16 $T=660560 155040 0 0 $X=660370 $Y=154800
X2737 1 2 541 2 341 1 sky130_fd_sc_hd__clkbuf_16 $T=690000 155040 0 0 $X=689810 $Y=154800
X2738 1 2 547 2 360 1 sky130_fd_sc_hd__clkbuf_16 $T=727720 160480 1 0 $X=727530 $Y=157520
X2739 1 2 641 29 680 680 654 38 ICV_59 $T=47840 144160 1 0 $X=47650 $Y=141200
X2740 1 2 745 5 763 757 760 40 ICV_59 $T=89700 155040 0 0 $X=89510 $Y=154800
X2741 1 2 729 26 793 792 752 20 ICV_59 $T=103960 176800 1 0 $X=103770 $Y=173840
X2742 1 2 782 27 819 819 798 37 ICV_59 $T=117760 155040 0 0 $X=117570 $Y=154800
X2743 1 2 837 8 846 846 851 21 ICV_59 $T=132020 144160 1 0 $X=131830 $Y=141200
X2744 1 2 125 29 959 955 128 32 ICV_59 $T=188140 171360 1 0 $X=187950 $Y=168400
X2745 1 2 941 5 986 986 969 20 ICV_59 $T=201940 138720 0 0 $X=201750 $Y=138480
X2746 1 2 941 28 987 987 969 40 ICV_59 $T=201940 144160 0 0 $X=201750 $Y=143920
X2747 1 2 125 28 988 988 128 40 ICV_59 $T=201940 171360 0 0 $X=201750 $Y=171120
X2748 1 2 125 9 990 990 128 11 ICV_59 $T=201940 176800 0 0 $X=201750 $Y=176560
X2749 1 2 1000 154 1013 1005 1004 166 ICV_59 $T=216200 133280 1 0 $X=216010 $Y=130320
X2750 1 2 1000 156 1011 1009 1014 166 ICV_59 $T=216200 138720 1 0 $X=216010 $Y=135760
X2751 1 2 1002 154 1016 1016 997 167 ICV_59 $T=216200 149600 1 0 $X=216010 $Y=146640
X2752 1 2 151 156 1018 1018 163 162 ICV_59 $T=216200 176800 1 0 $X=216010 $Y=173840
X2753 1 2 1000 179 1029 1029 1014 188 ICV_59 $T=230000 133280 0 0 $X=229810 $Y=133040
X2754 1 2 1001 175 1033 1033 995 185 ICV_59 $T=230000 171360 0 0 $X=229810 $Y=171120
X2755 1 2 1108 196 1137 1137 1117 207 ICV_59 $T=286120 149600 0 0 $X=285930 $Y=149360
X2756 1 2 1153 154 1168 1168 1163 167 ICV_59 $T=300380 155040 1 0 $X=300190 $Y=152080
X2757 1 2 230 155 1194 1190 231 166 ICV_59 $T=314180 176800 0 0 $X=313990 $Y=176560
X2758 1 2 1349 178 1380 1380 1360 189 ICV_59 $T=412620 155040 1 0 $X=412430 $Y=152080
X2759 1 2 1395 197 1402 1402 1400 203 ICV_59 $T=426420 133280 0 0 $X=426230 $Y=133040
X2760 1 2 392 395 1550 402 393 405 ICV_59 $T=510600 176800 0 0 $X=510410 $Y=176560
X2761 1 2 392 388 1584 1584 393 396 ICV_59 $T=524860 176800 1 0 $X=524670 $Y=173840
X2762 1 2 452 295 1648 1650 1639 320 ICV_59 $T=566720 116960 0 0 $X=566530 $Y=116720
X2763 1 2 1688 310 1711 1714 1679 325 ICV_59 $T=609040 149600 1 0 $X=608850 $Y=146640
X2764 1 2 1749 281 1766 1772 1763 309 ICV_59 $T=637100 133280 1 0 $X=636910 $Y=130320
X2765 1 2 1749 310 1791 1792 1763 304 ICV_59 $T=650900 127840 0 0 $X=650710 $Y=127600
X2766 1 2 529 360 1813 1815 531 371 ICV_59 $T=665160 122400 1 0 $X=664970 $Y=119440
X2767 1 2 1806 338 1823 1823 1824 345 ICV_59 $T=665160 133280 1 0 $X=664970 $Y=130320
X2768 1 2 1795 400 1814 1812 1804 396 ICV_59 $T=665160 165920 1 0 $X=664970 $Y=162960
X2769 1 2 1844 338 1876 1876 1866 345 ICV_59 $T=693220 133280 1 0 $X=693030 $Y=130320
X2770 1 2 1859 339 1877 1872 1868 356 ICV_59 $T=693220 138720 1 0 $X=693030 $Y=135760
X2771 1 2 1859 340 1906 1900 1868 365 ICV_59 $T=707020 133280 0 0 $X=706830 $Y=133040
X2772 1 2 664 29 673 678 683 19 ICV_60 $T=46920 171360 0 0 $X=46730 $Y=171120
X2773 1 2 641 6 677 677 654 19 ICV_60 $T=47380 138720 0 0 $X=47190 $Y=138480
X2774 1 2 73 9 767 773 754 37 ICV_60 $T=93840 127840 0 0 $X=93650 $Y=127600
X2775 1 2 941 27 964 963 969 21 ICV_60 $T=188600 144160 1 0 $X=188410 $Y=141200
X2776 1 2 1000 155 1007 1011 1014 162 ICV_60 $T=215280 138720 0 0 $X=215090 $Y=138480
X2777 1 2 1000 153 1009 1013 1014 167 ICV_60 $T=215740 133280 0 0 $X=215550 $Y=133040
X2778 1 2 1001 156 1010 1010 995 162 ICV_60 $T=215740 160480 0 0 $X=215550 $Y=160240
X2779 1 2 1044 194 1053 1026 997 189 ICV_60 $T=243800 144160 0 0 $X=243610 $Y=143920
X2780 1 2 1044 206 1078 1078 1042 216 ICV_60 $T=258060 144160 1 0 $X=257870 $Y=141200
X2781 1 2 1075 197 1086 1086 1094 203 ICV_60 $T=264040 122400 0 0 $X=263850 $Y=122160
X2782 1 2 1124 156 1136 1136 1118 162 ICV_60 $T=286120 176800 1 0 $X=285930 $Y=173840
X2783 1 2 1156 178 1193 1197 1161 162 ICV_60 $T=314180 165920 1 0 $X=313990 $Y=162960
X2784 1 2 1248 175 1289 1289 1261 185 ICV_60 $T=361100 138720 1 0 $X=360910 $Y=135760
X2785 1 2 1350 179 1378 1381 1367 186 ICV_60 $T=412160 160480 0 0 $X=411970 $Y=160240
X2786 1 2 1354 176 1388 1388 1372 186 ICV_60 $T=415380 138720 1 0 $X=415190 $Y=135760
X2787 1 2 314 283 1446 324 319 305 ICV_60 $T=448040 176800 1 0 $X=447850 $Y=173840
X2788 1 2 1476 343 1506 1506 1501 354 ICV_60 $T=482540 122400 1 0 $X=482350 $Y=119440
X2789 1 2 1548 295 1554 1561 1555 294 ICV_60 $T=510140 127840 1 0 $X=509950 $Y=124880
X2790 1 2 1547 295 1551 1562 1538 316 ICV_60 $T=510600 155040 1 0 $X=510410 $Y=152080
X2791 1 2 424 357 449 1629 433 371 ICV_60 $T=552460 116960 0 0 $X=552270 $Y=116720
X2792 1 2 1704 296 1737 1737 1719 304 ICV_60 $T=622840 127840 1 0 $X=622650 $Y=124880
X2793 1 2 1688 307 1738 1741 1707 305 ICV_60 $T=622840 160480 1 0 $X=622650 $Y=157520
X2794 1 2 1733 295 1751 1751 1756 320 ICV_60 $T=628820 133280 0 0 $X=628630 $Y=133040
X2795 1 2 1795 378 1810 1810 1804 391 ICV_60 $T=660100 165920 0 0 $X=659910 $Y=165680
X2796 1 2 1779 339 1817 1817 1794 344 ICV_60 $T=664240 138720 0 0 $X=664050 $Y=138480
X2797 1 2 1806 339 1820 1820 1824 344 ICV_60 $T=664700 133280 0 0 $X=664510 $Y=133040
X2798 1 2 1779 343 1821 1821 1794 354 ICV_60 $T=664700 144160 0 0 $X=664510 $Y=143920
X2799 1 2 1835 382 1840 1851 539 407 ICV_60 $T=678960 176800 1 0 $X=678770 $Y=173840
X2800 1 2 1806 357 1848 1847 1824 351 ICV_60 $T=679420 133280 0 0 $X=679230 $Y=133040
X2801 1 2 1859 341 1867 1875 1868 371 ICV_60 $T=692300 138720 0 0 $X=692110 $Y=138480
X2802 1 2 1844 357 1874 1874 1866 356 ICV_60 $T=692760 127840 0 0 $X=692570 $Y=127600
X2803 1 2 1869 339 1881 1856 1837 342 ICV_60 $T=697360 149600 1 0 $X=697170 $Y=146640
X2804 1 2 1871 380 1888 1883 1891 407 ICV_60 $T=699660 176800 1 0 $X=699470 $Y=173840
X2805 1 2 1919 382 1936 1941 1928 405 ICV_60 $T=720820 171360 0 0 $X=720630 $Y=171120
X2806 1 2 632 615 32 ICV_62 $T=39100 176800 1 0 $X=38910 $Y=173840
X2807 1 2 646 649 32 ICV_62 $T=42320 171360 0 0 $X=42130 $Y=171120
X2808 1 2 696 695 38 ICV_62 $T=64860 116960 1 0 $X=64670 $Y=114000
X2809 1 2 867 103 20 ICV_62 $T=147660 116960 0 0 $X=147470 $Y=116720
X2810 1 2 930 892 20 ICV_62 $T=180780 160480 0 0 $X=180590 $Y=160240
X2811 1 2 1051 1047 201 ICV_62 $T=256220 133280 1 0 $X=256030 $Y=130320
X2812 1 2 1132 1094 210 ICV_62 $T=291640 122400 1 0 $X=291450 $Y=119440
X2813 1 2 1155 227 162 ICV_62 $T=305440 116960 0 0 $X=305250 $Y=116720
X2814 1 2 1238 1205 214 ICV_62 $T=343160 122400 0 0 $X=342970 $Y=122160
X2815 1 2 1359 1360 150 ICV_62 $T=425500 149600 1 0 $X=425310 $Y=146640
X2816 1 2 1424 302 316 ICV_62 $T=445740 165920 0 0 $X=445550 $Y=165680
X2817 1 2 1459 1452 300 ICV_62 $T=464140 122400 1 0 $X=463950 $Y=119440
X2818 1 2 1531 1534 344 ICV_62 $T=505540 127840 1 0 $X=505350 $Y=124880
X2819 1 2 1565 386 407 ICV_62 $T=524860 171360 0 0 $X=524670 $Y=171120
X2820 1 2 1643 1639 316 ICV_62 $T=568100 127840 0 0 $X=567910 $Y=127600
X2821 1 2 1711 1707 325 ICV_62 $T=618240 149600 0 0 $X=618050 $Y=149360
X2822 1 2 1730 1707 300 ICV_62 $T=622380 149600 1 0 $X=622190 $Y=146640
X2823 1 2 1784 1743 325 ICV_62 $T=660560 149600 0 0 $X=660370 $Y=149360
X2824 1 2 1788 517 325 ICV_62 $T=677120 122400 1 0 $X=676930 $Y=119440
X2825 1 2 652 649 37 ICV_63 $T=42780 160480 1 0 $X=42590 $Y=157520
X2826 1 2 749 752 11 ICV_63 $T=88780 176800 1 0 $X=88590 $Y=173840
X2827 1 2 753 754 32 ICV_63 $T=90160 122400 0 0 $X=89970 $Y=122160
X2828 1 2 768 760 38 ICV_63 $T=98900 160480 1 0 $X=98710 $Y=157520
X2829 1 2 856 858 19 ICV_63 $T=139840 171360 1 0 $X=139650 $Y=168400
X2830 1 2 885 858 37 ICV_63 $T=156860 171360 0 0 $X=156670 $Y=171120
X2831 1 2 897 899 19 ICV_63 $T=160540 122400 1 0 $X=160350 $Y=119440
X2832 1 2 893 899 40 ICV_63 $T=160540 127840 1 0 $X=160350 $Y=124880
X2833 1 2 945 951 32 ICV_63 $T=188600 116960 1 0 $X=188410 $Y=114000
X2834 1 2 949 951 37 ICV_63 $T=188600 127840 1 0 $X=188410 $Y=124880
X2835 1 2 947 944 38 ICV_63 $T=188600 160480 1 0 $X=188410 $Y=157520
X2836 1 2 1230 1214 189 ICV_63 $T=337180 171360 0 0 $X=336990 $Y=171120
X2837 1 2 1331 1324 185 ICV_63 $T=391000 160480 0 0 $X=390810 $Y=160240
X2838 1 2 1393 293 186 ICV_63 $T=426880 122400 0 0 $X=426690 $Y=122160
X2839 1 2 1564 1555 309 ICV_63 $T=519340 122400 1 0 $X=519150 $Y=119440
X2840 1 2 1623 1604 351 ICV_63 $T=553380 127840 1 0 $X=553190 $Y=124880
X2841 1 2 1624 1604 371 ICV_63 $T=553380 133280 1 0 $X=553190 $Y=130320
X2842 1 2 1702 1707 320 ICV_63 $T=609500 155040 1 0 $X=609310 $Y=152080
X2843 1 2 1800 1794 365 ICV_63 $T=659640 133280 0 0 $X=659450 $Y=133040
X2844 1 2 1887 1892 351 ICV_63 $T=707480 149600 0 0 $X=707290 $Y=149360
X2845 1 2 745 29 768 ICV_66 $T=96600 155040 1 0 $X=96410 $Y=152080
X2846 1 2 876 9 891 ICV_66 $T=152720 155040 1 0 $X=152530 $Y=152080
X2847 1 2 1077 206 1090 ICV_66 $T=264960 138720 1 0 $X=264770 $Y=135760
X2848 1 2 1076 206 1093 ICV_66 $T=264960 160480 1 0 $X=264770 $Y=157520
X2849 1 2 1192 175 1210 ICV_66 $T=321080 138720 1 0 $X=320890 $Y=135760
X2850 1 2 1208 175 1236 ICV_66 $T=334880 149600 0 0 $X=334690 $Y=149360
X2851 1 2 1208 178 1237 ICV_66 $T=334880 155040 0 0 $X=334690 $Y=154800
X2852 1 2 1253 153 1266 ICV_66 $T=349140 155040 1 0 $X=348950 $Y=152080
X2853 1 2 1303 179 1344 ICV_66 $T=391000 133280 0 0 $X=390810 $Y=133040
X2854 1 2 1354 154 1371 ICV_66 $T=405260 138720 1 0 $X=405070 $Y=135760
X2855 1 2 279 281 1394 ICV_66 $T=419060 176800 0 0 $X=418870 $Y=176560
X2856 1 2 1377 178 1415 ICV_66 $T=433320 116960 1 0 $X=433130 $Y=114000
X2857 1 2 160 356 1522 ICV_66 $T=489440 160480 1 0 $X=489250 $Y=157520
X2858 1 2 1795 380 1807 ICV_66 $T=657800 171360 1 0 $X=657610 $Y=168400
X2859 1 2 1818 360 1832 ICV_66 $T=671600 149600 0 0 $X=671410 $Y=149360
X2860 1 2 1904 358 1922 ICV_66 $T=713920 122400 1 0 $X=713730 $Y=119440
X2861 1 2 544 395 1923 ICV_66 $T=713920 176800 1 0 $X=713730 $Y=173840
X2862 1 2 544 400 1947 ICV_66 $T=727720 176800 0 0 $X=727530 $Y=176560
X2863 1 2 88 14 138 141 2 132 1 sky130_fd_sc_hd__and4b_2 $T=199640 116960 1 0 $X=199450 $Y=114000
X2864 1 2 1553 1556 1552 1560 2 336 1 sky130_fd_sc_hd__and4b_2 $T=515200 138720 0 0 $X=515010 $Y=138480
X2865 1 2 1552 1556 1553 1557 2 404 1 sky130_fd_sc_hd__and4b_2 $T=518420 144160 0 0 $X=518230 $Y=143920
X2866 1 2 1553 1556 1552 1557 2 330 1 sky130_fd_sc_hd__and4b_2 $T=520720 149600 1 0 $X=520530 $Y=146640
X2867 1 2 1556 1553 1552 1557 2 410 1 sky130_fd_sc_hd__and4b_2 $T=522560 144160 0 0 $X=522370 $Y=143920
X2868 1 2 88 14 138 1572 2 1570 1 sky130_fd_sc_hd__and4b_2 $T=525320 133280 1 0 $X=525130 $Y=130320
X2869 1 2 138 88 14 1572 2 1589 1 sky130_fd_sc_hd__and4b_2 $T=533600 138720 0 0 $X=533410 $Y=138480
X2870 1 2 14 88 138 1572 2 1599 1 sky130_fd_sc_hd__and4b_2 $T=534980 149600 1 0 $X=534790 $Y=146640
X2871 1 2 1553 1556 1552 1586 2 427 1 sky130_fd_sc_hd__and4b_2 $T=539580 133280 0 0 $X=539390 $Y=133040
X2872 1 2 1556 1553 1552 1586 2 431 1 sky130_fd_sc_hd__and4b_2 $T=542800 133280 1 0 $X=542610 $Y=130320
X2873 1 2 1556 1553 1552 1579 2 432 1 sky130_fd_sc_hd__and4b_2 $T=544640 144160 0 0 $X=544450 $Y=143920
X2874 1 2 1552 1556 1553 1586 2 437 1 sky130_fd_sc_hd__and4b_2 $T=548320 133280 0 0 $X=548130 $Y=133040
X2875 1 2 1552 1556 1553 1560 2 384 1 sky130_fd_sc_hd__and4b_2 $T=548780 138720 1 0 $X=548590 $Y=135760
X2876 1 2 1553 1556 1552 1579 2 352 1 sky130_fd_sc_hd__and4b_2 $T=553380 144160 1 0 $X=553190 $Y=141200
X2877 1 2 1556 1553 1552 1560 2 447 1 sky130_fd_sc_hd__and4b_2 $T=554760 138720 0 0 $X=554570 $Y=138480
X2878 1 2 1552 1556 1553 1579 2 464 1 sky130_fd_sc_hd__and4b_2 $T=570860 138720 0 0 $X=570670 $Y=138480
X2879 1 2 1553 1556 1552 1570 2 474 1 sky130_fd_sc_hd__and4b_2 $T=579600 133280 0 0 $X=579410 $Y=133040
X2880 1 2 1556 1553 1552 1589 2 472 1 sky130_fd_sc_hd__and4b_2 $T=582360 138720 0 0 $X=582170 $Y=138480
X2881 1 2 1552 1556 1553 1589 2 461 1 sky130_fd_sc_hd__and4b_2 $T=588800 138720 1 0 $X=588610 $Y=135760
X2882 1 2 1553 1556 1552 1589 2 490 1 sky130_fd_sc_hd__and4b_2 $T=602140 138720 1 0 $X=601950 $Y=135760
X2883 1 2 1556 1553 1552 1570 2 495 1 sky130_fd_sc_hd__and4b_2 $T=604440 133280 0 0 $X=604250 $Y=133040
X2884 1 2 1552 1556 1553 1570 2 504 1 sky130_fd_sc_hd__and4b_2 $T=614100 133280 0 0 $X=613910 $Y=133040
X2885 1 2 1552 1556 1553 1592 2 489 1 sky130_fd_sc_hd__and4b_2 $T=617320 138720 0 0 $X=617130 $Y=138480
X2886 1 2 1553 1556 1552 1599 2 509 1 sky130_fd_sc_hd__and4b_2 $T=618700 144160 0 0 $X=618510 $Y=143920
X2887 1 2 1553 1556 1552 1592 2 511 1 sky130_fd_sc_hd__and4b_2 $T=621460 133280 1 0 $X=621270 $Y=130320
X2888 1 2 1552 1556 1553 1599 2 514 1 sky130_fd_sc_hd__and4b_2 $T=622840 144160 1 0 $X=622650 $Y=141200
X2889 1 2 1556 1553 1552 1592 2 513 1 sky130_fd_sc_hd__and4b_2 $T=623300 133280 0 0 $X=623110 $Y=133040
X2890 1 2 1556 1553 1552 1599 2 508 1 sky130_fd_sc_hd__and4b_2 $T=623300 144160 0 0 $X=623110 $Y=143920
X2891 1 2 1553 1556 1552 1557 2 406 1 sky130_fd_sc_hd__and4_2 $T=520260 133280 1 0 $X=520070 $Y=130320
X2892 1 2 14 88 138 1572 2 1592 1 sky130_fd_sc_hd__and4_2 $T=534980 133280 0 0 $X=534790 $Y=133040
X2893 1 2 1553 1556 1552 1586 2 438 1 sky130_fd_sc_hd__and4_2 $T=549240 149600 1 0 $X=549050 $Y=146640
X2894 1 2 1553 1556 1552 1579 2 457 1 sky130_fd_sc_hd__and4_2 $T=565800 149600 1 0 $X=565610 $Y=146640
X2895 1 2 1553 1556 1552 1560 2 460 1 sky130_fd_sc_hd__and4_2 $T=567180 138720 0 0 $X=566990 $Y=138480
X2896 1 2 1553 1556 1552 1589 2 468 1 sky130_fd_sc_hd__and4_2 $T=593400 133280 1 0 $X=593210 $Y=130320
X2897 1 2 1553 1556 1552 1570 2 507 1 sky130_fd_sc_hd__and4_2 $T=618240 133280 0 0 $X=618050 $Y=133040
X2898 1 2 1553 1556 1552 1592 2 516 1 sky130_fd_sc_hd__and4_2 $T=627440 127840 0 0 $X=627250 $Y=127600
X2899 1 2 1553 1556 1552 1599 2 521 1 sky130_fd_sc_hd__and4_2 $T=633420 149600 1 0 $X=633230 $Y=146640
X2900 1 2 954 956 2 32 1 sky130_fd_sc_hd__ebufn_4 $T=189980 149600 0 0 $X=189790 $Y=149360
X2901 1 2 954 956 2 37 1 sky130_fd_sc_hd__ebufn_4 $T=192740 155040 1 0 $X=192550 $Y=152080
X2902 1 2 954 956 2 38 1 sky130_fd_sc_hd__ebufn_4 $T=192740 155040 0 0 $X=192550 $Y=154800
X2903 1 2 954 956 2 21 1 sky130_fd_sc_hd__ebufn_4 $T=195960 149600 0 0 $X=195770 $Y=149360
X2904 1 2 954 956 2 19 1 sky130_fd_sc_hd__ebufn_4 $T=203780 149600 0 0 $X=203590 $Y=149360
X2905 1 2 954 956 2 40 1 sky130_fd_sc_hd__ebufn_4 $T=203780 155040 1 0 $X=203590 $Y=152080
X2906 1 2 954 956 2 20 1 sky130_fd_sc_hd__ebufn_4 $T=203780 155040 0 0 $X=203590 $Y=154800
X2907 1 2 954 956 2 152 1 sky130_fd_sc_hd__ebufn_4 $T=209760 160480 0 0 $X=209570 $Y=160240
X2908 1 2 954 956 2 95 1 sky130_fd_sc_hd__ebufn_4 $T=210220 155040 0 0 $X=210030 $Y=154800
X2909 1 2 954 956 2 11 1 sky130_fd_sc_hd__ebufn_4 $T=210220 160480 1 0 $X=210030 $Y=157520
X2910 1 2 954 956 2 71 1 sky130_fd_sc_hd__ebufn_4 $T=216200 155040 0 0 $X=216010 $Y=154800
X2911 1 2 954 956 2 47 1 sky130_fd_sc_hd__ebufn_4 $T=216660 155040 1 0 $X=216470 $Y=152080
X2912 1 2 954 956 2 167 1 sky130_fd_sc_hd__ebufn_4 $T=222640 155040 1 0 $X=222450 $Y=152080
X2913 1 2 954 956 2 174 1 sky130_fd_sc_hd__ebufn_4 $T=224020 155040 0 0 $X=223830 $Y=154800
X2914 1 2 954 956 2 161 1 sky130_fd_sc_hd__ebufn_4 $T=224020 160480 1 0 $X=223830 $Y=157520
X2915 1 2 954 956 2 182 1 sky130_fd_sc_hd__ebufn_4 $T=230460 155040 0 0 $X=230270 $Y=154800
X2916 1 2 954 956 2 162 1 sky130_fd_sc_hd__ebufn_4 $T=232300 160480 1 0 $X=232110 $Y=157520
X2917 1 2 954 956 2 150 1 sky130_fd_sc_hd__ebufn_4 $T=233680 160480 0 0 $X=233490 $Y=160240
X2918 1 2 954 956 2 186 1 sky130_fd_sc_hd__ebufn_4 $T=236440 155040 0 0 $X=236250 $Y=154800
X2919 1 2 954 956 2 189 1 sky130_fd_sc_hd__ebufn_4 $T=237820 155040 1 0 $X=237630 $Y=152080
X2920 1 2 954 956 2 166 1 sky130_fd_sc_hd__ebufn_4 $T=238280 160480 1 0 $X=238090 $Y=157520
X2921 1 2 954 956 2 201 1 sky130_fd_sc_hd__ebufn_4 $T=244260 149600 0 0 $X=244070 $Y=149360
X2922 1 2 954 956 2 188 1 sky130_fd_sc_hd__ebufn_4 $T=244720 155040 1 0 $X=244530 $Y=152080
X2923 1 2 954 956 2 203 1 sky130_fd_sc_hd__ebufn_4 $T=246100 160480 1 0 $X=245910 $Y=157520
X2924 1 2 954 956 2 202 1 sky130_fd_sc_hd__ebufn_4 $T=246560 155040 0 0 $X=246370 $Y=154800
X2925 1 2 954 956 2 207 1 sky130_fd_sc_hd__ebufn_4 $T=249780 160480 0 0 $X=249590 $Y=160240
X2926 1 2 954 956 2 210 1 sky130_fd_sc_hd__ebufn_4 $T=250700 149600 0 0 $X=250510 $Y=149360
X2927 1 2 954 956 2 214 1 sky130_fd_sc_hd__ebufn_4 $T=252540 160480 1 0 $X=252350 $Y=157520
X2928 1 2 954 956 2 200 1 sky130_fd_sc_hd__ebufn_4 $T=255760 155040 1 0 $X=255570 $Y=152080
X2929 1 2 954 956 2 216 1 sky130_fd_sc_hd__ebufn_4 $T=258520 149600 0 0 $X=258330 $Y=149360
X2930 1 2 954 956 2 185 1 sky130_fd_sc_hd__ebufn_4 $T=258520 155040 0 0 $X=258330 $Y=154800
X2931 1 2 954 956 2 211 1 sky130_fd_sc_hd__ebufn_4 $T=258520 160480 0 0 $X=258330 $Y=160240
X2932 1 2 459 456 2 316 1 sky130_fd_sc_hd__ebufn_4 $T=569020 155040 1 0 $X=568830 $Y=152080
X2933 1 2 459 456 2 351 1 sky130_fd_sc_hd__ebufn_4 $T=569480 149600 1 0 $X=569290 $Y=146640
X2934 1 2 459 456 2 356 1 sky130_fd_sc_hd__ebufn_4 $T=569480 149600 0 0 $X=569290 $Y=149360
X2935 1 2 459 456 2 305 1 sky130_fd_sc_hd__ebufn_4 $T=571780 155040 0 0 $X=571590 $Y=154800
X2936 1 2 459 456 2 304 1 sky130_fd_sc_hd__ebufn_4 $T=571780 160480 1 0 $X=571590 $Y=157520
X2937 1 2 459 456 2 465 1 sky130_fd_sc_hd__ebufn_4 $T=572240 176800 1 0 $X=572050 $Y=173840
X2938 1 2 459 456 2 396 1 sky130_fd_sc_hd__ebufn_4 $T=574540 160480 0 0 $X=574350 $Y=160240
X2939 1 2 459 456 2 300 1 sky130_fd_sc_hd__ebufn_4 $T=575000 155040 1 0 $X=574810 $Y=152080
X2940 1 2 459 456 2 405 1 sky130_fd_sc_hd__ebufn_4 $T=576380 176800 0 0 $X=576190 $Y=176560
X2941 1 2 459 456 2 342 1 sky130_fd_sc_hd__ebufn_4 $T=576840 144160 0 0 $X=576650 $Y=143920
X2942 1 2 459 456 2 345 1 sky130_fd_sc_hd__ebufn_4 $T=576840 149600 0 0 $X=576650 $Y=149360
X2943 1 2 459 456 2 320 1 sky130_fd_sc_hd__ebufn_4 $T=579600 155040 0 0 $X=579410 $Y=154800
X2944 1 2 459 456 2 397 1 sky130_fd_sc_hd__ebufn_4 $T=580520 160480 0 0 $X=580330 $Y=160240
X2945 1 2 459 456 2 344 1 sky130_fd_sc_hd__ebufn_4 $T=581440 149600 1 0 $X=581250 $Y=146640
X2946 1 2 459 456 2 371 1 sky130_fd_sc_hd__ebufn_4 $T=581440 155040 1 0 $X=581250 $Y=152080
X2947 1 2 459 456 2 444 1 sky130_fd_sc_hd__ebufn_4 $T=582360 171360 1 0 $X=582170 $Y=168400
X2948 1 2 459 456 2 354 1 sky130_fd_sc_hd__ebufn_4 $T=582820 149600 0 0 $X=582630 $Y=149360
X2949 1 2 459 456 2 423 1 sky130_fd_sc_hd__ebufn_4 $T=582820 165920 1 0 $X=582630 $Y=162960
X2950 1 2 459 456 2 407 1 sky130_fd_sc_hd__ebufn_4 $T=582820 176800 1 0 $X=582630 $Y=173840
X2951 1 2 459 456 2 409 1 sky130_fd_sc_hd__ebufn_4 $T=584200 171360 0 0 $X=584010 $Y=171120
X2952 1 2 459 456 2 391 1 sky130_fd_sc_hd__ebufn_4 $T=584660 165920 0 0 $X=584470 $Y=165680
X2953 1 2 459 456 2 294 1 sky130_fd_sc_hd__ebufn_4 $T=586040 155040 0 0 $X=585850 $Y=154800
X2954 1 2 459 456 2 309 1 sky130_fd_sc_hd__ebufn_4 $T=586500 160480 1 0 $X=586310 $Y=157520
X2955 1 2 459 456 2 365 1 sky130_fd_sc_hd__ebufn_4 $T=587420 155040 1 0 $X=587230 $Y=152080
X2956 1 2 459 456 2 325 1 sky130_fd_sc_hd__ebufn_4 $T=588800 149600 0 0 $X=588610 $Y=149360
X2957 1 2 1553 1556 1552 1557 2 308 1 sky130_fd_sc_hd__nor4b_2 $T=519340 138720 0 0 $X=519150 $Y=138480
X2958 1 2 1553 1556 1552 1570 2 408 1 sky130_fd_sc_hd__nor4b_2 $T=521180 133280 0 0 $X=520990 $Y=133040
X2959 1 2 1553 1556 1552 1560 2 312 1 sky130_fd_sc_hd__nor4b_2 $T=525320 138720 1 0 $X=525130 $Y=135760
X2960 1 2 14 88 138 1572 2 1557 1 sky130_fd_sc_hd__nor4b_2 $T=525320 144160 1 0 $X=525130 $Y=141200
X2961 1 2 1553 1556 1552 1586 2 337 1 sky130_fd_sc_hd__nor4b_2 $T=529460 133280 0 0 $X=529270 $Y=133040
X2962 1 2 1553 1556 1552 1589 2 419 1 sky130_fd_sc_hd__nor4b_2 $T=531300 138720 1 0 $X=531110 $Y=135760
X2963 1 2 1553 1556 1552 1592 2 289 1 sky130_fd_sc_hd__nor4b_2 $T=539120 138720 0 0 $X=538930 $Y=138480
X2964 1 2 1553 1556 1552 1599 2 350 1 sky130_fd_sc_hd__nor4b_2 $T=539120 144160 0 0 $X=538930 $Y=143920
X2965 1 2 1553 1556 1552 1579 2 430 1 sky130_fd_sc_hd__nor4b_2 $T=541420 144160 1 0 $X=541230 $Y=141200
X2966 1 2 130 131 132 133 2 78 1 sky130_fd_sc_hd__and4bb_2 $T=193660 116960 1 0 $X=193470 $Y=114000
X2967 1 2 1552 1553 1557 1556 2 398 1 sky130_fd_sc_hd__and4bb_2 $T=513360 144160 1 0 $X=513170 $Y=141200
X2968 1 2 1553 1552 1557 1556 2 366 1 sky130_fd_sc_hd__and4bb_2 $T=513820 144160 0 0 $X=513630 $Y=143920
X2969 1 2 1552 1556 1560 1553 2 306 1 sky130_fd_sc_hd__and4bb_2 $T=515200 138720 1 0 $X=515010 $Y=135760
X2970 1 2 1552 1556 1557 1553 2 401 1 sky130_fd_sc_hd__and4bb_2 $T=517960 144160 1 0 $X=517770 $Y=141200
X2971 1 2 1553 1552 1560 1556 2 322 1 sky130_fd_sc_hd__and4bb_2 $T=519800 138720 1 0 $X=519610 $Y=135760
X2972 1 2 138 88 1572 14 2 1560 1 sky130_fd_sc_hd__and4bb_2 $T=525780 138720 0 0 $X=525590 $Y=138480
X2973 1 2 1552 1556 1579 1553 2 333 1 sky130_fd_sc_hd__and4bb_2 $T=527160 144160 0 0 $X=526970 $Y=143920
X2974 1 2 1552 1556 1586 1553 2 413 1 sky130_fd_sc_hd__and4bb_2 $T=530380 133280 1 0 $X=530190 $Y=130320
X2975 1 2 138 14 1572 88 2 1579 1 sky130_fd_sc_hd__and4bb_2 $T=531300 144160 1 0 $X=531110 $Y=141200
X2976 1 2 1553 1552 1579 1556 2 416 1 sky130_fd_sc_hd__and4bb_2 $T=531760 144160 0 0 $X=531570 $Y=143920
X2977 1 2 14 138 1572 88 2 1586 1 sky130_fd_sc_hd__and4bb_2 $T=536820 138720 1 0 $X=536630 $Y=135760
X2978 1 2 1553 1552 1586 1556 2 426 1 sky130_fd_sc_hd__and4bb_2 $T=541420 138720 1 0 $X=541230 $Y=135760
X2979 1 2 1552 1553 1586 1556 2 429 1 sky130_fd_sc_hd__and4bb_2 $T=543720 133280 0 0 $X=543530 $Y=133040
X2980 1 2 1552 1553 1579 1556 2 421 1 sky130_fd_sc_hd__and4bb_2 $T=547400 144160 1 0 $X=547210 $Y=141200
X2981 1 2 1552 1553 1560 1556 2 434 1 sky130_fd_sc_hd__and4bb_2 $T=550160 138720 0 0 $X=549970 $Y=138480
X2982 1 2 1552 1556 1589 1553 2 453 1 sky130_fd_sc_hd__and4bb_2 $T=562120 138720 0 0 $X=561930 $Y=138480
X2983 1 2 1553 1552 1599 1556 2 470 1 sky130_fd_sc_hd__and4bb_2 $T=581440 144160 1 0 $X=581250 $Y=141200
X2984 1 2 1552 1553 1570 1556 2 476 1 sky130_fd_sc_hd__and4bb_2 $T=583740 138720 1 0 $X=583550 $Y=135760
X2985 1 2 1553 1552 1589 1556 2 482 1 sky130_fd_sc_hd__and4bb_2 $T=592940 138720 1 0 $X=592750 $Y=135760
X2986 1 2 1552 1553 1589 1556 2 487 1 sky130_fd_sc_hd__and4bb_2 $T=597540 138720 1 0 $X=597350 $Y=135760
X2987 1 2 1552 1556 1599 1553 2 479 1 sky130_fd_sc_hd__and4bb_2 $T=599840 138720 0 0 $X=599650 $Y=138480
X2988 1 2 1552 1556 1570 1553 2 496 1 sky130_fd_sc_hd__and4bb_2 $T=608580 133280 0 0 $X=608390 $Y=133040
X2989 1 2 1553 1552 1570 1556 2 499 1 sky130_fd_sc_hd__and4bb_2 $T=609500 138720 1 0 $X=609310 $Y=135760
X2990 1 2 1552 1556 1592 1553 2 501 1 sky130_fd_sc_hd__and4bb_2 $T=611340 138720 0 0 $X=611150 $Y=138480
X2991 1 2 1552 1553 1592 1556 2 502 1 sky130_fd_sc_hd__and4bb_2 $T=615480 138720 1 0 $X=615290 $Y=135760
X2992 1 2 1552 1553 1599 1556 2 505 1 sky130_fd_sc_hd__and4bb_2 $T=618240 144160 1 0 $X=618050 $Y=141200
X2993 1 2 1553 1552 1592 1556 2 510 1 sky130_fd_sc_hd__and4bb_2 $T=623300 138720 0 0 $X=623110 $Y=138480
X2994 1 2 141 2 956 1 sky130_fd_sc_hd__clkbuf_4 $T=209760 149600 0 0 $X=209570 $Y=149360
X2995 1 2 1572 2 456 1 sky130_fd_sc_hd__clkbuf_4 $T=565340 155040 1 0 $X=565150 $Y=152080
X2996 2 1 954 sky130_fd_sc_hd__conb_1 $T=191360 155040 0 0 $X=191170 $Y=154800
X2997 2 1 459 sky130_fd_sc_hd__conb_1 $T=575460 149600 0 0 $X=575270 $Y=149360
X2998 1 2 729 6 769 ICV_72 $T=93840 171360 1 0 $X=93650 $Y=168400
X2999 1 2 1040 179 1050 ICV_72 $T=241960 171360 0 0 $X=241770 $Y=171120
X3000 1 2 199 156 1085 ICV_72 $T=262660 176800 0 0 $X=262470 $Y=176560
X3001 1 2 1075 206 1087 ICV_72 $T=264500 122400 1 0 $X=264310 $Y=119440
X3002 1 2 1192 179 1229 ICV_72 $T=333040 133280 1 0 $X=332850 $Y=130320
X3003 1 2 255 175 1313 ICV_72 $T=373520 171360 0 0 $X=373330 $Y=171120
X3004 1 2 255 179 1314 ICV_72 $T=373520 176800 0 0 $X=373330 $Y=176560
X3005 1 2 1312 178 1335 ICV_72 $T=387780 122400 0 0 $X=387590 $Y=122160
X3006 1 2 1377 179 1399 ICV_72 $T=422280 122400 1 0 $X=422090 $Y=119440
X3007 1 2 1440 310 1451 ICV_72 $T=454020 144160 1 0 $X=453830 $Y=141200
X3008 1 2 160 201 334 ICV_72 $T=460920 155040 1 0 $X=460730 $Y=152080
X3009 1 2 1476 340 1526 ICV_72 $T=496340 122400 0 0 $X=496150 $Y=122160
X3010 1 2 1588 339 1605 ICV_72 $T=534980 133280 1 0 $X=534790 $Y=130320
X3011 1 2 477 295 494 ICV_72 $T=598460 116960 1 0 $X=598270 $Y=114000
X3012 1 2 477 281 1726 ICV_72 $T=615020 116960 0 0 $X=614830 $Y=116720
X3013 1 2 1904 343 1925 ICV_72 $T=715300 122400 0 0 $X=715110 $Y=122160
X3014 1 2 17 18 614 614 584 111 ICV_74 $T=17480 138720 0 0 $X=17290 $Y=138480
X3015 1 2 33 18 631 631 586 111 ICV_74 $T=29440 138720 1 0 $X=29250 $Y=135760
X3016 1 2 60 18 714 714 702 111 ICV_74 $T=69460 116960 0 0 $X=69270 $Y=116720
X3017 1 2 75 18 762 762 745 111 ICV_74 $T=94760 149600 0 0 $X=94570 $Y=149360
X3018 1 2 87 18 810 810 816 111 ICV_74 $T=116840 116960 1 0 $X=116650 $Y=114000
X3019 1 2 99 18 841 841 100 111 ICV_74 $T=132940 116960 1 0 $X=132750 $Y=114000
X3020 1 2 102 18 868 868 837 111 ICV_74 $T=146280 138720 1 0 $X=146090 $Y=135760
X3021 1 2 22 146 984 984 1000 111 ICV_74 $T=207460 133280 1 0 $X=207270 $Y=130320
X3022 1 2 31 146 989 989 151 111 ICV_74 $T=207460 176800 1 0 $X=207270 $Y=173840
X3023 1 2 17 146 1039 1039 1040 111 ICV_74 $T=239200 165920 0 0 $X=239010 $Y=165680
X3024 1 2 31 191 1046 1046 1041 111 ICV_74 $T=242420 122400 0 0 $X=242230 $Y=122160
X3025 1 2 217 191 1082 1082 1077 111 ICV_74 $T=264500 127840 0 0 $X=264310 $Y=127600
X3026 1 2 120 146 1308 1308 1303 111 ICV_74 $T=377660 138720 0 0 $X=377470 $Y=138480
X3027 1 2 101 146 1321 1321 263 111 ICV_74 $T=381340 176800 0 0 $X=381150 $Y=176560
X3028 1 2 136 146 1374 1374 1377 111 ICV_74 $T=413540 122400 1 0 $X=413350 $Y=119440
X3029 1 2 337 332 1474 1474 347 481 ICV_74 $T=469200 116960 1 0 $X=469010 $Y=114000
X3030 1 2 366 370 1514 1514 1524 481 ICV_74 $T=491280 171360 0 0 $X=491090 $Y=171120
X3031 1 2 430 332 1618 1618 1626 481 ICV_74 $T=549240 144160 0 0 $X=549050 $Y=143920
X3032 1 2 461 290 1652 1652 1628 481 ICV_74 $T=572700 127840 0 0 $X=572510 $Y=127600
X3033 1 2 479 469 1670 1670 484 481 ICV_74 $T=588800 176800 1 0 $X=588610 $Y=173840
X3034 1 2 490 290 1694 1694 1704 481 ICV_74 $T=602600 127840 0 0 $X=602410 $Y=127600
X3035 1 2 513 290 1732 1732 1749 481 ICV_74 $T=625600 133280 1 0 $X=625410 $Y=130320
X3036 1 2 501 370 1744 1744 1755 481 ICV_74 $T=628820 160480 0 0 $X=628630 $Y=160240
X3037 1 2 429 370 1750 1750 522 481 ICV_74 $T=633420 176800 0 0 $X=633230 $Y=176560
X3038 1 2 406 370 1786 1786 1795 481 ICV_74 $T=651820 160480 0 0 $X=651630 $Y=160240
X3039 1 2 432 332 1797 1797 1806 481 ICV_74 $T=656420 133280 1 0 $X=656230 $Y=130320
X3040 1 2 508 332 1861 1861 1869 481 ICV_74 $T=690000 149600 0 0 $X=689810 $Y=149360
X3041 1 2 513 332 1907 1907 1916 481 ICV_74 $T=712540 144160 1 0 $X=712350 $Y=141200
X3042 1 2 1479 348 168 353 1498 173 2 359 1 sky130_fd_sc_hd__mux4_1 $T=477020 155040 1 0 $X=476830 $Y=152080
X3043 1 2 1434 355 168 362 1499 173 2 369 1 sky130_fd_sc_hd__mux4_1 $T=483000 155040 0 0 $X=482810 $Y=154800
X3044 1 2 1441 363 168 368 1512 173 2 373 1 sky130_fd_sc_hd__mux4_1 $T=487140 155040 1 0 $X=486950 $Y=152080
X3045 1 2 1435 367 168 372 1522 173 2 376 1 sky130_fd_sc_hd__mux4_1 $T=490820 149600 0 0 $X=490630 $Y=149360
X3046 1 2 1421 375 168 381 1527 173 2 387 1 sky130_fd_sc_hd__mux4_1 $T=498640 155040 0 0 $X=498450 $Y=154800
X3047 1 2 1407 377 168 383 1530 173 2 389 1 sky130_fd_sc_hd__mux4_1 $T=499560 160480 0 0 $X=499370 $Y=160240
X3048 1 2 1445 412 168 414 1585 173 2 422 1 sky130_fd_sc_hd__mux4_1 $T=527620 149600 0 0 $X=527430 $Y=149360
X3049 1 2 1417 417 168 420 1590 173 2 425 1 sky130_fd_sc_hd__mux4_1 $T=531760 160480 1 0 $X=531570 $Y=157520
X3050 1 2 843 29 859 ICV_80 $T=137080 165920 0 0 $X=136890 $Y=165680
X3051 1 2 928 5 979 ICV_80 $T=198720 133280 1 0 $X=198530 $Y=130320
X3052 1 2 199 153 1064 ICV_80 $T=247940 176800 0 0 $X=247750 $Y=176560
X3053 1 2 1077 197 1110 ICV_80 $T=273240 127840 0 0 $X=273050 $Y=127600
X3054 1 2 1075 193 1127 ICV_80 $T=281060 127840 1 0 $X=280870 $Y=124880
X3055 1 2 1108 193 1144 ICV_80 $T=289340 149600 1 0 $X=289150 $Y=146640
X3056 1 2 1395 204 1432 ICV_80 $T=448500 133280 1 0 $X=448310 $Y=130320
X3057 1 2 1475 296 1486 ICV_80 $T=471500 165920 0 0 $X=471310 $Y=165680
X3058 1 2 1476 338 1496 ICV_80 $T=473800 122400 0 0 $X=473610 $Y=122160
X3059 1 2 347 343 1503 ICV_80 $T=477940 116960 1 0 $X=477750 $Y=114000
X3060 1 2 347 339 1518 ICV_80 $T=488060 116960 1 0 $X=487870 $Y=114000
X3061 1 2 1548 296 1578 ICV_80 $T=523480 116960 0 0 $X=523290 $Y=116720
X3062 1 2 1625 380 1662 ICV_80 $T=575460 171360 0 0 $X=575270 $Y=171120
X3063 1 2 1625 399 1663 ICV_80 $T=575920 165920 0 0 $X=575730 $Y=165680
X3064 1 2 1668 378 1699 ICV_80 $T=600300 165920 1 0 $X=600110 $Y=162960
X3065 1 2 1844 340 1895 ICV_80 $T=702880 122400 1 0 $X=702690 $Y=119440
X3066 1 2 ICV_81 $T=33580 155040 0 0 $X=33390 $Y=154800
X3067 1 2 ICV_81 $T=47840 127840 1 0 $X=47650 $Y=124880
X3068 1 2 ICV_81 $T=61640 127840 0 0 $X=61450 $Y=127600
X3069 1 2 ICV_81 $T=75900 138720 1 0 $X=75710 $Y=135760
X3070 1 2 ICV_81 $T=145820 138720 0 0 $X=145630 $Y=138480
X3071 1 2 ICV_81 $T=160080 138720 1 0 $X=159890 $Y=135760
X3072 1 2 ICV_81 $T=188140 176800 1 0 $X=187950 $Y=173840
X3073 1 2 ICV_81 $T=272320 165920 1 0 $X=272130 $Y=162960
X3074 1 2 ICV_81 $T=496800 171360 1 0 $X=496610 $Y=168400
X3075 1 2 ICV_81 $T=510600 144160 0 0 $X=510410 $Y=143920
X3076 1 2 ICV_81 $T=552920 138720 1 0 $X=552730 $Y=135760
X3077 1 2 ICV_81 $T=566720 133280 0 0 $X=566530 $Y=133040
X3078 1 2 ICV_81 $T=637100 155040 1 0 $X=636910 $Y=152080
X3079 1 2 ICV_81 $T=650900 165920 0 0 $X=650710 $Y=165680
X3080 1 2 ICV_81 $T=665160 127840 1 0 $X=664970 $Y=124880
X3081 1 2 ICV_81 $T=665160 160480 1 0 $X=664970 $Y=157520
X3099 1 2 168 170 173 2 141 1 sky130_fd_sc_hd__and3b_4 $T=225400 149600 0 0 $X=225210 $Y=149360
X3100 1 2 173 170 168 2 1572 1 sky130_fd_sc_hd__and3b_4 $T=525320 149600 1 0 $X=525130 $Y=146640
.ENDS
***************************************
.SUBCKT ICV_84 1 2 3 4 5 6 7 8 9 10 11
** N=11 EP=11 IP=15 FDC=48
*.SEEDPROM
X0 1 2 3 4 2 5 1 sky130_fd_sc_hd__ebufn_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 9 10 11 6 7 8 ICV_13 $T=4140 0 0 0 $X=3950 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_85 1 2 3 4 5
** N=5 EP=5 IP=9 FDC=26
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=7820 0 0 0 $X=7630 $Y=-240
X1 1 2 3 4 5 ICV_20 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_86 1 2 3 4 5
** N=5 EP=5 IP=11 FDC=20
*.SEEDPROM
X1 1 2 5 3 2 4 1 sky130_fd_sc_hd__dlclkp_1 $T=920 0 0 0 $X=730 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_87 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=14 FDC=18
*.SEEDPROM
X0 1 2 3 4 2 5 1 sky130_fd_sc_hd__ebufn_2 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 6 7 2 8 1 sky130_fd_sc_hd__and2_1 $T=4140 0 0 0 $X=3950 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_88 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 260
+ 261 262 263 264 265 266 267 268 269 270 271 272 273 274 275 276 277 278 279 280
+ 281 282 283 284 285 286 287 288 289 290 291 292 293 294 295 296 297 298 299 300
+ 301 302 303 304 305 306 307 308 309 310 311 312 313 314 315 316 317 318 319 320
+ 321 322 323 324 325 326 327 328 329 330 331 332 333 334 335 336 337 338 339 340
+ 341 342 343 344 345 346 347 348 349 350 351 352 353 354 355 356 357 358 359 360
+ 361 362 363 364 365 366 367 368 369 370 371 372 373 374 375 376 377 378 379 380
+ 381 382 383 384 385 386 387 388 389 390 391 392 393 394 395 396 397 398 399 400
+ 401 402 403 404 405 406 407 408 409 415
** N=1923 EP=410 IP=16464 FDC=47607
*.SEEDPROM
X0 1 2 Dpar a=2090.22 p=1485.84 m=1 $[nwdiode] $X=5330 $Y=52985 $D=191
X1 1 2 Dpar a=2091.12 p=1484.74 m=1 $[nwdiode] $X=5330 $Y=58425 $D=191
X2 1 2 Dpar a=2090.79 p=1485.14 m=1 $[nwdiode] $X=5330 $Y=63865 $D=191
X3 1 2 Dpar a=2091.03 p=1484.84 m=1 $[nwdiode] $X=5330 $Y=69305 $D=191
X4 1 2 Dpar a=2090.55 p=1485.44 m=1 $[nwdiode] $X=5330 $Y=74745 $D=191
X5 1 2 Dpar a=2091.03 p=1484.84 m=1 $[nwdiode] $X=5330 $Y=80185 $D=191
X6 1 2 Dpar a=2090.55 p=1485.44 m=1 $[nwdiode] $X=5330 $Y=85625 $D=191
X7 1 2 Dpar a=2090.47 p=1485.54 m=1 $[nwdiode] $X=5330 $Y=91065 $D=191
X8 1 2 Dpar a=2090.87 p=1485.04 m=1 $[nwdiode] $X=5330 $Y=96505 $D=191
X9 1 2 Dpar a=2091.03 p=1484.84 m=1 $[nwdiode] $X=5330 $Y=101945 $D=191
X10 1 2 Dpar a=2090.63 p=1485.34 m=1 $[nwdiode] $X=5330 $Y=107385 $D=191
X11 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=18400 62560 1 0 $X=18210 $Y=59600
X12 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=18400 78880 0 0 $X=18210 $Y=78640
X13 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=20240 51680 1 0 $X=20050 $Y=48720
X14 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=38180 73440 0 0 $X=37990 $Y=73200
X15 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=40480 78880 0 0 $X=40290 $Y=78640
X16 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=42320 57120 1 0 $X=42130 $Y=54160
X17 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=50600 68000 0 0 $X=50410 $Y=67760
X18 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=57960 84320 0 0 $X=57770 $Y=84080
X19 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=80500 51680 1 0 $X=80310 $Y=48720
X20 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=80960 57120 0 0 $X=80770 $Y=56880
X21 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=95220 84320 1 0 $X=95030 $Y=81360
X22 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=97520 78880 0 0 $X=97330 $Y=78640
X23 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=109020 89760 0 0 $X=108830 $Y=89520
X24 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=118220 51680 0 0 $X=118030 $Y=51440
X25 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=132480 111520 1 0 $X=132290 $Y=108560
X26 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=137080 95200 0 0 $X=136890 $Y=94960
X27 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=150420 106080 1 0 $X=150230 $Y=103120
X28 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=152260 73440 1 0 $X=152070 $Y=70480
X29 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=156400 111520 1 0 $X=156210 $Y=108560
X30 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=156860 111520 0 0 $X=156670 $Y=111280
X31 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=172500 100640 0 0 $X=172310 $Y=100400
X32 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=174340 62560 0 0 $X=174150 $Y=62320
X33 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=187220 57120 0 0 $X=187030 $Y=56880
X34 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=202400 84320 0 0 $X=202210 $Y=84080
X35 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=202400 95200 0 0 $X=202210 $Y=94960
X36 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=207460 57120 1 0 $X=207270 $Y=54160
X37 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=211140 100640 1 0 $X=210950 $Y=97680
X38 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=220800 106080 1 0 $X=220610 $Y=103120
X39 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=224020 106080 0 0 $X=223830 $Y=105840
X40 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=224480 111520 0 0 $X=224290 $Y=111280
X41 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=230460 89760 0 0 $X=230270 $Y=89520
X42 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=235520 111520 1 0 $X=235330 $Y=108560
X43 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=238740 95200 1 0 $X=238550 $Y=92240
X44 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=256680 89760 0 0 $X=256490 $Y=89520
X45 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=266340 111520 0 0 $X=266150 $Y=111280
X46 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=277840 78880 0 0 $X=277650 $Y=78640
X47 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=280600 89760 0 0 $X=280410 $Y=89520
X48 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=284740 106080 0 0 $X=284550 $Y=105840
X49 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=297620 111520 0 0 $X=297430 $Y=111280
X50 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=299000 73440 1 0 $X=298810 $Y=70480
X51 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=300840 51680 1 0 $X=300650 $Y=48720
X52 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=300840 57120 1 0 $X=300650 $Y=54160
X53 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=306360 89760 0 0 $X=306170 $Y=89520
X54 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=312800 62560 0 0 $X=312610 $Y=62320
X55 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=317400 84320 1 0 $X=317210 $Y=81360
X56 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=321080 100640 1 0 $X=320890 $Y=97680
X57 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=322000 73440 0 0 $X=321810 $Y=73200
X58 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=329820 106080 0 0 $X=329630 $Y=105840
X59 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=330280 57120 0 0 $X=330090 $Y=56880
X60 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=373980 51680 1 0 $X=373790 $Y=48720
X61 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=378120 106080 0 0 $X=377930 $Y=105840
X62 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=386400 84320 0 0 $X=386210 $Y=84080
X63 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=398820 68000 0 0 $X=398630 $Y=67760
X64 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=408940 111520 1 0 $X=408750 $Y=108560
X65 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=413080 106080 1 0 $X=412890 $Y=103120
X66 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=426880 100640 0 0 $X=426690 $Y=100400
X67 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=432400 57120 1 0 $X=432210 $Y=54160
X68 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=432400 95200 0 0 $X=432210 $Y=94960
X69 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=434240 57120 0 0 $X=434050 $Y=56880
X70 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=439300 73440 1 0 $X=439110 $Y=70480
X71 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=439300 89760 1 0 $X=439110 $Y=86800
X72 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=459080 62560 0 0 $X=458890 $Y=62320
X73 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=462300 84320 0 0 $X=462110 $Y=84080
X74 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=467360 62560 1 0 $X=467170 $Y=59600
X75 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=468740 111520 0 0 $X=468550 $Y=111280
X76 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=477480 73440 1 0 $X=477290 $Y=70480
X77 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=483000 84320 0 0 $X=482810 $Y=84080
X78 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=488520 95200 0 0 $X=488330 $Y=94960
X79 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=495420 106080 0 0 $X=495230 $Y=105840
X80 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=497260 73440 1 0 $X=497070 $Y=70480
X81 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=516120 78880 1 0 $X=515930 $Y=75920
X82 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=528080 78880 0 0 $X=527890 $Y=78640
X83 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=530840 100640 0 0 $X=530650 $Y=100400
X84 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=533600 57120 1 0 $X=533410 $Y=54160
X85 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=534980 78880 1 0 $X=534790 $Y=75920
X86 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=535900 84320 0 0 $X=535710 $Y=84080
X87 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=547860 57120 0 0 $X=547670 $Y=56880
X88 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=562120 100640 1 0 $X=561930 $Y=97680
X89 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=574540 111520 0 0 $X=574350 $Y=111280
X90 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=577300 89760 1 0 $X=577110 $Y=86800
X91 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=581440 95200 1 0 $X=581250 $Y=92240
X92 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=581440 111520 1 0 $X=581250 $Y=108560
X93 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=595240 73440 0 0 $X=595050 $Y=73200
X94 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=599380 106080 0 0 $X=599190 $Y=105840
X95 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=603060 111520 1 0 $X=602870 $Y=108560
X96 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=621460 78880 0 0 $X=621270 $Y=78640
X97 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=623300 73440 0 0 $X=623110 $Y=73200
X98 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=652740 106080 0 0 $X=652550 $Y=105840
X99 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=654580 68000 1 0 $X=654390 $Y=65040
X100 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=659640 84320 1 0 $X=659450 $Y=81360
X101 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=665160 78880 0 0 $X=664970 $Y=78640
X102 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=672980 89760 1 0 $X=672790 $Y=86800
X103 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=673440 100640 0 0 $X=673250 $Y=100400
X104 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=675280 78880 0 0 $X=675090 $Y=78640
X105 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=677120 95200 1 0 $X=676930 $Y=92240
X106 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=693680 84320 1 0 $X=693490 $Y=81360
X107 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=707480 73440 0 0 $X=707290 $Y=73200
X108 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=719900 89760 1 0 $X=719710 $Y=86800
X109 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=720360 51680 0 0 $X=720170 $Y=51440
X110 1 2 ICV_2 $T=5520 51680 1 0 $X=5330 $Y=48720
X111 1 2 ICV_2 $T=5520 62560 1 0 $X=5330 $Y=59600
X112 1 2 ICV_2 $T=5520 73440 1 0 $X=5330 $Y=70480
X113 1 2 ICV_2 $T=5520 84320 1 0 $X=5330 $Y=81360
X114 1 2 ICV_2 $T=5520 95200 1 0 $X=5330 $Y=92240
X115 1 2 ICV_2 $T=5520 106080 1 0 $X=5330 $Y=103120
X116 1 2 ICV_2 $T=744280 51680 0 180 $X=742710 $Y=48720
X117 1 2 ICV_2 $T=744280 62560 0 180 $X=742710 $Y=59600
X118 1 2 ICV_2 $T=744280 73440 0 180 $X=742710 $Y=70480
X119 1 2 ICV_2 $T=744280 84320 0 180 $X=742710 $Y=81360
X120 1 2 ICV_2 $T=744280 95200 0 180 $X=742710 $Y=92240
X121 1 2 ICV_2 $T=744280 106080 0 180 $X=742710 $Y=103120
X273 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=6900 95200 0 0 $X=6710 $Y=94960
X274 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17480 68000 0 0 $X=17290 $Y=67760
X275 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17480 111520 1 0 $X=17290 $Y=108560
X276 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 73440 1 0 $X=17750 $Y=70480
X277 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=38640 89760 1 0 $X=38450 $Y=86800
X278 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=43700 84320 0 0 $X=43510 $Y=84080
X279 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=59800 51680 0 0 $X=59610 $Y=51440
X280 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=62100 78880 0 0 $X=61910 $Y=78640
X281 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=76360 84320 1 0 $X=76170 $Y=81360
X282 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=88320 100640 1 0 $X=88130 $Y=97680
X283 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=94760 89760 1 0 $X=94570 $Y=86800
X284 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=102120 57120 0 0 $X=101930 $Y=56880
X285 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=104420 57120 1 0 $X=104230 $Y=54160
X286 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=129720 78880 1 0 $X=129530 $Y=75920
X287 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=129720 84320 1 0 $X=129530 $Y=81360
X288 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=146280 68000 0 0 $X=146090 $Y=67760
X289 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=155020 57120 0 0 $X=154830 $Y=56880
X290 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=160540 57120 1 0 $X=160350 $Y=54160
X291 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=160540 78880 1 0 $X=160350 $Y=75920
X292 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=160540 89760 1 0 $X=160350 $Y=86800
X293 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=164680 111520 0 0 $X=164490 $Y=111280
X294 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=181700 106080 0 0 $X=181510 $Y=105840
X295 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=186300 84320 1 0 $X=186110 $Y=81360
X296 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=192280 100640 0 0 $X=192090 $Y=100400
X297 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=202400 100640 0 0 $X=202210 $Y=100400
X298 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=206080 111520 1 0 $X=205890 $Y=108560
X299 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=208380 95200 0 0 $X=208190 $Y=94960
X300 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=214360 84320 1 0 $X=214170 $Y=81360
X301 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=214360 111520 0 0 $X=214170 $Y=111280
X302 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=216660 68000 1 0 $X=216470 $Y=65040
X303 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=219420 78880 0 0 $X=219230 $Y=78640
X304 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=283820 111520 0 0 $X=283630 $Y=111280
X305 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=333960 78880 0 0 $X=333770 $Y=78640
X306 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=339940 106080 0 0 $X=339750 $Y=105840
X307 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=350980 106080 0 0 $X=350790 $Y=105840
X308 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=368460 89760 0 0 $X=368270 $Y=89520
X309 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=370760 100640 0 0 $X=370570 $Y=100400
X310 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=385020 84320 1 0 $X=384830 $Y=81360
X311 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=398820 51680 0 0 $X=398630 $Y=51440
X312 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=406180 57120 0 0 $X=405990 $Y=56880
X313 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=406180 106080 0 0 $X=405990 $Y=105840
X314 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=415840 51680 0 0 $X=415650 $Y=51440
X315 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=417220 73440 0 0 $X=417030 $Y=73200
X316 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=426880 111520 0 0 $X=426690 $Y=111280
X317 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=452180 73440 0 0 $X=451990 $Y=73200
X318 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=454940 78880 0 0 $X=454750 $Y=78640
X319 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=459080 111520 0 0 $X=458890 $Y=111280
X320 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=464140 95200 0 0 $X=463950 $Y=94960
X321 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=469200 51680 1 0 $X=469010 $Y=48720
X322 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=490820 73440 1 0 $X=490630 $Y=70480
X323 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=494500 78880 1 0 $X=494310 $Y=75920
X324 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=497260 78880 1 0 $X=497070 $Y=75920
X325 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=533600 111520 1 0 $X=533410 $Y=108560
X326 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=536360 111520 0 0 $X=536170 $Y=111280
X327 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=596160 57120 1 0 $X=595970 $Y=54160
X328 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=603520 95200 0 0 $X=603330 $Y=94960
X329 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=607200 78880 1 0 $X=607010 $Y=75920
X330 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=635260 100640 1 0 $X=635070 $Y=97680
X331 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=644920 106080 1 0 $X=644730 $Y=103120
X332 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=658720 62560 0 0 $X=658530 $Y=62320
X333 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=658720 100640 0 0 $X=658530 $Y=100400
X334 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=659640 89760 0 0 $X=659450 $Y=89520
X335 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=704720 51680 0 0 $X=704530 $Y=51440
X336 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=704720 106080 0 0 $X=704530 $Y=105840
X337 1 2 ICV_3 $T=16100 95200 1 0 $X=15910 $Y=92240
X338 1 2 ICV_3 $T=17020 84320 0 0 $X=16830 $Y=84080
X339 1 2 ICV_3 $T=34040 106080 0 0 $X=33850 $Y=105840
X340 1 2 ICV_3 $T=48300 78880 1 0 $X=48110 $Y=75920
X341 1 2 ICV_3 $T=55200 106080 0 0 $X=55010 $Y=105840
X342 1 2 ICV_3 $T=81880 89760 0 0 $X=81690 $Y=89520
X343 1 2 ICV_3 $T=101660 73440 1 0 $X=101470 $Y=70480
X344 1 2 ICV_3 $T=132480 106080 1 0 $X=132290 $Y=103120
X345 1 2 ICV_3 $T=139380 84320 0 0 $X=139190 $Y=84080
X346 1 2 ICV_3 $T=168820 51680 1 0 $X=168630 $Y=48720
X347 1 2 ICV_3 $T=169280 111520 1 0 $X=169090 $Y=108560
X348 1 2 ICV_3 $T=181700 100640 0 0 $X=181510 $Y=100400
X349 1 2 ICV_3 $T=216660 89760 1 0 $X=216470 $Y=86800
X350 1 2 ICV_3 $T=291640 68000 1 0 $X=291450 $Y=65040
X351 1 2 ICV_3 $T=300380 68000 0 0 $X=300190 $Y=67760
X352 1 2 ICV_3 $T=304980 100640 1 0 $X=304790 $Y=97680
X353 1 2 ICV_3 $T=314640 51680 0 0 $X=314450 $Y=51440
X354 1 2 ICV_3 $T=354200 89760 1 0 $X=354010 $Y=86800
X355 1 2 ICV_3 $T=359260 106080 0 0 $X=359070 $Y=105840
X356 1 2 ICV_3 $T=373980 100640 1 0 $X=373790 $Y=97680
X357 1 2 ICV_3 $T=379960 111520 0 0 $X=379770 $Y=111280
X358 1 2 ICV_3 $T=396060 57120 0 0 $X=395870 $Y=56880
X359 1 2 ICV_3 $T=434240 95200 1 0 $X=434050 $Y=92240
X360 1 2 ICV_3 $T=465060 78880 0 0 $X=464870 $Y=78640
X361 1 2 ICV_3 $T=480240 100640 0 0 $X=480050 $Y=100400
X362 1 2 ICV_3 $T=490360 100640 0 0 $X=490170 $Y=100400
X363 1 2 ICV_3 $T=506000 57120 1 0 $X=505810 $Y=54160
X364 1 2 ICV_3 $T=543260 84320 0 0 $X=543070 $Y=84080
X365 1 2 ICV_3 $T=564420 68000 0 0 $X=564230 $Y=67760
X366 1 2 ICV_3 $T=564880 78880 1 0 $X=564690 $Y=75920
X367 1 2 ICV_3 $T=574540 100640 0 0 $X=574350 $Y=100400
X368 1 2 ICV_3 $T=580060 111520 0 0 $X=579870 $Y=111280
X369 1 2 ICV_3 $T=580980 89760 0 0 $X=580790 $Y=89520
X370 1 2 ICV_3 $T=591560 73440 1 0 $X=591370 $Y=70480
X371 1 2 ICV_3 $T=634800 73440 1 0 $X=634610 $Y=70480
X372 1 2 ICV_3 $T=634800 95200 1 0 $X=634610 $Y=92240
X373 1 2 ICV_3 $T=651360 57120 0 0 $X=651170 $Y=56880
X374 1 2 ICV_3 $T=653200 57120 1 0 $X=653010 $Y=54160
X375 1 2 ICV_3 $T=662860 68000 0 0 $X=662670 $Y=67760
X376 1 2 ICV_3 $T=662860 89760 1 0 $X=662670 $Y=86800
X377 1 2 ICV_3 $T=677120 111520 1 0 $X=676930 $Y=108560
X378 1 2 ICV_3 $T=693680 89760 1 0 $X=693490 $Y=86800
X379 1 2 ICV_3 $T=712540 51680 1 0 $X=712350 $Y=48720
X380 1 2 ICV_3 $T=718980 73440 1 0 $X=718790 $Y=70480
X381 1 2 ICV_3 $T=732780 62560 0 0 $X=732590 $Y=62320
X382 1 2 ICV_3 $T=732780 78880 0 0 $X=732590 $Y=78640
X383 1 2 ICV_3 $T=735540 51680 0 0 $X=735350 $Y=51440
X384 1 2 ICV_3 $T=735540 73440 0 0 $X=735350 $Y=73200
X385 1 2 ICV_3 $T=735540 106080 0 0 $X=735350 $Y=105840
X386 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=6900 84320 0 0 $X=6710 $Y=84080
X387 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=6900 106080 0 0 $X=6710 $Y=105840
X388 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=22540 73440 0 0 $X=22350 $Y=73200
X389 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=26680 73440 1 0 $X=26490 $Y=70480
X390 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=48300 106080 1 0 $X=48110 $Y=103120
X391 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=54280 73440 0 0 $X=54090 $Y=73200
X392 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=67160 84320 1 0 $X=66970 $Y=81360
X393 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=72680 62560 1 0 $X=72490 $Y=59600
X394 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=86480 95200 0 0 $X=86290 $Y=94960
X395 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=90160 84320 0 0 $X=89970 $Y=84080
X396 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=100740 78880 1 0 $X=100550 $Y=75920
X397 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=104420 78880 1 0 $X=104230 $Y=75920
X398 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=107180 73440 0 0 $X=106990 $Y=73200
X399 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=111780 106080 1 0 $X=111590 $Y=103120
X400 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=112700 57120 1 0 $X=112510 $Y=54160
X401 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=115000 51680 0 0 $X=114810 $Y=51440
X402 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=115000 100640 0 0 $X=114810 $Y=100400
X403 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=146280 100640 1 0 $X=146090 $Y=97680
X404 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=152720 51680 1 0 $X=152530 $Y=48720
X405 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=174340 89760 0 0 $X=174150 $Y=89520
X406 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=198720 100640 0 0 $X=198530 $Y=100400
X407 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=198720 106080 0 0 $X=198530 $Y=105840
X408 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=213440 62560 1 0 $X=213250 $Y=59600
X409 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=215280 73440 0 0 $X=215090 $Y=73200
X410 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=222640 73440 0 0 $X=222450 $Y=73200
X411 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=232300 106080 1 0 $X=232110 $Y=103120
X412 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=234600 78880 0 0 $X=234410 $Y=78640
X413 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=251160 68000 0 0 $X=250970 $Y=67760
X414 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=282900 68000 0 0 $X=282710 $Y=67760
X415 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=282900 95200 0 0 $X=282710 $Y=94960
X416 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=283360 57120 0 0 $X=283170 $Y=56880
X417 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=308200 73440 1 0 $X=308010 $Y=70480
X418 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=310960 68000 0 0 $X=310770 $Y=67760
X419 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=314640 68000 0 0 $X=314450 $Y=67760
X420 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=318780 106080 0 0 $X=318590 $Y=105840
X421 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=325680 51680 1 0 $X=325490 $Y=48720
X422 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=325680 73440 1 0 $X=325490 $Y=70480
X423 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=328900 68000 0 0 $X=328710 $Y=67760
X424 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=353280 95200 1 0 $X=353090 $Y=92240
X425 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=356960 73440 1 0 $X=356770 $Y=70480
X426 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=364320 106080 1 0 $X=364130 $Y=103120
X427 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=389160 100640 1 0 $X=388970 $Y=97680
X428 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=395600 106080 0 0 $X=395410 $Y=105840
X429 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=409400 84320 1 0 $X=409210 $Y=81360
X430 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=409860 62560 1 0 $X=409670 $Y=59600
X431 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=423200 62560 0 0 $X=423010 $Y=62320
X432 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=423660 57120 0 0 $X=423470 $Y=56880
X433 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=454940 73440 0 0 $X=454750 $Y=73200
X434 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=455860 95200 1 0 $X=455670 $Y=92240
X435 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=457240 62560 1 0 $X=457050 $Y=59600
X436 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=476560 89760 1 0 $X=476370 $Y=86800
X437 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=478860 57120 1 0 $X=478670 $Y=54160
X438 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=479320 106080 0 0 $X=479130 $Y=105840
X439 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=496340 95200 0 0 $X=496150 $Y=94960
X440 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=511060 111520 0 0 $X=510870 $Y=111280
X441 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=517040 95200 1 0 $X=516850 $Y=92240
X442 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=528080 89760 0 0 $X=527890 $Y=89520
X443 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=547400 78880 0 0 $X=547210 $Y=78640
X444 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=567180 84320 0 0 $X=566990 $Y=84080
X445 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=567180 111520 0 0 $X=566990 $Y=111280
X446 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=581440 51680 1 0 $X=581250 $Y=48720
X447 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=581440 68000 1 0 $X=581250 $Y=65040
X448 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=581440 73440 1 0 $X=581250 $Y=70480
X449 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=585580 84320 1 0 $X=585390 $Y=81360
X450 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=620080 62560 0 0 $X=619890 $Y=62320
X451 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=623300 68000 0 0 $X=623110 $Y=67760
X452 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=634340 84320 1 0 $X=634150 $Y=81360
X453 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=638940 62560 1 0 $X=638750 $Y=59600
X454 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=651360 95200 0 0 $X=651170 $Y=94960
X455 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=667000 62560 0 0 $X=666810 $Y=62320
X456 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=667000 100640 0 0 $X=666810 $Y=100400
X457 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=683560 111520 0 0 $X=683370 $Y=111280
X458 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=698740 62560 0 0 $X=698550 $Y=62320
X459 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=718060 68000 1 0 $X=717870 $Y=65040
X460 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=729100 73440 1 0 $X=728910 $Y=70480
X461 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=731860 73440 0 0 $X=731670 $Y=73200
X462 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=731860 106080 0 0 $X=731670 $Y=105840
X463 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=732320 111520 0 0 $X=732130 $Y=111280
X464 1 2 ICV_4 $T=34040 84320 0 0 $X=33850 $Y=84080
X465 1 2 ICV_4 $T=44620 68000 1 0 $X=44430 $Y=65040
X466 1 2 ICV_4 $T=62560 106080 1 0 $X=62370 $Y=103120
X467 1 2 ICV_4 $T=184920 111520 0 0 $X=184730 $Y=111280
X468 1 2 ICV_4 $T=202400 111520 0 0 $X=202210 $Y=111280
X469 1 2 ICV_4 $T=218040 89760 0 0 $X=217850 $Y=89520
X470 1 2 ICV_4 $T=221260 95200 1 0 $X=221070 $Y=92240
X471 1 2 ICV_4 $T=339020 73440 0 0 $X=338830 $Y=73200
X472 1 2 ICV_4 $T=340400 78880 1 0 $X=340210 $Y=75920
X473 1 2 ICV_4 $T=367080 78880 0 0 $X=366890 $Y=78640
X474 1 2 ICV_4 $T=406180 78880 0 0 $X=405990 $Y=78640
X475 1 2 ICV_4 $T=445280 57120 1 0 $X=445090 $Y=54160
X476 1 2 ICV_4 $T=462300 100640 0 0 $X=462110 $Y=100400
X477 1 2 ICV_4 $T=511060 100640 1 0 $X=510870 $Y=97680
X478 1 2 ICV_4 $T=527620 73440 0 0 $X=527430 $Y=73200
X479 1 2 ICV_4 $T=543260 106080 0 0 $X=543070 $Y=105840
X480 1 2 ICV_4 $T=549700 100640 1 0 $X=549510 $Y=97680
X481 1 2 ICV_4 $T=603520 89760 1 0 $X=603330 $Y=86800
X482 1 2 ICV_4 $T=627440 51680 1 0 $X=627250 $Y=48720
X483 1 2 ICV_4 $T=648140 51680 1 0 $X=647950 $Y=48720
X484 1 2 ICV_4 $T=675740 84320 0 0 $X=675550 $Y=84080
X485 1 2 ICV_4 $T=721740 95200 1 0 $X=721550 $Y=92240
X486 1 2 ICV_4 $T=731860 57120 0 0 $X=731670 $Y=56880
X487 1 2 ICV_4 $T=731860 68000 0 0 $X=731670 $Y=67760
X488 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 51680 0 0 $X=6710 $Y=51440
X489 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 57120 1 0 $X=6710 $Y=54160
X490 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 62560 1 0 $X=6710 $Y=59600
X491 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 62560 0 0 $X=6710 $Y=62320
X492 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 68000 1 0 $X=6710 $Y=65040
X493 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 73440 0 0 $X=6710 $Y=73200
X494 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 78880 1 0 $X=6710 $Y=75920
X495 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 78880 0 0 $X=6710 $Y=78640
X496 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 84320 1 0 $X=6710 $Y=81360
X497 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 89760 1 0 $X=6710 $Y=86800
X498 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 100640 0 0 $X=6710 $Y=100400
X499 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 106080 1 0 $X=6710 $Y=103120
X500 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=12420 57120 0 0 $X=12230 $Y=56880
X501 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=49220 95200 0 0 $X=49030 $Y=94960
X502 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=62100 106080 0 0 $X=61910 $Y=105840
X503 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=76360 62560 1 0 $X=76170 $Y=59600
X504 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=78200 51680 0 0 $X=78010 $Y=51440
X505 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=91080 57120 1 0 $X=90890 $Y=54160
X506 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=102580 68000 0 0 $X=102390 $Y=67760
X507 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=116840 100640 1 0 $X=116650 $Y=97680
X508 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=132480 84320 1 0 $X=132290 $Y=81360
X509 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=148120 57120 1 0 $X=147930 $Y=54160
X510 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=161000 73440 0 0 $X=160810 $Y=73200
X511 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=168820 100640 1 0 $X=168630 $Y=97680
X512 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=174340 73440 0 0 $X=174150 $Y=73200
X513 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=174800 73440 1 0 $X=174610 $Y=70480
X514 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=183540 95200 0 0 $X=183350 $Y=94960
X515 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=188600 106080 1 0 $X=188410 $Y=103120
X516 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=211600 89760 1 0 $X=211410 $Y=86800
X517 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=215740 57120 0 0 $X=215550 $Y=56880
X518 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=226320 62560 0 0 $X=226130 $Y=62320
X519 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=230460 68000 1 0 $X=230270 $Y=65040
X520 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=249780 51680 0 0 $X=249590 $Y=51440
X521 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=251620 89760 0 0 $X=251430 $Y=89520
X522 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=261280 68000 1 0 $X=261090 $Y=65040
X523 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=262660 62560 0 0 $X=262470 $Y=62320
X524 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=268640 78880 1 0 $X=268450 $Y=75920
X525 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=296700 62560 1 0 $X=296510 $Y=59600
X526 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=299920 106080 0 0 $X=299730 $Y=105840
X527 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=309120 62560 0 0 $X=308930 $Y=62320
X528 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=310500 73440 0 0 $X=310310 $Y=73200
X529 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=312800 106080 1 0 $X=312610 $Y=103120
X530 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=322460 78880 0 0 $X=322270 $Y=78640
X531 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=324760 106080 1 0 $X=324570 $Y=103120
X532 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=351900 78880 1 0 $X=351710 $Y=75920
X533 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=370300 51680 1 0 $X=370110 $Y=48720
X534 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=389160 57120 1 0 $X=388970 $Y=54160
X535 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=398820 95200 0 0 $X=398630 $Y=94960
X536 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=408940 100640 1 0 $X=408750 $Y=97680
X537 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=422280 68000 0 0 $X=422090 $Y=67760
X538 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=426880 68000 0 0 $X=426690 $Y=67760
X539 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=436080 78880 1 0 $X=435890 $Y=75920
X540 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=441140 51680 1 0 $X=440950 $Y=48720
X541 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=442980 78880 0 0 $X=442790 $Y=78640
X542 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=445280 84320 1 0 $X=445090 $Y=81360
X543 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=445280 106080 1 0 $X=445090 $Y=103120
X544 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=460000 73440 1 0 $X=459810 $Y=70480
X545 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=460920 100640 1 0 $X=460730 $Y=97680
X546 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=465060 73440 0 0 $X=464870 $Y=73200
X547 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=469200 73440 1 0 $X=469010 $Y=70480
X548 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=526700 62560 0 0 $X=526510 $Y=62320
X549 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=553380 95200 1 0 $X=553190 $Y=92240
X550 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=583740 73440 0 0 $X=583550 $Y=73200
X551 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=595240 84320 0 0 $X=595050 $Y=84080
X552 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=595240 95200 1 0 $X=595050 $Y=92240
X553 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=611800 111520 0 0 $X=611610 $Y=111280
X554 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=633420 111520 1 0 $X=633230 $Y=108560
X555 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=638940 106080 0 0 $X=638750 $Y=105840
X556 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=641700 111520 1 0 $X=641510 $Y=108560
X557 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=644920 73440 1 0 $X=644730 $Y=70480
X558 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=675280 95200 0 0 $X=675090 $Y=94960
X559 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=679420 57120 0 0 $X=679230 $Y=56880
X560 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=683560 68000 0 0 $X=683370 $Y=67760
X561 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=689080 51680 0 0 $X=688890 $Y=51440
X562 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=707480 62560 0 0 $X=707290 $Y=62320
X563 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=717600 62560 1 0 $X=717410 $Y=59600
X564 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=731400 100640 0 0 $X=731210 $Y=100400
X565 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=739220 73440 1 0 $X=739030 $Y=70480
X566 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=739220 89760 1 0 $X=739030 $Y=86800
X567 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 51680 1 0 $X=6710 $Y=48720
X568 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 57120 0 0 $X=6710 $Y=56880
X569 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 73440 1 0 $X=6710 $Y=70480
X570 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 100640 1 0 $X=6710 $Y=97680
X571 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=12420 73440 1 0 $X=12230 $Y=70480
X572 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=27140 57120 0 0 $X=26950 $Y=56880
X573 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=34960 106080 1 0 $X=34770 $Y=103120
X574 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=247020 100640 0 0 $X=246830 $Y=100400
X575 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=266800 95200 1 0 $X=266610 $Y=92240
X576 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=316940 78880 0 0 $X=316750 $Y=78640
X577 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=347760 95200 1 0 $X=347570 $Y=92240
X578 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=354660 89760 0 0 $X=354470 $Y=89520
X579 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=356960 95200 1 0 $X=356770 $Y=92240
X580 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=392840 78880 0 0 $X=392650 $Y=78640
X581 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=400660 89760 1 0 $X=400470 $Y=86800
X582 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=483000 95200 0 0 $X=482810 $Y=94960
X583 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=485760 57120 1 0 $X=485570 $Y=54160
X584 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=621000 106080 1 0 $X=620810 $Y=103120
X585 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=631120 89760 1 0 $X=630930 $Y=86800
X586 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=649060 68000 1 0 $X=648870 $Y=65040
X587 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=683560 51680 0 0 $X=683370 $Y=51440
X588 1 2 450 451 2 11 1 sky130_fd_sc_hd__ebufn_2 $T=8740 95200 0 0 $X=8550 $Y=94960
X589 1 2 480 9 2 18 1 sky130_fd_sc_hd__ebufn_2 $T=21620 51680 1 0 $X=21430 $Y=48720
X590 1 2 506 14 2 33 1 sky130_fd_sc_hd__ebufn_2 $T=36340 106080 0 0 $X=36150 $Y=105840
X591 1 2 491 476 2 30 1 sky130_fd_sc_hd__ebufn_2 $T=40480 68000 1 0 $X=40290 $Y=65040
X592 1 2 498 14 2 34 1 sky130_fd_sc_hd__ebufn_2 $T=40480 111520 0 0 $X=40290 $Y=111280
X593 1 2 546 508 2 30 1 sky130_fd_sc_hd__ebufn_2 $T=85560 78880 0 0 $X=85370 $Y=78640
X594 1 2 585 563 2 32 1 sky130_fd_sc_hd__ebufn_2 $T=90160 95200 0 0 $X=89970 $Y=94960
X595 1 2 625 586 2 30 1 sky130_fd_sc_hd__ebufn_2 $T=97520 73440 1 0 $X=97330 $Y=70480
X596 1 2 631 632 2 20 1 sky130_fd_sc_hd__ebufn_2 $T=99820 68000 1 0 $X=99630 $Y=65040
X597 1 2 657 658 2 30 1 sky130_fd_sc_hd__ebufn_2 $T=113620 84320 0 0 $X=113430 $Y=84080
X598 1 2 660 80 2 32 1 sky130_fd_sc_hd__ebufn_2 $T=119600 62560 1 0 $X=119410 $Y=59600
X599 1 2 749 748 2 32 1 sky130_fd_sc_hd__ebufn_2 $T=156860 73440 0 0 $X=156670 $Y=73200
X600 1 2 806 810 2 32 1 sky130_fd_sc_hd__ebufn_2 $T=201480 68000 1 0 $X=201290 $Y=65040
X601 1 2 815 817 2 11 1 sky130_fd_sc_hd__ebufn_2 $T=206080 89760 1 0 $X=205890 $Y=86800
X602 1 2 852 856 2 18 1 sky130_fd_sc_hd__ebufn_2 $T=218500 68000 1 0 $X=218310 $Y=65040
X603 1 2 869 857 2 30 1 sky130_fd_sc_hd__ebufn_2 $T=225860 78880 0 0 $X=225670 $Y=78640
X604 1 2 878 856 2 30 1 sky130_fd_sc_hd__ebufn_2 $T=231840 89760 0 0 $X=231650 $Y=89520
X605 1 2 889 891 2 170 1 sky130_fd_sc_hd__ebufn_2 $T=240120 95200 1 0 $X=239930 $Y=92240
X606 1 2 906 179 2 182 1 sky130_fd_sc_hd__ebufn_2 $T=245640 111520 1 0 $X=245450 $Y=108560
X607 1 2 954 201 2 177 1 sky130_fd_sc_hd__ebufn_2 $T=272780 51680 1 0 $X=272590 $Y=48720
X608 1 2 1002 988 2 171 1 sky130_fd_sc_hd__ebufn_2 $T=296240 78880 1 0 $X=296050 $Y=75920
X609 1 2 1007 977 2 171 1 sky130_fd_sc_hd__ebufn_2 $T=302220 84320 0 0 $X=302030 $Y=84080
X610 1 2 1019 1018 2 193 1 sky130_fd_sc_hd__ebufn_2 $T=304980 62560 0 0 $X=304790 $Y=62320
X611 1 2 1040 1018 2 195 1 sky130_fd_sc_hd__ebufn_2 $T=316940 51680 0 0 $X=316750 $Y=51440
X612 1 2 1077 1039 2 195 1 sky130_fd_sc_hd__ebufn_2 $T=333960 84320 1 0 $X=333770 $Y=81360
X613 1 2 1167 1149 2 193 1 sky130_fd_sc_hd__ebufn_2 $T=376740 62560 1 0 $X=376550 $Y=59600
X614 1 2 1197 233 2 180 1 sky130_fd_sc_hd__ebufn_2 $T=393760 57120 1 0 $X=393570 $Y=54160
X615 1 2 1203 1199 2 180 1 sky130_fd_sc_hd__ebufn_2 $T=396520 89760 1 0 $X=396330 $Y=86800
X616 1 2 1201 1168 2 191 1 sky130_fd_sc_hd__ebufn_2 $T=398360 106080 1 0 $X=398170 $Y=103120
X617 1 2 1241 1212 2 174 1 sky130_fd_sc_hd__ebufn_2 $T=414460 106080 1 0 $X=414270 $Y=103120
X618 1 2 254 256 2 174 1 sky130_fd_sc_hd__ebufn_2 $T=428720 111520 0 0 $X=428530 $Y=111280
X619 1 2 1285 1270 2 170 1 sky130_fd_sc_hd__ebufn_2 $T=436540 95200 1 0 $X=436350 $Y=92240
X620 1 2 1313 252 2 171 1 sky130_fd_sc_hd__ebufn_2 $T=454940 51680 0 0 $X=454750 $Y=51440
X621 1 2 1338 1333 2 277 1 sky130_fd_sc_hd__ebufn_2 $T=464600 89760 1 0 $X=464410 $Y=86800
X622 1 2 1373 1312 2 277 1 sky130_fd_sc_hd__ebufn_2 $T=478400 68000 0 0 $X=478210 $Y=67760
X623 1 2 1366 1331 2 275 1 sky130_fd_sc_hd__ebufn_2 $T=478400 89760 0 0 $X=478210 $Y=89520
X624 1 2 1372 1333 2 280 1 sky130_fd_sc_hd__ebufn_2 $T=478860 73440 1 0 $X=478670 $Y=70480
X625 1 2 1377 1333 2 275 1 sky130_fd_sc_hd__ebufn_2 $T=479320 89760 1 0 $X=479130 $Y=86800
X626 1 2 1379 1357 2 300 1 sky130_fd_sc_hd__ebufn_2 $T=481620 57120 1 0 $X=481430 $Y=54160
X627 1 2 1411 1386 2 296 1 sky130_fd_sc_hd__ebufn_2 $T=498180 68000 1 0 $X=497990 $Y=65040
X628 1 2 1414 1399 2 303 1 sky130_fd_sc_hd__ebufn_2 $T=500480 95200 0 0 $X=500290 $Y=94960
X629 1 2 1430 298 2 304 1 sky130_fd_sc_hd__ebufn_2 $T=506460 100640 0 0 $X=506270 $Y=100400
X630 1 2 1480 1446 2 304 1 sky130_fd_sc_hd__ebufn_2 $T=536820 100640 1 0 $X=536630 $Y=97680
X631 1 2 1516 334 2 300 1 sky130_fd_sc_hd__ebufn_2 $T=548780 57120 1 0 $X=548590 $Y=54160
X632 1 2 1523 1525 2 269 1 sky130_fd_sc_hd__ebufn_2 $T=552000 84320 0 0 $X=551810 $Y=84080
X633 1 2 1547 1551 2 268 1 sky130_fd_sc_hd__ebufn_2 $T=562580 100640 0 0 $X=562390 $Y=100400
X634 1 2 1539 333 2 304 1 sky130_fd_sc_hd__ebufn_2 $T=562580 106080 0 0 $X=562390 $Y=105840
X635 1 2 344 345 2 269 1 sky130_fd_sc_hd__ebufn_2 $T=575920 111520 0 0 $X=575730 $Y=111280
X636 1 2 1573 1565 2 273 1 sky130_fd_sc_hd__ebufn_2 $T=576840 89760 0 0 $X=576650 $Y=89520
X637 1 2 347 340 2 307 1 sky130_fd_sc_hd__ebufn_2 $T=579140 51680 0 0 $X=578950 $Y=51440
X638 1 2 1581 1582 2 269 1 sky130_fd_sc_hd__ebufn_2 $T=582360 62560 1 0 $X=582170 $Y=59600
X639 1 2 1606 1582 2 276 1 sky130_fd_sc_hd__ebufn_2 $T=593860 68000 1 0 $X=593670 $Y=65040
X640 1 2 1614 1600 2 273 1 sky130_fd_sc_hd__ebufn_2 $T=596160 100640 0 0 $X=595970 $Y=100400
X641 1 2 1609 1612 2 277 1 sky130_fd_sc_hd__ebufn_2 $T=599380 89760 1 0 $X=599190 $Y=86800
X642 1 2 1608 1612 2 275 1 sky130_fd_sc_hd__ebufn_2 $T=602600 78880 0 0 $X=602410 $Y=78640
X643 1 2 1693 1688 2 276 1 sky130_fd_sc_hd__ebufn_2 $T=634800 106080 0 0 $X=634610 $Y=105840
X644 1 2 1717 1697 2 267 1 sky130_fd_sc_hd__ebufn_2 $T=646760 100640 0 0 $X=646570 $Y=100400
X645 1 2 1728 1697 2 269 1 sky130_fd_sc_hd__ebufn_2 $T=654120 95200 0 0 $X=653930 $Y=94960
X646 1 2 1757 384 2 309 1 sky130_fd_sc_hd__ebufn_2 $T=669760 62560 0 0 $X=669570 $Y=62320
X647 1 2 1778 384 2 294 1 sky130_fd_sc_hd__ebufn_2 $T=679420 51680 0 0 $X=679230 $Y=51440
X648 1 2 1779 1748 2 304 1 sky130_fd_sc_hd__ebufn_2 $T=679420 68000 0 0 $X=679230 $Y=67760
X649 1 2 1793 1798 2 294 1 sky130_fd_sc_hd__ebufn_2 $T=687240 68000 0 0 $X=687050 $Y=67760
X650 1 2 1832 1824 2 304 1 sky130_fd_sc_hd__ebufn_2 $T=708400 51680 1 0 $X=708210 $Y=48720
X651 1 2 1843 1816 2 304 1 sky130_fd_sc_hd__ebufn_2 $T=710240 78880 1 0 $X=710050 $Y=75920
X763 1 2 466 476 18 ICV_6 $T=19780 62560 1 0 $X=19590 $Y=59600
X764 1 2 462 476 17 ICV_6 $T=19780 68000 1 0 $X=19590 $Y=65040
X765 1 2 471 477 11 ICV_6 $T=19780 73440 1 0 $X=19590 $Y=70480
X766 1 2 464 477 17 ICV_6 $T=19780 78880 1 0 $X=19590 $Y=75920
X767 1 2 468 477 18 ICV_6 $T=19780 84320 1 0 $X=19590 $Y=81360
X768 1 2 458 473 18 ICV_6 $T=19780 89760 1 0 $X=19590 $Y=86800
X769 1 2 465 451 20 ICV_6 $T=19780 100640 1 0 $X=19590 $Y=97680
X770 1 2 502 9 32 ICV_6 $T=33580 57120 0 0 $X=33390 $Y=56880
X771 1 2 487 477 33 ICV_6 $T=33580 73440 0 0 $X=33390 $Y=73200
X772 1 2 493 477 34 ICV_6 $T=33580 78880 0 0 $X=33390 $Y=78640
X773 1 2 529 534 11 ICV_6 $T=47840 100640 1 0 $X=47650 $Y=97680
X774 1 2 532 534 20 ICV_6 $T=47840 111520 1 0 $X=47650 $Y=108560
X775 1 2 519 525 30 ICV_6 $T=61640 62560 0 0 $X=61450 $Y=62320
X776 1 2 580 53 33 ICV_6 $T=75900 51680 1 0 $X=75710 $Y=48720
X777 1 2 637 615 18 ICV_6 $T=103960 84320 1 0 $X=103770 $Y=81360
X778 1 2 621 68 34 ICV_6 $T=103960 95200 1 0 $X=103770 $Y=92240
X779 1 2 659 80 33 ICV_6 $T=117760 57120 0 0 $X=117570 $Y=56880
X780 1 2 665 632 18 ICV_6 $T=117760 68000 0 0 $X=117570 $Y=67760
X781 1 2 668 632 32 ICV_6 $T=117760 73440 0 0 $X=117570 $Y=73200
X782 1 2 669 643 17 ICV_6 $T=117760 84320 0 0 $X=117570 $Y=84080
X783 1 2 662 643 18 ICV_6 $T=117760 95200 0 0 $X=117570 $Y=94960
X784 1 2 686 658 34 ICV_6 $T=132020 89760 1 0 $X=131830 $Y=86800
X785 1 2 711 658 17 ICV_6 $T=145820 78880 0 0 $X=145630 $Y=78640
X786 1 2 721 86 34 ICV_6 $T=145820 100640 0 0 $X=145630 $Y=100400
X787 1 2 720 95 96 ICV_6 $T=145820 111520 0 0 $X=145630 $Y=111280
X788 1 2 763 760 20 ICV_6 $T=173880 57120 0 0 $X=173690 $Y=56880
X789 1 2 774 760 30 ICV_6 $T=188140 62560 1 0 $X=187950 $Y=59600
X790 1 2 825 114 34 ICV_6 $T=201940 51680 0 0 $X=201750 $Y=51440
X791 1 2 812 810 17 ICV_6 $T=201940 57120 0 0 $X=201750 $Y=56880
X792 1 2 873 857 32 ICV_6 $T=230000 78880 0 0 $X=229810 $Y=78640
X793 1 2 874 857 17 ICV_6 $T=230000 84320 0 0 $X=229810 $Y=84080
X794 1 2 904 890 180 ICV_6 $T=244260 73440 1 0 $X=244070 $Y=70480
X795 1 2 900 886 177 ICV_6 $T=244260 89760 1 0 $X=244070 $Y=86800
X796 1 2 893 891 182 ICV_6 $T=244260 95200 1 0 $X=244070 $Y=92240
X797 1 2 927 176 192 ICV_6 $T=258060 51680 0 0 $X=257870 $Y=51440
X798 1 2 925 890 195 ICV_6 $T=258060 62560 0 0 $X=257870 $Y=62320
X799 1 2 955 923 177 ICV_6 $T=272320 95200 1 0 $X=272130 $Y=92240
X800 1 2 958 940 195 ICV_6 $T=286120 84320 0 0 $X=285930 $Y=84080
X801 1 2 973 943 174 ICV_6 $T=286120 106080 0 0 $X=285930 $Y=105840
X802 1 2 983 977 192 ICV_6 $T=300380 84320 1 0 $X=300190 $Y=81360
X803 1 2 1008 1005 188 ICV_6 $T=300380 100640 1 0 $X=300190 $Y=97680
X804 1 2 1037 1038 193 ICV_6 $T=314180 84320 0 0 $X=313990 $Y=84080
X805 1 2 1032 211 188 ICV_6 $T=314180 106080 0 0 $X=313990 $Y=105840
X806 1 2 1062 216 171 ICV_6 $T=328440 51680 1 0 $X=328250 $Y=48720
X807 1 2 1046 1053 170 ICV_6 $T=328440 100640 1 0 $X=328250 $Y=97680
X808 1 2 1058 1053 174 ICV_6 $T=328440 106080 1 0 $X=328250 $Y=103120
X809 1 2 1119 1101 194 ICV_6 $T=356500 51680 1 0 $X=356310 $Y=48720
X810 1 2 1141 1110 169 ICV_6 $T=370300 89760 0 0 $X=370110 $Y=89520
X811 1 2 1175 233 177 ICV_6 $T=384560 57120 1 0 $X=384370 $Y=54160
X812 1 2 1181 1149 192 ICV_6 $T=384560 68000 1 0 $X=384370 $Y=65040
X813 1 2 1177 1168 182 ICV_6 $T=384560 100640 1 0 $X=384370 $Y=97680
X814 1 2 1266 1270 182 ICV_6 $T=426420 95200 0 0 $X=426230 $Y=94960
X815 1 2 1294 252 180 ICV_6 $T=440680 57120 1 0 $X=440490 $Y=54160
X816 1 2 1296 1246 169 ICV_6 $T=440680 84320 1 0 $X=440490 $Y=81360
X817 1 2 1281 1246 180 ICV_6 $T=440680 89760 1 0 $X=440490 $Y=86800
X818 1 2 1293 1270 187 ICV_6 $T=440680 95200 1 0 $X=440490 $Y=92240
X819 1 2 1271 253 174 ICV_6 $T=440680 106080 1 0 $X=440490 $Y=103120
X820 1 2 1319 1312 275 ICV_6 $T=454480 57120 0 0 $X=454290 $Y=56880
X821 1 2 1324 1312 267 ICV_6 $T=454480 62560 0 0 $X=454290 $Y=62320
X822 1 2 1318 1312 276 ICV_6 $T=454480 68000 0 0 $X=454290 $Y=67760
X823 1 2 1328 271 269 ICV_6 $T=454480 111520 0 0 $X=454290 $Y=111280
X824 1 2 1351 1345 273 ICV_6 $T=468740 62560 1 0 $X=468550 $Y=59600
X825 1 2 1403 1399 304 ICV_6 $T=496800 84320 1 0 $X=496610 $Y=81360
X826 1 2 1437 1443 275 ICV_6 $T=510600 73440 0 0 $X=510410 $Y=73200
X827 1 2 1408 1386 288 ICV_6 $T=510600 78880 0 0 $X=510410 $Y=78640
X828 1 2 1441 1431 269 ICV_6 $T=510600 84320 0 0 $X=510410 $Y=84080
X829 1 2 1468 1431 267 ICV_6 $T=524860 84320 1 0 $X=524670 $Y=81360
X830 1 2 1488 1498 276 ICV_6 $T=538660 84320 0 0 $X=538470 $Y=84080
X831 1 2 1482 1461 277 ICV_6 $T=538660 106080 0 0 $X=538470 $Y=105840
X832 1 2 1570 1565 269 ICV_6 $T=580980 84320 1 0 $X=580790 $Y=81360
X833 1 2 1603 1600 276 ICV_6 $T=594780 106080 0 0 $X=594590 $Y=105840
X834 1 2 1629 1612 273 ICV_6 $T=609040 78880 1 0 $X=608850 $Y=75920
X835 1 2 1666 1657 273 ICV_6 $T=622840 78880 0 0 $X=622650 $Y=78640
X836 1 2 1653 1660 280 ICV_6 $T=622840 100640 0 0 $X=622650 $Y=100400
X837 1 2 1665 358 267 ICV_6 $T=622840 111520 0 0 $X=622650 $Y=111280
X838 1 2 1691 1688 269 ICV_6 $T=637100 111520 1 0 $X=636910 $Y=108560
X839 1 2 1724 1701 269 ICV_6 $T=650900 84320 0 0 $X=650710 $Y=84080
X840 1 2 390 391 307 ICV_6 $T=678960 111520 0 0 $X=678770 $Y=111280
X841 1 2 1837 1800 294 ICV_6 $T=707020 95200 0 0 $X=706830 $Y=94960
X993 1 2 449 6 2 458 1 sky130_fd_sc_hd__dfxtp_1 $T=9660 84320 0 0 $X=9470 $Y=84080
X994 1 2 3 6 2 459 1 sky130_fd_sc_hd__dfxtp_1 $T=9660 106080 0 0 $X=9470 $Y=105840
X995 1 2 453 4 2 463 1 sky130_fd_sc_hd__dfxtp_1 $T=10580 73440 0 0 $X=10390 $Y=73200
X996 1 2 454 4 2 465 1 sky130_fd_sc_hd__dfxtp_1 $T=10580 106080 1 0 $X=10390 $Y=103120
X997 1 2 454 8 2 450 1 sky130_fd_sc_hd__dfxtp_1 $T=12420 100640 1 0 $X=12230 $Y=97680
X998 1 2 453 25 2 487 1 sky130_fd_sc_hd__dfxtp_1 $T=25300 73440 0 0 $X=25110 $Y=73200
X999 1 2 452 26 2 488 1 sky130_fd_sc_hd__dfxtp_1 $T=25760 68000 0 0 $X=25570 $Y=67760
X1000 1 2 453 27 2 493 1 sky130_fd_sc_hd__dfxtp_1 $T=26220 78880 0 0 $X=26030 $Y=78640
X1001 1 2 454 26 2 504 1 sky130_fd_sc_hd__dfxtp_1 $T=27600 106080 1 0 $X=27410 $Y=103120
X1002 1 2 10 26 2 502 1 sky130_fd_sc_hd__dfxtp_1 $T=34960 57120 1 0 $X=34770 $Y=54160
X1003 1 2 509 4 2 518 1 sky130_fd_sc_hd__dfxtp_1 $T=38180 57120 0 0 $X=37990 $Y=56880
X1004 1 2 509 25 2 526 1 sky130_fd_sc_hd__dfxtp_1 $T=40020 73440 1 0 $X=39830 $Y=70480
X1005 1 2 510 8 2 547 1 sky130_fd_sc_hd__dfxtp_1 $T=50600 84320 0 0 $X=50410 $Y=84080
X1006 1 2 512 24 2 552 1 sky130_fd_sc_hd__dfxtp_1 $T=52440 100640 1 0 $X=52250 $Y=97680
X1007 1 2 512 8 2 554 1 sky130_fd_sc_hd__dfxtp_1 $T=52900 95200 0 0 $X=52710 $Y=94960
X1008 1 2 512 26 2 555 1 sky130_fd_sc_hd__dfxtp_1 $T=53360 89760 0 0 $X=53170 $Y=89520
X1009 1 2 45 26 2 564 1 sky130_fd_sc_hd__dfxtp_1 $T=57960 57120 1 0 $X=57770 $Y=54160
X1010 1 2 45 27 2 567 1 sky130_fd_sc_hd__dfxtp_1 $T=61640 51680 1 0 $X=61450 $Y=48720
X1011 1 2 591 5 2 604 1 sky130_fd_sc_hd__dfxtp_1 $T=80040 62560 1 0 $X=79850 $Y=59600
X1012 1 2 594 24 2 63 1 sky130_fd_sc_hd__dfxtp_1 $T=81880 51680 0 0 $X=81690 $Y=51440
X1013 1 2 594 25 2 611 1 sky130_fd_sc_hd__dfxtp_1 $T=83720 57120 1 0 $X=83530 $Y=54160
X1014 1 2 607 24 2 616 1 sky130_fd_sc_hd__dfxtp_1 $T=87860 84320 1 0 $X=87670 $Y=81360
X1015 1 2 610 24 2 70 1 sky130_fd_sc_hd__dfxtp_1 $T=94300 106080 1 0 $X=94110 $Y=103120
X1016 1 2 594 5 2 630 1 sky130_fd_sc_hd__dfxtp_1 $T=94760 57120 1 0 $X=94570 $Y=54160
X1017 1 2 649 25 2 661 1 sky130_fd_sc_hd__dfxtp_1 $T=109020 78880 0 0 $X=108830 $Y=78640
X1018 1 2 649 6 2 662 1 sky130_fd_sc_hd__dfxtp_1 $T=109480 95200 0 0 $X=109290 $Y=94960
X1019 1 2 72 6 2 674 1 sky130_fd_sc_hd__dfxtp_1 $T=115460 57120 1 0 $X=115270 $Y=54160
X1020 1 2 671 5 2 682 1 sky130_fd_sc_hd__dfxtp_1 $T=120980 73440 1 0 $X=120790 $Y=70480
X1021 1 2 675 8 2 707 1 sky130_fd_sc_hd__dfxtp_1 $T=136160 84320 1 0 $X=135970 $Y=81360
X1022 1 2 91 92 2 720 1 sky130_fd_sc_hd__dfxtp_1 $T=138460 111520 0 0 $X=138270 $Y=111280
X1023 1 2 708 4 2 724 1 sky130_fd_sc_hd__dfxtp_1 $T=140760 57120 1 0 $X=140570 $Y=54160
X1024 1 2 730 27 2 743 1 sky130_fd_sc_hd__dfxtp_1 $T=149040 100640 1 0 $X=148850 $Y=97680
X1025 1 2 97 25 2 745 1 sky130_fd_sc_hd__dfxtp_1 $T=151800 57120 1 0 $X=151610 $Y=54160
X1026 1 2 732 25 2 756 1 sky130_fd_sc_hd__dfxtp_1 $T=163300 84320 0 0 $X=163110 $Y=84080
X1027 1 2 741 5 2 787 1 sky130_fd_sc_hd__dfxtp_1 $T=173880 89760 1 0 $X=173690 $Y=86800
X1028 1 2 776 25 2 803 1 sky130_fd_sc_hd__dfxtp_1 $T=178020 111520 1 0 $X=177830 $Y=108560
X1029 1 2 775 26 2 805 1 sky130_fd_sc_hd__dfxtp_1 $T=179400 78880 1 0 $X=179210 $Y=75920
X1030 1 2 790 25 2 809 1 sky130_fd_sc_hd__dfxtp_1 $T=180780 62560 1 0 $X=180590 $Y=59600
X1031 1 2 790 24 2 830 1 sky130_fd_sc_hd__dfxtp_1 $T=194580 57120 0 0 $X=194390 $Y=56880
X1032 1 2 811 5 2 844 1 sky130_fd_sc_hd__dfxtp_1 $T=204700 68000 0 0 $X=204510 $Y=67760
X1033 1 2 837 6 2 849 1 sky130_fd_sc_hd__dfxtp_1 $T=207460 51680 1 0 $X=207270 $Y=48720
X1034 1 2 843 27 2 859 1 sky130_fd_sc_hd__dfxtp_1 $T=218960 62560 0 0 $X=218770 $Y=62320
X1035 1 2 847 26 2 873 1 sky130_fd_sc_hd__dfxtp_1 $T=224020 78880 1 0 $X=223830 $Y=75920
X1036 1 2 885 167 2 904 1 sky130_fd_sc_hd__dfxtp_1 $T=239660 73440 0 0 $X=239470 $Y=73200
X1037 1 2 883 186 2 950 1 sky130_fd_sc_hd__dfxtp_1 $T=261740 57120 1 0 $X=261550 $Y=54160
X1038 1 2 952 185 2 990 1 sky130_fd_sc_hd__dfxtp_1 $T=284280 68000 1 0 $X=284090 $Y=65040
X1039 1 2 984 185 2 986 1 sky130_fd_sc_hd__dfxtp_1 $T=287500 78880 1 0 $X=287310 $Y=75920
X1040 1 2 1009 184 2 1017 1 sky130_fd_sc_hd__dfxtp_1 $T=298080 57120 0 0 $X=297890 $Y=56880
X1041 1 2 207 158 2 1031 1 sky130_fd_sc_hd__dfxtp_1 $T=303600 106080 0 0 $X=303410 $Y=105840
X1042 1 2 1034 157 2 1052 1 sky130_fd_sc_hd__dfxtp_1 $T=324300 100640 0 0 $X=324110 $Y=100400
X1043 1 2 1049 185 2 1091 1 sky130_fd_sc_hd__dfxtp_1 $T=333500 62560 0 0 $X=333310 $Y=62320
X1044 1 2 1049 167 2 1092 1 sky130_fd_sc_hd__dfxtp_1 $T=333960 57120 0 0 $X=333770 $Y=56880
X1045 1 2 1078 181 2 1095 1 sky130_fd_sc_hd__dfxtp_1 $T=333960 100640 0 0 $X=333770 $Y=100400
X1046 1 2 1124 160 2 1158 1 sky130_fd_sc_hd__dfxtp_1 $T=367080 106080 1 0 $X=366890 $Y=103120
X1047 1 2 1162 158 2 1177 1 sky130_fd_sc_hd__dfxtp_1 $T=376280 95200 1 0 $X=376090 $Y=92240
X1048 1 2 1145 168 2 1182 1 sky130_fd_sc_hd__dfxtp_1 $T=379040 84320 0 0 $X=378850 $Y=84080
X1049 1 2 1162 165 2 1202 1 sky130_fd_sc_hd__dfxtp_1 $T=387320 95200 1 0 $X=387130 $Y=92240
X1050 1 2 1148 167 2 1183 1 sky130_fd_sc_hd__dfxtp_1 $T=387780 62560 0 0 $X=387590 $Y=62320
X1051 1 2 241 167 2 1233 1 sky130_fd_sc_hd__dfxtp_1 $T=404800 51680 1 0 $X=404610 $Y=48720
X1052 1 2 1256 184 2 1286 1 sky130_fd_sc_hd__dfxtp_1 $T=430560 68000 0 0 $X=430370 $Y=67760
X1053 1 2 1304 264 2 1329 1 sky130_fd_sc_hd__dfxtp_1 $T=448960 84320 1 0 $X=448770 $Y=81360
X1054 1 2 1292 264 2 1342 1 sky130_fd_sc_hd__dfxtp_1 $T=457700 73440 0 0 $X=457510 $Y=73200
X1055 1 2 1335 257 2 1343 1 sky130_fd_sc_hd__dfxtp_1 $T=460000 57120 1 0 $X=459810 $Y=54160
X1056 1 2 1335 262 2 1351 1 sky130_fd_sc_hd__dfxtp_1 $T=460000 62560 1 0 $X=459810 $Y=59600
X1057 1 2 1335 264 2 1354 1 sky130_fd_sc_hd__dfxtp_1 $T=460920 68000 1 0 $X=460730 $Y=65040
X1058 1 2 290 283 2 1380 1 sky130_fd_sc_hd__dfxtp_1 $T=475180 111520 0 0 $X=474990 $Y=111280
X1059 1 2 1381 301 2 1385 1 sky130_fd_sc_hd__dfxtp_1 $T=492660 78880 0 0 $X=492470 $Y=78640
X1060 1 2 1382 292 2 1415 1 sky130_fd_sc_hd__dfxtp_1 $T=494500 84320 0 0 $X=494310 $Y=84080
X1061 1 2 1420 258 2 1441 1 sky130_fd_sc_hd__dfxtp_1 $T=504620 89760 1 0 $X=504430 $Y=86800
X1062 1 2 1418 258 2 1449 1 sky130_fd_sc_hd__dfxtp_1 $T=510140 73440 1 0 $X=509950 $Y=70480
X1063 1 2 318 258 2 1463 1 sky130_fd_sc_hd__dfxtp_1 $T=513820 111520 0 0 $X=513630 $Y=111280
X1064 1 2 1418 262 2 1470 1 sky130_fd_sc_hd__dfxtp_1 $T=519340 62560 0 0 $X=519150 $Y=62320
X1065 1 2 1473 265 2 1499 1 sky130_fd_sc_hd__dfxtp_1 $T=530840 89760 0 0 $X=530650 $Y=89520
X1066 1 2 1473 257 2 1503 1 sky130_fd_sc_hd__dfxtp_1 $T=535900 89760 1 0 $X=535710 $Y=86800
X1067 1 2 331 292 2 1516 1 sky130_fd_sc_hd__dfxtp_1 $T=541880 51680 1 0 $X=541690 $Y=48720
X1068 1 2 1527 272 2 1552 1 sky130_fd_sc_hd__dfxtp_1 $T=557060 68000 0 0 $X=556870 $Y=67760
X1069 1 2 1506 259 2 1553 1 sky130_fd_sc_hd__dfxtp_1 $T=557060 95200 1 0 $X=556870 $Y=92240
X1070 1 2 338 262 2 1585 1 sky130_fd_sc_hd__dfxtp_1 $T=576840 106080 0 0 $X=576650 $Y=105840
X1071 1 2 1554 272 2 1586 1 sky130_fd_sc_hd__dfxtp_1 $T=579140 84320 0 0 $X=578950 $Y=84080
X1072 1 2 1569 266 2 1597 1 sky130_fd_sc_hd__dfxtp_1 $T=584200 73440 1 0 $X=584010 $Y=70480
X1073 1 2 1593 259 2 1599 1 sky130_fd_sc_hd__dfxtp_1 $T=587880 95200 1 0 $X=587690 $Y=92240
X1074 1 2 1592 262 2 1629 1 sky130_fd_sc_hd__dfxtp_1 $T=598920 73440 0 0 $X=598730 $Y=73200
X1075 1 2 1593 257 2 1633 1 sky130_fd_sc_hd__dfxtp_1 $T=598920 95200 1 0 $X=598730 $Y=92240
X1076 1 2 1640 272 2 1653 1 sky130_fd_sc_hd__dfxtp_1 $T=610420 100640 0 0 $X=610230 $Y=100400
X1077 1 2 361 259 2 1665 1 sky130_fd_sc_hd__dfxtp_1 $T=615480 111520 0 0 $X=615290 $Y=111280
X1078 1 2 1664 258 2 1691 1 sky130_fd_sc_hd__dfxtp_1 $T=626060 111520 1 0 $X=625870 $Y=108560
X1079 1 2 1694 265 2 1721 1 sky130_fd_sc_hd__dfxtp_1 $T=641700 62560 1 0 $X=641510 $Y=59600
X1080 1 2 1664 265 2 1725 1 sky130_fd_sc_hd__dfxtp_1 $T=645380 111520 1 0 $X=645190 $Y=108560
X1081 1 2 1753 292 2 1771 1 sky130_fd_sc_hd__dfxtp_1 $T=667920 78880 0 0 $X=667730 $Y=78640
X1082 1 2 1753 301 2 1779 1 sky130_fd_sc_hd__dfxtp_1 $T=670680 73440 0 0 $X=670490 $Y=73200
X1083 1 2 394 302 2 1809 1 sky130_fd_sc_hd__dfxtp_1 $T=686320 111520 0 0 $X=686130 $Y=111280
X1084 1 2 1817 292 2 1839 1 sky130_fd_sc_hd__dfxtp_1 $T=698740 100640 0 0 $X=698550 $Y=100400
X1085 1 2 1808 301 2 1843 1 sky130_fd_sc_hd__dfxtp_1 $T=711620 73440 1 0 $X=711430 $Y=70480
X1086 1 2 1867 301 2 1894 1 sky130_fd_sc_hd__dfxtp_1 $T=731860 73440 1 0 $X=731670 $Y=70480
X1087 1 2 499 9 33 10 25 499 ICV_13 $T=27140 51680 1 0 $X=26950 $Y=48720
X1088 1 2 516 14 30 3 24 516 ICV_13 $T=36340 111520 1 0 $X=36150 $Y=108560
X1089 1 2 518 525 20 509 24 519 ICV_13 $T=38640 62560 0 0 $X=38450 $Y=62320
X1090 1 2 521 525 18 509 6 521 ICV_13 $T=39100 68000 0 0 $X=38910 $Y=67760
X1091 1 2 530 533 18 512 6 530 ICV_13 $T=41860 89760 0 0 $X=41670 $Y=89520
X1092 1 2 537 40 34 35 27 537 ICV_13 $T=46000 51680 0 0 $X=45810 $Y=51440
X1093 1 2 542 525 17 509 5 542 ICV_13 $T=48300 62560 1 0 $X=48110 $Y=59600
X1094 1 2 553 534 34 39 27 553 ICV_13 $T=52440 111520 1 0 $X=52250 $Y=108560
X1095 1 2 568 47 18 540 6 568 ICV_13 $T=62560 73440 1 0 $X=62370 $Y=70480
X1096 1 2 571 573 20 560 4 571 ICV_13 $T=63940 78880 1 0 $X=63750 $Y=75920
X1097 1 2 579 563 18 566 5 578 ICV_13 $T=66700 95200 0 0 $X=66510 $Y=94960
X1098 1 2 577 54 32 566 24 561 ICV_13 $T=66700 100640 0 0 $X=66510 $Y=100400
X1099 1 2 583 573 11 566 26 585 ICV_13 $T=70380 89760 0 0 $X=70190 $Y=89520
X1100 1 2 593 573 32 560 26 593 ICV_13 $T=74060 78880 0 0 $X=73870 $Y=78640
X1101 1 2 595 573 17 560 5 595 ICV_13 $T=76360 78880 1 0 $X=76170 $Y=75920
X1102 1 2 596 54 11 51 8 596 ICV_13 $T=76360 106080 1 0 $X=76170 $Y=103120
X1103 1 2 599 54 17 51 5 599 ICV_13 $T=77740 111520 0 0 $X=77550 $Y=111280
X1104 1 2 608 64 20 591 8 587 ICV_13 $T=87400 62560 1 0 $X=87210 $Y=59600
X1105 1 2 628 64 18 594 6 628 ICV_13 $T=92000 51680 1 0 $X=91810 $Y=48720
X1106 1 2 635 615 11 610 26 639 ICV_13 $T=97520 89760 0 0 $X=97330 $Y=89520
X1107 1 2 651 644 18 633 6 651 ICV_13 $T=103500 100640 0 0 $X=103310 $Y=100400
X1108 1 2 695 692 33 671 25 695 ICV_13 $T=125120 62560 0 0 $X=124930 $Y=62320
X1109 1 2 699 700 33 678 25 699 ICV_13 $T=126040 89760 0 0 $X=125850 $Y=89520
X1110 1 2 709 86 33 679 25 709 ICV_13 $T=134320 100640 0 0 $X=134130 $Y=100400
X1111 1 2 728 725 30 708 6 726 ICV_13 $T=140760 73440 1 0 $X=140570 $Y=70480
X1112 1 2 750 748 34 732 26 749 ICV_13 $T=150420 78880 0 0 $X=150230 $Y=78640
X1113 1 2 756 748 33 741 24 735 ICV_13 $T=155020 89760 0 0 $X=154830 $Y=89520
X1114 1 2 757 760 34 738 4 763 ICV_13 $T=160540 62560 1 0 $X=160350 $Y=59600
X1115 1 2 767 102 17 97 5 767 ICV_13 $T=161000 51680 0 0 $X=160810 $Y=51440
X1116 1 2 771 748 17 732 24 769 ICV_13 $T=161920 78880 0 0 $X=161730 $Y=78640
X1117 1 2 753 760 11 112 5 795 ICV_13 $T=175720 57120 1 0 $X=175530 $Y=54160
X1118 1 2 833 817 18 802 6 833 ICV_13 $T=194580 89760 1 0 $X=194390 $Y=86800
X1119 1 2 835 810 20 790 4 835 ICV_13 $T=195960 57120 1 0 $X=195770 $Y=54160
X1120 1 2 842 826 34 811 27 842 ICV_13 $T=203780 73440 0 0 $X=203590 $Y=73200
X1121 1 2 858 857 18 847 4 854 ICV_13 $T=212060 84320 0 0 $X=211870 $Y=84080
X1122 1 2 863 139 32 149 26 875 ICV_13 $T=225400 51680 1 0 $X=225210 $Y=48720
X1123 1 2 884 857 11 847 8 884 ICV_13 $T=231380 78880 1 0 $X=231190 $Y=75920
X1124 1 2 908 890 171 885 164 887 ICV_13 $T=239660 68000 0 0 $X=239470 $Y=67760
X1125 1 2 934 892 193 883 183 934 ICV_13 $T=257140 62560 1 0 $X=256950 $Y=59600
X1126 1 2 939 176 194 161 185 939 ICV_13 $T=258980 51680 1 0 $X=258790 $Y=48720
X1127 1 2 941 940 171 928 185 937 ICV_13 $T=258980 73440 1 0 $X=258790 $Y=70480
X1128 1 2 942 923 180 909 167 942 ICV_13 $T=259440 89760 1 0 $X=259250 $Y=86800
X1129 1 2 960 940 177 928 168 960 ICV_13 $T=271400 68000 0 0 $X=271210 $Y=67760
X1130 1 2 961 967 192 952 184 961 ICV_13 $T=271860 57120 0 0 $X=271670 $Y=56880
X1131 1 2 963 967 169 952 164 963 ICV_13 $T=272780 62560 1 0 $X=272590 $Y=59600
X1132 1 2 964 967 171 952 166 964 ICV_13 $T=272780 68000 1 0 $X=272590 $Y=65040
X1133 1 2 965 940 180 928 167 965 ICV_13 $T=272780 73440 1 0 $X=272590 $Y=70480
X1134 1 2 972 923 171 909 166 972 ICV_13 $T=274620 84320 0 0 $X=274430 $Y=84080
X1135 1 2 981 977 177 959 168 981 ICV_13 $T=277380 89760 1 0 $X=277190 $Y=86800
X1136 1 2 962 940 169 959 184 983 ICV_13 $T=278300 84320 1 0 $X=278110 $Y=81360
X1137 1 2 997 988 195 984 183 995 ICV_13 $T=286580 68000 0 0 $X=286390 $Y=67760
X1138 1 2 999 1005 187 989 175 999 ICV_13 $T=288880 100640 1 0 $X=288690 $Y=97680
X1139 1 2 1003 977 180 959 166 1007 ICV_13 $T=290720 84320 0 0 $X=290530 $Y=84080
X1140 1 2 1013 212 193 208 166 213 ICV_13 $T=300840 51680 0 0 $X=300650 $Y=51440
X1141 1 2 1026 1005 174 989 160 1026 ICV_13 $T=300840 100640 0 0 $X=300650 $Y=100400
X1142 1 2 1041 1038 169 1020 164 1041 ICV_13 $T=309580 89760 1 0 $X=309390 $Y=86800
X1143 1 2 1055 217 189 215 181 1055 ICV_13 $T=316020 111520 0 0 $X=315830 $Y=111280
X1144 1 2 1069 1071 177 1049 168 1069 ICV_13 $T=322000 62560 0 0 $X=321810 $Y=62320
X1145 1 2 1067 1038 180 1020 186 1072 ICV_13 $T=323840 89760 0 0 $X=323650 $Y=89520
X1146 1 2 1065 1071 169 214 167 1075 ICV_13 $T=328900 51680 0 0 $X=328710 $Y=51440
X1147 1 2 1082 1039 194 1033 185 1082 ICV_13 $T=328900 78880 1 0 $X=328710 $Y=75920
X1148 1 2 1083 1038 194 1020 185 1083 ICV_13 $T=328900 89760 1 0 $X=328710 $Y=86800
X1149 1 2 1085 1074 191 215 160 218 ICV_13 $T=328900 111520 1 0 $X=328710 $Y=108560
X1150 1 2 1092 1071 180 1049 186 1093 ICV_13 $T=333960 62560 1 0 $X=333770 $Y=59600
X1151 1 2 1104 222 187 220 175 1104 ICV_13 $T=340400 111520 1 0 $X=340210 $Y=108560
X1152 1 2 1136 1100 177 1089 168 1136 ICV_13 $T=356960 78880 1 0 $X=356770 $Y=75920
X1153 1 2 1139 1133 178 220 165 229 ICV_13 $T=358340 111520 0 0 $X=358150 $Y=111280
X1154 1 2 1153 1110 177 1096 168 1153 ICV_13 $T=364320 89760 1 0 $X=364130 $Y=86800
X1155 1 2 1170 232 182 231 158 1170 ICV_13 $T=371680 111520 1 0 $X=371490 $Y=108560
X1156 1 2 1189 232 187 231 175 1189 ICV_13 $T=384100 106080 0 0 $X=383910 $Y=105840
X1157 1 2 1194 233 192 1159 167 1197 ICV_13 $T=386400 51680 0 0 $X=386210 $Y=51440
X1158 1 2 1208 233 194 1159 185 1208 ICV_13 $T=393300 51680 1 0 $X=393110 $Y=48720
X1159 1 2 1211 1210 177 1188 168 1211 ICV_13 $T=395600 68000 1 0 $X=395410 $Y=65040
X1160 1 2 242 243 178 1205 173 1218 ICV_13 $T=397440 111520 1 0 $X=397250 $Y=108560
X1161 1 2 1219 1199 171 1180 166 1219 ICV_13 $T=397900 95200 1 0 $X=397710 $Y=92240
X1162 1 2 1222 1228 180 1204 167 1222 ICV_13 $T=398820 62560 0 0 $X=398630 $Y=62320
X1163 1 2 1245 1212 187 1205 156 1243 ICV_13 $T=408940 95200 0 0 $X=408750 $Y=94960
X1164 1 2 1252 1228 171 1204 164 1247 ICV_13 $T=411700 62560 0 0 $X=411510 $Y=62320
X1165 1 2 1269 1270 174 1250 160 1269 ICV_13 $T=420440 100640 1 0 $X=420250 $Y=97680
X1166 1 2 1278 1261 171 1242 166 1278 ICV_13 $T=426880 78880 0 0 $X=426690 $Y=78640
X1167 1 2 1268 1246 177 1239 167 1281 ICV_13 $T=427800 89760 1 0 $X=427610 $Y=86800
X1168 1 2 1282 252 193 249 183 1282 ICV_13 $T=428720 51680 1 0 $X=428530 $Y=48720
X1169 1 2 1295 1270 189 1250 181 1295 ICV_13 $T=434240 100640 0 0 $X=434050 $Y=100400
X1170 1 2 1288 1246 195 1239 164 1296 ICV_13 $T=434700 84320 0 0 $X=434510 $Y=84080
X1171 1 2 1300 1262 194 1256 185 1300 ICV_13 $T=437920 68000 0 0 $X=437730 $Y=67760
X1172 1 2 1316 1312 273 1301 262 1316 ICV_13 $T=445740 62560 1 0 $X=445550 $Y=59600
X1173 1 2 1325 1311 273 1292 262 1325 ICV_13 $T=448500 73440 1 0 $X=448310 $Y=70480
X1174 1 2 278 252 195 249 185 1317 ICV_13 $T=452640 51680 1 0 $X=452450 $Y=48720
X1175 1 2 1361 1345 280 1335 266 1359 ICV_13 $T=466900 68000 0 0 $X=466710 $Y=67760
X1176 1 2 1360 1331 269 1305 258 1360 ICV_13 $T=466900 89760 0 0 $X=466710 $Y=89520
X1177 1 2 1365 1315 269 1306 272 1363 ICV_13 $T=467820 106080 0 0 $X=467630 $Y=105840
X1178 1 2 1398 1399 307 1382 299 1398 ICV_13 $T=483920 95200 1 0 $X=483730 $Y=92240
X1179 1 2 1397 1357 303 282 299 1402 ICV_13 $T=484380 57120 0 0 $X=484190 $Y=56880
X1180 1 2 1422 1428 294 1409 283 1422 ICV_13 $T=497260 62560 0 0 $X=497070 $Y=62320
X1181 1 2 1424 1399 309 1382 302 1424 ICV_13 $T=497260 95200 1 0 $X=497070 $Y=92240
X1182 1 2 1438 1431 268 1420 266 1429 ICV_13 $T=504620 78880 1 0 $X=504430 $Y=75920
X1183 1 2 1450 1446 300 1436 283 1456 ICV_13 $T=511980 95200 0 0 $X=511790 $Y=94960
X1184 1 2 1448 1428 304 1418 257 1459 ICV_13 $T=512900 68000 1 0 $X=512710 $Y=65040
X1185 1 2 1475 1461 275 318 265 1475 ICV_13 $T=522560 106080 0 0 $X=522370 $Y=105840
X1186 1 2 1476 1446 288 1436 301 1480 ICV_13 $T=525320 100640 1 0 $X=525130 $Y=97680
X1187 1 2 1493 1498 269 1473 258 1493 ICV_13 $T=529460 84320 1 0 $X=529270 $Y=81360
X1188 1 2 1495 1498 267 1473 259 1495 ICV_13 $T=529920 95200 1 0 $X=529730 $Y=92240
X1189 1 2 1496 1461 267 318 259 1496 ICV_13 $T=529920 106080 1 0 $X=529730 $Y=103120
X1190 1 2 1515 1513 269 1500 258 1515 ICV_13 $T=541420 106080 1 0 $X=541230 $Y=103120
X1191 1 2 1532 1513 276 1500 257 1531 ICV_13 $T=551080 106080 0 0 $X=550890 $Y=105840
X1192 1 2 1533 334 304 331 301 1533 ICV_13 $T=553380 51680 1 0 $X=553190 $Y=48720
X1193 1 2 1536 1512 273 1491 262 1536 ICV_13 $T=553380 78880 1 0 $X=553190 $Y=75920
X1194 1 2 335 333 307 329 301 1539 ICV_13 $T=553380 111520 0 0 $X=553190 $Y=111280
X1195 1 2 1540 1512 280 1491 272 1540 ICV_13 $T=553840 73440 0 0 $X=553650 $Y=73200
X1196 1 2 1613 1612 276 1592 265 1608 ICV_13 $T=587420 78880 1 0 $X=587230 $Y=75920
X1197 1 2 1624 1601 269 1593 258 1624 ICV_13 $T=597080 100640 1 0 $X=596890 $Y=97680
X1198 1 2 1652 1657 275 1637 265 1652 ICV_13 $T=609960 78880 0 0 $X=609770 $Y=78640
X1199 1 2 1656 1660 275 1640 265 1656 ICV_13 $T=610880 95200 0 0 $X=610690 $Y=94960
X1200 1 2 1672 365 309 364 305 1677 ICV_13 $T=623300 51680 0 0 $X=623110 $Y=51440
X1201 1 2 1683 1660 273 1640 266 1684 ICV_13 $T=623300 95200 0 0 $X=623110 $Y=94960
X1202 1 2 1667 1674 273 1646 265 1671 ICV_13 $T=624680 62560 1 0 $X=624490 $Y=59600
X1203 1 2 1707 1709 267 1694 272 1702 ICV_13 $T=634800 57120 0 0 $X=634610 $Y=56880
X1204 1 2 1703 1709 276 1694 264 1703 ICV_13 $T=634800 62560 0 0 $X=634610 $Y=62320
X1205 1 2 1704 1708 276 1692 264 1704 ICV_13 $T=634800 73440 0 0 $X=634610 $Y=73200
X1206 1 2 1705 1701 267 1690 259 1705 ICV_13 $T=634800 78880 0 0 $X=634610 $Y=78640
X1207 1 2 1710 1697 276 1695 272 1706 ICV_13 $T=635260 100640 0 0 $X=635070 $Y=100400
X1208 1 2 1715 1701 277 1692 266 1714 ICV_13 $T=637560 78880 1 0 $X=637370 $Y=75920
X1209 1 2 1698 1688 280 377 259 378 ICV_13 $T=638480 111520 0 0 $X=638290 $Y=111280
X1210 1 2 1719 379 300 376 301 1718 ICV_13 $T=639400 51680 0 0 $X=639210 $Y=51440
X1211 1 2 1732 1709 273 1694 262 1732 ICV_13 $T=649060 62560 1 0 $X=648870 $Y=59600
X1212 1 2 1739 1708 273 1692 262 1739 ICV_13 $T=651360 68000 0 0 $X=651170 $Y=67760
X1213 1 2 1751 1746 307 1731 299 1751 ICV_13 $T=655500 84320 0 0 $X=655310 $Y=84080
X1214 1 2 1763 1748 309 1753 302 1763 ICV_13 $T=665620 68000 1 0 $X=665430 $Y=65040
X1215 1 2 1758 1748 307 1753 305 1764 ICV_13 $T=665620 78880 1 0 $X=665430 $Y=75920
X1216 1 2 1767 386 300 1754 292 1767 ICV_13 $T=665620 106080 1 0 $X=665430 $Y=103120
X1217 1 2 1768 386 294 1754 283 1768 ICV_13 $T=665620 111520 1 0 $X=665430 $Y=108560
X1218 1 2 1770 1746 303 1731 297 1770 ICV_13 $T=666080 89760 0 0 $X=665890 $Y=89520
X1219 1 2 1785 386 296 1754 287 1785 ICV_13 $T=677120 106080 1 0 $X=676930 $Y=103120
X1220 1 2 1784 1800 300 1754 301 1789 ICV_13 $T=679420 100640 0 0 $X=679230 $Y=100400
X1221 1 2 1790 386 288 1754 305 1790 ICV_13 $T=679420 106080 0 0 $X=679230 $Y=105840
X1222 1 2 1795 1800 309 1776 302 1795 ICV_13 $T=680340 95200 0 0 $X=680150 $Y=94960
X1223 1 2 1797 1798 296 1782 287 1797 ICV_13 $T=680800 62560 1 0 $X=680610 $Y=59600
X1224 1 2 1801 1800 303 1776 301 1799 ICV_13 $T=680800 95200 1 0 $X=680610 $Y=92240
X1225 1 2 1810 1798 303 1782 297 1810 ICV_13 $T=687240 62560 0 0 $X=687050 $Y=62320
X1226 1 2 1818 1800 307 1776 305 1822 ICV_13 $T=693680 100640 1 0 $X=693490 $Y=97680
X1227 1 2 1809 400 309 394 283 399 ICV_13 $T=693680 111520 0 0 $X=693490 $Y=111280
X1228 1 2 1830 1824 307 1807 301 1832 ICV_13 $T=696900 51680 1 0 $X=696710 $Y=48720
X1229 1 2 1846 1824 296 1807 287 1846 ICV_13 $T=706100 62560 1 0 $X=705910 $Y=59600
X1230 1 2 1850 1816 309 1808 302 1850 ICV_13 $T=707480 68000 0 0 $X=707290 $Y=67760
X1231 1 2 1857 1838 288 1817 305 1857 ICV_13 $T=708860 111520 1 0 $X=708670 $Y=108560
X1232 1 2 1881 1883 300 1866 297 1875 ICV_13 $T=719900 62560 0 0 $X=719710 $Y=62320
X1233 1 2 1875 1883 303 1867 297 1888 ICV_13 $T=721740 68000 1 0 $X=721550 $Y=65040
X1234 1 2 1889 1882 303 1868 305 1891 ICV_13 $T=723120 89760 0 0 $X=722930 $Y=89520
X1235 1 2 1903 1882 307 1867 299 1880 ICV_13 $T=731400 78880 1 0 $X=731210 $Y=75920
X1236 1 2 591 27 624 624 586 34 ICV_14 $T=90160 68000 0 0 $X=89970 $Y=67760
X1237 1 2 633 4 652 652 644 20 ICV_14 $T=103040 106080 0 0 $X=102850 $Y=105840
X1238 1 2 85 25 722 722 90 33 ICV_14 $T=138920 51680 1 0 $X=138730 $Y=48720
X1239 1 2 811 25 822 822 826 33 ICV_14 $T=188600 73440 1 0 $X=188410 $Y=70480
X1240 1 2 811 4 845 845 826 20 ICV_14 $T=203780 78880 1 0 $X=203590 $Y=75920
X1241 1 2 837 25 136 849 139 18 ICV_14 $T=206540 51680 0 0 $X=206350 $Y=51440
X1242 1 2 881 165 910 910 891 188 ICV_14 $T=243800 95200 0 0 $X=243610 $Y=94960
X1243 1 2 928 166 941 920 886 194 ICV_14 $T=258520 73440 0 0 $X=258330 $Y=73200
X1244 1 2 952 186 991 991 967 195 ICV_14 $T=284280 62560 1 0 $X=284090 $Y=59600
X1245 1 2 984 166 1002 1022 988 192 ICV_14 $T=298080 78880 0 0 $X=297890 $Y=78640
X1246 1 2 1020 184 1035 1035 1038 192 ICV_14 $T=304980 84320 1 0 $X=304790 $Y=81360
X1247 1 2 1096 167 1108 1108 1110 180 ICV_14 $T=340400 89760 1 0 $X=340210 $Y=86800
X1248 1 2 1096 164 1141 1137 1110 193 ICV_14 $T=356960 84320 0 0 $X=356770 $Y=84080
X1249 1 2 1102 184 1142 1142 1101 192 ICV_14 $T=357420 57120 0 0 $X=357230 $Y=56880
X1250 1 2 1102 186 1143 1134 1101 171 ICV_14 $T=357420 62560 0 0 $X=357230 $Y=62320
X1251 1 2 231 156 1196 1196 232 170 ICV_14 $T=385020 111520 1 0 $X=384830 $Y=108560
X1252 1 2 1205 158 1216 1216 1212 182 ICV_14 $T=396520 100640 1 0 $X=396330 $Y=97680
X1253 1 2 1306 262 1332 1332 1315 273 ICV_14 $T=448500 100640 1 0 $X=448310 $Y=97680
X1254 1 2 1301 258 1384 1384 1312 269 ICV_14 $T=477480 68000 1 0 $X=477290 $Y=65040
X1255 1 2 1409 297 1426 1427 1428 309 ICV_14 $T=497260 57120 0 0 $X=497070 $Y=56880
X1256 1 2 1409 287 1454 1457 1428 307 ICV_14 $T=511060 57120 0 0 $X=510870 $Y=56880
X1257 1 2 1420 264 1466 1466 1431 276 ICV_14 $T=515200 84320 0 0 $X=515010 $Y=84080
X1258 1 2 1527 266 1562 1564 1546 276 ICV_14 $T=564880 73440 1 0 $X=564690 $Y=70480
X1259 1 2 1640 262 1683 1686 1660 276 ICV_14 $T=622380 95200 1 0 $X=622190 $Y=92240
X1260 1 2 1782 301 1794 1794 1798 304 ICV_14 $T=679420 73440 0 0 $X=679230 $Y=73200
X1261 1 2 1819 292 1853 1853 1829 300 ICV_14 $T=707480 89760 1 0 $X=707290 $Y=86800
X1262 1 2 1807 297 1856 1856 1824 303 ICV_14 $T=707940 57120 1 0 $X=707750 $Y=54160
X1263 1 2 1817 302 1862 1862 1838 309 ICV_14 $T=708400 106080 1 0 $X=708210 $Y=103120
X1264 1 2 1867 305 1870 1885 1869 300 ICV_14 $T=719440 73440 0 0 $X=719250 $Y=73200
X1265 1 2 1865 301 1872 1904 1874 294 ICV_14 $T=730480 100640 1 0 $X=730290 $Y=97680
X1266 1 2 452 8 467 460 476 20 ICV_16 $T=10580 62560 0 0 $X=10390 $Y=62320
X1267 1 2 449 26 500 500 473 32 ICV_16 $T=26680 89760 1 0 $X=26490 $Y=86800
X1268 1 2 449 25 505 495 473 34 ICV_16 $T=27600 95200 1 0 $X=27410 $Y=92240
X1269 1 2 35 6 543 543 40 18 ICV_16 $T=48300 51680 1 0 $X=48110 $Y=48720
X1270 1 2 566 25 597 597 563 33 ICV_16 $T=76360 100640 1 0 $X=76170 $Y=97680
X1271 1 2 72 8 74 634 64 32 ICV_16 $T=103040 51680 0 0 $X=102850 $Y=51440
X1272 1 2 679 4 702 703 86 11 ICV_16 $T=126500 111520 0 0 $X=126310 $Y=111280
X1273 1 2 708 26 727 727 725 32 ICV_16 $T=140760 62560 1 0 $X=140570 $Y=59600
X1274 1 2 775 4 793 793 792 20 ICV_16 $T=174340 78880 0 0 $X=174150 $Y=78640
X1275 1 2 775 8 794 794 792 11 ICV_16 $T=174340 84320 1 0 $X=174150 $Y=81360
X1276 1 2 775 5 799 799 792 17 ICV_16 $T=175720 68000 0 0 $X=175530 $Y=67760
X1277 1 2 775 25 804 804 792 33 ICV_16 $T=178020 73440 0 0 $X=177830 $Y=73200
X1278 1 2 802 4 813 780 734 11 ICV_16 $T=184000 89760 0 0 $X=183810 $Y=89520
X1279 1 2 811 8 824 824 826 11 ICV_16 $T=189980 73440 0 0 $X=189790 $Y=73200
X1280 1 2 843 25 860 860 856 33 ICV_16 $T=214360 68000 0 0 $X=214170 $Y=67760
X1281 1 2 843 4 877 880 856 32 ICV_16 $T=224940 62560 1 0 $X=224750 $Y=59600
X1282 1 2 881 160 895 894 891 178 ICV_16 $T=235060 100640 0 0 $X=234870 $Y=100400
X1283 1 2 871 164 896 901 886 180 ICV_16 $T=235980 84320 0 0 $X=235790 $Y=84080
X1284 1 2 161 168 903 897 176 171 ICV_16 $T=237820 51680 0 0 $X=237630 $Y=51440
X1285 1 2 952 183 968 968 967 193 ICV_16 $T=272780 62560 0 0 $X=272590 $Y=62320
X1286 1 2 196 158 969 969 198 182 ICV_16 $T=272780 106080 0 0 $X=272590 $Y=105840
X1287 1 2 196 156 970 970 198 170 ICV_16 $T=272780 111520 1 0 $X=272590 $Y=108560
X1288 1 2 984 164 996 996 988 169 ICV_16 $T=286580 73440 0 0 $X=286390 $Y=73200
X1289 1 2 984 167 1015 1021 988 177 ICV_16 $T=298540 73440 0 0 $X=298350 $Y=73200
X1290 1 2 989 157 1027 1027 1005 178 ICV_16 $T=300840 106080 1 0 $X=300650 $Y=103120
X1291 1 2 215 165 1054 1054 217 188 ICV_16 $T=315100 111520 1 0 $X=314910 $Y=108560
X1292 1 2 1049 183 1090 1090 1071 193 ICV_16 $T=332580 68000 1 0 $X=332390 $Y=65040
X1293 1 2 219 168 1099 1099 221 177 ICV_16 $T=337180 57120 1 0 $X=336990 $Y=54160
X1294 1 2 1096 186 1111 1111 1110 195 ICV_16 $T=342700 89760 0 0 $X=342510 $Y=89520
X1295 1 2 1145 186 1161 1164 1157 180 ICV_16 $T=370760 84320 1 0 $X=370570 $Y=81360
X1296 1 2 1204 184 1220 1220 1228 192 ICV_16 $T=397900 62560 1 0 $X=397710 $Y=59600
X1297 1 2 1180 186 1227 1214 1199 169 ICV_16 $T=398820 84320 0 0 $X=398630 $Y=84080
X1298 1 2 1188 184 1236 1236 1210 192 ICV_16 $T=405260 73440 0 0 $X=405070 $Y=73200
X1299 1 2 241 164 1255 1255 246 169 ICV_16 $T=413080 51680 1 0 $X=412890 $Y=48720
X1300 1 2 1242 183 1259 1259 1261 193 ICV_16 $T=415380 78880 1 0 $X=415190 $Y=75920
X1301 1 2 1242 167 1280 1280 1261 180 ICV_16 $T=427340 73440 1 0 $X=427150 $Y=70480
X1302 1 2 1248 181 1299 1299 253 189 ICV_16 $T=435160 106080 0 0 $X=434970 $Y=105840
X1303 1 2 1292 257 1307 1308 1311 267 ICV_16 $T=440220 73440 0 0 $X=440030 $Y=73200
X1304 1 2 1292 266 1368 1368 1311 277 ICV_16 $T=469200 78880 1 0 $X=469010 $Y=75920
X1305 1 2 1381 283 1391 1391 1386 294 ICV_16 $T=482540 78880 1 0 $X=482350 $Y=75920
X1306 1 2 282 297 1397 1393 1312 280 ICV_16 $T=483460 62560 1 0 $X=483270 $Y=59600
X1307 1 2 1409 292 1425 1425 1428 300 ICV_16 $T=497260 62560 1 0 $X=497070 $Y=59600
X1308 1 2 1436 287 1478 1478 1446 296 ICV_16 $T=523480 95200 0 0 $X=523290 $Y=94960
X1309 1 2 1500 259 1514 1514 1513 267 ICV_16 $T=540500 100640 0 0 $X=540310 $Y=100400
X1310 1 2 329 287 1541 1541 333 296 ICV_16 $T=553380 111520 1 0 $X=553190 $Y=108560
X1311 1 2 1591 258 1619 1619 1600 269 ICV_16 $T=591100 111520 1 0 $X=590910 $Y=108560
X1312 1 2 1640 257 1654 1654 1660 268 ICV_16 $T=610420 89760 0 0 $X=610230 $Y=89520
X1313 1 2 1640 264 1686 1684 1660 277 ICV_16 $T=623300 89760 0 0 $X=623110 $Y=89520
X1314 1 2 1692 265 1734 1734 1708 275 ICV_16 $T=649060 78880 1 0 $X=648870 $Y=75920
X1315 1 2 1753 297 1769 1769 1748 303 ICV_16 $T=665620 73440 1 0 $X=665430 $Y=70480
X1316 1 2 1753 287 1747 1765 1746 296 ICV_16 $T=665620 84320 1 0 $X=665430 $Y=81360
X1317 1 2 1807 302 1820 1820 1824 309 ICV_16 $T=692760 51680 0 0 $X=692570 $Y=51440
X1318 1 2 1817 287 1852 1852 1838 296 ICV_16 $T=707480 111520 0 0 $X=707290 $Y=111280
X1319 1 2 1865 302 1873 1873 1874 309 ICV_16 $T=718060 95200 0 0 $X=717870 $Y=94960
X1320 1 2 1868 292 1886 1886 1882 300 ICV_16 $T=720820 78880 0 0 $X=720630 $Y=78640
X1321 1 2 540 5 562 564 53 32 ICV_17 $T=59800 62560 1 0 $X=59610 $Y=59600
X1322 1 2 594 27 626 626 64 34 ICV_17 $T=90160 51680 0 0 $X=89970 $Y=51440
X1323 1 2 610 8 627 623 68 33 ICV_17 $T=90160 106080 0 0 $X=89970 $Y=105840
X1324 1 2 633 8 648 650 644 33 ICV_17 $T=99820 111520 0 0 $X=99630 $Y=111280
X1325 1 2 649 24 664 661 643 33 ICV_17 $T=108560 84320 1 0 $X=108370 $Y=81360
X1326 1 2 811 24 823 823 826 30 ICV_17 $T=188600 68000 1 0 $X=188410 $Y=65040
X1327 1 2 837 5 870 870 139 17 ICV_17 $T=218960 57120 1 0 $X=218770 $Y=54160
X1328 1 2 881 181 912 913 891 191 ICV_17 $T=244720 106080 1 0 $X=244530 $Y=103120
X1329 1 2 928 183 944 944 940 193 ICV_17 $T=258520 68000 0 0 $X=258330 $Y=67760
X1330 1 2 926 158 945 945 943 182 ICV_17 $T=258520 95200 0 0 $X=258330 $Y=94960
X1331 1 2 926 156 946 935 943 191 ICV_17 $T=259440 100640 1 0 $X=259250 $Y=97680
X1332 1 2 928 164 962 966 940 192 ICV_17 $T=270940 73440 0 0 $X=270750 $Y=73200
X1333 1 2 989 156 1025 1024 1005 182 ICV_17 $T=299460 95200 0 0 $X=299270 $Y=94960
X1334 1 2 1009 186 1040 1042 1018 169 ICV_17 $T=308200 62560 1 0 $X=308010 $Y=59600
X1335 1 2 1009 164 1042 1047 1018 171 ICV_17 $T=309580 68000 1 0 $X=309390 $Y=65040
X1336 1 2 219 183 1113 1113 221 193 ICV_17 $T=342700 51680 0 0 $X=342510 $Y=51440
X1337 1 2 1078 158 1114 1114 1074 182 ICV_17 $T=342700 95200 0 0 $X=342510 $Y=94960
X1338 1 2 1159 166 1198 1198 233 171 ICV_17 $T=385020 62560 1 0 $X=384830 $Y=59600
X1339 1 2 1205 157 1238 1243 1212 170 ICV_17 $T=406180 100640 0 0 $X=405990 $Y=100400
X1340 1 2 1256 168 1273 1274 1262 180 ICV_17 $T=420440 62560 1 0 $X=420250 $Y=59600
X1341 1 2 1304 258 1376 1376 1333 269 ICV_17 $T=471500 84320 1 0 $X=471310 $Y=81360
X1342 1 2 282 302 1401 1401 1357 309 ICV_17 $T=483000 51680 0 0 $X=482810 $Y=51440
X1343 1 2 1420 262 1467 1467 1431 273 ICV_17 $T=515200 78880 0 0 $X=515010 $Y=78640
X1344 1 2 1491 259 1505 1472 1443 277 ICV_17 $T=534980 73440 1 0 $X=534790 $Y=70480
X1345 1 2 331 283 1530 1530 334 294 ICV_17 $T=549700 51680 0 0 $X=549510 $Y=51440
X1346 1 2 1544 264 1557 1557 1551 276 ICV_17 $T=560740 106080 1 0 $X=560550 $Y=103120
X1347 1 2 1527 259 1568 1568 1546 267 ICV_17 $T=566720 62560 1 0 $X=566530 $Y=59600
X1348 1 2 1616 259 1643 1643 1625 267 ICV_17 $T=604440 57120 0 0 $X=604250 $Y=56880
X1349 1 2 1640 259 1655 1655 1660 267 ICV_17 $T=609500 95200 1 0 $X=609310 $Y=92240
X1350 1 2 1692 257 1735 1735 1708 268 ICV_17 $T=648600 73440 1 0 $X=648410 $Y=70480
X1351 1 2 1754 302 1760 1760 386 309 ICV_17 $T=662400 106080 0 0 $X=662210 $Y=105840
X1352 1 2 1781 302 1811 1814 1816 296 ICV_17 $T=686780 78880 0 0 $X=686590 $Y=78640
X1353 1 2 1781 297 1812 1812 1774 303 ICV_17 $T=687240 89760 0 0 $X=687050 $Y=89520
X1354 1 2 1807 292 1855 1855 1824 300 ICV_17 $T=707480 51680 0 0 $X=707290 $Y=51440
X1355 1 2 1866 305 1877 1884 1883 309 ICV_17 $T=718980 57120 0 0 $X=718790 $Y=56880
X1356 1 2 1867 302 1878 1878 1869 309 ICV_17 $T=718980 68000 0 0 $X=718790 $Y=67760
X1357 1 2 403 305 1845 407 397 309 ICV_17 $T=719440 111520 0 0 $X=719250 $Y=111280
X1374 1 2 452 25 489 489 476 33 ICV_19 $T=24380 62560 1 0 $X=24190 $Y=59600
X1375 1 2 560 6 589 589 573 18 ICV_19 $T=69920 84320 0 0 $X=69730 $Y=84080
X1376 1 2 671 24 691 691 692 30 ICV_19 $T=122360 68000 0 0 $X=122170 $Y=67760
X1377 1 2 708 25 731 731 725 33 ICV_19 $T=140760 68000 1 0 $X=140570 $Y=65040
X1378 1 2 112 25 798 798 114 33 ICV_19 $T=174340 51680 0 0 $X=174150 $Y=51440
X1379 1 2 811 6 821 821 826 18 ICV_19 $T=187680 68000 0 0 $X=187490 $Y=67760
X1380 1 2 1162 173 1201 1178 1168 189 ICV_19 $T=385020 106080 1 0 $X=384830 $Y=103120
X1381 1 2 1242 186 1284 1284 1261 195 ICV_19 $T=426880 73440 0 0 $X=426690 $Y=73200
X1382 1 2 1306 266 1370 1370 1315 277 ICV_19 $T=469200 100640 1 0 $X=469010 $Y=97680
X1383 1 2 282 301 1400 1400 1357 304 ICV_19 $T=482540 51680 1 0 $X=482350 $Y=48720
X1384 1 2 1471 262 1484 1484 1479 273 ICV_19 $T=525320 62560 1 0 $X=525130 $Y=59600
X1385 1 2 1471 257 1501 1507 1479 276 ICV_19 $T=539120 62560 0 0 $X=538930 $Y=62320
X1386 1 2 1527 262 1542 1542 1546 273 ICV_19 $T=553380 62560 1 0 $X=553190 $Y=59600
X1387 1 2 1646 258 1669 1671 1674 275 ICV_19 $T=616860 68000 1 0 $X=616670 $Y=65040
X1388 1 2 1690 257 1720 1729 1701 273 ICV_19 $T=644920 84320 1 0 $X=644730 $Y=81360
X1389 1 2 1782 305 1786 1786 1798 288 ICV_19 $T=677580 73440 1 0 $X=677390 $Y=70480
X1390 1 2 1819 287 1858 1858 1829 296 ICV_19 $T=707480 78880 0 0 $X=707290 $Y=78640
X1391 1 2 452 6 466 ICV_20 $T=10580 62560 1 0 $X=10390 $Y=59600
X1392 1 2 453 6 468 ICV_20 $T=10580 78880 0 0 $X=10390 $Y=78640
X1393 1 2 454 6 469 ICV_20 $T=10580 100640 0 0 $X=10390 $Y=100400
X1394 1 2 453 24 486 ICV_20 $T=24380 78880 1 0 $X=24190 $Y=75920
X1395 1 2 452 27 490 ICV_20 $T=25760 62560 0 0 $X=25570 $Y=62320
X1396 1 2 453 26 492 ICV_20 $T=25760 84320 1 0 $X=25570 $Y=81360
X1397 1 2 449 24 494 ICV_20 $T=25760 84320 0 0 $X=25570 $Y=84080
X1398 1 2 449 27 495 ICV_20 $T=25760 89760 0 0 $X=25570 $Y=89520
X1399 1 2 3 27 498 ICV_20 $T=25760 106080 0 0 $X=25570 $Y=105840
X1400 1 2 39 25 535 ICV_20 $T=43240 100640 0 0 $X=43050 $Y=100400
X1401 1 2 39 4 532 ICV_20 $T=44620 111520 0 0 $X=44430 $Y=111280
X1402 1 2 510 24 546 ICV_20 $T=50140 78880 0 0 $X=49950 $Y=78640
X1403 1 2 39 5 549 ICV_20 $T=53820 111520 0 0 $X=53630 $Y=111280
X1404 1 2 540 25 569 ICV_20 $T=62100 73440 0 0 $X=61910 $Y=73200
X1405 1 2 560 27 570 ICV_20 $T=62100 84320 0 0 $X=61910 $Y=84080
X1406 1 2 591 25 605 ICV_20 $T=79580 73440 1 0 $X=79390 $Y=70480
X1407 1 2 629 24 638 ICV_20 $T=99360 62560 0 0 $X=99170 $Y=62320
X1408 1 2 649 27 667 ICV_20 $T=110860 89760 1 0 $X=110670 $Y=86800
X1409 1 2 629 26 668 ICV_20 $T=111780 78880 1 0 $X=111590 $Y=75920
X1410 1 2 675 26 685 ICV_20 $T=121900 78880 1 0 $X=121710 $Y=75920
X1411 1 2 671 8 687 ICV_20 $T=122820 57120 1 0 $X=122630 $Y=54160
X1412 1 2 671 26 690 ICV_20 $T=123740 62560 1 0 $X=123550 $Y=59600
X1413 1 2 85 27 716 ICV_20 $T=137540 51680 0 0 $X=137350 $Y=51440
X1414 1 2 678 27 723 ICV_20 $T=141220 95200 1 0 $X=141030 $Y=92240
X1415 1 2 730 8 744 ICV_20 $T=148580 111520 1 0 $X=148390 $Y=108560
X1416 1 2 732 6 755 ICV_20 $T=155480 84320 0 0 $X=155290 $Y=84080
X1417 1 2 775 27 786 ICV_20 $T=171580 78880 1 0 $X=171390 $Y=75920
X1418 1 2 802 24 818 ICV_20 $T=186300 78880 0 0 $X=186110 $Y=78640
X1419 1 2 112 26 819 ICV_20 $T=187680 51680 0 0 $X=187490 $Y=51440
X1420 1 2 802 26 831 ICV_20 $T=194120 78880 0 0 $X=193930 $Y=78640
X1421 1 2 837 27 850 ICV_20 $T=207920 57120 0 0 $X=207730 $Y=56880
X1422 1 2 847 27 853 ICV_20 $T=211600 78880 0 0 $X=211410 $Y=78640
X1423 1 2 837 8 866 ICV_20 $T=218960 51680 0 0 $X=218770 $Y=51440
X1424 1 2 843 5 872 ICV_20 $T=222640 68000 1 0 $X=222450 $Y=65040
X1425 1 2 881 158 893 ICV_20 $T=234600 95200 0 0 $X=234410 $Y=94960
X1426 1 2 871 168 900 ICV_20 $T=236440 89760 1 0 $X=236250 $Y=86800
X1427 1 2 885 168 905 ICV_20 $T=240120 62560 0 0 $X=239930 $Y=62320
X1428 1 2 885 184 915 ICV_20 $T=248400 73440 0 0 $X=248210 $Y=73200
X1429 1 2 885 185 924 ICV_20 $T=249320 62560 1 0 $X=249130 $Y=59600
X1430 1 2 162 156 917 ICV_20 $T=249780 111520 1 0 $X=249590 $Y=108560
X1431 1 2 926 173 935 ICV_20 $T=257600 106080 1 0 $X=257410 $Y=103120
X1432 1 2 928 186 958 ICV_20 $T=270020 78880 0 0 $X=269830 $Y=78640
X1433 1 2 196 165 204 ICV_20 $T=276000 111520 0 0 $X=275810 $Y=111280
X1434 1 2 208 183 1013 ICV_20 $T=293020 51680 0 0 $X=292830 $Y=51440
X1435 1 2 1020 183 1037 ICV_20 $T=306360 84320 0 0 $X=306170 $Y=84080
X1436 1 2 1034 173 1048 ICV_20 $T=313260 100640 1 0 $X=313070 $Y=97680
X1437 1 2 1034 175 1056 ICV_20 $T=316020 89760 0 0 $X=315830 $Y=89520
X1438 1 2 214 184 1068 ICV_20 $T=321080 51680 0 0 $X=320890 $Y=51440
X1439 1 2 1033 186 1077 ICV_20 $T=326140 78880 0 0 $X=325950 $Y=78640
X1440 1 2 1078 173 1085 ICV_20 $T=333040 106080 1 0 $X=332850 $Y=103120
X1441 1 2 1078 175 1097 ICV_20 $T=334420 95200 0 0 $X=334230 $Y=94960
X1442 1 2 1089 183 1106 ICV_20 $T=340400 73440 1 0 $X=340210 $Y=70480
X1443 1 2 1089 166 1109 ICV_20 $T=342700 78880 0 0 $X=342510 $Y=78640
X1444 1 2 1102 164 1128 ICV_20 $T=353740 68000 0 0 $X=353550 $Y=67760
X1445 1 2 1145 167 1164 ICV_20 $T=368460 78880 1 0 $X=368270 $Y=75920
X1446 1 2 1188 166 1213 ICV_20 $T=396520 73440 1 0 $X=396330 $Y=70480
X1447 1 2 1248 158 1263 ICV_20 $T=418140 106080 0 0 $X=417950 $Y=105840
X1448 1 2 1248 165 1267 ICV_20 $T=419520 111520 1 0 $X=419330 $Y=108560
X1449 1 2 1256 186 1275 ICV_20 $T=424580 57120 1 0 $X=424390 $Y=54160
X1450 1 2 1239 185 1279 ICV_20 $T=426880 84320 0 0 $X=426690 $Y=84080
X1451 1 2 1250 156 1285 ICV_20 $T=431940 100640 1 0 $X=431750 $Y=97680
X1452 1 2 1239 186 1288 ICV_20 $T=432860 84320 1 0 $X=432670 $Y=81360
X1453 1 2 249 164 270 ICV_20 $T=444820 51680 1 0 $X=444630 $Y=48720
X1454 1 2 1301 257 1310 ICV_20 $T=445740 57120 0 0 $X=445550 $Y=56880
X1455 1 2 1301 265 1319 ICV_20 $T=446660 62560 0 0 $X=446470 $Y=62320
X1456 1 2 1304 259 1320 ICV_20 $T=446660 78880 0 0 $X=446470 $Y=78640
X1457 1 2 1305 262 1322 ICV_20 $T=446660 89760 0 0 $X=446470 $Y=89520
X1458 1 2 263 266 1323 ICV_20 $T=446660 111520 0 0 $X=446470 $Y=111280
X1459 1 2 263 258 1328 ICV_20 $T=448040 111520 1 0 $X=447850 $Y=108560
X1460 1 2 1292 272 1337 ICV_20 $T=454480 78880 1 0 $X=454290 $Y=75920
X1461 1 2 1335 259 1348 ICV_20 $T=459080 57120 0 0 $X=458890 $Y=56880
X1462 1 2 1335 258 1349 ICV_20 $T=459080 68000 0 0 $X=458890 $Y=67760
X1463 1 2 1301 272 1393 ICV_20 $T=483000 62560 0 0 $X=482810 $Y=62320
X1464 1 2 1381 297 1394 ICV_20 $T=483000 73440 1 0 $X=482810 $Y=70480
X1465 1 2 290 299 311 ICV_20 $T=490360 111520 0 0 $X=490170 $Y=111280
X1466 1 2 1409 301 1448 ICV_20 $T=509220 62560 1 0 $X=509030 $Y=59600
X1467 1 2 1420 259 1468 ICV_20 $T=516120 84320 1 0 $X=515930 $Y=81360
X1468 1 2 1471 264 1507 ICV_20 $T=537740 68000 1 0 $X=537550 $Y=65040
X1469 1 2 1500 265 1510 ICV_20 $T=539120 95200 0 0 $X=538930 $Y=94960
X1470 1 2 336 283 1558 ICV_20 $T=562120 57120 1 0 $X=561930 $Y=54160
X1471 1 2 1554 262 1573 ICV_20 $T=569480 89760 1 0 $X=569290 $Y=86800
X1472 1 2 1569 257 1588 ICV_20 $T=577300 57120 0 0 $X=577110 $Y=56880
X1473 1 2 1616 272 1636 ICV_20 $T=599840 73440 1 0 $X=599650 $Y=70480
X1474 1 2 1593 266 1626 ICV_20 $T=600300 100640 0 0 $X=600110 $Y=100400
X1475 1 2 1646 262 1667 ICV_20 $T=616860 62560 1 0 $X=616670 $Y=59600
X1476 1 2 1646 264 1668 ICV_20 $T=617780 73440 1 0 $X=617590 $Y=70480
X1477 1 2 1646 259 1673 ICV_20 $T=619620 57120 1 0 $X=619430 $Y=54160
X1478 1 2 1664 272 1698 ICV_20 $T=630660 111520 0 0 $X=630470 $Y=111280
X1479 1 2 1692 259 1700 ICV_20 $T=632960 68000 0 0 $X=632770 $Y=67760
X1480 1 2 1695 266 1696 ICV_20 $T=634800 95200 0 0 $X=634610 $Y=94960
X1481 1 2 1731 301 1749 ICV_20 $T=655040 89760 1 0 $X=654850 $Y=86800
X1482 1 2 383 305 385 ICV_20 $T=661020 111520 0 0 $X=660830 $Y=111280
X1483 1 2 1736 305 1756 ICV_20 $T=661940 51680 0 0 $X=661750 $Y=51440
X1484 1 2 1736 302 1757 ICV_20 $T=661940 57120 0 0 $X=661750 $Y=56880
X1485 1 2 1753 299 1758 ICV_20 $T=662860 73440 0 0 $X=662670 $Y=73200
X1486 1 2 1782 292 1792 ICV_20 $T=679420 62560 0 0 $X=679230 $Y=62320
X1487 1 2 393 301 395 ICV_20 $T=684480 51680 1 0 $X=684290 $Y=48720
X1488 1 2 1781 283 1803 ICV_20 $T=684480 84320 1 0 $X=684290 $Y=81360
X1489 1 2 1776 299 1818 ICV_20 $T=690920 100640 0 0 $X=690730 $Y=100400
X1490 1 2 1819 305 1860 ICV_20 $T=708860 89760 0 0 $X=708670 $Y=89520
X1491 1 2 452 4 460 ICV_21 $T=6900 68000 0 0 $X=6710 $Y=67760
X1492 1 2 3 8 461 ICV_21 $T=6900 111520 1 0 $X=6710 $Y=108560
X1493 1 2 512 4 531 ICV_21 $T=38640 95200 0 0 $X=38450 $Y=94960
X1494 1 2 512 5 550 ICV_21 $T=48300 89760 1 0 $X=48110 $Y=86800
X1495 1 2 39 24 557 ICV_21 $T=51060 100640 0 0 $X=50870 $Y=100400
X1496 1 2 540 8 57 ICV_21 $T=65320 68000 1 0 $X=65130 $Y=65040
X1497 1 2 678 24 693 ICV_21 $T=121440 95200 1 0 $X=121250 $Y=92240
X1498 1 2 741 8 780 ICV_21 $T=163300 95200 0 0 $X=163110 $Y=94960
X1499 1 2 776 8 783 ICV_21 $T=168820 106080 1 0 $X=168630 $Y=103120
X1500 1 2 790 6 828 ICV_21 $T=190440 62560 0 0 $X=190250 $Y=62320
X1501 1 2 909 164 929 ICV_21 $T=248860 89760 1 0 $X=248670 $Y=86800
X1502 1 2 1034 165 1061 ICV_21 $T=314640 95200 0 0 $X=314450 $Y=94960
X1503 1 2 1148 168 1160 ICV_21 $T=365240 68000 1 0 $X=365050 $Y=65040
X1504 1 2 1162 175 1195 ICV_21 $T=382720 95200 0 0 $X=382530 $Y=94960
X1505 1 2 1305 259 1326 ICV_21 $T=445280 89760 1 0 $X=445090 $Y=86800
X1506 1 2 1381 292 1413 ICV_21 $T=489440 73440 0 0 $X=489250 $Y=73200
X1507 1 2 290 301 1430 ICV_21 $T=498180 111520 0 0 $X=497990 $Y=111280
X1508 1 2 1418 265 1437 ICV_21 $T=500020 73440 0 0 $X=499830 $Y=73200
X1509 1 2 318 264 1490 ICV_21 $T=525780 111520 0 0 $X=525590 $Y=111280
X1510 1 2 331 302 1517 ICV_21 $T=539120 51680 0 0 $X=538930 $Y=51440
X1511 1 2 1491 264 1528 ICV_21 $T=546480 68000 0 0 $X=546290 $Y=67760
X1512 1 2 1569 264 1606 ICV_21 $T=584200 68000 0 0 $X=584010 $Y=67760
X1513 1 2 1637 272 1670 ICV_21 $T=615940 89760 1 0 $X=615750 $Y=86800
X1514 1 2 364 302 1672 ICV_21 $T=616860 51680 1 0 $X=616670 $Y=48720
X1515 1 2 1690 265 1722 ICV_21 $T=640320 84320 0 0 $X=640130 $Y=84080
X1516 1 2 1808 297 1844 ICV_21 $T=701040 73440 1 0 $X=700850 $Y=70480
X1517 1 2 730 24 768 768 740 30 ICV_22 $T=158700 100640 0 0 $X=158510 $Y=100400
X1518 1 2 732 4 772 772 748 20 ICV_22 $T=160540 84320 1 0 $X=160350 $Y=81360
X1519 1 2 1020 166 1066 1066 1038 171 ICV_22 $T=318780 84320 0 0 $X=318590 $Y=84080
X1520 1 2 1148 164 1184 1184 1149 169 ICV_22 $T=378120 73440 0 0 $X=377930 $Y=73200
X1521 1 2 1159 183 1190 1190 233 193 ICV_22 $T=382260 57120 0 0 $X=382070 $Y=56880
X1522 1 2 1248 160 1271 1267 253 188 ICV_22 $T=418600 106080 1 0 $X=418410 $Y=103120
X1523 1 2 1248 175 1298 1291 253 170 ICV_22 $T=432860 111520 0 0 $X=432670 $Y=111280
X1524 1 2 1527 258 1545 1526 1479 280 ICV_22 $T=553380 68000 1 0 $X=553190 $Y=65040
X1525 1 2 1781 299 1815 1803 1774 294 ICV_22 $T=686780 84320 0 0 $X=686590 $Y=84080
X1526 1 2 1819 297 1863 1863 1829 303 ICV_22 $T=707480 84320 0 0 $X=707290 $Y=84080
X1527 1 2 1817 283 1864 1864 1838 294 ICV_22 $T=707480 106080 0 0 $X=707290 $Y=105840
X1528 1 2 1866 283 1896 1896 1883 294 ICV_22 $T=729100 57120 1 0 $X=728910 $Y=54160
X1529 1 2 1866 287 1897 1897 1883 296 ICV_22 $T=729100 62560 1 0 $X=728910 $Y=59600
X1530 1 2 1868 283 1900 1900 1882 294 ICV_22 $T=729100 84320 1 0 $X=728910 $Y=81360
X1531 1 2 1865 287 1902 1905 1874 307 ICV_22 $T=729100 106080 1 0 $X=728910 $Y=103120
X1532 1 2 403 299 1871 409 397 294 ICV_22 $T=729100 111520 1 0 $X=728910 $Y=108560
X1533 1 2 ICV_23 $T=46460 84320 1 0 $X=46270 $Y=81360
X1534 1 2 ICV_23 $T=74520 95200 1 0 $X=74330 $Y=92240
X1535 1 2 ICV_23 $T=88320 62560 0 0 $X=88130 $Y=62320
X1536 1 2 ICV_23 $T=116380 78880 0 0 $X=116190 $Y=78640
X1537 1 2 ICV_23 $T=130640 57120 1 0 $X=130450 $Y=54160
X1538 1 2 ICV_23 $T=144440 68000 0 0 $X=144250 $Y=67760
X1539 1 2 ICV_23 $T=172500 51680 0 0 $X=172310 $Y=51440
X1540 1 2 ICV_23 $T=186760 51680 1 0 $X=186570 $Y=48720
X1541 1 2 ICV_23 $T=186760 111520 1 0 $X=186570 $Y=108560
X1542 1 2 ICV_23 $T=214820 51680 1 0 $X=214630 $Y=48720
X1543 1 2 ICV_23 $T=228620 51680 0 0 $X=228430 $Y=51440
X1544 1 2 ICV_23 $T=228620 95200 0 0 $X=228430 $Y=94960
X1545 1 2 ICV_23 $T=242880 78880 1 0 $X=242690 $Y=75920
X1546 1 2 ICV_23 $T=270940 89760 1 0 $X=270750 $Y=86800
X1547 1 2 ICV_23 $T=299000 51680 1 0 $X=298810 $Y=48720
X1548 1 2 ICV_23 $T=312800 78880 0 0 $X=312610 $Y=78640
X1549 1 2 ICV_23 $T=327060 111520 1 0 $X=326870 $Y=108560
X1550 1 2 ICV_23 $T=340860 62560 0 0 $X=340670 $Y=62320
X1551 1 2 ICV_23 $T=383180 111520 1 0 $X=382990 $Y=108560
X1552 1 2 ICV_23 $T=467360 57120 1 0 $X=467170 $Y=54160
X1553 1 2 ICV_23 $T=495420 62560 1 0 $X=495230 $Y=59600
X1554 1 2 ICV_23 $T=495420 95200 1 0 $X=495230 $Y=92240
X1555 1 2 ICV_23 $T=537280 73440 0 0 $X=537090 $Y=73200
X1556 1 2 ICV_23 $T=565340 73440 0 0 $X=565150 $Y=73200
X1557 1 2 ICV_23 $T=579600 51680 1 0 $X=579410 $Y=48720
X1558 1 2 ICV_23 $T=579600 62560 1 0 $X=579410 $Y=59600
X1559 1 2 ICV_23 $T=607660 73440 1 0 $X=607470 $Y=70480
X1560 1 2 ICV_23 $T=607660 95200 1 0 $X=607470 $Y=92240
X1561 1 2 ICV_23 $T=621460 51680 0 0 $X=621270 $Y=51440
X1562 1 2 ICV_23 $T=621460 73440 0 0 $X=621270 $Y=73200
X1563 1 2 ICV_23 $T=663780 106080 1 0 $X=663590 $Y=103120
X1564 1 2 ICV_23 $T=677580 89760 0 0 $X=677390 $Y=89520
X1565 1 2 ICV_23 $T=691840 68000 1 0 $X=691650 $Y=65040
X1566 1 2 ICV_24 $T=74060 73440 1 0 $X=73870 $Y=70480
X1567 1 2 ICV_24 $T=74060 100640 1 0 $X=73870 $Y=97680
X1568 1 2 ICV_24 $T=87860 68000 0 0 $X=87670 $Y=67760
X1569 1 2 ICV_24 $T=87860 100640 0 0 $X=87670 $Y=100400
X1570 1 2 ICV_24 $T=172040 84320 0 0 $X=171850 $Y=84080
X1571 1 2 ICV_24 $T=214360 106080 1 0 $X=214170 $Y=103120
X1572 1 2 ICV_24 $T=256220 73440 0 0 $X=256030 $Y=73200
X1573 1 2 ICV_24 $T=256220 95200 0 0 $X=256030 $Y=94960
X1574 1 2 ICV_24 $T=256220 111520 0 0 $X=256030 $Y=111280
X1575 1 2 ICV_24 $T=270480 73440 1 0 $X=270290 $Y=70480
X1576 1 2 ICV_24 $T=312340 51680 0 0 $X=312150 $Y=51440
X1577 1 2 ICV_24 $T=312340 95200 0 0 $X=312150 $Y=94960
X1578 1 2 ICV_24 $T=312340 100640 0 0 $X=312150 $Y=100400
X1579 1 2 ICV_24 $T=382720 84320 1 0 $X=382530 $Y=81360
X1580 1 2 ICV_24 $T=382720 106080 1 0 $X=382530 $Y=103120
X1581 1 2 ICV_24 $T=480700 95200 0 0 $X=480510 $Y=94960
X1582 1 2 ICV_24 $T=508760 62560 0 0 $X=508570 $Y=62320
X1583 1 2 ICV_24 $T=508760 111520 0 0 $X=508570 $Y=111280
X1584 1 2 ICV_24 $T=564880 89760 0 0 $X=564690 $Y=89520
X1585 1 2 ICV_24 $T=564880 111520 0 0 $X=564690 $Y=111280
X1586 1 2 ICV_24 $T=663320 68000 1 0 $X=663130 $Y=65040
X1587 1 2 ICV_24 $T=663320 78880 1 0 $X=663130 $Y=75920
X1588 1 2 ICV_24 $T=705180 111520 0 0 $X=704990 $Y=111280
X1589 1 2 15 2 473 1 sky130_fd_sc_hd__inv_1 $T=18400 95200 1 0 $X=18210 $Y=92240
X1590 1 2 16 2 451 1 sky130_fd_sc_hd__inv_1 $T=18400 106080 1 0 $X=18210 $Y=103120
X1591 1 2 22 2 477 1 sky130_fd_sc_hd__inv_1 $T=24380 84320 1 0 $X=24190 $Y=81360
X1592 1 2 12 2 9 1 sky130_fd_sc_hd__inv_1 $T=25760 51680 1 0 $X=25570 $Y=48720
X1593 1 2 23 2 14 1 sky130_fd_sc_hd__inv_1 $T=28520 111520 0 0 $X=28330 $Y=111280
X1594 1 2 43 2 44 1 sky130_fd_sc_hd__inv_1 $T=52440 111520 0 0 $X=52250 $Y=111280
X1595 1 2 28 2 525 1 sky130_fd_sc_hd__inv_1 $T=52900 73440 1 0 $X=52710 $Y=70480
X1596 1 2 41 2 40 1 sky130_fd_sc_hd__inv_1 $T=60260 51680 1 0 $X=60070 $Y=48720
X1597 1 2 37 2 533 1 sky130_fd_sc_hd__inv_1 $T=60260 95200 0 0 $X=60070 $Y=94960
X1598 1 2 50 2 534 1 sky130_fd_sc_hd__inv_1 $T=62100 111520 0 0 $X=61910 $Y=111280
X1599 1 2 46 2 53 1 sky130_fd_sc_hd__inv_1 $T=74520 57120 1 0 $X=74330 $Y=54160
X1600 1 2 42 2 47 1 sky130_fd_sc_hd__inv_1 $T=76360 68000 1 0 $X=76170 $Y=65040
X1601 1 2 48 2 573 1 sky130_fd_sc_hd__inv_1 $T=78200 84320 1 0 $X=78010 $Y=81360
X1602 1 2 49 2 563 1 sky130_fd_sc_hd__inv_1 $T=86480 100640 0 0 $X=86290 $Y=100400
X1603 1 2 58 2 586 1 sky130_fd_sc_hd__inv_1 $T=96140 73440 1 0 $X=95950 $Y=70480
X1604 1 2 65 2 68 1 sky130_fd_sc_hd__inv_1 $T=101660 106080 1 0 $X=101470 $Y=103120
X1605 1 2 60 2 64 1 sky130_fd_sc_hd__inv_1 $T=102120 57120 1 0 $X=101930 $Y=54160
X1606 1 2 61 2 615 1 sky130_fd_sc_hd__inv_1 $T=102580 84320 1 0 $X=102390 $Y=81360
X1607 1 2 79 2 632 1 sky130_fd_sc_hd__inv_1 $T=116380 73440 0 0 $X=116190 $Y=73200
X1608 1 2 76 2 644 1 sky130_fd_sc_hd__inv_1 $T=116380 106080 0 0 $X=116190 $Y=105840
X1609 1 2 78 2 80 1 sky130_fd_sc_hd__inv_1 $T=119600 51680 0 0 $X=119410 $Y=51440
X1610 1 2 77 2 692 1 sky130_fd_sc_hd__inv_1 $T=130640 68000 1 0 $X=130450 $Y=65040
X1611 1 2 94 2 700 1 sky130_fd_sc_hd__inv_1 $T=149040 95200 1 0 $X=148850 $Y=92240
X1612 1 2 83 2 90 1 sky130_fd_sc_hd__inv_1 $T=151340 51680 1 0 $X=151150 $Y=48720
X1613 1 2 104 2 740 1 sky130_fd_sc_hd__inv_1 $T=167900 111520 1 0 $X=167710 $Y=108560
X1614 1 2 99 2 748 1 sky130_fd_sc_hd__inv_1 $T=170660 84320 0 0 $X=170470 $Y=84080
X1615 1 2 100 2 760 1 sky130_fd_sc_hd__inv_1 $T=174340 68000 0 0 $X=174150 $Y=67760
X1616 1 2 103 2 734 1 sky130_fd_sc_hd__inv_1 $T=177100 95200 1 0 $X=176910 $Y=92240
X1617 1 2 111 2 784 1 sky130_fd_sc_hd__inv_1 $T=185380 111520 1 0 $X=185190 $Y=108560
X1618 1 2 106 2 792 1 sky130_fd_sc_hd__inv_1 $T=186760 78880 1 0 $X=186570 $Y=75920
X1619 1 2 127 2 826 1 sky130_fd_sc_hd__inv_1 $T=202400 73440 0 0 $X=202210 $Y=73200
X1620 1 2 109 2 810 1 sky130_fd_sc_hd__inv_1 $T=206540 57120 0 0 $X=206350 $Y=56880
X1621 1 2 115 2 817 1 sky130_fd_sc_hd__inv_1 $T=210220 89760 1 0 $X=210030 $Y=86800
X1622 1 2 140 2 139 1 sky130_fd_sc_hd__inv_1 $T=227240 51680 0 0 $X=227050 $Y=51440
X1623 1 2 129 2 857 1 sky130_fd_sc_hd__inv_1 $T=234600 84320 0 0 $X=234410 $Y=84080
X1624 1 2 22 2 886 1 sky130_fd_sc_hd__inv_1 $T=238740 84320 1 0 $X=238550 $Y=81360
X1625 1 2 151 2 891 1 sky130_fd_sc_hd__inv_1 $T=242420 95200 0 0 $X=242230 $Y=94960
X1626 1 2 131 2 179 1 sky130_fd_sc_hd__inv_1 $T=246560 111520 0 0 $X=246370 $Y=111280
X1627 1 2 28 2 890 1 sky130_fd_sc_hd__inv_1 $T=247020 73440 0 0 $X=246830 $Y=73200
X1628 1 2 41 2 176 1 sky130_fd_sc_hd__inv_1 $T=249320 51680 1 0 $X=249130 $Y=48720
X1629 1 2 15 2 923 1 sky130_fd_sc_hd__inv_1 $T=255300 89760 0 0 $X=255110 $Y=89520
X1630 1 2 43 2 198 1 sky130_fd_sc_hd__inv_1 $T=264960 111520 0 0 $X=264770 $Y=111280
X1631 1 2 142 2 943 1 sky130_fd_sc_hd__inv_1 $T=265880 106080 1 0 $X=265690 $Y=103120
X1632 1 2 12 2 201 1 sky130_fd_sc_hd__inv_1 $T=270480 51680 1 0 $X=270290 $Y=48720
X1633 1 2 42 2 967 1 sky130_fd_sc_hd__inv_1 $T=284740 62560 0 0 $X=284550 $Y=62320
X1634 1 2 61 2 977 1 sky130_fd_sc_hd__inv_1 $T=288880 89760 1 0 $X=288690 $Y=86800
X1635 1 2 48 2 988 1 sky130_fd_sc_hd__inv_1 $T=294860 78880 1 0 $X=294670 $Y=75920
X1636 1 2 67 2 1005 1 sky130_fd_sc_hd__inv_1 $T=298080 95200 0 0 $X=297890 $Y=94960
X1637 1 2 46 2 212 1 sky130_fd_sc_hd__inv_1 $T=302220 57120 1 0 $X=302030 $Y=54160
X1638 1 2 77 2 1018 1 sky130_fd_sc_hd__inv_1 $T=308200 68000 1 0 $X=308010 $Y=65040
X1639 1 2 94 2 1038 1 sky130_fd_sc_hd__inv_1 $T=314640 89760 0 0 $X=314450 $Y=89520
X1640 1 2 153 2 211 1 sky130_fd_sc_hd__inv_1 $T=314640 111520 0 0 $X=314450 $Y=111280
X1641 1 2 79 2 1039 1 sky130_fd_sc_hd__inv_1 $T=315560 78880 0 0 $X=315370 $Y=78640
X1642 1 2 133 2 1053 1 sky130_fd_sc_hd__inv_1 $T=322460 100640 1 0 $X=322270 $Y=97680
X1643 1 2 58 2 1071 1 sky130_fd_sc_hd__inv_1 $T=331200 68000 1 0 $X=331010 $Y=65040
X1644 1 2 148 2 1074 1 sky130_fd_sc_hd__inv_1 $T=332580 100640 0 0 $X=332390 $Y=100400
X1645 1 2 60 2 221 1 sky130_fd_sc_hd__inv_1 $T=340400 51680 0 0 $X=340210 $Y=51440
X1646 1 2 122 2 222 1 sky130_fd_sc_hd__inv_1 $T=340860 111520 0 0 $X=340670 $Y=111280
X1647 1 2 100 2 1101 1 sky130_fd_sc_hd__inv_1 $T=344540 68000 1 0 $X=344350 $Y=65040
X1648 1 2 87 2 1100 1 sky130_fd_sc_hd__inv_1 $T=346840 84320 1 0 $X=346650 $Y=81360
X1649 1 2 71 2 1110 1 sky130_fd_sc_hd__inv_1 $T=352820 89760 1 0 $X=352630 $Y=86800
X1650 1 2 78 2 226 1 sky130_fd_sc_hd__inv_1 $T=355120 51680 1 0 $X=354930 $Y=48720
X1651 1 2 106 2 1149 1 sky130_fd_sc_hd__inv_1 $T=368920 73440 0 0 $X=368730 $Y=73200
X1652 1 2 99 2 1157 1 sky130_fd_sc_hd__inv_1 $T=378120 78880 0 0 $X=377930 $Y=78640
X1653 1 2 145 2 232 1 sky130_fd_sc_hd__inv_1 $T=390540 111520 0 0 $X=390350 $Y=111280
X1654 1 2 103 2 1199 1 sky130_fd_sc_hd__inv_1 $T=396980 89760 0 0 $X=396790 $Y=89520
X1655 1 2 127 2 1210 1 sky130_fd_sc_hd__inv_1 $T=402040 78880 1 0 $X=401850 $Y=75920
X1656 1 2 143 2 1212 1 sky130_fd_sc_hd__inv_1 $T=402500 106080 1 0 $X=402310 $Y=103120
X1657 1 2 93 2 1228 1 sky130_fd_sc_hd__inv_1 $T=410320 62560 0 0 $X=410130 $Y=62320
X1658 1 2 115 2 1246 1 sky130_fd_sc_hd__inv_1 $T=419980 89760 0 0 $X=419790 $Y=89520
X1659 1 2 129 2 1261 1 sky130_fd_sc_hd__inv_1 $T=422280 84320 1 0 $X=422090 $Y=81360
X1660 1 2 134 2 1262 1 sky130_fd_sc_hd__inv_1 $T=424120 68000 1 0 $X=423930 $Y=65040
X1661 1 2 140 2 252 1 sky130_fd_sc_hd__inv_1 $T=427340 51680 1 0 $X=427150 $Y=48720
X1662 1 2 150 2 253 1 sky130_fd_sc_hd__inv_1 $T=427800 111520 1 0 $X=427610 $Y=108560
X1663 1 2 132 2 1270 1 sky130_fd_sc_hd__inv_1 $T=431020 95200 0 0 $X=430830 $Y=94960
X1664 1 2 281 2 271 1 sky130_fd_sc_hd__inv_1 $T=467360 111520 0 0 $X=467170 $Y=111280
X1665 1 2 260 2 1331 1 sky130_fd_sc_hd__inv_1 $T=472880 95200 0 0 $X=472690 $Y=94960
X1666 1 2 274 2 1345 1 sky130_fd_sc_hd__inv_1 $T=473340 62560 1 0 $X=473150 $Y=59600
X1667 1 2 285 2 1315 1 sky130_fd_sc_hd__inv_1 $T=476560 106080 1 0 $X=476370 $Y=103120
X1668 1 2 279 2 1333 1 sky130_fd_sc_hd__inv_1 $T=480700 84320 0 0 $X=480510 $Y=84080
X1669 1 2 284 2 1311 1 sky130_fd_sc_hd__inv_1 $T=481160 78880 1 0 $X=480970 $Y=75920
X1670 1 2 289 2 1312 1 sky130_fd_sc_hd__inv_1 $T=483000 57120 0 0 $X=482810 $Y=56880
X1671 1 2 291 2 1357 1 sky130_fd_sc_hd__inv_1 $T=495880 57120 0 0 $X=495690 $Y=56880
X1672 1 2 308 2 1389 1 sky130_fd_sc_hd__inv_1 $T=499100 95200 0 0 $X=498910 $Y=94960
X1673 1 2 284 2 1386 1 sky130_fd_sc_hd__inv_1 $T=500020 78880 0 0 $X=499830 $Y=78640
X1674 1 2 295 2 1399 1 sky130_fd_sc_hd__inv_1 $T=504620 95200 0 0 $X=504430 $Y=94960
X1675 1 2 317 2 1431 1 sky130_fd_sc_hd__inv_1 $T=512440 89760 1 0 $X=512250 $Y=86800
X1676 1 2 306 2 1428 1 sky130_fd_sc_hd__inv_1 $T=517040 62560 1 0 $X=516850 $Y=59600
X1677 1 2 312 2 1446 1 sky130_fd_sc_hd__inv_1 $T=522560 100640 1 0 $X=522370 $Y=97680
X1678 1 2 319 2 323 1 sky130_fd_sc_hd__inv_1 $T=536820 51680 0 0 $X=536630 $Y=51440
X1679 1 2 322 2 1498 1 sky130_fd_sc_hd__inv_1 $T=537280 84320 0 0 $X=537090 $Y=84080
X1680 1 2 316 2 1461 1 sky130_fd_sc_hd__inv_1 $T=539120 100640 0 0 $X=538930 $Y=100400
X1681 1 2 332 2 1479 1 sky130_fd_sc_hd__inv_1 $T=550620 62560 1 0 $X=550430 $Y=59600
X1682 1 2 324 2 1512 1 sky130_fd_sc_hd__inv_1 $T=552460 73440 0 0 $X=552270 $Y=73200
X1683 1 2 281 2 334 1 sky130_fd_sc_hd__inv_1 $T=560740 57120 1 0 $X=560550 $Y=54160
X1684 1 2 327 2 1513 1 sky130_fd_sc_hd__inv_1 $T=560740 100640 1 0 $X=560550 $Y=97680
X1685 1 2 330 2 1525 1 sky130_fd_sc_hd__inv_1 $T=568100 89760 1 0 $X=567910 $Y=86800
X1686 1 2 337 2 1546 1 sky130_fd_sc_hd__inv_1 $T=571780 68000 1 0 $X=571590 $Y=65040
X1687 1 2 337 2 340 1 sky130_fd_sc_hd__inv_1 $T=575920 57120 0 0 $X=575730 $Y=56880
X1688 1 2 348 2 1551 1 sky130_fd_sc_hd__inv_1 $T=579600 106080 1 0 $X=579410 $Y=103120
X1689 1 2 343 2 345 1 sky130_fd_sc_hd__inv_1 $T=584200 106080 0 0 $X=584010 $Y=105840
X1690 1 2 355 2 1582 1 sky130_fd_sc_hd__inv_1 $T=592480 68000 1 0 $X=592290 $Y=65040
X1691 1 2 289 2 354 1 sky130_fd_sc_hd__inv_1 $T=598000 57120 1 0 $X=597810 $Y=54160
X1692 1 2 359 2 1600 1 sky130_fd_sc_hd__inv_1 $T=603060 106080 1 0 $X=602870 $Y=103120
X1693 1 2 351 2 1601 1 sky130_fd_sc_hd__inv_1 $T=606280 95200 1 0 $X=606090 $Y=92240
X1694 1 2 360 2 1625 1 sky130_fd_sc_hd__inv_1 $T=607660 68000 1 0 $X=607470 $Y=65040
X1695 1 2 279 2 365 1 sky130_fd_sc_hd__inv_1 $T=609500 57120 1 0 $X=609310 $Y=54160
X1696 1 2 363 2 1657 1 sky130_fd_sc_hd__inv_1 $T=624680 73440 0 0 $X=624490 $Y=73200
X1697 1 2 369 2 1660 1 sky130_fd_sc_hd__inv_1 $T=627440 100640 1 0 $X=627250 $Y=97680
X1698 1 2 366 2 1674 1 sky130_fd_sc_hd__inv_1 $T=637560 62560 1 0 $X=637370 $Y=59600
X1699 1 2 368 2 1688 1 sky130_fd_sc_hd__inv_1 $T=651360 106080 0 0 $X=651170 $Y=105840
X1700 1 2 372 2 1709 1 sky130_fd_sc_hd__inv_1 $T=655500 57120 1 0 $X=655310 $Y=54160
X1701 1 2 375 2 1701 1 sky130_fd_sc_hd__inv_1 $T=658260 84320 1 0 $X=658070 $Y=81360
X1702 1 2 373 2 1697 1 sky130_fd_sc_hd__inv_1 $T=658260 95200 0 0 $X=658070 $Y=94960
X1703 1 2 322 2 1746 1 sky130_fd_sc_hd__inv_1 $T=663780 95200 1 0 $X=663590 $Y=92240
X1704 1 2 343 2 1748 1 sky130_fd_sc_hd__inv_1 $T=666540 78880 0 0 $X=666350 $Y=78640
X1705 1 2 348 2 386 1 sky130_fd_sc_hd__inv_1 $T=672060 100640 0 0 $X=671870 $Y=100400
X1706 1 2 356 2 384 1 sky130_fd_sc_hd__inv_1 $T=673900 62560 0 0 $X=673710 $Y=62320
X1707 1 2 317 2 1774 1 sky130_fd_sc_hd__inv_1 $T=685860 89760 0 0 $X=685670 $Y=89520
X1708 1 2 373 2 1800 1 sky130_fd_sc_hd__inv_1 $T=691380 100640 1 0 $X=691190 $Y=97680
X1709 1 2 308 2 1798 1 sky130_fd_sc_hd__inv_1 $T=691840 73440 0 0 $X=691650 $Y=73200
X1710 1 2 363 2 1816 1 sky130_fd_sc_hd__inv_1 $T=700120 78880 1 0 $X=699930 $Y=75920
X1711 1 2 346 2 1829 1 sky130_fd_sc_hd__inv_1 $T=707480 89760 0 0 $X=707290 $Y=89520
X1712 1 2 368 2 1838 1 sky130_fd_sc_hd__inv_1 $T=721280 106080 0 0 $X=721090 $Y=105840
X1713 1 2 372 2 404 1 sky130_fd_sc_hd__inv_1 $T=721740 51680 0 0 $X=721550 $Y=51440
X1714 1 2 375 2 1869 1 sky130_fd_sc_hd__inv_1 $T=721740 78880 1 0 $X=721550 $Y=75920
X1715 1 2 351 2 1882 1 sky130_fd_sc_hd__inv_1 $T=729100 89760 1 0 $X=728910 $Y=86800
X1716 1 2 369 2 1874 1 sky130_fd_sc_hd__inv_1 $T=729100 100640 1 0 $X=728910 $Y=97680
X1717 1 2 370 2 1883 1 sky130_fd_sc_hd__inv_1 $T=731400 62560 0 0 $X=731210 $Y=62320
X1718 1 2 463 477 20 ICV_26 $T=17940 73440 0 0 $X=17750 $Y=73200
X1719 1 2 469 451 18 ICV_26 $T=18400 100640 0 0 $X=18210 $Y=100400
X1720 1 2 494 473 30 ICV_26 $T=33580 84320 1 0 $X=33390 $Y=81360
X1721 1 2 501 9 34 ICV_26 $T=34040 51680 0 0 $X=33850 $Y=51440
X1722 1 2 503 451 33 ICV_26 $T=34040 95200 0 0 $X=33850 $Y=94960
X1723 1 2 548 47 30 ICV_26 $T=57040 73440 0 0 $X=56850 $Y=73200
X1724 1 2 617 615 34 ICV_26 $T=96140 78880 1 0 $X=95950 $Y=75920
X1725 1 2 647 632 34 ICV_26 $T=107180 78880 1 0 $X=106990 $Y=75920
X1726 1 2 663 643 20 ICV_26 $T=116840 95200 1 0 $X=116650 $Y=92240
X1727 1 2 667 643 34 ICV_26 $T=118220 89760 0 0 $X=118030 $Y=89520
X1728 1 2 745 102 33 ICV_26 $T=155480 51680 1 0 $X=155290 $Y=48720
X1729 1 2 853 857 34 ICV_26 $T=218040 73440 0 0 $X=217850 $Y=73200
X1730 1 2 868 856 11 ICV_26 $T=225400 73440 0 0 $X=225210 $Y=73200
X1731 1 2 887 890 169 ICV_26 $T=239660 73440 1 0 $X=239470 $Y=70480
X1732 1 2 903 176 177 ICV_26 $T=244720 51680 1 0 $X=244530 $Y=48720
X1733 1 2 902 892 177 ICV_26 $T=244720 62560 1 0 $X=244530 $Y=59600
X1734 1 2 911 891 187 ICV_26 $T=251160 95200 1 0 $X=250970 $Y=92240
X1735 1 2 914 892 171 ICV_26 $T=253460 51680 0 0 $X=253270 $Y=51440
X1736 1 2 917 179 170 ICV_26 $T=253460 106080 0 0 $X=253270 $Y=105840
X1737 1 2 1048 1053 191 ICV_26 $T=323840 100640 1 0 $X=323650 $Y=97680
X1738 1 2 1097 1074 187 ICV_26 $T=343160 95200 1 0 $X=342970 $Y=92240
X1739 1 2 1121 222 170 ICV_26 $T=351900 111520 1 0 $X=351710 $Y=108560
X1740 1 2 1128 1101 169 ICV_26 $T=359720 73440 1 0 $X=359530 $Y=70480
X1741 1 2 1186 1157 193 ICV_26 $T=388240 78880 0 0 $X=388050 $Y=78640
X1742 1 2 1195 1168 187 ICV_26 $T=391920 100640 1 0 $X=391730 $Y=97680
X1743 1 2 1223 1199 194 ICV_26 $T=404800 84320 1 0 $X=404610 $Y=81360
X1744 1 2 1279 1246 194 ICV_26 $T=438380 78880 0 0 $X=438190 $Y=78640
X1745 1 2 1297 1262 171 ICV_26 $T=441140 62560 1 0 $X=440950 $Y=59600
X1746 1 2 1341 271 273 ICV_26 $T=463220 106080 0 0 $X=463030 $Y=105840
X1747 1 2 1343 1345 268 ICV_26 $T=464140 51680 1 0 $X=463950 $Y=48720
X1748 1 2 1359 1345 277 ICV_26 $T=472880 73440 1 0 $X=472690 $Y=70480
X1749 1 2 1358 1357 294 ICV_26 $T=474260 51680 0 0 $X=474070 $Y=51440
X1750 1 2 1394 1386 303 ICV_26 $T=489900 68000 1 0 $X=489710 $Y=65040
X1751 1 2 1429 1431 277 ICV_26 $T=506000 95200 0 0 $X=505810 $Y=94960
X1752 1 2 1442 315 288 ICV_26 $T=511060 51680 0 0 $X=510870 $Y=51440
X1753 1 2 1465 1461 273 ICV_26 $T=521180 111520 0 0 $X=520990 $Y=111280
X1754 1 2 1560 1551 277 ICV_26 $T=569940 111520 0 0 $X=569750 $Y=111280
X1755 1 2 1626 1601 277 ICV_26 $T=604440 106080 1 0 $X=604250 $Y=103120
X1756 1 2 1675 1657 269 ICV_26 $T=626520 89760 1 0 $X=626330 $Y=86800
X1757 1 2 1687 1688 277 ICV_26 $T=630660 100640 0 0 $X=630470 $Y=100400
X1758 1 2 1720 1701 268 ICV_26 $T=646300 78880 0 0 $X=646110 $Y=78640
X1759 1 2 1725 1688 275 ICV_26 $T=652740 111520 1 0 $X=652550 $Y=108560
X1760 1 2 1894 1869 304 ICV_26 $T=737380 51680 1 0 $X=737190 $Y=48720
X1761 1 2 449 4 455 ICV_28 $T=6900 95200 1 0 $X=6710 $Y=92240
X1762 1 2 3 5 456 ICV_28 $T=6900 111520 0 0 $X=6710 $Y=111280
X1763 1 2 452 24 491 ICV_28 $T=24380 68000 1 0 $X=24190 $Y=65040
X1764 1 2 509 26 523 ICV_28 $T=37720 62560 1 0 $X=37530 $Y=59600
X1765 1 2 51 26 577 ICV_28 $T=63940 111520 1 0 $X=63750 $Y=108560
X1766 1 2 591 24 625 ICV_28 $T=90160 62560 0 0 $X=89970 $Y=62320
X1767 1 2 671 27 689 ICV_28 $T=121440 68000 1 0 $X=121250 $Y=65040
X1768 1 2 675 5 711 ICV_28 $T=133400 78880 0 0 $X=133210 $Y=78640
X1769 1 2 708 8 718 ICV_28 $T=136620 62560 0 0 $X=136430 $Y=62320
X1770 1 2 741 25 785 ICV_28 $T=167900 95200 1 0 $X=167710 $Y=92240
X1771 1 2 802 5 836 ICV_28 $T=195960 84320 1 0 $X=195770 $Y=81360
X1772 1 2 989 173 1001 ICV_28 $T=287500 106080 1 0 $X=287310 $Y=103120
X1773 1 2 959 185 992 ICV_28 $T=290260 89760 1 0 $X=290070 $Y=86800
X1774 1 2 207 175 1011 ICV_28 $T=290720 106080 0 0 $X=290530 $Y=105840
X1775 1 2 1124 181 1144 ICV_28 $T=357420 100640 0 0 $X=357230 $Y=100400
X1776 1 2 231 165 1171 ICV_28 $T=370760 111520 0 0 $X=370570 $Y=111280
X1777 1 2 1239 184 1244 ICV_28 $T=413080 84320 1 0 $X=412890 $Y=81360
X1778 1 2 1242 164 1276 ICV_28 $T=423660 84320 1 0 $X=423470 $Y=81360
X1779 1 2 1375 266 1388 ICV_28 $T=477940 106080 1 0 $X=477750 $Y=103120
X1780 1 2 1420 257 1438 ICV_28 $T=501400 78880 0 0 $X=501210 $Y=78640
X1781 1 2 1569 262 1605 ICV_28 $T=585120 62560 0 0 $X=584930 $Y=62320
X1782 1 2 1616 257 1622 ICV_28 $T=595240 57120 0 0 $X=595050 $Y=56880
X1783 1 2 1640 258 1658 ICV_28 $T=609500 100640 1 0 $X=609310 $Y=97680
X1784 1 2 1731 305 1743 ICV_28 $T=654580 95200 1 0 $X=654390 $Y=92240
X1785 1 2 1808 283 1826 ICV_28 $T=693680 68000 1 0 $X=693490 $Y=65040
X1786 1 2 449 5 457 ICV_29 $T=6900 89760 0 0 $X=6710 $Y=89520
X1787 1 2 3 25 506 ICV_29 $T=26680 111520 1 0 $X=26490 $Y=108560
X1788 1 2 540 27 565 ICV_29 $T=55660 68000 1 0 $X=55470 $Y=65040
X1789 1 2 566 27 581 ICV_29 $T=64860 95200 1 0 $X=64670 $Y=92240
X1790 1 2 540 4 582 ICV_29 $T=66240 62560 0 0 $X=66050 $Y=62320
X1791 1 2 560 8 583 ICV_29 $T=66240 89760 1 0 $X=66050 $Y=86800
X1792 1 2 566 4 598 ICV_29 $T=76360 95200 1 0 $X=76170 $Y=92240
X1793 1 2 591 6 606 ICV_29 $T=78200 68000 0 0 $X=78010 $Y=67760
X1794 1 2 629 25 645 ICV_29 $T=97520 73440 0 0 $X=97330 $Y=73200
X1795 1 2 629 8 670 ICV_29 $T=111780 68000 1 0 $X=111590 $Y=65040
X1796 1 2 802 8 815 ICV_29 $T=182620 84320 0 0 $X=182430 $Y=84080
X1797 1 2 112 27 825 ICV_29 $T=188600 51680 1 0 $X=188410 $Y=48720
X1798 1 2 802 27 832 ICV_29 $T=192280 84320 0 0 $X=192090 $Y=84080
X1799 1 2 1034 160 1058 ICV_29 $T=314640 100640 0 0 $X=314450 $Y=100400
X1800 1 2 1124 175 1155 ICV_29 $T=364320 100640 1 0 $X=364130 $Y=97680
X1801 1 2 1148 184 1181 ICV_29 $T=378120 62560 0 0 $X=377930 $Y=62320
X1802 1 2 1188 167 1209 ICV_29 $T=392380 78880 1 0 $X=392190 $Y=75920
X1803 1 2 1180 164 1214 ICV_29 $T=395140 84320 1 0 $X=394950 $Y=81360
X1804 1 2 263 262 1341 ICV_29 $T=455860 111520 1 0 $X=455670 $Y=108560
X1805 1 2 282 287 1371 ICV_29 $T=469200 57120 1 0 $X=469010 $Y=54160
X1806 1 2 1381 299 1404 ICV_29 $T=483000 78880 0 0 $X=482810 $Y=78640
X1807 1 2 1381 302 1412 ICV_29 $T=490360 68000 0 0 $X=490170 $Y=67760
X1808 1 2 1473 266 1486 ICV_29 $T=525320 78880 1 0 $X=525130 $Y=75920
X1809 1 2 1554 258 1570 ICV_29 $T=567180 78880 0 0 $X=566990 $Y=78640
X1810 1 2 1569 258 1581 ICV_29 $T=574540 68000 0 0 $X=574350 $Y=67760
X1811 1 2 1544 262 1584 ICV_29 $T=574540 95200 0 0 $X=574350 $Y=94960
X1812 1 2 1569 265 1589 ICV_29 $T=575460 62560 0 0 $X=575270 $Y=62320
X1813 1 2 1637 262 1666 ICV_29 $T=613640 78880 1 0 $X=613450 $Y=75920
X1814 1 2 1690 264 1699 ICV_29 $T=630660 84320 0 0 $X=630470 $Y=84080
X1815 1 2 1695 258 1728 ICV_29 $T=644920 95200 1 0 $X=644730 $Y=92240
X1816 1 2 457 473 17 455 473 20 ICV_30 $T=17480 89760 0 0 $X=17290 $Y=89520
X1817 1 2 467 476 11 474 9 17 ICV_30 $T=18860 57120 0 0 $X=18670 $Y=56880
X1818 1 2 486 477 30 507 508 32 ICV_30 $T=31740 73440 1 0 $X=31550 $Y=70480
X1819 1 2 504 451 32 497 451 30 ICV_30 $T=34960 100640 0 0 $X=34770 $Y=100400
X1820 1 2 515 508 20 520 508 34 ICV_30 $T=41860 78880 0 0 $X=41670 $Y=78640
X1821 1 2 528 533 33 527 533 34 ICV_30 $T=48300 95200 1 0 $X=48110 $Y=92240
X1822 1 2 541 525 11 551 47 32 ICV_30 $T=54280 73440 1 0 $X=54090 $Y=70480
X1823 1 2 531 533 20 555 533 32 ICV_30 $T=56580 95200 1 0 $X=56390 $Y=92240
X1824 1 2 552 533 30 544 508 18 ICV_30 $T=58880 84320 1 0 $X=58690 $Y=81360
X1825 1 2 550 533 17 554 533 11 ICV_30 $T=62100 89760 0 0 $X=61910 $Y=89520
X1826 1 2 581 563 34 578 563 17 ICV_30 $T=78200 95200 0 0 $X=78010 $Y=94960
X1827 1 2 592 573 33 547 508 11 ICV_30 $T=79580 84320 1 0 $X=79390 $Y=81360
X1828 1 2 639 68 32 627 68 11 ICV_30 $T=118220 111520 0 0 $X=118030 $Y=111280
X1829 1 2 687 692 11 89 90 11 ICV_30 $T=132480 57120 1 0 $X=132290 $Y=54160
X1830 1 2 690 692 32 704 90 30 ICV_30 $T=132480 62560 1 0 $X=132290 $Y=59600
X1831 1 2 689 692 34 685 658 32 ICV_30 $T=132480 68000 1 0 $X=132290 $Y=65040
X1832 1 2 682 692 17 705 658 20 ICV_30 $T=132480 73440 1 0 $X=132290 $Y=70480
X1833 1 2 707 658 11 713 700 17 ICV_30 $T=137540 89760 0 0 $X=137350 $Y=89520
X1834 1 2 726 725 18 739 725 17 ICV_30 $T=148120 68000 0 0 $X=147930 $Y=67760
X1835 1 2 737 740 32 743 740 34 ICV_30 $T=151800 106080 1 0 $X=151610 $Y=103120
X1836 1 2 752 102 18 105 102 11 ICV_30 $T=160540 51680 1 0 $X=160350 $Y=48720
X1837 1 2 751 740 33 759 734 18 ICV_30 $T=160540 100640 1 0 $X=160350 $Y=97680
X1838 1 2 758 760 32 769 748 30 ICV_30 $T=164680 73440 0 0 $X=164490 $Y=73200
X1839 1 2 778 734 34 787 734 17 ICV_30 $T=174340 84320 0 0 $X=174150 $Y=84080
X1840 1 2 783 784 11 791 784 17 ICV_30 $T=175260 95200 0 0 $X=175070 $Y=94960
X1841 1 2 113 114 30 795 114 17 ICV_30 $T=178480 51680 1 0 $X=178290 $Y=48720
X1842 1 2 786 792 34 796 792 30 ICV_30 $T=179400 73440 1 0 $X=179210 $Y=70480
X1843 1 2 803 784 33 807 784 34 ICV_30 $T=184000 100640 0 0 $X=183810 $Y=100400
X1844 1 2 805 792 32 816 817 33 ICV_30 $T=188600 78880 1 0 $X=188410 $Y=75920
X1845 1 2 828 810 18 820 810 11 ICV_30 $T=202400 62560 0 0 $X=202210 $Y=62320
X1846 1 2 831 817 32 818 817 30 ICV_30 $T=203320 78880 0 0 $X=203130 $Y=78640
X1847 1 2 832 817 34 836 817 17 ICV_30 $T=203780 84320 0 0 $X=203590 $Y=84080
X1848 1 2 850 139 34 851 139 30 ICV_30 $T=216660 62560 1 0 $X=216470 $Y=59600
X1849 1 2 844 826 17 859 856 34 ICV_30 $T=216660 73440 1 0 $X=216470 $Y=70480
X1850 1 2 872 856 17 877 856 20 ICV_30 $T=231380 68000 0 0 $X=231190 $Y=67760
X1851 1 2 916 886 193 921 886 195 ICV_30 $T=258520 78880 0 0 $X=258330 $Y=78640
X1852 1 2 199 198 187 202 198 178 ICV_30 $T=267720 111520 0 0 $X=267530 $Y=111280
X1853 1 2 950 892 195 203 201 169 ICV_30 $T=272780 57120 1 0 $X=272590 $Y=54160
X1854 1 2 980 201 180 982 201 171 ICV_30 $T=283820 57120 1 0 $X=283630 $Y=54160
X1855 1 2 1011 211 187 1010 211 170 ICV_30 $T=299000 111520 0 0 $X=298810 $Y=111280
X1856 1 2 1015 988 180 1023 1018 180 ICV_30 $T=302680 68000 0 0 $X=302490 $Y=67760
X1857 1 2 1017 1018 192 1012 212 180 ICV_30 $T=304520 57120 1 0 $X=304330 $Y=54160
X1858 1 2 1036 1018 194 1045 1018 177 ICV_30 $T=313720 57120 1 0 $X=313530 $Y=54160
X1859 1 2 1052 1053 178 1060 1053 189 ICV_30 $T=321540 106080 0 0 $X=321350 $Y=105840
X1860 1 2 1061 1053 188 1056 1053 187 ICV_30 $T=326140 95200 0 0 $X=325950 $Y=94960
X1861 1 2 1068 216 192 1075 216 180 ICV_30 $T=328900 57120 1 0 $X=328710 $Y=54160
X1862 1 2 1094 1074 170 1095 1074 189 ICV_30 $T=342700 100640 0 0 $X=342510 $Y=100400
X1863 1 2 1098 1100 195 1107 1100 180 ICV_30 $T=343620 78880 1 0 $X=343430 $Y=75920
X1864 1 2 1129 1133 191 1144 1133 189 ICV_30 $T=361560 106080 0 0 $X=361370 $Y=105840
X1865 1 2 228 226 192 1130 226 171 ICV_30 $T=362020 51680 1 0 $X=361830 $Y=48720
X1866 1 2 1146 1110 171 1161 1157 195 ICV_30 $T=370760 84320 0 0 $X=370570 $Y=84080
X1867 1 2 1166 1168 178 1174 1168 170 ICV_30 $T=376280 100640 1 0 $X=376090 $Y=97680
X1868 1 2 235 232 189 236 232 191 ICV_30 $T=382260 111520 0 0 $X=382070 $Y=111280
X1869 1 2 1182 1157 177 1185 1157 192 ICV_30 $T=386860 84320 1 0 $X=386670 $Y=81360
X1870 1 2 1217 1212 188 1225 1212 189 ICV_30 $T=403880 106080 1 0 $X=403690 $Y=103120
X1871 1 2 1247 1228 169 1273 1262 177 ICV_30 $T=426880 62560 0 0 $X=426690 $Y=62320
X1872 1 2 1218 1212 191 1263 253 182 ICV_30 $T=426880 106080 0 0 $X=426690 $Y=105840
X1873 1 2 1303 1270 191 1290 253 191 ICV_30 $T=445740 100640 0 0 $X=445550 $Y=100400
X1874 1 2 1310 1312 268 1317 252 194 ICV_30 $T=448500 57120 1 0 $X=448310 $Y=54160
X1875 1 2 1323 271 277 1330 1315 276 ICV_30 $T=454940 106080 0 0 $X=454750 $Y=105840
X1876 1 2 1327 1331 276 1336 1315 267 ICV_30 $T=455860 95200 0 0 $X=455670 $Y=94960
X1877 1 2 1320 1333 267 1337 1311 280 ICV_30 $T=456780 78880 0 0 $X=456590 $Y=78640
X1878 1 2 1348 1345 267 1352 1345 275 ICV_30 $T=467820 57120 0 0 $X=467630 $Y=56880
X1879 1 2 1354 1345 276 1349 1345 269 ICV_30 $T=469200 68000 1 0 $X=469010 $Y=65040
X1880 1 2 1347 1315 275 1363 1315 280 ICV_30 $T=471960 100640 0 0 $X=471770 $Y=100400
X1881 1 2 1390 1389 268 1388 1389 277 ICV_30 $T=488060 106080 1 0 $X=487870 $Y=103120
X1882 1 2 1435 1443 276 1434 1443 280 ICV_30 $T=511060 68000 0 0 $X=510870 $Y=67760
X1883 1 2 1445 1446 307 1452 1446 309 ICV_30 $T=514280 100640 1 0 $X=514090 $Y=97680
X1884 1 2 1462 1443 267 1470 1443 273 ICV_30 $T=520260 68000 0 0 $X=520070 $Y=67760
X1885 1 2 1454 1428 296 1474 323 309 ICV_30 $T=525320 57120 1 0 $X=525130 $Y=54160
X1886 1 2 1477 1479 277 1487 1479 269 ICV_30 $T=530380 62560 0 0 $X=530190 $Y=62320
X1887 1 2 1492 1498 273 1486 1498 277 ICV_30 $T=539120 78880 0 0 $X=538930 $Y=78640
X1888 1 2 1517 334 309 1520 1479 275 ICV_30 $T=549240 57120 0 0 $X=549050 $Y=56880
X1889 1 2 1522 1525 268 1524 1525 277 ICV_30 $T=550160 78880 0 0 $X=549970 $Y=78640
X1890 1 2 1521 1512 275 1535 1512 268 ICV_30 $T=558440 78880 0 0 $X=558250 $Y=78640
X1891 1 2 1563 1565 268 1572 1565 276 ICV_30 $T=572700 84320 1 0 $X=572510 $Y=81360
X1892 1 2 1574 340 288 1576 340 296 ICV_30 $T=581440 57120 1 0 $X=581250 $Y=54160
X1893 1 2 1585 345 273 352 345 275 ICV_30 $T=582820 111520 1 0 $X=582630 $Y=108560
X1894 1 2 1590 1565 275 1595 1565 277 ICV_30 $T=584200 68000 1 0 $X=584010 $Y=65040
X1895 1 2 1599 1601 267 1610 1601 273 ICV_30 $T=591100 89760 1 0 $X=590910 $Y=86800
X1896 1 2 1596 354 288 1618 354 296 ICV_30 $T=595240 51680 0 0 $X=595050 $Y=51440
X1897 1 2 1605 1582 273 1589 1582 275 ICV_30 $T=595240 62560 0 0 $X=595050 $Y=62320
X1898 1 2 1611 1601 276 1615 1601 280 ICV_30 $T=595240 95200 0 0 $X=595050 $Y=94960
X1899 1 2 1604 1600 280 357 358 276 ICV_30 $T=595240 111520 0 0 $X=595050 $Y=111280
X1900 1 2 1597 1582 277 1628 1625 269 ICV_30 $T=603520 62560 0 0 $X=603330 $Y=62320
X1901 1 2 1635 1612 268 1636 1625 280 ICV_30 $T=609500 73440 1 0 $X=609310 $Y=70480
X1902 1 2 1630 1612 269 1631 1612 280 ICV_30 $T=609500 84320 1 0 $X=609310 $Y=81360
X1903 1 2 1641 1625 273 1648 1625 277 ICV_30 $T=611800 62560 0 0 $X=611610 $Y=62320
X1904 1 2 1627 354 304 1647 365 296 ICV_30 $T=613180 51680 0 0 $X=612990 $Y=51440
X1905 1 2 1663 1657 276 1670 1657 280 ICV_30 $T=623760 84320 1 0 $X=623570 $Y=81360
X1906 1 2 1669 1674 269 1662 1674 277 ICV_30 $T=626520 73440 1 0 $X=626330 $Y=70480
X1907 1 2 1700 1708 267 1713 1708 280 ICV_30 $T=641700 68000 0 0 $X=641510 $Y=67760
X1908 1 2 1711 1688 267 380 381 280 ICV_30 $T=642620 106080 0 0 $X=642430 $Y=105840
X1909 1 2 1722 1701 275 1723 1697 275 ICV_30 $T=651360 89760 0 0 $X=651170 $Y=89520
X1910 1 2 1726 1709 268 1738 379 296 ICV_30 $T=653660 57120 0 0 $X=653470 $Y=56880
X1911 1 2 1727 1688 273 1742 1688 268 ICV_30 $T=654120 106080 0 0 $X=653930 $Y=105840
X1912 1 2 1764 1748 288 1787 1774 300 ICV_30 $T=684480 78880 1 0 $X=684290 $Y=75920
X1913 1 2 1823 397 296 1836 1838 304 ICV_30 $T=700120 106080 1 0 $X=699930 $Y=103120
X1914 1 2 1839 1838 300 1845 397 288 ICV_30 $T=707480 100640 0 0 $X=707290 $Y=100400
X1915 1 2 1844 1816 303 1805 1774 296 ICV_30 $T=711160 73440 0 0 $X=710970 $Y=73200
X1916 1 2 405 404 300 1877 1883 288 ICV_30 $T=723120 51680 0 0 $X=722930 $Y=51440
X1917 1 2 1870 1869 288 1880 1869 307 ICV_30 $T=723120 78880 1 0 $X=722930 $Y=75920
X1918 1 2 1871 397 307 1887 1874 288 ICV_30 $T=723580 106080 0 0 $X=723390 $Y=105840
X1919 1 2 1872 1874 304 1891 1882 288 ICV_30 $T=724960 95200 1 0 $X=724770 $Y=92240
X1920 1 2 1879 1882 309 1892 1869 296 ICV_30 $T=726800 84320 0 0 $X=726610 $Y=84080
X1921 1 2 12 13 2 470 1 sky130_fd_sc_hd__and2_1 $T=16560 57120 0 0 $X=16370 $Y=56880
X1922 1 2 16 13 2 483 1 sky130_fd_sc_hd__and2_1 $T=23000 100640 0 0 $X=22810 $Y=100400
X1923 1 2 21 13 2 479 1 sky130_fd_sc_hd__and2_1 $T=24380 73440 1 0 $X=24190 $Y=70480
X1924 1 2 15 13 2 482 1 sky130_fd_sc_hd__and2_1 $T=24380 89760 1 0 $X=24190 $Y=86800
X1925 1 2 28 13 2 485 1 sky130_fd_sc_hd__and2_1 $T=29440 73440 1 0 $X=29250 $Y=70480
X1926 1 2 36 13 2 511 1 sky130_fd_sc_hd__and2_1 $T=38180 78880 0 0 $X=37990 $Y=78640
X1927 1 2 41 13 2 514 1 sky130_fd_sc_hd__and2_1 $T=48300 57120 1 0 $X=48110 $Y=54160
X1928 1 2 46 13 2 538 1 sky130_fd_sc_hd__and2_1 $T=57500 51680 0 0 $X=57310 $Y=51440
X1929 1 2 48 13 2 556 1 sky130_fd_sc_hd__and2_1 $T=59340 84320 0 0 $X=59150 $Y=84080
X1930 1 2 49 13 2 558 1 sky130_fd_sc_hd__and2_1 $T=60260 100640 1 0 $X=60070 $Y=97680
X1931 1 2 55 13 2 56 1 sky130_fd_sc_hd__and2_1 $T=73140 111520 1 0 $X=72950 $Y=108560
X1932 1 2 58 13 2 588 1 sky130_fd_sc_hd__and2_1 $T=77280 73440 1 0 $X=77090 $Y=70480
X1933 1 2 60 13 2 590 1 sky130_fd_sc_hd__and2_1 $T=78660 57120 0 0 $X=78470 $Y=56880
X1934 1 2 61 13 2 600 1 sky130_fd_sc_hd__and2_1 $T=84180 89760 1 0 $X=83990 $Y=86800
X1935 1 2 67 69 2 612 1 sky130_fd_sc_hd__and2_1 $T=97520 111520 0 0 $X=97330 $Y=111280
X1936 1 2 71 13 2 636 1 sky130_fd_sc_hd__and2_1 $T=101660 95200 1 0 $X=101470 $Y=92240
X1937 1 2 78 13 2 646 1 sky130_fd_sc_hd__and2_1 $T=115460 57120 0 0 $X=115270 $Y=56880
X1938 1 2 79 13 2 653 1 sky130_fd_sc_hd__and2_1 $T=119600 78880 1 0 $X=119410 $Y=75920
X1939 1 2 83 13 2 681 1 sky130_fd_sc_hd__and2_1 $T=126040 51680 0 0 $X=125850 $Y=51440
X1940 1 2 84 13 2 680 1 sky130_fd_sc_hd__and2_1 $T=126040 106080 0 0 $X=125850 $Y=105840
X1941 1 2 93 13 2 706 1 sky130_fd_sc_hd__and2_1 $T=142140 68000 0 0 $X=141950 $Y=67760
X1942 1 2 94 13 2 710 1 sky130_fd_sc_hd__and2_1 $T=146280 95200 0 0 $X=146090 $Y=94960
X1943 1 2 99 13 2 729 1 sky130_fd_sc_hd__and2_1 $T=153180 84320 0 0 $X=152990 $Y=84080
X1944 1 2 100 13 2 742 1 sky130_fd_sc_hd__and2_1 $T=153640 73440 0 0 $X=153450 $Y=73200
X1945 1 2 103 13 2 736 1 sky130_fd_sc_hd__and2_1 $T=156860 95200 1 0 $X=156670 $Y=92240
X1946 1 2 104 13 2 754 1 sky130_fd_sc_hd__and2_1 $T=157780 111520 1 0 $X=157590 $Y=108560
X1947 1 2 106 13 2 773 1 sky130_fd_sc_hd__and2_1 $T=171120 68000 0 0 $X=170930 $Y=67760
X1948 1 2 108 13 2 777 1 sky130_fd_sc_hd__and2_1 $T=171580 57120 0 0 $X=171390 $Y=56880
X1949 1 2 111 13 2 781 1 sky130_fd_sc_hd__and2_1 $T=174340 111520 0 0 $X=174150 $Y=111280
X1950 1 2 115 13 2 800 1 sky130_fd_sc_hd__and2_1 $T=181700 89760 0 0 $X=181510 $Y=89520
X1951 1 2 127 13 2 827 1 sky130_fd_sc_hd__and2_1 $T=202400 68000 0 0 $X=202210 $Y=67760
X1952 1 2 134 13 2 838 1 sky130_fd_sc_hd__and2_1 $T=212060 68000 0 0 $X=211870 $Y=67760
X1953 1 2 140 13 2 840 1 sky130_fd_sc_hd__and2_1 $T=216660 57120 1 0 $X=216470 $Y=54160
X1954 1 2 22 154 2 864 1 sky130_fd_sc_hd__and2_1 $T=234140 89760 1 0 $X=233950 $Y=86800
X1955 1 2 21 154 2 882 1 sky130_fd_sc_hd__and2_1 $T=237820 62560 0 0 $X=237630 $Y=62320
X1956 1 2 15 154 2 907 1 sky130_fd_sc_hd__and2_1 $T=248860 95200 1 0 $X=248670 $Y=92240
X1957 1 2 142 152 2 919 1 sky130_fd_sc_hd__and2_1 $T=255760 95200 1 0 $X=255570 $Y=92240
X1958 1 2 43 152 2 930 1 sky130_fd_sc_hd__and2_1 $T=257600 111520 1 0 $X=257410 $Y=108560
X1959 1 2 12 154 2 200 1 sky130_fd_sc_hd__and2_1 $T=269100 57120 1 0 $X=268910 $Y=54160
X1960 1 2 61 154 2 953 1 sky130_fd_sc_hd__and2_1 $T=270020 84320 1 0 $X=269830 $Y=81360
X1961 1 2 46 154 2 979 1 sky130_fd_sc_hd__and2_1 $T=281520 57120 1 0 $X=281330 $Y=54160
X1962 1 2 48 154 2 976 1 sky130_fd_sc_hd__and2_1 $T=283820 73440 0 0 $X=283630 $Y=73200
X1963 1 2 67 152 2 987 1 sky130_fd_sc_hd__and2_1 $T=286580 89760 0 0 $X=286390 $Y=89520
X1964 1 2 153 152 2 985 1 sky130_fd_sc_hd__and2_1 $T=286580 111520 0 0 $X=286390 $Y=111280
X1965 1 2 77 154 2 998 1 sky130_fd_sc_hd__and2_1 $T=298080 68000 0 0 $X=297890 $Y=67760
X1966 1 2 133 152 2 1028 1 sky130_fd_sc_hd__and2_1 $T=308200 95200 1 0 $X=308010 $Y=92240
X1967 1 2 79 154 2 1030 1 sky130_fd_sc_hd__and2_1 $T=310500 78880 0 0 $X=310310 $Y=78640
X1968 1 2 146 152 2 1029 1 sky130_fd_sc_hd__and2_1 $T=310960 106080 0 0 $X=310770 $Y=105840
X1969 1 2 58 154 2 1059 1 sky130_fd_sc_hd__and2_1 $T=328900 68000 1 0 $X=328710 $Y=65040
X1970 1 2 60 154 2 1076 1 sky130_fd_sc_hd__and2_1 $T=331660 57120 0 0 $X=331470 $Y=56880
X1971 1 2 87 154 2 1086 1 sky130_fd_sc_hd__and2_1 $T=339020 84320 0 0 $X=338830 $Y=84080
X1972 1 2 148 152 2 1084 1 sky130_fd_sc_hd__and2_1 $T=340860 95200 1 0 $X=340670 $Y=92240
X1973 1 2 78 154 2 1123 1 sky130_fd_sc_hd__and2_1 $T=353740 57120 1 0 $X=353550 $Y=54160
X1974 1 2 106 154 2 1135 1 sky130_fd_sc_hd__and2_1 $T=362020 68000 0 0 $X=361830 $Y=67760
X1975 1 2 99 154 2 1131 1 sky130_fd_sc_hd__and2_1 $T=368460 84320 1 0 $X=368270 $Y=81360
X1976 1 2 109 154 2 1156 1 sky130_fd_sc_hd__and2_1 $T=371680 57120 1 0 $X=371490 $Y=54160
X1977 1 2 103 154 2 1172 1 sky130_fd_sc_hd__and2_1 $T=385020 95200 1 0 $X=384830 $Y=92240
X1978 1 2 93 154 2 1187 1 sky130_fd_sc_hd__and2_1 $T=395140 62560 0 0 $X=394950 $Y=62320
X1979 1 2 143 152 2 1215 1 sky130_fd_sc_hd__and2_1 $T=409400 95200 1 0 $X=409210 $Y=92240
X1980 1 2 150 152 2 1235 1 sky130_fd_sc_hd__and2_1 $T=410320 111520 1 0 $X=410130 $Y=108560
X1981 1 2 129 154 2 1231 1 sky130_fd_sc_hd__and2_1 $T=413080 78880 1 0 $X=412890 $Y=75920
X1982 1 2 132 152 2 1240 1 sky130_fd_sc_hd__and2_1 $T=413080 89760 1 0 $X=412890 $Y=86800
X1983 1 2 115 154 2 1237 1 sky130_fd_sc_hd__and2_1 $T=417680 89760 0 0 $X=417490 $Y=89520
X1984 1 2 141 154 2 251 1 sky130_fd_sc_hd__and2_1 $T=425040 51680 1 0 $X=424850 $Y=48720
X1985 1 2 260 261 2 1302 1 sky130_fd_sc_hd__and2_1 $T=445280 95200 1 0 $X=445090 $Y=92240
X1986 1 2 274 261 2 1334 1 sky130_fd_sc_hd__and2_1 $T=457700 57120 1 0 $X=457510 $Y=54160
X1987 1 2 281 261 2 1339 1 sky130_fd_sc_hd__and2_1 $T=465520 111520 1 0 $X=465330 $Y=108560
X1988 1 2 284 261 2 1340 1 sky130_fd_sc_hd__and2_1 $T=469200 84320 1 0 $X=469010 $Y=81360
X1989 1 2 291 293 2 1369 1 sky130_fd_sc_hd__and2_1 $T=476100 57120 0 0 $X=475910 $Y=56880
X1990 1 2 284 293 2 1378 1 sky130_fd_sc_hd__and2_1 $T=479320 78880 0 0 $X=479130 $Y=78640
X1991 1 2 306 293 2 1405 1 sky130_fd_sc_hd__and2_1 $T=494500 68000 1 0 $X=494310 $Y=65040
X1992 1 2 312 293 2 1416 1 sky130_fd_sc_hd__and2_1 $T=499560 100640 0 0 $X=499370 $Y=100400
X1993 1 2 314 293 2 1410 1 sky130_fd_sc_hd__and2_1 $T=504620 51680 1 0 $X=504430 $Y=48720
X1994 1 2 316 261 2 1444 1 sky130_fd_sc_hd__and2_1 $T=511060 106080 0 0 $X=510870 $Y=105840
X1995 1 2 319 293 2 1451 1 sky130_fd_sc_hd__and2_1 $T=515200 51680 1 0 $X=515010 $Y=48720
X1996 1 2 321 261 2 1458 1 sky130_fd_sc_hd__and2_1 $T=517500 78880 1 0 $X=517310 $Y=75920
X1997 1 2 317 261 2 1447 1 sky130_fd_sc_hd__and2_1 $T=525320 89760 1 0 $X=525130 $Y=86800
X1998 1 2 324 261 2 1481 1 sky130_fd_sc_hd__and2_1 $T=532680 73440 1 0 $X=532490 $Y=70480
X1999 1 2 327 261 2 1485 1 sky130_fd_sc_hd__and2_1 $T=536360 95200 0 0 $X=536170 $Y=94960
X2000 1 2 330 261 2 1504 1 sky130_fd_sc_hd__and2_1 $T=540960 84320 1 0 $X=540770 $Y=81360
X2001 1 2 332 261 2 1502 1 sky130_fd_sc_hd__and2_1 $T=545560 57120 0 0 $X=545370 $Y=56880
X2002 1 2 337 293 2 1555 1 sky130_fd_sc_hd__and2_1 $T=565800 51680 1 0 $X=565610 $Y=48720
X2003 1 2 337 261 2 1556 1 sky130_fd_sc_hd__and2_1 $T=573620 57120 0 0 $X=573430 $Y=56880
X2004 1 2 343 261 2 1571 1 sky130_fd_sc_hd__and2_1 $T=574540 106080 0 0 $X=574350 $Y=105840
X2005 1 2 289 293 2 1577 1 sky130_fd_sc_hd__and2_1 $T=578680 57120 1 0 $X=578490 $Y=54160
X2006 1 2 346 261 2 1578 1 sky130_fd_sc_hd__and2_1 $T=578680 89760 1 0 $X=578490 $Y=86800
X2007 1 2 351 261 2 1587 1 sky130_fd_sc_hd__and2_1 $T=584200 95200 0 0 $X=584010 $Y=94960
X2008 1 2 356 261 2 1617 1 sky130_fd_sc_hd__and2_1 $T=596620 73440 0 0 $X=596430 $Y=73200
X2009 1 2 360 261 2 1620 1 sky130_fd_sc_hd__and2_1 $T=603520 51680 0 0 $X=603330 $Y=51440
X2010 1 2 279 293 2 1638 1 sky130_fd_sc_hd__and2_1 $T=606740 57120 1 0 $X=606550 $Y=54160
X2011 1 2 363 261 2 1639 1 sky130_fd_sc_hd__and2_1 $T=606740 89760 1 0 $X=606550 $Y=86800
X2012 1 2 359 261 2 1621 1 sky130_fd_sc_hd__and2_1 $T=608120 100640 0 0 $X=607930 $Y=100400
X2013 1 2 368 261 2 1659 1 sky130_fd_sc_hd__and2_1 $T=623300 106080 0 0 $X=623110 $Y=105840
X2014 1 2 369 261 2 1661 1 sky130_fd_sc_hd__and2_1 $T=625140 100640 1 0 $X=624950 $Y=97680
X2015 1 2 373 261 2 1685 1 sky130_fd_sc_hd__and2_1 $T=628360 100640 0 0 $X=628170 $Y=100400
X2016 1 2 371 261 2 374 1 sky130_fd_sc_hd__and2_1 $T=628360 111520 0 0 $X=628170 $Y=111280
X2017 1 2 375 261 2 1682 1 sky130_fd_sc_hd__and2_1 $T=632040 84320 1 0 $X=631850 $Y=81360
X2018 1 2 274 293 2 1689 1 sky130_fd_sc_hd__and2_1 $T=637560 51680 1 0 $X=637370 $Y=48720
X2019 1 2 348 293 2 1744 1 sky130_fd_sc_hd__and2_1 $T=658720 111520 0 0 $X=658530 $Y=111280
X2020 1 2 356 293 2 1750 1 sky130_fd_sc_hd__and2_1 $T=661020 68000 1 0 $X=660830 $Y=65040
X2021 1 2 343 293 2 1745 1 sky130_fd_sc_hd__and2_1 $T=661020 78880 1 0 $X=660830 $Y=75920
X2022 1 2 322 293 2 1752 1 sky130_fd_sc_hd__and2_1 $T=661480 106080 1 0 $X=661290 $Y=103120
X2023 1 2 373 293 2 1761 1 sky130_fd_sc_hd__and2_1 $T=669760 100640 0 0 $X=669570 $Y=100400
X2024 1 2 308 293 2 1780 1 sky130_fd_sc_hd__and2_1 $T=676660 78880 0 0 $X=676470 $Y=78640
X2025 1 2 317 293 2 1783 1 sky130_fd_sc_hd__and2_1 $T=678500 95200 1 0 $X=678310 $Y=92240
X2026 1 2 355 293 2 392 1 sky130_fd_sc_hd__and2_1 $T=682180 51680 1 0 $X=681990 $Y=48720
X2027 1 2 363 293 2 1804 1 sky130_fd_sc_hd__and2_1 $T=690920 73440 1 0 $X=690730 $Y=70480
X2028 1 2 368 293 2 1806 1 sky130_fd_sc_hd__and2_1 $T=690920 106080 0 0 $X=690730 $Y=105840
X2029 1 2 346 293 2 1828 1 sky130_fd_sc_hd__and2_1 $T=700580 84320 0 0 $X=700390 $Y=84080
X2030 1 2 369 293 2 1841 1 sky130_fd_sc_hd__and2_1 $T=705640 100640 1 0 $X=705450 $Y=97680
X2031 1 2 375 293 2 1842 1 sky130_fd_sc_hd__and2_1 $T=708860 73440 0 0 $X=708670 $Y=73200
X2032 1 2 351 293 2 1854 1 sky130_fd_sc_hd__and2_1 $T=713460 95200 1 0 $X=713270 $Y=92240
X2033 1 2 81 479 2 452 1 sky130_fd_sc_hd__dlclkp_1 $T=19320 68000 0 0 $X=19130 $Y=67760
X2034 1 2 81 481 2 453 1 sky130_fd_sc_hd__dlclkp_1 $T=19780 78880 0 0 $X=19590 $Y=78640
X2035 1 2 81 470 2 10 1 sky130_fd_sc_hd__dlclkp_1 $T=20240 57120 1 0 $X=20050 $Y=54160
X2036 1 2 81 482 2 449 1 sky130_fd_sc_hd__dlclkp_1 $T=21160 95200 1 0 $X=20970 $Y=92240
X2037 1 2 81 483 2 454 1 sky130_fd_sc_hd__dlclkp_1 $T=21160 106080 1 0 $X=20970 $Y=103120
X2038 1 2 81 484 2 3 1 sky130_fd_sc_hd__dlclkp_1 $T=22080 111520 0 0 $X=21890 $Y=111280
X2039 1 2 81 485 2 509 1 sky130_fd_sc_hd__dlclkp_1 $T=34040 68000 1 0 $X=33850 $Y=65040
X2040 1 2 81 31 2 38 1 sky130_fd_sc_hd__dlclkp_1 $T=34040 111520 0 0 $X=33850 $Y=111280
X2041 1 2 81 511 2 510 1 sky130_fd_sc_hd__dlclkp_1 $T=37260 84320 0 0 $X=37070 $Y=84080
X2042 1 2 81 558 2 566 1 sky130_fd_sc_hd__dlclkp_1 $T=65780 106080 1 0 $X=65590 $Y=103120
X2043 1 2 81 588 2 591 1 sky130_fd_sc_hd__dlclkp_1 $T=76360 73440 0 0 $X=76170 $Y=73200
X2044 1 2 81 590 2 594 1 sky130_fd_sc_hd__dlclkp_1 $T=77280 57120 1 0 $X=77090 $Y=54160
X2045 1 2 81 600 2 607 1 sky130_fd_sc_hd__dlclkp_1 $T=83260 84320 0 0 $X=83070 $Y=84080
X2046 1 2 81 614 2 610 1 sky130_fd_sc_hd__dlclkp_1 $T=91540 111520 1 0 $X=91350 $Y=108560
X2047 1 2 81 636 2 649 1 sky130_fd_sc_hd__dlclkp_1 $T=104420 89760 1 0 $X=104230 $Y=86800
X2048 1 2 81 646 2 72 1 sky130_fd_sc_hd__dlclkp_1 $T=106260 57120 1 0 $X=106070 $Y=54160
X2049 1 2 81 653 2 629 1 sky130_fd_sc_hd__dlclkp_1 $T=109940 73440 0 0 $X=109750 $Y=73200
X2050 1 2 81 680 2 679 1 sky130_fd_sc_hd__dlclkp_1 $T=125580 111520 1 0 $X=125390 $Y=108560
X2051 1 2 81 681 2 85 1 sky130_fd_sc_hd__dlclkp_1 $T=132480 51680 1 0 $X=132290 $Y=48720
X2052 1 2 81 706 2 708 1 sky130_fd_sc_hd__dlclkp_1 $T=135700 68000 0 0 $X=135510 $Y=67760
X2053 1 2 81 710 2 678 1 sky130_fd_sc_hd__dlclkp_1 $T=139840 100640 1 0 $X=139650 $Y=97680
X2054 1 2 81 729 2 732 1 sky130_fd_sc_hd__dlclkp_1 $T=146740 84320 0 0 $X=146550 $Y=84080
X2055 1 2 81 736 2 741 1 sky130_fd_sc_hd__dlclkp_1 $T=150420 95200 1 0 $X=150230 $Y=92240
X2056 1 2 81 98 2 101 1 sky130_fd_sc_hd__dlclkp_1 $T=150420 111520 0 0 $X=150230 $Y=111280
X2057 1 2 81 742 2 738 1 sky130_fd_sc_hd__dlclkp_1 $T=153640 73440 1 0 $X=153450 $Y=70480
X2058 1 2 81 754 2 730 1 sky130_fd_sc_hd__dlclkp_1 $T=158240 111520 0 0 $X=158050 $Y=111280
X2059 1 2 81 773 2 775 1 sky130_fd_sc_hd__dlclkp_1 $T=168360 73440 1 0 $X=168170 $Y=70480
X2060 1 2 81 777 2 112 1 sky130_fd_sc_hd__dlclkp_1 $T=171120 51680 1 0 $X=170930 $Y=48720
X2061 1 2 81 781 2 776 1 sky130_fd_sc_hd__dlclkp_1 $T=171580 111520 1 0 $X=171390 $Y=108560
X2062 1 2 81 800 2 802 1 sky130_fd_sc_hd__dlclkp_1 $T=181240 89760 1 0 $X=181050 $Y=86800
X2063 1 2 81 827 2 811 1 sky130_fd_sc_hd__dlclkp_1 $T=197340 78880 1 0 $X=197150 $Y=75920
X2064 1 2 81 838 2 843 1 sky130_fd_sc_hd__dlclkp_1 $T=205620 68000 1 0 $X=205430 $Y=65040
X2065 1 2 81 840 2 837 1 sky130_fd_sc_hd__dlclkp_1 $T=207000 62560 1 0 $X=206810 $Y=59600
X2066 1 2 81 864 2 871 1 sky130_fd_sc_hd__dlclkp_1 $T=223560 84320 0 0 $X=223370 $Y=84080
X2067 1 2 81 882 2 883 1 sky130_fd_sc_hd__dlclkp_1 $T=234140 68000 1 0 $X=233950 $Y=65040
X2068 1 2 81 159 2 162 1 sky130_fd_sc_hd__dlclkp_1 $T=234600 106080 0 0 $X=234410 $Y=105840
X2069 1 2 81 907 2 909 1 sky130_fd_sc_hd__dlclkp_1 $T=245180 89760 0 0 $X=244990 $Y=89520
X2070 1 2 81 930 2 196 1 sky130_fd_sc_hd__dlclkp_1 $T=258520 111520 0 0 $X=258330 $Y=111280
X2071 1 2 81 947 2 952 1 sky130_fd_sc_hd__dlclkp_1 $T=266340 62560 0 0 $X=266150 $Y=62320
X2072 1 2 81 953 2 959 1 sky130_fd_sc_hd__dlclkp_1 $T=279220 78880 0 0 $X=279030 $Y=78640
X2073 1 2 81 985 2 207 1 sky130_fd_sc_hd__dlclkp_1 $T=284740 111520 1 0 $X=284550 $Y=108560
X2074 1 2 81 987 2 989 1 sky130_fd_sc_hd__dlclkp_1 $T=285200 95200 1 0 $X=285010 $Y=92240
X2075 1 2 81 979 2 208 1 sky130_fd_sc_hd__dlclkp_1 $T=286580 51680 0 0 $X=286390 $Y=51440
X2076 1 2 81 998 2 1009 1 sky130_fd_sc_hd__dlclkp_1 $T=293940 68000 1 0 $X=293750 $Y=65040
X2077 1 2 81 1028 2 1034 1 sky130_fd_sc_hd__dlclkp_1 $T=307740 89760 0 0 $X=307550 $Y=89520
X2078 1 2 81 1029 2 215 1 sky130_fd_sc_hd__dlclkp_1 $T=307740 111520 0 0 $X=307550 $Y=111280
X2079 1 2 81 1030 2 1033 1 sky130_fd_sc_hd__dlclkp_1 $T=308200 78880 1 0 $X=308010 $Y=75920
X2080 1 2 81 1059 2 1049 1 sky130_fd_sc_hd__dlclkp_1 $T=322460 68000 0 0 $X=322270 $Y=67760
X2081 1 2 81 1076 2 219 1 sky130_fd_sc_hd__dlclkp_1 $T=333040 51680 1 0 $X=332850 $Y=48720
X2082 1 2 81 1084 2 1078 1 sky130_fd_sc_hd__dlclkp_1 $T=334420 95200 1 0 $X=334230 $Y=92240
X2083 1 2 81 1086 2 1089 1 sky130_fd_sc_hd__dlclkp_1 $T=335800 78880 0 0 $X=335610 $Y=78640
X2084 1 2 81 1087 2 1096 1 sky130_fd_sc_hd__dlclkp_1 $T=335800 89760 0 0 $X=335610 $Y=89520
X2085 1 2 81 1105 2 1102 1 sky130_fd_sc_hd__dlclkp_1 $T=345920 68000 1 0 $X=345730 $Y=65040
X2086 1 2 81 1122 2 1124 1 sky130_fd_sc_hd__dlclkp_1 $T=352820 106080 0 0 $X=352630 $Y=105840
X2087 1 2 81 1123 2 225 1 sky130_fd_sc_hd__dlclkp_1 $T=356960 57120 1 0 $X=356770 $Y=54160
X2088 1 2 81 1131 2 1145 1 sky130_fd_sc_hd__dlclkp_1 $T=360640 78880 0 0 $X=360450 $Y=78640
X2089 1 2 81 1135 2 1148 1 sky130_fd_sc_hd__dlclkp_1 $T=364320 73440 1 0 $X=364130 $Y=70480
X2090 1 2 81 1156 2 1159 1 sky130_fd_sc_hd__dlclkp_1 $T=370300 62560 1 0 $X=370110 $Y=59600
X2091 1 2 81 1165 2 1162 1 sky130_fd_sc_hd__dlclkp_1 $T=374900 89760 0 0 $X=374710 $Y=89520
X2092 1 2 81 1187 2 1204 1 sky130_fd_sc_hd__dlclkp_1 $T=389160 68000 1 0 $X=388970 $Y=65040
X2093 1 2 81 1207 2 1188 1 sky130_fd_sc_hd__dlclkp_1 $T=398820 73440 0 0 $X=398630 $Y=73200
X2094 1 2 81 240 2 241 1 sky130_fd_sc_hd__dlclkp_1 $T=400660 51680 0 0 $X=400470 $Y=51440
X2095 1 2 81 1215 2 1205 1 sky130_fd_sc_hd__dlclkp_1 $T=402500 95200 0 0 $X=402310 $Y=94960
X2096 1 2 81 1231 2 1242 1 sky130_fd_sc_hd__dlclkp_1 $T=409400 78880 0 0 $X=409210 $Y=78640
X2097 1 2 81 1240 2 1250 1 sky130_fd_sc_hd__dlclkp_1 $T=413080 95200 1 0 $X=412890 $Y=92240
X2098 1 2 81 1235 2 1248 1 sky130_fd_sc_hd__dlclkp_1 $T=413080 111520 1 0 $X=412890 $Y=108560
X2099 1 2 81 1253 2 1256 1 sky130_fd_sc_hd__dlclkp_1 $T=417680 68000 1 0 $X=417490 $Y=65040
X2100 1 2 415 1302 2 1305 1 sky130_fd_sc_hd__dlclkp_1 $T=443900 95200 0 0 $X=443710 $Y=94960
X2101 1 2 415 1334 2 1335 1 sky130_fd_sc_hd__dlclkp_1 $T=459080 51680 0 0 $X=458890 $Y=51440
X2102 1 2 415 1339 2 263 1 sky130_fd_sc_hd__dlclkp_1 $T=460920 111520 0 0 $X=460730 $Y=111280
X2103 1 2 415 1340 2 1292 1 sky130_fd_sc_hd__dlclkp_1 $T=462300 78880 1 0 $X=462110 $Y=75920
X2104 1 2 415 1353 2 1306 1 sky130_fd_sc_hd__dlclkp_1 $T=465520 100640 0 0 $X=465330 $Y=100400
X2105 1 2 415 1378 2 1381 1 sky130_fd_sc_hd__dlclkp_1 $T=483000 73440 0 0 $X=482810 $Y=73200
X2106 1 2 415 1405 2 1409 1 sky130_fd_sc_hd__dlclkp_1 $T=490820 62560 0 0 $X=490630 $Y=62320
X2107 1 2 415 1406 2 1375 1 sky130_fd_sc_hd__dlclkp_1 $T=492660 100640 0 0 $X=492470 $Y=100400
X2108 1 2 415 1410 2 310 1 sky130_fd_sc_hd__dlclkp_1 $T=495880 51680 0 0 $X=495690 $Y=51440
X2109 1 2 415 1416 2 1436 1 sky130_fd_sc_hd__dlclkp_1 $T=504620 100640 1 0 $X=504430 $Y=97680
X2110 1 2 415 1447 2 1420 1 sky130_fd_sc_hd__dlclkp_1 $T=513820 89760 1 0 $X=513630 $Y=86800
X2111 1 2 415 1451 2 320 1 sky130_fd_sc_hd__dlclkp_1 $T=515660 51680 0 0 $X=515470 $Y=51440
X2112 1 2 415 1458 2 1418 1 sky130_fd_sc_hd__dlclkp_1 $T=517500 73440 1 0 $X=517310 $Y=70480
X2113 1 2 415 1444 2 318 1 sky130_fd_sc_hd__dlclkp_1 $T=518420 106080 1 0 $X=518230 $Y=103120
X2114 1 2 415 1481 2 1491 1 sky130_fd_sc_hd__dlclkp_1 $T=530840 73440 0 0 $X=530650 $Y=73200
X2115 1 2 415 1485 2 1500 1 sky130_fd_sc_hd__dlclkp_1 $T=532220 100640 0 0 $X=532030 $Y=100400
X2116 1 2 415 1502 2 1471 1 sky130_fd_sc_hd__dlclkp_1 $T=539120 57120 0 0 $X=538930 $Y=56880
X2117 1 2 415 1504 2 1506 1 sky130_fd_sc_hd__dlclkp_1 $T=545560 84320 0 0 $X=545370 $Y=84080
X2118 1 2 415 1555 2 336 1 sky130_fd_sc_hd__dlclkp_1 $T=567180 51680 0 0 $X=566990 $Y=51440
X2119 1 2 415 1556 2 1527 1 sky130_fd_sc_hd__dlclkp_1 $T=567180 57120 0 0 $X=566990 $Y=56880
X2120 1 2 415 1575 2 1544 1 sky130_fd_sc_hd__dlclkp_1 $T=576840 100640 0 0 $X=576650 $Y=100400
X2121 1 2 415 1578 2 1554 1 sky130_fd_sc_hd__dlclkp_1 $T=581440 89760 1 0 $X=581250 $Y=86800
X2122 1 2 415 1577 2 350 1 sky130_fd_sc_hd__dlclkp_1 $T=583280 51680 0 0 $X=583090 $Y=51440
X2123 1 2 415 1594 2 1569 1 sky130_fd_sc_hd__dlclkp_1 $T=586500 62560 1 0 $X=586310 $Y=59600
X2124 1 2 415 1617 2 1592 1 sky130_fd_sc_hd__dlclkp_1 $T=596160 78880 0 0 $X=595970 $Y=78640
X2125 1 2 415 1620 2 1616 1 sky130_fd_sc_hd__dlclkp_1 $T=599380 57120 1 0 $X=599190 $Y=54160
X2126 1 2 415 1621 2 1591 1 sky130_fd_sc_hd__dlclkp_1 $T=600760 106080 0 0 $X=600570 $Y=105840
X2127 1 2 415 1639 2 1637 1 sky130_fd_sc_hd__dlclkp_1 $T=609500 89760 1 0 $X=609310 $Y=86800
X2128 1 2 415 1659 2 1664 1 sky130_fd_sc_hd__dlclkp_1 $T=616400 106080 0 0 $X=616210 $Y=105840
X2129 1 2 415 1661 2 1640 1 sky130_fd_sc_hd__dlclkp_1 $T=618700 100640 1 0 $X=618510 $Y=97680
X2130 1 2 415 1685 2 1695 1 sky130_fd_sc_hd__dlclkp_1 $T=628820 100640 1 0 $X=628630 $Y=97680
X2131 1 2 415 1689 2 376 1 sky130_fd_sc_hd__dlclkp_1 $T=630660 51680 1 0 $X=630470 $Y=48720
X2132 1 2 415 1745 2 1753 1 sky130_fd_sc_hd__dlclkp_1 $T=658720 78880 0 0 $X=658530 $Y=78640
X2133 1 2 415 1750 2 1736 1 sky130_fd_sc_hd__dlclkp_1 $T=660560 62560 0 0 $X=660370 $Y=62320
X2134 1 2 415 1752 2 1731 1 sky130_fd_sc_hd__dlclkp_1 $T=660560 100640 0 0 $X=660370 $Y=100400
X2135 1 2 415 1761 2 1776 1 sky130_fd_sc_hd__dlclkp_1 $T=670220 100640 1 0 $X=670030 $Y=97680
X2136 1 2 415 1783 2 1781 1 sky130_fd_sc_hd__dlclkp_1 $T=679420 89760 0 0 $X=679230 $Y=89520
X2137 1 2 415 1804 2 1808 1 sky130_fd_sc_hd__dlclkp_1 $T=693680 78880 1 0 $X=693490 $Y=75920
X2138 1 2 415 1806 2 1817 1 sky130_fd_sc_hd__dlclkp_1 $T=693680 106080 1 0 $X=693490 $Y=103120
X2139 1 2 415 1828 2 1819 1 sky130_fd_sc_hd__dlclkp_1 $T=700580 89760 0 0 $X=700390 $Y=89520
X2140 1 2 415 1841 2 1865 1 sky130_fd_sc_hd__dlclkp_1 $T=711620 95200 0 0 $X=711430 $Y=94960
X2141 1 2 415 1842 2 1867 1 sky130_fd_sc_hd__dlclkp_1 $T=714380 78880 1 0 $X=714190 $Y=75920
X2142 1 2 415 401 2 402 1 sky130_fd_sc_hd__dlclkp_1 $T=714840 51680 1 0 $X=714650 $Y=48720
X2143 1 2 415 1854 2 1868 1 sky130_fd_sc_hd__dlclkp_1 $T=716680 89760 0 0 $X=716490 $Y=89520
X2144 1 2 ICV_32 $T=29900 111520 0 0 $X=29710 $Y=111280
X2145 1 2 ICV_32 $T=72220 106080 1 0 $X=72030 $Y=103120
X2146 1 2 ICV_32 $T=128340 73440 1 0 $X=128150 $Y=70480
X2147 1 2 ICV_32 $T=156400 100640 1 0 $X=156210 $Y=97680
X2148 1 2 ICV_32 $T=212520 73440 1 0 $X=212330 $Y=70480
X2149 1 2 ICV_32 $T=212520 111520 1 0 $X=212330 $Y=108560
X2150 1 2 ICV_32 $T=268640 62560 1 0 $X=268450 $Y=59600
X2151 1 2 ICV_32 $T=268640 111520 1 0 $X=268450 $Y=108560
X2152 1 2 ICV_32 $T=282440 100640 0 0 $X=282250 $Y=100400
X2153 1 2 ICV_32 $T=296700 106080 1 0 $X=296510 $Y=103120
X2154 1 2 ICV_32 $T=478860 51680 0 0 $X=478670 $Y=51440
X2155 1 2 ICV_32 $T=549240 51680 1 0 $X=549050 $Y=48720
X2156 1 2 ICV_32 $T=577300 73440 1 0 $X=577110 $Y=70480
X2157 1 2 ICV_32 $T=675280 62560 0 0 $X=675090 $Y=62320
X2158 1 2 ICV_32 $T=675280 106080 0 0 $X=675090 $Y=105840
X2159 1 2 ICV_32 $T=731400 51680 0 0 $X=731210 $Y=51440
X2160 1 2 453 8 471 ICV_35 $T=10580 78880 1 0 $X=10390 $Y=75920
X2161 1 2 449 8 472 ICV_35 $T=10580 89760 1 0 $X=10390 $Y=86800
X2162 1 2 454 24 497 ICV_35 $T=25300 100640 0 0 $X=25110 $Y=100400
X2163 1 2 10 27 501 ICV_35 $T=26680 57120 1 0 $X=26490 $Y=54160
X2164 1 2 510 25 522 ICV_35 $T=38180 84320 1 0 $X=37990 $Y=81360
X2165 1 2 512 25 528 ICV_35 $T=39560 95200 1 0 $X=39370 $Y=92240
X2166 1 2 566 8 601 ICV_35 $T=78200 100640 0 0 $X=78010 $Y=100400
X2167 1 2 607 4 613 ICV_35 $T=86480 89760 1 0 $X=86290 $Y=86800
X2168 1 2 607 27 617 ICV_35 $T=87860 78880 1 0 $X=87670 $Y=75920
X2169 1 2 649 8 641 ICV_35 $T=108560 95200 1 0 $X=108370 $Y=92240
X2170 1 2 675 27 686 ICV_35 $T=121440 84320 1 0 $X=121250 $Y=81360
X2171 1 2 671 6 688 ICV_35 $T=122360 57120 0 0 $X=122170 $Y=56880
X2172 1 2 675 24 657 ICV_35 $T=122360 84320 0 0 $X=122170 $Y=84080
X2173 1 2 730 25 751 ICV_35 $T=150420 100640 0 0 $X=150230 $Y=100400
X2174 1 2 730 5 766 ICV_35 $T=160540 106080 1 0 $X=160350 $Y=103120
X2175 1 2 776 6 801 ICV_35 $T=176640 111520 0 0 $X=176450 $Y=111280
X2176 1 2 776 24 808 ICV_35 $T=179400 106080 1 0 $X=179210 $Y=103120
X2177 1 2 843 6 852 ICV_35 $T=210680 62560 0 0 $X=210490 $Y=62320
X2178 1 2 162 158 906 ICV_35 $T=238280 111520 0 0 $X=238090 $Y=111280
X2179 1 2 162 175 190 ICV_35 $T=247940 111520 0 0 $X=247750 $Y=111280
X2180 1 2 161 184 927 ICV_35 $T=250700 51680 1 0 $X=250510 $Y=48720
X2181 1 2 883 184 931 ICV_35 $T=253460 57120 1 0 $X=253270 $Y=54160
X2182 1 2 926 175 971 ICV_35 $T=272780 100640 1 0 $X=272590 $Y=97680
X2183 1 2 959 183 974 ICV_35 $T=276920 95200 1 0 $X=276730 $Y=92240
X2184 1 2 208 167 1012 ICV_35 $T=292100 57120 1 0 $X=291910 $Y=54160
X2185 1 2 1034 156 1046 ICV_35 $T=310500 95200 1 0 $X=310310 $Y=92240
X2186 1 2 1034 181 1060 ICV_35 $T=316480 106080 1 0 $X=316290 $Y=103120
X2187 1 2 1049 184 1070 ICV_35 $T=322000 57120 0 0 $X=321810 $Y=56880
X2188 1 2 1078 156 1094 ICV_35 $T=333040 100640 1 0 $X=332850 $Y=97680
X2189 1 2 1078 157 1112 ICV_35 $T=342700 106080 0 0 $X=342510 $Y=105840
X2190 1 2 1089 185 1125 ICV_35 $T=348220 73440 1 0 $X=348030 $Y=70480
X2191 1 2 220 158 227 ICV_35 $T=350060 111520 0 0 $X=349870 $Y=111280
X2192 1 2 1102 168 1140 ICV_35 $T=356960 68000 1 0 $X=356770 $Y=65040
X2193 1 2 1096 185 1147 ICV_35 $T=360180 89760 0 0 $X=359990 $Y=89520
X2194 1 2 225 186 1152 ICV_35 $T=363400 57120 1 0 $X=363210 $Y=54160
X2195 1 2 1162 157 1166 ICV_35 $T=374440 106080 1 0 $X=374250 $Y=103120
X2196 1 2 1145 164 1179 ICV_35 $T=376280 78880 1 0 $X=376090 $Y=75920
X2197 1 2 1159 184 1194 ICV_35 $T=385020 51680 1 0 $X=384830 $Y=48720
X2198 1 2 1188 186 1234 ICV_35 $T=404340 73440 1 0 $X=404150 $Y=70480
X2199 1 2 1248 173 1290 ICV_35 $T=432400 106080 1 0 $X=432210 $Y=103120
X2200 1 2 1304 257 1321 ICV_35 $T=446200 84320 0 0 $X=446010 $Y=84080
X2201 1 2 1305 264 1327 ICV_35 $T=447580 95200 1 0 $X=447390 $Y=92240
X2202 1 2 1304 265 1377 ICV_35 $T=472420 84320 0 0 $X=472230 $Y=84080
X2203 1 2 310 301 1433 ICV_35 $T=502320 51680 0 0 $X=502130 $Y=51440
X2204 1 2 310 305 1442 ICV_35 $T=506920 51680 1 0 $X=506730 $Y=48720
X2205 1 2 1436 292 1450 ICV_35 $T=508760 95200 1 0 $X=508570 $Y=92240
X2206 1 2 1409 305 1455 ICV_35 $T=511060 62560 0 0 $X=510870 $Y=62320
X2207 1 2 318 266 1482 ICV_35 $T=525320 111520 1 0 $X=525130 $Y=108560
X2208 1 2 1473 264 1488 ICV_35 $T=527620 84320 0 0 $X=527430 $Y=84080
X2209 1 2 1473 272 1489 ICV_35 $T=527620 89760 1 0 $X=527430 $Y=86800
X2210 1 2 1544 258 1561 ICV_35 $T=564420 95200 1 0 $X=564230 $Y=92240
X2211 1 2 338 257 341 ICV_35 $T=565340 111520 1 0 $X=565150 $Y=108560
X2212 1 2 1527 265 1567 ICV_35 $T=567180 62560 0 0 $X=566990 $Y=62320
X2213 1 2 1554 257 1563 ICV_35 $T=567180 73440 0 0 $X=566990 $Y=73200
X2214 1 2 1544 272 1579 ICV_35 $T=572700 95200 1 0 $X=572510 $Y=92240
X2215 1 2 1569 272 1583 ICV_35 $T=575460 73440 0 0 $X=575270 $Y=73200
X2216 1 2 1591 264 1603 ICV_35 $T=585580 106080 0 0 $X=585390 $Y=105840
X2217 1 2 1592 266 1609 ICV_35 $T=586500 84320 0 0 $X=586310 $Y=84080
X2218 1 2 1593 264 1611 ICV_35 $T=586500 95200 0 0 $X=586310 $Y=94960
X2219 1 2 1593 272 1615 ICV_35 $T=588800 100640 1 0 $X=588610 $Y=97680
X2220 1 2 1592 257 1635 ICV_35 $T=598920 78880 1 0 $X=598730 $Y=75920
X2221 1 2 361 257 367 ICV_35 $T=603520 111520 0 0 $X=603330 $Y=111280
X2222 1 2 1664 266 1687 ICV_35 $T=625600 106080 0 0 $X=625410 $Y=105840
X2223 1 2 376 292 1719 ICV_35 $T=639860 51680 1 0 $X=639670 $Y=48720
X2224 1 2 1695 265 1723 ICV_35 $T=642620 95200 0 0 $X=642430 $Y=94960
X2225 1 2 1694 257 1726 ICV_35 $T=644920 57120 1 0 $X=644730 $Y=54160
X2226 1 2 1736 287 1755 ICV_35 $T=656880 57120 1 0 $X=656690 $Y=54160
X2227 1 2 402 287 408 ICV_35 $T=729100 51680 1 0 $X=728910 $Y=48720
X2228 1 2 509 8 541 ICV_37 $T=47840 68000 1 0 $X=47650 $Y=65040
X2229 1 2 45 8 52 ICV_37 $T=61640 51680 0 0 $X=61450 $Y=51440
X2230 1 2 540 26 551 ICV_37 $T=61640 68000 0 0 $X=61450 $Y=67760
X2231 1 2 560 25 592 ICV_37 $T=75900 89760 1 0 $X=75710 $Y=86800
X2232 1 2 607 26 619 ICV_37 $T=89700 73440 0 0 $X=89510 $Y=73200
X2233 1 2 607 5 620 ICV_37 $T=89700 78880 0 0 $X=89510 $Y=78640
X2234 1 2 610 27 621 ICV_37 $T=89700 89760 0 0 $X=89510 $Y=89520
X2235 1 2 72 4 75 ICV_37 $T=103960 51680 1 0 $X=103770 $Y=48720
X2236 1 2 629 4 631 ICV_37 $T=103960 68000 1 0 $X=103770 $Y=65040
X2237 1 2 629 27 647 ICV_37 $T=103960 73440 1 0 $X=103770 $Y=70480
X2238 1 2 633 24 642 ICV_37 $T=103960 106080 1 0 $X=103770 $Y=103120
X2239 1 2 633 25 650 ICV_37 $T=103960 111520 1 0 $X=103770 $Y=108560
X2240 1 2 633 27 677 ICV_37 $T=117760 100640 0 0 $X=117570 $Y=100400
X2241 1 2 633 5 673 ICV_37 $T=117760 106080 0 0 $X=117570 $Y=105840
X2242 1 2 679 26 683 ICV_37 $T=132020 100640 1 0 $X=131830 $Y=97680
X2243 1 2 708 24 728 ICV_37 $T=145820 62560 0 0 $X=145630 $Y=62320
X2244 1 2 708 5 739 ICV_37 $T=145820 73440 0 0 $X=145630 $Y=73200
X2245 1 2 738 25 765 ICV_37 $T=160080 73440 1 0 $X=159890 $Y=70480
X2246 1 2 741 6 759 ICV_37 $T=160080 95200 1 0 $X=159890 $Y=92240
X2247 1 2 730 6 762 ICV_37 $T=160080 111520 1 0 $X=159890 $Y=108560
X2248 1 2 776 5 791 ICV_37 $T=173880 100640 0 0 $X=173690 $Y=100400
X2249 1 2 776 4 788 ICV_37 $T=173880 106080 0 0 $X=173690 $Y=105840
X2250 1 2 790 8 820 ICV_37 $T=188140 57120 1 0 $X=187950 $Y=54160
X2251 1 2 802 25 816 ICV_37 $T=188140 84320 1 0 $X=187950 $Y=81360
X2252 1 2 847 25 861 ICV_37 $T=216200 78880 1 0 $X=216010 $Y=75920
X2253 1 2 847 6 858 ICV_37 $T=216200 84320 1 0 $X=216010 $Y=81360
X2254 1 2 843 26 880 ICV_37 $T=230000 62560 0 0 $X=229810 $Y=62320
X2255 1 2 881 175 911 ICV_37 $T=244260 100640 1 0 $X=244070 $Y=97680
X2256 1 2 909 184 938 ICV_37 $T=258060 84320 0 0 $X=257870 $Y=84080
X2257 1 2 909 186 933 ICV_37 $T=258060 89760 0 0 $X=257870 $Y=89520
X2258 1 2 928 184 966 ICV_37 $T=272320 78880 1 0 $X=272130 $Y=75920
X2259 1 2 1009 183 1019 ICV_37 $T=300380 62560 1 0 $X=300190 $Y=59600
X2260 1 2 1009 167 1023 ICV_37 $T=300380 68000 1 0 $X=300190 $Y=65040
X2261 1 2 984 168 1021 ICV_37 $T=300380 73440 1 0 $X=300190 $Y=70480
X2262 1 2 984 184 1022 ICV_37 $T=300380 78880 1 0 $X=300190 $Y=75920
X2263 1 2 989 158 1024 ICV_37 $T=300380 95200 1 0 $X=300190 $Y=92240
X2264 1 2 1009 168 1045 ICV_37 $T=314180 57120 0 0 $X=313990 $Y=56880
X2265 1 2 1009 166 1047 ICV_37 $T=314180 62560 0 0 $X=313990 $Y=62320
X2266 1 2 1033 167 1050 ICV_37 $T=314180 73440 0 0 $X=313990 $Y=73200
X2267 1 2 1089 167 1107 ICV_37 $T=342240 73440 0 0 $X=342050 $Y=73200
X2268 1 2 220 160 223 ICV_37 $T=342240 111520 0 0 $X=342050 $Y=111280
X2269 1 2 1096 183 1137 ICV_37 $T=356500 89760 1 0 $X=356310 $Y=86800
X2270 1 2 1124 165 1138 ICV_37 $T=356500 100640 1 0 $X=356310 $Y=97680
X2271 1 2 1124 157 1139 ICV_37 $T=356500 106080 1 0 $X=356310 $Y=103120
X2272 1 2 220 156 1121 ICV_37 $T=356500 111520 1 0 $X=356310 $Y=108560
X2273 1 2 1148 183 1167 ICV_37 $T=370300 62560 0 0 $X=370110 $Y=62320
X2274 1 2 1145 185 1154 ICV_37 $T=370300 73440 0 0 $X=370110 $Y=73200
X2275 1 2 1145 166 1169 ICV_37 $T=370300 78880 0 0 $X=370110 $Y=78640
X2276 1 2 1124 173 1129 ICV_37 $T=370300 106080 0 0 $X=370110 $Y=105840
X2277 1 2 1145 183 1186 ICV_37 $T=384560 78880 1 0 $X=384370 $Y=75920
X2278 1 2 1204 185 1221 ICV_37 $T=398360 57120 0 0 $X=398170 $Y=56880
X2279 1 2 1180 185 1223 ICV_37 $T=398360 78880 0 0 $X=398170 $Y=78640
X2280 1 2 1205 165 1217 ICV_37 $T=398360 100640 0 0 $X=398170 $Y=100400
X2281 1 2 1205 181 1225 ICV_37 $T=398360 106080 0 0 $X=398170 $Y=105840
X2282 1 2 1204 166 1252 ICV_37 $T=412620 62560 1 0 $X=412430 $Y=59600
X2283 1 2 1205 175 1245 ICV_37 $T=412620 100640 1 0 $X=412430 $Y=97680
X2284 1 2 249 184 1277 ICV_37 $T=426420 51680 0 0 $X=426230 $Y=51440
X2285 1 2 1256 167 1274 ICV_37 $T=426420 57120 0 0 $X=426230 $Y=56880
X2286 1 2 1292 259 1308 ICV_37 $T=440680 73440 1 0 $X=440490 $Y=70480
X2287 1 2 1250 173 1303 ICV_37 $T=440680 100640 1 0 $X=440490 $Y=97680
X2288 1 2 1304 266 1338 ICV_37 $T=454480 84320 0 0 $X=454290 $Y=84080
X2289 1 2 1306 259 1336 ICV_37 $T=454480 100640 0 0 $X=454290 $Y=100400
X2290 1 2 1305 265 1366 ICV_37 $T=468740 89760 1 0 $X=468550 $Y=86800
X2291 1 2 1305 272 1362 ICV_37 $T=468740 95200 1 0 $X=468550 $Y=92240
X2292 1 2 1306 258 1365 ICV_37 $T=468740 106080 1 0 $X=468550 $Y=103120
X2293 1 2 263 264 1356 ICV_37 $T=468740 111520 1 0 $X=468550 $Y=108560
X2294 1 2 1301 266 1373 ICV_37 $T=482540 68000 0 0 $X=482350 $Y=67760
X2295 1 2 1382 287 1392 ICV_37 $T=482540 89760 0 0 $X=482350 $Y=89520
X2296 1 2 1375 257 1390 ICV_37 $T=482540 100640 0 0 $X=482350 $Y=100400
X2297 1 2 290 297 1383 ICV_37 $T=482540 111520 0 0 $X=482350 $Y=111280
X2298 1 2 310 299 313 ICV_37 $T=496800 51680 1 0 $X=496610 $Y=48720
X2299 1 2 1382 305 1423 ICV_37 $T=496800 89760 1 0 $X=496610 $Y=86800
X2300 1 2 1375 259 1417 ICV_37 $T=496800 100640 1 0 $X=496610 $Y=97680
X2301 1 2 1375 265 1419 ICV_37 $T=496800 111520 1 0 $X=496610 $Y=108560
X2302 1 2 1436 299 1445 ICV_37 $T=510600 89760 0 0 $X=510410 $Y=89520
X2303 1 2 1436 302 1452 ICV_37 $T=510600 100640 0 0 $X=510410 $Y=100400
X2304 1 2 1418 259 1462 ICV_37 $T=524860 73440 1 0 $X=524670 $Y=70480
X2305 1 2 1491 266 1508 ICV_37 $T=538660 68000 0 0 $X=538470 $Y=67760
X2306 1 2 331 297 1534 ICV_37 $T=552920 57120 1 0 $X=552730 $Y=54160
X2307 1 2 1500 266 1538 ICV_37 $T=552920 100640 1 0 $X=552730 $Y=97680
X2308 1 2 1500 264 1532 ICV_37 $T=552920 106080 1 0 $X=552730 $Y=103120
X2309 1 2 1527 264 1564 ICV_37 $T=566720 68000 0 0 $X=566530 $Y=67760
X2310 1 2 1544 257 1547 ICV_37 $T=566720 95200 0 0 $X=566530 $Y=94960
X2311 1 2 1544 266 1560 ICV_37 $T=566720 100640 0 0 $X=566530 $Y=100400
X2312 1 2 338 272 342 ICV_37 $T=566720 106080 0 0 $X=566530 $Y=105840
X2313 1 2 364 287 1647 ICV_37 $T=609040 51680 1 0 $X=608850 $Y=48720
X2314 1 2 1616 262 1641 ICV_37 $T=609040 62560 1 0 $X=608850 $Y=59600
X2315 1 2 1616 266 1648 ICV_37 $T=609040 68000 1 0 $X=608850 $Y=65040
X2316 1 2 1637 258 1675 ICV_37 $T=622840 84320 0 0 $X=622650 $Y=84080
X2317 1 2 1694 259 1707 ICV_37 $T=637100 57120 1 0 $X=636910 $Y=54160
X2318 1 2 1692 272 1713 ICV_37 $T=637100 73440 1 0 $X=636910 $Y=70480
X2319 1 2 1690 266 1715 ICV_37 $T=637100 84320 1 0 $X=636910 $Y=81360
X2320 1 2 1690 272 1716 ICV_37 $T=637100 89760 1 0 $X=636910 $Y=86800
X2321 1 2 1695 264 1710 ICV_37 $T=637100 95200 1 0 $X=636910 $Y=92240
X2322 1 2 1695 259 1717 ICV_37 $T=637100 100640 1 0 $X=636910 $Y=97680
X2323 1 2 1664 259 1711 ICV_37 $T=637100 106080 1 0 $X=636910 $Y=103120
X2324 1 2 376 287 1738 ICV_37 $T=650900 51680 0 0 $X=650710 $Y=51440
X2325 1 2 1694 258 1733 ICV_37 $T=650900 62560 0 0 $X=650710 $Y=62320
X2326 1 2 1690 262 1729 ICV_37 $T=650900 78880 0 0 $X=650710 $Y=78640
X2327 1 2 1695 257 1741 ICV_37 $T=650900 100640 0 0 $X=650710 $Y=100400
X2328 1 2 377 258 382 ICV_37 $T=650900 111520 0 0 $X=650710 $Y=111280
X2329 1 2 1731 287 1765 ICV_37 $T=665160 89760 1 0 $X=664970 $Y=86800
X2330 1 2 1781 292 1787 ICV_37 $T=678960 78880 0 0 $X=678770 $Y=78640
X2331 1 2 1781 305 1788 ICV_37 $T=678960 84320 0 0 $X=678770 $Y=84080
X2332 1 2 1808 305 1821 ICV_37 $T=693220 73440 1 0 $X=693030 $Y=70480
X2333 1 2 402 297 406 ICV_37 $T=721280 51680 1 0 $X=721090 $Y=48720
X2334 1 2 1866 302 1884 ICV_37 $T=721280 57120 1 0 $X=721090 $Y=54160
X2335 1 2 1866 292 1881 ICV_37 $T=721280 62560 1 0 $X=721090 $Y=59600
X2336 1 2 1867 292 1885 ICV_37 $T=721280 73440 1 0 $X=721090 $Y=70480
X2337 1 2 1868 302 1879 ICV_37 $T=721280 84320 1 0 $X=721090 $Y=81360
X2338 1 2 1868 297 1889 ICV_37 $T=721280 89760 1 0 $X=721090 $Y=86800
X2339 1 2 1865 297 1890 ICV_37 $T=721280 100640 1 0 $X=721090 $Y=97680
X2340 1 2 1865 305 1887 ICV_37 $T=721280 106080 1 0 $X=721090 $Y=103120
X2341 1 2 403 297 1861 ICV_37 $T=721280 111520 1 0 $X=721090 $Y=108560
X2342 1 2 1866 299 1895 ICV_37 $T=735080 57120 0 0 $X=734890 $Y=56880
X2343 1 2 1866 301 1898 ICV_37 $T=735080 62560 0 0 $X=734890 $Y=62320
X2344 1 2 1867 283 1899 ICV_37 $T=735080 68000 0 0 $X=734890 $Y=67760
X2345 1 2 1867 287 1892 ICV_37 $T=735080 78880 0 0 $X=734890 $Y=78640
X2346 1 2 1868 299 1903 ICV_37 $T=735080 84320 0 0 $X=734890 $Y=84080
X2347 1 2 1868 287 1901 ICV_37 $T=735080 89760 0 0 $X=734890 $Y=89520
X2348 1 2 1865 283 1904 ICV_37 $T=735080 95200 0 0 $X=734890 $Y=94960
X2349 1 2 1865 299 1905 ICV_37 $T=735080 100640 0 0 $X=734890 $Y=100400
X2350 1 2 403 287 1823 ICV_37 $T=735080 111520 0 0 $X=734890 $Y=111280
X2351 1 2 510 5 524 510 26 507 ICV_38 $T=39560 73440 0 0 $X=39370 $Y=73200
X2352 1 2 678 26 714 678 8 712 ICV_38 $T=136620 89760 1 0 $X=136430 $Y=86800
X2353 1 2 730 26 737 741 26 733 ICV_38 $T=148580 95200 0 0 $X=148390 $Y=94960
X2354 1 2 738 27 757 738 24 774 ICV_38 $T=156860 57120 0 0 $X=156670 $Y=56880
X2355 1 2 776 26 789 776 27 807 ICV_38 $T=172500 100640 1 0 $X=172310 $Y=97680
X2356 1 2 775 24 796 790 5 812 ICV_38 $T=175720 62560 0 0 $X=175530 $Y=62320
X2357 1 2 847 5 874 847 24 869 ICV_38 $T=224020 84320 1 0 $X=223830 $Y=81360
X2358 1 2 843 8 868 843 24 878 ICV_38 $T=224940 73440 1 0 $X=224750 $Y=70480
X2359 1 2 909 168 955 909 185 956 ICV_38 $T=265880 89760 0 0 $X=265690 $Y=89520
X2360 1 2 214 168 1043 214 166 1062 ICV_38 $T=310960 51680 1 0 $X=310770 $Y=48720
X2361 1 2 1033 183 1044 1033 168 1057 ICV_38 $T=310960 73440 1 0 $X=310770 $Y=70480
X2362 1 2 225 166 1130 225 168 1150 ICV_38 $T=355580 51680 0 0 $X=355390 $Y=51440
X2363 1 2 1124 158 1132 1124 156 1151 ICV_38 $T=355580 95200 0 0 $X=355390 $Y=94960
X2364 1 2 1250 158 1266 1250 165 1272 ICV_38 $T=419520 95200 1 0 $X=419330 $Y=92240
X2365 1 2 1301 264 1318 1301 259 1324 ICV_38 $T=446200 68000 1 0 $X=446010 $Y=65040
X2366 1 2 1335 265 1352 1335 272 1361 ICV_38 $T=460460 62560 0 0 $X=460270 $Y=62320
X2367 1 2 320 302 1474 320 301 326 ICV_38 $T=522100 51680 0 0 $X=521910 $Y=51440
X2368 1 2 350 305 1596 350 287 1618 ICV_38 $T=584200 51680 1 0 $X=584010 $Y=48720
X2369 1 2 1591 262 1614 1591 266 1598 ICV_38 $T=588340 106080 1 0 $X=588150 $Y=103120
X2370 1 2 1637 266 1645 1637 264 1663 ICV_38 $T=608120 84320 0 0 $X=607930 $Y=84080
X2371 1 2 1664 262 1727 1664 257 1742 ICV_38 $T=646760 106080 1 0 $X=646570 $Y=103120
X2372 1 2 1776 292 1784 1776 297 1801 ICV_38 $T=676660 100640 1 0 $X=676470 $Y=97680
X2373 1 2 456 14 17 ICV_39 $T=17020 111520 0 0 $X=16830 $Y=111280
X2374 1 2 488 476 32 ICV_39 $T=34040 68000 0 0 $X=33850 $Y=67760
X2375 1 2 522 508 33 ICV_39 $T=45540 84320 0 0 $X=45350 $Y=84080
X2376 1 2 619 615 32 ICV_39 $T=108560 84320 0 0 $X=108370 $Y=84080
X2377 1 2 648 644 11 ICV_39 $T=112700 111520 0 0 $X=112510 $Y=111280
X2378 1 2 676 80 17 ICV_39 $T=126960 51680 1 0 $X=126770 $Y=48720
X2379 1 2 684 658 18 ICV_39 $T=132480 78880 1 0 $X=132290 $Y=75920
X2380 1 2 714 700 32 ICV_39 $T=144440 84320 1 0 $X=144250 $Y=81360
X2381 1 2 866 139 11 ICV_39 $T=231840 57120 1 0 $X=231650 $Y=54160
X2382 1 2 896 886 169 ICV_39 $T=259900 84320 1 0 $X=259710 $Y=81360
X2383 1 2 938 923 192 ICV_39 $T=264960 84320 1 0 $X=264770 $Y=81360
X2384 1 2 1044 1039 193 ICV_39 $T=317400 68000 0 0 $X=317210 $Y=67760
X2385 1 2 1063 1038 177 ICV_39 $T=328900 84320 1 0 $X=328710 $Y=81360
X2386 1 2 224 221 194 ICV_39 $T=350060 51680 1 0 $X=349870 $Y=48720
X2387 1 2 1151 1133 170 ICV_39 $T=371220 95200 1 0 $X=371030 $Y=92240
X2388 1 2 1169 1157 171 ICV_39 $T=379500 73440 1 0 $X=379310 $Y=70480
X2389 1 2 1257 1246 193 ICV_39 $T=421360 89760 0 0 $X=421170 $Y=89520
X2390 1 2 1286 1262 192 ICV_39 $T=441140 68000 1 0 $X=440950 $Y=65040
X2391 1 2 1307 1311 268 ICV_39 $T=449420 68000 0 0 $X=449230 $Y=67760
X2392 1 2 1356 271 276 ICV_39 $T=470120 111520 0 0 $X=469930 $Y=111280
X2393 1 2 1407 1389 276 ICV_39 $T=497260 106080 1 0 $X=497070 $Y=103120
X2394 1 2 1459 1443 268 ICV_39 $T=519800 78880 1 0 $X=519610 $Y=75920
X2395 1 2 1456 1446 294 ICV_39 $T=519800 95200 1 0 $X=519610 $Y=92240
X2396 1 2 1503 1498 268 ICV_39 $T=541420 95200 1 0 $X=541230 $Y=92240
X2397 1 2 1497 323 296 ICV_39 $T=543720 57120 1 0 $X=543530 $Y=54160
X2398 1 2 1505 1512 267 ICV_39 $T=547860 73440 1 0 $X=547670 $Y=70480
X2399 1 2 1518 1513 280 ICV_39 $T=552460 100640 0 0 $X=552270 $Y=100400
X2400 1 2 1531 1513 268 ICV_39 $T=557520 100640 0 0 $X=557330 $Y=100400
X2401 1 2 1561 1551 269 ICV_39 $T=571780 89760 0 0 $X=571590 $Y=89520
X2402 1 2 1584 1551 273 ICV_39 $T=582820 95200 1 0 $X=582630 $Y=92240
X2403 1 2 1634 1625 276 ICV_39 $T=610420 68000 0 0 $X=610230 $Y=67760
X2404 1 2 1649 1600 268 ICV_39 $T=621000 111520 1 0 $X=620810 $Y=108560
X2405 1 2 1733 1709 269 ICV_39 $T=655960 68000 1 0 $X=655770 $Y=65040
X2406 1 2 1834 1800 296 ICV_39 $T=708400 95200 1 0 $X=708210 $Y=92240
X2407 1 2 1890 1874 303 ICV_39 $T=730020 95200 0 0 $X=729830 $Y=94960
X2408 1 2 1895 1883 307 ICV_39 $T=737840 51680 0 0 $X=737650 $Y=51440
X2409 1 2 1898 1883 304 ICV_39 $T=737840 68000 1 0 $X=737650 $Y=65040
X2410 1 2 1899 1869 294 ICV_39 $T=737840 73440 0 0 $X=737650 $Y=73200
X2411 1 2 1902 1874 296 ICV_39 $T=737840 106080 0 0 $X=737650 $Y=105840
X2412 1 2 492 477 32 ICV_40 $T=32660 78880 1 0 $X=32470 $Y=75920
X2413 1 2 567 53 34 ICV_40 $T=69920 51680 1 0 $X=69730 $Y=48720
X2414 1 2 570 573 34 ICV_40 $T=69920 84320 1 0 $X=69730 $Y=81360
X2415 1 2 620 615 17 ICV_40 $T=96600 84320 1 0 $X=96410 $Y=81360
X2416 1 2 618 68 17 ICV_40 $T=97980 111520 1 0 $X=97790 $Y=108560
X2417 1 2 670 632 11 ICV_40 $T=119140 62560 0 0 $X=118950 $Y=62320
X2418 1 2 718 725 11 ICV_40 $T=154100 68000 1 0 $X=153910 $Y=65040
X2419 1 2 744 740 11 ICV_40 $T=161000 106080 0 0 $X=160810 $Y=105840
X2420 1 2 809 810 33 ICV_40 $T=188600 57120 0 0 $X=188410 $Y=56880
X2421 1 2 779 734 20 ICV_40 $T=188600 89760 1 0 $X=188410 $Y=86800
X2422 1 2 813 817 20 ICV_40 $T=195960 89760 0 0 $X=195770 $Y=89520
X2423 1 2 854 857 20 ICV_40 $T=218960 89760 1 0 $X=218770 $Y=86800
X2424 1 2 1025 1005 170 ICV_40 $T=307280 100640 1 0 $X=307090 $Y=97680
X2425 1 2 1043 216 177 ICV_40 $T=322000 57120 1 0 $X=321810 $Y=54160
X2426 1 2 1050 1039 180 ICV_40 $T=322460 68000 1 0 $X=322270 $Y=65040
X2427 1 2 1140 1101 177 ICV_40 $T=364320 68000 0 0 $X=364130 $Y=67760
X2428 1 2 1173 233 169 ICV_40 $T=380420 51680 0 0 $X=380230 $Y=51440
X2429 1 2 1227 1199 195 ICV_40 $T=406180 89760 1 0 $X=405990 $Y=86800
X2430 1 2 1238 1212 178 ICV_40 $T=420440 95200 0 0 $X=420250 $Y=94960
X2431 1 2 1265 1270 178 ICV_40 $T=428260 100640 0 0 $X=428070 $Y=100400
X2432 1 2 1298 253 187 ICV_40 $T=442060 111520 1 0 $X=441870 $Y=108560
X2433 1 2 1380 298 294 ICV_40 $T=490820 111520 1 0 $X=490630 $Y=108560
X2434 1 2 1455 1428 288 ICV_40 $T=518880 62560 1 0 $X=518690 $Y=59600
X2435 1 2 1510 1513 275 ICV_40 $T=546480 95200 1 0 $X=546290 $Y=92240
X2436 1 2 1559 1551 267 ICV_40 $T=573620 106080 1 0 $X=573430 $Y=103120
X2437 1 2 1566 1565 267 ICV_40 $T=581440 78880 1 0 $X=581250 $Y=75920
X2438 1 2 1579 1551 280 ICV_40 $T=582360 106080 1 0 $X=582170 $Y=103120
X2439 1 2 1607 1612 267 ICV_40 $T=593860 73440 1 0 $X=593670 $Y=70480
X2440 1 2 1645 1657 277 ICV_40 $T=617780 84320 1 0 $X=617590 $Y=81360
X2441 1 2 1799 1800 304 ICV_40 $T=691840 95200 0 0 $X=691650 $Y=94960
X2442 1 2 560 24 572 ICV_41 $T=63940 78880 0 0 $X=63750 $Y=78640
X2443 1 2 51 25 602 ICV_41 $T=79120 106080 0 0 $X=78930 $Y=105840
X2444 1 2 594 8 62 ICV_41 $T=81880 51680 1 0 $X=81690 $Y=48720
X2445 1 2 607 25 640 ICV_41 $T=98900 78880 0 0 $X=98710 $Y=78640
X2446 1 2 629 5 655 ICV_41 $T=107180 62560 0 0 $X=106990 $Y=62320
X2447 1 2 679 24 88 ICV_41 $T=128340 106080 0 0 $X=128150 $Y=105840
X2448 1 2 732 8 746 ICV_41 $T=149500 84320 1 0 $X=149310 $Y=81360
X2449 1 2 738 26 758 ICV_41 $T=156860 62560 0 0 $X=156670 $Y=62320
X2450 1 2 837 4 867 ICV_41 $T=219420 57120 0 0 $X=219230 $Y=56880
X2451 1 2 871 166 888 ICV_41 $T=237360 78880 0 0 $X=237170 $Y=78640
X2452 1 2 871 183 916 ICV_41 $T=247480 78880 0 0 $X=247290 $Y=78640
X2453 1 2 883 166 914 ICV_41 $T=247940 57120 0 0 $X=247750 $Y=56880
X2454 1 2 885 166 908 ICV_41 $T=247940 62560 0 0 $X=247750 $Y=62320
X2455 1 2 871 184 918 ICV_41 $T=247940 84320 0 0 $X=247750 $Y=84080
X2456 1 2 885 183 922 ICV_41 $T=248860 73440 1 0 $X=248670 $Y=70480
X2457 1 2 1049 166 1088 ICV_41 $T=331660 68000 0 0 $X=331470 $Y=67760
X2458 1 2 1089 164 1126 ICV_41 $T=350520 78880 0 0 $X=350330 $Y=78640
X2459 1 2 1180 167 1203 ICV_41 $T=387780 84320 0 0 $X=387590 $Y=84080
X2460 1 2 1205 160 1241 ICV_41 $T=408020 106080 0 0 $X=407830 $Y=105840
X2461 1 2 1242 168 1260 ICV_41 $T=415840 78880 0 0 $X=415650 $Y=78640
X2462 1 2 1250 175 1293 ICV_41 $T=433780 95200 0 0 $X=433590 $Y=94960
X2463 1 2 1256 166 1297 ICV_41 $T=435620 57120 0 0 $X=435430 $Y=56880
X2464 1 2 1305 266 1344 ICV_41 $T=458620 95200 1 0 $X=458430 $Y=92240
X2465 1 2 1382 301 1403 ICV_41 $T=484380 84320 0 0 $X=484190 $Y=84080
X2466 1 2 1381 287 1411 ICV_41 $T=500020 68000 0 0 $X=499830 $Y=67760
X2467 1 2 1471 266 1477 ICV_41 $T=528540 68000 0 0 $X=528350 $Y=67760
X2468 1 2 329 283 1519 ICV_41 $T=542340 111520 1 0 $X=542150 $Y=108560
X2469 1 2 1544 259 1559 ICV_41 $T=563500 100640 1 0 $X=563310 $Y=97680
X2470 1 2 1592 264 1613 ICV_41 $T=588340 84320 1 0 $X=588150 $Y=81360
X2471 1 2 350 301 1627 ICV_41 $T=598920 51680 1 0 $X=598730 $Y=48720
X2472 1 2 1690 258 1724 ICV_41 $T=644920 89760 1 0 $X=644730 $Y=86800
X2473 1 2 1754 297 387 ICV_41 $T=668840 111520 0 0 $X=668650 $Y=111280
X2474 1 2 459 14 18 461 14 11 ICV_44 $T=17020 106080 0 0 $X=16830 $Y=105840
X2475 1 2 569 47 33 565 47 34 ICV_44 $T=69460 68000 0 0 $X=69270 $Y=67760
X2476 1 2 606 586 18 609 586 20 ICV_44 $T=87400 73440 1 0 $X=87210 $Y=70480
X2477 1 2 698 700 18 693 700 30 ICV_44 $T=132480 95200 1 0 $X=132290 $Y=92240
X2478 1 2 717 725 34 724 725 20 ICV_44 $T=146280 57120 0 0 $X=146090 $Y=56880
X2479 1 2 723 700 34 733 734 32 ICV_44 $T=146280 89760 0 0 $X=146090 $Y=89520
X2480 1 2 735 734 30 746 748 11 ICV_44 $T=151340 89760 1 0 $X=151150 $Y=86800
X2481 1 2 788 784 20 789 784 32 ICV_44 $T=178480 95200 1 0 $X=178290 $Y=92240
X2482 1 2 898 892 180 899 892 169 ICV_44 $T=244720 57120 1 0 $X=244530 $Y=54160
X2483 1 2 929 923 169 933 923 195 ICV_44 $T=258060 95200 1 0 $X=257870 $Y=92240
X2484 1 2 992 977 194 1001 1005 191 ICV_44 $T=291640 95200 1 0 $X=291450 $Y=92240
X2485 1 2 1006 977 169 1004 977 195 ICV_44 $T=297620 89760 0 0 $X=297430 $Y=89520
X2486 1 2 1132 1133 182 1138 1133 188 ICV_44 $T=362480 95200 1 0 $X=362290 $Y=92240
X2487 1 2 1150 226 177 1152 226 195 ICV_44 $T=370760 51680 0 0 $X=370570 $Y=51440
X2488 1 2 1154 1157 194 1163 1149 171 ICV_44 $T=370760 73440 1 0 $X=370570 $Y=70480
X2489 1 2 1176 1149 195 1183 1149 180 ICV_44 $T=382260 68000 0 0 $X=382070 $Y=67760
X2490 1 2 245 246 171 1233 246 180 ICV_44 $T=407100 51680 0 0 $X=406910 $Y=51440
X2491 1 2 247 244 187 248 244 182 ICV_44 $T=410320 111520 0 0 $X=410130 $Y=111280
X2492 1 2 1264 1261 194 1276 1261 169 ICV_44 $T=427340 78880 1 0 $X=427150 $Y=75920
X2493 1 2 1326 1331 267 1321 1333 268 ICV_44 $T=455860 89760 1 0 $X=455670 $Y=86800
X2494 1 2 1696 1697 277 1699 1701 276 ICV_44 $T=635260 89760 0 0 $X=635070 $Y=89520
X2495 1 2 1827 1829 307 1840 1829 309 ICV_44 $T=701500 78880 1 0 $X=701310 $Y=75920
X2496 1 2 1893 1882 304 1901 1882 296 ICV_44 $T=733240 95200 1 0 $X=733050 $Y=92240
X2497 1 2 10 5 474 ICV_47 $T=10580 57120 1 0 $X=10390 $Y=54160
X2498 1 2 45 5 59 ICV_47 $T=69460 51680 0 0 $X=69270 $Y=51440
X2499 1 2 679 6 701 ICV_47 $T=125580 100640 0 0 $X=125390 $Y=100400
X2500 1 2 790 26 806 ICV_47 $T=178480 57120 0 0 $X=178290 $Y=56880
X2501 1 2 837 26 863 ICV_47 $T=216660 51680 1 0 $X=216470 $Y=48720
X2502 1 2 871 167 901 ICV_47 $T=235980 89760 0 0 $X=235790 $Y=89520
X2503 1 2 196 173 948 ICV_47 $T=259900 111520 1 0 $X=259710 $Y=108560
X2504 1 2 909 183 957 ICV_47 $T=265880 84320 0 0 $X=265690 $Y=84080
X2505 1 2 926 160 973 ICV_47 $T=273700 100640 0 0 $X=273510 $Y=100400
X2506 1 2 197 166 982 ICV_47 $T=276920 51680 0 0 $X=276730 $Y=51440
X2507 1 2 959 186 1004 ICV_47 $T=288880 89760 0 0 $X=288690 $Y=89520
X2508 1 2 207 157 209 ICV_47 $T=288880 111520 0 0 $X=288690 $Y=111280
X2509 1 2 1009 185 1036 ICV_47 $T=305440 57120 0 0 $X=305250 $Y=56880
X2510 1 2 1089 186 1098 ICV_47 $T=338100 84320 1 0 $X=337910 $Y=81360
X2511 1 2 1148 186 1176 ICV_47 $T=375820 68000 1 0 $X=375630 $Y=65040
X2512 1 2 1145 184 1185 ICV_47 $T=379500 78880 0 0 $X=379310 $Y=78640
X2513 1 2 1188 185 1232 ICV_47 $T=403420 78880 1 0 $X=403230 $Y=75920
X2514 1 2 282 283 1358 ICV_47 $T=465520 51680 0 0 $X=465330 $Y=51440
X2515 1 2 1409 302 1427 ICV_47 $T=497260 57120 1 0 $X=497070 $Y=54160
X2516 1 2 1420 265 1439 ICV_47 $T=501860 84320 0 0 $X=501670 $Y=84080
X2517 1 2 329 305 1511 ICV_47 $T=539120 111520 0 0 $X=538930 $Y=111280
X2518 1 2 1500 272 1518 ICV_47 $T=540960 100640 1 0 $X=540770 $Y=97680
X2519 1 2 336 305 1574 ICV_47 $T=569940 57120 1 0 $X=569750 $Y=54160
X2520 1 2 1554 265 1590 ICV_47 $T=576840 78880 0 0 $X=576650 $Y=78640
X2521 1 2 1569 259 1602 ICV_47 $T=585120 57120 0 0 $X=584930 $Y=56880
X2522 1 2 1616 264 1634 ICV_47 $T=598000 68000 1 0 $X=597810 $Y=65040
X2523 1 2 1731 292 1772 ICV_47 $T=667000 84320 0 0 $X=666810 $Y=84080
X2524 1 2 1736 299 389 ICV_47 $T=669760 51680 0 0 $X=669570 $Y=51440
X2525 1 2 1868 301 1893 ICV_47 $T=730480 89760 1 0 $X=730290 $Y=86800
X2526 1 2 517 40 32 ICV_48 $T=43700 57120 1 0 $X=43510 $Y=54160
X2527 1 2 549 534 17 ICV_48 $T=57500 106080 0 0 $X=57310 $Y=105840
X2528 1 2 630 64 17 ICV_48 $T=99820 62560 1 0 $X=99630 $Y=59600
X2529 1 2 683 86 32 ICV_48 $T=127880 106080 1 0 $X=127690 $Y=103120
X2530 1 2 712 700 11 ICV_48 $T=141680 84320 0 0 $X=141490 $Y=84080
X2531 1 2 846 826 32 ICV_48 $T=212060 68000 1 0 $X=211870 $Y=65040
X2532 1 2 888 886 171 ICV_48 $T=240120 84320 1 0 $X=239930 $Y=81360
X2533 1 2 915 890 192 ICV_48 $T=253920 68000 0 0 $X=253730 $Y=67760
X2534 1 2 974 977 193 ICV_48 $T=281980 89760 0 0 $X=281790 $Y=89520
X2535 1 2 1120 1101 193 ICV_48 $T=352360 68000 1 0 $X=352170 $Y=65040
X2536 1 2 1314 1315 268 ICV_48 $T=450340 95200 0 0 $X=450150 $Y=94960
X2537 1 2 1344 1331 277 ICV_48 $T=464600 100640 1 0 $X=464410 $Y=97680
X2538 1 2 1371 1357 296 ICV_48 $T=478400 57120 0 0 $X=478210 $Y=56880
X2539 1 2 1404 1386 307 ICV_48 $T=492660 73440 1 0 $X=492470 $Y=70480
X2540 1 2 1534 334 303 ICV_48 $T=562580 51680 0 0 $X=562390 $Y=51440
X2541 1 2 353 354 307 ICV_48 $T=590640 51680 0 0 $X=590450 $Y=51440
X2542 1 2 1598 1600 277 ICV_48 $T=590640 100640 0 0 $X=590450 $Y=100400
X2543 1 2 1747 1748 296 ICV_48 $T=661020 84320 1 0 $X=660830 $Y=81360
X2544 1 2 1773 1774 304 ICV_48 $T=674820 100640 0 0 $X=674630 $Y=100400
X2545 1 2 1831 1829 294 ICV_48 $T=702880 84320 0 0 $X=702690 $Y=84080
X2546 1 2 671 4 696 696 692 20 ICV_49 $T=122360 73440 0 0 $X=122170 $Y=73200
X2547 1 2 790 27 834 834 810 34 ICV_49 $T=192740 62560 1 0 $X=192550 $Y=59600
X2548 1 2 196 181 949 949 198 189 ICV_49 $T=258520 106080 0 0 $X=258330 $Y=105840
X2549 1 2 197 168 954 936 892 194 ICV_49 $T=262660 51680 0 0 $X=262470 $Y=51440
X2550 1 2 989 181 1000 1000 1005 189 ICV_49 $T=286580 100640 0 0 $X=286390 $Y=100400
X2551 1 2 207 165 1032 1031 211 182 ICV_49 $T=300840 111520 1 0 $X=300650 $Y=108560
X2552 1 2 1096 184 1117 1117 1110 192 ICV_49 $T=342700 84320 0 0 $X=342510 $Y=84080
X2553 1 2 1089 184 1127 1127 1100 192 ICV_49 $T=350060 73440 0 0 $X=349870 $Y=73200
X2554 1 2 1162 160 1200 1200 1168 174 ICV_49 $T=384100 100640 0 0 $X=383910 $Y=100400
X2555 1 2 1242 184 1258 1258 1261 192 ICV_49 $T=413080 73440 1 0 $X=412890 $Y=70480
X2556 1 2 1375 272 1387 1387 1389 280 ICV_49 $T=476560 111520 1 0 $X=476370 $Y=108560
X2557 1 2 1506 264 1537 1537 1525 276 ICV_49 $T=550620 89760 0 0 $X=550430 $Y=89520
X2558 1 2 1527 257 1543 1545 1546 269 ICV_49 $T=552460 62560 0 0 $X=552270 $Y=62320
X2559 1 2 1782 299 1796 1796 1798 307 ICV_49 $T=678040 57120 1 0 $X=677850 $Y=54160
X2560 1 2 1807 299 1830 1833 1824 294 ICV_49 $T=693680 57120 1 0 $X=693490 $Y=54160
X2561 1 2 1819 301 1859 1859 1829 304 ICV_49 $T=706560 84320 1 0 $X=706370 $Y=81360
X2562 1 2 509 27 545 545 525 34 ICV_50 $T=45540 57120 0 0 $X=45350 $Y=56880
X2563 1 2 610 5 618 616 615 30 ICV_50 $T=86020 95200 1 0 $X=85830 $Y=92240
X2564 1 2 610 4 73 641 643 11 ICV_50 $T=94300 95200 0 0 $X=94110 $Y=94960
X2565 1 2 72 26 660 655 632 17 ICV_50 $T=104420 62560 1 0 $X=104230 $Y=59600
X2566 1 2 72 5 676 82 80 34 ICV_50 $T=111780 51680 1 0 $X=111590 $Y=48720
X2567 1 2 675 6 684 664 643 30 ICV_50 $T=118220 78880 0 0 $X=118030 $Y=78640
X2568 1 2 775 6 797 797 792 18 ICV_50 $T=172040 68000 1 0 $X=171850 $Y=65040
X2569 1 2 871 185 920 922 890 193 ICV_50 $T=244720 78880 1 0 $X=244530 $Y=75920
X2570 1 2 871 186 921 918 886 192 ICV_50 $T=244720 84320 1 0 $X=244530 $Y=81360
X2571 1 2 926 181 951 951 943 189 ICV_50 $T=258520 100640 0 0 $X=258330 $Y=100400
X2572 1 2 1471 259 1483 1483 1479 267 ICV_50 $T=523480 57120 0 0 $X=523290 $Y=56880
X2573 1 2 1500 262 1529 1529 1513 273 ICV_50 $T=546940 95200 0 0 $X=546750 $Y=94960
X2574 1 2 1616 258 1628 1583 1582 280 ICV_50 $T=595240 68000 0 0 $X=595050 $Y=67760
X2575 1 2 1593 265 1632 1632 1601 275 ICV_50 $T=595240 89760 0 0 $X=595050 $Y=89520
X2576 1 2 1637 257 1651 1651 1657 268 ICV_50 $T=606280 73440 0 0 $X=606090 $Y=73200
X2577 1 2 1736 297 1775 1775 384 303 ICV_50 $T=665620 62560 1 0 $X=665430 $Y=59600
X2578 1 2 1808 299 1825 1826 1816 294 ICV_50 $T=691380 68000 0 0 $X=691190 $Y=67760
X2579 1 2 1817 301 1836 1835 1838 303 ICV_50 $T=693680 111520 1 0 $X=693490 $Y=108560
X2580 1 2 1808 292 1848 1848 1816 300 ICV_50 $T=702880 68000 1 0 $X=702690 $Y=65040
X2581 1 2 523 525 32 540 24 548 ICV_51 $T=50140 62560 0 0 $X=49950 $Y=62320
X2582 1 2 536 534 18 39 26 559 ICV_51 $T=51060 106080 1 0 $X=50870 $Y=103120
X2583 1 2 561 563 30 566 6 579 ICV_51 $T=62560 100640 1 0 $X=62370 $Y=97680
X2584 1 2 584 586 32 591 26 584 ICV_51 $T=76820 62560 0 0 $X=76630 $Y=62320
X2585 1 2 611 64 33 594 26 634 ICV_51 $T=90620 57120 0 0 $X=90430 $Y=56880
X2586 1 2 638 632 30 72 25 659 ICV_51 $T=103960 57120 0 0 $X=103770 $Y=56880
X2587 1 2 642 644 30 649 4 663 ICV_51 $T=105340 100640 1 0 $X=105150 $Y=97680
X2588 1 2 645 632 33 629 6 665 ICV_51 $T=106260 68000 0 0 $X=106070 $Y=67760
X2589 1 2 672 644 32 678 4 694 ICV_51 $T=120520 100640 1 0 $X=120330 $Y=97680
X2590 1 2 702 86 20 679 8 703 ICV_51 $T=133860 111520 1 0 $X=133670 $Y=108560
X2591 1 2 755 748 18 741 27 778 ICV_51 $T=162380 89760 1 0 $X=162190 $Y=86800
X2592 1 2 830 810 30 811 26 846 ICV_51 $T=201020 73440 1 0 $X=200830 $Y=70480
X2593 1 2 895 891 174 881 173 913 ICV_51 $T=241960 106080 0 0 $X=241770 $Y=105840
X2594 1 2 946 943 170 926 165 975 ICV_51 $T=271400 95200 0 0 $X=271210 $Y=94960
X2595 1 2 986 988 194 959 164 1006 ICV_51 $T=286580 78880 0 0 $X=286390 $Y=78640
X2596 1 2 978 943 178 989 165 1008 ICV_51 $T=286580 95200 0 0 $X=286390 $Y=94960
X2597 1 2 205 206 194 208 184 210 ICV_51 $T=287500 51680 1 0 $X=287310 $Y=48720
X2598 1 2 1126 1100 169 1096 166 1146 ICV_51 $T=356960 84320 1 0 $X=356770 $Y=81360
X2599 1 2 1143 1101 195 1159 168 1175 ICV_51 $T=370760 57120 0 0 $X=370570 $Y=56880
X2600 1 2 1155 1133 187 1162 156 1174 ICV_51 $T=371220 95200 0 0 $X=371030 $Y=94960
X2601 1 2 1158 1133 174 1162 181 1178 ICV_51 $T=372600 100640 0 0 $X=372410 $Y=100400
X2602 1 2 1244 1246 192 1239 168 1268 ICV_51 $T=416300 89760 1 0 $X=416110 $Y=86800
X2603 1 2 255 256 178 1248 156 1291 ICV_51 $T=429180 111520 1 0 $X=428990 $Y=108560
X2604 1 2 1322 1331 273 1305 257 1350 ICV_51 $T=455400 89760 0 0 $X=455210 $Y=89520
X2605 1 2 1329 1333 276 1304 262 1355 ICV_51 $T=457240 84320 1 0 $X=457050 $Y=81360
X2606 1 2 1355 1333 273 1304 272 1372 ICV_51 $T=467360 78880 0 0 $X=467170 $Y=78640
X2607 1 2 286 1357 288 282 292 1379 ICV_51 $T=471040 51680 1 0 $X=470850 $Y=48720
X2608 1 2 1383 298 303 1375 264 1407 ICV_51 $T=483920 106080 0 0 $X=483730 $Y=105840
X2609 1 2 1385 1386 304 1381 305 1408 ICV_51 $T=485300 84320 1 0 $X=485110 $Y=81360
X2610 1 2 1412 1386 309 1418 264 1435 ICV_51 $T=498640 73440 1 0 $X=498450 $Y=70480
X2611 1 2 1432 298 296 1436 297 1453 ICV_51 $T=506920 106080 1 0 $X=506730 $Y=103120
X2612 1 2 1449 1443 269 1418 266 1472 ICV_51 $T=516120 73440 0 0 $X=515930 $Y=73200
X2613 1 2 1460 1461 268 1436 305 1476 ICV_51 $T=519340 100640 0 0 $X=519150 $Y=100400
X2614 1 2 1501 1479 268 1471 265 1520 ICV_51 $T=539120 62560 1 0 $X=538930 $Y=59600
X2615 1 2 1499 1498 275 1506 266 1524 ICV_51 $T=539120 89760 0 0 $X=538930 $Y=89520
X2616 1 2 339 340 309 336 287 1576 ICV_51 $T=568100 51680 1 0 $X=567910 $Y=48720
X2617 1 2 349 345 276 1591 272 1604 ICV_51 $T=582360 111520 0 0 $X=582170 $Y=111280
X2618 1 2 1586 1565 280 1593 262 1610 ICV_51 $T=583280 89760 0 0 $X=583090 $Y=89520
X2619 1 2 1755 384 296 1736 283 1778 ICV_51 $T=666540 57120 1 0 $X=666350 $Y=54160
X2620 1 2 1772 1746 300 1781 301 1773 ICV_51 $T=674360 89760 1 0 $X=674170 $Y=86800
X2621 1 2 396 397 304 1817 297 1835 ICV_51 $T=693220 106080 0 0 $X=693030 $Y=105840
X2622 1 2 1811 1774 309 1819 299 1827 ICV_51 $T=695060 84320 1 0 $X=694870 $Y=81360
X2623 1 2 1815 1774 307 1819 283 1831 ICV_51 $T=695980 89760 1 0 $X=695790 $Y=86800
X2624 1 2 572 573 30 ICV_52 $T=70840 73440 0 0 $X=70650 $Y=73200
X2625 1 2 598 563 20 ICV_52 $T=84180 89760 0 0 $X=83990 $Y=89520
X2626 1 2 604 586 17 ICV_52 $T=94300 68000 1 0 $X=94110 $Y=65040
X2627 1 2 716 90 34 ICV_52 $T=146280 51680 0 0 $X=146090 $Y=51440
X2628 1 2 801 784 18 ICV_52 $T=183540 106080 0 0 $X=183350 $Y=105840
X2629 1 2 819 114 32 ICV_52 $T=196420 51680 0 0 $X=196230 $Y=51440
X2630 1 2 808 784 30 ICV_52 $T=196420 95200 0 0 $X=196230 $Y=94960
X2631 1 2 912 891 189 ICV_52 $T=252540 100640 0 0 $X=252350 $Y=100400
X2632 1 2 1064 1053 182 ICV_52 $T=328900 95200 1 0 $X=328710 $Y=92240
X2633 1 2 1213 1210 171 ICV_52 $T=407100 68000 1 0 $X=406910 $Y=65040
X2634 1 2 1272 1270 188 ICV_52 $T=427800 89760 0 0 $X=427610 $Y=89520
X2635 1 2 1402 1357 307 ICV_52 $T=491280 57120 1 0 $X=491090 $Y=54160
X2636 1 2 1413 1386 300 ICV_52 $T=499100 78880 1 0 $X=498910 $Y=75920
X2637 1 2 1423 1399 288 ICV_52 $T=505080 89760 0 0 $X=504890 $Y=89520
X2638 1 2 1558 340 294 ICV_52 $T=573620 51680 0 0 $X=573430 $Y=51440
X2639 1 2 1633 1601 268 ICV_52 $T=605360 95200 0 0 $X=605170 $Y=94960
X2640 1 2 1622 1625 268 ICV_52 $T=617320 57120 0 0 $X=617130 $Y=56880
X2641 1 2 1706 1697 280 ICV_52 $T=659640 100640 1 0 $X=659450 $Y=97680
X2642 1 2 1825 1816 307 ICV_52 $T=701500 62560 0 0 $X=701310 $Y=62320
X2643 1 2 1860 1829 288 ICV_52 $T=715760 95200 1 0 $X=715570 $Y=92240
X2644 1 2 1788 1774 288 ICV_52 $T=721280 84320 0 0 $X=721090 $Y=84080
X2645 1 2 116 2 120 1 sky130_fd_sc_hd__clkbuf_16 $T=187220 95200 0 0 $X=187030 $Y=94960
X2646 1 2 118 2 119 1 sky130_fd_sc_hd__clkbuf_16 $T=188600 95200 1 0 $X=188410 $Y=92240
X2647 1 2 147 2 117 1 sky130_fd_sc_hd__clkbuf_16 $T=224940 89760 1 0 $X=224750 $Y=86800
X2648 1 2 505 473 33 ICV_56 $T=34960 89760 0 0 $X=34770 $Y=89520
X2649 1 2 582 47 20 ICV_56 $T=82800 73440 0 0 $X=82610 $Y=73200
X2650 1 2 688 692 18 ICV_56 $T=131560 57120 0 0 $X=131370 $Y=56880
X2651 1 2 764 760 17 ICV_56 $T=166980 62560 0 0 $X=166790 $Y=62320
X2652 1 2 766 740 17 ICV_56 $T=166980 106080 0 0 $X=166790 $Y=105840
X2653 1 2 867 139 20 ICV_56 $T=230460 57120 0 0 $X=230270 $Y=56880
X2654 1 2 975 943 188 ICV_56 $T=281980 100640 1 0 $X=281790 $Y=97680
X2655 1 2 990 967 194 ICV_56 $T=298080 62560 0 0 $X=297890 $Y=62320
X2656 1 2 1109 1100 171 ICV_56 $T=349140 84320 1 0 $X=348950 $Y=81360
X2657 1 2 1277 252 192 ICV_56 $T=433780 57120 1 0 $X=433590 $Y=54160
X2658 1 2 1287 1262 169 ICV_56 $T=439760 62560 0 0 $X=439570 $Y=62320
X2659 1 2 1490 1461 276 ICV_56 $T=535440 111520 1 0 $X=535250 $Y=108560
X2660 1 2 1489 1498 280 ICV_56 $T=536360 78880 1 0 $X=536170 $Y=75920
X2661 1 2 1567 1546 275 ICV_56 $T=574080 68000 1 0 $X=573890 $Y=65040
X2662 1 2 1668 1674 276 ICV_56 $T=626060 68000 0 0 $X=625870 $Y=67760
X2663 1 2 1679 1674 268 ICV_56 $T=630200 68000 1 0 $X=630010 $Y=65040
X2664 1 2 1716 1701 280 ICV_56 $T=644000 89760 0 0 $X=643810 $Y=89520
X2665 1 2 1771 1748 300 ICV_56 $T=677580 84320 1 0 $X=677390 $Y=81360
X2666 1 2 454 25 503 496 451 34 ICV_58 $T=24380 100640 1 0 $X=24190 $Y=97680
X2667 1 2 39 6 536 535 534 33 ICV_58 $T=40480 106080 0 0 $X=40290 $Y=105840
X2668 1 2 51 24 603 602 54 33 ICV_58 $T=76360 111520 1 0 $X=76170 $Y=108560
X2669 1 2 678 6 698 694 700 20 ICV_58 $T=122360 95200 0 0 $X=122170 $Y=94960
X2670 1 2 730 4 747 747 740 20 ICV_58 $T=146280 106080 0 0 $X=146090 $Y=105840
X2671 1 2 738 6 761 761 760 18 ICV_58 $T=156400 68000 0 0 $X=156210 $Y=67760
X2672 1 2 926 157 978 971 943 187 ICV_58 $T=272780 106080 1 0 $X=272590 $Y=103120
X2673 1 2 984 186 997 995 988 193 ICV_58 $T=284280 73440 1 0 $X=284090 $Y=70480
X2674 1 2 1078 160 1115 1115 1074 174 ICV_58 $T=340860 106080 1 0 $X=340670 $Y=103120
X2675 1 2 1078 165 1116 1116 1074 188 ICV_58 $T=341320 100640 1 0 $X=341130 $Y=97680
X2676 1 2 1102 167 1118 1093 1071 195 ICV_58 $T=342700 57120 0 0 $X=342510 $Y=56880
X2677 1 2 1102 183 1120 1091 1071 194 ICV_58 $T=342700 62560 0 0 $X=342510 $Y=62320
X2678 1 2 1204 186 1229 1221 1228 194 ICV_58 $T=397900 57120 1 0 $X=397710 $Y=54160
X2679 1 2 1256 183 1283 1283 1262 193 ICV_58 $T=425500 68000 1 0 $X=425310 $Y=65040
X2680 1 2 1382 297 1414 1415 1399 300 ICV_58 $T=490360 89760 0 0 $X=490170 $Y=89520
X2681 1 2 1420 272 1440 1440 1431 280 ICV_58 $T=501400 84320 1 0 $X=501210 $Y=81360
X2682 1 2 1506 262 1548 1549 1525 275 ICV_58 $T=553380 84320 1 0 $X=553190 $Y=81360
X2683 1 2 1506 272 1550 1548 1525 273 ICV_58 $T=553380 89760 1 0 $X=553190 $Y=86800
X2684 1 2 1695 262 1730 1730 1697 273 ICV_58 $T=644920 100640 1 0 $X=644730 $Y=97680
X2685 1 2 1782 283 1793 1792 1798 300 ICV_58 $T=677120 68000 1 0 $X=676930 $Y=65040
X2686 1 2 1776 287 1834 1822 1800 288 ICV_58 $T=693680 95200 1 0 $X=693490 $Y=92240
X2687 1 2 738 5 764 765 760 33 ICV_59 $T=160080 68000 1 0 $X=159890 $Y=65040
X2688 1 2 952 167 993 993 967 180 ICV_59 $T=286120 57120 0 0 $X=285930 $Y=56880
X2689 1 2 952 168 994 994 967 177 ICV_59 $T=286120 62560 0 0 $X=285930 $Y=62320
X2690 1 2 1033 166 1081 1081 1039 171 ICV_59 $T=328440 73440 1 0 $X=328250 $Y=70480
X2691 1 2 1148 166 1163 1160 1149 177 ICV_59 $T=370300 68000 0 0 $X=370110 $Y=67760
X2692 1 2 1148 185 1191 1191 1149 194 ICV_59 $T=384560 73440 1 0 $X=384370 $Y=70480
X2693 1 2 1180 183 1192 1192 1199 193 ICV_59 $T=384560 89760 1 0 $X=384370 $Y=86800
X2694 1 2 1180 168 1224 1224 1199 177 ICV_59 $T=398360 89760 0 0 $X=398170 $Y=89520
X2695 1 2 239 156 1226 1226 244 170 ICV_59 $T=398360 111520 0 0 $X=398170 $Y=111280
X2696 1 2 1204 183 1254 1254 1228 193 ICV_59 $T=412620 57120 1 0 $X=412430 $Y=54160
X2697 1 2 1491 257 1535 1528 1512 276 ICV_59 $T=552920 73440 1 0 $X=552730 $Y=70480
X2698 1 2 1591 257 1649 1650 1600 275 ICV_59 $T=609040 106080 1 0 $X=608850 $Y=103120
X2699 1 2 1591 265 1650 1644 1600 267 ICV_59 $T=609040 111520 1 0 $X=608850 $Y=108560
X2700 1 2 1646 257 1679 1673 1674 267 ICV_59 $T=622840 57120 0 0 $X=622650 $Y=56880
X2701 1 2 1646 272 1680 1680 1674 280 ICV_59 $T=622840 62560 0 0 $X=622650 $Y=62320
X2702 1 2 1694 266 1712 1712 1709 277 ICV_59 $T=637100 68000 1 0 $X=636910 $Y=65040
X2703 1 2 1692 258 1740 1740 1708 269 ICV_59 $T=650900 73440 0 0 $X=650710 $Y=73200
X2704 1 2 1731 302 1766 1766 1746 309 ICV_59 $T=665160 95200 1 0 $X=664970 $Y=92240
X2705 1 2 1807 305 1849 1849 1824 288 ICV_59 $T=707020 57120 0 0 $X=706830 $Y=56880
X2706 1 2 21 476 ICV_61 $T=22540 62560 0 0 $X=22350 $Y=62320
X2707 1 2 36 508 ICV_61 $T=57960 78880 0 0 $X=57770 $Y=78640
X2708 1 2 71 643 ICV_61 $T=122820 89760 0 0 $X=122630 $Y=89520
X2709 1 2 87 658 ICV_61 $T=142600 78880 0 0 $X=142410 $Y=78640
X2710 1 2 84 86 ICV_61 $T=145360 111520 1 0 $X=145170 $Y=108560
X2711 1 2 93 725 ICV_61 $T=153640 62560 0 0 $X=153450 $Y=62320
X2712 1 2 134 856 ICV_61 $T=226320 68000 0 0 $X=226130 $Y=67760
X2713 1 2 21 892 ICV_61 $T=240580 68000 1 0 $X=240390 $Y=65040
X2714 1 2 36 940 ICV_61 $T=266800 78880 0 0 $X=266610 $Y=78640
X2715 1 2 138 1133 ICV_61 $T=366620 100640 0 0 $X=366430 $Y=100400
X2716 1 2 109 233 ICV_61 $T=380880 62560 1 0 $X=380690 $Y=59600
X2717 1 2 137 1168 ICV_61 $T=394680 95200 1 0 $X=394490 $Y=92240
X2718 1 2 321 1443 ICV_61 $T=525320 68000 1 0 $X=525130 $Y=65040
X2719 1 2 346 1565 ICV_61 $T=587880 89760 1 0 $X=587690 $Y=86800
X2720 1 2 356 1612 ICV_61 $T=606740 78880 0 0 $X=606550 $Y=78640
X2721 1 2 274 379 ICV_61 $T=658720 51680 0 0 $X=658530 $Y=51440
X2722 1 2 370 1708 ICV_61 $T=661480 73440 1 0 $X=661290 $Y=70480
X2723 1 2 355 398 ICV_61 $T=693680 51680 1 0 $X=693490 $Y=48720
X2724 1 2 321 1824 ICV_61 $T=702880 62560 1 0 $X=702690 $Y=59600
X2725 1 2 490 476 34 ICV_62 $T=34040 62560 0 0 $X=33850 $Y=62320
X2726 1 2 526 525 33 ICV_62 $T=48300 73440 1 0 $X=48110 $Y=70480
X2727 1 2 557 534 30 ICV_62 $T=62100 95200 0 0 $X=61910 $Y=94960
X2728 1 2 559 534 32 ICV_62 $T=62100 100640 0 0 $X=61910 $Y=100400
X2729 1 2 673 644 17 ICV_62 $T=120980 111520 1 0 $X=120790 $Y=108560
X2730 1 2 674 80 18 ICV_62 $T=121440 51680 0 0 $X=121250 $Y=51440
X2731 1 2 785 734 33 ICV_62 $T=177100 89760 0 0 $X=176910 $Y=89520
X2732 1 2 861 857 33 ICV_62 $T=221260 78880 0 0 $X=221070 $Y=78640
X2733 1 2 948 198 191 ICV_62 $T=267720 106080 1 0 $X=267530 $Y=103120
X2734 1 2 956 923 194 ICV_62 $T=272780 89760 1 0 $X=272590 $Y=86800
X2735 1 2 957 923 193 ICV_62 $T=273700 84320 1 0 $X=273510 $Y=81360
X2736 1 2 1070 1071 192 ICV_62 $T=329360 62560 1 0 $X=329170 $Y=59600
X2737 1 2 1088 1071 171 ICV_62 $T=342700 68000 0 0 $X=342510 $Y=67760
X2738 1 2 1103 221 171 ICV_62 $T=349140 57120 1 0 $X=348950 $Y=54160
X2739 1 2 1125 1100 194 ICV_62 $T=364320 73440 0 0 $X=364130 $Y=73200
X2740 1 2 1171 232 188 ICV_62 $T=379500 106080 0 0 $X=379310 $Y=105840
X2741 1 2 1202 1168 188 ICV_62 $T=393760 95200 0 0 $X=393570 $Y=94960
X2742 1 2 1206 1210 169 ICV_62 $T=413080 68000 1 0 $X=412890 $Y=65040
X2743 1 2 1275 1262 195 ICV_62 $T=435160 62560 0 0 $X=434970 $Y=62320
X2744 1 2 1342 1311 276 ICV_62 $T=464140 73440 1 0 $X=463950 $Y=70480
X2745 1 2 1417 1389 267 ICV_62 $T=501860 100640 0 0 $X=501670 $Y=100400
X2746 1 2 1419 1389 275 ICV_62 $T=502320 106080 1 0 $X=502130 $Y=103120
X2747 1 2 1439 1431 275 ICV_62 $T=520260 89760 1 0 $X=520070 $Y=86800
X2748 1 2 1453 1446 303 ICV_62 $T=525320 95200 1 0 $X=525130 $Y=92240
X2749 1 2 1463 1461 269 ICV_62 $T=525320 106080 1 0 $X=525130 $Y=103120
X2750 1 2 325 1461 280 ICV_62 $T=534060 106080 0 0 $X=533870 $Y=105840
X2751 1 2 1511 333 288 ICV_62 $T=546480 106080 0 0 $X=546290 $Y=105840
X2752 1 2 1519 333 294 ICV_62 $T=548780 111520 0 0 $X=548590 $Y=111280
X2753 1 2 1508 1512 277 ICV_62 $T=557520 57120 0 0 $X=557330 $Y=56880
X2754 1 2 1543 1546 268 ICV_62 $T=562120 57120 0 0 $X=561930 $Y=56880
X2755 1 2 1538 1513 277 ICV_62 $T=562120 95200 0 0 $X=561930 $Y=94960
X2756 1 2 1552 1546 280 ICV_62 $T=567180 68000 1 0 $X=566990 $Y=65040
X2757 1 2 1553 1525 267 ICV_62 $T=567180 89760 0 0 $X=566990 $Y=89520
X2758 1 2 1550 1525 280 ICV_62 $T=568100 84320 1 0 $X=567910 $Y=81360
X2759 1 2 362 358 277 ICV_62 $T=604440 111520 1 0 $X=604250 $Y=108560
X2760 1 2 1658 1660 269 ICV_62 $T=618240 100640 0 0 $X=618050 $Y=100400
X2761 1 2 1677 365 288 ICV_62 $T=634800 51680 0 0 $X=634610 $Y=51440
X2762 1 2 1718 379 304 ICV_62 $T=646300 57120 0 0 $X=646110 $Y=56880
X2763 1 2 1702 1709 280 ICV_62 $T=646300 62560 0 0 $X=646110 $Y=62320
X2764 1 2 1714 1708 277 ICV_62 $T=646300 73440 0 0 $X=646110 $Y=73200
X2765 1 2 1721 1709 275 ICV_62 $T=660560 62560 1 0 $X=660370 $Y=59600
X2766 1 2 1749 1746 304 ICV_62 $T=661480 89760 0 0 $X=661290 $Y=89520
X2767 1 2 1741 1697 268 ICV_62 $T=665620 100640 1 0 $X=665430 $Y=97680
X2768 1 2 1789 386 304 ICV_62 $T=688620 106080 1 0 $X=688430 $Y=103120
X2769 1 2 1888 1869 303 ICV_62 $T=733240 68000 1 0 $X=733050 $Y=65040
X2770 1 2 10 4 475 ICV_66 $T=12420 51680 1 0 $X=12230 $Y=48720
X2771 1 2 10 24 29 ICV_66 $T=26220 51680 0 0 $X=26030 $Y=51440
X2772 1 2 454 27 496 ICV_66 $T=26220 95200 0 0 $X=26030 $Y=94960
X2773 1 2 512 27 527 ICV_66 $T=40480 89760 1 0 $X=40290 $Y=86800
X2774 1 2 39 8 529 ICV_66 $T=40480 106080 1 0 $X=40290 $Y=103120
X2775 1 2 594 4 608 ICV_66 $T=82340 57120 0 0 $X=82150 $Y=56880
X2776 1 2 607 8 635 ICV_66 $T=96600 89760 1 0 $X=96410 $Y=86800
X2777 1 2 649 26 666 ICV_66 $T=110400 89760 0 0 $X=110210 $Y=89520
X2778 1 2 708 27 717 ICV_66 $T=138460 57120 0 0 $X=138270 $Y=56880
X2779 1 2 678 5 713 ICV_66 $T=138460 95200 0 0 $X=138270 $Y=94960
X2780 1 2 679 5 719 ICV_66 $T=138460 106080 0 0 $X=138270 $Y=105840
X2781 1 2 738 8 753 ICV_66 $T=152720 62560 1 0 $X=152530 $Y=59600
X2782 1 2 741 4 779 ICV_66 $T=166520 89760 0 0 $X=166330 $Y=89520
X2783 1 2 837 24 851 ICV_66 $T=208840 57120 1 0 $X=208650 $Y=54160
X2784 1 2 161 166 897 ICV_66 $T=236900 51680 1 0 $X=236710 $Y=48720
X2785 1 2 883 167 898 ICV_66 $T=236900 57120 1 0 $X=236710 $Y=54160
X2786 1 2 883 164 899 ICV_66 $T=236900 62560 1 0 $X=236710 $Y=59600
X2787 1 2 162 165 172 ICV_66 $T=236900 111520 1 0 $X=236710 $Y=108560
X2788 1 2 1049 164 1065 ICV_66 $T=321080 62560 1 0 $X=320890 $Y=59600
X2789 1 2 1020 167 1067 ICV_66 $T=321080 89760 1 0 $X=320890 $Y=86800
X2790 1 2 1188 164 1206 ICV_66 $T=391000 68000 0 0 $X=390810 $Y=67760
X2791 1 2 1242 185 1264 ICV_66 $T=419060 73440 0 0 $X=418870 $Y=73200
X2792 1 2 1250 157 1265 ICV_66 $T=419060 100640 0 0 $X=418870 $Y=100400
X2793 1 2 1248 157 250 ICV_66 $T=419060 111520 0 0 $X=418870 $Y=111280
X2794 1 2 1256 164 1287 ICV_66 $T=433320 62560 1 0 $X=433130 $Y=59600
X2795 1 2 1306 257 1314 ICV_66 $T=447120 106080 0 0 $X=446930 $Y=105840
X2796 1 2 320 305 1469 ICV_66 $T=517500 51680 1 0 $X=517310 $Y=48720
X2797 1 2 1471 272 1526 ICV_66 $T=545560 68000 1 0 $X=545370 $Y=65040
X2798 1 2 1544 265 1580 ICV_66 $T=573620 100640 1 0 $X=573430 $Y=97680
X2799 1 2 1592 259 1607 ICV_66 $T=587420 73440 0 0 $X=587230 $Y=73200
X2800 1 2 1646 266 1662 ICV_66 $T=615480 68000 0 0 $X=615290 $Y=67760
X2801 1 2 1781 287 1805 ICV_66 $T=685860 89760 1 0 $X=685670 $Y=86800
X2802 1 2 1819 302 1840 ICV_66 $T=699660 78880 0 0 $X=699470 $Y=78640
X2803 1 2 117 119 120 121 2 111 1 sky130_fd_sc_hd__and4b_2 $T=188140 111520 0 0 $X=187950 $Y=111280
X2804 1 2 117 119 120 814 2 65 1 sky130_fd_sc_hd__and4b_2 $T=189060 106080 0 0 $X=188870 $Y=105840
X2805 1 2 120 119 117 814 2 49 1 sky130_fd_sc_hd__and4b_2 $T=192280 106080 1 0 $X=192090 $Y=103120
X2806 1 2 119 117 120 121 2 50 1 sky130_fd_sc_hd__and4b_2 $T=197800 111520 0 0 $X=197610 $Y=111280
X2807 1 2 119 117 120 829 2 115 1 sky130_fd_sc_hd__and4b_2 $T=198260 95200 1 0 $X=198070 $Y=92240
X2808 1 2 120 119 117 121 2 99 1 sky130_fd_sc_hd__and4b_2 $T=198260 111520 1 0 $X=198070 $Y=108560
X2809 1 2 119 117 120 814 2 61 1 sky130_fd_sc_hd__and4b_2 $T=198720 100640 1 0 $X=198530 $Y=97680
X2810 1 2 123 124 125 126 2 829 1 sky130_fd_sc_hd__and4b_2 $T=203320 106080 0 0 $X=203130 $Y=105840
X2811 1 2 120 119 117 841 2 133 1 sky130_fd_sc_hd__and4b_2 $T=207000 100640 1 0 $X=206810 $Y=97680
X2812 1 2 120 119 117 829 2 84 1 sky130_fd_sc_hd__and4b_2 $T=207460 106080 0 0 $X=207270 $Y=105840
X2813 1 2 117 119 120 829 2 94 1 sky130_fd_sc_hd__and4b_2 $T=207920 89760 0 0 $X=207730 $Y=89520
X2814 1 2 117 119 120 848 2 48 1 sky130_fd_sc_hd__and4b_2 $T=210220 95200 0 0 $X=210030 $Y=94960
X2815 1 2 117 119 120 841 2 15 1 sky130_fd_sc_hd__and4b_2 $T=210220 106080 1 0 $X=210030 $Y=103120
X2816 1 2 119 117 120 841 2 23 1 sky130_fd_sc_hd__and4b_2 $T=210220 111520 0 0 $X=210030 $Y=111280
X2817 1 2 119 117 120 848 2 60 1 sky130_fd_sc_hd__and4b_2 $T=216660 100640 1 0 $X=216470 $Y=97680
X2818 1 2 119 117 120 855 2 87 1 sky130_fd_sc_hd__and4b_2 $T=216660 106080 1 0 $X=216470 $Y=103120
X2819 1 2 120 119 117 848 2 144 1 sky130_fd_sc_hd__and4b_2 $T=218960 95200 0 0 $X=218770 $Y=94960
X2820 1 2 120 119 117 855 2 100 1 sky130_fd_sc_hd__and4b_2 $T=220800 100640 0 0 $X=220610 $Y=100400
X2821 1 2 117 119 120 862 2 146 1 sky130_fd_sc_hd__and4b_2 $T=221260 89760 0 0 $X=221070 $Y=89520
X2822 1 2 117 119 120 855 2 109 1 sky130_fd_sc_hd__and4b_2 $T=224940 100640 0 0 $X=224750 $Y=100400
X2823 1 2 120 119 117 862 2 77 1 sky130_fd_sc_hd__and4b_2 $T=225400 89760 0 0 $X=225210 $Y=89520
X2824 1 2 117 119 120 865 2 76 1 sky130_fd_sc_hd__and4b_2 $T=225860 111520 0 0 $X=225670 $Y=111280
X2825 1 2 119 117 120 862 2 79 1 sky130_fd_sc_hd__and4b_2 $T=230460 95200 0 0 $X=230270 $Y=94960
X2826 1 2 125 124 123 126 2 865 1 sky130_fd_sc_hd__and4b_2 $T=230460 106080 0 0 $X=230270 $Y=105840
X2827 1 2 120 119 117 865 2 55 1 sky130_fd_sc_hd__and4b_2 $T=230460 111520 0 0 $X=230270 $Y=111280
X2828 1 2 119 117 120 865 2 129 1 sky130_fd_sc_hd__and4b_2 $T=231380 111520 1 0 $X=231190 $Y=108560
X2829 1 2 117 119 120 829 2 71 1 sky130_fd_sc_hd__and4_2 $T=201940 106080 1 0 $X=201750 $Y=103120
X2830 1 2 117 119 120 121 2 103 1 sky130_fd_sc_hd__and4_2 $T=202400 111520 1 0 $X=202210 $Y=108560
X2831 1 2 117 119 120 814 2 130 1 sky130_fd_sc_hd__and4_2 $T=202860 100640 1 0 $X=202670 $Y=97680
X2832 1 2 117 119 120 841 2 67 1 sky130_fd_sc_hd__and4_2 $T=211600 106080 0 0 $X=211410 $Y=105840
X2833 1 2 117 119 120 848 2 107 1 sky130_fd_sc_hd__and4_2 $T=212520 100640 1 0 $X=212330 $Y=97680
X2834 1 2 123 124 125 126 2 855 1 sky130_fd_sc_hd__and4_2 $T=220340 106080 0 0 $X=220150 $Y=105840
X2835 1 2 117 119 120 862 2 145 1 sky130_fd_sc_hd__and4_2 $T=220800 100640 1 0 $X=220610 $Y=97680
X2836 1 2 117 119 120 855 2 83 1 sky130_fd_sc_hd__and4_2 $T=220800 111520 0 0 $X=220610 $Y=111280
X2837 1 2 117 119 120 865 2 93 1 sky130_fd_sc_hd__and4_2 $T=234600 111520 0 0 $X=234410 $Y=111280
X2838 1 2 117 119 120 121 2 104 1 sky130_fd_sc_hd__nor4b_2 $T=192280 111520 0 0 $X=192090 $Y=111280
X2839 1 2 117 119 120 814 2 106 1 sky130_fd_sc_hd__nor4b_2 $T=193200 106080 0 0 $X=193010 $Y=105840
X2840 1 2 123 124 125 126 2 814 1 sky130_fd_sc_hd__nor4b_2 $T=196420 106080 1 0 $X=196230 $Y=103120
X2841 1 2 117 119 120 829 2 127 1 sky130_fd_sc_hd__nor4b_2 $T=202400 89760 0 0 $X=202210 $Y=89520
X2842 1 2 117 119 120 841 2 132 1 sky130_fd_sc_hd__nor4b_2 $T=204240 100640 0 0 $X=204050 $Y=100400
X2843 1 2 117 119 120 848 2 137 1 sky130_fd_sc_hd__nor4b_2 $T=212520 89760 0 0 $X=212330 $Y=89520
X2844 1 2 117 119 120 855 2 134 1 sky130_fd_sc_hd__nor4b_2 $T=215280 100640 0 0 $X=215090 $Y=100400
X2845 1 2 117 119 120 862 2 150 1 sky130_fd_sc_hd__nor4b_2 $T=224480 95200 1 0 $X=224290 $Y=92240
X2846 1 2 117 119 120 865 2 140 1 sky130_fd_sc_hd__nor4b_2 $T=226780 106080 1 0 $X=226590 $Y=103120
X2847 1 2 117 120 121 119 2 58 1 sky130_fd_sc_hd__and4bb_2 $T=189060 111520 1 0 $X=188870 $Y=108560
X2848 1 2 117 120 814 119 2 22 1 sky130_fd_sc_hd__and4bb_2 $T=189520 100640 1 0 $X=189330 $Y=97680
X2849 1 2 120 117 121 119 2 122 1 sky130_fd_sc_hd__and4bb_2 $T=193660 111520 1 0 $X=193470 $Y=108560
X2850 1 2 120 117 814 119 2 21 1 sky130_fd_sc_hd__and4bb_2 $T=194120 100640 1 0 $X=193930 $Y=97680
X2851 1 2 120 119 814 117 2 28 1 sky130_fd_sc_hd__and4bb_2 $T=194120 100640 0 0 $X=193930 $Y=100400
X2852 1 2 120 117 829 119 2 42 1 sky130_fd_sc_hd__and4bb_2 $T=202400 95200 1 0 $X=202210 $Y=92240
X2853 1 2 120 119 829 117 2 37 1 sky130_fd_sc_hd__and4bb_2 $T=203780 95200 0 0 $X=203590 $Y=94960
X2854 1 2 120 119 841 117 2 43 1 sky130_fd_sc_hd__and4bb_2 $T=205620 106080 1 0 $X=205430 $Y=103120
X2855 1 2 117 120 841 119 2 131 1 sky130_fd_sc_hd__and4bb_2 $T=205620 111520 0 0 $X=205430 $Y=111280
X2856 1 2 117 120 829 119 2 36 1 sky130_fd_sc_hd__and4bb_2 $T=207000 95200 1 0 $X=206810 $Y=92240
X2857 1 2 125 124 126 123 2 841 1 sky130_fd_sc_hd__and4bb_2 $T=207920 111520 1 0 $X=207730 $Y=108560
X2858 1 2 120 117 841 119 2 41 1 sky130_fd_sc_hd__and4bb_2 $T=209760 100640 0 0 $X=209570 $Y=100400
X2859 1 2 117 120 848 119 2 135 1 sky130_fd_sc_hd__and4bb_2 $T=211600 95200 1 0 $X=211410 $Y=92240
X2860 1 2 120 119 848 117 2 138 1 sky130_fd_sc_hd__and4bb_2 $T=214360 95200 0 0 $X=214170 $Y=94960
X2861 1 2 123 125 126 124 2 848 1 sky130_fd_sc_hd__and4bb_2 $T=215740 106080 0 0 $X=215550 $Y=105840
X2862 1 2 120 119 855 117 2 141 1 sky130_fd_sc_hd__and4bb_2 $T=216200 111520 0 0 $X=216010 $Y=111280
X2863 1 2 120 117 848 119 2 142 1 sky130_fd_sc_hd__and4bb_2 $T=216660 95200 1 0 $X=216470 $Y=92240
X2864 1 2 120 117 855 119 2 143 1 sky130_fd_sc_hd__and4bb_2 $T=216660 111520 1 0 $X=216470 $Y=108560
X2865 1 2 117 120 855 119 2 108 1 sky130_fd_sc_hd__and4bb_2 $T=221260 111520 1 0 $X=221070 $Y=108560
X2866 1 2 117 120 865 119 2 46 1 sky130_fd_sc_hd__and4bb_2 $T=222180 106080 1 0 $X=221990 $Y=103120
X2867 1 2 117 120 862 119 2 148 1 sky130_fd_sc_hd__and4bb_2 $T=224020 95200 0 0 $X=223830 $Y=94960
X2868 1 2 120 117 862 119 2 12 1 sky130_fd_sc_hd__and4bb_2 $T=224480 100640 1 0 $X=224290 $Y=97680
X2869 1 2 125 123 126 124 2 862 1 sky130_fd_sc_hd__and4bb_2 $T=225400 106080 0 0 $X=225210 $Y=105840
X2870 1 2 120 119 865 117 2 16 1 sky130_fd_sc_hd__and4bb_2 $T=226780 111520 1 0 $X=226590 $Y=108560
X2871 1 2 120 119 862 117 2 151 1 sky130_fd_sc_hd__and4bb_2 $T=229080 100640 1 0 $X=228890 $Y=97680
X2872 1 2 120 117 865 119 2 153 1 sky130_fd_sc_hd__and4bb_2 $T=230460 100640 0 0 $X=230270 $Y=100400
X2873 1 2 454 5 478 478 451 17 ICV_68 $T=12880 95200 0 0 $X=12690 $Y=94960
X2874 1 2 510 4 515 524 508 17 ICV_68 $T=50600 78880 1 0 $X=50410 $Y=75920
X2875 1 2 51 27 574 574 54 34 ICV_68 $T=64400 111520 0 0 $X=64210 $Y=111280
X2876 1 2 51 6 576 576 54 18 ICV_68 $T=65780 106080 0 0 $X=65590 $Y=105840
X2877 1 2 610 6 622 601 563 11 ICV_68 $T=90160 100640 1 0 $X=89970 $Y=97680
X2878 1 2 610 25 623 622 68 18 ICV_68 $T=90160 100640 0 0 $X=89970 $Y=100400
X2879 1 2 633 26 672 677 644 34 ICV_68 $T=114540 106080 1 0 $X=114350 $Y=103120
X2880 1 2 649 5 669 666 643 32 ICV_68 $T=118680 89760 1 0 $X=118490 $Y=86800
X2881 1 2 675 25 715 715 658 33 ICV_68 $T=137540 78880 1 0 $X=137350 $Y=75920
X2882 1 2 97 26 770 770 102 32 ICV_68 $T=162380 57120 1 0 $X=162190 $Y=54160
X2883 1 2 883 185 936 931 892 192 ICV_68 $T=258520 57120 0 0 $X=258330 $Y=56880
X2884 1 2 1033 184 1051 1051 1039 192 ICV_68 $T=314640 78880 1 0 $X=314450 $Y=75920
X2885 1 2 215 175 1080 1080 217 187 ICV_68 $T=327520 111520 0 0 $X=327330 $Y=111280
X2886 1 2 1102 166 1134 1118 1101 180 ICV_68 $T=356960 62560 1 0 $X=356770 $Y=59600
X2887 1 2 1239 166 1289 1289 1246 171 ICV_68 $T=433320 89760 0 0 $X=433130 $Y=89520
X2888 1 2 1292 258 1309 1309 1311 269 ICV_68 $T=441140 78880 1 0 $X=440950 $Y=75920
X2889 1 2 1292 265 1364 1364 1311 275 ICV_68 $T=468740 73440 0 0 $X=468550 $Y=73200
X2890 1 2 1382 283 1395 1395 1399 294 ICV_68 $T=483460 89760 1 0 $X=483270 $Y=86800
X2891 1 2 1375 258 1396 1396 1389 269 ICV_68 $T=483460 100640 1 0 $X=483270 $Y=97680
X2892 1 2 1375 262 1421 1421 1389 273 ICV_68 $T=496800 106080 0 0 $X=496610 $Y=105840
X2893 1 2 1491 258 1509 1509 1512 269 ICV_68 $T=539120 73440 0 0 $X=538930 $Y=73200
X2894 1 2 1554 259 1566 1562 1546 277 ICV_68 $T=567180 78880 1 0 $X=566990 $Y=75920
X2895 1 2 1637 259 1681 1681 1657 267 ICV_68 $T=623300 78880 1 0 $X=623110 $Y=75920
X2896 1 2 376 305 1737 1737 379 288 ICV_68 $T=651360 51680 1 0 $X=651170 $Y=48720
X2897 1 2 1753 283 1762 1762 1748 294 ICV_68 $T=665160 68000 0 0 $X=664970 $Y=67760
X2898 1 2 1754 299 1791 1791 386 307 ICV_68 $T=679420 111520 1 0 $X=679230 $Y=108560
X2899 1 2 1782 302 1802 1802 1798 309 ICV_68 $T=683100 57120 0 0 $X=682910 $Y=56880
X2900 1 2 1808 287 1814 1821 1816 288 ICV_68 $T=693220 73440 0 0 $X=693030 $Y=73200
X2901 1 2 1817 299 1851 1851 1838 307 ICV_68 $T=707940 100640 1 0 $X=707750 $Y=97680
X2902 1 2 452 5 462 ICV_69 $T=10580 68000 1 0 $X=10390 $Y=65040
X2903 1 2 453 5 464 ICV_69 $T=10580 84320 1 0 $X=10390 $Y=81360
X2904 1 2 35 26 517 ICV_69 $T=38640 51680 1 0 $X=38450 $Y=48720
X2905 1 2 510 27 520 ICV_69 $T=38640 78880 1 0 $X=38450 $Y=75920
X2906 1 2 45 6 575 ICV_69 $T=65320 57120 1 0 $X=65130 $Y=54160
X2907 1 2 85 24 704 ICV_69 $T=128340 51680 0 0 $X=128150 $Y=51440
X2908 1 2 675 4 705 ICV_69 $T=136620 73440 0 0 $X=136430 $Y=73200
X2909 1 2 732 27 750 ICV_69 $T=150880 78880 1 0 $X=150690 $Y=75920
X2910 1 2 97 6 752 ICV_69 $T=151800 51680 0 0 $X=151610 $Y=51440
X2911 1 2 732 5 771 ICV_69 $T=162380 78880 1 0 $X=162190 $Y=75920
X2912 1 2 112 8 128 ICV_69 $T=198260 51680 1 0 $X=198070 $Y=48720
X2913 1 2 881 157 894 ICV_69 $T=235060 106080 1 0 $X=234870 $Y=103120
X2914 1 2 207 156 1010 ICV_69 $T=291180 111520 1 0 $X=290990 $Y=108560
X2915 1 2 1020 168 1063 ICV_69 $T=318780 84320 1 0 $X=318590 $Y=81360
X2916 1 2 1034 158 1064 ICV_69 $T=318780 95200 1 0 $X=318590 $Y=92240
X2917 1 2 1159 186 234 ICV_69 $T=375360 51680 1 0 $X=375170 $Y=48720
X2918 1 2 249 167 1294 ICV_69 $T=434240 51680 0 0 $X=434050 $Y=51440
X2919 1 2 1306 264 1330 ICV_69 $T=448960 106080 1 0 $X=448770 $Y=103120
X2920 1 2 290 287 1432 ICV_69 $T=504620 111520 1 0 $X=504430 $Y=108560
X2921 1 2 318 257 1460 ICV_69 $T=513360 106080 0 0 $X=513170 $Y=105840
X2922 1 2 1471 258 1487 ICV_69 $T=528540 68000 1 0 $X=528350 $Y=65040
X2923 1 2 1473 262 1492 ICV_69 $T=529460 78880 0 0 $X=529270 $Y=78640
X2924 1 2 1491 265 1521 ICV_69 $T=543260 78880 1 0 $X=543070 $Y=75920
X2925 1 2 1506 257 1522 ICV_69 $T=543260 84320 1 0 $X=543070 $Y=81360
X2926 1 2 1506 258 1523 ICV_69 $T=543260 89760 1 0 $X=543070 $Y=86800
X2927 1 2 1554 264 1572 ICV_69 $T=569940 84320 0 0 $X=569750 $Y=84080
X2928 1 2 1554 266 1595 ICV_69 $T=585580 78880 0 0 $X=585390 $Y=78640
X2929 1 2 1592 272 1631 ICV_69 $T=598920 84320 0 0 $X=598730 $Y=84080
X2930 1 2 1591 259 1644 ICV_69 $T=607200 106080 0 0 $X=607010 $Y=105840
X2931 1 2 1736 301 388 ICV_69 $T=669760 57120 0 0 $X=669570 $Y=56880
X2932 1 2 1776 283 1837 ICV_69 $T=697820 95200 0 0 $X=697630 $Y=94960
X2933 1 2 37 13 513 513 512 81 ICV_74 $T=39100 100640 1 0 $X=38910 $Y=97680
X2934 1 2 42 13 539 539 540 81 ICV_74 $T=51980 68000 0 0 $X=51790 $Y=67760
X2935 1 2 76 13 654 654 633 81 ICV_74 $T=111780 111520 1 0 $X=111590 $Y=108560
X2936 1 2 77 13 656 656 671 81 ICV_74 $T=112240 73440 1 0 $X=112050 $Y=70480
X2937 1 2 87 13 697 697 675 81 ICV_74 $T=130640 84320 0 0 $X=130450 $Y=84080
X2938 1 2 109 13 782 782 790 81 ICV_74 $T=172040 62560 1 0 $X=171850 $Y=59600
X2939 1 2 129 13 839 839 847 81 ICV_74 $T=205620 84320 1 0 $X=205430 $Y=81360
X2940 1 2 151 152 876 876 881 81 ICV_74 $T=230000 95200 1 0 $X=229810 $Y=92240
X2941 1 2 28 154 879 879 885 81 ICV_74 $T=230920 73440 0 0 $X=230730 $Y=73200
X2942 1 2 36 154 932 932 928 81 ICV_74 $T=259900 78880 1 0 $X=259710 $Y=75920
X2943 1 2 94 154 1014 1014 1020 81 ICV_74 $T=300840 89760 1 0 $X=300650 $Y=86800
X2944 1 2 146 154 1016 1016 214 81 ICV_74 $T=302220 51680 1 0 $X=302030 $Y=48720
X2945 1 2 122 152 1073 1073 220 81 ICV_74 $T=331200 106080 0 0 $X=331010 $Y=105840
X2946 1 2 137 152 1165 1172 1180 81 ICV_74 $T=375820 89760 1 0 $X=375630 $Y=86800
X2947 1 2 140 154 1251 1251 249 81 ICV_74 $T=417680 51680 0 0 $X=417490 $Y=51440
X2948 1 2 279 261 1346 1346 1304 415 ICV_74 $T=463680 84320 0 0 $X=463490 $Y=84080
X2949 1 2 289 261 1367 1369 282 415 ICV_74 $T=474720 62560 1 0 $X=474530 $Y=59600
X2950 1 2 322 261 1464 1464 1473 415 ICV_74 $T=519340 89760 0 0 $X=519150 $Y=89520
X2951 1 2 281 293 1494 1494 331 415 ICV_74 $T=534980 57120 1 0 $X=534790 $Y=54160
X2952 1 2 366 261 1642 1642 1646 415 ICV_74 $T=610880 57120 1 0 $X=610690 $Y=54160
X2953 1 2 370 261 1676 1676 1692 415 ICV_74 $T=626060 73440 0 0 $X=625870 $Y=73200
X2954 1 2 372 261 1678 1678 1694 415 ICV_74 $T=628360 57120 1 0 $X=628170 $Y=54160
X2955 1 2 321 293 1813 1813 1807 415 ICV_74 $T=694140 62560 1 0 $X=693950 $Y=59600
X2956 1 2 370 293 1847 1847 1866 415 ICV_74 $T=711160 62560 0 0 $X=710970 $Y=62320
X2957 1 2 7 9 11 10 6 480 475 9 20 ICV_84 $T=10580 51680 0 0 $X=10390 $Y=51440
X2958 1 2 562 47 17 45 25 580 575 53 18 ICV_84 $T=63020 57120 0 0 $X=62830 $Y=56880
X2959 1 2 587 586 11 591 4 609 605 586 33 ICV_84 $T=78660 68000 1 0 $X=78470 $Y=65040
X2960 1 2 613 615 20 607 6 637 640 615 33 ICV_84 $T=92920 84320 0 0 $X=92730 $Y=84080
X2961 1 2 701 86 18 679 27 721 719 86 17 ICV_84 $T=134780 106080 1 0 $X=134590 $Y=103120
X2962 1 2 905 890 177 885 186 925 924 890 194 ICV_84 $T=245640 68000 1 0 $X=245450 $Y=65040
X2963 1 2 1057 1039 177 1033 164 1079 1079 1039 169 ICV_84 $T=323380 73440 0 0 $X=323190 $Y=73200
X2964 1 2 1147 1110 194 1180 184 1193 1193 1199 192 ICV_84 $T=381340 89760 0 0 $X=381150 $Y=89520
X2965 1 2 1209 1210 180 1188 183 1230 1230 1210 193 ICV_84 $T=400200 68000 0 0 $X=400010 $Y=67760
X2966 1 2 1229 1228 195 1204 168 1249 1249 1228 177 ICV_84 $T=408020 57120 0 0 $X=407830 $Y=56880
X2967 1 2 1232 1210 194 1239 183 1257 1260 1261 177 ICV_84 $T=410780 84320 0 0 $X=410590 $Y=84080
X2968 1 2 1433 315 304 1409 299 1457 1426 1428 303 ICV_84 $T=508300 57120 1 0 $X=508110 $Y=54160
X2969 1 2 1469 323 288 320 287 1497 328 323 307 ICV_84 $T=526240 51680 1 0 $X=526050 $Y=48720
X2970 1 2 1602 1582 267 1616 265 1623 1623 1625 275 ICV_84 $T=592940 62560 1 0 $X=592750 $Y=59600
X2971 1 2 1743 1746 288 1731 283 1759 1759 1746 294 ICV_84 $T=659640 95200 0 0 $X=659450 $Y=94960
X2972 1 2 1756 384 288 1736 292 1777 1777 384 300 ICV_84 $T=666540 51680 1 0 $X=666350 $Y=48720
X2973 1 2 1861 397 303 1865 292 1876 1876 1874 300 ICV_84 $T=715760 100640 0 0 $X=715570 $Y=100400
X2974 1 2 510 6 544 ICV_85 $T=48300 84320 1 0 $X=48110 $Y=81360
X2975 1 2 881 156 889 ICV_85 $T=233680 100640 1 0 $X=233490 $Y=97680
X2976 1 2 883 168 902 ICV_85 $T=237360 57120 0 0 $X=237170 $Y=56880
X2977 1 2 197 167 980 ICV_85 $T=276920 51680 1 0 $X=276730 $Y=48720
X2978 1 2 959 167 1003 ICV_85 $T=289800 84320 1 0 $X=289610 $Y=81360
X2979 1 2 219 166 1103 ICV_85 $T=339480 51680 1 0 $X=339290 $Y=48720
X2980 1 2 1102 185 1119 ICV_85 $T=345460 62560 1 0 $X=345270 $Y=59600
X2981 1 2 1159 164 1173 ICV_85 $T=373980 57120 1 0 $X=373790 $Y=54160
X2982 1 2 249 166 1313 ICV_85 $T=443440 51680 0 0 $X=443250 $Y=51440
X2983 1 2 1306 265 1347 ICV_85 $T=458160 106080 1 0 $X=457970 $Y=103120
X2984 1 2 1418 272 1434 ICV_85 $T=502320 68000 1 0 $X=502130 $Y=65040
X2985 1 2 318 262 1465 ICV_85 $T=513820 111520 1 0 $X=513630 $Y=108560
X2986 1 2 1506 265 1549 ICV_85 $T=556140 84320 0 0 $X=555950 $Y=84080
X2987 1 2 1592 258 1630 ICV_85 $T=598460 84320 1 0 $X=598270 $Y=81360
X2988 1 2 1664 264 1693 ICV_85 $T=626520 106080 1 0 $X=626330 $Y=103120
X2989 1 2 1807 283 1833 ICV_85 $T=696440 57120 0 0 $X=696250 $Y=56880
X2990 1 2 514 35 81 ICV_86 $T=38640 51680 0 0 $X=38450 $Y=51440
X2991 1 2 538 45 81 ICV_86 $T=50600 57120 1 0 $X=50410 $Y=54160
X2992 1 2 556 560 81 ICV_86 $T=58880 89760 1 0 $X=58690 $Y=86800
X2993 1 2 612 66 81 ICV_86 $T=90160 111520 0 0 $X=89970 $Y=111280
X2994 1 2 919 926 81 ICV_86 $T=252080 100640 1 0 $X=251890 $Y=97680
X2995 1 2 976 984 81 ICV_86 $T=280140 78880 1 0 $X=279950 $Y=75920
X2996 1 2 230 231 81 ICV_86 $T=364320 111520 1 0 $X=364130 $Y=108560
X2997 1 2 1237 1239 81 ICV_86 $T=410320 89760 0 0 $X=410130 $Y=89520
X2998 1 2 1367 1301 415 ICV_86 $T=475180 62560 0 0 $X=474990 $Y=62320
X2999 1 2 1374 1382 415 ICV_86 $T=476560 95200 1 0 $X=476370 $Y=92240
X3000 1 2 1571 338 415 ICV_86 $T=573620 111520 1 0 $X=573430 $Y=108560
X3001 1 2 1587 1593 415 ICV_86 $T=581440 100640 1 0 $X=581250 $Y=97680
X3002 1 2 1638 364 415 ICV_86 $T=605820 51680 0 0 $X=605630 $Y=51440
X3003 1 2 1682 1690 415 ICV_86 $T=627440 78880 0 0 $X=627250 $Y=78640
X3004 1 2 1744 1754 415 ICV_86 $T=657340 111520 1 0 $X=657150 $Y=108560
X3005 1 2 1780 1782 415 ICV_86 $T=677120 78880 1 0 $X=676930 $Y=75920
X3006 1 2 472 473 11 22 13 481 ICV_87 $T=19320 84320 0 0 $X=19130 $Y=84080
X3007 1 2 19 14 20 23 13 484 ICV_87 $T=20240 111520 1 0 $X=20050 $Y=108560
X3008 1 2 603 54 30 65 13 614 ICV_87 $T=87860 106080 1 0 $X=87670 $Y=103120
X3009 1 2 762 740 18 107 69 110 ICV_87 $T=166520 111520 0 0 $X=166330 $Y=111280
X3010 1 2 875 155 32 41 154 163 ICV_87 $T=231380 51680 0 0 $X=231190 $Y=51440
X3011 1 2 937 940 194 42 154 947 ICV_87 $T=264960 68000 1 0 $X=264770 $Y=65040
X3012 1 2 1072 1038 195 71 154 1087 ICV_87 $T=332580 84320 0 0 $X=332390 $Y=84080
X3013 1 2 1106 1100 193 100 154 1105 ICV_87 $T=347300 68000 0 0 $X=347110 $Y=67760
X3014 1 2 1112 1074 178 138 152 1122 ICV_87 $T=350980 100640 0 0 $X=350790 $Y=100400
X3015 1 2 1179 1157 169 127 154 1207 ICV_87 $T=391920 73440 0 0 $X=391730 $Y=73200
X3016 1 2 237 232 178 140 152 238 ICV_87 $T=391920 111520 0 0 $X=391730 $Y=111280
X3017 1 2 1234 1210 195 134 154 1253 ICV_87 $T=415840 68000 0 0 $X=415650 $Y=67760
X3018 1 2 1350 1331 268 285 261 1353 ICV_87 $T=465980 95200 0 0 $X=465790 $Y=94960
X3019 1 2 1362 1331 280 295 293 1374 ICV_87 $T=474260 95200 0 0 $X=474070 $Y=94960
X3020 1 2 1392 1399 296 308 261 1406 ICV_87 $T=489900 95200 0 0 $X=489710 $Y=94960
X3021 1 2 1580 1551 275 348 261 1575 ICV_87 $T=583280 100640 0 0 $X=583090 $Y=100400
X3022 1 2 1588 1582 268 355 261 1594 ICV_87 $T=589720 57120 1 0 $X=589530 $Y=54160
.ENDS
***************************************
.SUBCKT ICV_89 1 2
** N=2 EP=2 IP=4 FDC=6
*.SEEDPROM
X0 1 2 ICV_10 $T=11040 0 0 0 $X=10850 $Y=-240
X1 1 2 ICV_11 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_90 1 2
** N=2 EP=2 IP=4 FDC=8
*.SEEDPROM
X0 1 2 ICV_11 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 ICV_11 $T=11040 0 0 0 $X=10850 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_91 1 2
** N=2 EP=2 IP=6 FDC=2
*.SEEDPROM
X0 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=0 0 0 0 $X=-190 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_92 1 2
** N=2 EP=2 IP=4 FDC=10
*.SEEDPROM
X0 1 2 ICV_90 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 ICV_91 $T=22080 0 0 0 $X=21890 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_93 1 2
** N=2 EP=2 IP=4 FDC=20
*.SEEDPROM
X0 1 2 ICV_92 $T=0 0 0 0 $X=-190 $Y=-240
X1 1 2 ICV_92 $T=28060 0 0 0 $X=27870 $Y=-240
.ENDS
***************************************
.SUBCKT ICV_94 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 253
** N=967 EP=247 IP=8822 FDC=23185
*.SEEDPROM
X0 1 2 Dpar a=1186.32 p=1481.49 m=1 $[nwdiode] $X=5330 $Y=10690 $D=191
X1 1 2 Dpar a=2091.77 p=1483.94 m=1 $[nwdiode] $X=5330 $Y=14905 $D=191
X2 1 2 Dpar a=2090.95 p=1484.94 m=1 $[nwdiode] $X=5330 $Y=20345 $D=191
X3 1 2 Dpar a=2090.95 p=1484.94 m=1 $[nwdiode] $X=5330 $Y=25785 $D=191
X4 1 2 Dpar a=2091.12 p=1484.74 m=1 $[nwdiode] $X=5330 $Y=31225 $D=191
X5 1 2 Dpar a=2090.55 p=1485.44 m=1 $[nwdiode] $X=5330 $Y=36665 $D=191
X6 1 2 Dpar a=2090.95 p=1484.94 m=1 $[nwdiode] $X=5330 $Y=42105 $D=191
X7 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 13600 1 0 $X=5330 $Y=10640
X8 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 13600 0 0 $X=5330 $Y=13360
X9 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 19040 1 0 $X=5330 $Y=16080
X10 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 19040 0 0 $X=5330 $Y=18800
X11 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 24480 1 0 $X=5330 $Y=21520
X12 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 24480 0 0 $X=5330 $Y=24240
X13 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 29920 1 0 $X=5330 $Y=26960
X14 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 29920 0 0 $X=5330 $Y=29680
X15 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 35360 1 0 $X=5330 $Y=32400
X16 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 35360 0 0 $X=5330 $Y=35120
X17 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 40800 1 0 $X=5330 $Y=37840
X18 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 40800 0 0 $X=5330 $Y=40560
X19 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 46240 1 0 $X=5330 $Y=43280
X20 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=5520 46240 0 0 $X=5330 $Y=46000
X21 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=34040 13600 0 0 $X=33850 $Y=13360
X22 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=68080 40800 1 0 $X=67890 $Y=37840
X23 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=76360 24480 1 0 $X=76170 $Y=21520
X24 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=88320 29920 0 0 $X=88130 $Y=29680
X25 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=114080 46240 1 0 $X=113890 $Y=43280
X26 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=121440 40800 1 0 $X=121250 $Y=37840
X27 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=175260 46240 1 0 $X=175070 $Y=43280
X28 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=196880 13600 1 0 $X=196690 $Y=10640
X29 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=200560 35360 0 0 $X=200370 $Y=35120
X30 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=202400 19040 0 0 $X=202210 $Y=18800
X31 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=214820 35360 1 0 $X=214630 $Y=32400
X32 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=230460 19040 0 0 $X=230270 $Y=18800
X33 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=250240 24480 0 0 $X=250050 $Y=24240
X34 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=264040 29920 0 0 $X=263850 $Y=29680
X35 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=284740 19040 0 0 $X=284550 $Y=18800
X36 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=293940 29920 0 0 $X=293750 $Y=29680
X37 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=300840 35360 1 0 $X=300650 $Y=32400
X38 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=340400 29920 1 0 $X=340210 $Y=26960
X39 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=341320 35360 1 0 $X=341130 $Y=32400
X40 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=342700 40800 1 0 $X=342510 $Y=37840
X41 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=351440 35360 0 0 $X=351250 $Y=35120
X42 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=354660 19040 0 0 $X=354470 $Y=18800
X43 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=368920 13600 0 0 $X=368730 $Y=13360
X44 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=369840 35360 1 0 $X=369650 $Y=32400
X45 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=383180 35360 1 0 $X=382990 $Y=32400
X46 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=396980 40800 0 0 $X=396790 $Y=40560
X47 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=410320 29920 0 0 $X=410130 $Y=29680
X48 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=453100 46240 0 0 $X=452910 $Y=46000
X49 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=462300 40800 1 0 $X=462110 $Y=37840
X50 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=483000 29920 0 0 $X=482810 $Y=29680
X51 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=506460 29920 1 0 $X=506270 $Y=26960
X52 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=516120 40800 1 0 $X=515930 $Y=37840
X53 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=549240 46240 1 0 $X=549050 $Y=43280
X54 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=558900 29920 1 0 $X=558710 $Y=26960
X55 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=561660 46240 1 0 $X=561470 $Y=43280
X56 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=565340 40800 0 0 $X=565150 $Y=40560
X57 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=608120 40800 0 0 $X=607930 $Y=40560
X58 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=620540 40800 1 0 $X=620350 $Y=37840
X59 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=621460 35360 0 0 $X=621270 $Y=35120
X60 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=663780 40800 1 0 $X=663590 $Y=37840
X61 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=677580 46240 0 0 $X=677390 $Y=46000
X62 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=690000 29920 0 0 $X=689810 $Y=29680
X63 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=713000 24480 0 0 $X=712810 $Y=24240
X64 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=718980 46240 0 0 $X=718790 $Y=46000
X65 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=733700 35360 0 0 $X=733510 $Y=35120
X66 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 13600 0 180 $X=742710 $Y=10640
X67 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 13600 1 180 $X=742710 $Y=13360
X68 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 19040 0 180 $X=742710 $Y=16080
X69 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 19040 1 180 $X=742710 $Y=18800
X70 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 24480 0 180 $X=742710 $Y=21520
X71 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 24480 1 180 $X=742710 $Y=24240
X72 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 29920 0 180 $X=742710 $Y=26960
X73 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 29920 1 180 $X=742710 $Y=29680
X74 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 35360 0 180 $X=742710 $Y=32400
X75 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 35360 1 180 $X=742710 $Y=35120
X76 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 40800 0 180 $X=742710 $Y=37840
X77 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 40800 1 180 $X=742710 $Y=40560
X78 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 46240 0 180 $X=742710 $Y=43280
X79 1 2 1 2 sky130_fd_sc_hd__decap_3 $T=744280 46240 1 180 $X=742710 $Y=46000
X164 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 24480 1 0 $X=17750 $Y=21520
X165 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=17940 29920 1 0 $X=17750 $Y=26960
X166 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=50600 40800 0 0 $X=50410 $Y=40560
X167 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=67620 40800 0 0 $X=67430 $Y=40560
X168 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=73600 40800 0 0 $X=73410 $Y=40560
X169 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=83720 19040 1 0 $X=83530 $Y=16080
X170 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=91540 46240 1 0 $X=91350 $Y=43280
X171 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=96600 24480 1 0 $X=96410 $Y=21520
X172 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=118220 29920 0 0 $X=118030 $Y=29680
X173 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=125580 13600 0 0 $X=125390 $Y=13360
X174 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=159620 40800 0 0 $X=159430 $Y=40560
X175 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=169280 24480 1 0 $X=169090 $Y=21520
X176 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=184920 24480 1 0 $X=184730 $Y=21520
X177 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=186300 29920 1 0 $X=186110 $Y=26960
X178 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=186300 35360 1 0 $X=186110 $Y=32400
X179 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=188140 29920 0 0 $X=187950 $Y=29680
X180 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=214360 19040 1 0 $X=214170 $Y=16080
X181 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=230460 46240 0 0 $X=230270 $Y=46000
X182 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=239660 19040 1 0 $X=239470 $Y=16080
X183 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=244720 46240 1 0 $X=244530 $Y=43280
X184 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=248860 19040 1 0 $X=248670 $Y=16080
X185 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=256220 35360 1 0 $X=256030 $Y=32400
X186 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=266340 19040 1 0 $X=266150 $Y=16080
X187 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=270480 13600 1 0 $X=270290 $Y=10640
X188 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=284280 24480 0 0 $X=284090 $Y=24240
X189 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=284280 29920 0 0 $X=284090 $Y=29680
X190 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=298540 19040 1 0 $X=298350 $Y=16080
X191 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=298540 40800 1 0 $X=298350 $Y=37840
X192 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=304980 19040 1 0 $X=304790 $Y=16080
X193 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=327060 40800 0 0 $X=326870 $Y=40560
X194 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=340400 29920 0 0 $X=340210 $Y=29680
X195 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=364320 24480 1 0 $X=364130 $Y=21520
X196 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=380420 40800 0 0 $X=380230 $Y=40560
X197 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=382260 46240 0 0 $X=382070 $Y=46000
X198 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=392380 40800 1 0 $X=392190 $Y=37840
X199 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=396520 13600 0 0 $X=396330 $Y=13360
X200 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=396980 29920 1 0 $X=396790 $Y=26960
X201 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=406180 35360 0 0 $X=405990 $Y=35120
X202 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=412620 46240 0 0 $X=412430 $Y=46000
X203 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=413080 46240 1 0 $X=412890 $Y=43280
X204 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=426880 40800 0 0 $X=426690 $Y=40560
X205 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=448500 19040 1 0 $X=448310 $Y=16080
X206 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=459080 13600 0 0 $X=458890 $Y=13360
X207 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=465060 46240 0 0 $X=464870 $Y=46000
X208 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=475640 24480 0 0 $X=475450 $Y=24240
X209 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=521640 35360 0 0 $X=521450 $Y=35120
X210 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=525320 29920 0 0 $X=525130 $Y=29680
X211 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=525320 35360 1 0 $X=525130 $Y=32400
X212 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=525320 46240 1 0 $X=525130 $Y=43280
X213 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=536360 24480 1 0 $X=536170 $Y=21520
X214 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=539120 35360 0 0 $X=538930 $Y=35120
X215 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=598920 35360 1 0 $X=598730 $Y=32400
X216 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=640320 40800 0 0 $X=640130 $Y=40560
X217 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=651360 24480 0 0 $X=651170 $Y=24240
X218 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=665620 35360 0 0 $X=665430 $Y=35120
X219 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=683560 46240 0 0 $X=683370 $Y=46000
X220 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=712540 35360 0 0 $X=712350 $Y=35120
X221 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=729100 46240 1 0 $X=728910 $Y=43280
X222 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 13600 0 0 $X=740870 $Y=13360
X223 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 19040 0 0 $X=740870 $Y=18800
X224 1 2 1 2 sky130_fd_sc_hd__decap_4 $T=741060 24480 0 0 $X=740870 $Y=24240
X225 1 2 ICV_3 $T=31280 46240 0 0 $X=31090 $Y=46000
X226 1 2 ICV_3 $T=74060 46240 0 0 $X=73870 $Y=46000
X227 1 2 ICV_3 $T=101660 29920 1 0 $X=101470 $Y=26960
X228 1 2 ICV_3 $T=123280 29920 1 0 $X=123090 $Y=26960
X229 1 2 ICV_3 $T=138000 24480 1 0 $X=137810 $Y=21520
X230 1 2 ICV_3 $T=155940 35360 0 0 $X=155750 $Y=35120
X231 1 2 ICV_3 $T=171580 40800 1 0 $X=171390 $Y=37840
X232 1 2 ICV_3 $T=174340 29920 0 0 $X=174150 $Y=29680
X233 1 2 ICV_3 $T=198260 40800 0 0 $X=198070 $Y=40560
X234 1 2 ICV_3 $T=216660 40800 1 0 $X=216470 $Y=37840
X235 1 2 ICV_3 $T=230460 40800 0 0 $X=230270 $Y=40560
X236 1 2 ICV_3 $T=276920 13600 1 0 $X=276730 $Y=10640
X237 1 2 ICV_3 $T=281060 35360 1 0 $X=280870 $Y=32400
X238 1 2 ICV_3 $T=300840 46240 1 0 $X=300650 $Y=43280
X239 1 2 ICV_3 $T=306820 29920 0 0 $X=306630 $Y=29680
X240 1 2 ICV_3 $T=319700 13600 1 0 $X=319510 $Y=10640
X241 1 2 ICV_3 $T=340400 19040 1 0 $X=340210 $Y=16080
X242 1 2 ICV_3 $T=354200 19040 1 0 $X=354010 $Y=16080
X243 1 2 ICV_3 $T=356960 40800 1 0 $X=356770 $Y=37840
X244 1 2 ICV_3 $T=382260 19040 1 0 $X=382070 $Y=16080
X245 1 2 ICV_3 $T=382260 29920 1 0 $X=382070 $Y=26960
X246 1 2 ICV_3 $T=382260 35360 0 0 $X=382070 $Y=35120
X247 1 2 ICV_3 $T=396060 35360 0 0 $X=395870 $Y=35120
X248 1 2 ICV_3 $T=410320 29920 1 0 $X=410130 $Y=26960
X249 1 2 ICV_3 $T=420440 29920 1 0 $X=420250 $Y=26960
X250 1 2 ICV_3 $T=434700 24480 0 0 $X=434510 $Y=24240
X251 1 2 ICV_3 $T=441140 24480 1 0 $X=440950 $Y=21520
X252 1 2 ICV_3 $T=441140 29920 1 0 $X=440950 $Y=26960
X253 1 2 ICV_3 $T=452180 40800 0 0 $X=451990 $Y=40560
X254 1 2 ICV_3 $T=508300 40800 0 0 $X=508110 $Y=40560
X255 1 2 ICV_3 $T=518420 40800 0 0 $X=518230 $Y=40560
X256 1 2 ICV_3 $T=532220 40800 0 0 $X=532030 $Y=40560
X257 1 2 ICV_3 $T=564420 46240 0 0 $X=564230 $Y=46000
X258 1 2 ICV_3 $T=579140 24480 0 0 $X=578950 $Y=24240
X259 1 2 ICV_3 $T=581440 46240 1 0 $X=581250 $Y=43280
X260 1 2 ICV_3 $T=634800 29920 0 0 $X=634610 $Y=29680
X261 1 2 ICV_3 $T=634800 40800 1 0 $X=634610 $Y=37840
X262 1 2 ICV_3 $T=646300 40800 1 0 $X=646110 $Y=37840
X263 1 2 ICV_3 $T=649060 35360 1 0 $X=648870 $Y=32400
X264 1 2 ICV_3 $T=661940 13600 1 0 $X=661750 $Y=10640
X265 1 2 ICV_3 $T=662860 46240 0 0 $X=662670 $Y=46000
X266 1 2 ICV_3 $T=667460 46240 0 0 $X=667270 $Y=46000
X267 1 2 ICV_3 $T=679420 29920 0 0 $X=679230 $Y=29680
X268 1 2 ICV_3 $T=693680 35360 1 0 $X=693490 $Y=32400
X269 1 2 ICV_3 $T=735540 40800 0 0 $X=735350 $Y=40560
X270 1 2 ICV_3 $T=740600 35360 1 0 $X=740410 $Y=32400
X271 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=33120 35360 1 0 $X=32930 $Y=32400
X272 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=34960 46240 1 0 $X=34770 $Y=43280
X273 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=48300 19040 1 0 $X=48110 $Y=16080
X274 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=58420 29920 0 0 $X=58230 $Y=29680
X275 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=73140 46240 1 0 $X=72950 $Y=43280
X276 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=86020 24480 1 0 $X=85830 $Y=21520
X277 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=90160 19040 0 0 $X=89970 $Y=18800
X278 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=101660 29920 0 0 $X=101470 $Y=29680
X279 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=115000 35360 0 0 $X=114810 $Y=35120
X280 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=125580 46240 0 0 $X=125390 $Y=46000
X281 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=142600 24480 0 0 $X=142410 $Y=24240
X282 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=146740 35360 1 0 $X=146550 $Y=32400
X283 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=155480 19040 0 0 $X=155290 $Y=18800
X284 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=170660 13600 0 0 $X=170470 $Y=13360
X285 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=182620 35360 0 0 $X=182430 $Y=35120
X286 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=185380 24480 0 0 $X=185190 $Y=24240
X287 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=205620 13600 1 0 $X=205430 $Y=10640
X288 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=209760 13600 0 0 $X=209570 $Y=13360
X289 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=212520 13600 1 0 $X=212330 $Y=10640
X290 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=226780 13600 0 0 $X=226590 $Y=13360
X291 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=228160 46240 1 0 $X=227970 $Y=43280
X292 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=230460 35360 0 0 $X=230270 $Y=35120
X293 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=251160 46240 0 0 $X=250970 $Y=46000
X294 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=254840 40800 0 0 $X=254650 $Y=40560
X295 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=282900 46240 0 0 $X=282710 $Y=46000
X296 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=284280 40800 1 0 $X=284090 $Y=37840
X297 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=286580 40800 0 0 $X=286390 $Y=40560
X298 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=298540 35360 0 0 $X=298350 $Y=35120
X299 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=300840 29920 1 0 $X=300650 $Y=26960
X300 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=302220 13600 1 0 $X=302030 $Y=10640
X301 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=356960 29920 1 0 $X=356770 $Y=26960
X302 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=395140 29920 0 0 $X=394950 $Y=29680
X303 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=409860 40800 1 0 $X=409670 $Y=37840
X304 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=415840 13600 0 0 $X=415650 $Y=13360
X305 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=438380 19040 0 0 $X=438190 $Y=18800
X306 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=441140 24480 0 0 $X=440950 $Y=24240
X307 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=441140 35360 1 0 $X=440950 $Y=32400
X308 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=451260 29920 0 0 $X=451070 $Y=29680
X309 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=451720 24480 0 0 $X=451530 $Y=24240
X310 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=465520 19040 1 0 $X=465330 $Y=16080
X311 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=465980 40800 1 0 $X=465790 $Y=37840
X312 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=483000 24480 0 0 $X=482810 $Y=24240
X313 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=497260 24480 1 0 $X=497070 $Y=21520
X314 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=536820 29920 1 0 $X=536630 $Y=26960
X315 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=538660 46240 1 0 $X=538470 $Y=43280
X316 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=549700 24480 1 0 $X=549510 $Y=21520
X317 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=553380 35360 1 0 $X=553190 $Y=32400
X318 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=577760 46240 1 0 $X=577570 $Y=43280
X319 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=578220 24480 1 0 $X=578030 $Y=21520
X320 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=578220 35360 0 0 $X=578030 $Y=35120
X321 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=590180 29920 1 0 $X=589990 $Y=26960
X322 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=596620 24480 1 0 $X=596430 $Y=21520
X323 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=606740 24480 0 0 $X=606550 $Y=24240
X324 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=620080 40800 0 0 $X=619890 $Y=40560
X325 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=632960 24480 0 0 $X=632770 $Y=24240
X326 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=633880 46240 1 0 $X=633690 $Y=43280
X327 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=651360 35360 0 0 $X=651170 $Y=35120
X328 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=672520 13600 1 0 $X=672330 $Y=10640
X329 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=683560 40800 0 0 $X=683370 $Y=40560
X330 1 2 1 2 sky130_fd_sc_hd__decap_6 $T=697820 29920 1 0 $X=697630 $Y=26960
X331 1 2 ICV_4 $T=24380 40800 1 0 $X=24190 $Y=37840
X332 1 2 ICV_4 $T=73140 13600 0 0 $X=72950 $Y=13360
X333 1 2 ICV_4 $T=114540 46240 0 0 $X=114350 $Y=46000
X334 1 2 ICV_4 $T=142600 29920 1 0 $X=142410 $Y=26960
X335 1 2 ICV_4 $T=160540 46240 1 0 $X=160350 $Y=43280
X336 1 2 ICV_4 $T=162840 13600 1 0 $X=162650 $Y=10640
X337 1 2 ICV_4 $T=195960 46240 1 0 $X=195770 $Y=43280
X338 1 2 ICV_4 $T=258520 19040 0 0 $X=258330 $Y=18800
X339 1 2 ICV_4 $T=325680 29920 0 0 $X=325490 $Y=29680
X340 1 2 ICV_4 $T=411700 40800 0 0 $X=411510 $Y=40560
X341 1 2 ICV_4 $T=460460 35360 0 0 $X=460270 $Y=35120
X342 1 2 ICV_4 $T=480700 46240 1 0 $X=480510 $Y=43280
X343 1 2 ICV_4 $T=481160 35360 1 0 $X=480970 $Y=32400
X344 1 2 ICV_4 $T=493580 40800 0 0 $X=493390 $Y=40560
X345 1 2 ICV_4 $T=553380 40800 1 0 $X=553190 $Y=37840
X346 1 2 ICV_4 $T=591560 29920 0 0 $X=591370 $Y=29680
X347 1 2 ICV_4 $T=662860 29920 0 0 $X=662670 $Y=29680
X348 1 2 ICV_4 $T=739680 29920 0 0 $X=739490 $Y=29680
X349 1 2 ICV_4 $T=739680 35360 0 0 $X=739490 $Y=35120
X350 1 2 ICV_4 $T=739680 46240 0 0 $X=739490 $Y=46000
X351 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=6900 46240 0 0 $X=6710 $Y=46000
X352 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=12420 29920 0 0 $X=12230 $Y=29680
X353 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=15640 13600 1 0 $X=15450 $Y=10640
X354 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=17940 24480 0 0 $X=17750 $Y=24240
X355 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=20240 19040 1 0 $X=20050 $Y=16080
X356 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=28980 13600 0 0 $X=28790 $Y=13360
X357 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=57960 46240 1 0 $X=57770 $Y=43280
X358 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=57960 46240 0 0 $X=57770 $Y=46000
X359 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=63940 19040 1 0 $X=63750 $Y=16080
X360 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=64400 24480 1 0 $X=64210 $Y=21520
X361 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=84640 13600 0 0 $X=84450 $Y=13360
X362 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=90160 13600 0 0 $X=89970 $Y=13360
X363 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=94300 46240 0 0 $X=94110 $Y=46000
X364 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=100280 19040 1 0 $X=100090 $Y=16080
X365 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=113620 24480 1 0 $X=113430 $Y=21520
X366 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=132480 35360 1 0 $X=132290 $Y=32400
X367 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=134780 19040 0 0 $X=134590 $Y=18800
X368 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=150880 46240 0 0 $X=150690 $Y=46000
X369 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=165600 40800 0 0 $X=165410 $Y=40560
X370 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=174340 19040 0 0 $X=174150 $Y=18800
X371 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=174340 24480 0 0 $X=174150 $Y=24240
X372 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=188600 40800 1 0 $X=188410 $Y=37840
X373 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=195040 24480 1 0 $X=194850 $Y=21520
X374 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=195960 35360 1 0 $X=195770 $Y=32400
X375 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=201020 40800 1 0 $X=200830 $Y=37840
X376 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=206540 35360 0 0 $X=206350 $Y=35120
X377 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=211140 35360 1 0 $X=210950 $Y=32400
X378 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=211140 46240 0 0 $X=210950 $Y=46000
X379 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=211600 29920 1 0 $X=211410 $Y=26960
X380 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=218960 46240 0 0 $X=218770 $Y=46000
X381 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=226320 35360 0 0 $X=226130 $Y=35120
X382 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=234140 13600 1 0 $X=233950 $Y=10640
X383 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=234600 13600 0 0 $X=234410 $Y=13360
X384 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=261280 29920 1 0 $X=261090 $Y=26960
X385 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=290720 46240 0 0 $X=290530 $Y=46000
X386 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=306360 24480 0 0 $X=306170 $Y=24240
X387 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=314640 29920 0 0 $X=314450 $Y=29680
X388 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=333040 40800 0 0 $X=332850 $Y=40560
X389 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=344080 13600 1 0 $X=343890 $Y=10640
X390 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=352820 46240 1 0 $X=352630 $Y=43280
X391 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=354660 40800 0 0 $X=354470 $Y=40560
X392 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=364320 46240 1 0 $X=364130 $Y=43280
X393 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=371220 29920 1 0 $X=371030 $Y=26960
X394 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=379500 35360 1 0 $X=379310 $Y=32400
X395 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=408940 19040 1 0 $X=408750 $Y=16080
X396 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=417220 19040 1 0 $X=417030 $Y=16080
X397 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=426880 13600 0 0 $X=426690 $Y=13360
X398 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=427340 24480 1 0 $X=427150 $Y=21520
X399 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=437000 46240 1 0 $X=436810 $Y=43280
X400 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=450800 13600 0 0 $X=450610 $Y=13360
X401 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=458620 46240 1 0 $X=458430 $Y=43280
X402 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=459080 46240 0 0 $X=458890 $Y=46000
X403 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=464600 29920 1 0 $X=464410 $Y=26960
X404 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=465060 35360 1 0 $X=464870 $Y=32400
X405 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=478860 35360 0 0 $X=478670 $Y=35120
X406 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=497260 35360 1 0 $X=497070 $Y=32400
X407 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=512440 40800 1 0 $X=512250 $Y=37840
X408 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=513820 35360 1 0 $X=513630 $Y=32400
X409 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=515200 35360 0 0 $X=515010 $Y=35120
X410 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=519340 13600 1 0 $X=519150 $Y=10640
X411 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=520720 46240 1 0 $X=520530 $Y=43280
X412 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=549240 46240 0 0 $X=549050 $Y=46000
X413 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=567180 29920 0 0 $X=566990 $Y=29680
X414 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=575920 35360 1 0 $X=575730 $Y=32400
X415 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=591100 40800 0 0 $X=590910 $Y=40560
X416 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=591100 46240 0 0 $X=590910 $Y=46000
X417 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=603980 24480 1 0 $X=603790 $Y=21520
X418 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=604440 40800 0 0 $X=604250 $Y=40560
X419 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=619160 24480 0 0 $X=618970 $Y=24240
X420 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=630660 35360 0 0 $X=630470 $Y=35120
X421 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=632500 35360 1 0 $X=632310 $Y=32400
X422 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=634800 46240 0 0 $X=634610 $Y=46000
X423 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=642160 13600 1 0 $X=641970 $Y=10640
X424 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=647220 24480 0 0 $X=647030 $Y=24240
X425 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=649060 29920 1 0 $X=648870 $Y=26960
X426 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=660100 24480 1 0 $X=659910 $Y=21520
X427 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=671140 35360 1 0 $X=670950 $Y=32400
X428 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=673900 46240 0 0 $X=673710 $Y=46000
X429 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=675280 40800 0 0 $X=675090 $Y=40560
X430 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=681720 13600 1 0 $X=681530 $Y=10640
X431 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=682180 29920 1 0 $X=681990 $Y=26960
X432 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=682180 35360 1 0 $X=681990 $Y=32400
X433 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=697820 40800 1 0 $X=697630 $Y=37840
X434 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=702880 29920 0 0 $X=702690 $Y=29680
X435 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=713460 13600 1 0 $X=713270 $Y=10640
X436 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=731400 24480 0 0 $X=731210 $Y=24240
X437 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=738300 19040 1 0 $X=738110 $Y=16080
X438 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=738300 24480 1 0 $X=738110 $Y=21520
X439 1 2 1 2 sky130_fd_sc_hd__decap_8 $T=738760 29920 1 0 $X=738570 $Y=26960
X440 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 13600 1 0 $X=6710 $Y=10640
X441 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 29920 0 0 $X=6710 $Y=29680
X442 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 35360 0 0 $X=6710 $Y=35120
X443 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 40800 1 0 $X=6710 $Y=37840
X444 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=6900 40800 0 0 $X=6710 $Y=40560
X445 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=20240 35360 1 0 $X=20050 $Y=32400
X446 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=33120 19040 1 0 $X=32930 $Y=16080
X447 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=34040 24480 0 0 $X=33850 $Y=24240
X448 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=34960 24480 1 0 $X=34770 $Y=21520
X449 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=62100 40800 0 0 $X=61910 $Y=40560
X450 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=71300 19040 0 0 $X=71110 $Y=18800
X451 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=97980 40800 1 0 $X=97790 $Y=37840
X452 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=138920 13600 0 0 $X=138730 $Y=13360
X453 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=148580 13600 1 0 $X=148390 $Y=10640
X454 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=151340 13600 0 0 $X=151150 $Y=13360
X455 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=191360 13600 1 0 $X=191170 $Y=10640
X456 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=212060 19040 0 0 $X=211870 $Y=18800
X457 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=221720 29920 1 0 $X=221530 $Y=26960
X458 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=336260 24480 0 0 $X=336070 $Y=24240
X459 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=374900 40800 0 0 $X=374710 $Y=40560
X460 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=391460 29920 1 0 $X=391270 $Y=26960
X461 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=438840 46240 0 0 $X=438650 $Y=46000
X462 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=453100 46240 1 0 $X=452910 $Y=43280
X463 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=454940 35360 0 0 $X=454750 $Y=35120
X464 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=456780 40800 1 0 $X=456590 $Y=37840
X465 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=459080 29920 1 0 $X=458890 $Y=26960
X466 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=459540 35360 1 0 $X=459350 $Y=32400
X467 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=470120 24480 0 0 $X=469930 $Y=24240
X468 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=474720 13600 0 0 $X=474530 $Y=13360
X469 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=493580 13600 1 0 $X=493390 $Y=10640
X470 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=505080 13600 1 0 $X=504890 $Y=10640
X471 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=505080 29920 0 0 $X=504890 $Y=29680
X472 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=515200 24480 0 0 $X=515010 $Y=24240
X473 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=526700 13600 1 0 $X=526510 $Y=10640
X474 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=544640 40800 0 0 $X=544450 $Y=40560
X475 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=552920 24480 0 0 $X=552730 $Y=24240
X476 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=553380 29920 1 0 $X=553190 $Y=26960
X477 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=593400 35360 1 0 $X=593210 $Y=32400
X478 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=613640 24480 0 0 $X=613450 $Y=24240
X479 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=613640 35360 1 0 $X=613450 $Y=32400
X480 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=627440 24480 0 0 $X=627250 $Y=24240
X481 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=633420 13600 1 0 $X=633230 $Y=10640
X482 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=665620 35360 1 0 $X=665430 $Y=32400
X483 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=667000 13600 1 0 $X=666810 $Y=10640
X484 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=676200 13600 1 0 $X=676010 $Y=10640
X485 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=701040 40800 0 0 $X=700850 $Y=40560
X486 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=704720 13600 1 0 $X=704530 $Y=10640
X487 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=707480 24480 0 0 $X=707290 $Y=24240
X488 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=707480 35360 1 0 $X=707290 $Y=32400
X489 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=715300 29920 1 0 $X=715110 $Y=26960
X490 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=725880 24480 0 0 $X=725690 $Y=24240
X491 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=730020 35360 1 0 $X=729830 $Y=32400
X492 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=732780 19040 1 0 $X=732590 $Y=16080
X493 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=732780 24480 1 0 $X=732590 $Y=21520
X494 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 13600 0 0 $X=735350 $Y=13360
X495 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 19040 0 0 $X=735350 $Y=18800
X496 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=735540 24480 0 0 $X=735350 $Y=24240
X497 1 2 1 2 sky130_fd_sc_hd__decap_12 $T=736460 13600 1 0 $X=736270 $Y=10640
X498 1 2 293 291 2 13 1 sky130_fd_sc_hd__ebufn_2 $T=51060 19040 1 0 $X=50870 $Y=16080
X499 1 2 308 37 2 25 1 sky130_fd_sc_hd__ebufn_2 $T=69460 40800 0 0 $X=69270 $Y=40560
X500 1 2 334 336 2 30 1 sky130_fd_sc_hd__ebufn_2 $T=98440 24480 1 0 $X=98250 $Y=21520
X501 1 2 339 49 2 25 1 sky130_fd_sc_hd__ebufn_2 $T=99820 46240 1 0 $X=99630 $Y=43280
X502 1 2 361 362 2 27 1 sky130_fd_sc_hd__ebufn_2 $T=120060 29920 0 0 $X=119870 $Y=29680
X503 1 2 368 362 2 25 1 sky130_fd_sc_hd__ebufn_2 $T=126960 24480 1 0 $X=126770 $Y=21520
X504 1 2 372 362 2 14 1 sky130_fd_sc_hd__ebufn_2 $T=142600 35360 1 0 $X=142410 $Y=32400
X505 1 2 393 394 2 27 1 sky130_fd_sc_hd__ebufn_2 $T=149500 35360 1 0 $X=149310 $Y=32400
X506 1 2 406 65 2 13 1 sky130_fd_sc_hd__ebufn_2 $T=161460 40800 0 0 $X=161270 $Y=40560
X507 1 2 412 404 2 30 1 sky130_fd_sc_hd__ebufn_2 $T=174340 13600 0 0 $X=174150 $Y=13360
X508 1 2 445 442 2 14 1 sky130_fd_sc_hd__ebufn_2 $T=196420 29920 0 0 $X=196230 $Y=29680
X509 1 2 449 452 2 25 1 sky130_fd_sc_hd__ebufn_2 $T=201020 13600 1 0 $X=200830 $Y=10640
X510 1 2 461 452 2 13 1 sky130_fd_sc_hd__ebufn_2 $T=208380 13600 1 0 $X=208190 $Y=10640
X511 1 2 80 81 2 28 1 sky130_fd_sc_hd__ebufn_2 $T=214820 46240 0 0 $X=214630 $Y=46000
X512 1 2 466 468 2 27 1 sky130_fd_sc_hd__ebufn_2 $T=215280 13600 1 0 $X=215090 $Y=10640
X513 1 2 471 82 2 16 1 sky130_fd_sc_hd__ebufn_2 $T=218960 40800 1 0 $X=218770 $Y=37840
X514 1 2 467 82 2 27 1 sky130_fd_sc_hd__ebufn_2 $T=222180 35360 0 0 $X=221990 $Y=35120
X515 1 2 485 468 2 14 1 sky130_fd_sc_hd__ebufn_2 $T=230460 13600 0 0 $X=230270 $Y=13360
X516 1 2 482 473 2 30 1 sky130_fd_sc_hd__ebufn_2 $T=230460 29920 1 0 $X=230270 $Y=26960
X517 1 2 483 82 2 15 1 sky130_fd_sc_hd__ebufn_2 $T=230920 46240 1 0 $X=230730 $Y=43280
X518 1 2 490 473 2 13 1 sky130_fd_sc_hd__ebufn_2 $T=233220 35360 0 0 $X=233030 $Y=35120
X519 1 2 508 96 2 97 1 sky130_fd_sc_hd__ebufn_2 $T=246560 46240 1 0 $X=246370 $Y=43280
X520 1 2 514 103 2 104 1 sky130_fd_sc_hd__ebufn_2 $T=253920 46240 0 0 $X=253730 $Y=46000
X521 1 2 530 524 2 97 1 sky130_fd_sc_hd__ebufn_2 $T=268180 19040 1 0 $X=267990 $Y=16080
X522 1 2 538 524 2 107 1 sky130_fd_sc_hd__ebufn_2 $T=272320 13600 1 0 $X=272130 $Y=10640
X523 1 2 529 103 2 107 1 sky130_fd_sc_hd__ebufn_2 $T=278760 46240 0 0 $X=278570 $Y=46000
X524 1 2 549 543 2 94 1 sky130_fd_sc_hd__ebufn_2 $T=282900 19040 1 0 $X=282710 $Y=16080
X525 1 2 552 113 2 104 1 sky130_fd_sc_hd__ebufn_2 $T=286580 46240 0 0 $X=286390 $Y=46000
X526 1 2 564 563 2 104 1 sky130_fd_sc_hd__ebufn_2 $T=296240 29920 1 0 $X=296050 $Y=26960
X527 1 2 578 563 2 93 1 sky130_fd_sc_hd__ebufn_2 $T=309120 29920 0 0 $X=308930 $Y=29680
X528 1 2 579 563 2 94 1 sky130_fd_sc_hd__ebufn_2 $T=310040 24480 0 0 $X=309850 $Y=24240
X529 1 2 554 103 2 108 1 sky130_fd_sc_hd__ebufn_2 $T=322920 40800 0 0 $X=322730 $Y=40560
X530 1 2 597 589 2 104 1 sky130_fd_sc_hd__ebufn_2 $T=323840 35360 1 0 $X=323650 $Y=32400
X531 1 2 602 124 2 104 1 sky130_fd_sc_hd__ebufn_2 $T=328900 40800 0 0 $X=328710 $Y=40560
X532 1 2 608 589 2 94 1 sky130_fd_sc_hd__ebufn_2 $T=337180 35360 1 0 $X=336990 $Y=32400
X533 1 2 623 618 2 107 1 sky130_fd_sc_hd__ebufn_2 $T=350980 35360 1 0 $X=350790 $Y=32400
X534 1 2 635 618 2 97 1 sky130_fd_sc_hd__ebufn_2 $T=359260 40800 1 0 $X=359070 $Y=37840
X535 1 2 648 132 2 108 1 sky130_fd_sc_hd__ebufn_2 $T=370760 40800 0 0 $X=370570 $Y=40560
X536 1 2 669 652 2 106 1 sky130_fd_sc_hd__ebufn_2 $T=385020 24480 1 0 $X=384830 $Y=21520
X537 1 2 666 652 2 108 1 sky130_fd_sc_hd__ebufn_2 $T=392380 24480 0 0 $X=392190 $Y=24240
X538 1 2 676 670 2 94 1 sky130_fd_sc_hd__ebufn_2 $T=392840 40800 0 0 $X=392650 $Y=40560
X539 1 2 695 685 2 108 1 sky130_fd_sc_hd__ebufn_2 $T=408020 35360 0 0 $X=407830 $Y=35120
X540 1 2 733 732 2 106 1 sky130_fd_sc_hd__ebufn_2 $T=437000 24480 0 0 $X=436810 $Y=24240
X541 1 2 741 732 2 104 1 sky130_fd_sc_hd__ebufn_2 $T=450340 19040 1 0 $X=450150 $Y=16080
X542 1 2 744 723 2 94 1 sky130_fd_sc_hd__ebufn_2 $T=454940 29920 0 0 $X=454750 $Y=29680
X543 1 2 759 760 2 167 1 sky130_fd_sc_hd__ebufn_2 $T=477480 24480 0 0 $X=477290 $Y=24240
X544 1 2 794 795 2 178 1 sky130_fd_sc_hd__ebufn_2 $T=532680 24480 0 0 $X=532490 $Y=24240
X545 1 2 196 195 2 179 1 sky130_fd_sc_hd__ebufn_2 $T=534520 40800 0 0 $X=534330 $Y=40560
X546 1 2 798 795 2 179 1 sky130_fd_sc_hd__ebufn_2 $T=535440 35360 1 0 $X=535250 $Y=32400
X547 1 2 852 846 2 167 1 sky130_fd_sc_hd__ebufn_2 $T=609500 24480 0 0 $X=609310 $Y=24240
X548 1 2 857 215 2 167 1 sky130_fd_sc_hd__ebufn_2 $T=615940 40800 0 0 $X=615750 $Y=40560
X549 1 2 866 861 2 179 1 sky130_fd_sc_hd__ebufn_2 $T=628360 35360 1 0 $X=628170 $Y=32400
X550 1 2 864 215 2 179 1 sky130_fd_sc_hd__ebufn_2 $T=636180 40800 0 0 $X=635990 $Y=40560
X551 1 2 882 220 2 168 1 sky130_fd_sc_hd__ebufn_2 $T=651360 40800 0 0 $X=651170 $Y=40560
X552 1 2 225 226 2 179 1 sky130_fd_sc_hd__ebufn_2 $T=669760 46240 0 0 $X=669570 $Y=46000
X553 1 2 913 909 2 168 1 sky130_fd_sc_hd__ebufn_2 $T=693680 40800 1 0 $X=693490 $Y=37840
X554 1 2 937 928 2 168 1 sky130_fd_sc_hd__ebufn_2 $T=735540 29920 0 0 $X=735350 $Y=29680
X555 1 2 941 241 2 168 1 sky130_fd_sc_hd__ebufn_2 $T=737840 40800 0 0 $X=737650 $Y=40560
X630 1 2 258 261 13 ICV_6 $T=19780 40800 1 0 $X=19590 $Y=37840
X631 1 2 275 261 28 ICV_6 $T=33580 40800 0 0 $X=33390 $Y=40560
X632 1 2 22 23 25 ICV_6 $T=33580 46240 0 0 $X=33390 $Y=46000
X633 1 2 327 318 25 ICV_6 $T=89700 29920 0 0 $X=89510 $Y=29680
X634 1 2 328 318 14 ICV_6 $T=89700 35360 0 0 $X=89510 $Y=35120
X635 1 2 46 44 14 ICV_6 $T=89700 46240 0 0 $X=89510 $Y=46000
X636 1 2 341 336 28 ICV_6 $T=103960 19040 1 0 $X=103770 $Y=16080
X637 1 2 343 346 25 ICV_6 $T=103960 29920 1 0 $X=103770 $Y=26960
X638 1 2 429 438 28 ICV_6 $T=188140 19040 1 0 $X=187950 $Y=16080
X639 1 2 435 438 16 ICV_6 $T=188140 24480 1 0 $X=187950 $Y=21520
X640 1 2 432 438 15 ICV_6 $T=188140 29920 1 0 $X=187950 $Y=26960
X641 1 2 451 452 15 ICV_6 $T=201940 24480 0 0 $X=201750 $Y=24240
X642 1 2 448 442 25 ICV_6 $T=201940 35360 0 0 $X=201750 $Y=35120
X643 1 2 504 502 94 ICV_6 $T=244260 19040 1 0 $X=244070 $Y=16080
X644 1 2 515 502 107 ICV_6 $T=258060 13600 0 0 $X=257870 $Y=13360
X645 1 2 509 498 98 ICV_6 $T=258060 24480 0 0 $X=257870 $Y=24240
X646 1 2 522 96 106 ICV_6 $T=258060 46240 0 0 $X=257870 $Y=46000
X647 1 2 535 498 104 ICV_6 $T=272320 29920 1 0 $X=272130 $Y=26960
X648 1 2 520 500 108 ICV_6 $T=272320 40800 1 0 $X=272130 $Y=37840
X649 1 2 544 524 104 ICV_6 $T=286120 24480 0 0 $X=285930 $Y=24240
X650 1 2 568 543 106 ICV_6 $T=300380 19040 1 0 $X=300190 $Y=16080
X651 1 2 603 124 106 ICV_6 $T=328440 46240 1 0 $X=328250 $Y=43280
X652 1 2 630 631 94 ICV_6 $T=356500 19040 1 0 $X=356310 $Y=16080
X653 1 2 649 645 104 ICV_6 $T=370300 29920 0 0 $X=370110 $Y=29680
X654 1 2 668 652 98 ICV_6 $T=384560 19040 1 0 $X=384370 $Y=16080
X655 1 2 661 645 107 ICV_6 $T=384560 29920 1 0 $X=384370 $Y=26960
X656 1 2 682 670 93 ICV_6 $T=398360 40800 0 0 $X=398170 $Y=40560
X657 1 2 691 679 104 ICV_6 $T=412620 19040 1 0 $X=412430 $Y=16080
X658 1 2 698 145 104 ICV_6 $T=412620 40800 1 0 $X=412430 $Y=37840
X659 1 2 714 703 106 ICV_6 $T=426420 19040 0 0 $X=426230 $Y=18800
X660 1 2 737 732 108 ICV_6 $T=454480 13600 0 0 $X=454290 $Y=13360
X661 1 2 746 723 104 ICV_6 $T=454480 24480 0 0 $X=454290 $Y=24240
X662 1 2 739 725 108 ICV_6 $T=454480 40800 0 0 $X=454290 $Y=40560
X663 1 2 152 148 94 ICV_6 $T=454480 46240 0 0 $X=454290 $Y=46000
X664 1 2 784 782 178 ICV_6 $T=510600 24480 0 0 $X=510410 $Y=24240
X665 1 2 777 782 168 ICV_6 $T=510600 29920 0 0 $X=510410 $Y=29680
X666 1 2 781 782 174 ICV_6 $T=510600 35360 0 0 $X=510410 $Y=35120
X667 1 2 802 195 173 ICV_6 $T=538660 40800 0 0 $X=538470 $Y=40560
X668 1 2 824 820 178 ICV_6 $T=566720 24480 0 0 $X=566530 $Y=24240
X669 1 2 821 820 179 ICV_6 $T=566720 40800 0 0 $X=566530 $Y=40560
X670 1 2 832 834 167 ICV_6 $T=580980 24480 1 0 $X=580790 $Y=21520
X671 1 2 841 211 168 ICV_6 $T=594780 40800 0 0 $X=594590 $Y=40560
X672 1 2 853 846 177 ICV_6 $T=609040 29920 1 0 $X=608850 $Y=26960
X673 1 2 854 846 169 ICV_6 $T=609040 35360 1 0 $X=608850 $Y=32400
X674 1 2 863 861 177 ICV_6 $T=622840 24480 0 0 $X=622650 $Y=24240
X675 1 2 860 861 168 ICV_6 $T=622840 40800 0 0 $X=622650 $Y=40560
X676 1 2 895 886 173 ICV_6 $T=665160 40800 1 0 $X=664970 $Y=37840
X677 1 2 903 900 173 ICV_6 $T=678960 40800 0 0 $X=678770 $Y=40560
X678 1 2 227 226 177 ICV_6 $T=678960 46240 0 0 $X=678770 $Y=46000
X679 1 2 912 909 177 ICV_6 $T=693220 29920 1 0 $X=693030 $Y=26960
X680 1 2 935 928 174 ICV_6 $T=735080 35360 0 0 $X=734890 $Y=35120
X681 1 2 245 241 167 ICV_6 $T=735080 46240 0 0 $X=734890 $Y=46000
X754 1 2 ICV_10 $T=58880 35360 0 0 $X=58690 $Y=35120
X755 1 2 ICV_10 $T=86940 24480 0 0 $X=86750 $Y=24240
X756 1 2 ICV_10 $T=86940 40800 0 0 $X=86750 $Y=40560
X757 1 2 ICV_10 $T=157320 29920 1 0 $X=157130 $Y=26960
X758 1 2 ICV_10 $T=185380 40800 1 0 $X=185190 $Y=37840
X759 1 2 ICV_10 $T=269560 35360 1 0 $X=269370 $Y=32400
X760 1 2 ICV_10 $T=367540 46240 0 0 $X=367350 $Y=46000
X761 1 2 ICV_10 $T=416300 13600 1 0 $X=416110 $Y=10640
X762 1 2 ICV_10 $T=423660 35360 0 0 $X=423470 $Y=35120
X763 1 2 ICV_10 $T=444820 13600 1 0 $X=444630 $Y=10640
X764 1 2 ICV_10 $T=634340 29920 1 0 $X=634150 $Y=26960
X765 1 2 ICV_11 $T=6900 19040 1 0 $X=6710 $Y=16080
X766 1 2 ICV_11 $T=6900 19040 0 0 $X=6710 $Y=18800
X767 1 2 ICV_11 $T=6900 24480 1 0 $X=6710 $Y=21520
X768 1 2 ICV_11 $T=6900 24480 0 0 $X=6710 $Y=24240
X769 1 2 ICV_11 $T=6900 29920 1 0 $X=6710 $Y=26960
X770 1 2 ICV_11 $T=6900 35360 1 0 $X=6710 $Y=32400
X771 1 2 ICV_11 $T=6900 46240 1 0 $X=6710 $Y=43280
X772 1 2 ICV_11 $T=62100 13600 0 0 $X=61910 $Y=13360
X773 1 2 ICV_11 $T=105800 13600 0 0 $X=105610 $Y=13360
X774 1 2 ICV_11 $T=454480 19040 1 0 $X=454290 $Y=16080
X775 1 2 ICV_11 $T=459080 24480 0 0 $X=458890 $Y=24240
X776 1 2 ICV_11 $T=459080 29920 0 0 $X=458890 $Y=29680
X777 1 2 ICV_11 $T=459080 40800 0 0 $X=458890 $Y=40560
X778 1 2 ICV_11 $T=463680 13600 0 0 $X=463490 $Y=13360
X779 1 2 ICV_11 $T=479320 13600 1 0 $X=479130 $Y=10640
X780 1 2 ICV_11 $T=512440 24480 1 0 $X=512250 $Y=21520
X781 1 2 ICV_11 $T=525320 24480 1 0 $X=525130 $Y=21520
X782 1 2 ICV_11 $T=550620 13600 1 0 $X=550430 $Y=10640
X783 1 2 ICV_11 $T=567180 24480 1 0 $X=566990 $Y=21520
X784 1 2 ICV_11 $T=585580 24480 1 0 $X=585390 $Y=21520
X785 1 2 ICV_11 $T=649060 24480 1 0 $X=648870 $Y=21520
X786 1 2 ICV_11 $T=667920 24480 0 0 $X=667730 $Y=24240
X787 1 2 ICV_11 $T=721740 19040 1 0 $X=721550 $Y=16080
X788 1 2 ICV_11 $T=721740 24480 1 0 $X=721550 $Y=21520
X789 1 2 256 6 2 258 1 sky130_fd_sc_hd__dfxtp_1 $T=12420 40800 1 0 $X=12230 $Y=37840
X790 1 2 257 6 2 266 1 sky130_fd_sc_hd__dfxtp_1 $T=17940 19040 0 0 $X=17750 $Y=18800
X791 1 2 256 4 2 260 1 sky130_fd_sc_hd__dfxtp_1 $T=22080 40800 0 0 $X=21890 $Y=40560
X792 1 2 256 17 2 270 1 sky130_fd_sc_hd__dfxtp_1 $T=25760 35360 1 0 $X=25570 $Y=32400
X793 1 2 257 18 2 273 1 sky130_fd_sc_hd__dfxtp_1 $T=27600 24480 1 0 $X=27410 $Y=21520
X794 1 2 257 19 2 279 1 sky130_fd_sc_hd__dfxtp_1 $T=35880 29920 1 0 $X=35690 $Y=26960
X795 1 2 280 20 2 288 1 sky130_fd_sc_hd__dfxtp_1 $T=40480 24480 1 0 $X=40290 $Y=21520
X796 1 2 281 6 2 289 1 sky130_fd_sc_hd__dfxtp_1 $T=40480 35360 1 0 $X=40290 $Y=32400
X797 1 2 281 17 2 297 1 sky130_fd_sc_hd__dfxtp_1 $T=50600 35360 1 0 $X=50410 $Y=32400
X798 1 2 281 4 2 277 1 sky130_fd_sc_hd__dfxtp_1 $T=51060 29920 0 0 $X=50870 $Y=29680
X799 1 2 280 19 2 303 1 sky130_fd_sc_hd__dfxtp_1 $T=57040 24480 1 0 $X=56850 $Y=21520
X800 1 2 306 19 2 313 1 sky130_fd_sc_hd__dfxtp_1 $T=68540 29920 1 0 $X=68350 $Y=26960
X801 1 2 332 17 2 343 1 sky130_fd_sc_hd__dfxtp_1 $T=94300 29920 0 0 $X=94110 $Y=29680
X802 1 2 332 4 2 345 1 sky130_fd_sc_hd__dfxtp_1 $T=94300 35360 0 0 $X=94110 $Y=35120
X803 1 2 349 4 2 356 1 sky130_fd_sc_hd__dfxtp_1 $T=109480 19040 0 0 $X=109290 $Y=18800
X804 1 2 370 4 2 386 1 sky130_fd_sc_hd__dfxtp_1 $T=138460 19040 0 0 $X=138270 $Y=18800
X805 1 2 370 6 2 392 1 sky130_fd_sc_hd__dfxtp_1 $T=147660 19040 1 0 $X=147470 $Y=16080
X806 1 2 60 6 2 406 1 sky130_fd_sc_hd__dfxtp_1 $T=154560 46240 0 0 $X=154370 $Y=46000
X807 1 2 408 9 2 420 1 sky130_fd_sc_hd__dfxtp_1 $T=164680 35360 0 0 $X=164490 $Y=35120
X808 1 2 401 17 2 421 1 sky130_fd_sc_hd__dfxtp_1 $T=166060 19040 0 0 $X=165870 $Y=18800
X809 1 2 414 19 2 431 1 sky130_fd_sc_hd__dfxtp_1 $T=177560 24480 1 0 $X=177370 $Y=21520
X810 1 2 414 9 2 435 1 sky130_fd_sc_hd__dfxtp_1 $T=178020 24480 0 0 $X=177830 $Y=24240
X811 1 2 437 17 2 448 1 sky130_fd_sc_hd__dfxtp_1 $T=193200 35360 0 0 $X=193010 $Y=35120
X812 1 2 444 8 2 451 1 sky130_fd_sc_hd__dfxtp_1 $T=194580 24480 0 0 $X=194390 $Y=24240
X813 1 2 463 19 2 482 1 sky130_fd_sc_hd__dfxtp_1 $T=222640 29920 0 0 $X=222450 $Y=29680
X814 1 2 78 8 2 483 1 sky130_fd_sc_hd__dfxtp_1 $T=222640 46240 0 0 $X=222450 $Y=46000
X815 1 2 465 8 2 486 1 sky130_fd_sc_hd__dfxtp_1 $T=224020 24480 1 0 $X=223830 $Y=21520
X816 1 2 492 89 2 505 1 sky130_fd_sc_hd__dfxtp_1 $T=238280 19040 0 0 $X=238090 $Y=18800
X817 1 2 501 100 2 535 1 sky130_fd_sc_hd__dfxtp_1 $T=264960 29920 1 0 $X=264770 $Y=26960
X818 1 2 540 102 2 550 1 sky130_fd_sc_hd__dfxtp_1 $T=276460 35360 0 0 $X=276270 $Y=35120
X819 1 2 540 88 2 551 1 sky130_fd_sc_hd__dfxtp_1 $T=276920 29920 1 0 $X=276730 $Y=26960
X820 1 2 540 100 2 552 1 sky130_fd_sc_hd__dfxtp_1 $T=276920 29920 0 0 $X=276730 $Y=29680
X821 1 2 540 99 2 553 1 sky130_fd_sc_hd__dfxtp_1 $T=276920 40800 1 0 $X=276730 $Y=37840
X822 1 2 548 99 2 570 1 sky130_fd_sc_hd__dfxtp_1 $T=294860 13600 1 0 $X=294670 $Y=10640
X823 1 2 572 99 2 581 1 sky130_fd_sc_hd__dfxtp_1 $T=306360 13600 0 0 $X=306170 $Y=13360
X824 1 2 586 101 2 588 1 sky130_fd_sc_hd__dfxtp_1 $T=318320 29920 1 0 $X=318130 $Y=26960
X825 1 2 586 100 2 597 1 sky130_fd_sc_hd__dfxtp_1 $T=318320 29920 0 0 $X=318130 $Y=29680
X826 1 2 586 89 2 600 1 sky130_fd_sc_hd__dfxtp_1 $T=319240 35360 0 0 $X=319050 $Y=35120
X827 1 2 121 100 2 602 1 sky130_fd_sc_hd__dfxtp_1 $T=321080 46240 1 0 $X=320890 $Y=43280
X828 1 2 586 88 2 608 1 sky130_fd_sc_hd__dfxtp_1 $T=328900 24480 0 0 $X=328710 $Y=24240
X829 1 2 599 102 2 613 1 sky130_fd_sc_hd__dfxtp_1 $T=332580 19040 0 0 $X=332390 $Y=18800
X830 1 2 599 89 2 619 1 sky130_fd_sc_hd__dfxtp_1 $T=337640 24480 1 0 $X=337450 $Y=21520
X831 1 2 638 99 2 661 1 sky130_fd_sc_hd__dfxtp_1 $T=374900 29920 1 0 $X=374710 $Y=26960
X832 1 2 643 101 2 666 1 sky130_fd_sc_hd__dfxtp_1 $T=378120 13600 0 0 $X=377930 $Y=13360
X833 1 2 643 89 2 668 1 sky130_fd_sc_hd__dfxtp_1 $T=385940 19040 0 0 $X=385750 $Y=18800
X834 1 2 673 90 2 680 1 sky130_fd_sc_hd__dfxtp_1 $T=389160 13600 0 0 $X=388970 $Y=13360
X835 1 2 665 102 2 686 1 sky130_fd_sc_hd__dfxtp_1 $T=393760 46240 1 0 $X=393570 $Y=43280
X836 1 2 678 101 2 695 1 sky130_fd_sc_hd__dfxtp_1 $T=403880 35360 1 0 $X=403690 $Y=32400
X837 1 2 694 100 2 702 1 sky130_fd_sc_hd__dfxtp_1 $T=408940 13600 1 0 $X=408750 $Y=10640
X838 1 2 720 102 2 733 1 sky130_fd_sc_hd__dfxtp_1 $T=431020 19040 0 0 $X=430830 $Y=18800
X839 1 2 720 89 2 730 1 sky130_fd_sc_hd__dfxtp_1 $T=431020 24480 1 0 $X=430830 $Y=21520
X840 1 2 717 88 2 744 1 sky130_fd_sc_hd__dfxtp_1 $T=443900 29920 0 0 $X=443710 $Y=29680
X841 1 2 718 100 2 747 1 sky130_fd_sc_hd__dfxtp_1 $T=446200 35360 0 0 $X=446010 $Y=35120
X842 1 2 751 161 2 757 1 sky130_fd_sc_hd__dfxtp_1 $T=470120 40800 0 0 $X=469930 $Y=40560
X843 1 2 752 170 2 770 1 sky130_fd_sc_hd__dfxtp_1 $T=487140 29920 1 0 $X=486950 $Y=26960
X844 1 2 786 159 2 790 1 sky130_fd_sc_hd__dfxtp_1 $T=517500 35360 1 0 $X=517310 $Y=32400
X845 1 2 815 160 2 822 1 sky130_fd_sc_hd__dfxtp_1 $T=557980 29920 0 0 $X=557790 $Y=29680
X846 1 2 828 159 2 831 1 sky130_fd_sc_hd__dfxtp_1 $T=570860 35360 0 0 $X=570670 $Y=35120
X847 1 2 828 165 2 833 1 sky130_fd_sc_hd__dfxtp_1 $T=571780 29920 1 0 $X=571590 $Y=26960
X848 1 2 204 172 2 208 1 sky130_fd_sc_hd__dfxtp_1 $T=574540 46240 0 0 $X=574350 $Y=46000
X849 1 2 209 170 2 840 1 sky130_fd_sc_hd__dfxtp_1 $T=583740 40800 0 0 $X=583550 $Y=40560
X850 1 2 885 165 2 895 1 sky130_fd_sc_hd__dfxtp_1 $T=656420 40800 1 0 $X=656230 $Y=37840
X851 1 2 897 170 2 905 1 sky130_fd_sc_hd__dfxtp_1 $T=674820 35360 1 0 $X=674630 $Y=32400
X852 1 2 908 172 2 912 1 sky130_fd_sc_hd__dfxtp_1 $T=685860 29920 1 0 $X=685670 $Y=26960
X853 1 2 908 160 2 913 1 sky130_fd_sc_hd__dfxtp_1 $T=685860 35360 1 0 $X=685670 $Y=32400
X854 1 2 270 261 25 256 19 274 ICV_13 $T=27600 40800 1 0 $X=27410 $Y=37840
X855 1 2 298 278 28 281 9 302 ICV_13 $T=56580 40800 1 0 $X=56390 $Y=37840
X856 1 2 307 37 13 35 6 307 ICV_13 $T=61640 46240 1 0 $X=61450 $Y=43280
X857 1 2 314 316 16 306 9 314 ICV_13 $T=69000 29920 0 0 $X=68810 $Y=29680
X858 1 2 321 318 16 309 9 321 ICV_13 $T=75440 40800 0 0 $X=75250 $Y=40560
X859 1 2 324 318 15 309 8 324 ICV_13 $T=78200 35360 0 0 $X=78010 $Y=35120
X860 1 2 329 318 30 309 19 329 ICV_13 $T=84180 40800 1 0 $X=83990 $Y=37840
X861 1 2 335 336 13 325 6 335 ICV_13 $T=91540 13600 1 0 $X=91350 $Y=10640
X862 1 2 52 49 13 50 17 339 ICV_13 $T=103040 46240 0 0 $X=102850 $Y=46000
X863 1 2 353 346 30 332 8 350 ICV_13 $T=103500 40800 0 0 $X=103310 $Y=40560
X864 1 2 351 346 13 332 6 351 ICV_13 $T=104420 29920 0 0 $X=104230 $Y=29680
X865 1 2 369 359 27 349 18 369 ICV_13 $T=120060 13600 1 0 $X=119870 $Y=10640
X866 1 2 373 362 15 354 4 372 ICV_13 $T=124200 29920 0 0 $X=124010 $Y=29680
X867 1 2 374 362 13 354 6 374 ICV_13 $T=125580 35360 0 0 $X=125390 $Y=35120
X868 1 2 376 379 25 370 17 376 ICV_13 $T=127420 13600 0 0 $X=127230 $Y=13360
X869 1 2 396 394 16 383 9 396 ICV_13 $T=145820 29920 1 0 $X=145630 $Y=26960
X870 1 2 398 394 25 383 17 398 ICV_13 $T=146280 24480 0 0 $X=146090 $Y=24240
X871 1 2 400 394 28 383 8 402 ICV_13 $T=148120 40800 1 0 $X=147930 $Y=37840
X872 1 2 417 65 27 60 18 417 ICV_13 $T=163760 46240 1 0 $X=163570 $Y=43280
X873 1 2 426 423 15 408 8 426 ICV_13 $T=173880 40800 1 0 $X=173690 $Y=37840
X874 1 2 421 404 25 414 20 429 ICV_13 $T=176640 19040 1 0 $X=176450 $Y=16080
X875 1 2 425 423 14 408 17 428 ICV_13 $T=176640 29920 0 0 $X=176450 $Y=29680
X876 1 2 430 69 13 67 6 430 ICV_13 $T=176640 46240 1 0 $X=176450 $Y=43280
X877 1 2 436 438 13 414 6 436 ICV_13 $T=178480 13600 0 0 $X=178290 $Y=13360
X878 1 2 460 442 16 437 19 457 ICV_13 $T=199180 46240 1 0 $X=198990 $Y=43280
X879 1 2 458 442 15 437 8 458 ICV_13 $T=199640 35360 1 0 $X=199450 $Y=32400
X880 1 2 462 452 27 444 6 461 ICV_13 $T=202860 19040 1 0 $X=202670 $Y=16080
X881 1 2 476 468 28 465 18 466 ICV_13 $T=212520 13600 0 0 $X=212330 $Y=13360
X882 1 2 477 82 28 78 20 477 ICV_13 $T=216660 46240 1 0 $X=216470 $Y=43280
X883 1 2 478 82 13 78 6 478 ICV_13 $T=218500 40800 0 0 $X=218310 $Y=40560
X884 1 2 493 468 30 465 19 493 ICV_13 $T=231380 24480 1 0 $X=231190 $Y=21520
X885 1 2 488 82 14 78 17 495 ICV_13 $T=231840 40800 1 0 $X=231650 $Y=37840
X886 1 2 506 502 93 492 88 504 ICV_13 $T=238280 13600 0 0 $X=238090 $Y=13360
X887 1 2 510 500 98 496 89 510 ICV_13 $T=244720 35360 1 0 $X=244530 $Y=32400
X888 1 2 511 500 97 496 91 511 ICV_13 $T=244720 40800 1 0 $X=244530 $Y=37840
X889 1 2 512 502 97 492 91 512 ICV_13 $T=245640 19040 0 0 $X=245450 $Y=18800
X890 1 2 527 500 104 496 99 526 ICV_13 $T=258060 35360 1 0 $X=257870 $Y=32400
X891 1 2 526 500 107 496 100 527 ICV_13 $T=258520 35360 0 0 $X=258330 $Y=35120
X892 1 2 528 96 104 87 100 528 ICV_13 $T=258980 46240 1 0 $X=258790 $Y=43280
X893 1 2 531 524 98 518 89 531 ICV_13 $T=261740 19040 0 0 $X=261550 $Y=18800
X894 1 2 534 498 97 501 91 534 ICV_13 $T=264500 24480 0 0 $X=264310 $Y=24240
X895 1 2 537 498 106 501 102 537 ICV_13 $T=265420 29920 0 0 $X=265230 $Y=29680
X896 1 2 545 524 106 518 102 545 ICV_13 $T=273240 19040 0 0 $X=273050 $Y=18800
X897 1 2 551 113 94 105 101 554 ICV_13 $T=278300 46240 1 0 $X=278110 $Y=43280
X898 1 2 557 543 93 548 88 549 ICV_13 $T=287040 19040 1 0 $X=286850 $Y=16080
X899 1 2 559 113 97 540 91 559 ICV_13 $T=287040 40800 1 0 $X=286850 $Y=37840
X900 1 2 118 119 107 114 101 569 ICV_13 $T=294400 46240 0 0 $X=294210 $Y=46000
X901 1 2 569 119 108 114 88 576 ICV_13 $T=300840 40800 0 0 $X=300650 $Y=40560
X902 1 2 577 563 98 565 89 577 ICV_13 $T=301300 35360 0 0 $X=301110 $Y=35120
X903 1 2 575 563 107 565 90 578 ICV_13 $T=302220 35360 1 0 $X=302030 $Y=32400
X904 1 2 591 574 97 572 91 591 ICV_13 $T=314640 24480 0 0 $X=314450 $Y=24240
X905 1 2 594 574 93 572 101 592 ICV_13 $T=315100 19040 1 0 $X=314910 $Y=16080
X906 1 2 596 574 98 572 89 596 ICV_13 $T=316020 24480 1 0 $X=315830 $Y=21520
X907 1 2 605 595 93 599 90 605 ICV_13 $T=328440 13600 0 0 $X=328250 $Y=13360
X908 1 2 607 595 94 599 100 598 ICV_13 $T=328900 19040 1 0 $X=328710 $Y=16080
X909 1 2 610 589 97 586 99 609 ICV_13 $T=328900 29920 1 0 $X=328710 $Y=26960
X910 1 2 609 589 107 586 91 610 ICV_13 $T=328900 29920 0 0 $X=328710 $Y=29680
X911 1 2 606 589 106 586 90 604 ICV_13 $T=328900 40800 1 0 $X=328710 $Y=37840
X912 1 2 614 126 97 125 91 614 ICV_13 $T=333040 46240 1 0 $X=332850 $Y=43280
X913 1 2 627 618 98 615 89 627 ICV_13 $T=344080 40800 1 0 $X=343890 $Y=37840
X914 1 2 624 618 94 599 91 620 ICV_13 $T=345000 24480 1 0 $X=344810 $Y=21520
X915 1 2 632 631 104 621 100 632 ICV_13 $T=348220 13600 1 0 $X=348030 $Y=10640
X916 1 2 639 631 106 621 89 637 ICV_13 $T=356040 19040 0 0 $X=355850 $Y=18800
X917 1 2 641 132 106 130 99 131 ICV_13 $T=356040 46240 0 0 $X=355850 $Y=46000
X918 1 2 642 631 107 621 99 642 ICV_13 $T=357420 13600 0 0 $X=357230 $Y=13360
X919 1 2 647 631 108 621 101 647 ICV_13 $T=362480 13600 1 0 $X=362290 $Y=10640
X920 1 2 654 132 97 130 91 654 ICV_13 $T=368000 46240 1 0 $X=367810 $Y=43280
X921 1 2 656 645 98 638 89 656 ICV_13 $T=370760 35360 0 0 $X=370570 $Y=35120
X922 1 2 657 132 94 130 88 657 ICV_13 $T=370760 46240 0 0 $X=370570 $Y=46000
X923 1 2 658 645 97 638 91 658 ICV_13 $T=372140 40800 1 0 $X=371950 $Y=37840
X924 1 2 659 652 97 643 91 659 ICV_13 $T=372600 24480 1 0 $X=372410 $Y=21520
X925 1 2 660 645 94 638 88 660 ICV_13 $T=374440 24480 0 0 $X=374250 $Y=24240
X926 1 2 662 645 93 638 90 662 ICV_13 $T=374900 29920 0 0 $X=374710 $Y=29680
X927 1 2 675 670 97 665 91 675 ICV_13 $T=384560 35360 0 0 $X=384370 $Y=35120
X928 1 2 680 679 93 673 101 689 ICV_13 $T=397440 19040 1 0 $X=397250 $Y=16080
X929 1 2 690 679 98 673 89 690 ICV_13 $T=398360 24480 1 0 $X=398170 $Y=21520
X930 1 2 692 685 93 678 90 692 ICV_13 $T=398820 29920 0 0 $X=398630 $Y=29680
X931 1 2 706 685 97 678 100 704 ICV_13 $T=411700 29920 0 0 $X=411510 $Y=29680
X932 1 2 705 685 107 678 99 705 ICV_13 $T=412160 35360 0 0 $X=411970 $Y=35120
X933 1 2 707 685 98 678 89 707 ICV_13 $T=413080 35360 1 0 $X=412890 $Y=32400
X934 1 2 708 145 107 141 99 708 ICV_13 $T=414460 46240 0 0 $X=414270 $Y=46000
X935 1 2 709 145 106 141 102 709 ICV_13 $T=414920 40800 0 0 $X=414730 $Y=40560
X936 1 2 710 145 98 141 89 710 ICV_13 $T=414920 46240 1 0 $X=414730 $Y=43280
X937 1 2 715 703 107 694 99 715 ICV_13 $T=419520 13600 1 0 $X=419330 $Y=10640
X938 1 2 716 703 98 694 101 719 ICV_13 $T=420900 19040 1 0 $X=420710 $Y=16080
X939 1 2 722 725 106 718 102 722 ICV_13 $T=426880 35360 0 0 $X=426690 $Y=35120
X940 1 2 728 725 98 718 89 728 ICV_13 $T=428720 40800 0 0 $X=428530 $Y=40560
X941 1 2 729 723 106 717 102 729 ICV_13 $T=429180 29920 1 0 $X=428990 $Y=26960
X942 1 2 731 732 107 720 99 731 ICV_13 $T=430560 13600 0 0 $X=430370 $Y=13360
X943 1 2 738 732 97 720 91 738 ICV_13 $T=441140 19040 0 0 $X=440950 $Y=18800
X944 1 2 742 732 94 720 88 742 ICV_13 $T=443440 24480 1 0 $X=443250 $Y=21520
X945 1 2 748 732 93 720 90 748 ICV_13 $T=448040 13600 1 0 $X=447850 $Y=10640
X946 1 2 754 758 168 751 160 754 ICV_13 $T=469200 46240 1 0 $X=469010 $Y=43280
X947 1 2 765 758 178 751 170 765 ICV_13 $T=483920 46240 1 0 $X=483730 $Y=43280
X948 1 2 770 760 178 752 172 767 ICV_13 $T=484380 29920 0 0 $X=484190 $Y=29680
X949 1 2 768 760 179 752 171 768 ICV_13 $T=484380 35360 1 0 $X=484190 $Y=32400
X950 1 2 769 758 177 751 172 769 ICV_13 $T=484380 40800 1 0 $X=484190 $Y=37840
X951 1 2 775 185 178 180 170 775 ICV_13 $T=496800 40800 0 0 $X=496610 $Y=40560
X952 1 2 776 185 167 180 161 776 ICV_13 $T=497260 46240 1 0 $X=497070 $Y=43280
X953 1 2 793 195 167 192 160 792 ICV_13 $T=520720 40800 0 0 $X=520530 $Y=40560
X954 1 2 790 795 169 786 162 796 ICV_13 $T=523480 35360 0 0 $X=523290 $Y=35120
X955 1 2 797 795 177 786 172 797 ICV_13 $T=525320 29920 1 0 $X=525130 $Y=26960
X956 1 2 799 795 167 786 161 799 ICV_13 $T=527160 29920 0 0 $X=526970 $Y=29680
X957 1 2 804 803 167 801 161 804 ICV_13 $T=538200 24480 1 0 $X=538010 $Y=21520
X958 1 2 814 803 168 801 160 814 ICV_13 $T=546480 29920 0 0 $X=546290 $Y=29680
X959 1 2 816 203 169 199 159 816 ICV_13 $T=552920 46240 0 0 $X=552730 $Y=46000
X960 1 2 818 820 173 815 165 818 ICV_13 $T=556140 35360 1 0 $X=555950 $Y=32400
X961 1 2 825 820 177 815 172 825 ICV_13 $T=560280 29920 1 0 $X=560090 $Y=26960
X962 1 2 837 834 179 828 171 837 ICV_13 $T=580980 35360 0 0 $X=580790 $Y=35120
X963 1 2 839 834 177 828 170 836 ICV_13 $T=581440 24480 0 0 $X=581250 $Y=24240
X964 1 2 840 211 178 209 160 841 ICV_13 $T=583740 46240 1 0 $X=583550 $Y=43280
X965 1 2 845 846 173 843 170 844 ICV_13 $T=595240 24480 0 0 $X=595050 $Y=24240
X966 1 2 849 211 173 209 165 849 ICV_13 $T=595240 46240 1 0 $X=595050 $Y=43280
X967 1 2 850 211 167 209 161 850 ICV_13 $T=595240 46240 0 0 $X=595050 $Y=46000
X968 1 2 858 215 173 213 165 858 ICV_13 $T=609500 46240 1 0 $X=609310 $Y=43280
X969 1 2 869 861 174 856 171 866 ICV_13 $T=621920 40800 1 0 $X=621730 $Y=37840
X970 1 2 868 861 178 856 161 870 ICV_13 $T=623300 29920 0 0 $X=623110 $Y=29680
X971 1 2 871 215 177 213 172 871 ICV_13 $T=623300 46240 0 0 $X=623110 $Y=46000
X972 1 2 874 875 178 872 170 874 ICV_13 $T=635720 24480 0 0 $X=635530 $Y=24240
X973 1 2 876 875 173 872 165 876 ICV_13 $T=637100 29920 0 0 $X=636910 $Y=29680
X974 1 2 877 875 167 872 161 877 ICV_13 $T=637560 24480 1 0 $X=637370 $Y=21520
X975 1 2 878 875 177 872 172 878 ICV_13 $T=637560 29920 1 0 $X=637370 $Y=26960
X976 1 2 879 875 168 872 160 879 ICV_13 $T=637560 35360 1 0 $X=637370 $Y=32400
X977 1 2 881 220 178 217 160 882 ICV_13 $T=638480 46240 0 0 $X=638290 $Y=46000
X978 1 2 887 886 168 885 160 887 ICV_13 $T=651360 29920 0 0 $X=651170 $Y=29680
X979 1 2 888 886 169 885 159 888 ICV_13 $T=651360 35360 1 0 $X=651170 $Y=32400
X980 1 2 889 220 167 217 161 889 ICV_13 $T=651360 46240 0 0 $X=651170 $Y=46000
X981 1 2 893 886 179 885 171 893 ICV_13 $T=654120 35360 0 0 $X=653930 $Y=35120
X982 1 2 901 900 167 897 161 901 ICV_13 $T=666080 29920 0 0 $X=665890 $Y=29680
X983 1 2 902 900 169 897 159 902 ICV_13 $T=667460 35360 0 0 $X=667270 $Y=35120
X984 1 2 911 234 167 229 161 911 ICV_13 $T=685400 46240 0 0 $X=685210 $Y=46000
X985 1 2 915 909 178 908 170 915 ICV_13 $T=691380 29920 0 0 $X=691190 $Y=29680
X986 1 2 918 909 179 908 171 918 ICV_13 $T=695980 35360 1 0 $X=695790 $Y=32400
X987 1 2 919 234 174 229 159 922 ICV_13 $T=707480 46240 0 0 $X=707290 $Y=46000
X988 1 2 930 928 167 925 161 930 ICV_13 $T=714380 24480 0 0 $X=714190 $Y=24240
X989 1 2 931 928 169 925 159 931 ICV_13 $T=714380 35360 0 0 $X=714190 $Y=35120
X990 1 2 938 928 177 925 160 937 ICV_13 $T=727260 29920 1 0 $X=727070 $Y=26960
X991 1 2 939 241 177 238 160 941 ICV_13 $T=730940 46240 1 0 $X=730750 $Y=43280
X992 1 2 29 17 286 285 31 15 ICV_14 $T=38180 40800 0 0 $X=37990 $Y=40560
X993 1 2 306 18 323 323 316 27 ICV_14 $T=76820 19040 0 0 $X=76630 $Y=18800
X994 1 2 414 18 433 433 438 27 ICV_14 $T=177100 13600 1 0 $X=176910 $Y=10640
X995 1 2 465 6 480 480 468 13 ICV_14 $T=219880 13600 1 0 $X=219690 $Y=10640
X996 1 2 87 91 508 503 96 94 ICV_14 $T=238740 46240 0 0 $X=238550 $Y=46000
X997 1 2 548 89 560 560 543 98 ICV_14 $T=286580 24480 1 0 $X=286390 $Y=21520
X998 1 2 548 100 541 570 543 107 ICV_14 $T=293940 13600 0 0 $X=293750 $Y=13360
X999 1 2 643 90 664 664 652 93 ICV_14 $T=376740 13600 1 0 $X=376550 $Y=10640
X1000 1 2 718 99 724 724 725 107 ICV_14 $T=426420 40800 1 0 $X=426230 $Y=37840
X1001 1 2 752 161 759 756 760 168 ICV_14 $T=470120 29920 0 0 $X=469930 $Y=29680
X1002 1 2 751 171 766 766 758 179 ICV_14 $T=483000 46240 0 0 $X=482810 $Y=46000
X1003 1 2 801 159 810 810 803 169 ICV_14 $T=540040 40800 1 0 $X=539850 $Y=37840
X1004 1 2 204 165 835 835 206 173 ICV_14 $T=571320 40800 0 0 $X=571130 $Y=40560
X1005 1 2 856 170 868 870 861 167 ICV_14 $T=621920 29920 1 0 $X=621730 $Y=26960
X1006 1 2 217 170 881 883 875 179 ICV_14 $T=637560 46240 1 0 $X=637370 $Y=43280
X1007 1 2 217 172 892 892 220 177 ICV_14 $T=652280 46240 1 0 $X=652090 $Y=43280
X1008 1 2 297 278 25 281 18 305 305 278 27 ICV_15 $T=57960 35360 1 0 $X=57770 $Y=32400
X1009 1 2 367 359 13 349 20 364 364 359 28 ICV_15 $T=116380 19040 1 0 $X=116190 $Y=16080
X1010 1 2 399 394 14 383 4 399 387 394 13 ICV_15 $T=147200 29920 0 0 $X=147010 $Y=29680
X1011 1 2 418 423 27 401 8 413 413 404 15 ICV_15 $T=160540 29920 1 0 $X=160350 $Y=26960
X1012 1 2 428 423 25 408 4 425 415 423 13 ICV_15 $T=170660 35360 1 0 $X=170470 $Y=32400
X1013 1 2 434 438 14 414 4 434 431 438 30 ICV_15 $T=178020 19040 0 0 $X=177830 $Y=18800
X1014 1 2 481 468 25 465 4 485 486 468 15 ICV_15 $T=224020 19040 1 0 $X=223830 $Y=16080
X1015 1 2 495 82 25 496 90 507 507 500 93 ICV_15 $T=239200 40800 0 0 $X=239010 $Y=40560
X1016 1 2 517 502 108 492 101 517 521 502 106 ICV_15 $T=250700 19040 1 0 $X=250510 $Y=16080
X1017 1 2 651 652 94 643 88 651 653 652 107 ICV_15 $T=366620 19040 1 0 $X=366430 $Y=16080
X1018 1 2 693 670 108 665 99 687 687 670 107 ICV_15 $T=394220 40800 1 0 $X=394030 $Y=37840
X1019 1 2 696 685 106 673 91 688 689 679 108 ICV_15 $T=398820 24480 0 0 $X=398630 $Y=24240
X1020 1 2 747 725 104 718 101 739 735 725 97 ICV_15 $T=441140 40800 1 0 $X=440950 $Y=37840
X1021 1 2 743 723 93 717 90 743 734 723 97 ICV_15 $T=443440 29920 1 0 $X=443250 $Y=26960
X1022 1 2 745 723 108 717 101 745 721 723 107 ICV_15 $T=443900 35360 1 0 $X=443710 $Y=32400
X1023 1 2 809 803 179 801 171 809 807 803 174 ICV_15 $T=540960 35360 0 0 $X=540770 $Y=35120
X1024 1 2 823 820 174 815 159 819 819 820 169 ICV_15 $T=556600 40800 1 0 $X=556410 $Y=37840
X1025 1 2 830 834 168 828 160 830 833 834 173 ICV_15 $T=570860 29920 0 0 $X=570670 $Y=29680
X1026 1 2 906 900 174 897 162 906 907 900 168 ICV_15 $T=674820 40800 1 0 $X=674630 $Y=37840
X1027 1 2 926 234 178 229 165 923 923 234 173 ICV_15 $T=702880 46240 1 0 $X=702690 $Y=43280
X1028 1 2 246 241 174 925 171 936 936 928 179 ICV_15 $T=726340 40800 1 0 $X=726150 $Y=37840
X1029 1 2 256 8 259 259 261 15 ICV_16 $T=12420 35360 0 0 $X=12230 $Y=35120
X1030 1 2 29 8 285 284 31 28 ICV_16 $T=38180 46240 0 0 $X=37990 $Y=46000
X1031 1 2 280 8 301 303 291 30 ICV_16 $T=56580 29920 1 0 $X=56390 $Y=26960
X1032 1 2 35 17 308 38 37 14 ICV_16 $T=62100 46240 0 0 $X=61910 $Y=46000
X1033 1 2 306 4 315 313 316 30 ICV_16 $T=69460 24480 0 0 $X=69270 $Y=24240
X1034 1 2 325 20 341 337 336 27 ICV_16 $T=93840 13600 0 0 $X=93650 $Y=13360
X1035 1 2 54 8 391 391 58 15 ICV_16 $T=139840 46240 1 0 $X=139650 $Y=43280
X1036 1 2 408 19 427 427 423 30 ICV_16 $T=174340 40800 0 0 $X=174150 $Y=40560
X1037 1 2 437 20 443 443 442 28 ICV_16 $T=186300 40800 0 0 $X=186110 $Y=40560
X1038 1 2 444 19 454 454 452 30 ICV_16 $T=195040 29920 1 0 $X=194850 $Y=26960
X1039 1 2 463 18 470 470 473 27 ICV_16 $T=210220 35360 0 0 $X=210030 $Y=35120
X1040 1 2 463 17 472 472 473 25 ICV_16 $T=211140 24480 0 0 $X=210950 $Y=24240
X1041 1 2 540 89 558 558 113 98 ICV_16 $T=286580 35360 0 0 $X=286390 $Y=35120
X1042 1 2 125 101 129 625 126 94 ICV_16 $T=342700 40800 0 0 $X=342510 $Y=40560
X1043 1 2 621 90 629 629 631 93 ICV_16 $T=345460 13600 0 0 $X=345270 $Y=13360
X1044 1 2 718 88 736 736 725 94 ICV_16 $T=440220 40800 0 0 $X=440030 $Y=40560
X1045 1 2 718 90 740 740 725 93 ICV_16 $T=441140 46240 1 0 $X=440950 $Y=43280
X1046 1 2 752 159 755 753 758 169 ICV_16 $T=469200 35360 1 0 $X=469010 $Y=32400
X1047 1 2 180 160 785 787 185 173 ICV_16 $T=508760 46240 1 0 $X=508570 $Y=43280
X1048 1 2 786 170 794 789 795 173 ICV_16 $T=520720 24480 0 0 $X=520530 $Y=24240
X1049 1 2 801 162 807 805 803 173 ICV_16 $T=539580 35360 1 0 $X=539390 $Y=32400
X1050 1 2 828 162 838 838 834 174 ICV_16 $T=581440 35360 1 0 $X=581250 $Y=32400
X1051 1 2 885 162 894 894 886 174 ICV_16 $T=655500 40800 0 0 $X=655310 $Y=40560
X1052 1 2 908 159 917 917 909 169 ICV_16 $T=694600 35360 0 0 $X=694410 $Y=35120
X1053 1 2 908 162 921 922 234 169 ICV_16 $T=701500 40800 1 0 $X=701310 $Y=37840
X1054 1 2 257 8 264 ICV_20 $T=16100 29920 0 0 $X=15910 $Y=29680
X1055 1 2 29 20 284 ICV_20 $T=37720 46240 1 0 $X=37530 $Y=43280
X1056 1 2 29 4 295 ICV_20 $T=50140 46240 0 0 $X=49950 $Y=46000
X1057 1 2 306 17 312 ICV_20 $T=68080 24480 1 0 $X=67890 $Y=21520
X1058 1 2 306 8 322 ICV_20 $T=76360 29920 1 0 $X=76170 $Y=26960
X1059 1 2 309 17 327 ICV_20 $T=80500 29920 0 0 $X=80310 $Y=29680
X1060 1 2 309 6 330 ICV_20 $T=83720 46240 1 0 $X=83530 $Y=43280
X1061 1 2 325 19 334 ICV_20 $T=88780 24480 1 0 $X=88590 $Y=21520
X1062 1 2 325 4 338 ICV_20 $T=92920 19040 0 0 $X=92730 $Y=18800
X1063 1 2 332 9 352 ICV_20 $T=104420 35360 1 0 $X=104230 $Y=32400
X1064 1 2 349 17 355 ICV_20 $T=108560 19040 1 0 $X=108370 $Y=16080
X1065 1 2 349 9 357 ICV_20 $T=109940 24480 0 0 $X=109750 $Y=24240
X1066 1 2 54 6 380 ICV_20 $T=128340 46240 0 0 $X=128150 $Y=46000
X1067 1 2 401 4 403 ICV_20 $T=158240 19040 0 0 $X=158050 $Y=18800
X1068 1 2 437 18 441 ICV_20 $T=185380 35360 0 0 $X=185190 $Y=35120
X1069 1 2 444 4 450 ICV_20 $T=193660 19040 0 0 $X=193470 $Y=18800
X1070 1 2 87 88 503 ICV_20 $T=236440 46240 1 0 $X=236250 $Y=43280
X1071 1 2 518 90 532 ICV_20 $T=262660 13600 1 0 $X=262470 $Y=10640
X1072 1 2 518 100 544 ICV_20 $T=272780 19040 1 0 $X=272590 $Y=16080
X1073 1 2 586 102 606 ICV_20 $T=327980 35360 0 0 $X=327790 $Y=35120
X1074 1 2 643 102 669 ICV_20 $T=378120 19040 0 0 $X=377930 $Y=18800
X1075 1 2 665 90 682 ICV_20 $T=390540 46240 0 0 $X=390350 $Y=46000
X1076 1 2 141 101 697 ICV_20 $T=403420 46240 1 0 $X=403230 $Y=43280
X1077 1 2 694 90 713 ICV_20 $T=418600 13600 0 0 $X=418410 $Y=13360
X1078 1 2 694 89 716 ICV_20 $T=419520 24480 1 0 $X=419330 $Y=21520
X1079 1 2 717 91 734 ICV_20 $T=436080 29920 0 0 $X=435890 $Y=29680
X1080 1 2 718 91 735 ICV_20 $T=438380 35360 0 0 $X=438190 $Y=35120
X1081 1 2 717 100 746 ICV_20 $T=443900 24480 0 0 $X=443710 $Y=24240
X1082 1 2 751 165 763 ICV_20 $T=476560 40800 1 0 $X=476370 $Y=37840
X1083 1 2 772 171 779 ICV_20 $T=499560 40800 1 0 $X=499370 $Y=37840
X1084 1 2 772 172 780 ICV_20 $T=500020 24480 1 0 $X=499830 $Y=21520
X1085 1 2 801 172 806 ICV_20 $T=539580 29920 1 0 $X=539390 $Y=26960
X1086 1 2 199 172 811 ICV_20 $T=541420 46240 1 0 $X=541230 $Y=43280
X1087 1 2 828 161 832 ICV_20 $T=571320 24480 0 0 $X=571130 $Y=24240
X1088 1 2 843 165 845 ICV_20 $T=592940 29920 1 0 $X=592750 $Y=26960
X1089 1 2 843 172 853 ICV_20 $T=602600 29920 0 0 $X=602410 $Y=29680
X1090 1 2 843 159 854 ICV_20 $T=602600 35360 0 0 $X=602410 $Y=35120
X1091 1 2 213 161 857 ICV_20 $T=606740 46240 0 0 $X=606550 $Y=46000
X1092 1 2 213 160 865 ICV_20 $T=621000 46240 1 0 $X=620810 $Y=43280
X1093 1 2 885 161 891 ICV_20 $T=652740 29920 1 0 $X=652550 $Y=26960
X1094 1 2 897 165 903 ICV_20 $T=667460 40800 0 0 $X=667270 $Y=40560
X1095 1 2 925 162 935 ICV_20 $T=725880 35360 0 0 $X=725690 $Y=35120
X1096 1 2 ICV_23 $T=32200 24480 0 0 $X=32010 $Y=24240
X1097 1 2 ICV_23 $T=60260 13600 0 0 $X=60070 $Y=13360
X1098 1 2 ICV_23 $T=88320 13600 0 0 $X=88130 $Y=13360
X1099 1 2 ICV_23 $T=144440 13600 0 0 $X=144250 $Y=13360
X1100 1 2 ICV_23 $T=158700 35360 1 0 $X=158510 $Y=32400
X1101 1 2 ICV_23 $T=189520 13600 1 0 $X=189330 $Y=10640
X1102 1 2 ICV_23 $T=200560 29920 0 0 $X=200370 $Y=29680
X1103 1 2 ICV_23 $T=232300 13600 1 0 $X=232110 $Y=10640
X1104 1 2 ICV_23 $T=299000 24480 1 0 $X=298810 $Y=21520
X1105 1 2 ICV_23 $T=312800 19040 0 0 $X=312610 $Y=18800
X1106 1 2 ICV_23 $T=312800 35360 0 0 $X=312610 $Y=35120
X1107 1 2 ICV_23 $T=327060 29920 1 0 $X=326870 $Y=26960
X1108 1 2 ICV_23 $T=355120 35360 1 0 $X=354930 $Y=32400
X1109 1 2 ICV_23 $T=389160 13600 1 0 $X=388970 $Y=10640
X1110 1 2 ICV_23 $T=411240 35360 1 0 $X=411050 $Y=32400
X1111 1 2 ICV_23 $T=411240 46240 1 0 $X=411050 $Y=43280
X1112 1 2 ICV_23 $T=439300 35360 1 0 $X=439110 $Y=32400
X1113 1 2 ICV_23 $T=495420 46240 1 0 $X=495230 $Y=43280
X1114 1 2 ICV_23 $T=523480 24480 1 0 $X=523290 $Y=21520
X1115 1 2 ICV_23 $T=551540 35360 1 0 $X=551350 $Y=32400
X1116 1 2 ICV_23 $T=565340 29920 0 0 $X=565150 $Y=29680
X1117 1 2 ICV_23 $T=579600 35360 1 0 $X=579410 $Y=32400
X1118 1 2 ICV_23 $T=607660 24480 1 0 $X=607470 $Y=21520
X1119 1 2 ICV_23 $T=607660 40800 1 0 $X=607470 $Y=37840
X1120 1 2 ICV_23 $T=645840 13600 1 0 $X=645650 $Y=10640
X1121 1 2 ICV_23 $T=663780 24480 1 0 $X=663590 $Y=21520
X1122 1 2 ICV_23 $T=677580 29920 0 0 $X=677390 $Y=29680
X1123 1 2 ICV_23 $T=717140 13600 1 0 $X=716950 $Y=10640
X1124 1 2 ICV_24 $T=17940 19040 1 0 $X=17750 $Y=16080
X1125 1 2 ICV_24 $T=17940 35360 1 0 $X=17750 $Y=32400
X1126 1 2 ICV_24 $T=17940 46240 1 0 $X=17750 $Y=43280
X1127 1 2 ICV_24 $T=31740 29920 0 0 $X=31550 $Y=29680
X1128 1 2 ICV_24 $T=46000 40800 1 0 $X=45810 $Y=37840
X1129 1 2 ICV_24 $T=115920 29920 0 0 $X=115730 $Y=29680
X1130 1 2 ICV_24 $T=143980 40800 0 0 $X=143790 $Y=40560
X1131 1 2 ICV_24 $T=172040 35360 0 0 $X=171850 $Y=35120
X1132 1 2 ICV_24 $T=246100 13600 1 0 $X=245910 $Y=10640
X1133 1 2 ICV_24 $T=270480 46240 1 0 $X=270290 $Y=43280
X1134 1 2 ICV_24 $T=312340 40800 0 0 $X=312150 $Y=40560
X1135 1 2 ICV_24 $T=326600 19040 1 0 $X=326410 $Y=16080
X1136 1 2 ICV_24 $T=340400 46240 0 0 $X=340210 $Y=46000
X1137 1 2 ICV_24 $T=438840 40800 1 0 $X=438650 $Y=37840
X1138 1 2 ICV_24 $T=452640 19040 0 0 $X=452450 $Y=18800
X1139 1 2 ICV_24 $T=536820 24480 0 0 $X=536630 $Y=24240
X1140 1 2 ICV_24 $T=564880 35360 0 0 $X=564690 $Y=35120
X1141 1 2 ICV_24 $T=579140 29920 1 0 $X=578950 $Y=26960
X1142 1 2 ICV_24 $T=579140 40800 1 0 $X=578950 $Y=37840
X1143 1 2 ICV_24 $T=592940 24480 0 0 $X=592750 $Y=24240
X1144 1 2 ICV_24 $T=649060 35360 0 0 $X=648870 $Y=35120
X1145 1 2 ICV_24 $T=688160 13600 1 0 $X=687970 $Y=10640
X1146 1 2 11 2 267 1 sky130_fd_sc_hd__inv_1 $T=30360 29920 0 0 $X=30170 $Y=29680
X1147 1 2 21 2 261 1 sky130_fd_sc_hd__inv_1 $T=32200 40800 0 0 $X=32010 $Y=40560
X1148 1 2 33 2 291 1 sky130_fd_sc_hd__inv_1 $T=57960 24480 0 0 $X=57770 $Y=24240
X1149 1 2 32 2 278 1 sky130_fd_sc_hd__inv_1 $T=67160 35360 0 0 $X=66970 $Y=35120
X1150 1 2 36 2 316 1 sky130_fd_sc_hd__inv_1 $T=84180 29920 1 0 $X=83990 $Y=26960
X1151 1 2 39 2 318 1 sky130_fd_sc_hd__inv_1 $T=90620 35360 1 0 $X=90430 $Y=32400
X1152 1 2 45 2 336 1 sky130_fd_sc_hd__inv_1 $T=102580 24480 1 0 $X=102390 $Y=21520
X1153 1 2 47 2 346 1 sky130_fd_sc_hd__inv_1 $T=112700 46240 1 0 $X=112510 $Y=43280
X1154 1 2 51 2 359 1 sky130_fd_sc_hd__inv_1 $T=117300 24480 1 0 $X=117110 $Y=21520
X1155 1 2 53 2 362 1 sky130_fd_sc_hd__inv_1 $T=133860 40800 0 0 $X=133670 $Y=40560
X1156 1 2 56 2 379 1 sky130_fd_sc_hd__inv_1 $T=148580 24480 1 0 $X=148390 $Y=21520
X1157 1 2 59 2 394 1 sky130_fd_sc_hd__inv_1 $T=154560 35360 0 0 $X=154370 $Y=35120
X1158 1 2 61 2 404 1 sky130_fd_sc_hd__inv_1 $T=167900 24480 1 0 $X=167710 $Y=21520
X1159 1 2 62 2 65 1 sky130_fd_sc_hd__inv_1 $T=171580 46240 0 0 $X=171390 $Y=46000
X1160 1 2 64 2 423 1 sky130_fd_sc_hd__inv_1 $T=184920 29920 1 0 $X=184730 $Y=26960
X1161 1 2 66 2 438 1 sky130_fd_sc_hd__inv_1 $T=186760 24480 1 0 $X=186570 $Y=21520
X1162 1 2 72 2 442 1 sky130_fd_sc_hd__inv_1 $T=200560 40800 0 0 $X=200370 $Y=40560
X1163 1 2 75 2 69 1 sky130_fd_sc_hd__inv_1 $T=200560 46240 0 0 $X=200370 $Y=46000
X1164 1 2 71 2 452 1 sky130_fd_sc_hd__inv_1 $T=214360 24480 1 0 $X=214170 $Y=21520
X1165 1 2 79 2 468 1 sky130_fd_sc_hd__inv_1 $T=223100 24480 0 0 $X=222910 $Y=24240
X1166 1 2 77 2 473 1 sky130_fd_sc_hd__inv_1 $T=234600 29920 1 0 $X=234410 $Y=26960
X1167 1 2 76 2 82 1 sky130_fd_sc_hd__inv_1 $T=235060 46240 1 0 $X=234870 $Y=43280
X1168 1 2 33 2 502 1 sky130_fd_sc_hd__inv_1 $T=242880 24480 1 0 $X=242690 $Y=21520
X1169 1 2 11 2 498 1 sky130_fd_sc_hd__inv_1 $T=242880 29920 1 0 $X=242690 $Y=26960
X1170 1 2 21 2 500 1 sky130_fd_sc_hd__inv_1 $T=259440 40800 0 0 $X=259250 $Y=40560
X1171 1 2 39 2 524 1 sky130_fd_sc_hd__inv_1 $T=263120 24480 0 0 $X=262930 $Y=24240
X1172 1 2 32 2 113 1 sky130_fd_sc_hd__inv_1 $T=291640 35360 1 0 $X=291450 $Y=32400
X1173 1 2 45 2 543 1 sky130_fd_sc_hd__inv_1 $T=296240 24480 0 0 $X=296050 $Y=24240
X1174 1 2 36 2 563 1 sky130_fd_sc_hd__inv_1 $T=314180 35360 1 0 $X=313990 $Y=32400
X1175 1 2 47 2 124 1 sky130_fd_sc_hd__inv_1 $T=319700 46240 1 0 $X=319510 $Y=43280
X1176 1 2 56 2 574 1 sky130_fd_sc_hd__inv_1 $T=325680 29920 1 0 $X=325490 $Y=26960
X1177 1 2 53 2 589 1 sky130_fd_sc_hd__inv_1 $T=326600 35360 0 0 $X=326410 $Y=35120
X1178 1 2 51 2 595 1 sky130_fd_sc_hd__inv_1 $T=336260 24480 1 0 $X=336070 $Y=21520
X1179 1 2 62 2 618 1 sky130_fd_sc_hd__inv_1 $T=350060 35360 0 0 $X=349870 $Y=35120
X1180 1 2 61 2 631 1 sky130_fd_sc_hd__inv_1 $T=353280 19040 0 0 $X=353090 $Y=18800
X1181 1 2 59 2 645 1 sky130_fd_sc_hd__inv_1 $T=368460 35360 1 0 $X=368270 $Y=32400
X1182 1 2 66 2 652 1 sky130_fd_sc_hd__inv_1 $T=373060 24480 0 0 $X=372870 $Y=24240
X1183 1 2 75 2 670 1 sky130_fd_sc_hd__inv_1 $T=392380 46240 1 0 $X=392190 $Y=43280
X1184 1 2 72 2 679 1 sky130_fd_sc_hd__inv_1 $T=396520 24480 0 0 $X=396330 $Y=24240
X1185 1 2 77 2 685 1 sky130_fd_sc_hd__inv_1 $T=402500 35360 1 0 $X=402310 $Y=32400
X1186 1 2 139 2 145 1 sky130_fd_sc_hd__inv_1 $T=411240 46240 0 0 $X=411050 $Y=46000
X1187 1 2 71 2 703 1 sky130_fd_sc_hd__inv_1 $T=416300 19040 0 0 $X=416110 $Y=18800
X1188 1 2 79 2 723 1 sky130_fd_sc_hd__inv_1 $T=433320 24480 0 0 $X=433130 $Y=24240
X1189 1 2 76 2 725 1 sky130_fd_sc_hd__inv_1 $T=435620 46240 1 0 $X=435430 $Y=43280
X1190 1 2 64 2 732 1 sky130_fd_sc_hd__inv_1 $T=438380 24480 1 0 $X=438190 $Y=21520
X1191 1 2 156 2 760 1 sky130_fd_sc_hd__inv_1 $T=491280 35360 0 0 $X=491090 $Y=35120
X1192 1 2 155 2 758 1 sky130_fd_sc_hd__inv_1 $T=492200 40800 0 0 $X=492010 $Y=40560
X1193 1 2 181 2 782 1 sky130_fd_sc_hd__inv_1 $T=509220 35360 0 0 $X=509030 $Y=35120
X1194 1 2 186 2 185 1 sky130_fd_sc_hd__inv_1 $T=509220 46240 0 0 $X=509030 $Y=46000
X1195 1 2 191 2 795 1 sky130_fd_sc_hd__inv_1 $T=537280 35360 0 0 $X=537090 $Y=35120
X1196 1 2 197 2 803 1 sky130_fd_sc_hd__inv_1 $T=543260 40800 0 0 $X=543070 $Y=40560
X1197 1 2 202 2 820 1 sky130_fd_sc_hd__inv_1 $T=567180 35360 0 0 $X=566990 $Y=35120
X1198 1 2 205 2 834 1 sky130_fd_sc_hd__inv_1 $T=589720 40800 1 0 $X=589530 $Y=37840
X1199 1 2 212 2 846 1 sky130_fd_sc_hd__inv_1 $T=610420 35360 0 0 $X=610230 $Y=35120
X1200 1 2 214 2 861 1 sky130_fd_sc_hd__inv_1 $T=633420 40800 1 0 $X=633230 $Y=37840
X1201 1 2 216 2 875 1 sky130_fd_sc_hd__inv_1 $T=644920 40800 1 0 $X=644730 $Y=37840
X1202 1 2 221 2 886 1 sky130_fd_sc_hd__inv_1 $T=655040 40800 1 0 $X=654850 $Y=37840
X1203 1 2 223 2 900 1 sky130_fd_sc_hd__inv_1 $T=672060 46240 1 0 $X=671870 $Y=43280
X1204 1 2 231 2 909 1 sky130_fd_sc_hd__inv_1 $T=686780 35360 0 0 $X=686590 $Y=35120
X1205 1 2 237 2 928 1 sky130_fd_sc_hd__inv_1 $T=719900 40800 1 0 $X=719710 $Y=37840
X1206 1 2 277 278 14 ICV_26 $T=35880 35360 1 0 $X=35690 $Y=32400
X1207 1 2 283 278 30 ICV_26 $T=43240 29920 1 0 $X=43050 $Y=26960
X1208 1 2 330 318 13 ICV_26 $T=90160 40800 0 0 $X=89970 $Y=40560
X1209 1 2 352 346 16 ICV_26 $T=110400 35360 0 0 $X=110210 $Y=35120
X1210 1 2 357 359 16 ICV_26 $T=118680 29920 1 0 $X=118490 $Y=26960
X1211 1 2 375 362 30 ICV_26 $T=132480 40800 1 0 $X=132290 $Y=37840
X1212 1 2 388 394 30 ICV_26 $T=146280 40800 0 0 $X=146090 $Y=40560
X1213 1 2 389 58 30 ICV_26 $T=146280 46240 0 0 $X=146090 $Y=46000
X1214 1 2 416 65 25 ICV_26 $T=169280 40800 0 0 $X=169090 $Y=40560
X1215 1 2 447 69 16 ICV_26 $T=195960 46240 0 0 $X=195770 $Y=46000
X1216 1 2 459 452 16 ICV_26 $T=206540 24480 0 0 $X=206350 $Y=24240
X1217 1 2 475 473 28 ICV_26 $T=218040 29920 0 0 $X=217850 $Y=29680
X1218 1 2 487 473 15 ICV_26 $T=230460 29920 0 0 $X=230270 $Y=29680
X1219 1 2 525 500 106 ICV_26 $T=264960 40800 1 0 $X=264770 $Y=37840
X1220 1 2 584 563 97 ICV_26 $T=314640 35360 0 0 $X=314450 $Y=35120
X1221 1 2 757 758 167 ICV_26 $T=477480 40800 0 0 $X=477290 $Y=40560
X1222 1 2 764 760 173 ICV_26 $T=485760 24480 0 0 $X=485570 $Y=24240
X1223 1 2 767 760 177 ICV_26 $T=490360 24480 0 0 $X=490170 $Y=24240
X1224 1 2 184 185 177 ICV_26 $T=503700 46240 0 0 $X=503510 $Y=46000
X1225 1 2 773 782 167 ICV_26 $T=507840 24480 1 0 $X=507650 $Y=21520
X1226 1 2 783 782 169 ICV_26 $T=509220 35360 1 0 $X=509030 $Y=32400
X1227 1 2 806 803 177 ICV_26 $T=547400 29920 1 0 $X=547210 $Y=26960
X1228 1 2 808 803 178 ICV_26 $T=548320 24480 0 0 $X=548130 $Y=24240
X1229 1 2 817 820 167 ICV_26 $T=562580 24480 1 0 $X=562390 $Y=21520
X1230 1 2 844 846 178 ICV_26 $T=599380 24480 1 0 $X=599190 $Y=21520
X1231 1 2 890 886 178 ICV_26 $T=660560 29920 1 0 $X=660370 $Y=26960
X1232 1 2 233 234 179 ICV_26 $T=688620 46240 1 0 $X=688430 $Y=43280
X1233 1 2 932 241 178 ICV_26 $T=721740 40800 1 0 $X=721550 $Y=37840
X1234 1 2 256 18 272 ICV_28 $T=24380 35360 0 0 $X=24190 $Y=35120
X1235 1 2 280 9 290 ICV_28 $T=39560 24480 0 0 $X=39370 $Y=24240
X1236 1 2 325 8 342 ICV_28 $T=92460 29920 1 0 $X=92270 $Y=26960
X1237 1 2 354 18 361 ICV_28 $T=112240 35360 1 0 $X=112050 $Y=32400
X1238 1 2 67 17 68 ICV_28 $T=174340 46240 0 0 $X=174150 $Y=46000
X1239 1 2 501 99 523 ICV_28 $T=252080 29920 1 0 $X=251890 $Y=26960
X1240 1 2 540 90 555 ICV_28 $T=284280 29920 1 0 $X=284090 $Y=26960
X1241 1 2 621 91 636 ICV_28 $T=355580 24480 0 0 $X=355390 $Y=24240
X1242 1 2 673 102 681 ICV_28 $T=389160 24480 1 0 $X=388970 $Y=21520
X1243 1 2 146 89 726 ICV_28 $T=426420 46240 1 0 $X=426230 $Y=43280
X1244 1 2 717 89 727 ICV_28 $T=426880 29920 0 0 $X=426690 $Y=29680
X1245 1 2 772 160 777 ICV_28 $T=495880 29920 0 0 $X=495690 $Y=29680
X1246 1 2 772 165 778 ICV_28 $T=497260 29920 1 0 $X=497070 $Y=26960
X1247 1 2 772 162 781 ICV_28 $T=499100 35360 0 0 $X=498910 $Y=35120
X1248 1 2 801 170 808 ICV_28 $T=539120 24480 0 0 $X=538930 $Y=24240
X1249 1 2 815 161 817 ICV_28 $T=553380 24480 1 0 $X=553190 $Y=21520
X1250 1 2 209 172 210 ICV_28 $T=581900 46240 0 0 $X=581710 $Y=46000
X1251 1 2 238 172 939 ICV_28 $T=725880 40800 0 0 $X=725690 $Y=40560
X1252 1 2 256 9 262 ICV_29 $T=12420 40800 0 0 $X=12230 $Y=40560
X1253 1 2 256 20 275 ICV_29 $T=25300 46240 1 0 $X=25110 $Y=43280
X1254 1 2 29 6 296 ICV_29 $T=48300 46240 1 0 $X=48110 $Y=43280
X1255 1 2 309 18 317 ICV_29 $T=68540 35360 0 0 $X=68350 $Y=35120
X1256 1 2 332 18 344 ICV_29 $T=92000 35360 1 0 $X=91810 $Y=32400
X1257 1 2 354 20 363 ICV_29 $T=111780 40800 1 0 $X=111590 $Y=37840
X1258 1 2 54 19 389 ICV_29 $T=136160 46240 0 0 $X=135970 $Y=46000
X1259 1 2 370 18 390 ICV_29 $T=138000 19040 1 0 $X=137810 $Y=16080
X1260 1 2 60 17 416 ICV_29 $T=161920 46240 0 0 $X=161730 $Y=46000
X1261 1 2 105 88 111 ICV_29 $T=262660 46240 0 0 $X=262470 $Y=46000
X1262 1 2 518 99 538 ICV_29 $T=270940 13600 0 0 $X=270750 $Y=13360
X1263 1 2 105 100 514 ICV_29 $T=275540 40800 0 0 $X=275350 $Y=40560
X1264 1 2 114 100 566 ICV_29 $T=289800 46240 1 0 $X=289610 $Y=43280
X1265 1 2 565 91 584 ICV_29 $T=308200 40800 1 0 $X=308010 $Y=37840
X1266 1 2 678 88 684 ICV_29 $T=392380 35360 1 0 $X=392190 $Y=32400
X1267 1 2 694 88 700 ICV_29 $T=406180 13600 0 0 $X=405990 $Y=13360
X1268 1 2 717 99 721 ICV_29 $T=424580 35360 1 0 $X=424390 $Y=32400
X1269 1 2 752 165 764 ICV_29 $T=477480 29920 1 0 $X=477290 $Y=26960
X1270 1 2 856 159 862 ICV_29 $T=611800 35360 0 0 $X=611610 $Y=35120
X1271 1 2 229 162 919 ICV_29 $T=696900 46240 0 0 $X=696710 $Y=46000
X1272 1 2 265 267 16 264 267 15 ICV_30 $T=23920 24480 0 0 $X=23730 $Y=24240
X1273 1 2 266 267 13 269 267 14 ICV_30 $T=24840 19040 1 0 $X=24650 $Y=16080
X1274 1 2 272 261 27 274 261 30 ICV_30 $T=34040 35360 0 0 $X=33850 $Y=35120
X1275 1 2 273 267 27 271 267 25 ICV_30 $T=34500 19040 0 0 $X=34310 $Y=18800
X1276 1 2 276 267 28 279 267 30 ICV_30 $T=34500 29920 0 0 $X=34310 $Y=29680
X1277 1 2 290 291 16 289 278 13 ICV_30 $T=48300 29920 1 0 $X=48110 $Y=26960
X1278 1 2 286 31 25 292 278 15 ICV_30 $T=48300 40800 1 0 $X=48110 $Y=37840
X1279 1 2 288 291 28 287 291 25 ICV_30 $T=48760 24480 1 0 $X=48570 $Y=21520
X1280 1 2 295 31 14 296 31 13 ICV_30 $T=52440 40800 0 0 $X=52250 $Y=40560
X1281 1 2 299 291 27 300 291 14 ICV_30 $T=63020 19040 0 0 $X=62830 $Y=18800
X1282 1 2 311 316 28 320 316 13 ICV_30 $T=76360 13600 0 0 $X=76170 $Y=13360
X1283 1 2 40 37 15 41 42 14 ICV_30 $T=76360 46240 0 0 $X=76170 $Y=46000
X1284 1 2 315 316 14 312 316 25 ICV_30 $T=77740 24480 1 0 $X=77550 $Y=21520
X1285 1 2 338 336 14 331 336 25 ICV_30 $T=101200 19040 0 0 $X=101010 $Y=18800
X1286 1 2 340 336 16 342 336 15 ICV_30 $T=101660 24480 0 0 $X=101470 $Y=24240
X1287 1 2 344 346 27 345 346 14 ICV_30 $T=102120 35360 0 0 $X=101930 $Y=35120
X1288 1 2 347 346 28 350 346 15 ICV_30 $T=104420 46240 1 0 $X=104230 $Y=43280
X1289 1 2 356 359 14 355 359 25 ICV_30 $T=118220 19040 0 0 $X=118030 $Y=18800
X1290 1 2 360 359 30 365 359 15 ICV_30 $T=118680 24480 1 0 $X=118490 $Y=21520
X1291 1 2 366 362 16 363 362 28 ICV_30 $T=122820 40800 1 0 $X=122630 $Y=37840
X1292 1 2 381 58 16 380 58 13 ICV_30 $T=135700 40800 0 0 $X=135510 $Y=40560
X1293 1 2 384 379 15 385 379 30 ICV_30 $T=140300 24480 1 0 $X=140110 $Y=21520
X1294 1 2 390 379 27 386 379 14 ICV_30 $T=147200 19040 0 0 $X=147010 $Y=18800
X1295 1 2 409 404 27 407 404 13 ICV_30 $T=166060 13600 1 0 $X=165870 $Y=10640
X1296 1 2 420 423 16 419 423 28 ICV_30 $T=174340 35360 0 0 $X=174150 $Y=35120
X1297 1 2 441 442 27 446 442 13 ICV_30 $T=192740 40800 1 0 $X=192550 $Y=37840
X1298 1 2 453 452 28 450 452 14 ICV_30 $T=203780 19040 0 0 $X=203590 $Y=18800
X1299 1 2 519 498 108 533 524 108 ICV_30 $T=272780 35360 1 0 $X=272590 $Y=32400
X1300 1 2 532 524 93 542 524 94 ICV_30 $T=276000 24480 0 0 $X=275810 $Y=24240
X1301 1 2 550 113 106 553 113 107 ICV_30 $T=283360 35360 1 0 $X=283170 $Y=32400
X1302 1 2 567 119 98 576 119 94 ICV_30 $T=303140 46240 1 0 $X=302950 $Y=43280
X1303 1 2 120 119 93 566 119 104 ICV_30 $T=305900 46240 0 0 $X=305710 $Y=46000
X1304 1 2 573 574 104 580 574 94 ICV_30 $T=306820 19040 1 0 $X=306630 $Y=16080
X1305 1 2 582 124 108 587 124 94 ICV_30 $T=314640 40800 0 0 $X=314450 $Y=40560
X1306 1 2 585 563 106 588 589 108 ICV_30 $T=315560 35360 1 0 $X=315370 $Y=32400
X1307 1 2 583 574 106 592 574 108 ICV_30 $T=317400 19040 0 0 $X=317210 $Y=18800
X1308 1 2 600 589 98 604 589 93 ICV_30 $T=328900 35360 1 0 $X=328710 $Y=32400
X1309 1 2 613 595 106 619 595 98 ICV_30 $T=342700 19040 0 0 $X=342510 $Y=18800
X1310 1 2 617 618 108 622 618 106 ICV_30 $T=342700 35360 1 0 $X=342510 $Y=32400
X1311 1 2 650 645 106 655 652 104 ICV_30 $T=371220 35360 1 0 $X=371030 $Y=32400
X1312 1 2 667 670 104 674 670 98 ICV_30 $T=384560 40800 0 0 $X=384370 $Y=40560
X1313 1 2 681 679 106 688 679 97 ICV_30 $T=399280 19040 0 0 $X=399090 $Y=18800
X1314 1 2 701 703 97 700 703 94 ICV_30 $T=414920 24480 0 0 $X=414730 $Y=24240
X1315 1 2 704 685 104 697 145 108 ICV_30 $T=418140 40800 1 0 $X=417950 $Y=37840
X1316 1 2 713 703 93 730 732 98 ICV_30 $T=432400 19040 1 0 $X=432210 $Y=16080
X1317 1 2 702 703 104 719 703 108 ICV_30 $T=433780 13600 1 0 $X=433590 $Y=10640
X1318 1 2 755 760 169 761 760 174 ICV_30 $T=483000 35360 0 0 $X=482810 $Y=35120
X1319 1 2 763 758 173 762 758 174 ICV_30 $T=483920 40800 0 0 $X=483730 $Y=40560
X1320 1 2 778 782 173 780 782 177 ICV_30 $T=507840 29920 1 0 $X=507650 $Y=26960
X1321 1 2 774 185 174 785 185 168 ICV_30 $T=511060 46240 0 0 $X=510870 $Y=46000
X1322 1 2 791 795 168 796 795 174 ICV_30 $T=527160 35360 1 0 $X=526970 $Y=32400
X1323 1 2 811 203 177 812 203 174 ICV_30 $T=553380 46240 1 0 $X=553190 $Y=43280
X1324 1 2 822 820 168 826 206 167 ICV_30 $T=567640 35360 1 0 $X=567450 $Y=32400
X1325 1 2 831 834 169 829 206 179 ICV_30 $T=581440 40800 1 0 $X=581250 $Y=37840
X1326 1 2 848 846 168 851 846 179 ICV_30 $T=600760 35360 1 0 $X=600570 $Y=32400
X1327 1 2 859 861 173 862 861 169 ICV_30 $T=620080 35360 1 0 $X=619890 $Y=32400
X1328 1 2 873 875 169 880 875 174 ICV_30 $T=642160 40800 0 0 $X=641970 $Y=40560
X1329 1 2 896 886 177 891 886 167 ICV_30 $T=665620 29920 1 0 $X=665430 $Y=26960
X1330 1 2 905 900 178 904 900 177 ICV_30 $T=681720 29920 0 0 $X=681530 $Y=29680
X1331 1 2 914 234 168 916 234 177 ICV_30 $T=693680 46240 1 0 $X=693490 $Y=43280
X1332 1 2 920 909 173 924 909 167 ICV_30 $T=707480 29920 0 0 $X=707290 $Y=29680
X1333 1 2 929 928 173 934 241 169 ICV_30 $T=721740 35360 1 0 $X=721550 $Y=32400
X1334 1 2 11 12 2 263 1 sky130_fd_sc_hd__and2_1 $T=21620 24480 0 0 $X=21430 $Y=24240
X1335 1 2 21 12 2 268 1 sky130_fd_sc_hd__and2_1 $T=29440 40800 0 0 $X=29250 $Y=40560
X1336 1 2 32 12 2 282 1 sky130_fd_sc_hd__and2_1 $T=48300 35360 1 0 $X=48110 $Y=32400
X1337 1 2 33 12 2 294 1 sky130_fd_sc_hd__and2_1 $T=49220 24480 0 0 $X=49030 $Y=24240
X1338 1 2 36 12 2 304 1 sky130_fd_sc_hd__and2_1 $T=67160 24480 0 0 $X=66970 $Y=24240
X1339 1 2 39 12 2 310 1 sky130_fd_sc_hd__and2_1 $T=76360 40800 1 0 $X=76170 $Y=37840
X1340 1 2 45 12 2 326 1 sky130_fd_sc_hd__and2_1 $T=90160 24480 0 0 $X=89970 $Y=24240
X1341 1 2 47 12 2 333 1 sky130_fd_sc_hd__and2_1 $T=95680 40800 1 0 $X=95490 $Y=37840
X1342 1 2 51 12 2 348 1 sky130_fd_sc_hd__and2_1 $T=104880 24480 1 0 $X=104690 $Y=21520
X1343 1 2 53 12 2 358 1 sky130_fd_sc_hd__and2_1 $T=115460 40800 0 0 $X=115270 $Y=40560
X1344 1 2 56 12 2 371 1 sky130_fd_sc_hd__and2_1 $T=125580 24480 0 0 $X=125390 $Y=24240
X1345 1 2 59 12 2 382 1 sky130_fd_sc_hd__and2_1 $T=137080 40800 1 0 $X=136890 $Y=37840
X1346 1 2 61 12 2 395 1 sky130_fd_sc_hd__and2_1 $T=156860 24480 1 0 $X=156670 $Y=21520
X1347 1 2 62 12 2 397 1 sky130_fd_sc_hd__and2_1 $T=157320 40800 0 0 $X=157130 $Y=40560
X1348 1 2 64 12 2 405 1 sky130_fd_sc_hd__and2_1 $T=160540 40800 1 0 $X=160350 $Y=37840
X1349 1 2 66 12 2 422 1 sky130_fd_sc_hd__and2_1 $T=171580 24480 0 0 $X=171390 $Y=24240
X1350 1 2 71 12 2 439 1 sky130_fd_sc_hd__and2_1 $T=192740 24480 1 0 $X=192550 $Y=21520
X1351 1 2 72 12 2 440 1 sky130_fd_sc_hd__and2_1 $T=192740 29920 1 0 $X=192550 $Y=26960
X1352 1 2 76 12 2 455 1 sky130_fd_sc_hd__and2_1 $T=202400 46240 0 0 $X=202210 $Y=46000
X1353 1 2 77 12 2 456 1 sky130_fd_sc_hd__and2_1 $T=207000 29920 1 0 $X=206810 $Y=26960
X1354 1 2 79 12 2 464 1 sky130_fd_sc_hd__and2_1 $T=209300 29920 1 0 $X=209110 $Y=26960
X1355 1 2 11 85 2 484 1 sky130_fd_sc_hd__and2_1 $T=228160 29920 1 0 $X=227970 $Y=26960
X1356 1 2 33 85 2 489 1 sky130_fd_sc_hd__and2_1 $T=235060 29920 0 0 $X=234870 $Y=29680
X1357 1 2 21 85 2 491 1 sky130_fd_sc_hd__and2_1 $T=237360 35360 0 0 $X=237170 $Y=35120
X1358 1 2 39 85 2 513 1 sky130_fd_sc_hd__and2_1 $T=258520 24480 1 0 $X=258330 $Y=21520
X1359 1 2 32 85 2 536 1 sky130_fd_sc_hd__and2_1 $T=270020 40800 1 0 $X=269830 $Y=37840
X1360 1 2 45 85 2 546 1 sky130_fd_sc_hd__and2_1 $T=280600 19040 1 0 $X=280410 $Y=16080
X1361 1 2 36 85 2 561 1 sky130_fd_sc_hd__and2_1 $T=293940 29920 1 0 $X=293750 $Y=26960
X1362 1 2 56 85 2 571 1 sky130_fd_sc_hd__and2_1 $T=302220 19040 0 0 $X=302030 $Y=18800
X1363 1 2 53 85 2 590 1 sky130_fd_sc_hd__and2_1 $T=325220 40800 1 0 $X=325030 $Y=37840
X1364 1 2 51 85 2 601 1 sky130_fd_sc_hd__and2_1 $T=326600 24480 0 0 $X=326410 $Y=24240
X1365 1 2 62 85 2 611 1 sky130_fd_sc_hd__and2_1 $T=340400 40800 1 0 $X=340210 $Y=37840
X1366 1 2 61 85 2 626 1 sky130_fd_sc_hd__and2_1 $T=350980 19040 0 0 $X=350790 $Y=18800
X1367 1 2 59 85 2 640 1 sky130_fd_sc_hd__and2_1 $T=367540 35360 0 0 $X=367350 $Y=35120
X1368 1 2 66 85 2 646 1 sky130_fd_sc_hd__and2_1 $T=370760 24480 0 0 $X=370570 $Y=24240
X1369 1 2 75 85 2 663 1 sky130_fd_sc_hd__and2_1 $T=382260 40800 0 0 $X=382070 $Y=40560
X1370 1 2 77 85 2 672 1 sky130_fd_sc_hd__and2_1 $T=386400 29920 0 0 $X=386210 $Y=29680
X1371 1 2 72 85 2 671 1 sky130_fd_sc_hd__and2_1 $T=389160 29920 1 0 $X=388970 $Y=26960
X1372 1 2 139 85 2 140 1 sky130_fd_sc_hd__and2_1 $T=401120 46240 1 0 $X=400930 $Y=43280
X1373 1 2 71 85 2 699 1 sky130_fd_sc_hd__and2_1 $T=409860 24480 1 0 $X=409670 $Y=21520
X1374 1 2 64 85 2 712 1 sky130_fd_sc_hd__and2_1 $T=423200 24480 0 0 $X=423010 $Y=24240
X1375 1 2 79 85 2 711 1 sky130_fd_sc_hd__and2_1 $T=423200 29920 0 0 $X=423010 $Y=29680
X1376 1 2 155 157 2 749 1 sky130_fd_sc_hd__and2_1 $T=462760 46240 0 0 $X=462570 $Y=46000
X1377 1 2 156 157 2 750 1 sky130_fd_sc_hd__and2_1 $T=463680 40800 1 0 $X=463490 $Y=37840
X1378 1 2 181 157 2 771 1 sky130_fd_sc_hd__and2_1 $T=497260 40800 1 0 $X=497070 $Y=37840
X1379 1 2 191 157 2 788 1 sky130_fd_sc_hd__and2_1 $T=519340 35360 0 0 $X=519150 $Y=35120
X1380 1 2 197 157 2 800 1 sky130_fd_sc_hd__and2_1 $T=534980 35360 0 0 $X=534790 $Y=35120
X1381 1 2 202 157 2 813 1 sky130_fd_sc_hd__and2_1 $T=550620 46240 1 0 $X=550430 $Y=43280
X1382 1 2 205 157 2 827 1 sky130_fd_sc_hd__and2_1 $T=568560 35360 0 0 $X=568370 $Y=35120
X1383 1 2 212 157 2 842 1 sky130_fd_sc_hd__and2_1 $T=592480 35360 0 0 $X=592290 $Y=35120
X1384 1 2 214 157 2 855 1 sky130_fd_sc_hd__and2_1 $T=609500 40800 1 0 $X=609310 $Y=37840
X1385 1 2 216 157 2 867 1 sky130_fd_sc_hd__and2_1 $T=627440 40800 0 0 $X=627250 $Y=40560
X1386 1 2 221 157 2 884 1 sky130_fd_sc_hd__and2_1 $T=649980 46240 1 0 $X=649790 $Y=43280
X1387 1 2 223 157 2 898 1 sky130_fd_sc_hd__and2_1 $T=665160 46240 0 0 $X=664970 $Y=46000
X1388 1 2 231 157 2 910 1 sky130_fd_sc_hd__and2_1 $T=690460 40800 1 0 $X=690270 $Y=37840
X1389 1 2 237 157 2 927 1 sky130_fd_sc_hd__and2_1 $T=714840 40800 0 0 $X=714650 $Y=40560
X1390 1 2 239 157 2 240 1 sky130_fd_sc_hd__and2_1 $T=718520 46240 1 0 $X=718330 $Y=43280
X1391 1 2 ICV_31 $T=45540 46240 1 0 $X=45350 $Y=43280
X1392 1 2 ICV_31 $T=59340 24480 0 0 $X=59150 $Y=24240
X1393 1 2 ICV_31 $T=73600 35360 1 0 $X=73410 $Y=32400
X1394 1 2 ICV_31 $T=101660 35360 1 0 $X=101470 $Y=32400
X1395 1 2 ICV_31 $T=103040 13600 1 0 $X=102850 $Y=10640
X1396 1 2 ICV_31 $T=131560 13600 1 0 $X=131370 $Y=10640
X1397 1 2 ICV_31 $T=171580 29920 0 0 $X=171390 $Y=29680
X1398 1 2 ICV_31 $T=174340 13600 1 0 $X=174150 $Y=10640
X1399 1 2 ICV_31 $T=283820 35360 0 0 $X=283630 $Y=35120
X1400 1 2 ICV_31 $T=339940 13600 0 0 $X=339750 $Y=13360
X1401 1 2 ICV_31 $T=339940 19040 0 0 $X=339750 $Y=18800
X1402 1 2 ICV_31 $T=359720 13600 1 0 $X=359530 $Y=10640
X1403 1 2 ICV_31 $T=373980 13600 1 0 $X=373790 $Y=10640
X1404 1 2 ICV_31 $T=431020 13600 1 0 $X=430830 $Y=10640
X1405 1 2 ICV_31 $T=459540 13600 1 0 $X=459350 $Y=10640
X1406 1 2 ICV_31 $T=480240 13600 0 0 $X=480050 $Y=13360
X1407 1 2 ICV_31 $T=494500 29920 1 0 $X=494310 $Y=26960
X1408 1 2 ICV_31 $T=502320 13600 1 0 $X=502130 $Y=10640
X1409 1 2 ICV_31 $T=516580 13600 1 0 $X=516390 $Y=10640
X1410 1 2 ICV_31 $T=606740 46240 1 0 $X=606550 $Y=43280
X1411 1 2 ICV_31 $T=620540 29920 0 0 $X=620350 $Y=29680
X1412 1 2 ICV_31 $T=648600 29920 0 0 $X=648410 $Y=29680
X1413 1 2 ICV_31 $T=662860 35360 1 0 $X=662670 $Y=32400
X1414 1 2 34 263 2 257 1 sky130_fd_sc_hd__dlclkp_1 $T=23920 29920 0 0 $X=23730 $Y=29680
X1415 1 2 34 268 2 256 1 sky130_fd_sc_hd__dlclkp_1 $T=24840 46240 0 0 $X=24650 $Y=46000
X1416 1 2 34 282 2 281 1 sky130_fd_sc_hd__dlclkp_1 $T=39560 40800 1 0 $X=39370 $Y=37840
X1417 1 2 34 294 2 280 1 sky130_fd_sc_hd__dlclkp_1 $T=51520 24480 0 0 $X=51330 $Y=24240
X1418 1 2 34 304 2 306 1 sky130_fd_sc_hd__dlclkp_1 $T=62560 29920 0 0 $X=62370 $Y=29680
X1419 1 2 34 310 2 309 1 sky130_fd_sc_hd__dlclkp_1 $T=69460 40800 1 0 $X=69270 $Y=37840
X1420 1 2 34 326 2 325 1 sky130_fd_sc_hd__dlclkp_1 $T=86020 29920 1 0 $X=85830 $Y=26960
X1421 1 2 34 333 2 332 1 sky130_fd_sc_hd__dlclkp_1 $T=93380 46240 1 0 $X=93190 $Y=43280
X1422 1 2 34 348 2 349 1 sky130_fd_sc_hd__dlclkp_1 $T=107180 24480 1 0 $X=106990 $Y=21520
X1423 1 2 34 358 2 354 1 sky130_fd_sc_hd__dlclkp_1 $T=115460 46240 1 0 $X=115270 $Y=43280
X1424 1 2 34 371 2 370 1 sky130_fd_sc_hd__dlclkp_1 $T=125580 29920 1 0 $X=125390 $Y=26960
X1425 1 2 34 382 2 383 1 sky130_fd_sc_hd__dlclkp_1 $T=136160 35360 1 0 $X=135970 $Y=32400
X1426 1 2 34 395 2 401 1 sky130_fd_sc_hd__dlclkp_1 $T=150420 24480 1 0 $X=150230 $Y=21520
X1427 1 2 34 397 2 60 1 sky130_fd_sc_hd__dlclkp_1 $T=150880 40800 0 0 $X=150690 $Y=40560
X1428 1 2 34 405 2 408 1 sky130_fd_sc_hd__dlclkp_1 $T=158240 35360 0 0 $X=158050 $Y=35120
X1429 1 2 34 422 2 414 1 sky130_fd_sc_hd__dlclkp_1 $T=171120 24480 1 0 $X=170930 $Y=21520
X1430 1 2 34 439 2 444 1 sky130_fd_sc_hd__dlclkp_1 $T=188140 24480 0 0 $X=187950 $Y=24240
X1431 1 2 34 440 2 437 1 sky130_fd_sc_hd__dlclkp_1 $T=189980 29920 0 0 $X=189790 $Y=29680
X1432 1 2 34 456 2 463 1 sky130_fd_sc_hd__dlclkp_1 $T=203320 29920 0 0 $X=203130 $Y=29680
X1433 1 2 34 455 2 78 1 sky130_fd_sc_hd__dlclkp_1 $T=204700 46240 0 0 $X=204510 $Y=46000
X1434 1 2 34 464 2 465 1 sky130_fd_sc_hd__dlclkp_1 $T=207920 24480 1 0 $X=207730 $Y=21520
X1435 1 2 34 489 2 492 1 sky130_fd_sc_hd__dlclkp_1 $T=231840 19040 0 0 $X=231650 $Y=18800
X1436 1 2 34 86 2 87 1 sky130_fd_sc_hd__dlclkp_1 $T=232300 46240 0 0 $X=232110 $Y=46000
X1437 1 2 34 491 2 496 1 sky130_fd_sc_hd__dlclkp_1 $T=232760 40800 0 0 $X=232570 $Y=40560
X1438 1 2 34 484 2 501 1 sky130_fd_sc_hd__dlclkp_1 $T=235980 29920 1 0 $X=235790 $Y=26960
X1439 1 2 34 513 2 518 1 sky130_fd_sc_hd__dlclkp_1 $T=251620 24480 0 0 $X=251430 $Y=24240
X1440 1 2 34 536 2 540 1 sky130_fd_sc_hd__dlclkp_1 $T=270020 35360 0 0 $X=269830 $Y=35120
X1441 1 2 34 112 2 105 1 sky130_fd_sc_hd__dlclkp_1 $T=272320 46240 0 0 $X=272130 $Y=46000
X1442 1 2 34 546 2 548 1 sky130_fd_sc_hd__dlclkp_1 $T=280140 24480 1 0 $X=279950 $Y=21520
X1443 1 2 34 561 2 565 1 sky130_fd_sc_hd__dlclkp_1 $T=293940 35360 1 0 $X=293750 $Y=32400
X1444 1 2 34 571 2 572 1 sky130_fd_sc_hd__dlclkp_1 $T=301300 24480 1 0 $X=301110 $Y=21520
X1445 1 2 34 590 2 586 1 sky130_fd_sc_hd__dlclkp_1 $T=318780 40800 1 0 $X=318590 $Y=37840
X1446 1 2 34 601 2 599 1 sky130_fd_sc_hd__dlclkp_1 $T=326140 19040 0 0 $X=325950 $Y=18800
X1447 1 2 34 611 2 615 1 sky130_fd_sc_hd__dlclkp_1 $T=335800 35360 0 0 $X=335610 $Y=35120
X1448 1 2 34 626 2 621 1 sky130_fd_sc_hd__dlclkp_1 $T=349140 24480 0 0 $X=348950 $Y=24240
X1449 1 2 34 640 2 638 1 sky130_fd_sc_hd__dlclkp_1 $T=362020 35360 1 0 $X=361830 $Y=32400
X1450 1 2 34 646 2 643 1 sky130_fd_sc_hd__dlclkp_1 $T=366160 24480 1 0 $X=365970 $Y=21520
X1451 1 2 34 663 2 665 1 sky130_fd_sc_hd__dlclkp_1 $T=384100 46240 0 0 $X=383910 $Y=46000
X1452 1 2 34 671 2 673 1 sky130_fd_sc_hd__dlclkp_1 $T=385940 24480 0 0 $X=385750 $Y=24240
X1453 1 2 34 672 2 678 1 sky130_fd_sc_hd__dlclkp_1 $T=388700 29920 0 0 $X=388510 $Y=29680
X1454 1 2 34 699 2 694 1 sky130_fd_sc_hd__dlclkp_1 $T=413080 24480 1 0 $X=412890 $Y=21520
X1455 1 2 34 711 2 717 1 sky130_fd_sc_hd__dlclkp_1 $T=422740 29920 1 0 $X=422550 $Y=26960
X1456 1 2 34 712 2 720 1 sky130_fd_sc_hd__dlclkp_1 $T=426880 24480 0 0 $X=426690 $Y=24240
X1457 1 2 34 147 2 718 1 sky130_fd_sc_hd__dlclkp_1 $T=426880 46240 0 0 $X=426690 $Y=46000
X1458 1 2 253 749 2 751 1 sky130_fd_sc_hd__dlclkp_1 $T=462300 46240 1 0 $X=462110 $Y=43280
X1459 1 2 253 750 2 752 1 sky130_fd_sc_hd__dlclkp_1 $T=463680 35360 0 0 $X=463490 $Y=35120
X1460 1 2 253 771 2 772 1 sky130_fd_sc_hd__dlclkp_1 $T=492660 35360 0 0 $X=492470 $Y=35120
X1461 1 2 253 788 2 786 1 sky130_fd_sc_hd__dlclkp_1 $T=517500 40800 1 0 $X=517310 $Y=37840
X1462 1 2 253 800 2 801 1 sky130_fd_sc_hd__dlclkp_1 $T=533600 40800 1 0 $X=533410 $Y=37840
X1463 1 2 253 813 2 815 1 sky130_fd_sc_hd__dlclkp_1 $T=550620 40800 0 0 $X=550430 $Y=40560
X1464 1 2 253 827 2 828 1 sky130_fd_sc_hd__dlclkp_1 $T=572700 40800 1 0 $X=572510 $Y=37840
X1465 1 2 253 842 2 843 1 sky130_fd_sc_hd__dlclkp_1 $T=591100 40800 1 0 $X=590910 $Y=37840
X1466 1 2 253 855 2 856 1 sky130_fd_sc_hd__dlclkp_1 $T=609500 40800 0 0 $X=609310 $Y=40560
X1467 1 2 253 867 2 872 1 sky130_fd_sc_hd__dlclkp_1 $T=629740 40800 0 0 $X=629550 $Y=40560
X1468 1 2 253 884 2 885 1 sky130_fd_sc_hd__dlclkp_1 $T=648600 40800 1 0 $X=648410 $Y=37840
X1469 1 2 253 898 2 897 1 sky130_fd_sc_hd__dlclkp_1 $T=665620 46240 1 0 $X=665430 $Y=43280
X1470 1 2 253 228 2 229 1 sky130_fd_sc_hd__dlclkp_1 $T=682180 46240 1 0 $X=681990 $Y=43280
X1471 1 2 253 910 2 908 1 sky130_fd_sc_hd__dlclkp_1 $T=688160 35360 0 0 $X=687970 $Y=35120
X1472 1 2 253 927 2 925 1 sky130_fd_sc_hd__dlclkp_1 $T=713460 40800 1 0 $X=713270 $Y=37840
X1473 1 2 257 17 271 ICV_35 $T=25300 19040 0 0 $X=25110 $Y=18800
X1474 1 2 257 20 276 ICV_35 $T=27600 29920 1 0 $X=27410 $Y=26960
X1475 1 2 281 8 292 ICV_35 $T=42320 35360 0 0 $X=42130 $Y=35120
X1476 1 2 281 19 283 ICV_35 $T=42780 29920 0 0 $X=42590 $Y=29680
X1477 1 2 281 20 298 ICV_35 $T=50600 35360 0 0 $X=50410 $Y=35120
X1478 1 2 306 20 311 ICV_35 $T=67620 19040 1 0 $X=67430 $Y=16080
X1479 1 2 354 19 375 ICV_35 $T=125580 40800 0 0 $X=125390 $Y=40560
X1480 1 2 370 20 377 ICV_35 $T=126500 19040 0 0 $X=126310 $Y=18800
X1481 1 2 383 20 400 ICV_35 $T=146280 35360 0 0 $X=146090 $Y=35120
X1482 1 2 60 4 63 ICV_35 $T=151800 46240 1 0 $X=151610 $Y=43280
X1483 1 2 401 6 407 ICV_35 $T=154100 13600 1 0 $X=153910 $Y=10640
X1484 1 2 401 9 410 ICV_35 $T=157780 24480 0 0 $X=157590 $Y=24240
X1485 1 2 463 9 469 ICV_35 $T=209760 29920 0 0 $X=209570 $Y=29680
X1486 1 2 492 90 506 ICV_35 $T=237820 13600 1 0 $X=237630 $Y=10640
X1487 1 2 496 88 499 ICV_35 $T=239660 35360 0 0 $X=239470 $Y=35120
X1488 1 2 492 99 515 ICV_35 $T=248400 13600 1 0 $X=248210 $Y=10640
X1489 1 2 492 100 516 ICV_35 $T=249780 13600 0 0 $X=249590 $Y=13360
X1490 1 2 501 101 519 ICV_35 $T=249780 29920 0 0 $X=249590 $Y=29680
X1491 1 2 87 102 522 ICV_35 $T=250700 46240 1 0 $X=250510 $Y=43280
X1492 1 2 518 91 530 ICV_35 $T=260820 24480 1 0 $X=260630 $Y=21520
X1493 1 2 518 101 533 ICV_35 $T=262660 13600 0 0 $X=262470 $Y=13360
X1494 1 2 548 102 568 ICV_35 $T=293940 19040 0 0 $X=293750 $Y=18800
X1495 1 2 572 88 580 ICV_35 $T=304520 19040 0 0 $X=304330 $Y=18800
X1496 1 2 572 102 583 ICV_35 $T=307740 24480 1 0 $X=307550 $Y=21520
X1497 1 2 121 88 587 ICV_35 $T=311420 46240 1 0 $X=311230 $Y=43280
X1498 1 2 572 90 594 ICV_35 $T=314640 13600 0 0 $X=314450 $Y=13360
X1499 1 2 121 102 603 ICV_35 $T=322000 46240 0 0 $X=321810 $Y=46000
X1500 1 2 125 88 625 ICV_35 $T=342700 46240 0 0 $X=342510 $Y=46000
X1501 1 2 125 99 628 ICV_35 $T=344540 46240 1 0 $X=344350 $Y=43280
X1502 1 2 673 88 677 ICV_35 $T=389160 19040 1 0 $X=388970 $Y=16080
X1503 1 2 673 99 683 ICV_35 $T=391000 13600 1 0 $X=390810 $Y=10640
X1504 1 2 752 160 756 ICV_35 $T=469200 29920 1 0 $X=469010 $Y=26960
X1505 1 2 180 162 774 ICV_35 $T=495420 46240 0 0 $X=495230 $Y=46000
X1506 1 2 772 159 783 ICV_35 $T=500940 35360 1 0 $X=500750 $Y=32400
X1507 1 2 786 165 789 ICV_35 $T=516120 29920 1 0 $X=515930 $Y=26960
X1508 1 2 815 171 821 ICV_35 $T=556600 35360 0 0 $X=556410 $Y=35120
X1509 1 2 815 162 823 ICV_35 $T=557060 40800 0 0 $X=556870 $Y=40560
X1510 1 2 815 170 824 ICV_35 $T=558440 24480 0 0 $X=558250 $Y=24240
X1511 1 2 843 161 852 ICV_35 $T=600760 29920 1 0 $X=600570 $Y=26960
X1512 1 2 856 172 863 ICV_35 $T=613640 29920 1 0 $X=613450 $Y=26960
X1513 1 2 213 171 864 ICV_35 $T=614560 46240 0 0 $X=614370 $Y=46000
X1514 1 2 897 172 904 ICV_35 $T=673900 29920 1 0 $X=673710 $Y=26960
X1515 1 2 925 165 929 ICV_35 $T=713000 35360 1 0 $X=712810 $Y=32400
X1516 1 2 280 18 299 ICV_36 $T=51520 19040 0 0 $X=51330 $Y=18800
X1517 1 2 349 19 360 ICV_36 $T=108560 29920 1 0 $X=108370 $Y=26960
X1518 1 2 354 8 373 ICV_36 $T=121440 35360 1 0 $X=121250 $Y=32400
X1519 1 2 54 4 57 ICV_36 $T=121900 46240 1 0 $X=121710 $Y=43280
X1520 1 2 370 19 385 ICV_36 $T=132480 29920 1 0 $X=132290 $Y=26960
X1521 1 2 383 6 387 ICV_36 $T=135700 29920 0 0 $X=135510 $Y=29680
X1522 1 2 408 6 415 ICV_36 $T=160540 35360 1 0 $X=160350 $Y=32400
X1523 1 2 444 20 453 ICV_36 $T=192740 19040 1 0 $X=192550 $Y=16080
X1524 1 2 496 101 520 ICV_36 $T=247940 35360 0 0 $X=247750 $Y=35120
X1525 1 2 125 100 612 ICV_36 $T=330280 46240 0 0 $X=330090 $Y=46000
X1526 1 2 599 99 616 ICV_36 $T=333960 13600 1 0 $X=333770 $Y=10640
X1527 1 2 615 100 633 ICV_36 $T=350060 29920 0 0 $X=349870 $Y=29680
X1528 1 2 638 101 644 ICV_36 $T=360180 29920 0 0 $X=359990 $Y=29680
X1529 1 2 786 160 791 ICV_36 $T=515200 29920 0 0 $X=515010 $Y=29680
X1530 1 2 192 172 198 ICV_36 $T=528080 46240 0 0 $X=527890 $Y=46000
X1531 1 2 199 162 812 ICV_36 $T=539120 46240 0 0 $X=538930 $Y=46000
X1532 1 2 843 171 851 ICV_36 $T=597540 40800 1 0 $X=597350 $Y=37840
X1533 1 2 856 165 859 ICV_36 $T=610420 29920 0 0 $X=610230 $Y=29680
X1534 1 2 925 172 938 ICV_36 $T=724500 29920 0 0 $X=724310 $Y=29680
X1535 1 2 257 4 269 ICV_37 $T=19780 24480 1 0 $X=19590 $Y=21520
X1536 1 2 257 9 265 ICV_37 $T=19780 29920 1 0 $X=19590 $Y=26960
X1537 1 2 306 6 320 ICV_37 $T=75900 19040 1 0 $X=75710 $Y=16080
X1538 1 2 309 20 319 ICV_37 $T=75900 46240 1 0 $X=75710 $Y=43280
X1539 1 2 332 19 353 ICV_37 $T=103960 40800 1 0 $X=103770 $Y=37840
X1540 1 2 349 6 367 ICV_37 $T=117760 13600 0 0 $X=117570 $Y=13360
X1541 1 2 349 8 365 ICV_37 $T=117760 24480 0 0 $X=117570 $Y=24240
X1542 1 2 354 17 368 ICV_37 $T=117760 35360 0 0 $X=117570 $Y=35120
X1543 1 2 354 9 366 ICV_37 $T=117760 40800 0 0 $X=117570 $Y=40560
X1544 1 2 50 18 55 ICV_37 $T=117760 46240 0 0 $X=117570 $Y=46000
X1545 1 2 54 9 381 ICV_37 $T=132020 46240 1 0 $X=131830 $Y=43280
X1546 1 2 401 20 411 ICV_37 $T=160080 19040 1 0 $X=159890 $Y=16080
X1547 1 2 401 19 412 ICV_37 $T=160080 24480 1 0 $X=159890 $Y=21520
X1548 1 2 437 4 445 ICV_37 $T=188140 35360 1 0 $X=187950 $Y=32400
X1549 1 2 437 6 446 ICV_37 $T=188140 46240 1 0 $X=187950 $Y=43280
X1550 1 2 444 18 462 ICV_37 $T=201940 13600 0 0 $X=201750 $Y=13360
X1551 1 2 437 9 460 ICV_37 $T=201940 40800 0 0 $X=201750 $Y=40560
X1552 1 2 465 20 476 ICV_37 $T=216200 19040 1 0 $X=216010 $Y=16080
X1553 1 2 465 9 474 ICV_37 $T=216200 24480 1 0 $X=216010 $Y=21520
X1554 1 2 463 20 475 ICV_37 $T=216200 35360 1 0 $X=216010 $Y=32400
X1555 1 2 463 4 479 ICV_37 $T=230000 24480 0 0 $X=229810 $Y=24240
X1556 1 2 501 88 497 ICV_37 $T=244260 29920 1 0 $X=244070 $Y=26960
X1557 1 2 518 88 542 ICV_37 $T=272320 24480 1 0 $X=272130 $Y=21520
X1558 1 2 548 90 557 ICV_37 $T=286120 13600 0 0 $X=285930 $Y=13360
X1559 1 2 548 91 556 ICV_37 $T=286120 19040 0 0 $X=285930 $Y=18800
X1560 1 2 540 101 117 ICV_37 $T=286120 29920 0 0 $X=285930 $Y=29680
X1561 1 2 565 99 575 ICV_37 $T=300380 40800 1 0 $X=300190 $Y=37840
X1562 1 2 572 100 573 ICV_37 $T=304980 13600 1 0 $X=304790 $Y=10640
X1563 1 2 121 101 582 ICV_37 $T=314180 46240 0 0 $X=313990 $Y=46000
X1564 1 2 599 88 607 ICV_37 $T=328440 24480 1 0 $X=328250 $Y=21520
X1565 1 2 615 88 624 ICV_37 $T=342240 29920 0 0 $X=342050 $Y=29680
X1566 1 2 615 102 622 ICV_37 $T=342240 35360 0 0 $X=342050 $Y=35120
X1567 1 2 621 102 639 ICV_37 $T=356500 24480 1 0 $X=356310 $Y=21520
X1568 1 2 130 102 641 ICV_37 $T=356500 46240 1 0 $X=356310 $Y=43280
X1569 1 2 643 99 653 ICV_37 $T=370300 13600 0 0 $X=370110 $Y=13360
X1570 1 2 643 100 655 ICV_37 $T=370300 19040 0 0 $X=370110 $Y=18800
X1571 1 2 665 100 667 ICV_37 $T=384560 35360 1 0 $X=384370 $Y=32400
X1572 1 2 665 88 676 ICV_37 $T=384560 40800 1 0 $X=384370 $Y=37840
X1573 1 2 665 89 674 ICV_37 $T=384560 46240 1 0 $X=384370 $Y=43280
X1574 1 2 673 100 691 ICV_37 $T=398360 13600 0 0 $X=398170 $Y=13360
X1575 1 2 665 101 693 ICV_37 $T=398360 35360 0 0 $X=398170 $Y=35120
X1576 1 2 678 91 706 ICV_37 $T=412620 29920 1 0 $X=412430 $Y=26960
X1577 1 2 720 101 737 ICV_37 $T=440680 19040 1 0 $X=440490 $Y=16080
X1578 1 2 751 159 753 ICV_37 $T=468740 40800 1 0 $X=468550 $Y=37840
X1579 1 2 180 165 787 ICV_37 $T=510600 40800 0 0 $X=510410 $Y=40560
X1580 1 2 786 171 798 ICV_37 $T=524860 40800 1 0 $X=524670 $Y=37840
X1581 1 2 801 165 805 ICV_37 $T=538660 29920 0 0 $X=538470 $Y=29680
X1582 1 2 204 170 207 ICV_37 $T=566720 46240 0 0 $X=566530 $Y=46000
X1583 1 2 843 160 848 ICV_37 $T=594780 29920 0 0 $X=594590 $Y=29680
X1584 1 2 843 162 847 ICV_37 $T=594780 35360 0 0 $X=594590 $Y=35120
X1585 1 2 856 162 869 ICV_37 $T=622840 35360 0 0 $X=622650 $Y=35120
X1586 1 2 872 162 880 ICV_37 $T=637100 40800 1 0 $X=636910 $Y=37840
X1587 1 2 897 171 899 ICV_37 $T=678960 35360 0 0 $X=678770 $Y=35120
X1588 1 2 229 170 926 ICV_37 $T=707020 40800 0 0 $X=706830 $Y=40560
X1589 1 2 238 159 934 ICV_37 $T=721280 46240 1 0 $X=721090 $Y=43280
X1590 1 2 325 17 331 325 18 337 ICV_38 $T=85560 19040 1 0 $X=85370 $Y=16080
X1591 1 2 370 9 378 370 8 384 ICV_38 $T=127880 24480 0 0 $X=127690 $Y=24240
X1592 1 2 463 8 487 463 6 490 ICV_38 $T=224020 35360 1 0 $X=223830 $Y=32400
X1593 1 2 105 99 529 105 102 539 ICV_38 $T=260820 40800 0 0 $X=260630 $Y=40560
X1594 1 2 565 88 579 565 102 585 ICV_38 $T=303600 29920 1 0 $X=303410 $Y=26960
X1595 1 2 615 99 623 615 101 617 ICV_38 $T=341780 29920 1 0 $X=341590 $Y=26960
X1596 1 2 615 91 635 615 90 634 ICV_38 $T=352820 35360 0 0 $X=352630 $Y=35120
X1597 1 2 158 159 163 751 162 762 ICV_38 $T=466900 46240 0 0 $X=466710 $Y=46000
X1598 1 2 772 161 773 772 170 784 ICV_38 $T=494960 24480 0 0 $X=494770 $Y=24240
X1599 1 2 204 161 826 204 171 829 ICV_38 $T=563040 46240 1 0 $X=562850 $Y=43280
X1600 1 2 872 159 873 872 171 883 ICV_38 $T=634340 35360 0 0 $X=634150 $Y=35120
X1601 1 2 885 170 890 885 172 896 ICV_38 $T=653200 24480 0 0 $X=653010 $Y=24240
X1602 1 2 229 160 914 229 172 916 ICV_38 $T=686320 40800 0 0 $X=686130 $Y=40560
X1603 1 2 908 165 920 908 161 924 ICV_38 $T=700580 29920 1 0 $X=700390 $Y=26960
X1604 1 2 238 165 242 238 171 940 ICV_38 $T=720360 46240 0 0 $X=720170 $Y=46000
X1605 1 2 3 4 10 ICV_47 $T=10580 46240 0 0 $X=10390 $Y=46000
X1606 1 2 280 17 287 ICV_47 $T=38640 19040 1 0 $X=38450 $Y=16080
X1607 1 2 280 6 293 ICV_47 $T=42780 19040 0 0 $X=42590 $Y=18800
X1608 1 2 280 4 300 ICV_47 $T=55200 19040 1 0 $X=55010 $Y=16080
X1609 1 2 309 4 328 ICV_47 $T=81880 35360 1 0 $X=81690 $Y=32400
X1610 1 2 325 9 340 ICV_47 $T=92460 24480 0 0 $X=92270 $Y=24240
X1611 1 2 332 20 347 ICV_47 $T=94760 40800 0 0 $X=94570 $Y=40560
X1612 1 2 383 19 388 ICV_47 $T=137080 35360 0 0 $X=136890 $Y=35120
X1613 1 2 383 18 393 ICV_47 $T=139380 40800 1 0 $X=139190 $Y=37840
X1614 1 2 401 18 409 ICV_47 $T=156860 13600 0 0 $X=156670 $Y=13360
X1615 1 2 408 18 418 ICV_47 $T=162840 29920 0 0 $X=162650 $Y=29680
X1616 1 2 408 20 419 ICV_47 $T=162840 40800 1 0 $X=162650 $Y=37840
X1617 1 2 414 17 424 ICV_47 $T=167900 19040 1 0 $X=167710 $Y=16080
X1618 1 2 414 8 432 ICV_47 $T=176180 29920 1 0 $X=175990 $Y=26960
X1619 1 2 444 9 459 ICV_47 $T=198720 24480 1 0 $X=198530 $Y=21520
X1620 1 2 78 9 471 ICV_47 $T=209760 40800 0 0 $X=209570 $Y=40560
X1621 1 2 78 4 488 ICV_47 $T=223100 40800 1 0 $X=222910 $Y=37840
X1622 1 2 492 102 521 ICV_47 $T=249780 24480 1 0 $X=249590 $Y=21520
X1623 1 2 496 102 525 ICV_47 $T=256220 40800 1 0 $X=256030 $Y=37840
X1624 1 2 565 101 562 ICV_47 $T=297620 24480 0 0 $X=297430 $Y=24240
X1625 1 2 638 102 650 ICV_47 $T=363400 40800 1 0 $X=363210 $Y=37840
X1626 1 2 141 100 698 ICV_47 $T=402960 40800 0 0 $X=402770 $Y=40560
X1627 1 2 694 91 701 ICV_47 $T=407560 19040 0 0 $X=407370 $Y=18800
X1628 1 2 694 102 714 ICV_47 $T=417680 19040 0 0 $X=417490 $Y=18800
X1629 1 2 720 100 741 ICV_47 $T=442060 13600 0 0 $X=441870 $Y=13360
X1630 1 2 146 100 151 ICV_47 $T=444360 46240 0 0 $X=444170 $Y=46000
X1631 1 2 752 162 761 ICV_47 $T=470120 35360 0 0 $X=469930 $Y=35120
X1632 1 2 192 161 793 ICV_47 $T=519340 46240 0 0 $X=519150 $Y=46000
X1633 1 2 828 172 839 ICV_47 $T=581440 29920 1 0 $X=581250 $Y=26960
X1634 1 2 856 160 860 ICV_47 $T=611800 40800 1 0 $X=611610 $Y=37840
X1635 1 2 897 160 907 ICV_47 $T=673440 46240 1 0 $X=673250 $Y=43280
X1636 1 2 925 170 933 ICV_47 $T=715760 29920 0 0 $X=715570 $Y=29680
X1637 1 2 238 170 932 ICV_47 $T=717140 40800 0 0 $X=716950 $Y=40560
X1638 1 2 70 69 14 67 9 447 ICV_51 $T=184460 46240 0 0 $X=184270 $Y=46000
X1639 1 2 424 438 25 444 17 449 ICV_51 $T=189980 13600 0 0 $X=189790 $Y=13360
X1640 1 2 457 442 30 78 18 467 ICV_51 $T=204700 40800 1 0 $X=204510 $Y=37840
X1641 1 2 474 468 16 465 17 481 ICV_51 $T=218500 19040 0 0 $X=218310 $Y=18800
X1642 1 2 494 498 93 501 90 494 ICV_51 $T=238280 29920 0 0 $X=238090 $Y=29680
X1643 1 2 497 498 94 501 89 509 ICV_51 $T=238740 24480 0 0 $X=238550 $Y=24240
X1644 1 2 541 543 104 548 101 547 ICV_51 $T=279220 13600 1 0 $X=279030 $Y=10640
X1645 1 2 555 113 93 114 89 567 ICV_51 $T=289340 40800 0 0 $X=289150 $Y=40560
X1646 1 2 562 563 108 565 100 564 ICV_51 $T=295320 29920 0 0 $X=295130 $Y=29680
X1647 1 2 593 595 108 599 101 593 ICV_51 $T=322000 13600 1 0 $X=321810 $Y=10640
X1648 1 2 616 595 107 621 88 630 ICV_51 $T=342700 19040 1 0 $X=342510 $Y=16080
X1649 1 2 634 618 93 130 101 648 ICV_51 $T=358340 40800 0 0 $X=358150 $Y=40560
X1650 1 2 636 631 97 638 100 649 ICV_51 $T=359720 29920 1 0 $X=359530 $Y=26960
X1651 1 2 684 685 94 678 102 696 ICV_51 $T=398820 29920 1 0 $X=398630 $Y=26960
X1652 1 2 686 670 106 141 90 144 ICV_51 $T=399740 46240 0 0 $X=399550 $Y=46000
X1653 1 2 792 195 168 192 165 802 ICV_51 $T=527160 46240 1 0 $X=526970 $Y=43280
X1654 1 2 317 318 27 ICV_53 $T=76360 35360 1 0 $X=76170 $Y=32400
X1655 1 2 319 318 28 ICV_53 $T=78660 40800 1 0 $X=78470 $Y=37840
X1656 1 2 322 316 15 ICV_53 $T=81420 24480 0 0 $X=81230 $Y=24240
X1657 1 2 377 379 28 ICV_53 $T=132480 19040 1 0 $X=132290 $Y=16080
X1658 1 2 378 379 16 ICV_53 $T=132480 24480 1 0 $X=132290 $Y=21520
X1659 1 2 479 473 14 ICV_53 $T=224480 24480 0 0 $X=224290 $Y=24240
X1660 1 2 499 500 94 ICV_53 $T=238740 35360 1 0 $X=238550 $Y=32400
X1661 1 2 523 498 107 ICV_53 $T=258520 29920 0 0 $X=258330 $Y=29680
X1662 1 2 539 103 106 ICV_53 $T=272780 46240 1 0 $X=272590 $Y=43280
X1663 1 2 547 543 108 ICV_53 $T=280600 13600 0 0 $X=280410 $Y=13360
X1664 1 2 556 543 97 ICV_53 $T=290720 24480 0 0 $X=290530 $Y=24240
X1665 1 2 581 574 107 ICV_53 $T=312800 13600 1 0 $X=312610 $Y=10640
X1666 1 2 598 595 104 ICV_53 $T=322920 13600 0 0 $X=322730 $Y=13360
X1667 1 2 612 126 104 ICV_53 $T=336720 40800 0 0 $X=336530 $Y=40560
X1668 1 2 620 595 97 ICV_53 $T=342700 24480 0 0 $X=342510 $Y=24240
X1669 1 2 637 631 98 ICV_53 $T=361100 19040 1 0 $X=360910 $Y=16080
X1670 1 2 644 645 108 ICV_53 $T=364780 24480 0 0 $X=364590 $Y=24240
X1671 1 2 726 148 98 ICV_53 $T=433320 46240 0 0 $X=433130 $Y=46000
X1672 1 2 933 928 178 ICV_53 $T=721740 29920 1 0 $X=721550 $Y=26960
X1673 1 2 260 261 14 ICV_63 $T=19320 46240 0 0 $X=19130 $Y=46000
X1674 1 2 262 261 16 ICV_63 $T=20240 46240 1 0 $X=20050 $Y=43280
X1675 1 2 301 291 15 ICV_63 $T=62100 24480 0 0 $X=61910 $Y=24240
X1676 1 2 302 278 16 ICV_63 $T=62100 35360 0 0 $X=61910 $Y=35120
X1677 1 2 43 44 25 ICV_63 $T=84640 46240 0 0 $X=84450 $Y=46000
X1678 1 2 48 49 14 ICV_63 $T=97980 46240 0 0 $X=97790 $Y=46000
X1679 1 2 392 379 13 ICV_63 $T=146280 13600 0 0 $X=146090 $Y=13360
X1680 1 2 402 394 15 ICV_63 $T=153640 35360 1 0 $X=153450 $Y=32400
X1681 1 2 403 404 14 ICV_63 $T=155020 19040 1 0 $X=154830 $Y=16080
X1682 1 2 411 404 28 ICV_63 $T=165600 13600 0 0 $X=165410 $Y=13360
X1683 1 2 410 404 16 ICV_63 $T=166060 24480 0 0 $X=165870 $Y=24240
X1684 1 2 469 473 16 ICV_63 $T=216660 29920 1 0 $X=216470 $Y=26960
X1685 1 2 505 502 98 ICV_63 $T=244720 24480 1 0 $X=244530 $Y=21520
X1686 1 2 516 502 104 ICV_63 $T=256680 13600 1 0 $X=256490 $Y=10640
X1687 1 2 628 126 107 ICV_63 $T=350980 46240 0 0 $X=350790 $Y=46000
X1688 1 2 633 618 104 ICV_63 $T=356960 35360 1 0 $X=356770 $Y=32400
X1689 1 2 135 136 104 ICV_63 $T=379500 46240 1 0 $X=379310 $Y=43280
X1690 1 2 677 679 94 ICV_63 $T=393300 19040 0 0 $X=393110 $Y=18800
X1691 1 2 683 679 107 ICV_63 $T=399280 13600 1 0 $X=399090 $Y=10640
X1692 1 2 727 723 98 ICV_63 $T=434240 35360 1 0 $X=434050 $Y=32400
X1693 1 2 779 782 179 ICV_63 $T=507380 40800 1 0 $X=507190 $Y=37840
X1694 1 2 836 834 178 ICV_63 $T=586500 29920 0 0 $X=586310 $Y=29680
X1695 1 2 847 846 174 ICV_63 $T=599380 40800 0 0 $X=599190 $Y=40560
X1696 1 2 865 215 168 ICV_63 $T=628820 46240 1 0 $X=628630 $Y=43280
X1697 1 2 899 900 179 ICV_63 $T=669760 40800 1 0 $X=669570 $Y=37840
X1698 1 2 921 909 174 ICV_63 $T=707480 35360 0 0 $X=707290 $Y=35120
X1699 1 2 940 241 179 ICV_63 $T=735540 35360 1 0 $X=735350 $Y=32400
X1700 1 2 5 2 7 1 sky130_fd_sc_hd__clkbuf_4 $T=12880 13600 1 0 $X=12690 $Y=10640
X1701 1 2 24 2 26 1 sky130_fd_sc_hd__clkbuf_4 $T=35420 13600 0 0 $X=35230 $Y=13360
X1702 1 2 73 2 74 1 sky130_fd_sc_hd__clkbuf_4 $T=198260 13600 1 0 $X=198070 $Y=10640
X1703 1 2 83 2 84 1 sky130_fd_sc_hd__clkbuf_4 $T=224020 13600 0 0 $X=223830 $Y=13360
X1704 1 2 92 2 95 1 sky130_fd_sc_hd__clkbuf_4 $T=241500 19040 1 0 $X=241310 $Y=16080
X1705 1 2 109 2 110 1 sky130_fd_sc_hd__clkbuf_4 $T=269100 24480 1 0 $X=268910 $Y=21520
X1706 1 2 115 2 116 1 sky130_fd_sc_hd__clkbuf_4 $T=292100 13600 1 0 $X=291910 $Y=10640
X1707 1 2 122 2 123 1 sky130_fd_sc_hd__clkbuf_4 $T=314640 19040 0 0 $X=314450 $Y=18800
X1708 1 2 127 2 128 1 sky130_fd_sc_hd__clkbuf_4 $T=342700 13600 0 0 $X=342510 $Y=13360
X1709 1 2 133 2 134 1 sky130_fd_sc_hd__clkbuf_4 $T=367540 19040 0 0 $X=367350 $Y=18800
X1710 1 2 137 2 138 1 sky130_fd_sc_hd__clkbuf_4 $T=386400 13600 0 0 $X=386210 $Y=13360
X1711 1 2 142 2 143 1 sky130_fd_sc_hd__clkbuf_4 $T=406180 13600 1 0 $X=405990 $Y=10640
X1712 1 2 149 2 150 1 sky130_fd_sc_hd__clkbuf_4 $T=442060 13600 1 0 $X=441870 $Y=10640
X1713 1 2 153 2 154 1 sky130_fd_sc_hd__clkbuf_4 $T=460920 13600 0 0 $X=460730 $Y=13360
X1714 1 2 164 2 166 1 sky130_fd_sc_hd__clkbuf_4 $T=476560 13600 1 0 $X=476370 $Y=10640
X1715 1 2 175 2 176 1 sky130_fd_sc_hd__clkbuf_4 $T=490820 13600 1 0 $X=490630 $Y=10640
X1716 1 2 182 2 183 1 sky130_fd_sc_hd__clkbuf_4 $T=499560 13600 1 0 $X=499370 $Y=10640
X1717 1 2 187 2 188 1 sky130_fd_sc_hd__clkbuf_4 $T=511060 13600 1 0 $X=510870 $Y=10640
X1718 1 2 189 2 190 1 sky130_fd_sc_hd__clkbuf_4 $T=513820 13600 1 0 $X=513630 $Y=10640
X1719 1 2 193 2 194 1 sky130_fd_sc_hd__clkbuf_4 $T=523940 13600 1 0 $X=523750 $Y=10640
X1720 1 2 200 2 201 1 sky130_fd_sc_hd__clkbuf_4 $T=547860 13600 1 0 $X=547670 $Y=10640
X1721 1 2 218 2 219 1 sky130_fd_sc_hd__clkbuf_4 $T=639400 13600 1 0 $X=639210 $Y=10640
X1722 1 2 222 2 224 1 sky130_fd_sc_hd__clkbuf_4 $T=664240 13600 1 0 $X=664050 $Y=10640
X1723 1 2 230 2 232 1 sky130_fd_sc_hd__clkbuf_4 $T=685400 13600 1 0 $X=685210 $Y=10640
X1724 1 2 235 2 236 1 sky130_fd_sc_hd__clkbuf_4 $T=710700 13600 1 0 $X=710510 $Y=10640
X1725 1 2 243 2 244 1 sky130_fd_sc_hd__clkbuf_4 $T=733700 13600 1 0 $X=733510 $Y=10640
X1726 1 2 ICV_89 $T=20240 13600 1 0 $X=20050 $Y=10640
X1727 1 2 ICV_89 $T=34500 13600 1 0 $X=34310 $Y=10640
X1728 1 2 ICV_89 $T=48760 13600 1 0 $X=48570 $Y=10640
X1729 1 2 ICV_89 $T=63020 13600 1 0 $X=62830 $Y=10640
X1730 1 2 ICV_89 $T=77280 13600 1 0 $X=77090 $Y=10640
X1731 1 2 ICV_89 $T=105800 13600 1 0 $X=105610 $Y=10640
X1732 1 2 ICV_89 $T=134320 13600 1 0 $X=134130 $Y=10640
X1733 1 2 ICV_89 $T=454940 24480 1 0 $X=454750 $Y=21520
X1734 1 2 ICV_89 $T=462300 13600 1 0 $X=462110 $Y=10640
X1735 1 2 ICV_89 $T=533600 13600 1 0 $X=533410 $Y=10640
X1736 1 2 ICV_89 $T=562120 13600 1 0 $X=561930 $Y=10640
X1737 1 2 ICV_89 $T=576380 13600 1 0 $X=576190 $Y=10640
X1738 1 2 ICV_89 $T=590640 13600 1 0 $X=590450 $Y=10640
X1739 1 2 ICV_89 $T=604900 13600 1 0 $X=604710 $Y=10640
X1740 1 2 ICV_89 $T=619160 13600 1 0 $X=618970 $Y=10640
X1741 1 2 ICV_89 $T=647680 13600 1 0 $X=647490 $Y=10640
X1742 1 2 ICV_89 $T=690460 13600 1 0 $X=690270 $Y=10640
X1743 1 2 ICV_89 $T=718980 13600 1 0 $X=718790 $Y=10640
X1744 1 2 ICV_90 $T=6900 13600 0 0 $X=6710 $Y=13360
X1745 1 2 ICV_90 $T=38180 13600 0 0 $X=37990 $Y=13360
X1746 1 2 ICV_91 $T=210680 46240 1 0 $X=210490 $Y=43280
X1747 1 2 ICV_92 $T=469200 24480 1 0 $X=469010 $Y=21520
X1748 1 2 ICV_92 $T=609500 24480 1 0 $X=609310 $Y=21520
X1749 1 2 ICV_92 $T=679420 24480 0 0 $X=679230 $Y=24240
X1750 1 2 ICV_92 $T=693680 19040 1 0 $X=693490 $Y=16080
X1751 1 2 ICV_92 $T=707480 13600 0 0 $X=707290 $Y=13360
X1752 1 2 ICV_93 $T=454940 19040 0 0 $X=454750 $Y=18800
X1753 1 2 ICV_93 $T=469200 19040 1 0 $X=469010 $Y=16080
X1754 1 2 ICV_93 $T=483000 13600 0 0 $X=482810 $Y=13360
X1755 1 2 ICV_93 $T=511060 19040 0 0 $X=510870 $Y=18800
X1756 1 2 ICV_93 $T=525320 19040 1 0 $X=525130 $Y=16080
X1757 1 2 ICV_93 $T=539120 13600 0 0 $X=538930 $Y=13360
X1758 1 2 ICV_93 $T=567180 19040 0 0 $X=566990 $Y=18800
X1759 1 2 ICV_93 $T=581440 19040 1 0 $X=581250 $Y=16080
X1760 1 2 ICV_93 $T=595240 13600 0 0 $X=595050 $Y=13360
X1761 1 2 ICV_93 $T=623300 19040 0 0 $X=623110 $Y=18800
X1762 1 2 ICV_93 $T=637560 19040 1 0 $X=637370 $Y=16080
X1763 1 2 ICV_93 $T=651360 13600 0 0 $X=651170 $Y=13360
X1764 1 2 ICV_93 $T=665620 24480 1 0 $X=665430 $Y=21520
X1765 1 2 ICV_93 $T=679420 19040 0 0 $X=679230 $Y=18800
.ENDS
***************************************
.SUBCKT DFFRAM VGND VPWR EN Di[0] Di[1] Di[2] Di[3] Di[4] Di[5] Di[6] Di[7] Di[8] Di[9] Di[10] Di[11] Di[12] Di[13] Di[14] Di[15] Di[16]
+ Di[17] Di[18] Di[19] Di[20] Di[21] Di[22] Di[23] Di[24] Di[25] Di[26] Di[27] Di[28] Di[29] Di[30] Di[31] A[0] A[2] A[6] A[7] A[1]
+ Do[2] Do[3] Do[4] Do[7] Do[6] Do[5] Do[0] Do[1] Do[8] Do[9] Do[10] Do[11] Do[12] Do[13] Do[14] Do[15] Do[16] Do[17] Do[18] Do[19]
+ Do[20] Do[21] Do[22] Do[23] Do[24] Do[25] Do[26] Do[27] Do[28] Do[29] Do[30] Do[31] WE[3] WE[1] WE[2] CLK WE[0] A[5] A[3] A[4]
** N=1516 EP=80 IP=3742 FDC=358817
X0 VGND VPWR Dpar a=2090.79 p=1485.14 m=1 $[nwdiode] $X=5330 $Y=47545 $D=191
X1 VGND VPWR Dpar a=2090.3 p=1485.74 m=1 $[nwdiode] $X=5330 $Y=112825 $D=191
X2 VGND VPWR Dpar a=2090.38 p=1485.64 m=1 $[nwdiode] $X=5330 $Y=178105 $D=191
X3 VGND VPWR Dpar a=2090.3 p=1485.74 m=1 $[nwdiode] $X=5330 $Y=243385 $D=191
X4 VGND VPWR 3 57 WE[3] 22 4 26 6 59 56 7 12 14 28 9 Di[0] 11 15 36
+ 13 23 17 31 16 20 19 21 18 25 66 32 27 67 30 Di[1] 29 35 68 39
+ 33 37 38 Di[2] 42 52 40 44 72 41 60 Di[3] 83 573 51 71 45 49 46 47
+ 48 89 Di[4] 55 53 65 54 128 58 61 82 64 62 70 Di[5] 646 69 81 76 74
+ 79 75 78 73 98 105 Di[6] 92 95 80 84 85 86 87 113 104 90 91 88 99
+ 93 103 94 96 Di[7] 100 101 102 106 109 108 107 111 112 Di[8] 120 124 114 119 115
+ 133 164 Di[9] 116 118 156 137 131 121 122 Di[10] 126 125 130 127 Di[11] 132 134 135 136
+ Di[12] 139 140 158 141 153 Di[13] 143 145 146 162 169 144 150 165 157 149 147 148 159
+ 167 163 175 180 174 151 188 152 171 173 170 Di[14] 154 160 161 182 195 177 168 Di[15]
+ 181 172 179 178 196 184 186 194 185 183 Di[16] 189 190 191 192 193 202 198 197 203
+ 200 Di[17] 201 204 209 210 206 205 274 208 Di[18] 218 215 212 219 213 211 214 216 Di[19]
+ 236 231 223 220 221 222 238 234 225 235 224 230 226 232 Di[20] 237 229 228 233 247
+ 166 239 248 244 240 Di[21] 243 245 242 246 250 249 251 Di[22] 261 254 256 257 252 255
+ 280 258 263 268 259 260 262 272 270 264 265 266 273 Di[23] 271 267 275 Di[24] 278 277
+ 279 Di[25] 284 282 281 285 287 286 291 Di[26] 289 292 293 295 Di[27] 296 297 300 298 299
+ 305 Di[28] 301 303 304 307 Di[29] 310 306 311 308 312 313 Di[30] 315 316 317 Di[31] 319 10
+ ICV_55 $T=0 0 0 0 $X=0 $Y=443100
X5 VGND VPWR 320 WE[1] 3 324 349 22 4 26 6 344 12 321 9 36 28 323 WE[2] 11
+ 322 326 16 23 13 14 402 15 31 20 19 348 325 21 18 25 32 27 340 342
+ 327 362 30 328 329 351 330 33 331 347 332 38 339 37 363 40 361 41 333 365
+ 334 587 335 45 355 336 337 338 122 46 47 134 343 341 49 352 366 54 360 357
+ 364 723 345 346 350 135 64 55 58 56 59 35 353 354 62 356 368 358 359 51
+ 65 66 48 67 367 69 76 73 75 74 78 98 105 109 370 373 79 86 87 84
+ 369 104 85 113 88 90 91 103 93 94 95 96 372 101 371 52 106 375 107 111
+ 108 374 376 377 378 380 118 116 379 82 381 119 70 121 384 120 127 385 126 387
+ 125 132 102 386 389 114 130 390 391 393 392 136 397 395 139 140 89 141 398 169
+ 17 394 157 400 399 143 149 162 401 423 404 173 144 396 165 145 382 388 150 418
+ 411 146 403 153 415 409 383 29 405 406 407 416 148 408 161 147 413 160 412 188
+ 437 435 152 158 414 151 174 167 154 442 417 175 159 410 426 427 424 189 180 422
+ 419 420 421 168 177 242 425 172 433 431 178 163 184 428 429 183 430 185 432 438
+ 434 191 290 193 192 202 436 439 440 200 197 198 441 443 454 204 444 206 457 445
+ 446 448 447 453 274 205 450 451 452 208 461 211 458 455 456 214 213 216 459 222
+ 473 223 462 465 221 226 234 469 464 468 470 467 463 238 475 224 225 471 229 232
+ 230 233 480 472 235 476 460 487 239 247 477 240 243 244 482 246 245 478 479 484
+ 481 483 258 236 271 485 203 210 249 181 215 511 251 486 268 449 257 252 256 254
+ 488 190 272 186 280 270 261 260 466 231 264 259 218 489 492 474 490 263 209 194
+ 262 491 237 171 265 501 506 504 505 493 510 502 496 498 499 250 508 494 266 497
+ 273 500 507 495 503 516 509 195 275 512 277 513 278 514 515 517 518 285 281 284
+ 519 522 520 289 286 287 521 523 292 524 291 296 525 295 526 293 527 297 528 298
+ 300 301 299 303 529 304 532 530 306 307 305 531 533 308 310 534 535 311 312 313
+ 536 317 316 538 537 10 166
+ ICV_67 $T=0 0 0 0 $X=0 $Y=377800
X6 VGND VPWR 624 A[6] A[7] 359 488 WE[0] 320 4 6 EN 539 542 544 326 57 543 541 12
+ 540 321 14 553 549 59 323 556 585 56 22 322 23 545 15 554 547 13 546 20
+ 548 558 550 551 28 31 19 325 21 552 555 559 329 563 25 342 557 66 32 561
+ 327 67 16 560 562 566 328 68 35 26 565 567 564 351 36 331 332 39 381 568
+ 42 569 334 333 570 571 572 71 60 335 83 588 51 574 337 575 336 338 576 341
+ 578 61 A[0] 579 345 89 350 360 135 346 A[2] 339 347 A[1] 581 349 353 582 128 65
+ 358 356 354 340 70 586 52 355 723 134 122 81 587 357 361 363 365 324 589 362
+ 109 119 92 76 590 72 120 367 102 591 114 75 593 82 592 98 343 113 CLK 369
+ 78 99 88 594 398 611 87 595 370 599 598 597 596 85 105 86 90 600 603 103
+ 91 601 602 604 93 605 606 104 609 607 608 376 94 95 371 610 612 616 613 10
+ 614 372 373 615 375 374 618 617 619 377 385 378 620 380 379 621 623 622 625 626
+ 627 628 629 743 384 630 631 632 386 389 634 633 635 387 638 640 636 637 395 390
+ 639 391 392 641 642 393 397 80 643 645 53 644 400 647 100 646 399 573 44 423
+ 408 401 435 404 416 407 409 415 405 648 151 414 412 406 427 166 442 649 650 424
+ 194 411 170 413 171 196 418 163 654 651 212 422 419 420 181 437 179 653 655 652
+ 228 656 267 201 255 657 658 660 659 426 661 428 662 182 665 433 186 663 432 434
+ 190 664 430 431 666 667 436 668 439 195 290 440 446 441 203 202 445 454 444 209
+ 220 669 451 452 218 447 448 210 670 215 450 219 457 461 214 671 455 456 458 672
+ 459 673 236 231 674 469 462 464 463 467 675 468 470 471 237 676 472 677 250 478
+ 678 476 477 7 482 248 498 473 247 483 479 429 480 481 485 484 499 500 496 497
+ 680 453 417 425 511 682 502 501 508 507 487 503 681 516 509 438 506 510 443 683
+ 492 505 684 504 465 513 685 495 494 686 493 514 512 515 687 517 518 688 689 690
+ 519 520 521 522 691 692 524 523 525 526 527 693 528 529 530 695 534 533 532 238
+ 531 535 694 696 697 698 536 538 699 537
+ ICV_75 $T=0 0 0 0 $X=0 $Y=312560
X7 VGND VPWR 344 542 539 585 541 349 540 544 543 700 546 549 324 545 554 547 556 348
+ 548 701 702 558 551 550 552 561 555 557 703 706 563 559 362 326 553 704 560 330
+ 705 566 562 14 707 564 568 347 570 565 567 708 340 351 709 710 365 52 711 363
+ A[6] 569 72 361 571 572 355 712 713 574 714 122 134 721 576 343 575 716 715 48
+ 717 578 352 718 579 587 719 135 592 366 720 582 581 364 722 586 591 82 81 589
+ 590 92 99 102 10 114 594 598 596 595 599 597 593 726 724 727 611 602 600 601
+ 603 604 605 725 606 609 607 608 731 610 616 729 728 614 612 613 617 615 623 730
+ 734 621 733 618 732 738 736 633 83 735 619 620 622 625 740 741 629 748 750 70
+ 746 634 744 632 631 635 636 637 745 747 641 642 749 644 643 751 398 437 645 427
+ 752 739 753 754 435 409 755 415 647 756 737 405 757 648 760 758 759 442 630 788
+ 424 410 321 A[7] 761 414 649 763 416 762 417 404 407 777 423 401 399 412 764 663
+ 400 765 766 156 742 767 639 786 772 768 769 771 421 770 776 652 790 783 319 773
+ 774 164 775 655 425 782 654 289 785 779 780 781 431 658 315 784 787 301 778 659
+ 793 789 429 792 662 791 296 796 665 664 279 438 282 666 794 797 798 795 668 808
+ 657 306 799 490 816 801 661 443 800 804 491 803 812 805 802 822 669 806 840 453
+ 670 857 807 656 867 809 449 829 813 811 810 823 671 465 815 864 672 820 814 667
+ 842 460 673 818 674 877 846 475 821 817 819 651 675 466 824 841 825 827 832 845
+ 830 828 473 676 831 677 872 653 870 851 474 833 834 678 869 868 839 835 487 502
+ 836 855 847 837 498 849 871 843 505 844 856 501 660 504 511 489 838 680 848 850
+ 854 852 826 499 853 650 497 506 500 508 486 860 682 858 681 859 865 516 510 509
+ 861 862 507 863 683 503 684 685 866 686 873 874 880 878 876 875 496 879 881 882
+ 687 886 883 884 885 888 887 688 689 889 690 892 890 891 898 692 893 908 691 894
+ 895 896 897 693 900 899 902 901 903 919 694 904 905 695 697 696 910 698 906 907
+ 909 912 699 913 911 914 918 916 915 917 166
+ ICV_78 $T=0 0 0 0 $X=0 $Y=244560
X8 VGND VPWR 702 700 544 539 542 546 928 920 923 922 921 549 926 924 701 554 925 550
+ 551 935 939 543 558 938 941 934 17 927 933 545 930 932 937 936 929 940 559 557
+ 563 340 541 949 957 547 704 942 944 945 703 561 705 951 707 706 947 946 948 708
+ 29 950 952 339 Do[2] 556 956 709 710 711 954 381 713 955 960 962 963 961 712 959
+ 44 573 588 966 Do[3] 714 716 964 967 717 965 972 970 715 A[5] 553 718 721 354 969
+ 977 723 719 971 53 973 70 720 722 976 974 978 975 980 368 979 646 984 982 80
+ 983 981 992 100 987 585 398 594 991 598 985 595 989 986 605 724 597 599 A[6] 761
+ A[7] 604 990 Do[5] 726 607 608 609 606 758 603 616 611 993 614 613 612 995 730 725
+ 762 729 728 727 996 731 994 943 1000 732 756 755 997 Do[6] 1019 733 999 1002 1001 1004
+ 1003 1007 1005 736 1012 735 738 1006 734 Do[4] 757 737 1009 1105 1010 1013 1008 1011 1016 1018
+ 1017 1015 Do[7] 739 1029 626 1014 627 382 396 1021 1023 1022 741 1020 1033 740 1028 1026 1024
+ 1025 1032 1027 1037 742 628 759 1030 383 1031 1086 1085 1034 1035 1038 743 1036 778 388 744
+ 1039 1041 1040 1087 7 745 746 640 780 747 793 1089 394 1092 789 748 1042 1043 749 750
+ 1076 1044 1098 751 638 931 1101 1045 403 753 771 752 1046 754 1084 112 137 1097 1077 1073
+ 1048 1078 1047 1091 784 785 10 779 115 131 133 1049 124 760 1053 1079 767 769 765 766
+ 1122 1081 1051 1050 764 1052 774 777 768 1056 1055 770 782 772 775 776 790 781 1054 1058
+ 1066 315 1062 1057 1059 1060 1063 1064 786 788 787 1061 1065 1069 792 791 1067 783 1068 1120
+ 319 797 1074 279 794 796 306 1070 1071 795 1072 289 798 799 803 1117 189 804 805 1075
+ 806 1080 1111 1082 808 809 816 1088 1083 810 1090 811 1093 1094 1096 1095 1099 1106 1100 1147
+ 1109 1103 1102 815 817 819 820 1104 824 1112 1107 1108 828 842 827 1110 1121 851 830 1113
+ 833 829 835 839 869 868 228 836 855 1114 1115 845 841 846 872 1116 212 255 201 843
+ 849 847 871 857 1118 1119 856 1124 854 867 1130 1125 1126 1123 1129 860 862 861 1127 866
+ 1128 1133 1131 1132 1134 1136 1135 1139 1137 874 1140 1141 873 1138 1149 875 1160 876 1144 878
+ 1146 1156 1145 1143 879 882 883 1148 901 1172 1153 1142 1150 884 885 1154 886 1151 888 1152
+ 1155 1157 890 891 1158 1159 1163 1161 899 893 1171 1164 1165 1162 894 1167 1166 1169 1168 897
+ 1170 900 1173 902 1174 1176 1175 903 904 905 1177 906 1178 907 910 911 909 1179 912 913
+ 914 915 1180 916 918 917 919
+ ICV_79 $T=0 0 0 0 $X=0 $Y=179280
X9 VGND VPWR A[3] 1181 921 920 1182 922 923 321 925 1183 924 358 926 1187 1185 938 933 941
+ 934 1190 927 1188 1184 932 930 936 937 928 935 957 1198 1186 940 1189 949 945 1191 942
+ 1194 1197 1032 1193 1192 944 1040 1195 946 950 947 951 1203 1196 1200 1205 954 1202 952 1207
+ 1201 955 1199 1204 960 962 959 1209 961 1206 1036 963 1208 964 1228 1213 1211 1215 1214 967
+ 1217 A[4] 1212 970 1210 969 1218 356 971 1224 1230 1216 976 1220 1020 1221 975 1234 1225 1222
+ 978 1231 1223 1053 1232 979 1229 1226 1227 981 931 982 1238 1233 986 985 991 1237 987 1244
+ 1235 989 990 965 994 1247 993 995 1240 1239 1241 1243 1242 1411 1254 1248 1001 354 996 997
+ 1246 999 1255 112 124 1002 1236 1245 115 1013 1004 1252 1006 1003 1005 1007 133 1249 164 398
+ 1250 1012 1009 156 1251 1010 1011 A[6] 1253 624 137 1015 A[7] 1028 1016 1029 1014 1017 1018 1256
+ 131 1025 1258 1257 1021 1033 402 1023 1026 948 1262 1027 1280 1274 1261 1259 1267 1260 1030 1276
+ 1264 1031 1270 1271 1080 1266 1286 1263 956 1279 1289 1035 1283 1074 1265 1291 929 1038 1037 1268
+ 1269 1041 1273 1272 1275 1277 1278 973 1043 1044 1045 1281 1282 972 1047 1048 974 1284 1049 1285
+ 1287 1288 1054 1055 1051 1290 1059 1056 1292 1058 1293 1060 1000 1062 1065 201 1294 1067 1299 1296
+ 1295 212 1068 1297 1298 992 1302 1071 1301 1072 1300 1019 801 1305 282 296 1303 301 1075 1304
+ 1073 220 1097 242 1308 807 267 255 1083 1081 1082 1307 1306 1076 1077 1079 228 1078 1100 1085
+ 1095 1096 1091 1086 1087 1088 1084 822 1089 1101 1090 812 1310 1093 1094 1092 1311 1309 1103 1098
+ 1312 1106 814 1099 1105 7 853 1102 821 816 844 1314 775 831 1104 840 829 1313 1342 1315
+ 1329 1320 1328 1331 1321 1107 1318 1050 1108 1069 1330 832 826 1338 1057 1323 1322 1334 1317 1327
+ 1316 850 1052 1110 1333 1111 1066 858 1319 851 1335 848 1324 1326 1064 1325 1063 839 868 869
+ 837 835 838 817 1114 1115 1336 855 1332 A[2] 846 1116 1119 A[0] 847 857 856 774 849 871
+ 798 1118 A[1] 842 867 1133 845 1120 841 808 1337 1070 1117 859 1123 1124 1061 1340 1122 863
+ 1128 1339 854 1343 1341 1136 864 1135 1127 796 830 823 1344 1109 1126 1130 1112 1143 1129 1125
+ 1138 1132 1131 872 784 786 1121 1134 1345 279 789 1346 870 1137 788 1141 1146 1348 1140 1139
+ 896 1347 1351 877 793 1349 1350 1142 777 1147 1144 881 1145 892 790 880 1353 1352 1356 1148
+ 783 1113 1149 1150 1354 785 901 1355 887 1172 1153 1152 1151 1357 889 1156 289 1359 1154 1155
+ 1358 1163 1159 899 1157 1158 1167 895 898 1360 1169 1161 908 1160 1361 1162 1365 1164 1362 1165
+ 1166 1168 1170 1363 1364 306 1171 1366 1367 1368 1372 1369 1370 1173 1371 1174 1374 1373 1176 1175
+ 315 1177 1375 1178 1376 1179 319 1377 1378 1180 1380 1379
+ ICV_83 $T=0 0 0 0 $X=0 $Y=114000
X10 VGND VPWR 1181 1182 1251 1236 1382 1256 1384 1381 1025 1185 1184 1192 939 935 1031 1250 1183 1036
+ 1190 1188 929 1253 1249 1186 1245 1194 1383 1020 1191 1040 1252 1028 1385 1032 948 1193 1196 1386
+ 1197 1202 1189 1195 1387 1203 1392 954 956 951 1199 1388 1389 1206 963 1201 1391 1209 1390 1204
+ 966 1394 1393 1395 965 1208 1211 1210 938 1216 972 1396 1212 1397 1398 973 1217 1215 977 1399
+ 931 1400 1228 974 1401 1221 980 1220 1402 1403 1222 937 978 983 1223 945 1404 1227 984 1234
+ 1226 1405 1232 992 1406 1238 1235 1244 1053 1233 989 1407 1408 1409 1237 A[2] 1242 A[1] 1241 1239
+ 1243 1231 358 356 354 1246 1000 1410 1019 1198 1187 1229 1224 1001 1205 1412 1411 1225 1413 1255
+ 1248 1207 1247 1230 1240 1213 A[0] 1214 1414 1254 1200 1002 1218 1262 1415 1016 1005 1029 1257 1006
+ 1417 1258 1416 1280 1018 1274 1259 1267 1264 1021 1279 1260 1017 1010 1003 1418 1270 1013 1261 1286
+ 1007 1033 1080 1266 1271 1283 1011 1023 1012 1263 1026 1291 1074 1276 1289 1265 1419 1272 1268 1420
+ 1422 1269 1421 1273 1424 1423 1275 1425 1277 1426 1278 1427 1428 1429 1281 1430 1282 1284 1431 1285
+ 1432 1287 1288 1433 1434 1436 1290 1435 1292 1293 1294 1298 1438 1437 1295 1296 1297 1300 1301 1439
+ 1440 1302 1299 1305 1441 1442 1303 1304 1444 1311 1443 1445 1309 1307 1308 1306 1101 1097 1091 823
+ 1081 1079 1310 1078 1084 1077 1092 1105 1076 1446 1312 1073 1086 1147 1089 1087 1098 1447 864 1085
+ 1109 1448 1313 1112 1121 1449 1329 1331 830 1318 1088 1328 1314 1321 774 1320 1315 1316 1322 1338
+ 1327 1334 1330 1333 1342 1122 1323 1113 1335 1450 1326 1120 1451 1106 1452 870 1133 1337 1083 1453
+ 1143 877 1454 1128 1340 1455 1124 1456 1343 1127 1457 1136 1344 1458 1345 1459 880 1346 1460 1462
+ 1350 1347 1160 1349 1351 1156 1461 892 1352 1463 1139 1348 1464 1465 1356 901 1354 1355 1154 1358
+ 1353 1357 1167 1466 1467 1163 1359 1146 1157 1142 1169 1360 1162 1361 1166 1468 1362 1364 1469 1363
+ 1365 1366 1367 1471 1368 1370 1369 1470 1472 1371 1372 1473 1474 1373 1475 1379 1378 1476 1375 1374
+ 1477 1478 1376 1479 1480 1481 1377 1482 1380 783
+ ICV_88 $T=0 0 0 0 $X=0 $Y=48720
X11 VGND VPWR 1381 1256 1008 1182 Do[0] 1251 1236 1382 1187 1184 1036 1025 1031 1250 1253 1245 1186 1249
+ 1189 1383 1384 943 1020 Do[1] 1028 1252 1385 1040 1386 1198 1200 931 1387 1205 1389 1388 1207 1390
+ 1391 1392 1393 1395 1211 1394 1213 1397 1399 1396 1214 1398 1218 1401 1400 1224 1402 1403 1225 1404
+ 1230 1231 1406 1229 1405 1235 1407 1408 1409 1410 1411 1240 1022 Do[8] 1244 1248 1247 1414 1254 1412
+ 1413 1415 1024 Do[9] 1262 1416 1417 1280 1267 1274 1259 1034 1279 1264 Do[10] 1418 1286 1270 1266 1283
+ 1271 1080 1422 1289 1419 1074 1291 1276 1039 Do[11] 1421 1420 1423 1425 1042 Do[12] 1424 1426 1427 1428
+ 1429 1046 Do[13] 1430 1431 1432 763 Do[14] 1433 1434 1435 1436 773 Do[15] 1437 1438 800 Do[16] 1228 1439
+ 1440 802 Do[17] 1441 1442 1444 1443 1445 813 Do[18] 1447 1446 818 Do[19] 798 1111 1314 1448 1342 1313
+ 1315 1329 1449 825 1328 Do[20] 1330 1321 1331 1334 1327 1322 1338 1320 1319 Do[26] 1323 1335 1333 1450
+ 1117 834 Do[21] 1451 1452 1106 1332 Do[24] 1336 Do[25] 1128 1453 852 Do[22] 1454 1455 1069 1456 1457 865
+ Do[23] 1121 1458 1459 1124 1462 1460 1461 1463 1464 1465 870 1466 817 1467 1127 1468 1325 Do[27] 1469
+ 1154 1339 1358 Do[28] 1470 1471 1472 1473 1474 1317 1136 Do[29] 1475 1476 1324 Do[30] 1163 1478 1360 1477
+ 1479 1480 1341 Do[31] 1481 1482 783
+ ICV_94 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
