magic
tech sky130A
magscale 1 2
timestamp 1606612150
<< error_s >>
rect 4601 2768 4659 2774
rect 4719 2768 4777 2774
rect 4837 2768 4895 2774
rect 4955 2768 5013 2774
rect 5073 2768 5131 2774
rect 5191 2768 5249 2774
rect 5309 2768 5367 2774
rect 5427 2768 5485 2774
rect 5545 2768 5603 2774
rect 5663 2768 5721 2774
rect 5781 2768 5839 2774
rect 5899 2768 5957 2774
rect 6017 2768 6075 2774
rect 6135 2768 6193 2774
rect 6253 2768 6311 2774
rect 6599 2768 6657 2774
rect 6717 2768 6775 2774
rect 6835 2768 6893 2774
rect 6953 2768 7011 2774
rect 7071 2768 7129 2774
rect 7189 2768 7247 2774
rect 7307 2768 7365 2774
rect 7425 2768 7483 2774
rect 7543 2768 7601 2774
rect 7661 2768 7719 2774
rect 7779 2768 7837 2774
rect 7897 2768 7955 2774
rect 8015 2768 8073 2774
rect 8133 2768 8191 2774
rect 8251 2768 8309 2774
rect 8597 2768 8655 2774
rect 8715 2768 8773 2774
rect 8833 2768 8891 2774
rect 8951 2768 9009 2774
rect 9069 2768 9127 2774
rect 9187 2768 9245 2774
rect 9305 2768 9363 2774
rect 9423 2768 9481 2774
rect 9541 2768 9599 2774
rect 9659 2768 9717 2774
rect 9777 2768 9835 2774
rect 9895 2768 9953 2774
rect 10013 2768 10071 2774
rect 10131 2768 10189 2774
rect 10249 2768 10307 2774
rect 4601 2734 4613 2768
rect 4719 2734 4731 2768
rect 4837 2734 4849 2768
rect 4955 2734 4967 2768
rect 5073 2734 5085 2768
rect 5191 2734 5203 2768
rect 5309 2734 5321 2768
rect 5427 2734 5439 2768
rect 5545 2734 5557 2768
rect 5663 2734 5675 2768
rect 5781 2734 5793 2768
rect 5899 2734 5911 2768
rect 6017 2734 6029 2768
rect 6135 2734 6147 2768
rect 6253 2734 6265 2768
rect 6599 2734 6611 2768
rect 6717 2734 6729 2768
rect 6835 2734 6847 2768
rect 6953 2734 6965 2768
rect 7071 2734 7083 2768
rect 7189 2734 7201 2768
rect 7307 2734 7319 2768
rect 7425 2734 7437 2768
rect 7543 2734 7555 2768
rect 7661 2734 7673 2768
rect 7779 2734 7791 2768
rect 7897 2734 7909 2768
rect 8015 2734 8027 2768
rect 8133 2734 8145 2768
rect 8251 2734 8263 2768
rect 8597 2734 8609 2768
rect 8715 2734 8727 2768
rect 8833 2734 8845 2768
rect 8951 2734 8963 2768
rect 9069 2734 9081 2768
rect 9187 2734 9199 2768
rect 9305 2734 9317 2768
rect 9423 2734 9435 2768
rect 9541 2734 9553 2768
rect 9659 2734 9671 2768
rect 9777 2734 9789 2768
rect 9895 2734 9907 2768
rect 10013 2734 10025 2768
rect 10131 2734 10143 2768
rect 10249 2734 10261 2768
rect 12547 2767 12605 2773
rect 12665 2767 12723 2773
rect 12783 2767 12841 2773
rect 12901 2767 12959 2773
rect 13019 2767 13077 2773
rect 13137 2767 13195 2773
rect 13255 2767 13313 2773
rect 13373 2767 13431 2773
rect 13491 2767 13549 2773
rect 13609 2767 13667 2773
rect 13727 2767 13785 2773
rect 13845 2767 13903 2773
rect 13963 2767 14021 2773
rect 14081 2767 14139 2773
rect 14199 2767 14257 2773
rect 14317 2767 14375 2773
rect 14435 2767 14493 2773
rect 14553 2767 14611 2773
rect 14671 2767 14729 2773
rect 14789 2767 14847 2773
rect 14907 2767 14965 2773
rect 15025 2767 15083 2773
rect 15143 2767 15201 2773
rect 15261 2767 15319 2773
rect 15379 2767 15437 2773
rect 15497 2767 15555 2773
rect 15615 2767 15673 2773
rect 15733 2767 15791 2773
rect 15851 2767 15909 2773
rect 15969 2767 16027 2773
rect 16087 2767 16145 2773
rect 16205 2767 16263 2773
rect 16323 2767 16381 2773
rect 16441 2767 16499 2773
rect 16559 2767 16617 2773
rect 16677 2767 16735 2773
rect 16795 2767 16853 2773
rect 16913 2767 16971 2773
rect 17031 2767 17089 2773
rect 17149 2767 17207 2773
rect 17267 2767 17325 2773
rect 17385 2767 17443 2773
rect 17503 2767 17561 2773
rect 17621 2767 17679 2773
rect 17739 2767 17797 2773
rect 17857 2767 17915 2773
rect 17975 2767 18033 2773
rect 18093 2767 18151 2773
rect 18211 2767 18269 2773
rect 18329 2767 18387 2773
rect 18447 2767 18505 2773
rect 18565 2767 18623 2773
rect 18683 2767 18741 2773
rect 18801 2767 18859 2773
rect 18919 2767 18977 2773
rect 19037 2767 19095 2773
rect 19155 2767 19213 2773
rect 19273 2767 19331 2773
rect 19391 2767 19449 2773
rect 19509 2767 19567 2773
rect 19627 2767 19685 2773
rect 19745 2767 19803 2773
rect 19863 2767 19921 2773
rect 19981 2767 20039 2773
rect 20099 2767 20157 2773
rect 20217 2767 20275 2773
rect 20335 2767 20393 2773
rect 20453 2767 20511 2773
rect 20571 2767 20629 2773
rect 20689 2767 20747 2773
rect 20807 2767 20865 2773
rect 20925 2767 20983 2773
rect 21043 2767 21101 2773
rect 21161 2767 21219 2773
rect 21279 2767 21337 2773
rect 4601 2728 4659 2734
rect 4719 2728 4777 2734
rect 4837 2728 4895 2734
rect 4955 2728 5013 2734
rect 5073 2728 5131 2734
rect 5191 2728 5249 2734
rect 5309 2728 5367 2734
rect 5427 2728 5485 2734
rect 5545 2728 5603 2734
rect 5663 2728 5721 2734
rect 5781 2728 5839 2734
rect 5899 2728 5957 2734
rect 6017 2728 6075 2734
rect 6135 2728 6193 2734
rect 6253 2728 6311 2734
rect 6599 2728 6657 2734
rect 6717 2728 6775 2734
rect 6835 2728 6893 2734
rect 6953 2728 7011 2734
rect 7071 2728 7129 2734
rect 7189 2728 7247 2734
rect 7307 2728 7365 2734
rect 7425 2728 7483 2734
rect 7543 2728 7601 2734
rect 7661 2728 7719 2734
rect 7779 2728 7837 2734
rect 7897 2728 7955 2734
rect 8015 2728 8073 2734
rect 8133 2728 8191 2734
rect 8251 2728 8309 2734
rect 8597 2728 8655 2734
rect 8715 2728 8773 2734
rect 8833 2728 8891 2734
rect 8951 2728 9009 2734
rect 9069 2728 9127 2734
rect 9187 2728 9245 2734
rect 9305 2728 9363 2734
rect 9423 2728 9481 2734
rect 9541 2728 9599 2734
rect 9659 2728 9717 2734
rect 9777 2728 9835 2734
rect 9895 2728 9953 2734
rect 10013 2728 10071 2734
rect 10131 2728 10189 2734
rect 10249 2728 10307 2734
rect 12547 2733 12559 2767
rect 12665 2733 12677 2767
rect 12783 2733 12795 2767
rect 12901 2733 12913 2767
rect 13019 2733 13031 2767
rect 13137 2733 13149 2767
rect 13255 2733 13267 2767
rect 13373 2733 13385 2767
rect 13491 2733 13503 2767
rect 13609 2733 13621 2767
rect 13727 2733 13739 2767
rect 13845 2733 13857 2767
rect 13963 2733 13975 2767
rect 14081 2733 14093 2767
rect 14199 2733 14211 2767
rect 14317 2733 14329 2767
rect 14435 2733 14447 2767
rect 14553 2733 14565 2767
rect 14671 2733 14683 2767
rect 14789 2733 14801 2767
rect 14907 2733 14919 2767
rect 15025 2733 15037 2767
rect 15143 2733 15155 2767
rect 15261 2733 15273 2767
rect 15379 2733 15391 2767
rect 15497 2733 15509 2767
rect 15615 2733 15627 2767
rect 15733 2733 15745 2767
rect 15851 2733 15863 2767
rect 15969 2733 15981 2767
rect 16087 2733 16099 2767
rect 16205 2733 16217 2767
rect 16323 2733 16335 2767
rect 16441 2733 16453 2767
rect 16559 2733 16571 2767
rect 16677 2733 16689 2767
rect 16795 2733 16807 2767
rect 16913 2733 16925 2767
rect 17031 2733 17043 2767
rect 17149 2733 17161 2767
rect 17267 2733 17279 2767
rect 17385 2733 17397 2767
rect 17503 2733 17515 2767
rect 17621 2733 17633 2767
rect 17739 2733 17751 2767
rect 17857 2733 17869 2767
rect 17975 2733 17987 2767
rect 18093 2733 18105 2767
rect 18211 2733 18223 2767
rect 18329 2733 18341 2767
rect 18447 2733 18459 2767
rect 18565 2733 18577 2767
rect 18683 2733 18695 2767
rect 18801 2733 18813 2767
rect 18919 2733 18931 2767
rect 19037 2733 19049 2767
rect 19155 2733 19167 2767
rect 19273 2733 19285 2767
rect 19391 2733 19403 2767
rect 19509 2733 19521 2767
rect 19627 2733 19639 2767
rect 19745 2733 19757 2767
rect 19863 2733 19875 2767
rect 19981 2733 19993 2767
rect 20099 2733 20111 2767
rect 20217 2733 20229 2767
rect 20335 2733 20347 2767
rect 20453 2733 20465 2767
rect 20571 2733 20583 2767
rect 20689 2733 20701 2767
rect 20807 2733 20819 2767
rect 20925 2733 20937 2767
rect 21043 2733 21055 2767
rect 21161 2733 21173 2767
rect 21279 2733 21291 2767
rect 12547 2727 12605 2733
rect 12665 2727 12723 2733
rect 12783 2727 12841 2733
rect 12901 2727 12959 2733
rect 13019 2727 13077 2733
rect 13137 2727 13195 2733
rect 13255 2727 13313 2733
rect 13373 2727 13431 2733
rect 13491 2727 13549 2733
rect 13609 2727 13667 2733
rect 13727 2727 13785 2733
rect 13845 2727 13903 2733
rect 13963 2727 14021 2733
rect 14081 2727 14139 2733
rect 14199 2727 14257 2733
rect 14317 2727 14375 2733
rect 14435 2727 14493 2733
rect 14553 2727 14611 2733
rect 14671 2727 14729 2733
rect 14789 2727 14847 2733
rect 14907 2727 14965 2733
rect 15025 2727 15083 2733
rect 15143 2727 15201 2733
rect 15261 2727 15319 2733
rect 15379 2727 15437 2733
rect 15497 2727 15555 2733
rect 15615 2727 15673 2733
rect 15733 2727 15791 2733
rect 15851 2727 15909 2733
rect 15969 2727 16027 2733
rect 16087 2727 16145 2733
rect 16205 2727 16263 2733
rect 16323 2727 16381 2733
rect 16441 2727 16499 2733
rect 16559 2727 16617 2733
rect 16677 2727 16735 2733
rect 16795 2727 16853 2733
rect 16913 2727 16971 2733
rect 17031 2727 17089 2733
rect 17149 2727 17207 2733
rect 17267 2727 17325 2733
rect 17385 2727 17443 2733
rect 17503 2727 17561 2733
rect 17621 2727 17679 2733
rect 17739 2727 17797 2733
rect 17857 2727 17915 2733
rect 17975 2727 18033 2733
rect 18093 2727 18151 2733
rect 18211 2727 18269 2733
rect 18329 2727 18387 2733
rect 18447 2727 18505 2733
rect 18565 2727 18623 2733
rect 18683 2727 18741 2733
rect 18801 2727 18859 2733
rect 18919 2727 18977 2733
rect 19037 2727 19095 2733
rect 19155 2727 19213 2733
rect 19273 2727 19331 2733
rect 19391 2727 19449 2733
rect 19509 2727 19567 2733
rect 19627 2727 19685 2733
rect 19745 2727 19803 2733
rect 19863 2727 19921 2733
rect 19981 2727 20039 2733
rect 20099 2727 20157 2733
rect 20217 2727 20275 2733
rect 20335 2727 20393 2733
rect 20453 2727 20511 2733
rect 20571 2727 20629 2733
rect 20689 2727 20747 2733
rect 20807 2727 20865 2733
rect 20925 2727 20983 2733
rect 21043 2727 21101 2733
rect 21161 2727 21219 2733
rect 21279 2727 21337 2733
rect 6530 2077 6582 2082
rect 6766 2077 6818 2082
rect 6502 2049 6610 2054
rect 6738 2049 6846 2054
rect 12547 1203 12605 1209
rect 12665 1203 12723 1209
rect 12783 1203 12841 1209
rect 12901 1203 12959 1209
rect 13019 1203 13077 1209
rect 13137 1203 13195 1209
rect 13255 1203 13313 1209
rect 13373 1203 13431 1209
rect 13491 1203 13549 1209
rect 13609 1203 13667 1209
rect 13727 1203 13785 1209
rect 13845 1203 13903 1209
rect 13963 1203 14021 1209
rect 14081 1203 14139 1209
rect 14199 1203 14257 1209
rect 14317 1203 14375 1209
rect 14435 1203 14493 1209
rect 14553 1203 14611 1209
rect 14671 1203 14729 1209
rect 14789 1203 14847 1209
rect 14907 1203 14965 1209
rect 15025 1203 15083 1209
rect 15143 1203 15201 1209
rect 15261 1203 15319 1209
rect 15379 1203 15437 1209
rect 15497 1203 15555 1209
rect 15615 1203 15673 1209
rect 15733 1203 15791 1209
rect 15851 1203 15909 1209
rect 15969 1203 16027 1209
rect 16087 1203 16145 1209
rect 16205 1203 16263 1209
rect 16323 1203 16381 1209
rect 16441 1203 16499 1209
rect 16559 1203 16617 1209
rect 16677 1203 16735 1209
rect 16795 1203 16853 1209
rect 16913 1203 16971 1209
rect 17031 1203 17089 1209
rect 17149 1203 17207 1209
rect 17267 1203 17325 1209
rect 17385 1203 17443 1209
rect 17503 1203 17561 1209
rect 17621 1203 17679 1209
rect 17739 1203 17797 1209
rect 17857 1203 17915 1209
rect 17975 1203 18033 1209
rect 18093 1203 18151 1209
rect 18211 1203 18269 1209
rect 18329 1203 18387 1209
rect 18447 1203 18505 1209
rect 18565 1203 18623 1209
rect 18683 1203 18741 1209
rect 18801 1203 18859 1209
rect 18919 1203 18977 1209
rect 19037 1203 19095 1209
rect 19155 1203 19213 1209
rect 19273 1203 19331 1209
rect 19391 1203 19449 1209
rect 19509 1203 19567 1209
rect 19627 1203 19685 1209
rect 19745 1203 19803 1209
rect 19863 1203 19921 1209
rect 19981 1203 20039 1209
rect 20099 1203 20157 1209
rect 20217 1203 20275 1209
rect 20335 1203 20393 1209
rect 20453 1203 20511 1209
rect 20571 1203 20629 1209
rect 20689 1203 20747 1209
rect 20807 1203 20865 1209
rect 20925 1203 20983 1209
rect 21043 1203 21101 1209
rect 21161 1203 21219 1209
rect 21279 1203 21337 1209
rect 12547 1169 12559 1203
rect 12665 1169 12677 1203
rect 12783 1169 12795 1203
rect 12901 1169 12913 1203
rect 13019 1169 13031 1203
rect 13137 1169 13149 1203
rect 13255 1169 13267 1203
rect 13373 1169 13385 1203
rect 13491 1169 13503 1203
rect 13609 1169 13621 1203
rect 13727 1169 13739 1203
rect 13845 1169 13857 1203
rect 13963 1169 13975 1203
rect 14081 1169 14093 1203
rect 14199 1169 14211 1203
rect 14317 1169 14329 1203
rect 14435 1169 14447 1203
rect 14553 1169 14565 1203
rect 14671 1169 14683 1203
rect 14789 1169 14801 1203
rect 14907 1169 14919 1203
rect 15025 1169 15037 1203
rect 15143 1169 15155 1203
rect 15261 1169 15273 1203
rect 15379 1169 15391 1203
rect 15497 1169 15509 1203
rect 15615 1169 15627 1203
rect 15733 1169 15745 1203
rect 15851 1169 15863 1203
rect 15969 1169 15981 1203
rect 16087 1169 16099 1203
rect 16205 1169 16217 1203
rect 16323 1169 16335 1203
rect 16441 1169 16453 1203
rect 16559 1169 16571 1203
rect 16677 1169 16689 1203
rect 16795 1169 16807 1203
rect 16913 1169 16925 1203
rect 17031 1169 17043 1203
rect 17149 1169 17161 1203
rect 17267 1169 17279 1203
rect 17385 1169 17397 1203
rect 17503 1169 17515 1203
rect 17621 1169 17633 1203
rect 17739 1169 17751 1203
rect 17857 1169 17869 1203
rect 17975 1169 17987 1203
rect 18093 1169 18105 1203
rect 18211 1169 18223 1203
rect 18329 1169 18341 1203
rect 18447 1169 18459 1203
rect 18565 1169 18577 1203
rect 18683 1169 18695 1203
rect 18801 1169 18813 1203
rect 18919 1169 18931 1203
rect 19037 1169 19049 1203
rect 19155 1169 19167 1203
rect 19273 1169 19285 1203
rect 19391 1169 19403 1203
rect 19509 1169 19521 1203
rect 19627 1169 19639 1203
rect 19745 1169 19757 1203
rect 19863 1169 19875 1203
rect 19981 1169 19993 1203
rect 20099 1169 20111 1203
rect 20217 1169 20229 1203
rect 20335 1169 20347 1203
rect 20453 1169 20465 1203
rect 20571 1169 20583 1203
rect 20689 1169 20701 1203
rect 20807 1169 20819 1203
rect 20925 1169 20937 1203
rect 21043 1169 21055 1203
rect 21161 1169 21173 1203
rect 21279 1169 21291 1203
rect 12547 1163 12605 1169
rect 12665 1163 12723 1169
rect 12783 1163 12841 1169
rect 12901 1163 12959 1169
rect 13019 1163 13077 1169
rect 13137 1163 13195 1169
rect 13255 1163 13313 1169
rect 13373 1163 13431 1169
rect 13491 1163 13549 1169
rect 13609 1163 13667 1169
rect 13727 1163 13785 1169
rect 13845 1163 13903 1169
rect 13963 1163 14021 1169
rect 14081 1163 14139 1169
rect 14199 1163 14257 1169
rect 14317 1163 14375 1169
rect 14435 1163 14493 1169
rect 14553 1163 14611 1169
rect 14671 1163 14729 1169
rect 14789 1163 14847 1169
rect 14907 1163 14965 1169
rect 15025 1163 15083 1169
rect 15143 1163 15201 1169
rect 15261 1163 15319 1169
rect 15379 1163 15437 1169
rect 15497 1163 15555 1169
rect 15615 1163 15673 1169
rect 15733 1163 15791 1169
rect 15851 1163 15909 1169
rect 15969 1163 16027 1169
rect 16087 1163 16145 1169
rect 16205 1163 16263 1169
rect 16323 1163 16381 1169
rect 16441 1163 16499 1169
rect 16559 1163 16617 1169
rect 16677 1163 16735 1169
rect 16795 1163 16853 1169
rect 16913 1163 16971 1169
rect 17031 1163 17089 1169
rect 17149 1163 17207 1169
rect 17267 1163 17325 1169
rect 17385 1163 17443 1169
rect 17503 1163 17561 1169
rect 17621 1163 17679 1169
rect 17739 1163 17797 1169
rect 17857 1163 17915 1169
rect 17975 1163 18033 1169
rect 18093 1163 18151 1169
rect 18211 1163 18269 1169
rect 18329 1163 18387 1169
rect 18447 1163 18505 1169
rect 18565 1163 18623 1169
rect 18683 1163 18741 1169
rect 18801 1163 18859 1169
rect 18919 1163 18977 1169
rect 19037 1163 19095 1169
rect 19155 1163 19213 1169
rect 19273 1163 19331 1169
rect 19391 1163 19449 1169
rect 19509 1163 19567 1169
rect 19627 1163 19685 1169
rect 19745 1163 19803 1169
rect 19863 1163 19921 1169
rect 19981 1163 20039 1169
rect 20099 1163 20157 1169
rect 20217 1163 20275 1169
rect 20335 1163 20393 1169
rect 20453 1163 20511 1169
rect 20571 1163 20629 1169
rect 20689 1163 20747 1169
rect 20807 1163 20865 1169
rect 20925 1163 20983 1169
rect 21043 1163 21101 1169
rect 21161 1163 21219 1169
rect 21279 1163 21337 1169
rect 1337 580 1395 586
rect 1455 580 1513 586
rect 1573 580 1631 586
rect 1691 580 1749 586
rect 1809 580 1867 586
rect 1927 580 1985 586
rect 2045 580 2103 586
rect 2163 580 2221 586
rect 2281 580 2339 586
rect 2399 580 2457 586
rect 2517 580 2575 586
rect 2635 580 2693 586
rect 2753 580 2811 586
rect 2871 580 2929 586
rect 2989 580 3047 586
rect 3107 580 3165 586
rect 3225 580 3283 586
rect 3343 580 3401 586
rect 3461 580 3519 586
rect 3579 580 3637 586
rect 3697 580 3755 586
rect 3815 580 3873 586
rect 3933 580 3991 586
rect 4051 580 4109 586
rect 4169 580 4227 586
rect 4287 580 4345 586
rect 4405 580 4463 586
rect 4523 580 4581 586
rect 4641 580 4699 586
rect 4759 580 4817 586
rect 4877 580 4935 586
rect 4995 580 5053 586
rect 5113 580 5171 586
rect 5231 580 5289 586
rect 5349 580 5407 586
rect 5467 580 5525 586
rect 5585 580 5643 586
rect 5703 580 5761 586
rect 5821 580 5879 586
rect 5939 580 5997 586
rect 6057 580 6115 586
rect 6175 580 6233 586
rect 6293 580 6351 586
rect 6411 580 6469 586
rect 6529 580 6587 586
rect 6647 580 6705 586
rect 6765 580 6823 586
rect 6883 580 6941 586
rect 7001 580 7059 586
rect 7119 580 7177 586
rect 1337 546 1349 580
rect 1455 546 1467 580
rect 1573 546 1585 580
rect 1691 546 1703 580
rect 1809 546 1821 580
rect 1927 546 1939 580
rect 2045 546 2057 580
rect 2163 546 2175 580
rect 2281 546 2293 580
rect 2399 546 2411 580
rect 2517 546 2529 580
rect 2635 546 2647 580
rect 2753 546 2765 580
rect 2871 546 2883 580
rect 2989 546 3001 580
rect 3107 546 3119 580
rect 3225 546 3237 580
rect 3343 546 3355 580
rect 3461 546 3473 580
rect 3579 546 3591 580
rect 3697 546 3709 580
rect 3815 546 3827 580
rect 3933 546 3945 580
rect 4051 546 4063 580
rect 4169 546 4181 580
rect 4287 546 4299 580
rect 4405 546 4417 580
rect 4523 546 4535 580
rect 4641 546 4653 580
rect 4759 546 4771 580
rect 4877 546 4889 580
rect 4995 546 5007 580
rect 5113 546 5125 580
rect 5231 546 5243 580
rect 5349 546 5361 580
rect 5467 546 5479 580
rect 5585 546 5597 580
rect 5703 546 5715 580
rect 5821 546 5833 580
rect 5939 546 5951 580
rect 6057 546 6069 580
rect 6175 546 6187 580
rect 6293 546 6305 580
rect 6411 546 6423 580
rect 6529 546 6541 580
rect 6647 546 6659 580
rect 6765 546 6777 580
rect 6883 546 6895 580
rect 7001 546 7013 580
rect 7119 546 7131 580
rect 1337 540 1395 546
rect 1455 540 1513 546
rect 1573 540 1631 546
rect 1691 540 1749 546
rect 1809 540 1867 546
rect 1927 540 1985 546
rect 2045 540 2103 546
rect 2163 540 2221 546
rect 2281 540 2339 546
rect 2399 540 2457 546
rect 2517 540 2575 546
rect 2635 540 2693 546
rect 2753 540 2811 546
rect 2871 540 2929 546
rect 2989 540 3047 546
rect 3107 540 3165 546
rect 3225 540 3283 546
rect 3343 540 3401 546
rect 3461 540 3519 546
rect 3579 540 3637 546
rect 3697 540 3755 546
rect 3815 540 3873 546
rect 3933 540 3991 546
rect 4051 540 4109 546
rect 4169 540 4227 546
rect 4287 540 4345 546
rect 4405 540 4463 546
rect 4523 540 4581 546
rect 4641 540 4699 546
rect 4759 540 4817 546
rect 4877 540 4935 546
rect 4995 540 5053 546
rect 5113 540 5171 546
rect 5231 540 5289 546
rect 5349 540 5407 546
rect 5467 540 5525 546
rect 5585 540 5643 546
rect 5703 540 5761 546
rect 5821 540 5879 546
rect 5939 540 5997 546
rect 6057 540 6115 546
rect 6175 540 6233 546
rect 6293 540 6351 546
rect 6411 540 6469 546
rect 6529 540 6587 546
rect 6647 540 6705 546
rect 6765 540 6823 546
rect 6883 540 6941 546
rect 7001 540 7059 546
rect 7119 540 7177 546
rect 7607 -165 7626 -149
rect 7725 -165 7744 -149
rect 7591 -181 7642 -165
rect 7709 -181 7760 -165
rect 7607 -183 7641 -181
rect 7725 -183 7759 -181
rect 7591 -199 7642 -183
rect 7709 -199 7760 -183
rect 7607 -215 7626 -199
rect 7725 -215 7744 -199
rect 7607 -273 7626 -257
rect 7725 -273 7744 -257
rect 7591 -289 7642 -273
rect 7709 -289 7760 -273
rect 7607 -291 7641 -289
rect 7725 -291 7759 -289
rect 7591 -307 7642 -291
rect 7709 -307 7760 -291
rect 7607 -323 7626 -307
rect 7725 -323 7744 -307
rect 1337 -984 1395 -978
rect 1455 -984 1513 -978
rect 1573 -984 1631 -978
rect 1691 -984 1749 -978
rect 1809 -984 1867 -978
rect 1927 -984 1985 -978
rect 2045 -984 2103 -978
rect 2163 -984 2221 -978
rect 2281 -984 2339 -978
rect 2399 -984 2457 -978
rect 2517 -984 2575 -978
rect 2635 -984 2693 -978
rect 2753 -984 2811 -978
rect 2871 -984 2929 -978
rect 2989 -984 3047 -978
rect 3107 -984 3165 -978
rect 3225 -984 3283 -978
rect 3343 -984 3401 -978
rect 3461 -984 3519 -978
rect 3579 -984 3637 -978
rect 3697 -984 3755 -978
rect 3815 -984 3873 -978
rect 3933 -984 3991 -978
rect 4051 -984 4109 -978
rect 4169 -984 4227 -978
rect 4287 -984 4345 -978
rect 4405 -984 4463 -978
rect 4523 -984 4581 -978
rect 4641 -984 4699 -978
rect 4759 -984 4817 -978
rect 4877 -984 4935 -978
rect 4995 -984 5053 -978
rect 5113 -984 5171 -978
rect 5231 -984 5289 -978
rect 5349 -984 5407 -978
rect 5467 -984 5525 -978
rect 5585 -984 5643 -978
rect 5703 -984 5761 -978
rect 5821 -984 5879 -978
rect 5939 -984 5997 -978
rect 6057 -984 6115 -978
rect 6175 -984 6233 -978
rect 6293 -984 6351 -978
rect 6411 -984 6469 -978
rect 6529 -984 6587 -978
rect 6647 -984 6705 -978
rect 6765 -984 6823 -978
rect 6883 -984 6941 -978
rect 7001 -984 7059 -978
rect 7119 -984 7177 -978
rect 1337 -1018 1349 -984
rect 1455 -1018 1467 -984
rect 1573 -1018 1585 -984
rect 1691 -1018 1703 -984
rect 1809 -1018 1821 -984
rect 1927 -1018 1939 -984
rect 2045 -1018 2057 -984
rect 2163 -1018 2175 -984
rect 2281 -1018 2293 -984
rect 2399 -1018 2411 -984
rect 2517 -1018 2529 -984
rect 2635 -1018 2647 -984
rect 2753 -1018 2765 -984
rect 2871 -1018 2883 -984
rect 2989 -1018 3001 -984
rect 3107 -1018 3119 -984
rect 3225 -1018 3237 -984
rect 3343 -1018 3355 -984
rect 3461 -1018 3473 -984
rect 3579 -1018 3591 -984
rect 3697 -1018 3709 -984
rect 3815 -1018 3827 -984
rect 3933 -1018 3945 -984
rect 4051 -1018 4063 -984
rect 4169 -1018 4181 -984
rect 4287 -1018 4299 -984
rect 4405 -1018 4417 -984
rect 4523 -1018 4535 -984
rect 4641 -1018 4653 -984
rect 4759 -1018 4771 -984
rect 4877 -1018 4889 -984
rect 4995 -1018 5007 -984
rect 5113 -1018 5125 -984
rect 5231 -1018 5243 -984
rect 5349 -1018 5361 -984
rect 5467 -1018 5479 -984
rect 5585 -1018 5597 -984
rect 5703 -1018 5715 -984
rect 5821 -1018 5833 -984
rect 5939 -1018 5951 -984
rect 6057 -1018 6069 -984
rect 6175 -1018 6187 -984
rect 6293 -1018 6305 -984
rect 6411 -1018 6423 -984
rect 6529 -1018 6541 -984
rect 6647 -1018 6659 -984
rect 6765 -1018 6777 -984
rect 6883 -1018 6895 -984
rect 7001 -1018 7013 -984
rect 7119 -1018 7131 -984
rect 1337 -1024 1395 -1018
rect 1455 -1024 1513 -1018
rect 1573 -1024 1631 -1018
rect 1691 -1024 1749 -1018
rect 1809 -1024 1867 -1018
rect 1927 -1024 1985 -1018
rect 2045 -1024 2103 -1018
rect 2163 -1024 2221 -1018
rect 2281 -1024 2339 -1018
rect 2399 -1024 2457 -1018
rect 2517 -1024 2575 -1018
rect 2635 -1024 2693 -1018
rect 2753 -1024 2811 -1018
rect 2871 -1024 2929 -1018
rect 2989 -1024 3047 -1018
rect 3107 -1024 3165 -1018
rect 3225 -1024 3283 -1018
rect 3343 -1024 3401 -1018
rect 3461 -1024 3519 -1018
rect 3579 -1024 3637 -1018
rect 3697 -1024 3755 -1018
rect 3815 -1024 3873 -1018
rect 3933 -1024 3991 -1018
rect 4051 -1024 4109 -1018
rect 4169 -1024 4227 -1018
rect 4287 -1024 4345 -1018
rect 4405 -1024 4463 -1018
rect 4523 -1024 4581 -1018
rect 4641 -1024 4699 -1018
rect 4759 -1024 4817 -1018
rect 4877 -1024 4935 -1018
rect 4995 -1024 5053 -1018
rect 5113 -1024 5171 -1018
rect 5231 -1024 5289 -1018
rect 5349 -1024 5407 -1018
rect 5467 -1024 5525 -1018
rect 5585 -1024 5643 -1018
rect 5703 -1024 5761 -1018
rect 5821 -1024 5879 -1018
rect 5939 -1024 5997 -1018
rect 6057 -1024 6115 -1018
rect 6175 -1024 6233 -1018
rect 6293 -1024 6351 -1018
rect 6411 -1024 6469 -1018
rect 6529 -1024 6587 -1018
rect 6647 -1024 6705 -1018
rect 6765 -1024 6823 -1018
rect 6883 -1024 6941 -1018
rect 7001 -1024 7059 -1018
rect 7119 -1024 7177 -1018
rect 1337 -1188 1395 -1182
rect 1455 -1188 1513 -1182
rect 1573 -1188 1631 -1182
rect 1691 -1188 1749 -1182
rect 1809 -1188 1867 -1182
rect 1927 -1188 1985 -1182
rect 2045 -1188 2103 -1182
rect 2163 -1188 2221 -1182
rect 2281 -1188 2339 -1182
rect 2399 -1188 2457 -1182
rect 2517 -1188 2575 -1182
rect 2635 -1188 2693 -1182
rect 2753 -1188 2811 -1182
rect 2871 -1188 2929 -1182
rect 2989 -1188 3047 -1182
rect 3107 -1188 3165 -1182
rect 3225 -1188 3283 -1182
rect 3343 -1188 3401 -1182
rect 3461 -1188 3519 -1182
rect 3579 -1188 3637 -1182
rect 3697 -1188 3755 -1182
rect 3815 -1188 3873 -1182
rect 3933 -1188 3991 -1182
rect 4051 -1188 4109 -1182
rect 4169 -1188 4227 -1182
rect 4287 -1188 4345 -1182
rect 4405 -1188 4463 -1182
rect 4523 -1188 4581 -1182
rect 4641 -1188 4699 -1182
rect 4759 -1188 4817 -1182
rect 4877 -1188 4935 -1182
rect 4995 -1188 5053 -1182
rect 5113 -1188 5171 -1182
rect 5231 -1188 5289 -1182
rect 5349 -1188 5407 -1182
rect 5467 -1188 5525 -1182
rect 5585 -1188 5643 -1182
rect 5703 -1188 5761 -1182
rect 5821 -1188 5879 -1182
rect 5939 -1188 5997 -1182
rect 6057 -1188 6115 -1182
rect 6175 -1188 6233 -1182
rect 6293 -1188 6351 -1182
rect 6411 -1188 6469 -1182
rect 6529 -1188 6587 -1182
rect 6647 -1188 6705 -1182
rect 6765 -1188 6823 -1182
rect 6883 -1188 6941 -1182
rect 7001 -1188 7059 -1182
rect 7119 -1188 7177 -1182
rect 1337 -1222 1349 -1188
rect 1455 -1222 1467 -1188
rect 1573 -1222 1585 -1188
rect 1691 -1222 1703 -1188
rect 1809 -1222 1821 -1188
rect 1927 -1222 1939 -1188
rect 2045 -1222 2057 -1188
rect 2163 -1222 2175 -1188
rect 2281 -1222 2293 -1188
rect 2399 -1222 2411 -1188
rect 2517 -1222 2529 -1188
rect 2635 -1222 2647 -1188
rect 2753 -1222 2765 -1188
rect 2871 -1222 2883 -1188
rect 2989 -1222 3001 -1188
rect 3107 -1222 3119 -1188
rect 3225 -1222 3237 -1188
rect 3343 -1222 3355 -1188
rect 3461 -1222 3473 -1188
rect 3579 -1222 3591 -1188
rect 3697 -1222 3709 -1188
rect 3815 -1222 3827 -1188
rect 3933 -1222 3945 -1188
rect 4051 -1222 4063 -1188
rect 4169 -1222 4181 -1188
rect 4287 -1222 4299 -1188
rect 4405 -1222 4417 -1188
rect 4523 -1222 4535 -1188
rect 4641 -1222 4653 -1188
rect 4759 -1222 4771 -1188
rect 4877 -1222 4889 -1188
rect 4995 -1222 5007 -1188
rect 5113 -1222 5125 -1188
rect 5231 -1222 5243 -1188
rect 5349 -1222 5361 -1188
rect 5467 -1222 5479 -1188
rect 5585 -1222 5597 -1188
rect 5703 -1222 5715 -1188
rect 5821 -1222 5833 -1188
rect 5939 -1222 5951 -1188
rect 6057 -1222 6069 -1188
rect 6175 -1222 6187 -1188
rect 6293 -1222 6305 -1188
rect 6411 -1222 6423 -1188
rect 6529 -1222 6541 -1188
rect 6647 -1222 6659 -1188
rect 6765 -1222 6777 -1188
rect 6883 -1222 6895 -1188
rect 7001 -1222 7013 -1188
rect 7119 -1222 7131 -1188
rect 1337 -1228 1395 -1222
rect 1455 -1228 1513 -1222
rect 1573 -1228 1631 -1222
rect 1691 -1228 1749 -1222
rect 1809 -1228 1867 -1222
rect 1927 -1228 1985 -1222
rect 2045 -1228 2103 -1222
rect 2163 -1228 2221 -1222
rect 2281 -1228 2339 -1222
rect 2399 -1228 2457 -1222
rect 2517 -1228 2575 -1222
rect 2635 -1228 2693 -1222
rect 2753 -1228 2811 -1222
rect 2871 -1228 2929 -1222
rect 2989 -1228 3047 -1222
rect 3107 -1228 3165 -1222
rect 3225 -1228 3283 -1222
rect 3343 -1228 3401 -1222
rect 3461 -1228 3519 -1222
rect 3579 -1228 3637 -1222
rect 3697 -1228 3755 -1222
rect 3815 -1228 3873 -1222
rect 3933 -1228 3991 -1222
rect 4051 -1228 4109 -1222
rect 4169 -1228 4227 -1222
rect 4287 -1228 4345 -1222
rect 4405 -1228 4463 -1222
rect 4523 -1228 4581 -1222
rect 4641 -1228 4699 -1222
rect 4759 -1228 4817 -1222
rect 4877 -1228 4935 -1222
rect 4995 -1228 5053 -1222
rect 5113 -1228 5171 -1222
rect 5231 -1228 5289 -1222
rect 5349 -1228 5407 -1222
rect 5467 -1228 5525 -1222
rect 5585 -1228 5643 -1222
rect 5703 -1228 5761 -1222
rect 5821 -1228 5879 -1222
rect 5939 -1228 5997 -1222
rect 6057 -1228 6115 -1222
rect 6175 -1228 6233 -1222
rect 6293 -1228 6351 -1222
rect 6411 -1228 6469 -1222
rect 6529 -1228 6587 -1222
rect 6647 -1228 6705 -1222
rect 6765 -1228 6823 -1222
rect 6883 -1228 6941 -1222
rect 7001 -1228 7059 -1222
rect 7119 -1228 7177 -1222
rect 1337 -2752 1395 -2746
rect 1455 -2752 1513 -2746
rect 1573 -2752 1631 -2746
rect 1691 -2752 1749 -2746
rect 1809 -2752 1867 -2746
rect 1927 -2752 1985 -2746
rect 2045 -2752 2103 -2746
rect 2163 -2752 2221 -2746
rect 2281 -2752 2339 -2746
rect 2399 -2752 2457 -2746
rect 2517 -2752 2575 -2746
rect 2635 -2752 2693 -2746
rect 2753 -2752 2811 -2746
rect 2871 -2752 2929 -2746
rect 2989 -2752 3047 -2746
rect 3107 -2752 3165 -2746
rect 3225 -2752 3283 -2746
rect 3343 -2752 3401 -2746
rect 3461 -2752 3519 -2746
rect 3579 -2752 3637 -2746
rect 3697 -2752 3755 -2746
rect 3815 -2752 3873 -2746
rect 3933 -2752 3991 -2746
rect 4051 -2752 4109 -2746
rect 4169 -2752 4227 -2746
rect 4287 -2752 4345 -2746
rect 4405 -2752 4463 -2746
rect 4523 -2752 4581 -2746
rect 4641 -2752 4699 -2746
rect 4759 -2752 4817 -2746
rect 4877 -2752 4935 -2746
rect 4995 -2752 5053 -2746
rect 5113 -2752 5171 -2746
rect 5231 -2752 5289 -2746
rect 5349 -2752 5407 -2746
rect 5467 -2752 5525 -2746
rect 5585 -2752 5643 -2746
rect 5703 -2752 5761 -2746
rect 5821 -2752 5879 -2746
rect 5939 -2752 5997 -2746
rect 6057 -2752 6115 -2746
rect 6175 -2752 6233 -2746
rect 6293 -2752 6351 -2746
rect 6411 -2752 6469 -2746
rect 6529 -2752 6587 -2746
rect 6647 -2752 6705 -2746
rect 6765 -2752 6823 -2746
rect 6883 -2752 6941 -2746
rect 7001 -2752 7059 -2746
rect 7119 -2752 7177 -2746
rect 1337 -2786 1349 -2752
rect 1455 -2786 1467 -2752
rect 1573 -2786 1585 -2752
rect 1691 -2786 1703 -2752
rect 1809 -2786 1821 -2752
rect 1927 -2786 1939 -2752
rect 2045 -2786 2057 -2752
rect 2163 -2786 2175 -2752
rect 2281 -2786 2293 -2752
rect 2399 -2786 2411 -2752
rect 2517 -2786 2529 -2752
rect 2635 -2786 2647 -2752
rect 2753 -2786 2765 -2752
rect 2871 -2786 2883 -2752
rect 2989 -2786 3001 -2752
rect 3107 -2786 3119 -2752
rect 3225 -2786 3237 -2752
rect 3343 -2786 3355 -2752
rect 3461 -2786 3473 -2752
rect 3579 -2786 3591 -2752
rect 3697 -2786 3709 -2752
rect 3815 -2786 3827 -2752
rect 3933 -2786 3945 -2752
rect 4051 -2786 4063 -2752
rect 4169 -2786 4181 -2752
rect 4287 -2786 4299 -2752
rect 4405 -2786 4417 -2752
rect 4523 -2786 4535 -2752
rect 4641 -2786 4653 -2752
rect 4759 -2786 4771 -2752
rect 4877 -2786 4889 -2752
rect 4995 -2786 5007 -2752
rect 5113 -2786 5125 -2752
rect 5231 -2786 5243 -2752
rect 5349 -2786 5361 -2752
rect 5467 -2786 5479 -2752
rect 5585 -2786 5597 -2752
rect 5703 -2786 5715 -2752
rect 5821 -2786 5833 -2752
rect 5939 -2786 5951 -2752
rect 6057 -2786 6069 -2752
rect 6175 -2786 6187 -2752
rect 6293 -2786 6305 -2752
rect 6411 -2786 6423 -2752
rect 6529 -2786 6541 -2752
rect 6647 -2786 6659 -2752
rect 6765 -2786 6777 -2752
rect 6883 -2786 6895 -2752
rect 7001 -2786 7013 -2752
rect 7119 -2786 7131 -2752
rect 1337 -2792 1395 -2786
rect 1455 -2792 1513 -2786
rect 1573 -2792 1631 -2786
rect 1691 -2792 1749 -2786
rect 1809 -2792 1867 -2786
rect 1927 -2792 1985 -2786
rect 2045 -2792 2103 -2786
rect 2163 -2792 2221 -2786
rect 2281 -2792 2339 -2786
rect 2399 -2792 2457 -2786
rect 2517 -2792 2575 -2786
rect 2635 -2792 2693 -2786
rect 2753 -2792 2811 -2786
rect 2871 -2792 2929 -2786
rect 2989 -2792 3047 -2786
rect 3107 -2792 3165 -2786
rect 3225 -2792 3283 -2786
rect 3343 -2792 3401 -2786
rect 3461 -2792 3519 -2786
rect 3579 -2792 3637 -2786
rect 3697 -2792 3755 -2786
rect 3815 -2792 3873 -2786
rect 3933 -2792 3991 -2786
rect 4051 -2792 4109 -2786
rect 4169 -2792 4227 -2786
rect 4287 -2792 4345 -2786
rect 4405 -2792 4463 -2786
rect 4523 -2792 4581 -2786
rect 4641 -2792 4699 -2786
rect 4759 -2792 4817 -2786
rect 4877 -2792 4935 -2786
rect 4995 -2792 5053 -2786
rect 5113 -2792 5171 -2786
rect 5231 -2792 5289 -2786
rect 5349 -2792 5407 -2786
rect 5467 -2792 5525 -2786
rect 5585 -2792 5643 -2786
rect 5703 -2792 5761 -2786
rect 5821 -2792 5879 -2786
rect 5939 -2792 5997 -2786
rect 6057 -2792 6115 -2786
rect 6175 -2792 6233 -2786
rect 6293 -2792 6351 -2786
rect 6411 -2792 6469 -2786
rect 6529 -2792 6587 -2786
rect 6647 -2792 6705 -2786
rect 6765 -2792 6823 -2786
rect 6883 -2792 6941 -2786
rect 7001 -2792 7059 -2786
rect 7119 -2792 7177 -2786
rect 1337 -2956 1395 -2950
rect 1455 -2956 1513 -2950
rect 1573 -2956 1631 -2950
rect 1691 -2956 1749 -2950
rect 1809 -2956 1867 -2950
rect 1927 -2956 1985 -2950
rect 2045 -2956 2103 -2950
rect 2163 -2956 2221 -2950
rect 2281 -2956 2339 -2950
rect 2399 -2956 2457 -2950
rect 2517 -2956 2575 -2950
rect 2635 -2956 2693 -2950
rect 2753 -2956 2811 -2950
rect 2871 -2956 2929 -2950
rect 2989 -2956 3047 -2950
rect 3107 -2956 3165 -2950
rect 3225 -2956 3283 -2950
rect 3343 -2956 3401 -2950
rect 3461 -2956 3519 -2950
rect 3579 -2956 3637 -2950
rect 3697 -2956 3755 -2950
rect 3815 -2956 3873 -2950
rect 3933 -2956 3991 -2950
rect 4051 -2956 4109 -2950
rect 4169 -2956 4227 -2950
rect 4287 -2956 4345 -2950
rect 4405 -2956 4463 -2950
rect 4523 -2956 4581 -2950
rect 4641 -2956 4699 -2950
rect 4759 -2956 4817 -2950
rect 4877 -2956 4935 -2950
rect 4995 -2956 5053 -2950
rect 5113 -2956 5171 -2950
rect 5231 -2956 5289 -2950
rect 5349 -2956 5407 -2950
rect 5467 -2956 5525 -2950
rect 5585 -2956 5643 -2950
rect 5703 -2956 5761 -2950
rect 5821 -2956 5879 -2950
rect 5939 -2956 5997 -2950
rect 6057 -2956 6115 -2950
rect 6175 -2956 6233 -2950
rect 6293 -2956 6351 -2950
rect 6411 -2956 6469 -2950
rect 6529 -2956 6587 -2950
rect 6647 -2956 6705 -2950
rect 6765 -2956 6823 -2950
rect 6883 -2956 6941 -2950
rect 7001 -2956 7059 -2950
rect 7119 -2956 7177 -2950
rect 1337 -2990 1349 -2956
rect 1455 -2990 1467 -2956
rect 1573 -2990 1585 -2956
rect 1691 -2990 1703 -2956
rect 1809 -2990 1821 -2956
rect 1927 -2990 1939 -2956
rect 2045 -2990 2057 -2956
rect 2163 -2990 2175 -2956
rect 2281 -2990 2293 -2956
rect 2399 -2990 2411 -2956
rect 2517 -2990 2529 -2956
rect 2635 -2990 2647 -2956
rect 2753 -2990 2765 -2956
rect 2871 -2990 2883 -2956
rect 2989 -2990 3001 -2956
rect 3107 -2990 3119 -2956
rect 3225 -2990 3237 -2956
rect 3343 -2990 3355 -2956
rect 3461 -2990 3473 -2956
rect 3579 -2990 3591 -2956
rect 3697 -2990 3709 -2956
rect 3815 -2990 3827 -2956
rect 3933 -2990 3945 -2956
rect 4051 -2990 4063 -2956
rect 4169 -2990 4181 -2956
rect 4287 -2990 4299 -2956
rect 4405 -2990 4417 -2956
rect 4523 -2990 4535 -2956
rect 4641 -2990 4653 -2956
rect 4759 -2990 4771 -2956
rect 4877 -2990 4889 -2956
rect 4995 -2990 5007 -2956
rect 5113 -2990 5125 -2956
rect 5231 -2990 5243 -2956
rect 5349 -2990 5361 -2956
rect 5467 -2990 5479 -2956
rect 5585 -2990 5597 -2956
rect 5703 -2990 5715 -2956
rect 5821 -2990 5833 -2956
rect 5939 -2990 5951 -2956
rect 6057 -2990 6069 -2956
rect 6175 -2990 6187 -2956
rect 6293 -2990 6305 -2956
rect 6411 -2990 6423 -2956
rect 6529 -2990 6541 -2956
rect 6647 -2990 6659 -2956
rect 6765 -2990 6777 -2956
rect 6883 -2990 6895 -2956
rect 7001 -2990 7013 -2956
rect 7119 -2990 7131 -2956
rect 1337 -2996 1395 -2990
rect 1455 -2996 1513 -2990
rect 1573 -2996 1631 -2990
rect 1691 -2996 1749 -2990
rect 1809 -2996 1867 -2990
rect 1927 -2996 1985 -2990
rect 2045 -2996 2103 -2990
rect 2163 -2996 2221 -2990
rect 2281 -2996 2339 -2990
rect 2399 -2996 2457 -2990
rect 2517 -2996 2575 -2990
rect 2635 -2996 2693 -2990
rect 2753 -2996 2811 -2990
rect 2871 -2996 2929 -2990
rect 2989 -2996 3047 -2990
rect 3107 -2996 3165 -2990
rect 3225 -2996 3283 -2990
rect 3343 -2996 3401 -2990
rect 3461 -2996 3519 -2990
rect 3579 -2996 3637 -2990
rect 3697 -2996 3755 -2990
rect 3815 -2996 3873 -2990
rect 3933 -2996 3991 -2990
rect 4051 -2996 4109 -2990
rect 4169 -2996 4227 -2990
rect 4287 -2996 4345 -2990
rect 4405 -2996 4463 -2990
rect 4523 -2996 4581 -2990
rect 4641 -2996 4699 -2990
rect 4759 -2996 4817 -2990
rect 4877 -2996 4935 -2990
rect 4995 -2996 5053 -2990
rect 5113 -2996 5171 -2990
rect 5231 -2996 5289 -2990
rect 5349 -2996 5407 -2990
rect 5467 -2996 5525 -2990
rect 5585 -2996 5643 -2990
rect 5703 -2996 5761 -2990
rect 5821 -2996 5879 -2990
rect 5939 -2996 5997 -2990
rect 6057 -2996 6115 -2990
rect 6175 -2996 6233 -2990
rect 6293 -2996 6351 -2990
rect 6411 -2996 6469 -2990
rect 6529 -2996 6587 -2990
rect 6647 -2996 6705 -2990
rect 6765 -2996 6823 -2990
rect 6883 -2996 6941 -2990
rect 7001 -2996 7059 -2990
rect 7119 -2996 7177 -2990
rect 1337 -4520 1395 -4514
rect 1455 -4520 1513 -4514
rect 1573 -4520 1631 -4514
rect 1691 -4520 1749 -4514
rect 1809 -4520 1867 -4514
rect 1927 -4520 1985 -4514
rect 2045 -4520 2103 -4514
rect 2163 -4520 2221 -4514
rect 2281 -4520 2339 -4514
rect 2399 -4520 2457 -4514
rect 2517 -4520 2575 -4514
rect 2635 -4520 2693 -4514
rect 2753 -4520 2811 -4514
rect 2871 -4520 2929 -4514
rect 2989 -4520 3047 -4514
rect 3107 -4520 3165 -4514
rect 3225 -4520 3283 -4514
rect 3343 -4520 3401 -4514
rect 3461 -4520 3519 -4514
rect 3579 -4520 3637 -4514
rect 3697 -4520 3755 -4514
rect 3815 -4520 3873 -4514
rect 3933 -4520 3991 -4514
rect 4051 -4520 4109 -4514
rect 4169 -4520 4227 -4514
rect 4287 -4520 4345 -4514
rect 4405 -4520 4463 -4514
rect 4523 -4520 4581 -4514
rect 4641 -4520 4699 -4514
rect 4759 -4520 4817 -4514
rect 4877 -4520 4935 -4514
rect 4995 -4520 5053 -4514
rect 5113 -4520 5171 -4514
rect 5231 -4520 5289 -4514
rect 5349 -4520 5407 -4514
rect 5467 -4520 5525 -4514
rect 5585 -4520 5643 -4514
rect 5703 -4520 5761 -4514
rect 5821 -4520 5879 -4514
rect 5939 -4520 5997 -4514
rect 6057 -4520 6115 -4514
rect 6175 -4520 6233 -4514
rect 6293 -4520 6351 -4514
rect 6411 -4520 6469 -4514
rect 6529 -4520 6587 -4514
rect 6647 -4520 6705 -4514
rect 6765 -4520 6823 -4514
rect 6883 -4520 6941 -4514
rect 7001 -4520 7059 -4514
rect 7119 -4520 7177 -4514
rect 1337 -4554 1349 -4520
rect 1455 -4554 1467 -4520
rect 1573 -4554 1585 -4520
rect 1691 -4554 1703 -4520
rect 1809 -4554 1821 -4520
rect 1927 -4554 1939 -4520
rect 2045 -4554 2057 -4520
rect 2163 -4554 2175 -4520
rect 2281 -4554 2293 -4520
rect 2399 -4554 2411 -4520
rect 2517 -4554 2529 -4520
rect 2635 -4554 2647 -4520
rect 2753 -4554 2765 -4520
rect 2871 -4554 2883 -4520
rect 2989 -4554 3001 -4520
rect 3107 -4554 3119 -4520
rect 3225 -4554 3237 -4520
rect 3343 -4554 3355 -4520
rect 3461 -4554 3473 -4520
rect 3579 -4554 3591 -4520
rect 3697 -4554 3709 -4520
rect 3815 -4554 3827 -4520
rect 3933 -4554 3945 -4520
rect 4051 -4554 4063 -4520
rect 4169 -4554 4181 -4520
rect 4287 -4554 4299 -4520
rect 4405 -4554 4417 -4520
rect 4523 -4554 4535 -4520
rect 4641 -4554 4653 -4520
rect 4759 -4554 4771 -4520
rect 4877 -4554 4889 -4520
rect 4995 -4554 5007 -4520
rect 5113 -4554 5125 -4520
rect 5231 -4554 5243 -4520
rect 5349 -4554 5361 -4520
rect 5467 -4554 5479 -4520
rect 5585 -4554 5597 -4520
rect 5703 -4554 5715 -4520
rect 5821 -4554 5833 -4520
rect 5939 -4554 5951 -4520
rect 6057 -4554 6069 -4520
rect 6175 -4554 6187 -4520
rect 6293 -4554 6305 -4520
rect 6411 -4554 6423 -4520
rect 6529 -4554 6541 -4520
rect 6647 -4554 6659 -4520
rect 6765 -4554 6777 -4520
rect 6883 -4554 6895 -4520
rect 7001 -4554 7013 -4520
rect 7119 -4554 7131 -4520
rect 1337 -4560 1395 -4554
rect 1455 -4560 1513 -4554
rect 1573 -4560 1631 -4554
rect 1691 -4560 1749 -4554
rect 1809 -4560 1867 -4554
rect 1927 -4560 1985 -4554
rect 2045 -4560 2103 -4554
rect 2163 -4560 2221 -4554
rect 2281 -4560 2339 -4554
rect 2399 -4560 2457 -4554
rect 2517 -4560 2575 -4554
rect 2635 -4560 2693 -4554
rect 2753 -4560 2811 -4554
rect 2871 -4560 2929 -4554
rect 2989 -4560 3047 -4554
rect 3107 -4560 3165 -4554
rect 3225 -4560 3283 -4554
rect 3343 -4560 3401 -4554
rect 3461 -4560 3519 -4554
rect 3579 -4560 3637 -4554
rect 3697 -4560 3755 -4554
rect 3815 -4560 3873 -4554
rect 3933 -4560 3991 -4554
rect 4051 -4560 4109 -4554
rect 4169 -4560 4227 -4554
rect 4287 -4560 4345 -4554
rect 4405 -4560 4463 -4554
rect 4523 -4560 4581 -4554
rect 4641 -4560 4699 -4554
rect 4759 -4560 4817 -4554
rect 4877 -4560 4935 -4554
rect 4995 -4560 5053 -4554
rect 5113 -4560 5171 -4554
rect 5231 -4560 5289 -4554
rect 5349 -4560 5407 -4554
rect 5467 -4560 5525 -4554
rect 5585 -4560 5643 -4554
rect 5703 -4560 5761 -4554
rect 5821 -4560 5879 -4554
rect 5939 -4560 5997 -4554
rect 6057 -4560 6115 -4554
rect 6175 -4560 6233 -4554
rect 6293 -4560 6351 -4554
rect 6411 -4560 6469 -4554
rect 6529 -4560 6587 -4554
rect 6647 -4560 6705 -4554
rect 6765 -4560 6823 -4554
rect 6883 -4560 6941 -4554
rect 7001 -4560 7059 -4554
rect 7119 -4560 7177 -4554
rect 1337 -4724 1395 -4718
rect 1455 -4724 1513 -4718
rect 1573 -4724 1631 -4718
rect 1691 -4724 1749 -4718
rect 1809 -4724 1867 -4718
rect 1927 -4724 1985 -4718
rect 2045 -4724 2103 -4718
rect 2163 -4724 2221 -4718
rect 2281 -4724 2339 -4718
rect 2399 -4724 2457 -4718
rect 2517 -4724 2575 -4718
rect 2635 -4724 2693 -4718
rect 2753 -4724 2811 -4718
rect 2871 -4724 2929 -4718
rect 2989 -4724 3047 -4718
rect 3107 -4724 3165 -4718
rect 3225 -4724 3283 -4718
rect 3343 -4724 3401 -4718
rect 3461 -4724 3519 -4718
rect 3579 -4724 3637 -4718
rect 3697 -4724 3755 -4718
rect 3815 -4724 3873 -4718
rect 3933 -4724 3991 -4718
rect 4051 -4724 4109 -4718
rect 4169 -4724 4227 -4718
rect 4287 -4724 4345 -4718
rect 4405 -4724 4463 -4718
rect 4523 -4724 4581 -4718
rect 4641 -4724 4699 -4718
rect 4759 -4724 4817 -4718
rect 4877 -4724 4935 -4718
rect 4995 -4724 5053 -4718
rect 5113 -4724 5171 -4718
rect 5231 -4724 5289 -4718
rect 5349 -4724 5407 -4718
rect 5467 -4724 5525 -4718
rect 5585 -4724 5643 -4718
rect 5703 -4724 5761 -4718
rect 5821 -4724 5879 -4718
rect 5939 -4724 5997 -4718
rect 6057 -4724 6115 -4718
rect 6175 -4724 6233 -4718
rect 6293 -4724 6351 -4718
rect 6411 -4724 6469 -4718
rect 6529 -4724 6587 -4718
rect 6647 -4724 6705 -4718
rect 6765 -4724 6823 -4718
rect 6883 -4724 6941 -4718
rect 7001 -4724 7059 -4718
rect 7119 -4724 7177 -4718
rect 1337 -4758 1349 -4724
rect 1455 -4758 1467 -4724
rect 1573 -4758 1585 -4724
rect 1691 -4758 1703 -4724
rect 1809 -4758 1821 -4724
rect 1927 -4758 1939 -4724
rect 2045 -4758 2057 -4724
rect 2163 -4758 2175 -4724
rect 2281 -4758 2293 -4724
rect 2399 -4758 2411 -4724
rect 2517 -4758 2529 -4724
rect 2635 -4758 2647 -4724
rect 2753 -4758 2765 -4724
rect 2871 -4758 2883 -4724
rect 2989 -4758 3001 -4724
rect 3107 -4758 3119 -4724
rect 3225 -4758 3237 -4724
rect 3343 -4758 3355 -4724
rect 3461 -4758 3473 -4724
rect 3579 -4758 3591 -4724
rect 3697 -4758 3709 -4724
rect 3815 -4758 3827 -4724
rect 3933 -4758 3945 -4724
rect 4051 -4758 4063 -4724
rect 4169 -4758 4181 -4724
rect 4287 -4758 4299 -4724
rect 4405 -4758 4417 -4724
rect 4523 -4758 4535 -4724
rect 4641 -4758 4653 -4724
rect 4759 -4758 4771 -4724
rect 4877 -4758 4889 -4724
rect 4995 -4758 5007 -4724
rect 5113 -4758 5125 -4724
rect 5231 -4758 5243 -4724
rect 5349 -4758 5361 -4724
rect 5467 -4758 5479 -4724
rect 5585 -4758 5597 -4724
rect 5703 -4758 5715 -4724
rect 5821 -4758 5833 -4724
rect 5939 -4758 5951 -4724
rect 6057 -4758 6069 -4724
rect 6175 -4758 6187 -4724
rect 6293 -4758 6305 -4724
rect 6411 -4758 6423 -4724
rect 6529 -4758 6541 -4724
rect 6647 -4758 6659 -4724
rect 6765 -4758 6777 -4724
rect 6883 -4758 6895 -4724
rect 7001 -4758 7013 -4724
rect 7119 -4758 7131 -4724
rect 1337 -4764 1395 -4758
rect 1455 -4764 1513 -4758
rect 1573 -4764 1631 -4758
rect 1691 -4764 1749 -4758
rect 1809 -4764 1867 -4758
rect 1927 -4764 1985 -4758
rect 2045 -4764 2103 -4758
rect 2163 -4764 2221 -4758
rect 2281 -4764 2339 -4758
rect 2399 -4764 2457 -4758
rect 2517 -4764 2575 -4758
rect 2635 -4764 2693 -4758
rect 2753 -4764 2811 -4758
rect 2871 -4764 2929 -4758
rect 2989 -4764 3047 -4758
rect 3107 -4764 3165 -4758
rect 3225 -4764 3283 -4758
rect 3343 -4764 3401 -4758
rect 3461 -4764 3519 -4758
rect 3579 -4764 3637 -4758
rect 3697 -4764 3755 -4758
rect 3815 -4764 3873 -4758
rect 3933 -4764 3991 -4758
rect 4051 -4764 4109 -4758
rect 4169 -4764 4227 -4758
rect 4287 -4764 4345 -4758
rect 4405 -4764 4463 -4758
rect 4523 -4764 4581 -4758
rect 4641 -4764 4699 -4758
rect 4759 -4764 4817 -4758
rect 4877 -4764 4935 -4758
rect 4995 -4764 5053 -4758
rect 5113 -4764 5171 -4758
rect 5231 -4764 5289 -4758
rect 5349 -4764 5407 -4758
rect 5467 -4764 5525 -4758
rect 5585 -4764 5643 -4758
rect 5703 -4764 5761 -4758
rect 5821 -4764 5879 -4758
rect 5939 -4764 5997 -4758
rect 6057 -4764 6115 -4758
rect 6175 -4764 6233 -4758
rect 6293 -4764 6351 -4758
rect 6411 -4764 6469 -4758
rect 6529 -4764 6587 -4758
rect 6647 -4764 6705 -4758
rect 6765 -4764 6823 -4758
rect 6883 -4764 6941 -4758
rect 7001 -4764 7059 -4758
rect 7119 -4764 7177 -4758
rect 23119 -6093 23135 -6077
rect 23137 -6093 23153 -6077
rect 23103 -6109 23119 -6093
rect 23153 -6109 23169 -6093
rect 1337 -6288 1395 -6282
rect 1455 -6288 1513 -6282
rect 1573 -6288 1631 -6282
rect 1691 -6288 1749 -6282
rect 1809 -6288 1867 -6282
rect 1927 -6288 1985 -6282
rect 2045 -6288 2103 -6282
rect 2163 -6288 2221 -6282
rect 2281 -6288 2339 -6282
rect 2399 -6288 2457 -6282
rect 2517 -6288 2575 -6282
rect 2635 -6288 2693 -6282
rect 2753 -6288 2811 -6282
rect 2871 -6288 2929 -6282
rect 2989 -6288 3047 -6282
rect 3107 -6288 3165 -6282
rect 3225 -6288 3283 -6282
rect 3343 -6288 3401 -6282
rect 3461 -6288 3519 -6282
rect 3579 -6288 3637 -6282
rect 3697 -6288 3755 -6282
rect 3815 -6288 3873 -6282
rect 3933 -6288 3991 -6282
rect 4051 -6288 4109 -6282
rect 4169 -6288 4227 -6282
rect 4287 -6288 4345 -6282
rect 4405 -6288 4463 -6282
rect 4523 -6288 4581 -6282
rect 4641 -6288 4699 -6282
rect 4759 -6288 4817 -6282
rect 4877 -6288 4935 -6282
rect 4995 -6288 5053 -6282
rect 5113 -6288 5171 -6282
rect 5231 -6288 5289 -6282
rect 5349 -6288 5407 -6282
rect 5467 -6288 5525 -6282
rect 5585 -6288 5643 -6282
rect 5703 -6288 5761 -6282
rect 5821 -6288 5879 -6282
rect 5939 -6288 5997 -6282
rect 6057 -6288 6115 -6282
rect 6175 -6288 6233 -6282
rect 6293 -6288 6351 -6282
rect 6411 -6288 6469 -6282
rect 6529 -6288 6587 -6282
rect 6647 -6288 6705 -6282
rect 6765 -6288 6823 -6282
rect 6883 -6288 6941 -6282
rect 7001 -6288 7059 -6282
rect 7119 -6288 7177 -6282
rect 1337 -6322 1349 -6288
rect 1455 -6322 1467 -6288
rect 1573 -6322 1585 -6288
rect 1691 -6322 1703 -6288
rect 1809 -6322 1821 -6288
rect 1927 -6322 1939 -6288
rect 2045 -6322 2057 -6288
rect 2163 -6322 2175 -6288
rect 2281 -6322 2293 -6288
rect 2399 -6322 2411 -6288
rect 2517 -6322 2529 -6288
rect 2635 -6322 2647 -6288
rect 2753 -6322 2765 -6288
rect 2871 -6322 2883 -6288
rect 2989 -6322 3001 -6288
rect 3107 -6322 3119 -6288
rect 3225 -6322 3237 -6288
rect 3343 -6322 3355 -6288
rect 3461 -6322 3473 -6288
rect 3579 -6322 3591 -6288
rect 3697 -6322 3709 -6288
rect 3815 -6322 3827 -6288
rect 3933 -6322 3945 -6288
rect 4051 -6322 4063 -6288
rect 4169 -6322 4181 -6288
rect 4287 -6322 4299 -6288
rect 4405 -6322 4417 -6288
rect 4523 -6322 4535 -6288
rect 4641 -6322 4653 -6288
rect 4759 -6322 4771 -6288
rect 4877 -6322 4889 -6288
rect 4995 -6322 5007 -6288
rect 5113 -6322 5125 -6288
rect 5231 -6322 5243 -6288
rect 5349 -6322 5361 -6288
rect 5467 -6322 5479 -6288
rect 5585 -6322 5597 -6288
rect 5703 -6322 5715 -6288
rect 5821 -6322 5833 -6288
rect 5939 -6322 5951 -6288
rect 6057 -6322 6069 -6288
rect 6175 -6322 6187 -6288
rect 6293 -6322 6305 -6288
rect 6411 -6322 6423 -6288
rect 6529 -6322 6541 -6288
rect 6647 -6322 6659 -6288
rect 6765 -6322 6777 -6288
rect 6883 -6322 6895 -6288
rect 7001 -6322 7013 -6288
rect 7119 -6322 7131 -6288
rect 1337 -6328 1395 -6322
rect 1455 -6328 1513 -6322
rect 1573 -6328 1631 -6322
rect 1691 -6328 1749 -6322
rect 1809 -6328 1867 -6322
rect 1927 -6328 1985 -6322
rect 2045 -6328 2103 -6322
rect 2163 -6328 2221 -6322
rect 2281 -6328 2339 -6322
rect 2399 -6328 2457 -6322
rect 2517 -6328 2575 -6322
rect 2635 -6328 2693 -6322
rect 2753 -6328 2811 -6322
rect 2871 -6328 2929 -6322
rect 2989 -6328 3047 -6322
rect 3107 -6328 3165 -6322
rect 3225 -6328 3283 -6322
rect 3343 -6328 3401 -6322
rect 3461 -6328 3519 -6322
rect 3579 -6328 3637 -6322
rect 3697 -6328 3755 -6322
rect 3815 -6328 3873 -6322
rect 3933 -6328 3991 -6322
rect 4051 -6328 4109 -6322
rect 4169 -6328 4227 -6322
rect 4287 -6328 4345 -6322
rect 4405 -6328 4463 -6322
rect 4523 -6328 4581 -6322
rect 4641 -6328 4699 -6322
rect 4759 -6328 4817 -6322
rect 4877 -6328 4935 -6322
rect 4995 -6328 5053 -6322
rect 5113 -6328 5171 -6322
rect 5231 -6328 5289 -6322
rect 5349 -6328 5407 -6322
rect 5467 -6328 5525 -6322
rect 5585 -6328 5643 -6322
rect 5703 -6328 5761 -6322
rect 5821 -6328 5879 -6322
rect 5939 -6328 5997 -6322
rect 6057 -6328 6115 -6322
rect 6175 -6328 6233 -6322
rect 6293 -6328 6351 -6322
rect 6411 -6328 6469 -6322
rect 6529 -6328 6587 -6322
rect 6647 -6328 6705 -6322
rect 6765 -6328 6823 -6322
rect 6883 -6328 6941 -6322
rect 7001 -6328 7059 -6322
rect 7119 -6328 7177 -6322
rect 9735 -6513 9793 -6507
rect 9853 -6513 9911 -6507
rect 9735 -6547 9747 -6513
rect 9853 -6547 9865 -6513
rect 9735 -6553 9793 -6547
rect 9853 -6553 9911 -6547
rect 23103 -6969 23119 -6953
rect 23153 -6969 23169 -6953
rect 23119 -6985 23135 -6969
rect 23137 -6985 23153 -6969
rect 3063 -7057 3121 -7051
rect 3181 -7057 3239 -7051
rect 3299 -7057 3357 -7051
rect 3417 -7057 3475 -7051
rect 3535 -7057 3593 -7051
rect 3653 -7057 3711 -7051
rect 3771 -7057 3829 -7051
rect 3889 -7057 3947 -7051
rect 4007 -7057 4065 -7051
rect 4125 -7057 4183 -7051
rect 4243 -7057 4301 -7051
rect 4361 -7057 4419 -7051
rect 4479 -7057 4537 -7051
rect 4597 -7057 4655 -7051
rect 4715 -7057 4773 -7051
rect 5061 -7057 5119 -7051
rect 5179 -7057 5237 -7051
rect 5297 -7057 5355 -7051
rect 5415 -7057 5473 -7051
rect 5533 -7057 5591 -7051
rect 5651 -7057 5709 -7051
rect 5769 -7057 5827 -7051
rect 5887 -7057 5945 -7051
rect 6005 -7057 6063 -7051
rect 6123 -7057 6181 -7051
rect 6241 -7057 6299 -7051
rect 6359 -7057 6417 -7051
rect 6477 -7057 6535 -7051
rect 6595 -7057 6653 -7051
rect 6713 -7057 6771 -7051
rect 3063 -7091 3075 -7057
rect 3181 -7091 3193 -7057
rect 3299 -7091 3311 -7057
rect 3417 -7091 3429 -7057
rect 3535 -7091 3547 -7057
rect 3653 -7091 3665 -7057
rect 3771 -7091 3783 -7057
rect 3889 -7091 3901 -7057
rect 4007 -7091 4019 -7057
rect 4125 -7091 4137 -7057
rect 4243 -7091 4255 -7057
rect 4361 -7091 4373 -7057
rect 4479 -7091 4491 -7057
rect 4597 -7091 4609 -7057
rect 4715 -7091 4727 -7057
rect 5061 -7091 5073 -7057
rect 5179 -7091 5191 -7057
rect 5297 -7091 5309 -7057
rect 5415 -7091 5427 -7057
rect 5533 -7091 5545 -7057
rect 5651 -7091 5663 -7057
rect 5769 -7091 5781 -7057
rect 5887 -7091 5899 -7057
rect 6005 -7091 6017 -7057
rect 6123 -7091 6135 -7057
rect 6241 -7091 6253 -7057
rect 6359 -7091 6371 -7057
rect 6477 -7091 6489 -7057
rect 6595 -7091 6607 -7057
rect 6713 -7091 6725 -7057
rect 3063 -7097 3121 -7091
rect 3181 -7097 3239 -7091
rect 3299 -7097 3357 -7091
rect 3417 -7097 3475 -7091
rect 3535 -7097 3593 -7091
rect 3653 -7097 3711 -7091
rect 3771 -7097 3829 -7091
rect 3889 -7097 3947 -7091
rect 4007 -7097 4065 -7091
rect 4125 -7097 4183 -7091
rect 4243 -7097 4301 -7091
rect 4361 -7097 4419 -7091
rect 4479 -7097 4537 -7091
rect 4597 -7097 4655 -7091
rect 4715 -7097 4773 -7091
rect 5061 -7097 5119 -7091
rect 5179 -7097 5237 -7091
rect 5297 -7097 5355 -7091
rect 5415 -7097 5473 -7091
rect 5533 -7097 5591 -7091
rect 5651 -7097 5709 -7091
rect 5769 -7097 5827 -7091
rect 5887 -7097 5945 -7091
rect 6005 -7097 6063 -7091
rect 6123 -7097 6181 -7091
rect 6241 -7097 6299 -7091
rect 6359 -7097 6417 -7091
rect 6477 -7097 6535 -7091
rect 6595 -7097 6653 -7091
rect 6713 -7097 6771 -7091
rect 9735 -7223 9793 -7217
rect 9853 -7223 9911 -7217
rect 9735 -7257 9747 -7223
rect 9853 -7257 9865 -7223
rect 9735 -7263 9793 -7257
rect 9853 -7263 9911 -7257
rect 3063 -8585 3121 -8579
rect 3181 -8585 3239 -8579
rect 3299 -8585 3357 -8579
rect 3417 -8585 3475 -8579
rect 3535 -8585 3593 -8579
rect 3653 -8585 3711 -8579
rect 3771 -8585 3829 -8579
rect 3889 -8585 3947 -8579
rect 4007 -8585 4065 -8579
rect 4125 -8585 4183 -8579
rect 4243 -8585 4301 -8579
rect 4361 -8585 4419 -8579
rect 4479 -8585 4537 -8579
rect 4597 -8585 4655 -8579
rect 4715 -8585 4773 -8579
rect 5061 -8585 5119 -8579
rect 5179 -8585 5237 -8579
rect 5297 -8585 5355 -8579
rect 5415 -8585 5473 -8579
rect 5533 -8585 5591 -8579
rect 5651 -8585 5709 -8579
rect 5769 -8585 5827 -8579
rect 5887 -8585 5945 -8579
rect 6005 -8585 6063 -8579
rect 6123 -8585 6181 -8579
rect 6241 -8585 6299 -8579
rect 6359 -8585 6417 -8579
rect 6477 -8585 6535 -8579
rect 6595 -8585 6653 -8579
rect 6713 -8585 6771 -8579
rect 3063 -8619 3075 -8585
rect 3181 -8619 3193 -8585
rect 3299 -8619 3311 -8585
rect 3417 -8619 3429 -8585
rect 3535 -8619 3547 -8585
rect 3653 -8619 3665 -8585
rect 3771 -8619 3783 -8585
rect 3889 -8619 3901 -8585
rect 4007 -8619 4019 -8585
rect 4125 -8619 4137 -8585
rect 4243 -8619 4255 -8585
rect 4361 -8619 4373 -8585
rect 4479 -8619 4491 -8585
rect 4597 -8619 4609 -8585
rect 4715 -8619 4727 -8585
rect 5061 -8619 5073 -8585
rect 5179 -8619 5191 -8585
rect 5297 -8619 5309 -8585
rect 5415 -8619 5427 -8585
rect 5533 -8619 5545 -8585
rect 5651 -8619 5663 -8585
rect 5769 -8619 5781 -8585
rect 5887 -8619 5899 -8585
rect 6005 -8619 6017 -8585
rect 6123 -8619 6135 -8585
rect 6241 -8619 6253 -8585
rect 6359 -8619 6371 -8585
rect 6477 -8619 6489 -8585
rect 6595 -8619 6607 -8585
rect 6713 -8619 6725 -8585
rect 3063 -8625 3121 -8619
rect 3181 -8625 3239 -8619
rect 3299 -8625 3357 -8619
rect 3417 -8625 3475 -8619
rect 3535 -8625 3593 -8619
rect 3653 -8625 3711 -8619
rect 3771 -8625 3829 -8619
rect 3889 -8625 3947 -8619
rect 4007 -8625 4065 -8619
rect 4125 -8625 4183 -8619
rect 4243 -8625 4301 -8619
rect 4361 -8625 4419 -8619
rect 4479 -8625 4537 -8619
rect 4597 -8625 4655 -8619
rect 4715 -8625 4773 -8619
rect 5061 -8625 5119 -8619
rect 5179 -8625 5237 -8619
rect 5297 -8625 5355 -8619
rect 5415 -8625 5473 -8619
rect 5533 -8625 5591 -8619
rect 5651 -8625 5709 -8619
rect 5769 -8625 5827 -8619
rect 5887 -8625 5945 -8619
rect 6005 -8625 6063 -8619
rect 6123 -8625 6181 -8619
rect 6241 -8625 6299 -8619
rect 6359 -8625 6417 -8619
rect 6477 -8625 6535 -8619
rect 6595 -8625 6653 -8619
rect 6713 -8625 6771 -8619
<< nwell >>
rect 7530 1942 8351 2054
rect 8587 1942 10349 2054
rect 12350 1884 12531 2058
rect 12571 1884 13003 2058
rect 13043 1884 13947 2058
rect 13987 1884 15835 2058
rect 15875 1884 19611 2058
rect 19651 1884 20940 2058
<< ndiffc >>
rect 12647 -7518 12681 -6642
rect 12795 -7518 12829 -6642
rect 12943 -7518 12977 -6642
rect 13091 -7518 13125 -6642
rect 13239 -7518 13273 -6642
rect 13387 -7518 13421 -6642
rect 13535 -7518 13569 -6642
rect 13683 -7518 13717 -6642
rect 13831 -7518 13865 -6642
rect 13979 -7518 14013 -6642
rect 14127 -7518 14161 -6642
rect 14275 -7518 14309 -6642
rect 14423 -7518 14457 -6642
rect 14571 -7518 14605 -6642
rect 14719 -7518 14753 -6642
rect 14867 -7518 14901 -6642
rect 15015 -7518 15049 -6642
rect 15163 -7518 15197 -6642
rect 15311 -7518 15345 -6642
rect 15459 -7518 15493 -6642
rect 15607 -7518 15641 -6642
rect 15755 -7518 15789 -6642
rect 15903 -7518 15937 -6642
rect 16051 -7518 16085 -6642
rect 16199 -7518 16233 -6642
rect 16347 -7518 16381 -6642
rect 16495 -7518 16529 -6642
rect 16643 -7518 16677 -6642
rect 16791 -7518 16825 -6642
rect 16939 -7518 16973 -6642
rect 17087 -7518 17121 -6642
rect 17235 -7518 17269 -6642
rect 17383 -7518 17417 -6642
rect 17531 -7518 17565 -6642
rect 17679 -7518 17713 -6642
rect 17827 -7518 17861 -6642
rect 17975 -7518 18009 -6642
rect 18123 -7518 18157 -6642
rect 18271 -7518 18305 -6642
rect 18419 -7518 18453 -6642
rect 18567 -7518 18601 -6642
rect 18715 -7518 18749 -6642
rect 18863 -7518 18897 -6642
rect 19011 -7518 19045 -6642
rect 19159 -7518 19193 -6642
rect 19307 -7518 19341 -6642
rect 19455 -7518 19489 -6642
rect 19603 -7518 19637 -6642
rect 19751 -7518 19785 -6642
rect 19899 -7518 19933 -6642
rect 20047 -7518 20081 -6642
rect 20195 -7518 20229 -6642
rect 20343 -7518 20377 -6642
rect 20491 -7518 20525 -6642
rect 20639 -7518 20673 -6642
rect 20787 -7518 20821 -6642
rect 20935 -7518 20969 -6642
rect 21083 -7518 21117 -6642
rect 21231 -7518 21265 -6642
rect 21379 -7518 21413 -6642
rect 21527 -7518 21561 -6642
rect 21675 -7518 21709 -6642
rect 21823 -7518 21857 -6642
rect 21971 -7518 22005 -6642
rect 20343 -8636 20377 -7760
rect 20491 -8636 20525 -7760
rect 20639 -8636 20673 -7760
rect 20787 -8636 20821 -7760
rect 20935 -8636 20969 -7760
rect 21083 -8636 21117 -7760
rect 21231 -8636 21265 -7760
rect 21379 -8636 21413 -7760
<< poly >>
rect 7539 2040 7605 2054
rect 7539 2006 7555 2040
rect 7589 2006 7605 2040
rect 7539 1990 7605 2006
rect 7657 2040 7723 2054
rect 7657 2006 7673 2040
rect 7707 2006 7723 2040
rect 7657 1990 7723 2006
rect 7775 2040 7841 2054
rect 7775 2006 7791 2040
rect 7825 2006 7841 2040
rect 7775 1990 7841 2006
rect 7893 2040 7959 2054
rect 7893 2006 7909 2040
rect 7943 2006 7959 2040
rect 7893 1990 7959 2006
rect 8011 2040 8077 2054
rect 8011 2006 8027 2040
rect 8061 2006 8077 2040
rect 8011 1990 8077 2006
rect 8129 2040 8195 2054
rect 8129 2006 8145 2040
rect 8179 2006 8195 2040
rect 8129 1990 8195 2006
rect 8247 2040 8313 2054
rect 8247 2006 8263 2040
rect 8297 2006 8313 2040
rect 8247 1990 8313 2006
rect 8593 2040 8659 2054
rect 8593 2006 8609 2040
rect 8643 2006 8659 2040
rect 8593 1990 8659 2006
rect 8711 2040 8777 2054
rect 8711 2006 8727 2040
rect 8761 2006 8777 2040
rect 8711 1990 8777 2006
rect 8829 2040 8895 2054
rect 8829 2006 8845 2040
rect 8879 2006 8895 2040
rect 8829 1990 8895 2006
rect 8947 2040 9013 2054
rect 8947 2006 8963 2040
rect 8997 2006 9013 2040
rect 8947 1990 9013 2006
rect 9065 2040 9131 2054
rect 9065 2006 9081 2040
rect 9115 2006 9131 2040
rect 9065 1990 9131 2006
rect 9183 2040 9249 2054
rect 9183 2006 9199 2040
rect 9233 2006 9249 2040
rect 9183 1990 9249 2006
rect 9301 2040 9367 2054
rect 9301 2006 9317 2040
rect 9351 2006 9367 2040
rect 9301 1990 9367 2006
rect 9419 2040 9485 2054
rect 9419 2006 9435 2040
rect 9469 2006 9485 2040
rect 9419 1990 9485 2006
rect 9537 2040 9603 2054
rect 9537 2006 9553 2040
rect 9587 2006 9603 2040
rect 9537 1990 9603 2006
rect 9655 2040 9721 2054
rect 9655 2006 9671 2040
rect 9705 2006 9721 2040
rect 9655 1990 9721 2006
rect 9773 2040 9839 2054
rect 9773 2006 9789 2040
rect 9823 2006 9839 2040
rect 9773 1990 9839 2006
rect 9891 2040 9957 2054
rect 9891 2006 9907 2040
rect 9941 2006 9957 2040
rect 9891 1990 9957 2006
rect 10009 2040 10075 2054
rect 10009 2006 10025 2040
rect 10059 2006 10075 2040
rect 10009 1990 10075 2006
rect 10127 2040 10193 2054
rect 10127 2006 10143 2040
rect 10177 2006 10193 2040
rect 10127 1990 10193 2006
rect 10245 2040 10311 2054
rect 10245 2006 10261 2040
rect 10295 2006 10311 2040
rect 10245 1990 10311 2006
rect 12665 2039 12723 2045
rect 12665 2005 12677 2039
rect 12711 2005 12723 2039
rect 12665 1989 12723 2005
rect 12779 2039 12845 2055
rect 12779 2005 12795 2039
rect 12829 2005 12845 2039
rect 12779 1989 12845 2005
rect 12897 2039 12963 2055
rect 12897 2005 12913 2039
rect 12947 2005 12963 2039
rect 12897 1989 12963 2005
rect 13015 2039 13081 2055
rect 13015 2005 13031 2039
rect 13065 2005 13081 2039
rect 13015 1989 13081 2005
rect 13133 2039 13199 2055
rect 13133 2005 13149 2039
rect 13183 2005 13199 2039
rect 13133 1989 13199 2005
rect 13251 2039 13317 2055
rect 13251 2005 13267 2039
rect 13301 2005 13317 2039
rect 13251 1989 13317 2005
rect 13369 2039 13435 2055
rect 13369 2005 13385 2039
rect 13419 2005 13435 2039
rect 13369 1989 13435 2005
rect 13487 2039 13553 2055
rect 13487 2005 13503 2039
rect 13537 2005 13553 2039
rect 13487 1989 13553 2005
rect 13605 2039 13671 2055
rect 13605 2005 13621 2039
rect 13655 2005 13671 2039
rect 13605 1989 13671 2005
rect 13723 2039 13789 2055
rect 13723 2005 13739 2039
rect 13773 2005 13789 2039
rect 13723 1989 13789 2005
rect 13841 2039 13907 2055
rect 13841 2005 13857 2039
rect 13891 2005 13907 2039
rect 13841 1989 13907 2005
rect 13959 2039 14025 2055
rect 13959 2005 13975 2039
rect 14009 2005 14025 2039
rect 13959 1989 14025 2005
rect 14077 2039 14143 2055
rect 14077 2005 14093 2039
rect 14127 2005 14143 2039
rect 14077 1989 14143 2005
rect 14195 2039 14261 2055
rect 14195 2005 14211 2039
rect 14245 2005 14261 2039
rect 14195 1989 14261 2005
rect 14313 2039 14379 2055
rect 14313 2005 14329 2039
rect 14363 2005 14379 2039
rect 14313 1989 14379 2005
rect 14431 2039 14497 2055
rect 14431 2005 14447 2039
rect 14481 2005 14497 2039
rect 14431 1989 14497 2005
rect 14549 2039 14615 2055
rect 14549 2005 14565 2039
rect 14599 2005 14615 2039
rect 14549 1989 14615 2005
rect 14667 2039 14733 2055
rect 14667 2005 14683 2039
rect 14717 2005 14733 2039
rect 14667 1989 14733 2005
rect 14785 2039 14851 2055
rect 14785 2005 14801 2039
rect 14835 2005 14851 2039
rect 14785 1989 14851 2005
rect 14903 2039 14969 2055
rect 14903 2005 14919 2039
rect 14953 2005 14969 2039
rect 14903 1989 14969 2005
rect 15021 2039 15087 2055
rect 15021 2005 15037 2039
rect 15071 2005 15087 2039
rect 15021 1989 15087 2005
rect 15139 2039 15205 2055
rect 15139 2005 15155 2039
rect 15189 2005 15205 2039
rect 15139 1989 15205 2005
rect 15257 2039 15323 2055
rect 15257 2005 15273 2039
rect 15307 2005 15323 2039
rect 15257 1989 15323 2005
rect 15375 2039 15441 2055
rect 15375 2005 15391 2039
rect 15425 2005 15441 2039
rect 15375 1989 15441 2005
rect 15493 2039 15559 2055
rect 15493 2005 15509 2039
rect 15543 2005 15559 2039
rect 15493 1989 15559 2005
rect 15611 2039 15677 2055
rect 15611 2005 15627 2039
rect 15661 2005 15677 2039
rect 15611 1989 15677 2005
rect 15729 2039 15795 2055
rect 15729 2005 15745 2039
rect 15779 2005 15795 2039
rect 15729 1989 15795 2005
rect 15847 2039 15913 2055
rect 15847 2005 15863 2039
rect 15897 2005 15913 2039
rect 15847 1989 15913 2005
rect 15965 2039 16031 2055
rect 15965 2005 15981 2039
rect 16015 2005 16031 2039
rect 15965 1989 16031 2005
rect 16083 2039 16149 2055
rect 16083 2005 16099 2039
rect 16133 2005 16149 2039
rect 16083 1989 16149 2005
rect 16201 2039 16267 2055
rect 16201 2005 16217 2039
rect 16251 2005 16267 2039
rect 16201 1989 16267 2005
rect 16319 2039 16385 2055
rect 16319 2005 16335 2039
rect 16369 2005 16385 2039
rect 16319 1989 16385 2005
rect 16437 2039 16503 2055
rect 16437 2005 16453 2039
rect 16487 2005 16503 2039
rect 16437 1989 16503 2005
rect 16555 2039 16621 2055
rect 16555 2005 16571 2039
rect 16605 2005 16621 2039
rect 16555 1989 16621 2005
rect 16673 2039 16739 2055
rect 16673 2005 16689 2039
rect 16723 2005 16739 2039
rect 16673 1989 16739 2005
rect 16791 2039 16857 2055
rect 16791 2005 16807 2039
rect 16841 2005 16857 2039
rect 16791 1989 16857 2005
rect 16909 2039 16975 2055
rect 16909 2005 16925 2039
rect 16959 2005 16975 2039
rect 16909 1989 16975 2005
rect 17027 2039 17093 2055
rect 17027 2005 17043 2039
rect 17077 2005 17093 2039
rect 17027 1989 17093 2005
rect 17145 2039 17211 2055
rect 17145 2005 17161 2039
rect 17195 2005 17211 2039
rect 17145 1989 17211 2005
rect 17263 2039 17329 2055
rect 17263 2005 17279 2039
rect 17313 2005 17329 2039
rect 17263 1989 17329 2005
rect 17381 2039 17447 2055
rect 17381 2005 17397 2039
rect 17431 2005 17447 2039
rect 17381 1989 17447 2005
rect 17499 2039 17565 2055
rect 17499 2005 17515 2039
rect 17549 2005 17565 2039
rect 17499 1989 17565 2005
rect 17617 2039 17683 2055
rect 17617 2005 17633 2039
rect 17667 2005 17683 2039
rect 17617 1989 17683 2005
rect 17735 2039 17801 2055
rect 17735 2005 17751 2039
rect 17785 2005 17801 2039
rect 17735 1989 17801 2005
rect 17853 2039 17919 2055
rect 17853 2005 17869 2039
rect 17903 2005 17919 2039
rect 17853 1989 17919 2005
rect 17971 2039 18037 2055
rect 17971 2005 17987 2039
rect 18021 2005 18037 2039
rect 17971 1989 18037 2005
rect 18089 2039 18155 2055
rect 18089 2005 18105 2039
rect 18139 2005 18155 2039
rect 18089 1989 18155 2005
rect 18207 2039 18273 2055
rect 18207 2005 18223 2039
rect 18257 2005 18273 2039
rect 18207 1989 18273 2005
rect 18325 2039 18391 2055
rect 18325 2005 18341 2039
rect 18375 2005 18391 2039
rect 18325 1989 18391 2005
rect 18443 2039 18509 2055
rect 18443 2005 18459 2039
rect 18493 2005 18509 2039
rect 18443 1989 18509 2005
rect 18561 2039 18627 2055
rect 18561 2005 18577 2039
rect 18611 2005 18627 2039
rect 18561 1989 18627 2005
rect 18679 2039 18745 2055
rect 18679 2005 18695 2039
rect 18729 2005 18745 2039
rect 18679 1989 18745 2005
rect 18797 2039 18863 2055
rect 18797 2005 18813 2039
rect 18847 2005 18863 2039
rect 18797 1989 18863 2005
rect 18915 2039 18981 2055
rect 18915 2005 18931 2039
rect 18965 2005 18981 2039
rect 18915 1989 18981 2005
rect 19033 2039 19099 2055
rect 19033 2005 19049 2039
rect 19083 2005 19099 2039
rect 19033 1989 19099 2005
rect 19151 2039 19217 2055
rect 19151 2005 19167 2039
rect 19201 2005 19217 2039
rect 19151 1989 19217 2005
rect 19269 2039 19335 2055
rect 19269 2005 19285 2039
rect 19319 2005 19335 2039
rect 19269 1989 19335 2005
rect 19387 2039 19453 2055
rect 19387 2005 19403 2039
rect 19437 2005 19453 2039
rect 19387 1989 19453 2005
rect 19505 2039 19571 2055
rect 19505 2005 19521 2039
rect 19555 2005 19571 2039
rect 19505 1989 19571 2005
rect 19623 2039 19689 2055
rect 19623 2005 19639 2039
rect 19673 2005 19689 2039
rect 19623 1989 19689 2005
rect 19741 2039 19807 2055
rect 19741 2005 19757 2039
rect 19791 2005 19807 2039
rect 19741 1989 19807 2005
rect 19859 2039 19925 2055
rect 19859 2005 19875 2039
rect 19909 2005 19925 2039
rect 19859 1989 19925 2005
rect 19977 2039 20043 2055
rect 19977 2005 19993 2039
rect 20027 2005 20043 2039
rect 19977 1989 20043 2005
rect 20095 2039 20161 2055
rect 20095 2005 20111 2039
rect 20145 2005 20161 2039
rect 20095 1989 20161 2005
rect 20213 2039 20279 2055
rect 20213 2005 20229 2039
rect 20263 2005 20279 2039
rect 20213 1989 20279 2005
rect 20331 2039 20397 2055
rect 20331 2005 20347 2039
rect 20381 2005 20397 2039
rect 20331 1989 20397 2005
rect 20449 2039 20515 2055
rect 20449 2005 20465 2039
rect 20499 2005 20515 2039
rect 20449 1989 20515 2005
rect 20567 2039 20633 2055
rect 20567 2005 20583 2039
rect 20617 2005 20633 2039
rect 20567 1989 20633 2005
rect 20685 2039 20751 2055
rect 20685 2005 20701 2039
rect 20735 2005 20751 2039
rect 20685 1989 20751 2005
rect 20803 2039 20869 2055
rect 20803 2005 20819 2039
rect 20853 2005 20869 2039
rect 20803 1989 20869 2005
rect 20921 2039 20987 2055
rect 20921 2005 20937 2039
rect 20971 2005 20987 2039
rect 20921 1989 20987 2005
rect 21039 2039 21105 2055
rect 21039 2005 21055 2039
rect 21089 2005 21105 2039
rect 21039 1989 21105 2005
rect 21157 2039 21223 2055
rect 21157 2005 21173 2039
rect 21207 2005 21223 2039
rect 21157 1989 21223 2005
rect 21275 2039 21341 2055
rect 21275 2005 21291 2039
rect 21325 2005 21341 2039
rect 21275 1989 21341 2005
rect 12665 1931 12723 1947
rect 12665 1897 12677 1931
rect 12711 1897 12723 1931
rect 12665 1891 12723 1897
rect 12779 1931 12845 1947
rect 12779 1897 12795 1931
rect 12829 1897 12845 1931
rect 12779 1881 12845 1897
rect 12897 1931 12963 1947
rect 12897 1897 12913 1931
rect 12947 1897 12963 1931
rect 12897 1881 12963 1897
rect 13015 1931 13081 1947
rect 13015 1897 13031 1931
rect 13065 1897 13081 1931
rect 13015 1881 13081 1897
rect 13133 1931 13199 1947
rect 13133 1897 13149 1931
rect 13183 1897 13199 1931
rect 13133 1881 13199 1897
rect 13251 1931 13317 1947
rect 13251 1897 13267 1931
rect 13301 1897 13317 1931
rect 13251 1881 13317 1897
rect 13369 1931 13435 1947
rect 13369 1897 13385 1931
rect 13419 1897 13435 1931
rect 13369 1881 13435 1897
rect 13487 1931 13553 1947
rect 13487 1897 13503 1931
rect 13537 1897 13553 1931
rect 13487 1881 13553 1897
rect 13605 1931 13671 1947
rect 13605 1897 13621 1931
rect 13655 1897 13671 1931
rect 13605 1881 13671 1897
rect 13723 1931 13789 1947
rect 13723 1897 13739 1931
rect 13773 1897 13789 1931
rect 13723 1881 13789 1897
rect 13841 1931 13907 1947
rect 13841 1897 13857 1931
rect 13891 1897 13907 1931
rect 13841 1881 13907 1897
rect 13959 1931 14025 1947
rect 13959 1897 13975 1931
rect 14009 1897 14025 1931
rect 13959 1881 14025 1897
rect 14077 1931 14143 1947
rect 14077 1897 14093 1931
rect 14127 1897 14143 1931
rect 14077 1881 14143 1897
rect 14195 1931 14261 1947
rect 14195 1897 14211 1931
rect 14245 1897 14261 1931
rect 14195 1881 14261 1897
rect 14313 1931 14379 1947
rect 14313 1897 14329 1931
rect 14363 1897 14379 1931
rect 14313 1881 14379 1897
rect 14431 1931 14497 1947
rect 14431 1897 14447 1931
rect 14481 1897 14497 1931
rect 14431 1881 14497 1897
rect 14549 1931 14615 1947
rect 14549 1897 14565 1931
rect 14599 1897 14615 1931
rect 14549 1881 14615 1897
rect 14667 1931 14733 1947
rect 14667 1897 14683 1931
rect 14717 1897 14733 1931
rect 14667 1881 14733 1897
rect 14785 1931 14851 1947
rect 14785 1897 14801 1931
rect 14835 1897 14851 1931
rect 14785 1881 14851 1897
rect 14903 1931 14969 1947
rect 14903 1897 14919 1931
rect 14953 1897 14969 1931
rect 14903 1881 14969 1897
rect 15021 1931 15087 1947
rect 15021 1897 15037 1931
rect 15071 1897 15087 1931
rect 15021 1881 15087 1897
rect 15139 1931 15205 1947
rect 15139 1897 15155 1931
rect 15189 1897 15205 1931
rect 15139 1881 15205 1897
rect 15257 1931 15323 1947
rect 15257 1897 15273 1931
rect 15307 1897 15323 1931
rect 15257 1881 15323 1897
rect 15375 1931 15441 1947
rect 15375 1897 15391 1931
rect 15425 1897 15441 1931
rect 15375 1881 15441 1897
rect 15493 1931 15559 1947
rect 15493 1897 15509 1931
rect 15543 1897 15559 1931
rect 15493 1881 15559 1897
rect 15611 1931 15677 1947
rect 15611 1897 15627 1931
rect 15661 1897 15677 1931
rect 15611 1881 15677 1897
rect 15729 1931 15795 1947
rect 15729 1897 15745 1931
rect 15779 1897 15795 1931
rect 15729 1881 15795 1897
rect 15847 1931 15913 1947
rect 15847 1897 15863 1931
rect 15897 1897 15913 1931
rect 15847 1881 15913 1897
rect 15965 1931 16031 1947
rect 15965 1897 15981 1931
rect 16015 1897 16031 1931
rect 15965 1881 16031 1897
rect 16083 1931 16149 1947
rect 16083 1897 16099 1931
rect 16133 1897 16149 1931
rect 16083 1881 16149 1897
rect 16201 1931 16267 1947
rect 16201 1897 16217 1931
rect 16251 1897 16267 1931
rect 16201 1881 16267 1897
rect 16319 1931 16385 1947
rect 16319 1897 16335 1931
rect 16369 1897 16385 1931
rect 16319 1881 16385 1897
rect 16437 1931 16503 1947
rect 16437 1897 16453 1931
rect 16487 1897 16503 1931
rect 16437 1881 16503 1897
rect 16555 1931 16621 1947
rect 16555 1897 16571 1931
rect 16605 1897 16621 1931
rect 16555 1881 16621 1897
rect 16673 1931 16739 1947
rect 16673 1897 16689 1931
rect 16723 1897 16739 1931
rect 16673 1881 16739 1897
rect 16791 1931 16857 1947
rect 16791 1897 16807 1931
rect 16841 1897 16857 1931
rect 16791 1881 16857 1897
rect 16909 1931 16975 1947
rect 16909 1897 16925 1931
rect 16959 1897 16975 1931
rect 16909 1881 16975 1897
rect 17027 1931 17093 1947
rect 17027 1897 17043 1931
rect 17077 1897 17093 1931
rect 17027 1881 17093 1897
rect 17145 1931 17211 1947
rect 17145 1897 17161 1931
rect 17195 1897 17211 1931
rect 17145 1881 17211 1897
rect 17263 1931 17329 1947
rect 17263 1897 17279 1931
rect 17313 1897 17329 1931
rect 17263 1881 17329 1897
rect 17381 1931 17447 1947
rect 17381 1897 17397 1931
rect 17431 1897 17447 1931
rect 17381 1881 17447 1897
rect 17499 1931 17565 1947
rect 17499 1897 17515 1931
rect 17549 1897 17565 1931
rect 17499 1881 17565 1897
rect 17617 1931 17683 1947
rect 17617 1897 17633 1931
rect 17667 1897 17683 1931
rect 17617 1881 17683 1897
rect 17735 1931 17801 1947
rect 17735 1897 17751 1931
rect 17785 1897 17801 1931
rect 17735 1881 17801 1897
rect 17853 1931 17919 1947
rect 17853 1897 17869 1931
rect 17903 1897 17919 1931
rect 17853 1881 17919 1897
rect 17971 1931 18037 1947
rect 17971 1897 17987 1931
rect 18021 1897 18037 1931
rect 17971 1881 18037 1897
rect 18089 1931 18155 1947
rect 18089 1897 18105 1931
rect 18139 1897 18155 1931
rect 18089 1881 18155 1897
rect 18207 1931 18273 1947
rect 18207 1897 18223 1931
rect 18257 1897 18273 1931
rect 18207 1881 18273 1897
rect 18325 1931 18391 1947
rect 18325 1897 18341 1931
rect 18375 1897 18391 1931
rect 18325 1881 18391 1897
rect 18443 1931 18509 1947
rect 18443 1897 18459 1931
rect 18493 1897 18509 1931
rect 18443 1881 18509 1897
rect 18561 1931 18627 1947
rect 18561 1897 18577 1931
rect 18611 1897 18627 1931
rect 18561 1881 18627 1897
rect 18679 1931 18745 1947
rect 18679 1897 18695 1931
rect 18729 1897 18745 1931
rect 18679 1881 18745 1897
rect 18797 1931 18863 1947
rect 18797 1897 18813 1931
rect 18847 1897 18863 1931
rect 18797 1881 18863 1897
rect 18915 1931 18981 1947
rect 18915 1897 18931 1931
rect 18965 1897 18981 1931
rect 18915 1881 18981 1897
rect 19033 1931 19099 1947
rect 19033 1897 19049 1931
rect 19083 1897 19099 1931
rect 19033 1881 19099 1897
rect 19151 1931 19217 1947
rect 19151 1897 19167 1931
rect 19201 1897 19217 1931
rect 19151 1881 19217 1897
rect 19269 1931 19335 1947
rect 19269 1897 19285 1931
rect 19319 1897 19335 1931
rect 19269 1881 19335 1897
rect 19387 1931 19453 1947
rect 19387 1897 19403 1931
rect 19437 1897 19453 1931
rect 19387 1881 19453 1897
rect 19505 1931 19571 1947
rect 19505 1897 19521 1931
rect 19555 1897 19571 1931
rect 19505 1881 19571 1897
rect 19623 1931 19689 1947
rect 19623 1897 19639 1931
rect 19673 1897 19689 1931
rect 19623 1881 19689 1897
rect 19741 1931 19807 1947
rect 19741 1897 19757 1931
rect 19791 1897 19807 1931
rect 19741 1881 19807 1897
rect 19859 1931 19925 1947
rect 19859 1897 19875 1931
rect 19909 1897 19925 1931
rect 19859 1881 19925 1897
rect 19977 1931 20043 1947
rect 19977 1897 19993 1931
rect 20027 1897 20043 1931
rect 19977 1881 20043 1897
rect 20095 1931 20161 1947
rect 20095 1897 20111 1931
rect 20145 1897 20161 1931
rect 20095 1881 20161 1897
rect 20213 1931 20279 1947
rect 20213 1897 20229 1931
rect 20263 1897 20279 1931
rect 20213 1881 20279 1897
rect 20331 1931 20397 1947
rect 20331 1897 20347 1931
rect 20381 1897 20397 1931
rect 20331 1881 20397 1897
rect 20449 1931 20515 1947
rect 20449 1897 20465 1931
rect 20499 1897 20515 1931
rect 20449 1881 20515 1897
rect 20567 1931 20633 1947
rect 20567 1897 20583 1931
rect 20617 1897 20633 1931
rect 20567 1881 20633 1897
rect 20685 1931 20751 1947
rect 20685 1897 20701 1931
rect 20735 1897 20751 1931
rect 20685 1881 20751 1897
rect 20803 1931 20869 1947
rect 20803 1897 20819 1931
rect 20853 1897 20869 1931
rect 20803 1881 20869 1897
rect 20921 1931 20987 1947
rect 20921 1897 20937 1931
rect 20971 1897 20987 1931
rect 20921 1881 20987 1897
rect 21039 1931 21105 1947
rect 21039 1897 21055 1931
rect 21089 1897 21105 1931
rect 21039 1881 21105 1897
rect 21157 1931 21223 1947
rect 21157 1897 21173 1931
rect 21207 1897 21223 1931
rect 21157 1881 21223 1897
rect 21275 1931 21341 1947
rect 21275 1897 21291 1931
rect 21325 1897 21341 1931
rect 21275 1881 21341 1897
rect 1451 -148 1517 -132
rect 1451 -182 1467 -148
rect 1501 -182 1517 -148
rect 1333 -240 1399 -198
rect 1451 -256 1517 -182
rect 1451 -290 1467 -256
rect 1501 -290 1517 -256
rect 1451 -306 1517 -290
rect 1569 -148 1635 -132
rect 1569 -182 1585 -148
rect 1619 -182 1635 -148
rect 1569 -256 1635 -182
rect 1569 -290 1585 -256
rect 1619 -290 1635 -256
rect 1569 -306 1635 -290
rect 1687 -148 1753 -132
rect 1687 -182 1703 -148
rect 1737 -182 1753 -148
rect 1687 -256 1753 -182
rect 1687 -290 1703 -256
rect 1737 -290 1753 -256
rect 1687 -306 1753 -290
rect 1805 -148 1871 -132
rect 1805 -182 1821 -148
rect 1855 -182 1871 -148
rect 1805 -256 1871 -182
rect 1805 -290 1821 -256
rect 1855 -290 1871 -256
rect 1805 -306 1871 -290
rect 1923 -148 1989 -132
rect 1923 -182 1939 -148
rect 1973 -182 1989 -148
rect 1923 -256 1989 -182
rect 1923 -290 1939 -256
rect 1973 -290 1989 -256
rect 1923 -306 1989 -290
rect 2041 -148 2107 -132
rect 2041 -182 2057 -148
rect 2091 -182 2107 -148
rect 2041 -256 2107 -182
rect 2041 -290 2057 -256
rect 2091 -290 2107 -256
rect 2041 -306 2107 -290
rect 2159 -148 2225 -132
rect 2159 -182 2175 -148
rect 2209 -182 2225 -148
rect 2159 -256 2225 -182
rect 2159 -290 2175 -256
rect 2209 -290 2225 -256
rect 2159 -306 2225 -290
rect 2277 -148 2343 -132
rect 2277 -182 2293 -148
rect 2327 -182 2343 -148
rect 2277 -256 2343 -182
rect 2277 -290 2293 -256
rect 2327 -290 2343 -256
rect 2277 -306 2343 -290
rect 2395 -148 2461 -132
rect 2395 -182 2411 -148
rect 2445 -182 2461 -148
rect 2395 -256 2461 -182
rect 2395 -290 2411 -256
rect 2445 -290 2461 -256
rect 2395 -306 2461 -290
rect 2513 -148 2579 -132
rect 2513 -182 2529 -148
rect 2563 -182 2579 -148
rect 2513 -256 2579 -182
rect 2513 -290 2529 -256
rect 2563 -290 2579 -256
rect 2513 -306 2579 -290
rect 2631 -148 2697 -132
rect 2631 -182 2647 -148
rect 2681 -182 2697 -148
rect 2631 -256 2697 -182
rect 2631 -290 2647 -256
rect 2681 -290 2697 -256
rect 2631 -306 2697 -290
rect 2749 -148 2815 -132
rect 2749 -182 2765 -148
rect 2799 -182 2815 -148
rect 2749 -256 2815 -182
rect 2749 -290 2765 -256
rect 2799 -290 2815 -256
rect 2749 -306 2815 -290
rect 2867 -148 2933 -132
rect 2867 -182 2883 -148
rect 2917 -182 2933 -148
rect 2867 -256 2933 -182
rect 2867 -290 2883 -256
rect 2917 -290 2933 -256
rect 2867 -306 2933 -290
rect 2985 -148 3051 -132
rect 2985 -182 3001 -148
rect 3035 -182 3051 -148
rect 2985 -256 3051 -182
rect 2985 -290 3001 -256
rect 3035 -290 3051 -256
rect 2985 -306 3051 -290
rect 3103 -148 3169 -132
rect 3103 -182 3119 -148
rect 3153 -182 3169 -148
rect 3103 -256 3169 -182
rect 3103 -290 3119 -256
rect 3153 -290 3169 -256
rect 3103 -306 3169 -290
rect 3221 -148 3287 -132
rect 3221 -182 3237 -148
rect 3271 -182 3287 -148
rect 3221 -256 3287 -182
rect 3221 -290 3237 -256
rect 3271 -290 3287 -256
rect 3221 -306 3287 -290
rect 3339 -148 3405 -132
rect 3339 -182 3355 -148
rect 3389 -182 3405 -148
rect 3339 -256 3405 -182
rect 3339 -290 3355 -256
rect 3389 -290 3405 -256
rect 3339 -306 3405 -290
rect 3457 -148 3523 -132
rect 3457 -182 3473 -148
rect 3507 -182 3523 -148
rect 3457 -256 3523 -182
rect 3457 -290 3473 -256
rect 3507 -290 3523 -256
rect 3457 -306 3523 -290
rect 3575 -148 3641 -132
rect 3575 -182 3591 -148
rect 3625 -182 3641 -148
rect 3575 -256 3641 -182
rect 3575 -290 3591 -256
rect 3625 -290 3641 -256
rect 3575 -306 3641 -290
rect 3693 -148 3759 -132
rect 3693 -182 3709 -148
rect 3743 -182 3759 -148
rect 3693 -256 3759 -182
rect 3693 -290 3709 -256
rect 3743 -290 3759 -256
rect 3693 -306 3759 -290
rect 3811 -148 3877 -132
rect 3811 -182 3827 -148
rect 3861 -182 3877 -148
rect 3811 -256 3877 -182
rect 3811 -290 3827 -256
rect 3861 -290 3877 -256
rect 3811 -306 3877 -290
rect 3929 -148 3995 -132
rect 3929 -182 3945 -148
rect 3979 -182 3995 -148
rect 3929 -256 3995 -182
rect 3929 -290 3945 -256
rect 3979 -290 3995 -256
rect 3929 -306 3995 -290
rect 4047 -148 4113 -132
rect 4047 -182 4063 -148
rect 4097 -182 4113 -148
rect 4047 -256 4113 -182
rect 4047 -290 4063 -256
rect 4097 -290 4113 -256
rect 4047 -306 4113 -290
rect 4165 -148 4231 -132
rect 4165 -182 4181 -148
rect 4215 -182 4231 -148
rect 4165 -256 4231 -182
rect 4165 -290 4181 -256
rect 4215 -290 4231 -256
rect 4165 -306 4231 -290
rect 4283 -148 4349 -132
rect 4283 -182 4299 -148
rect 4333 -182 4349 -148
rect 4283 -256 4349 -182
rect 4283 -290 4299 -256
rect 4333 -290 4349 -256
rect 4283 -306 4349 -290
rect 4401 -148 4467 -132
rect 4401 -182 4417 -148
rect 4451 -182 4467 -148
rect 4401 -256 4467 -182
rect 4401 -290 4417 -256
rect 4451 -290 4467 -256
rect 4401 -306 4467 -290
rect 4519 -148 4585 -132
rect 4519 -182 4535 -148
rect 4569 -182 4585 -148
rect 4519 -256 4585 -182
rect 4519 -290 4535 -256
rect 4569 -290 4585 -256
rect 4519 -306 4585 -290
rect 4637 -148 4703 -132
rect 4637 -182 4653 -148
rect 4687 -182 4703 -148
rect 4637 -256 4703 -182
rect 4637 -290 4653 -256
rect 4687 -290 4703 -256
rect 4637 -306 4703 -290
rect 4755 -148 4821 -132
rect 4755 -182 4771 -148
rect 4805 -182 4821 -148
rect 4755 -256 4821 -182
rect 4755 -290 4771 -256
rect 4805 -290 4821 -256
rect 4755 -306 4821 -290
rect 4873 -148 4939 -132
rect 4873 -182 4889 -148
rect 4923 -182 4939 -148
rect 4873 -256 4939 -182
rect 4873 -290 4889 -256
rect 4923 -290 4939 -256
rect 4873 -306 4939 -290
rect 4991 -148 5057 -132
rect 4991 -182 5007 -148
rect 5041 -182 5057 -148
rect 4991 -256 5057 -182
rect 4991 -290 5007 -256
rect 5041 -290 5057 -256
rect 4991 -306 5057 -290
rect 5109 -148 5175 -132
rect 5109 -182 5125 -148
rect 5159 -182 5175 -148
rect 5109 -256 5175 -182
rect 5109 -290 5125 -256
rect 5159 -290 5175 -256
rect 5109 -306 5175 -290
rect 5227 -148 5293 -132
rect 5227 -182 5243 -148
rect 5277 -182 5293 -148
rect 5227 -256 5293 -182
rect 5227 -290 5243 -256
rect 5277 -290 5293 -256
rect 5227 -306 5293 -290
rect 5345 -148 5411 -132
rect 5345 -182 5361 -148
rect 5395 -182 5411 -148
rect 5345 -256 5411 -182
rect 5345 -290 5361 -256
rect 5395 -290 5411 -256
rect 5345 -306 5411 -290
rect 5463 -148 5529 -132
rect 5463 -182 5479 -148
rect 5513 -182 5529 -148
rect 5463 -256 5529 -182
rect 5463 -290 5479 -256
rect 5513 -290 5529 -256
rect 5463 -306 5529 -290
rect 5581 -148 5647 -132
rect 5581 -182 5597 -148
rect 5631 -182 5647 -148
rect 5581 -256 5647 -182
rect 5581 -290 5597 -256
rect 5631 -290 5647 -256
rect 5581 -306 5647 -290
rect 5699 -148 5765 -132
rect 5699 -182 5715 -148
rect 5749 -182 5765 -148
rect 5699 -256 5765 -182
rect 5699 -290 5715 -256
rect 5749 -290 5765 -256
rect 5699 -306 5765 -290
rect 5817 -148 5883 -132
rect 5817 -182 5833 -148
rect 5867 -182 5883 -148
rect 5817 -256 5883 -182
rect 5817 -290 5833 -256
rect 5867 -290 5883 -256
rect 5817 -306 5883 -290
rect 5935 -148 6001 -132
rect 5935 -182 5951 -148
rect 5985 -182 6001 -148
rect 5935 -256 6001 -182
rect 5935 -290 5951 -256
rect 5985 -290 6001 -256
rect 5935 -306 6001 -290
rect 6053 -148 6119 -132
rect 6053 -182 6069 -148
rect 6103 -182 6119 -148
rect 6053 -256 6119 -182
rect 6053 -290 6069 -256
rect 6103 -290 6119 -256
rect 6053 -306 6119 -290
rect 6171 -148 6237 -132
rect 6171 -182 6187 -148
rect 6221 -182 6237 -148
rect 6171 -256 6237 -182
rect 6171 -290 6187 -256
rect 6221 -290 6237 -256
rect 6171 -306 6237 -290
rect 6289 -148 6355 -132
rect 6289 -182 6305 -148
rect 6339 -182 6355 -148
rect 6289 -256 6355 -182
rect 6289 -290 6305 -256
rect 6339 -290 6355 -256
rect 6289 -306 6355 -290
rect 6407 -148 6473 -132
rect 6407 -182 6423 -148
rect 6457 -182 6473 -148
rect 6407 -256 6473 -182
rect 6407 -290 6423 -256
rect 6457 -290 6473 -256
rect 6407 -306 6473 -290
rect 6525 -148 6591 -132
rect 6525 -182 6541 -148
rect 6575 -182 6591 -148
rect 6525 -256 6591 -182
rect 6525 -290 6541 -256
rect 6575 -290 6591 -256
rect 6525 -306 6591 -290
rect 6643 -148 6709 -132
rect 6643 -182 6659 -148
rect 6693 -182 6709 -148
rect 6643 -256 6709 -182
rect 6643 -290 6659 -256
rect 6693 -290 6709 -256
rect 6643 -306 6709 -290
rect 6761 -148 6827 -132
rect 6761 -182 6777 -148
rect 6811 -182 6827 -148
rect 6761 -256 6827 -182
rect 6761 -290 6777 -256
rect 6811 -290 6827 -256
rect 6761 -306 6827 -290
rect 6879 -148 6945 -132
rect 6879 -182 6895 -148
rect 6929 -182 6945 -148
rect 6879 -256 6945 -182
rect 6879 -290 6895 -256
rect 6929 -290 6945 -256
rect 6879 -306 6945 -290
rect 6997 -148 7063 -132
rect 6997 -182 7013 -148
rect 7047 -182 7063 -148
rect 6997 -256 7063 -182
rect 6997 -290 7013 -256
rect 7047 -290 7063 -256
rect 6997 -306 7063 -290
rect 7115 -148 7181 -132
rect 7115 -182 7131 -148
rect 7165 -182 7181 -148
rect 7115 -256 7181 -182
rect 7115 -290 7131 -256
rect 7165 -290 7181 -256
rect 7115 -306 7181 -290
rect 1333 -1916 1399 -1900
rect 1333 -1950 1349 -1916
rect 1383 -1950 1399 -1916
rect 1333 -2024 1399 -1950
rect 1333 -2058 1349 -2024
rect 1383 -2058 1399 -2024
rect 1333 -2074 1399 -2058
rect 1451 -1916 1517 -1900
rect 1451 -1950 1467 -1916
rect 1501 -1950 1517 -1916
rect 1451 -2024 1517 -1950
rect 1451 -2058 1467 -2024
rect 1501 -2058 1517 -2024
rect 1451 -2074 1517 -2058
rect 1569 -1916 1635 -1900
rect 1569 -1950 1585 -1916
rect 1619 -1950 1635 -1916
rect 1569 -2024 1635 -1950
rect 1569 -2058 1585 -2024
rect 1619 -2058 1635 -2024
rect 1569 -2074 1635 -2058
rect 1687 -1916 1753 -1900
rect 1687 -1950 1703 -1916
rect 1737 -1950 1753 -1916
rect 1687 -2024 1753 -1950
rect 1687 -2058 1703 -2024
rect 1737 -2058 1753 -2024
rect 1687 -2074 1753 -2058
rect 1805 -1916 1871 -1900
rect 1805 -1950 1821 -1916
rect 1855 -1950 1871 -1916
rect 1805 -2024 1871 -1950
rect 1805 -2058 1821 -2024
rect 1855 -2058 1871 -2024
rect 1805 -2074 1871 -2058
rect 1923 -1916 1989 -1900
rect 1923 -1950 1939 -1916
rect 1973 -1950 1989 -1916
rect 1923 -2024 1989 -1950
rect 1923 -2058 1939 -2024
rect 1973 -2058 1989 -2024
rect 1923 -2074 1989 -2058
rect 2041 -1916 2107 -1900
rect 2041 -1950 2057 -1916
rect 2091 -1950 2107 -1916
rect 2041 -2024 2107 -1950
rect 2041 -2058 2057 -2024
rect 2091 -2058 2107 -2024
rect 2041 -2074 2107 -2058
rect 2159 -1916 2225 -1900
rect 2159 -1950 2175 -1916
rect 2209 -1950 2225 -1916
rect 2159 -2024 2225 -1950
rect 2159 -2058 2175 -2024
rect 2209 -2058 2225 -2024
rect 2159 -2074 2225 -2058
rect 2277 -1916 2343 -1900
rect 2277 -1950 2293 -1916
rect 2327 -1950 2343 -1916
rect 2277 -2024 2343 -1950
rect 2277 -2058 2293 -2024
rect 2327 -2058 2343 -2024
rect 2277 -2074 2343 -2058
rect 2395 -1916 2461 -1900
rect 2395 -1950 2411 -1916
rect 2445 -1950 2461 -1916
rect 2395 -2024 2461 -1950
rect 2395 -2058 2411 -2024
rect 2445 -2058 2461 -2024
rect 2395 -2074 2461 -2058
rect 2513 -1916 2579 -1900
rect 2513 -1950 2529 -1916
rect 2563 -1950 2579 -1916
rect 2513 -2024 2579 -1950
rect 2513 -2058 2529 -2024
rect 2563 -2058 2579 -2024
rect 2513 -2074 2579 -2058
rect 2631 -1916 2697 -1900
rect 2631 -1950 2647 -1916
rect 2681 -1950 2697 -1916
rect 2631 -2024 2697 -1950
rect 2631 -2058 2647 -2024
rect 2681 -2058 2697 -2024
rect 2631 -2074 2697 -2058
rect 2749 -1916 2815 -1900
rect 2749 -1950 2765 -1916
rect 2799 -1950 2815 -1916
rect 2749 -2024 2815 -1950
rect 2749 -2058 2765 -2024
rect 2799 -2058 2815 -2024
rect 2749 -2074 2815 -2058
rect 2867 -1916 2933 -1900
rect 2867 -1950 2883 -1916
rect 2917 -1950 2933 -1916
rect 2867 -2024 2933 -1950
rect 2867 -2058 2883 -2024
rect 2917 -2058 2933 -2024
rect 2867 -2074 2933 -2058
rect 2985 -1916 3051 -1900
rect 2985 -1950 3001 -1916
rect 3035 -1950 3051 -1916
rect 2985 -2024 3051 -1950
rect 2985 -2058 3001 -2024
rect 3035 -2058 3051 -2024
rect 2985 -2074 3051 -2058
rect 3103 -1916 3169 -1900
rect 3103 -1950 3119 -1916
rect 3153 -1950 3169 -1916
rect 3103 -2024 3169 -1950
rect 3103 -2058 3119 -2024
rect 3153 -2058 3169 -2024
rect 3103 -2074 3169 -2058
rect 3221 -1916 3287 -1900
rect 3221 -1950 3237 -1916
rect 3271 -1950 3287 -1916
rect 3221 -2024 3287 -1950
rect 3221 -2058 3237 -2024
rect 3271 -2058 3287 -2024
rect 3221 -2074 3287 -2058
rect 3339 -1916 3405 -1900
rect 3339 -1950 3355 -1916
rect 3389 -1950 3405 -1916
rect 3339 -2024 3405 -1950
rect 3339 -2058 3355 -2024
rect 3389 -2058 3405 -2024
rect 3339 -2074 3405 -2058
rect 3457 -1916 3523 -1900
rect 3457 -1950 3473 -1916
rect 3507 -1950 3523 -1916
rect 3457 -2024 3523 -1950
rect 3457 -2058 3473 -2024
rect 3507 -2058 3523 -2024
rect 3457 -2074 3523 -2058
rect 3575 -1916 3641 -1900
rect 3575 -1950 3591 -1916
rect 3625 -1950 3641 -1916
rect 3575 -2024 3641 -1950
rect 3575 -2058 3591 -2024
rect 3625 -2058 3641 -2024
rect 3575 -2074 3641 -2058
rect 3693 -1916 3759 -1900
rect 3693 -1950 3709 -1916
rect 3743 -1950 3759 -1916
rect 3693 -2024 3759 -1950
rect 3693 -2058 3709 -2024
rect 3743 -2058 3759 -2024
rect 3693 -2074 3759 -2058
rect 3811 -1916 3877 -1900
rect 3811 -1950 3827 -1916
rect 3861 -1950 3877 -1916
rect 3811 -2024 3877 -1950
rect 3811 -2058 3827 -2024
rect 3861 -2058 3877 -2024
rect 3811 -2074 3877 -2058
rect 3929 -1916 3995 -1900
rect 3929 -1950 3945 -1916
rect 3979 -1950 3995 -1916
rect 3929 -2024 3995 -1950
rect 3929 -2058 3945 -2024
rect 3979 -2058 3995 -2024
rect 3929 -2074 3995 -2058
rect 4047 -1916 4113 -1900
rect 4047 -1950 4063 -1916
rect 4097 -1950 4113 -1916
rect 4047 -2024 4113 -1950
rect 4047 -2058 4063 -2024
rect 4097 -2058 4113 -2024
rect 4047 -2074 4113 -2058
rect 4165 -1916 4231 -1900
rect 4165 -1950 4181 -1916
rect 4215 -1950 4231 -1916
rect 4165 -2024 4231 -1950
rect 4165 -2058 4181 -2024
rect 4215 -2058 4231 -2024
rect 4165 -2074 4231 -2058
rect 4283 -1916 4349 -1900
rect 4283 -1950 4299 -1916
rect 4333 -1950 4349 -1916
rect 4283 -2024 4349 -1950
rect 4283 -2058 4299 -2024
rect 4333 -2058 4349 -2024
rect 4283 -2074 4349 -2058
rect 4401 -1916 4467 -1900
rect 4401 -1950 4417 -1916
rect 4451 -1950 4467 -1916
rect 4401 -2024 4467 -1950
rect 4401 -2058 4417 -2024
rect 4451 -2058 4467 -2024
rect 4401 -2074 4467 -2058
rect 4519 -1916 4585 -1900
rect 4519 -1950 4535 -1916
rect 4569 -1950 4585 -1916
rect 4519 -2024 4585 -1950
rect 4519 -2058 4535 -2024
rect 4569 -2058 4585 -2024
rect 4519 -2074 4585 -2058
rect 4637 -1916 4703 -1900
rect 4637 -1950 4653 -1916
rect 4687 -1950 4703 -1916
rect 4637 -2024 4703 -1950
rect 4637 -2058 4653 -2024
rect 4687 -2058 4703 -2024
rect 4637 -2074 4703 -2058
rect 4755 -1916 4821 -1900
rect 4755 -1950 4771 -1916
rect 4805 -1950 4821 -1916
rect 4755 -2024 4821 -1950
rect 4755 -2058 4771 -2024
rect 4805 -2058 4821 -2024
rect 4755 -2074 4821 -2058
rect 4873 -1916 4939 -1900
rect 4873 -1950 4889 -1916
rect 4923 -1950 4939 -1916
rect 4873 -2024 4939 -1950
rect 4873 -2058 4889 -2024
rect 4923 -2058 4939 -2024
rect 4873 -2074 4939 -2058
rect 4991 -1916 5057 -1900
rect 4991 -1950 5007 -1916
rect 5041 -1950 5057 -1916
rect 4991 -2024 5057 -1950
rect 4991 -2058 5007 -2024
rect 5041 -2058 5057 -2024
rect 4991 -2074 5057 -2058
rect 5109 -1916 5175 -1900
rect 5109 -1950 5125 -1916
rect 5159 -1950 5175 -1916
rect 5109 -2024 5175 -1950
rect 5109 -2058 5125 -2024
rect 5159 -2058 5175 -2024
rect 5109 -2074 5175 -2058
rect 5227 -1916 5293 -1900
rect 5227 -1950 5243 -1916
rect 5277 -1950 5293 -1916
rect 5227 -2024 5293 -1950
rect 5227 -2058 5243 -2024
rect 5277 -2058 5293 -2024
rect 5227 -2074 5293 -2058
rect 5345 -1916 5411 -1900
rect 5345 -1950 5361 -1916
rect 5395 -1950 5411 -1916
rect 5345 -2024 5411 -1950
rect 5345 -2058 5361 -2024
rect 5395 -2058 5411 -2024
rect 5345 -2074 5411 -2058
rect 5463 -1916 5529 -1900
rect 5463 -1950 5479 -1916
rect 5513 -1950 5529 -1916
rect 5463 -2024 5529 -1950
rect 5463 -2058 5479 -2024
rect 5513 -2058 5529 -2024
rect 5463 -2074 5529 -2058
rect 5581 -1916 5647 -1900
rect 5581 -1950 5597 -1916
rect 5631 -1950 5647 -1916
rect 5581 -2024 5647 -1950
rect 5581 -2058 5597 -2024
rect 5631 -2058 5647 -2024
rect 5581 -2074 5647 -2058
rect 5699 -1916 5765 -1900
rect 5699 -1950 5715 -1916
rect 5749 -1950 5765 -1916
rect 5699 -2024 5765 -1950
rect 5699 -2058 5715 -2024
rect 5749 -2058 5765 -2024
rect 5699 -2074 5765 -2058
rect 5817 -1916 5883 -1900
rect 5817 -1950 5833 -1916
rect 5867 -1950 5883 -1916
rect 5817 -2024 5883 -1950
rect 5817 -2058 5833 -2024
rect 5867 -2058 5883 -2024
rect 5817 -2074 5883 -2058
rect 5935 -1916 6001 -1900
rect 5935 -1950 5951 -1916
rect 5985 -1950 6001 -1916
rect 5935 -2024 6001 -1950
rect 5935 -2058 5951 -2024
rect 5985 -2058 6001 -2024
rect 5935 -2074 6001 -2058
rect 6053 -1916 6119 -1900
rect 6053 -1950 6069 -1916
rect 6103 -1950 6119 -1916
rect 6053 -2024 6119 -1950
rect 6053 -2058 6069 -2024
rect 6103 -2058 6119 -2024
rect 6053 -2074 6119 -2058
rect 6171 -1916 6237 -1900
rect 6171 -1950 6187 -1916
rect 6221 -1950 6237 -1916
rect 6171 -2024 6237 -1950
rect 6171 -2058 6187 -2024
rect 6221 -2058 6237 -2024
rect 6171 -2074 6237 -2058
rect 6289 -1916 6355 -1900
rect 6289 -1950 6305 -1916
rect 6339 -1950 6355 -1916
rect 6289 -2024 6355 -1950
rect 6289 -2058 6305 -2024
rect 6339 -2058 6355 -2024
rect 6289 -2074 6355 -2058
rect 6407 -1916 6473 -1900
rect 6407 -1950 6423 -1916
rect 6457 -1950 6473 -1916
rect 6407 -2024 6473 -1950
rect 6407 -2058 6423 -2024
rect 6457 -2058 6473 -2024
rect 6407 -2074 6473 -2058
rect 6525 -1916 6591 -1900
rect 6525 -1950 6541 -1916
rect 6575 -1950 6591 -1916
rect 6525 -2024 6591 -1950
rect 6525 -2058 6541 -2024
rect 6575 -2058 6591 -2024
rect 6525 -2074 6591 -2058
rect 6643 -1916 6709 -1900
rect 6643 -1950 6659 -1916
rect 6693 -1950 6709 -1916
rect 6643 -2024 6709 -1950
rect 6643 -2058 6659 -2024
rect 6693 -2058 6709 -2024
rect 6643 -2074 6709 -2058
rect 6761 -1916 6827 -1900
rect 6761 -1950 6777 -1916
rect 6811 -1950 6827 -1916
rect 6761 -2024 6827 -1950
rect 6761 -2058 6777 -2024
rect 6811 -2058 6827 -2024
rect 6761 -2074 6827 -2058
rect 6879 -1916 6945 -1900
rect 6879 -1950 6895 -1916
rect 6929 -1950 6945 -1916
rect 6879 -2024 6945 -1950
rect 6879 -2058 6895 -2024
rect 6929 -2058 6945 -2024
rect 6879 -2074 6945 -2058
rect 6997 -1916 7063 -1900
rect 6997 -1950 7013 -1916
rect 7047 -1950 7063 -1916
rect 6997 -2024 7063 -1950
rect 6997 -2058 7013 -2024
rect 7047 -2058 7063 -2024
rect 6997 -2074 7063 -2058
rect 7115 -1916 7181 -1900
rect 7115 -1950 7131 -1916
rect 7165 -1950 7181 -1916
rect 7115 -2024 7181 -1950
rect 7115 -2058 7131 -2024
rect 7165 -2058 7181 -2024
rect 7115 -2074 7181 -2058
rect 1333 -3684 1399 -3668
rect 1333 -3718 1349 -3684
rect 1383 -3718 1399 -3684
rect 1333 -3792 1399 -3718
rect 1333 -3826 1349 -3792
rect 1383 -3826 1399 -3792
rect 1333 -3842 1399 -3826
rect 1451 -3684 1517 -3668
rect 1451 -3718 1467 -3684
rect 1501 -3718 1517 -3684
rect 1451 -3792 1517 -3718
rect 1451 -3826 1467 -3792
rect 1501 -3826 1517 -3792
rect 1451 -3842 1517 -3826
rect 1569 -3684 1635 -3668
rect 1569 -3718 1585 -3684
rect 1619 -3718 1635 -3684
rect 1569 -3792 1635 -3718
rect 1569 -3826 1585 -3792
rect 1619 -3826 1635 -3792
rect 1569 -3842 1635 -3826
rect 1687 -3684 1753 -3668
rect 1687 -3718 1703 -3684
rect 1737 -3718 1753 -3684
rect 1687 -3792 1753 -3718
rect 1687 -3826 1703 -3792
rect 1737 -3826 1753 -3792
rect 1687 -3842 1753 -3826
rect 1805 -3684 1871 -3668
rect 1805 -3718 1821 -3684
rect 1855 -3718 1871 -3684
rect 1805 -3792 1871 -3718
rect 1805 -3826 1821 -3792
rect 1855 -3826 1871 -3792
rect 1805 -3842 1871 -3826
rect 1923 -3684 1989 -3668
rect 1923 -3718 1939 -3684
rect 1973 -3718 1989 -3684
rect 1923 -3792 1989 -3718
rect 1923 -3826 1939 -3792
rect 1973 -3826 1989 -3792
rect 1923 -3842 1989 -3826
rect 2041 -3684 2107 -3668
rect 2041 -3718 2057 -3684
rect 2091 -3718 2107 -3684
rect 2041 -3792 2107 -3718
rect 2041 -3826 2057 -3792
rect 2091 -3826 2107 -3792
rect 2041 -3842 2107 -3826
rect 2159 -3684 2225 -3668
rect 2159 -3718 2175 -3684
rect 2209 -3718 2225 -3684
rect 2159 -3792 2225 -3718
rect 2159 -3826 2175 -3792
rect 2209 -3826 2225 -3792
rect 2159 -3842 2225 -3826
rect 2277 -3684 2343 -3668
rect 2277 -3718 2293 -3684
rect 2327 -3718 2343 -3684
rect 2277 -3792 2343 -3718
rect 2277 -3826 2293 -3792
rect 2327 -3826 2343 -3792
rect 2277 -3842 2343 -3826
rect 2395 -3684 2461 -3668
rect 2395 -3718 2411 -3684
rect 2445 -3718 2461 -3684
rect 2395 -3792 2461 -3718
rect 2395 -3826 2411 -3792
rect 2445 -3826 2461 -3792
rect 2395 -3842 2461 -3826
rect 2513 -3684 2579 -3668
rect 2513 -3718 2529 -3684
rect 2563 -3718 2579 -3684
rect 2513 -3792 2579 -3718
rect 2513 -3826 2529 -3792
rect 2563 -3826 2579 -3792
rect 2513 -3842 2579 -3826
rect 2631 -3684 2697 -3668
rect 2631 -3718 2647 -3684
rect 2681 -3718 2697 -3684
rect 2631 -3792 2697 -3718
rect 2631 -3826 2647 -3792
rect 2681 -3826 2697 -3792
rect 2631 -3842 2697 -3826
rect 2749 -3684 2815 -3668
rect 2749 -3718 2765 -3684
rect 2799 -3718 2815 -3684
rect 2749 -3792 2815 -3718
rect 2749 -3826 2765 -3792
rect 2799 -3826 2815 -3792
rect 2749 -3842 2815 -3826
rect 2867 -3684 2933 -3668
rect 2867 -3718 2883 -3684
rect 2917 -3718 2933 -3684
rect 2867 -3792 2933 -3718
rect 2867 -3826 2883 -3792
rect 2917 -3826 2933 -3792
rect 2867 -3842 2933 -3826
rect 2985 -3684 3051 -3668
rect 2985 -3718 3001 -3684
rect 3035 -3718 3051 -3684
rect 2985 -3792 3051 -3718
rect 2985 -3826 3001 -3792
rect 3035 -3826 3051 -3792
rect 2985 -3842 3051 -3826
rect 3103 -3684 3169 -3668
rect 3103 -3718 3119 -3684
rect 3153 -3718 3169 -3684
rect 3103 -3792 3169 -3718
rect 3103 -3826 3119 -3792
rect 3153 -3826 3169 -3792
rect 3103 -3842 3169 -3826
rect 3221 -3684 3287 -3668
rect 3221 -3718 3237 -3684
rect 3271 -3718 3287 -3684
rect 3221 -3792 3287 -3718
rect 3221 -3826 3237 -3792
rect 3271 -3826 3287 -3792
rect 3221 -3842 3287 -3826
rect 3339 -3684 3405 -3668
rect 3339 -3718 3355 -3684
rect 3389 -3718 3405 -3684
rect 3339 -3792 3405 -3718
rect 3339 -3826 3355 -3792
rect 3389 -3826 3405 -3792
rect 3339 -3842 3405 -3826
rect 3457 -3684 3523 -3668
rect 3457 -3718 3473 -3684
rect 3507 -3718 3523 -3684
rect 3457 -3792 3523 -3718
rect 3457 -3826 3473 -3792
rect 3507 -3826 3523 -3792
rect 3457 -3842 3523 -3826
rect 3575 -3684 3641 -3668
rect 3575 -3718 3591 -3684
rect 3625 -3718 3641 -3684
rect 3575 -3792 3641 -3718
rect 3575 -3826 3591 -3792
rect 3625 -3826 3641 -3792
rect 3575 -3842 3641 -3826
rect 3693 -3684 3759 -3668
rect 3693 -3718 3709 -3684
rect 3743 -3718 3759 -3684
rect 3693 -3792 3759 -3718
rect 3693 -3826 3709 -3792
rect 3743 -3826 3759 -3792
rect 3693 -3842 3759 -3826
rect 3811 -3684 3877 -3668
rect 3811 -3718 3827 -3684
rect 3861 -3718 3877 -3684
rect 3811 -3792 3877 -3718
rect 3811 -3826 3827 -3792
rect 3861 -3826 3877 -3792
rect 3811 -3842 3877 -3826
rect 3929 -3684 3995 -3668
rect 3929 -3718 3945 -3684
rect 3979 -3718 3995 -3684
rect 3929 -3792 3995 -3718
rect 3929 -3826 3945 -3792
rect 3979 -3826 3995 -3792
rect 3929 -3842 3995 -3826
rect 4047 -3684 4113 -3668
rect 4047 -3718 4063 -3684
rect 4097 -3718 4113 -3684
rect 4047 -3792 4113 -3718
rect 4047 -3826 4063 -3792
rect 4097 -3826 4113 -3792
rect 4047 -3842 4113 -3826
rect 4165 -3684 4231 -3668
rect 4165 -3718 4181 -3684
rect 4215 -3718 4231 -3684
rect 4165 -3792 4231 -3718
rect 4165 -3826 4181 -3792
rect 4215 -3826 4231 -3792
rect 4165 -3842 4231 -3826
rect 4283 -3684 4349 -3668
rect 4283 -3718 4299 -3684
rect 4333 -3718 4349 -3684
rect 4283 -3792 4349 -3718
rect 4283 -3826 4299 -3792
rect 4333 -3826 4349 -3792
rect 4283 -3842 4349 -3826
rect 4401 -3684 4467 -3668
rect 4401 -3718 4417 -3684
rect 4451 -3718 4467 -3684
rect 4401 -3792 4467 -3718
rect 4401 -3826 4417 -3792
rect 4451 -3826 4467 -3792
rect 4401 -3842 4467 -3826
rect 4519 -3684 4585 -3668
rect 4519 -3718 4535 -3684
rect 4569 -3718 4585 -3684
rect 4519 -3792 4585 -3718
rect 4519 -3826 4535 -3792
rect 4569 -3826 4585 -3792
rect 4519 -3842 4585 -3826
rect 4637 -3684 4703 -3668
rect 4637 -3718 4653 -3684
rect 4687 -3718 4703 -3684
rect 4637 -3792 4703 -3718
rect 4637 -3826 4653 -3792
rect 4687 -3826 4703 -3792
rect 4637 -3842 4703 -3826
rect 4755 -3684 4821 -3668
rect 4755 -3718 4771 -3684
rect 4805 -3718 4821 -3684
rect 4755 -3792 4821 -3718
rect 4755 -3826 4771 -3792
rect 4805 -3826 4821 -3792
rect 4755 -3842 4821 -3826
rect 4873 -3684 4939 -3668
rect 4873 -3718 4889 -3684
rect 4923 -3718 4939 -3684
rect 4873 -3792 4939 -3718
rect 4873 -3826 4889 -3792
rect 4923 -3826 4939 -3792
rect 4873 -3842 4939 -3826
rect 4991 -3684 5057 -3668
rect 4991 -3718 5007 -3684
rect 5041 -3718 5057 -3684
rect 4991 -3792 5057 -3718
rect 4991 -3826 5007 -3792
rect 5041 -3826 5057 -3792
rect 4991 -3842 5057 -3826
rect 5109 -3684 5175 -3668
rect 5109 -3718 5125 -3684
rect 5159 -3718 5175 -3684
rect 5109 -3792 5175 -3718
rect 5109 -3826 5125 -3792
rect 5159 -3826 5175 -3792
rect 5109 -3842 5175 -3826
rect 5227 -3684 5293 -3668
rect 5227 -3718 5243 -3684
rect 5277 -3718 5293 -3684
rect 5227 -3792 5293 -3718
rect 5227 -3826 5243 -3792
rect 5277 -3826 5293 -3792
rect 5227 -3842 5293 -3826
rect 5345 -3684 5411 -3668
rect 5345 -3718 5361 -3684
rect 5395 -3718 5411 -3684
rect 5345 -3792 5411 -3718
rect 5345 -3826 5361 -3792
rect 5395 -3826 5411 -3792
rect 5345 -3842 5411 -3826
rect 5463 -3684 5529 -3668
rect 5463 -3718 5479 -3684
rect 5513 -3718 5529 -3684
rect 5463 -3792 5529 -3718
rect 5463 -3826 5479 -3792
rect 5513 -3826 5529 -3792
rect 5463 -3842 5529 -3826
rect 5581 -3684 5647 -3668
rect 5581 -3718 5597 -3684
rect 5631 -3718 5647 -3684
rect 5581 -3792 5647 -3718
rect 5581 -3826 5597 -3792
rect 5631 -3826 5647 -3792
rect 5581 -3842 5647 -3826
rect 5699 -3684 5765 -3668
rect 5699 -3718 5715 -3684
rect 5749 -3718 5765 -3684
rect 5699 -3792 5765 -3718
rect 5699 -3826 5715 -3792
rect 5749 -3826 5765 -3792
rect 5699 -3842 5765 -3826
rect 5817 -3684 5883 -3668
rect 5817 -3718 5833 -3684
rect 5867 -3718 5883 -3684
rect 5817 -3792 5883 -3718
rect 5817 -3826 5833 -3792
rect 5867 -3826 5883 -3792
rect 5817 -3842 5883 -3826
rect 5935 -3684 6001 -3668
rect 5935 -3718 5951 -3684
rect 5985 -3718 6001 -3684
rect 5935 -3792 6001 -3718
rect 5935 -3826 5951 -3792
rect 5985 -3826 6001 -3792
rect 5935 -3842 6001 -3826
rect 6053 -3684 6119 -3668
rect 6053 -3718 6069 -3684
rect 6103 -3718 6119 -3684
rect 6053 -3792 6119 -3718
rect 6053 -3826 6069 -3792
rect 6103 -3826 6119 -3792
rect 6053 -3842 6119 -3826
rect 6171 -3684 6237 -3668
rect 6171 -3718 6187 -3684
rect 6221 -3718 6237 -3684
rect 6171 -3792 6237 -3718
rect 6171 -3826 6187 -3792
rect 6221 -3826 6237 -3792
rect 6171 -3842 6237 -3826
rect 6289 -3684 6355 -3668
rect 6289 -3718 6305 -3684
rect 6339 -3718 6355 -3684
rect 6289 -3792 6355 -3718
rect 6289 -3826 6305 -3792
rect 6339 -3826 6355 -3792
rect 6289 -3842 6355 -3826
rect 6407 -3684 6473 -3668
rect 6407 -3718 6423 -3684
rect 6457 -3718 6473 -3684
rect 6407 -3792 6473 -3718
rect 6407 -3826 6423 -3792
rect 6457 -3826 6473 -3792
rect 6407 -3842 6473 -3826
rect 6525 -3684 6591 -3668
rect 6525 -3718 6541 -3684
rect 6575 -3718 6591 -3684
rect 6525 -3792 6591 -3718
rect 6525 -3826 6541 -3792
rect 6575 -3826 6591 -3792
rect 6525 -3842 6591 -3826
rect 6643 -3684 6709 -3668
rect 6643 -3718 6659 -3684
rect 6693 -3718 6709 -3684
rect 6643 -3792 6709 -3718
rect 6643 -3826 6659 -3792
rect 6693 -3826 6709 -3792
rect 6643 -3842 6709 -3826
rect 6761 -3684 6827 -3668
rect 6761 -3718 6777 -3684
rect 6811 -3718 6827 -3684
rect 6761 -3792 6827 -3718
rect 6761 -3826 6777 -3792
rect 6811 -3826 6827 -3792
rect 6761 -3842 6827 -3826
rect 6879 -3684 6945 -3668
rect 6879 -3718 6895 -3684
rect 6929 -3718 6945 -3684
rect 6879 -3792 6945 -3718
rect 6879 -3826 6895 -3792
rect 6929 -3826 6945 -3792
rect 6879 -3842 6945 -3826
rect 6997 -3684 7063 -3668
rect 6997 -3718 7013 -3684
rect 7047 -3718 7063 -3684
rect 6997 -3792 7063 -3718
rect 6997 -3826 7013 -3792
rect 7047 -3826 7063 -3792
rect 6997 -3842 7063 -3826
rect 7115 -3684 7181 -3668
rect 7115 -3718 7131 -3684
rect 7165 -3718 7181 -3684
rect 7115 -3792 7181 -3718
rect 7115 -3826 7131 -3792
rect 7165 -3826 7181 -3792
rect 7115 -3842 7181 -3826
rect 1333 -5452 1399 -5436
rect 1333 -5486 1349 -5452
rect 1383 -5486 1399 -5452
rect 1333 -5560 1399 -5486
rect 1333 -5594 1349 -5560
rect 1383 -5594 1399 -5560
rect 1333 -5610 1399 -5594
rect 1451 -5452 1517 -5436
rect 1451 -5486 1467 -5452
rect 1501 -5486 1517 -5452
rect 1451 -5560 1517 -5486
rect 1451 -5594 1467 -5560
rect 1501 -5594 1517 -5560
rect 1451 -5610 1517 -5594
rect 1569 -5452 1635 -5436
rect 1569 -5486 1585 -5452
rect 1619 -5486 1635 -5452
rect 1569 -5560 1635 -5486
rect 1569 -5594 1585 -5560
rect 1619 -5594 1635 -5560
rect 1569 -5610 1635 -5594
rect 1687 -5452 1753 -5436
rect 1687 -5486 1703 -5452
rect 1737 -5486 1753 -5452
rect 1687 -5560 1753 -5486
rect 1687 -5594 1703 -5560
rect 1737 -5594 1753 -5560
rect 1687 -5610 1753 -5594
rect 1805 -5452 1871 -5436
rect 1805 -5486 1821 -5452
rect 1855 -5486 1871 -5452
rect 1805 -5560 1871 -5486
rect 1805 -5594 1821 -5560
rect 1855 -5594 1871 -5560
rect 1805 -5610 1871 -5594
rect 1923 -5452 1989 -5436
rect 1923 -5486 1939 -5452
rect 1973 -5486 1989 -5452
rect 1923 -5560 1989 -5486
rect 1923 -5594 1939 -5560
rect 1973 -5594 1989 -5560
rect 1923 -5610 1989 -5594
rect 2041 -5452 2107 -5436
rect 2041 -5486 2057 -5452
rect 2091 -5486 2107 -5452
rect 2041 -5560 2107 -5486
rect 2041 -5594 2057 -5560
rect 2091 -5594 2107 -5560
rect 2041 -5610 2107 -5594
rect 2159 -5452 2225 -5436
rect 2159 -5486 2175 -5452
rect 2209 -5486 2225 -5452
rect 2159 -5560 2225 -5486
rect 2159 -5594 2175 -5560
rect 2209 -5594 2225 -5560
rect 2159 -5610 2225 -5594
rect 2277 -5452 2343 -5436
rect 2277 -5486 2293 -5452
rect 2327 -5486 2343 -5452
rect 2277 -5560 2343 -5486
rect 2277 -5594 2293 -5560
rect 2327 -5594 2343 -5560
rect 2277 -5610 2343 -5594
rect 2395 -5452 2461 -5436
rect 2395 -5486 2411 -5452
rect 2445 -5486 2461 -5452
rect 2395 -5560 2461 -5486
rect 2395 -5594 2411 -5560
rect 2445 -5594 2461 -5560
rect 2395 -5610 2461 -5594
rect 2513 -5452 2579 -5436
rect 2513 -5486 2529 -5452
rect 2563 -5486 2579 -5452
rect 2513 -5560 2579 -5486
rect 2513 -5594 2529 -5560
rect 2563 -5594 2579 -5560
rect 2513 -5610 2579 -5594
rect 2631 -5452 2697 -5436
rect 2631 -5486 2647 -5452
rect 2681 -5486 2697 -5452
rect 2631 -5560 2697 -5486
rect 2631 -5594 2647 -5560
rect 2681 -5594 2697 -5560
rect 2631 -5610 2697 -5594
rect 2749 -5452 2815 -5436
rect 2749 -5486 2765 -5452
rect 2799 -5486 2815 -5452
rect 2749 -5560 2815 -5486
rect 2749 -5594 2765 -5560
rect 2799 -5594 2815 -5560
rect 2749 -5610 2815 -5594
rect 2867 -5452 2933 -5436
rect 2867 -5486 2883 -5452
rect 2917 -5486 2933 -5452
rect 2867 -5560 2933 -5486
rect 2867 -5594 2883 -5560
rect 2917 -5594 2933 -5560
rect 2867 -5610 2933 -5594
rect 2985 -5452 3051 -5436
rect 2985 -5486 3001 -5452
rect 3035 -5486 3051 -5452
rect 2985 -5560 3051 -5486
rect 2985 -5594 3001 -5560
rect 3035 -5594 3051 -5560
rect 2985 -5610 3051 -5594
rect 3103 -5452 3169 -5436
rect 3103 -5486 3119 -5452
rect 3153 -5486 3169 -5452
rect 3103 -5560 3169 -5486
rect 3103 -5594 3119 -5560
rect 3153 -5594 3169 -5560
rect 3103 -5610 3169 -5594
rect 3221 -5452 3287 -5436
rect 3221 -5486 3237 -5452
rect 3271 -5486 3287 -5452
rect 3221 -5560 3287 -5486
rect 3221 -5594 3237 -5560
rect 3271 -5594 3287 -5560
rect 3221 -5610 3287 -5594
rect 3339 -5452 3405 -5436
rect 3339 -5486 3355 -5452
rect 3389 -5486 3405 -5452
rect 3339 -5560 3405 -5486
rect 3339 -5594 3355 -5560
rect 3389 -5594 3405 -5560
rect 3339 -5610 3405 -5594
rect 3457 -5452 3523 -5436
rect 3457 -5486 3473 -5452
rect 3507 -5486 3523 -5452
rect 3457 -5560 3523 -5486
rect 3457 -5594 3473 -5560
rect 3507 -5594 3523 -5560
rect 3457 -5610 3523 -5594
rect 3575 -5452 3641 -5436
rect 3575 -5486 3591 -5452
rect 3625 -5486 3641 -5452
rect 3575 -5560 3641 -5486
rect 3575 -5594 3591 -5560
rect 3625 -5594 3641 -5560
rect 3575 -5610 3641 -5594
rect 3693 -5452 3759 -5436
rect 3693 -5486 3709 -5452
rect 3743 -5486 3759 -5452
rect 3693 -5560 3759 -5486
rect 3693 -5594 3709 -5560
rect 3743 -5594 3759 -5560
rect 3693 -5610 3759 -5594
rect 3811 -5452 3877 -5436
rect 3811 -5486 3827 -5452
rect 3861 -5486 3877 -5452
rect 3811 -5560 3877 -5486
rect 3811 -5594 3827 -5560
rect 3861 -5594 3877 -5560
rect 3811 -5610 3877 -5594
rect 3929 -5452 3995 -5436
rect 3929 -5486 3945 -5452
rect 3979 -5486 3995 -5452
rect 3929 -5560 3995 -5486
rect 3929 -5594 3945 -5560
rect 3979 -5594 3995 -5560
rect 3929 -5610 3995 -5594
rect 4047 -5452 4113 -5436
rect 4047 -5486 4063 -5452
rect 4097 -5486 4113 -5452
rect 4047 -5560 4113 -5486
rect 4047 -5594 4063 -5560
rect 4097 -5594 4113 -5560
rect 4047 -5610 4113 -5594
rect 4165 -5452 4231 -5436
rect 4165 -5486 4181 -5452
rect 4215 -5486 4231 -5452
rect 4165 -5560 4231 -5486
rect 4165 -5594 4181 -5560
rect 4215 -5594 4231 -5560
rect 4165 -5610 4231 -5594
rect 4283 -5452 4349 -5436
rect 4283 -5486 4299 -5452
rect 4333 -5486 4349 -5452
rect 4283 -5560 4349 -5486
rect 4283 -5594 4299 -5560
rect 4333 -5594 4349 -5560
rect 4283 -5610 4349 -5594
rect 4401 -5452 4467 -5436
rect 4401 -5486 4417 -5452
rect 4451 -5486 4467 -5452
rect 4401 -5560 4467 -5486
rect 4401 -5594 4417 -5560
rect 4451 -5594 4467 -5560
rect 4401 -5610 4467 -5594
rect 4519 -5452 4585 -5436
rect 4519 -5486 4535 -5452
rect 4569 -5486 4585 -5452
rect 4519 -5560 4585 -5486
rect 4519 -5594 4535 -5560
rect 4569 -5594 4585 -5560
rect 4519 -5610 4585 -5594
rect 4637 -5452 4703 -5436
rect 4637 -5486 4653 -5452
rect 4687 -5486 4703 -5452
rect 4637 -5560 4703 -5486
rect 4637 -5594 4653 -5560
rect 4687 -5594 4703 -5560
rect 4637 -5610 4703 -5594
rect 4755 -5452 4821 -5436
rect 4755 -5486 4771 -5452
rect 4805 -5486 4821 -5452
rect 4755 -5560 4821 -5486
rect 4755 -5594 4771 -5560
rect 4805 -5594 4821 -5560
rect 4755 -5610 4821 -5594
rect 4873 -5452 4939 -5436
rect 4873 -5486 4889 -5452
rect 4923 -5486 4939 -5452
rect 4873 -5560 4939 -5486
rect 4873 -5594 4889 -5560
rect 4923 -5594 4939 -5560
rect 4873 -5610 4939 -5594
rect 4991 -5452 5057 -5436
rect 4991 -5486 5007 -5452
rect 5041 -5486 5057 -5452
rect 4991 -5560 5057 -5486
rect 4991 -5594 5007 -5560
rect 5041 -5594 5057 -5560
rect 4991 -5610 5057 -5594
rect 5109 -5452 5175 -5436
rect 5109 -5486 5125 -5452
rect 5159 -5486 5175 -5452
rect 5109 -5560 5175 -5486
rect 5109 -5594 5125 -5560
rect 5159 -5594 5175 -5560
rect 5109 -5610 5175 -5594
rect 5227 -5452 5293 -5436
rect 5227 -5486 5243 -5452
rect 5277 -5486 5293 -5452
rect 5227 -5560 5293 -5486
rect 5227 -5594 5243 -5560
rect 5277 -5594 5293 -5560
rect 5227 -5610 5293 -5594
rect 5345 -5452 5411 -5436
rect 5345 -5486 5361 -5452
rect 5395 -5486 5411 -5452
rect 5345 -5560 5411 -5486
rect 5345 -5594 5361 -5560
rect 5395 -5594 5411 -5560
rect 5345 -5610 5411 -5594
rect 5463 -5452 5529 -5436
rect 5463 -5486 5479 -5452
rect 5513 -5486 5529 -5452
rect 5463 -5560 5529 -5486
rect 5463 -5594 5479 -5560
rect 5513 -5594 5529 -5560
rect 5463 -5610 5529 -5594
rect 5581 -5452 5647 -5436
rect 5581 -5486 5597 -5452
rect 5631 -5486 5647 -5452
rect 5581 -5560 5647 -5486
rect 5581 -5594 5597 -5560
rect 5631 -5594 5647 -5560
rect 5581 -5610 5647 -5594
rect 5699 -5452 5765 -5436
rect 5699 -5486 5715 -5452
rect 5749 -5486 5765 -5452
rect 5699 -5560 5765 -5486
rect 5699 -5594 5715 -5560
rect 5749 -5594 5765 -5560
rect 5699 -5610 5765 -5594
rect 5817 -5452 5883 -5436
rect 5817 -5486 5833 -5452
rect 5867 -5486 5883 -5452
rect 5817 -5560 5883 -5486
rect 5817 -5594 5833 -5560
rect 5867 -5594 5883 -5560
rect 5817 -5610 5883 -5594
rect 5935 -5452 6001 -5436
rect 5935 -5486 5951 -5452
rect 5985 -5486 6001 -5452
rect 5935 -5560 6001 -5486
rect 5935 -5594 5951 -5560
rect 5985 -5594 6001 -5560
rect 5935 -5610 6001 -5594
rect 6053 -5452 6119 -5436
rect 6053 -5486 6069 -5452
rect 6103 -5486 6119 -5452
rect 6053 -5560 6119 -5486
rect 6053 -5594 6069 -5560
rect 6103 -5594 6119 -5560
rect 6053 -5610 6119 -5594
rect 6171 -5452 6237 -5436
rect 6171 -5486 6187 -5452
rect 6221 -5486 6237 -5452
rect 6171 -5560 6237 -5486
rect 6171 -5594 6187 -5560
rect 6221 -5594 6237 -5560
rect 6171 -5610 6237 -5594
rect 6289 -5452 6355 -5436
rect 6289 -5486 6305 -5452
rect 6339 -5486 6355 -5452
rect 6289 -5560 6355 -5486
rect 6289 -5594 6305 -5560
rect 6339 -5594 6355 -5560
rect 6289 -5610 6355 -5594
rect 6407 -5452 6473 -5436
rect 6407 -5486 6423 -5452
rect 6457 -5486 6473 -5452
rect 6407 -5560 6473 -5486
rect 6407 -5594 6423 -5560
rect 6457 -5594 6473 -5560
rect 6407 -5610 6473 -5594
rect 6525 -5452 6591 -5436
rect 6525 -5486 6541 -5452
rect 6575 -5486 6591 -5452
rect 6525 -5560 6591 -5486
rect 6525 -5594 6541 -5560
rect 6575 -5594 6591 -5560
rect 6525 -5610 6591 -5594
rect 6643 -5452 6709 -5436
rect 6643 -5486 6659 -5452
rect 6693 -5486 6709 -5452
rect 6643 -5560 6709 -5486
rect 6643 -5594 6659 -5560
rect 6693 -5594 6709 -5560
rect 6643 -5610 6709 -5594
rect 6761 -5452 6827 -5436
rect 6761 -5486 6777 -5452
rect 6811 -5486 6827 -5452
rect 6761 -5560 6827 -5486
rect 6761 -5594 6777 -5560
rect 6811 -5594 6827 -5560
rect 6761 -5610 6827 -5594
rect 6879 -5452 6945 -5436
rect 6879 -5486 6895 -5452
rect 6929 -5486 6945 -5452
rect 6879 -5560 6945 -5486
rect 6879 -5594 6895 -5560
rect 6929 -5594 6945 -5560
rect 6879 -5610 6945 -5594
rect 6997 -5452 7063 -5436
rect 6997 -5486 7013 -5452
rect 7047 -5486 7063 -5452
rect 6997 -5560 7063 -5486
rect 6997 -5594 7013 -5560
rect 7047 -5594 7063 -5560
rect 6997 -5610 7063 -5594
rect 7115 -5452 7181 -5436
rect 7115 -5486 7131 -5452
rect 7165 -5486 7181 -5452
rect 7115 -5560 7181 -5486
rect 7115 -5594 7131 -5560
rect 7165 -5594 7181 -5560
rect 7115 -5610 7181 -5594
rect 11509 -7716 11599 -7562
rect 11657 -7726 11747 -7552
rect 11805 -7726 11895 -7552
rect 11953 -7726 12043 -7552
rect 12101 -7568 12191 -7552
rect 12101 -7602 12117 -7568
rect 12175 -7602 12191 -7568
rect 12101 -7676 12191 -7602
rect 12101 -7710 12117 -7676
rect 12175 -7710 12191 -7676
rect 12101 -7726 12191 -7710
rect 12249 -7568 12339 -7552
rect 12249 -7602 12265 -7568
rect 12323 -7602 12339 -7568
rect 12249 -7676 12339 -7602
rect 12249 -7710 12265 -7676
rect 12323 -7710 12339 -7676
rect 12249 -7726 12339 -7710
rect 12397 -7568 12487 -7552
rect 12397 -7602 12413 -7568
rect 12471 -7602 12487 -7568
rect 12397 -7676 12487 -7602
rect 12397 -7710 12413 -7676
rect 12471 -7710 12487 -7676
rect 12397 -7726 12487 -7710
rect 12545 -7568 12635 -7552
rect 12545 -7602 12561 -7568
rect 12619 -7602 12635 -7568
rect 12545 -7676 12635 -7602
rect 12545 -7710 12561 -7676
rect 12619 -7710 12635 -7676
rect 12545 -7726 12635 -7710
rect 12693 -7568 12783 -7552
rect 12693 -7602 12709 -7568
rect 12767 -7602 12783 -7568
rect 12693 -7676 12783 -7602
rect 12693 -7710 12709 -7676
rect 12767 -7710 12783 -7676
rect 12693 -7726 12783 -7710
rect 12841 -7568 12931 -7552
rect 12841 -7602 12857 -7568
rect 12915 -7602 12931 -7568
rect 12841 -7676 12931 -7602
rect 12841 -7710 12857 -7676
rect 12915 -7710 12931 -7676
rect 12841 -7726 12931 -7710
rect 12989 -7726 13079 -7552
rect 13137 -7726 13227 -7552
rect 13285 -7726 13375 -7552
rect 13433 -7726 13523 -7552
rect 13581 -7568 13671 -7552
rect 13581 -7602 13597 -7568
rect 13655 -7602 13671 -7568
rect 13581 -7676 13671 -7602
rect 13581 -7710 13597 -7676
rect 13655 -7710 13671 -7676
rect 13581 -7726 13671 -7710
rect 13729 -7568 13819 -7552
rect 13729 -7602 13745 -7568
rect 13803 -7602 13819 -7568
rect 13729 -7676 13819 -7602
rect 13729 -7710 13745 -7676
rect 13803 -7710 13819 -7676
rect 13729 -7726 13819 -7710
rect 13877 -7568 13967 -7552
rect 13877 -7602 13893 -7568
rect 13951 -7602 13967 -7568
rect 13877 -7676 13967 -7602
rect 13877 -7710 13893 -7676
rect 13951 -7710 13967 -7676
rect 13877 -7726 13967 -7710
rect 14025 -7568 14115 -7552
rect 14025 -7602 14041 -7568
rect 14099 -7602 14115 -7568
rect 14025 -7676 14115 -7602
rect 14025 -7710 14041 -7676
rect 14099 -7710 14115 -7676
rect 14025 -7726 14115 -7710
rect 14173 -7568 14263 -7552
rect 14173 -7602 14189 -7568
rect 14247 -7602 14263 -7568
rect 14173 -7676 14263 -7602
rect 14173 -7710 14189 -7676
rect 14247 -7710 14263 -7676
rect 14173 -7726 14263 -7710
rect 14321 -7568 14411 -7552
rect 14321 -7602 14337 -7568
rect 14395 -7602 14411 -7568
rect 14321 -7676 14411 -7602
rect 14321 -7710 14337 -7676
rect 14395 -7710 14411 -7676
rect 14321 -7726 14411 -7710
rect 14469 -7568 14559 -7552
rect 14469 -7602 14485 -7568
rect 14543 -7602 14559 -7568
rect 14469 -7676 14559 -7602
rect 14469 -7710 14485 -7676
rect 14543 -7710 14559 -7676
rect 14469 -7726 14559 -7710
rect 14617 -7568 14707 -7552
rect 14617 -7602 14633 -7568
rect 14691 -7602 14707 -7568
rect 14617 -7676 14707 -7602
rect 14617 -7710 14633 -7676
rect 14691 -7710 14707 -7676
rect 14617 -7726 14707 -7710
rect 14765 -7568 14855 -7552
rect 14765 -7602 14781 -7568
rect 14839 -7602 14855 -7568
rect 14765 -7676 14855 -7602
rect 14765 -7710 14781 -7676
rect 14839 -7710 14855 -7676
rect 14765 -7726 14855 -7710
rect 14913 -7568 15003 -7552
rect 14913 -7602 14929 -7568
rect 14987 -7602 15003 -7568
rect 14913 -7676 15003 -7602
rect 14913 -7710 14929 -7676
rect 14987 -7710 15003 -7676
rect 14913 -7726 15003 -7710
rect 15061 -7568 15151 -7552
rect 15061 -7602 15077 -7568
rect 15135 -7602 15151 -7568
rect 15061 -7676 15151 -7602
rect 15061 -7710 15077 -7676
rect 15135 -7710 15151 -7676
rect 15061 -7726 15151 -7710
rect 15209 -7568 15299 -7552
rect 15209 -7602 15225 -7568
rect 15283 -7602 15299 -7568
rect 15209 -7676 15299 -7602
rect 15209 -7710 15225 -7676
rect 15283 -7710 15299 -7676
rect 15209 -7726 15299 -7710
rect 15357 -7568 15447 -7552
rect 15357 -7602 15373 -7568
rect 15431 -7602 15447 -7568
rect 15357 -7676 15447 -7602
rect 15357 -7710 15373 -7676
rect 15431 -7710 15447 -7676
rect 15357 -7726 15447 -7710
rect 15505 -7568 15595 -7552
rect 15505 -7602 15521 -7568
rect 15579 -7602 15595 -7568
rect 15505 -7676 15595 -7602
rect 15505 -7710 15521 -7676
rect 15579 -7710 15595 -7676
rect 15505 -7726 15595 -7710
rect 15653 -7568 15743 -7552
rect 15653 -7602 15669 -7568
rect 15727 -7602 15743 -7568
rect 15653 -7676 15743 -7602
rect 15653 -7710 15669 -7676
rect 15727 -7710 15743 -7676
rect 15653 -7726 15743 -7710
rect 15801 -7568 15891 -7552
rect 15801 -7602 15817 -7568
rect 15875 -7602 15891 -7568
rect 15801 -7676 15891 -7602
rect 15801 -7710 15817 -7676
rect 15875 -7710 15891 -7676
rect 15801 -7726 15891 -7710
rect 15949 -7568 16039 -7552
rect 15949 -7602 15965 -7568
rect 16023 -7602 16039 -7568
rect 15949 -7676 16039 -7602
rect 15949 -7710 15965 -7676
rect 16023 -7710 16039 -7676
rect 15949 -7726 16039 -7710
rect 16097 -7568 16187 -7552
rect 16097 -7602 16113 -7568
rect 16171 -7602 16187 -7568
rect 16097 -7676 16187 -7602
rect 16097 -7710 16113 -7676
rect 16171 -7710 16187 -7676
rect 16097 -7726 16187 -7710
rect 16245 -7568 16335 -7552
rect 16245 -7602 16261 -7568
rect 16319 -7602 16335 -7568
rect 16245 -7676 16335 -7602
rect 16245 -7710 16261 -7676
rect 16319 -7710 16335 -7676
rect 16245 -7726 16335 -7710
rect 16393 -7568 16483 -7552
rect 16393 -7602 16409 -7568
rect 16467 -7602 16483 -7568
rect 16393 -7676 16483 -7602
rect 16393 -7710 16409 -7676
rect 16467 -7710 16483 -7676
rect 16393 -7726 16483 -7710
rect 16541 -7568 16631 -7552
rect 16541 -7602 16557 -7568
rect 16615 -7602 16631 -7568
rect 16541 -7676 16631 -7602
rect 16541 -7710 16557 -7676
rect 16615 -7710 16631 -7676
rect 16541 -7726 16631 -7710
rect 16689 -7568 16779 -7552
rect 16689 -7602 16705 -7568
rect 16763 -7602 16779 -7568
rect 16689 -7676 16779 -7602
rect 16689 -7710 16705 -7676
rect 16763 -7710 16779 -7676
rect 16689 -7726 16779 -7710
rect 16837 -7568 16927 -7552
rect 16837 -7602 16853 -7568
rect 16911 -7602 16927 -7568
rect 16837 -7676 16927 -7602
rect 16837 -7710 16853 -7676
rect 16911 -7710 16927 -7676
rect 16837 -7726 16927 -7710
rect 16985 -7568 17075 -7552
rect 16985 -7602 17001 -7568
rect 17059 -7602 17075 -7568
rect 16985 -7676 17075 -7602
rect 16985 -7710 17001 -7676
rect 17059 -7710 17075 -7676
rect 16985 -7726 17075 -7710
rect 17133 -7568 17223 -7552
rect 17133 -7602 17149 -7568
rect 17207 -7602 17223 -7568
rect 17133 -7676 17223 -7602
rect 17133 -7710 17149 -7676
rect 17207 -7710 17223 -7676
rect 17133 -7726 17223 -7710
rect 17281 -7568 17371 -7552
rect 17281 -7602 17297 -7568
rect 17355 -7602 17371 -7568
rect 17281 -7676 17371 -7602
rect 17281 -7710 17297 -7676
rect 17355 -7710 17371 -7676
rect 17281 -7726 17371 -7710
rect 17429 -7568 17519 -7552
rect 17429 -7602 17445 -7568
rect 17503 -7602 17519 -7568
rect 17429 -7676 17519 -7602
rect 17429 -7710 17445 -7676
rect 17503 -7710 17519 -7676
rect 17429 -7726 17519 -7710
rect 17577 -7568 17667 -7552
rect 17577 -7602 17593 -7568
rect 17651 -7602 17667 -7568
rect 17577 -7676 17667 -7602
rect 17577 -7710 17593 -7676
rect 17651 -7710 17667 -7676
rect 17577 -7726 17667 -7710
rect 17725 -7568 17815 -7552
rect 17725 -7602 17741 -7568
rect 17799 -7602 17815 -7568
rect 17725 -7676 17815 -7602
rect 17725 -7710 17741 -7676
rect 17799 -7710 17815 -7676
rect 17725 -7726 17815 -7710
rect 17873 -7568 17963 -7552
rect 17873 -7602 17889 -7568
rect 17947 -7602 17963 -7568
rect 17873 -7676 17963 -7602
rect 17873 -7710 17889 -7676
rect 17947 -7710 17963 -7676
rect 17873 -7726 17963 -7710
rect 18021 -7568 18111 -7552
rect 18021 -7602 18037 -7568
rect 18095 -7602 18111 -7568
rect 18021 -7676 18111 -7602
rect 18021 -7710 18037 -7676
rect 18095 -7710 18111 -7676
rect 18021 -7726 18111 -7710
rect 18169 -7726 18259 -7552
rect 18317 -7726 18407 -7552
rect 18465 -7726 18555 -7552
rect 18613 -7726 18703 -7552
rect 18761 -7568 18851 -7552
rect 18761 -7602 18777 -7568
rect 18835 -7602 18851 -7568
rect 18761 -7676 18851 -7602
rect 18761 -7710 18777 -7676
rect 18835 -7710 18851 -7676
rect 18761 -7726 18851 -7710
rect 18909 -7568 18999 -7552
rect 18909 -7602 18925 -7568
rect 18983 -7602 18999 -7568
rect 18909 -7676 18999 -7602
rect 18909 -7710 18925 -7676
rect 18983 -7710 18999 -7676
rect 18909 -7726 18999 -7710
rect 19057 -7568 19147 -7552
rect 19057 -7602 19073 -7568
rect 19131 -7602 19147 -7568
rect 19057 -7676 19147 -7602
rect 19057 -7710 19073 -7676
rect 19131 -7710 19147 -7676
rect 19057 -7726 19147 -7710
rect 19205 -7568 19295 -7552
rect 19205 -7602 19221 -7568
rect 19279 -7602 19295 -7568
rect 19205 -7676 19295 -7602
rect 19205 -7710 19221 -7676
rect 19279 -7710 19295 -7676
rect 19205 -7726 19295 -7710
rect 19353 -7568 19443 -7552
rect 19353 -7602 19369 -7568
rect 19427 -7602 19443 -7568
rect 19353 -7676 19443 -7602
rect 19353 -7710 19369 -7676
rect 19427 -7710 19443 -7676
rect 19353 -7726 19443 -7710
rect 19501 -7568 19591 -7552
rect 19501 -7602 19517 -7568
rect 19575 -7602 19591 -7568
rect 19501 -7676 19591 -7602
rect 19501 -7710 19517 -7676
rect 19575 -7710 19591 -7676
rect 19501 -7726 19591 -7710
rect 19649 -7568 19739 -7552
rect 19649 -7602 19665 -7568
rect 19723 -7602 19739 -7568
rect 19649 -7676 19739 -7602
rect 19649 -7710 19665 -7676
rect 19723 -7710 19739 -7676
rect 19649 -7726 19739 -7710
rect 19797 -7568 19887 -7552
rect 19797 -7602 19813 -7568
rect 19871 -7602 19887 -7568
rect 19797 -7676 19887 -7602
rect 19797 -7710 19813 -7676
rect 19871 -7710 19887 -7676
rect 19797 -7726 19887 -7710
rect 19945 -7568 20035 -7552
rect 19945 -7602 19961 -7568
rect 20019 -7602 20035 -7568
rect 19945 -7676 20035 -7602
rect 19945 -7710 19961 -7676
rect 20019 -7710 20035 -7676
rect 19945 -7726 20035 -7710
rect 20093 -7568 20183 -7552
rect 20093 -7602 20109 -7568
rect 20167 -7602 20183 -7568
rect 20093 -7676 20183 -7602
rect 20093 -7710 20109 -7676
rect 20167 -7710 20183 -7676
rect 20093 -7726 20183 -7710
rect 20241 -7568 20331 -7552
rect 20241 -7602 20257 -7568
rect 20315 -7602 20331 -7568
rect 20241 -7676 20331 -7602
rect 20241 -7710 20257 -7676
rect 20315 -7710 20331 -7676
rect 20241 -7726 20331 -7710
rect 20389 -7568 20479 -7552
rect 20389 -7602 20405 -7568
rect 20463 -7602 20479 -7568
rect 20389 -7676 20479 -7602
rect 20389 -7710 20405 -7676
rect 20463 -7710 20479 -7676
rect 20389 -7726 20479 -7710
rect 20537 -7568 20627 -7552
rect 20537 -7602 20553 -7568
rect 20611 -7602 20627 -7568
rect 20537 -7676 20627 -7602
rect 20537 -7710 20553 -7676
rect 20611 -7710 20627 -7676
rect 20537 -7726 20627 -7710
rect 20685 -7568 20775 -7552
rect 20685 -7602 20701 -7568
rect 20759 -7602 20775 -7568
rect 20685 -7676 20775 -7602
rect 20685 -7710 20701 -7676
rect 20759 -7710 20775 -7676
rect 20685 -7726 20775 -7710
rect 20833 -7568 20923 -7552
rect 20833 -7602 20849 -7568
rect 20907 -7602 20923 -7568
rect 20833 -7676 20923 -7602
rect 20833 -7710 20849 -7676
rect 20907 -7710 20923 -7676
rect 20833 -7726 20923 -7710
rect 20981 -7568 21071 -7552
rect 20981 -7602 20997 -7568
rect 21055 -7602 21071 -7568
rect 20981 -7676 21071 -7602
rect 20981 -7710 20997 -7676
rect 21055 -7710 21071 -7676
rect 20981 -7726 21071 -7710
rect 21129 -7568 21219 -7552
rect 21129 -7602 21145 -7568
rect 21203 -7602 21219 -7568
rect 21129 -7676 21219 -7602
rect 21129 -7710 21145 -7676
rect 21203 -7710 21219 -7676
rect 21129 -7726 21219 -7710
rect 21277 -7568 21367 -7552
rect 21277 -7602 21293 -7568
rect 21351 -7602 21367 -7568
rect 21277 -7676 21367 -7602
rect 21277 -7710 21293 -7676
rect 21351 -7710 21367 -7676
rect 21277 -7726 21367 -7710
rect 21425 -7568 21515 -7552
rect 21425 -7602 21441 -7568
rect 21499 -7602 21515 -7568
rect 21425 -7676 21515 -7602
rect 21425 -7710 21441 -7676
rect 21499 -7710 21515 -7676
rect 21425 -7726 21515 -7710
rect 21573 -7568 21663 -7552
rect 21573 -7602 21589 -7568
rect 21647 -7602 21663 -7568
rect 21573 -7676 21663 -7602
rect 21573 -7710 21589 -7676
rect 21647 -7710 21663 -7676
rect 21573 -7726 21663 -7710
rect 21721 -7568 21811 -7552
rect 21721 -7602 21737 -7568
rect 21795 -7602 21811 -7568
rect 21721 -7676 21811 -7602
rect 21721 -7710 21737 -7676
rect 21795 -7710 21811 -7676
rect 21721 -7726 21811 -7710
rect 21869 -7568 21959 -7552
rect 21869 -7602 21885 -7568
rect 21943 -7602 21959 -7568
rect 21869 -7676 21959 -7602
rect 21869 -7710 21885 -7676
rect 21943 -7710 21959 -7676
rect 21869 -7726 21959 -7710
rect 22017 -7568 22107 -7552
rect 22017 -7602 22033 -7568
rect 22091 -7602 22107 -7568
rect 22017 -7676 22107 -7602
rect 22017 -7710 22033 -7676
rect 22091 -7710 22107 -7676
rect 22017 -7726 22107 -7710
rect 22165 -7568 22255 -7552
rect 22165 -7602 22181 -7568
rect 22239 -7602 22255 -7568
rect 22165 -7676 22255 -7602
rect 22165 -7710 22181 -7676
rect 22239 -7710 22255 -7676
rect 22165 -7726 22255 -7710
rect 22313 -7568 22403 -7552
rect 22313 -7602 22329 -7568
rect 22387 -7602 22403 -7568
rect 22313 -7676 22403 -7602
rect 22313 -7710 22329 -7676
rect 22387 -7710 22403 -7676
rect 22313 -7726 22403 -7710
rect 22461 -7568 22551 -7552
rect 22461 -7602 22477 -7568
rect 22535 -7602 22551 -7568
rect 22461 -7676 22551 -7602
rect 22461 -7710 22477 -7676
rect 22535 -7710 22551 -7676
rect 22461 -7726 22551 -7710
rect 3059 -7767 3125 -7751
rect 3059 -7801 3075 -7767
rect 3109 -7801 3125 -7767
rect 3059 -7875 3125 -7801
rect 3059 -7909 3075 -7875
rect 3109 -7909 3125 -7875
rect 3059 -7925 3125 -7909
rect 3177 -7767 3243 -7751
rect 3177 -7801 3193 -7767
rect 3227 -7801 3243 -7767
rect 3177 -7875 3243 -7801
rect 3177 -7909 3193 -7875
rect 3227 -7909 3243 -7875
rect 3177 -7925 3243 -7909
rect 3295 -7767 3361 -7751
rect 3295 -7801 3311 -7767
rect 3345 -7801 3361 -7767
rect 3295 -7875 3361 -7801
rect 3295 -7909 3311 -7875
rect 3345 -7909 3361 -7875
rect 3295 -7925 3361 -7909
rect 3413 -7767 3479 -7751
rect 3413 -7801 3429 -7767
rect 3463 -7801 3479 -7767
rect 3413 -7875 3479 -7801
rect 3413 -7909 3429 -7875
rect 3463 -7909 3479 -7875
rect 3413 -7925 3479 -7909
rect 3531 -7767 3597 -7751
rect 3531 -7801 3547 -7767
rect 3581 -7801 3597 -7767
rect 3531 -7875 3597 -7801
rect 3531 -7909 3547 -7875
rect 3581 -7909 3597 -7875
rect 3531 -7925 3597 -7909
rect 3649 -7767 3715 -7751
rect 3649 -7801 3665 -7767
rect 3699 -7801 3715 -7767
rect 3649 -7875 3715 -7801
rect 3649 -7909 3665 -7875
rect 3699 -7909 3715 -7875
rect 3649 -7925 3715 -7909
rect 3767 -7767 3833 -7751
rect 3767 -7801 3783 -7767
rect 3817 -7801 3833 -7767
rect 3767 -7875 3833 -7801
rect 3767 -7909 3783 -7875
rect 3817 -7909 3833 -7875
rect 3767 -7925 3833 -7909
rect 3885 -7767 3951 -7751
rect 3885 -7801 3901 -7767
rect 3935 -7801 3951 -7767
rect 3885 -7875 3951 -7801
rect 3885 -7909 3901 -7875
rect 3935 -7909 3951 -7875
rect 3885 -7925 3951 -7909
rect 4003 -7767 4069 -7751
rect 4003 -7801 4019 -7767
rect 4053 -7801 4069 -7767
rect 4003 -7875 4069 -7801
rect 4003 -7909 4019 -7875
rect 4053 -7909 4069 -7875
rect 4003 -7925 4069 -7909
rect 4121 -7767 4187 -7751
rect 4121 -7801 4137 -7767
rect 4171 -7801 4187 -7767
rect 4121 -7875 4187 -7801
rect 4121 -7909 4137 -7875
rect 4171 -7909 4187 -7875
rect 4121 -7925 4187 -7909
rect 4239 -7767 4305 -7751
rect 4239 -7801 4255 -7767
rect 4289 -7801 4305 -7767
rect 4239 -7875 4305 -7801
rect 4239 -7909 4255 -7875
rect 4289 -7909 4305 -7875
rect 4239 -7925 4305 -7909
rect 4357 -7767 4423 -7751
rect 4357 -7801 4373 -7767
rect 4407 -7801 4423 -7767
rect 4357 -7875 4423 -7801
rect 4357 -7909 4373 -7875
rect 4407 -7909 4423 -7875
rect 4357 -7925 4423 -7909
rect 4475 -7767 4541 -7751
rect 4475 -7801 4491 -7767
rect 4525 -7801 4541 -7767
rect 4475 -7875 4541 -7801
rect 4475 -7909 4491 -7875
rect 4525 -7909 4541 -7875
rect 4475 -7925 4541 -7909
rect 4593 -7767 4659 -7751
rect 4593 -7801 4609 -7767
rect 4643 -7801 4659 -7767
rect 4593 -7875 4659 -7801
rect 4593 -7909 4609 -7875
rect 4643 -7909 4659 -7875
rect 4593 -7925 4659 -7909
rect 4711 -7767 4777 -7751
rect 4711 -7801 4727 -7767
rect 4761 -7801 4777 -7767
rect 4711 -7875 4777 -7801
rect 4711 -7909 4727 -7875
rect 4761 -7909 4777 -7875
rect 4711 -7925 4777 -7909
rect 5057 -7767 5123 -7751
rect 5057 -7801 5073 -7767
rect 5107 -7801 5123 -7767
rect 5057 -7875 5123 -7801
rect 5057 -7909 5073 -7875
rect 5107 -7909 5123 -7875
rect 5057 -7925 5123 -7909
rect 5175 -7767 5241 -7751
rect 5175 -7801 5191 -7767
rect 5225 -7801 5241 -7767
rect 5175 -7875 5241 -7801
rect 5175 -7909 5191 -7875
rect 5225 -7909 5241 -7875
rect 5175 -7925 5241 -7909
rect 5293 -7767 5359 -7751
rect 5293 -7801 5309 -7767
rect 5343 -7801 5359 -7767
rect 5293 -7875 5359 -7801
rect 5293 -7909 5309 -7875
rect 5343 -7909 5359 -7875
rect 5293 -7925 5359 -7909
rect 5411 -7767 5477 -7751
rect 5411 -7801 5427 -7767
rect 5461 -7801 5477 -7767
rect 5411 -7875 5477 -7801
rect 5411 -7909 5427 -7875
rect 5461 -7909 5477 -7875
rect 5411 -7925 5477 -7909
rect 5529 -7767 5595 -7751
rect 5529 -7801 5545 -7767
rect 5579 -7801 5595 -7767
rect 5529 -7875 5595 -7801
rect 5529 -7909 5545 -7875
rect 5579 -7909 5595 -7875
rect 5529 -7925 5595 -7909
rect 5647 -7767 5713 -7751
rect 5647 -7801 5663 -7767
rect 5697 -7801 5713 -7767
rect 5647 -7875 5713 -7801
rect 5647 -7909 5663 -7875
rect 5697 -7909 5713 -7875
rect 5647 -7925 5713 -7909
rect 5765 -7767 5831 -7751
rect 5765 -7801 5781 -7767
rect 5815 -7801 5831 -7767
rect 5765 -7875 5831 -7801
rect 5765 -7909 5781 -7875
rect 5815 -7909 5831 -7875
rect 5765 -7925 5831 -7909
rect 5883 -7767 5949 -7751
rect 5883 -7801 5899 -7767
rect 5933 -7801 5949 -7767
rect 5883 -7875 5949 -7801
rect 5883 -7909 5899 -7875
rect 5933 -7909 5949 -7875
rect 5883 -7925 5949 -7909
rect 6001 -7767 6067 -7751
rect 6001 -7801 6017 -7767
rect 6051 -7801 6067 -7767
rect 6001 -7875 6067 -7801
rect 6001 -7909 6017 -7875
rect 6051 -7909 6067 -7875
rect 6001 -7925 6067 -7909
rect 6119 -7767 6185 -7751
rect 6119 -7801 6135 -7767
rect 6169 -7801 6185 -7767
rect 6119 -7875 6185 -7801
rect 6119 -7909 6135 -7875
rect 6169 -7909 6185 -7875
rect 6119 -7925 6185 -7909
rect 6237 -7767 6303 -7751
rect 6237 -7801 6253 -7767
rect 6287 -7801 6303 -7767
rect 6237 -7875 6303 -7801
rect 6237 -7909 6253 -7875
rect 6287 -7909 6303 -7875
rect 6237 -7925 6303 -7909
rect 6355 -7767 6421 -7751
rect 6355 -7801 6371 -7767
rect 6405 -7801 6421 -7767
rect 6355 -7875 6421 -7801
rect 6355 -7909 6371 -7875
rect 6405 -7909 6421 -7875
rect 6355 -7925 6421 -7909
rect 6473 -7767 6539 -7751
rect 6473 -7801 6489 -7767
rect 6523 -7801 6539 -7767
rect 6473 -7875 6539 -7801
rect 6473 -7909 6489 -7875
rect 6523 -7909 6539 -7875
rect 6473 -7925 6539 -7909
rect 6591 -7767 6657 -7751
rect 6591 -7801 6607 -7767
rect 6641 -7801 6657 -7767
rect 6591 -7875 6657 -7801
rect 6591 -7909 6607 -7875
rect 6641 -7909 6657 -7875
rect 6591 -7925 6657 -7909
rect 6709 -7767 6775 -7751
rect 6709 -7801 6725 -7767
rect 6759 -7801 6775 -7767
rect 6709 -7875 6775 -7801
rect 6709 -7909 6725 -7875
rect 6759 -7909 6775 -7875
rect 6709 -7925 6775 -7909
<< polycont >>
rect 7555 2006 7589 2040
rect 7673 2006 7707 2040
rect 7791 2006 7825 2040
rect 7909 2006 7943 2040
rect 8027 2006 8061 2040
rect 8145 2006 8179 2040
rect 8263 2006 8297 2040
rect 8609 2006 8643 2040
rect 8727 2006 8761 2040
rect 8845 2006 8879 2040
rect 8963 2006 8997 2040
rect 9081 2006 9115 2040
rect 9199 2006 9233 2040
rect 9317 2006 9351 2040
rect 9435 2006 9469 2040
rect 9553 2006 9587 2040
rect 9671 2006 9705 2040
rect 9789 2006 9823 2040
rect 9907 2006 9941 2040
rect 10025 2006 10059 2040
rect 10143 2006 10177 2040
rect 10261 2006 10295 2040
rect 12677 2005 12711 2039
rect 12795 2005 12829 2039
rect 12913 2005 12947 2039
rect 13031 2005 13065 2039
rect 13149 2005 13183 2039
rect 13267 2005 13301 2039
rect 13385 2005 13419 2039
rect 13503 2005 13537 2039
rect 13621 2005 13655 2039
rect 13739 2005 13773 2039
rect 13857 2005 13891 2039
rect 13975 2005 14009 2039
rect 14093 2005 14127 2039
rect 14211 2005 14245 2039
rect 14329 2005 14363 2039
rect 14447 2005 14481 2039
rect 14565 2005 14599 2039
rect 14683 2005 14717 2039
rect 14801 2005 14835 2039
rect 14919 2005 14953 2039
rect 15037 2005 15071 2039
rect 15155 2005 15189 2039
rect 15273 2005 15307 2039
rect 15391 2005 15425 2039
rect 15509 2005 15543 2039
rect 15627 2005 15661 2039
rect 15745 2005 15779 2039
rect 15863 2005 15897 2039
rect 15981 2005 16015 2039
rect 16099 2005 16133 2039
rect 16217 2005 16251 2039
rect 16335 2005 16369 2039
rect 16453 2005 16487 2039
rect 16571 2005 16605 2039
rect 16689 2005 16723 2039
rect 16807 2005 16841 2039
rect 16925 2005 16959 2039
rect 17043 2005 17077 2039
rect 17161 2005 17195 2039
rect 17279 2005 17313 2039
rect 17397 2005 17431 2039
rect 17515 2005 17549 2039
rect 17633 2005 17667 2039
rect 17751 2005 17785 2039
rect 17869 2005 17903 2039
rect 17987 2005 18021 2039
rect 18105 2005 18139 2039
rect 18223 2005 18257 2039
rect 18341 2005 18375 2039
rect 18459 2005 18493 2039
rect 18577 2005 18611 2039
rect 18695 2005 18729 2039
rect 18813 2005 18847 2039
rect 18931 2005 18965 2039
rect 19049 2005 19083 2039
rect 19167 2005 19201 2039
rect 19285 2005 19319 2039
rect 19403 2005 19437 2039
rect 19521 2005 19555 2039
rect 19639 2005 19673 2039
rect 19757 2005 19791 2039
rect 19875 2005 19909 2039
rect 19993 2005 20027 2039
rect 20111 2005 20145 2039
rect 20229 2005 20263 2039
rect 20347 2005 20381 2039
rect 20465 2005 20499 2039
rect 20583 2005 20617 2039
rect 20701 2005 20735 2039
rect 20819 2005 20853 2039
rect 20937 2005 20971 2039
rect 21055 2005 21089 2039
rect 21173 2005 21207 2039
rect 21291 2005 21325 2039
rect 12677 1897 12711 1931
rect 12795 1897 12829 1931
rect 12913 1897 12947 1931
rect 13031 1897 13065 1931
rect 13149 1897 13183 1931
rect 13267 1897 13301 1931
rect 13385 1897 13419 1931
rect 13503 1897 13537 1931
rect 13621 1897 13655 1931
rect 13739 1897 13773 1931
rect 13857 1897 13891 1931
rect 13975 1897 14009 1931
rect 14093 1897 14127 1931
rect 14211 1897 14245 1931
rect 14329 1897 14363 1931
rect 14447 1897 14481 1931
rect 14565 1897 14599 1931
rect 14683 1897 14717 1931
rect 14801 1897 14835 1931
rect 14919 1897 14953 1931
rect 15037 1897 15071 1931
rect 15155 1897 15189 1931
rect 15273 1897 15307 1931
rect 15391 1897 15425 1931
rect 15509 1897 15543 1931
rect 15627 1897 15661 1931
rect 15745 1897 15779 1931
rect 15863 1897 15897 1931
rect 15981 1897 16015 1931
rect 16099 1897 16133 1931
rect 16217 1897 16251 1931
rect 16335 1897 16369 1931
rect 16453 1897 16487 1931
rect 16571 1897 16605 1931
rect 16689 1897 16723 1931
rect 16807 1897 16841 1931
rect 16925 1897 16959 1931
rect 17043 1897 17077 1931
rect 17161 1897 17195 1931
rect 17279 1897 17313 1931
rect 17397 1897 17431 1931
rect 17515 1897 17549 1931
rect 17633 1897 17667 1931
rect 17751 1897 17785 1931
rect 17869 1897 17903 1931
rect 17987 1897 18021 1931
rect 18105 1897 18139 1931
rect 18223 1897 18257 1931
rect 18341 1897 18375 1931
rect 18459 1897 18493 1931
rect 18577 1897 18611 1931
rect 18695 1897 18729 1931
rect 18813 1897 18847 1931
rect 18931 1897 18965 1931
rect 19049 1897 19083 1931
rect 19167 1897 19201 1931
rect 19285 1897 19319 1931
rect 19403 1897 19437 1931
rect 19521 1897 19555 1931
rect 19639 1897 19673 1931
rect 19757 1897 19791 1931
rect 19875 1897 19909 1931
rect 19993 1897 20027 1931
rect 20111 1897 20145 1931
rect 20229 1897 20263 1931
rect 20347 1897 20381 1931
rect 20465 1897 20499 1931
rect 20583 1897 20617 1931
rect 20701 1897 20735 1931
rect 20819 1897 20853 1931
rect 20937 1897 20971 1931
rect 21055 1897 21089 1931
rect 21173 1897 21207 1931
rect 21291 1897 21325 1931
rect 2293 -182 2327 -148
rect 2293 -290 2327 -256
rect 2411 -182 2445 -148
rect 2411 -290 2445 -256
rect 2529 -182 2563 -148
rect 2529 -290 2563 -256
rect 2647 -182 2681 -148
rect 2647 -290 2681 -256
rect 1349 -3718 1383 -3684
rect 1349 -3826 1383 -3792
rect 1467 -3718 1501 -3684
rect 1467 -3826 1501 -3792
rect 1585 -3718 1619 -3684
rect 1585 -3826 1619 -3792
rect 1703 -3718 1737 -3684
rect 1703 -3826 1737 -3792
rect 1821 -3718 1855 -3684
rect 1821 -3826 1855 -3792
rect 1939 -3718 1973 -3684
rect 1939 -3826 1973 -3792
rect 2057 -3718 2091 -3684
rect 2057 -3826 2091 -3792
rect 2175 -3718 2209 -3684
rect 2175 -3826 2209 -3792
rect 2293 -3718 2327 -3684
rect 2293 -3826 2327 -3792
rect 2411 -3718 2445 -3684
rect 2411 -3826 2445 -3792
rect 2529 -3718 2563 -3684
rect 2529 -3826 2563 -3792
rect 2647 -3718 2681 -3684
rect 2647 -3826 2681 -3792
rect 2765 -3718 2799 -3684
rect 2765 -3826 2799 -3792
rect 2883 -3718 2917 -3684
rect 2883 -3826 2917 -3792
rect 3001 -3718 3035 -3684
rect 3001 -3826 3035 -3792
rect 3119 -3718 3153 -3684
rect 3119 -3826 3153 -3792
rect 3237 -3718 3271 -3684
rect 3237 -3826 3271 -3792
rect 3355 -3718 3389 -3684
rect 3355 -3826 3389 -3792
rect 3473 -3718 3507 -3684
rect 3473 -3826 3507 -3792
rect 3591 -3718 3625 -3684
rect 3591 -3826 3625 -3792
rect 3709 -3718 3743 -3684
rect 3709 -3826 3743 -3792
rect 3827 -3718 3861 -3684
rect 3827 -3826 3861 -3792
rect 3945 -3718 3979 -3684
rect 3945 -3826 3979 -3792
rect 4063 -3718 4097 -3684
rect 4063 -3826 4097 -3792
rect 4181 -3718 4215 -3684
rect 4181 -3826 4215 -3792
rect 4299 -3718 4333 -3684
rect 4299 -3826 4333 -3792
rect 4417 -3718 4451 -3684
rect 4417 -3826 4451 -3792
rect 4535 -3718 4569 -3684
rect 4535 -3826 4569 -3792
rect 4653 -3718 4687 -3684
rect 4653 -3826 4687 -3792
rect 4771 -3718 4805 -3684
rect 4771 -3826 4805 -3792
rect 4889 -3718 4923 -3684
rect 4889 -3826 4923 -3792
rect 5007 -3718 5041 -3684
rect 5007 -3826 5041 -3792
rect 5125 -3718 5159 -3684
rect 5125 -3826 5159 -3792
rect 5243 -3718 5277 -3684
rect 5243 -3826 5277 -3792
rect 5361 -3718 5395 -3684
rect 5361 -3826 5395 -3792
rect 5479 -3718 5513 -3684
rect 5479 -3826 5513 -3792
rect 5597 -3718 5631 -3684
rect 5597 -3826 5631 -3792
rect 5715 -3718 5749 -3684
rect 5715 -3826 5749 -3792
rect 5833 -3718 5867 -3684
rect 5833 -3826 5867 -3792
rect 5951 -3718 5985 -3684
rect 5951 -3826 5985 -3792
rect 6069 -3718 6103 -3684
rect 6069 -3826 6103 -3792
rect 6187 -3718 6221 -3684
rect 6187 -3826 6221 -3792
rect 6305 -3718 6339 -3684
rect 6305 -3826 6339 -3792
rect 6423 -3718 6457 -3684
rect 6423 -3826 6457 -3792
rect 6541 -3718 6575 -3684
rect 6541 -3826 6575 -3792
rect 6659 -3718 6693 -3684
rect 6659 -3826 6693 -3792
rect 6777 -3718 6811 -3684
rect 6777 -3826 6811 -3792
rect 6895 -3718 6929 -3684
rect 6895 -3826 6929 -3792
rect 7013 -3718 7047 -3684
rect 7013 -3826 7047 -3792
rect 7131 -3718 7165 -3684
rect 7131 -3826 7165 -3792
rect 1349 -5486 1383 -5452
rect 1349 -5594 1383 -5560
rect 1467 -5486 1501 -5452
rect 1467 -5594 1501 -5560
rect 1585 -5486 1619 -5452
rect 1585 -5594 1619 -5560
rect 1703 -5486 1737 -5452
rect 1703 -5594 1737 -5560
rect 1821 -5486 1855 -5452
rect 1821 -5594 1855 -5560
rect 1939 -5486 1973 -5452
rect 1939 -5594 1973 -5560
rect 2057 -5486 2091 -5452
rect 2057 -5594 2091 -5560
rect 2175 -5486 2209 -5452
rect 2175 -5594 2209 -5560
rect 2293 -5486 2327 -5452
rect 2293 -5594 2327 -5560
rect 2411 -5486 2445 -5452
rect 2411 -5594 2445 -5560
rect 2529 -5486 2563 -5452
rect 2529 -5594 2563 -5560
rect 2647 -5486 2681 -5452
rect 2647 -5594 2681 -5560
rect 2765 -5486 2799 -5452
rect 2765 -5594 2799 -5560
rect 2883 -5486 2917 -5452
rect 2883 -5594 2917 -5560
rect 3001 -5486 3035 -5452
rect 3001 -5594 3035 -5560
rect 3119 -5486 3153 -5452
rect 3119 -5594 3153 -5560
rect 3237 -5486 3271 -5452
rect 3237 -5594 3271 -5560
rect 3355 -5486 3389 -5452
rect 3355 -5594 3389 -5560
rect 3473 -5486 3507 -5452
rect 3473 -5594 3507 -5560
rect 3591 -5486 3625 -5452
rect 3591 -5594 3625 -5560
rect 3709 -5486 3743 -5452
rect 3709 -5594 3743 -5560
rect 3827 -5486 3861 -5452
rect 3827 -5594 3861 -5560
rect 3945 -5486 3979 -5452
rect 3945 -5594 3979 -5560
rect 4063 -5486 4097 -5452
rect 4063 -5594 4097 -5560
rect 4181 -5486 4215 -5452
rect 4181 -5594 4215 -5560
rect 4299 -5486 4333 -5452
rect 4299 -5594 4333 -5560
rect 4417 -5486 4451 -5452
rect 4417 -5594 4451 -5560
rect 4535 -5486 4569 -5452
rect 4535 -5594 4569 -5560
rect 4653 -5486 4687 -5452
rect 4653 -5594 4687 -5560
rect 4771 -5486 4805 -5452
rect 4771 -5594 4805 -5560
rect 4889 -5486 4923 -5452
rect 4889 -5594 4923 -5560
rect 5007 -5486 5041 -5452
rect 5007 -5594 5041 -5560
rect 5125 -5486 5159 -5452
rect 5125 -5594 5159 -5560
rect 5243 -5486 5277 -5452
rect 5243 -5594 5277 -5560
rect 5361 -5486 5395 -5452
rect 5361 -5594 5395 -5560
rect 5479 -5486 5513 -5452
rect 5479 -5594 5513 -5560
rect 5597 -5486 5631 -5452
rect 5597 -5594 5631 -5560
rect 5715 -5486 5749 -5452
rect 5715 -5594 5749 -5560
rect 5833 -5486 5867 -5452
rect 5833 -5594 5867 -5560
rect 5951 -5486 5985 -5452
rect 5951 -5594 5985 -5560
rect 6069 -5486 6103 -5452
rect 6069 -5594 6103 -5560
rect 6187 -5486 6221 -5452
rect 6187 -5594 6221 -5560
rect 6305 -5486 6339 -5452
rect 6305 -5594 6339 -5560
rect 6423 -5486 6457 -5452
rect 6423 -5594 6457 -5560
rect 6541 -5486 6575 -5452
rect 6541 -5594 6575 -5560
rect 6659 -5486 6693 -5452
rect 6659 -5594 6693 -5560
rect 6777 -5486 6811 -5452
rect 6777 -5594 6811 -5560
rect 6895 -5486 6929 -5452
rect 6895 -5594 6929 -5560
rect 7013 -5486 7047 -5452
rect 7013 -5594 7047 -5560
rect 7131 -5486 7165 -5452
rect 7131 -5594 7165 -5560
rect 12117 -7602 12175 -7568
rect 12117 -7710 12175 -7676
rect 12265 -7602 12323 -7568
rect 12265 -7710 12323 -7676
rect 12413 -7602 12471 -7568
rect 12413 -7710 12471 -7676
rect 12561 -7602 12619 -7568
rect 12561 -7710 12619 -7676
rect 12709 -7602 12767 -7568
rect 12709 -7710 12767 -7676
rect 12857 -7602 12915 -7568
rect 12857 -7710 12915 -7676
rect 14485 -7602 14543 -7568
rect 14485 -7710 14543 -7676
rect 14633 -7602 14691 -7568
rect 14633 -7710 14691 -7676
rect 14781 -7602 14839 -7568
rect 14781 -7710 14839 -7676
rect 14929 -7602 14987 -7568
rect 14929 -7710 14987 -7676
rect 15077 -7602 15135 -7568
rect 15077 -7710 15135 -7676
rect 15225 -7602 15283 -7568
rect 15225 -7710 15283 -7676
rect 15373 -7602 15431 -7568
rect 15373 -7710 15431 -7676
rect 15521 -7602 15579 -7568
rect 15521 -7710 15579 -7676
rect 15669 -7602 15727 -7568
rect 15669 -7710 15727 -7676
rect 15817 -7602 15875 -7568
rect 15817 -7710 15875 -7676
rect 15965 -7602 16023 -7568
rect 15965 -7710 16023 -7676
rect 16113 -7602 16171 -7568
rect 16113 -7710 16171 -7676
rect 16261 -7602 16319 -7568
rect 16261 -7710 16319 -7676
rect 16409 -7602 16467 -7568
rect 16409 -7710 16467 -7676
rect 16557 -7602 16615 -7568
rect 16557 -7710 16615 -7676
rect 16705 -7602 16763 -7568
rect 16705 -7710 16763 -7676
rect 16853 -7602 16911 -7568
rect 16853 -7710 16911 -7676
rect 17001 -7602 17059 -7568
rect 17001 -7710 17059 -7676
rect 17149 -7602 17207 -7568
rect 17149 -7710 17207 -7676
rect 17297 -7602 17355 -7568
rect 17297 -7710 17355 -7676
rect 3075 -7801 3109 -7767
rect 3075 -7909 3109 -7875
rect 3193 -7801 3227 -7767
rect 3193 -7909 3227 -7875
rect 3311 -7801 3345 -7767
rect 3311 -7909 3345 -7875
rect 3429 -7801 3463 -7767
rect 3429 -7909 3463 -7875
rect 3547 -7801 3581 -7767
rect 3547 -7909 3581 -7875
rect 3665 -7801 3699 -7767
rect 3665 -7909 3699 -7875
rect 3783 -7801 3817 -7767
rect 3783 -7909 3817 -7875
rect 3901 -7801 3935 -7767
rect 3901 -7909 3935 -7875
rect 4019 -7801 4053 -7767
rect 4019 -7909 4053 -7875
rect 4137 -7801 4171 -7767
rect 4137 -7909 4171 -7875
rect 4255 -7801 4289 -7767
rect 4255 -7909 4289 -7875
rect 4373 -7801 4407 -7767
rect 4373 -7909 4407 -7875
rect 4491 -7801 4525 -7767
rect 4491 -7909 4525 -7875
rect 4609 -7801 4643 -7767
rect 4609 -7909 4643 -7875
rect 4727 -7801 4761 -7767
rect 4727 -7909 4761 -7875
<< locali >>
rect 7539 2006 7555 2040
rect 7589 2006 7605 2040
rect 7657 2006 7673 2040
rect 7707 2006 7723 2040
rect 7775 2006 7791 2040
rect 7825 2006 7841 2040
rect 7893 2006 7909 2040
rect 7943 2006 7959 2040
rect 8011 2006 8027 2040
rect 8061 2006 8077 2040
rect 8129 2006 8145 2040
rect 8179 2006 8195 2040
rect 8247 2006 8263 2040
rect 8297 2006 8313 2040
rect 8593 2006 8609 2040
rect 8643 2006 8659 2040
rect 8711 2006 8727 2040
rect 8761 2006 8777 2040
rect 8829 2006 8845 2040
rect 8879 2006 8895 2040
rect 8947 2006 8963 2040
rect 8997 2006 9013 2040
rect 9065 2006 9081 2040
rect 9115 2006 9131 2040
rect 9183 2006 9199 2040
rect 9233 2006 9249 2040
rect 9301 2006 9317 2040
rect 9351 2006 9367 2040
rect 9419 2006 9435 2040
rect 9469 2006 9485 2040
rect 9537 2006 9553 2040
rect 9587 2006 9603 2040
rect 9655 2006 9671 2040
rect 9705 2006 9721 2040
rect 9773 2006 9789 2040
rect 9823 2006 9839 2040
rect 9891 2006 9907 2040
rect 9941 2006 9957 2040
rect 10009 2006 10025 2040
rect 10059 2006 10075 2040
rect 10127 2006 10143 2040
rect 10177 2006 10193 2040
rect 10245 2006 10261 2040
rect 10295 2006 10311 2040
rect 12665 2005 12677 2039
rect 12711 2005 12723 2039
rect 12779 2005 12795 2039
rect 12829 2005 12845 2039
rect 12897 2005 12913 2039
rect 12947 2005 12963 2039
rect 13015 2005 13031 2039
rect 13065 2005 13081 2039
rect 13133 2005 13149 2039
rect 13183 2005 13199 2039
rect 13251 2005 13267 2039
rect 13301 2005 13317 2039
rect 13369 2005 13385 2039
rect 13419 2005 13435 2039
rect 13487 2005 13503 2039
rect 13537 2005 13553 2039
rect 13605 2005 13621 2039
rect 13655 2005 13671 2039
rect 13723 2005 13739 2039
rect 13773 2005 13789 2039
rect 13841 2005 13857 2039
rect 13891 2005 13907 2039
rect 13959 2005 13975 2039
rect 14009 2005 14025 2039
rect 14077 2005 14093 2039
rect 14127 2005 14143 2039
rect 14195 2005 14211 2039
rect 14245 2005 14261 2039
rect 14313 2005 14329 2039
rect 14363 2005 14379 2039
rect 14431 2005 14447 2039
rect 14481 2005 14497 2039
rect 14549 2005 14565 2039
rect 14599 2005 14615 2039
rect 14667 2005 14683 2039
rect 14717 2005 14733 2039
rect 14785 2005 14801 2039
rect 14835 2005 14851 2039
rect 14903 2005 14919 2039
rect 14953 2005 14969 2039
rect 15021 2005 15037 2039
rect 15071 2005 15087 2039
rect 15139 2005 15155 2039
rect 15189 2005 15205 2039
rect 15257 2005 15273 2039
rect 15307 2005 15323 2039
rect 15375 2005 15391 2039
rect 15425 2005 15441 2039
rect 15493 2005 15509 2039
rect 15543 2005 15559 2039
rect 15611 2005 15627 2039
rect 15661 2005 15677 2039
rect 15729 2005 15745 2039
rect 15779 2005 15795 2039
rect 15847 2005 15863 2039
rect 15897 2005 15913 2039
rect 15965 2005 15981 2039
rect 16015 2005 16031 2039
rect 16083 2005 16099 2039
rect 16133 2005 16149 2039
rect 16201 2005 16217 2039
rect 16251 2005 16267 2039
rect 16319 2005 16335 2039
rect 16369 2005 16385 2039
rect 16437 2005 16453 2039
rect 16487 2005 16503 2039
rect 16555 2005 16571 2039
rect 16605 2005 16621 2039
rect 16673 2005 16689 2039
rect 16723 2005 16739 2039
rect 16791 2005 16807 2039
rect 16841 2005 16857 2039
rect 16909 2005 16925 2039
rect 16959 2005 16975 2039
rect 17027 2005 17043 2039
rect 17077 2005 17093 2039
rect 17145 2005 17161 2039
rect 17195 2005 17211 2039
rect 17263 2005 17279 2039
rect 17313 2005 17329 2039
rect 17381 2005 17397 2039
rect 17431 2005 17447 2039
rect 17499 2005 17515 2039
rect 17549 2005 17565 2039
rect 17617 2005 17633 2039
rect 17667 2005 17683 2039
rect 17735 2005 17751 2039
rect 17785 2005 17801 2039
rect 17853 2005 17869 2039
rect 17903 2005 17919 2039
rect 17971 2005 17987 2039
rect 18021 2005 18037 2039
rect 18089 2005 18105 2039
rect 18139 2005 18155 2039
rect 18207 2005 18223 2039
rect 18257 2005 18273 2039
rect 18325 2005 18341 2039
rect 18375 2005 18391 2039
rect 18443 2005 18459 2039
rect 18493 2005 18509 2039
rect 18561 2005 18577 2039
rect 18611 2005 18627 2039
rect 18679 2005 18695 2039
rect 18729 2005 18745 2039
rect 18797 2005 18813 2039
rect 18847 2005 18863 2039
rect 18915 2005 18931 2039
rect 18965 2005 18981 2039
rect 19033 2005 19049 2039
rect 19083 2005 19099 2039
rect 19151 2005 19167 2039
rect 19201 2005 19217 2039
rect 19269 2005 19285 2039
rect 19319 2005 19335 2039
rect 19387 2005 19403 2039
rect 19437 2005 19453 2039
rect 19505 2005 19521 2039
rect 19555 2005 19571 2039
rect 19623 2005 19639 2039
rect 19673 2005 19689 2039
rect 19741 2005 19757 2039
rect 19791 2005 19807 2039
rect 19859 2005 19875 2039
rect 19909 2005 19925 2039
rect 19977 2005 19993 2039
rect 20027 2005 20043 2039
rect 20095 2005 20111 2039
rect 20145 2005 20161 2039
rect 20213 2005 20229 2039
rect 20263 2005 20279 2039
rect 20331 2005 20347 2039
rect 20381 2005 20397 2039
rect 20449 2005 20465 2039
rect 20499 2005 20515 2039
rect 20567 2005 20583 2039
rect 20617 2005 20633 2039
rect 20685 2005 20701 2039
rect 20735 2005 20751 2039
rect 20803 2005 20819 2039
rect 20853 2005 20869 2039
rect 20921 2005 20937 2039
rect 20971 2005 20987 2039
rect 21039 2005 21055 2039
rect 21089 2005 21105 2039
rect 21157 2005 21173 2039
rect 21207 2005 21223 2039
rect 21275 2005 21291 2039
rect 21325 2005 21341 2039
rect 12665 1897 12677 1931
rect 12711 1897 12723 1931
rect 12779 1897 12795 1931
rect 12829 1897 12845 1931
rect 12897 1897 12913 1931
rect 12947 1897 12963 1931
rect 13015 1897 13031 1931
rect 13065 1897 13081 1931
rect 13133 1897 13149 1931
rect 13183 1897 13199 1931
rect 13251 1897 13267 1931
rect 13301 1897 13317 1931
rect 13369 1897 13385 1931
rect 13419 1897 13435 1931
rect 13487 1897 13503 1931
rect 13537 1897 13553 1931
rect 13605 1897 13621 1931
rect 13655 1897 13671 1931
rect 13723 1897 13739 1931
rect 13773 1897 13789 1931
rect 13841 1897 13857 1931
rect 13891 1897 13907 1931
rect 13959 1897 13975 1931
rect 14009 1897 14025 1931
rect 14077 1897 14093 1931
rect 14127 1897 14143 1931
rect 14195 1897 14211 1931
rect 14245 1897 14261 1931
rect 14313 1897 14329 1931
rect 14363 1897 14379 1931
rect 14431 1897 14447 1931
rect 14481 1897 14497 1931
rect 14549 1897 14565 1931
rect 14599 1897 14615 1931
rect 14667 1897 14683 1931
rect 14717 1897 14733 1931
rect 14785 1897 14801 1931
rect 14835 1897 14851 1931
rect 14903 1897 14919 1931
rect 14953 1897 14969 1931
rect 15021 1897 15037 1931
rect 15071 1897 15087 1931
rect 15139 1897 15155 1931
rect 15189 1897 15205 1931
rect 15257 1897 15273 1931
rect 15307 1897 15323 1931
rect 15375 1897 15391 1931
rect 15425 1897 15441 1931
rect 15493 1897 15509 1931
rect 15543 1897 15559 1931
rect 15611 1897 15627 1931
rect 15661 1897 15677 1931
rect 15729 1897 15745 1931
rect 15779 1897 15795 1931
rect 15847 1897 15863 1931
rect 15897 1897 15913 1931
rect 15965 1897 15981 1931
rect 16015 1897 16031 1931
rect 16083 1897 16099 1931
rect 16133 1897 16149 1931
rect 16201 1897 16217 1931
rect 16251 1897 16267 1931
rect 16319 1897 16335 1931
rect 16369 1897 16385 1931
rect 16437 1897 16453 1931
rect 16487 1897 16503 1931
rect 16555 1897 16571 1931
rect 16605 1897 16621 1931
rect 16673 1897 16689 1931
rect 16723 1897 16739 1931
rect 16791 1897 16807 1931
rect 16841 1897 16857 1931
rect 16909 1897 16925 1931
rect 16959 1897 16975 1931
rect 17027 1897 17043 1931
rect 17077 1897 17093 1931
rect 17145 1897 17161 1931
rect 17195 1897 17211 1931
rect 17263 1897 17279 1931
rect 17313 1897 17329 1931
rect 17381 1897 17397 1931
rect 17431 1897 17447 1931
rect 17499 1897 17515 1931
rect 17549 1897 17565 1931
rect 17617 1897 17633 1931
rect 17667 1897 17683 1931
rect 17735 1897 17751 1931
rect 17785 1897 17801 1931
rect 17853 1897 17869 1931
rect 17903 1897 17919 1931
rect 17971 1897 17987 1931
rect 18021 1897 18037 1931
rect 18089 1897 18105 1931
rect 18139 1897 18155 1931
rect 18207 1897 18223 1931
rect 18257 1897 18273 1931
rect 18325 1897 18341 1931
rect 18375 1897 18391 1931
rect 18443 1897 18459 1931
rect 18493 1897 18509 1931
rect 18561 1897 18577 1931
rect 18611 1897 18627 1931
rect 18679 1897 18695 1931
rect 18729 1897 18745 1931
rect 18797 1897 18813 1931
rect 18847 1897 18863 1931
rect 18915 1897 18931 1931
rect 18965 1897 18981 1931
rect 19033 1897 19049 1931
rect 19083 1897 19099 1931
rect 19151 1897 19167 1931
rect 19201 1897 19217 1931
rect 19269 1897 19285 1931
rect 19319 1897 19335 1931
rect 19387 1897 19403 1931
rect 19437 1897 19453 1931
rect 19505 1897 19521 1931
rect 19555 1897 19571 1931
rect 19623 1897 19639 1931
rect 19673 1897 19689 1931
rect 19741 1897 19757 1931
rect 19791 1897 19807 1931
rect 19859 1897 19875 1931
rect 19909 1897 19925 1931
rect 19977 1897 19993 1931
rect 20027 1897 20043 1931
rect 20095 1897 20111 1931
rect 20145 1897 20161 1931
rect 20213 1897 20229 1931
rect 20263 1897 20279 1931
rect 20331 1897 20347 1931
rect 20381 1897 20397 1931
rect 20449 1897 20465 1931
rect 20499 1897 20515 1931
rect 20567 1897 20583 1931
rect 20617 1897 20633 1931
rect 20685 1897 20701 1931
rect 20735 1897 20751 1931
rect 20803 1897 20819 1931
rect 20853 1897 20869 1931
rect 20921 1897 20937 1931
rect 20971 1897 20987 1931
rect 21039 1897 21055 1931
rect 21089 1897 21105 1931
rect 21157 1897 21173 1931
rect 21207 1897 21223 1931
rect 21275 1897 21291 1931
rect 21325 1897 21341 1931
rect 1451 -182 1467 -148
rect 1501 -182 1517 -148
rect 1569 -182 1585 -148
rect 1619 -182 1635 -148
rect 1687 -182 1703 -148
rect 1737 -182 1753 -148
rect 1805 -182 1821 -148
rect 1855 -182 1871 -148
rect 1923 -182 1939 -148
rect 1973 -182 1989 -148
rect 2041 -182 2057 -148
rect 2091 -182 2107 -148
rect 2159 -182 2175 -148
rect 2209 -182 2225 -148
rect 2277 -182 2293 -148
rect 2327 -182 2343 -148
rect 2395 -182 2411 -148
rect 2445 -182 2461 -148
rect 2513 -182 2529 -148
rect 2563 -182 2579 -148
rect 2631 -182 2647 -148
rect 2681 -182 2697 -148
rect 2749 -182 2765 -148
rect 2799 -182 2815 -148
rect 2867 -182 2883 -148
rect 2917 -182 2933 -148
rect 2985 -182 3001 -148
rect 3035 -182 3051 -148
rect 3103 -182 3119 -148
rect 3153 -182 3169 -148
rect 3221 -182 3237 -148
rect 3271 -182 3287 -148
rect 3339 -182 3355 -148
rect 3389 -182 3405 -148
rect 3457 -182 3473 -148
rect 3507 -182 3523 -148
rect 3575 -182 3591 -148
rect 3625 -182 3641 -148
rect 3693 -182 3709 -148
rect 3743 -182 3759 -148
rect 3811 -182 3827 -148
rect 3861 -182 3877 -148
rect 3929 -182 3945 -148
rect 3979 -182 3995 -148
rect 4047 -182 4063 -148
rect 4097 -182 4113 -148
rect 4165 -182 4181 -148
rect 4215 -182 4231 -148
rect 4283 -182 4299 -148
rect 4333 -182 4349 -148
rect 4401 -182 4417 -148
rect 4451 -182 4467 -148
rect 4519 -182 4535 -148
rect 4569 -182 4585 -148
rect 4637 -182 4653 -148
rect 4687 -182 4703 -148
rect 4755 -182 4771 -148
rect 4805 -182 4821 -148
rect 4873 -182 4889 -148
rect 4923 -182 4939 -148
rect 4991 -182 5007 -148
rect 5041 -182 5057 -148
rect 5109 -182 5125 -148
rect 5159 -182 5175 -148
rect 5227 -182 5243 -148
rect 5277 -182 5293 -148
rect 5345 -182 5361 -148
rect 5395 -182 5411 -148
rect 5463 -182 5479 -148
rect 5513 -182 5529 -148
rect 5581 -182 5597 -148
rect 5631 -182 5647 -148
rect 5699 -182 5715 -148
rect 5749 -182 5765 -148
rect 5817 -182 5833 -148
rect 5867 -182 5883 -148
rect 5935 -182 5951 -148
rect 5985 -182 6001 -148
rect 6053 -182 6069 -148
rect 6103 -182 6119 -148
rect 6171 -182 6187 -148
rect 6221 -182 6237 -148
rect 6289 -182 6305 -148
rect 6339 -182 6355 -148
rect 6407 -182 6423 -148
rect 6457 -182 6473 -148
rect 6525 -182 6541 -148
rect 6575 -182 6591 -148
rect 6643 -182 6659 -148
rect 6693 -182 6709 -148
rect 6761 -182 6777 -148
rect 6811 -182 6827 -148
rect 6879 -182 6895 -148
rect 6929 -182 6945 -148
rect 6997 -182 7001 -148
rect 7012 -182 7013 -148
rect 7047 -182 7063 -148
rect 7130 -182 7131 -148
rect 7165 -182 7181 -148
rect 1451 -290 1467 -256
rect 1501 -290 1517 -256
rect 1569 -290 1585 -256
rect 1619 -290 1635 -256
rect 1687 -290 1703 -256
rect 1737 -290 1753 -256
rect 1805 -290 1821 -256
rect 1855 -290 1871 -256
rect 1923 -290 1939 -256
rect 1973 -290 1989 -256
rect 2041 -290 2057 -256
rect 2091 -290 2107 -256
rect 2159 -290 2175 -256
rect 2209 -290 2225 -256
rect 2277 -290 2293 -256
rect 2327 -290 2343 -256
rect 2395 -290 2411 -256
rect 2445 -290 2461 -256
rect 2513 -290 2529 -256
rect 2563 -290 2579 -256
rect 2631 -290 2647 -256
rect 2681 -290 2697 -256
rect 2749 -290 2765 -256
rect 2799 -290 2815 -256
rect 2867 -290 2883 -256
rect 2917 -290 2933 -256
rect 2985 -290 3001 -256
rect 3035 -290 3051 -256
rect 3103 -290 3119 -256
rect 3153 -290 3169 -256
rect 3221 -290 3237 -256
rect 3271 -290 3287 -256
rect 3339 -290 3355 -256
rect 3389 -290 3405 -256
rect 3457 -290 3473 -256
rect 3507 -290 3523 -256
rect 3575 -290 3591 -256
rect 3625 -290 3641 -256
rect 3693 -290 3709 -256
rect 3743 -290 3759 -256
rect 3811 -290 3827 -256
rect 3861 -290 3877 -256
rect 3929 -290 3945 -256
rect 3979 -290 3995 -256
rect 4047 -290 4063 -256
rect 4097 -290 4113 -256
rect 4165 -290 4181 -256
rect 4215 -290 4231 -256
rect 4283 -290 4299 -256
rect 4333 -290 4349 -256
rect 4401 -290 4417 -256
rect 4451 -290 4467 -256
rect 4519 -290 4535 -256
rect 4569 -290 4585 -256
rect 4637 -290 4653 -256
rect 4687 -290 4703 -256
rect 4755 -290 4771 -256
rect 4805 -290 4821 -256
rect 4873 -290 4889 -256
rect 4923 -290 4939 -256
rect 4991 -290 5007 -256
rect 5041 -290 5057 -256
rect 5109 -290 5125 -256
rect 5159 -290 5175 -256
rect 5227 -290 5243 -256
rect 5277 -290 5293 -256
rect 5345 -290 5361 -256
rect 5395 -290 5411 -256
rect 5463 -290 5479 -256
rect 5513 -290 5529 -256
rect 5581 -290 5597 -256
rect 5631 -290 5647 -256
rect 5699 -290 5715 -256
rect 5749 -290 5765 -256
rect 5817 -290 5833 -256
rect 5867 -290 5883 -256
rect 5935 -290 5951 -256
rect 5985 -290 6001 -256
rect 6053 -290 6069 -256
rect 6103 -290 6119 -256
rect 6171 -290 6187 -256
rect 6221 -290 6237 -256
rect 6289 -290 6305 -256
rect 6339 -290 6355 -256
rect 6407 -290 6423 -256
rect 6457 -290 6473 -256
rect 6525 -290 6541 -256
rect 6575 -290 6591 -256
rect 6643 -290 6659 -256
rect 6693 -290 6709 -256
rect 6761 -290 6777 -256
rect 6811 -290 6827 -256
rect 6879 -290 6895 -256
rect 6929 -290 6945 -256
rect 6997 -290 7001 -256
rect 7012 -290 7013 -256
rect 7047 -290 7063 -256
rect 7130 -290 7131 -256
rect 7165 -290 7181 -256
rect 1333 -1950 1349 -1916
rect 1383 -1950 1399 -1916
rect 1451 -1950 1467 -1916
rect 1501 -1950 1517 -1916
rect 1569 -1950 1585 -1916
rect 1619 -1950 1635 -1916
rect 1687 -1950 1703 -1916
rect 1737 -1950 1753 -1916
rect 1805 -1950 1821 -1916
rect 1855 -1950 1871 -1916
rect 1923 -1950 1939 -1916
rect 1973 -1950 1989 -1916
rect 2041 -1950 2057 -1916
rect 2091 -1950 2107 -1916
rect 2159 -1950 2175 -1916
rect 2209 -1950 2225 -1916
rect 2277 -1950 2293 -1916
rect 2327 -1950 2343 -1916
rect 2395 -1950 2411 -1916
rect 2445 -1950 2461 -1916
rect 2513 -1950 2529 -1916
rect 2563 -1950 2579 -1916
rect 2631 -1950 2647 -1916
rect 2681 -1950 2697 -1916
rect 2749 -1950 2765 -1916
rect 2799 -1950 2815 -1916
rect 2867 -1950 2883 -1916
rect 2917 -1950 2933 -1916
rect 2985 -1950 3001 -1916
rect 3035 -1950 3051 -1916
rect 3103 -1950 3119 -1916
rect 3153 -1950 3169 -1916
rect 3221 -1950 3237 -1916
rect 3271 -1950 3287 -1916
rect 3339 -1950 3355 -1916
rect 3389 -1950 3405 -1916
rect 3457 -1950 3473 -1916
rect 3507 -1950 3523 -1916
rect 3575 -1950 3591 -1916
rect 3625 -1950 3641 -1916
rect 3693 -1950 3709 -1916
rect 3743 -1950 3759 -1916
rect 3811 -1950 3827 -1916
rect 3861 -1950 3877 -1916
rect 3929 -1950 3945 -1916
rect 3979 -1950 3995 -1916
rect 4047 -1950 4063 -1916
rect 4097 -1950 4113 -1916
rect 4165 -1950 4181 -1916
rect 4215 -1950 4231 -1916
rect 4283 -1950 4299 -1916
rect 4333 -1950 4349 -1916
rect 4401 -1950 4417 -1916
rect 4451 -1950 4467 -1916
rect 4519 -1950 4535 -1916
rect 4569 -1950 4585 -1916
rect 4637 -1950 4653 -1916
rect 4687 -1950 4703 -1916
rect 4755 -1950 4771 -1916
rect 4805 -1950 4821 -1916
rect 4873 -1950 4889 -1916
rect 4923 -1950 4939 -1916
rect 4991 -1950 5007 -1916
rect 5041 -1950 5057 -1916
rect 5109 -1950 5125 -1916
rect 5159 -1950 5175 -1916
rect 5227 -1950 5243 -1916
rect 5277 -1950 5293 -1916
rect 5345 -1950 5361 -1916
rect 5395 -1950 5411 -1916
rect 5463 -1950 5479 -1916
rect 5513 -1950 5529 -1916
rect 5581 -1950 5597 -1916
rect 5631 -1950 5647 -1916
rect 5699 -1950 5715 -1916
rect 5749 -1950 5765 -1916
rect 5817 -1950 5833 -1916
rect 5867 -1950 5883 -1916
rect 5935 -1950 5951 -1916
rect 5985 -1950 6001 -1916
rect 6053 -1950 6069 -1916
rect 6103 -1950 6119 -1916
rect 6171 -1950 6187 -1916
rect 6221 -1950 6237 -1916
rect 6289 -1950 6305 -1916
rect 6339 -1950 6355 -1916
rect 6407 -1950 6423 -1916
rect 6457 -1950 6473 -1916
rect 6525 -1950 6541 -1916
rect 6575 -1950 6591 -1916
rect 6643 -1950 6659 -1916
rect 6693 -1950 6709 -1916
rect 6761 -1950 6777 -1916
rect 6811 -1950 6827 -1916
rect 6879 -1950 6895 -1916
rect 6929 -1950 6945 -1916
rect 6997 -1950 7013 -1916
rect 7047 -1950 7063 -1916
rect 7115 -1950 7131 -1916
rect 7165 -1950 7181 -1916
rect 1333 -2058 1349 -2024
rect 1383 -2058 1399 -2024
rect 1451 -2058 1467 -2024
rect 1501 -2058 1517 -2024
rect 1569 -2058 1585 -2024
rect 1619 -2058 1635 -2024
rect 1687 -2058 1703 -2024
rect 1737 -2058 1753 -2024
rect 1805 -2058 1821 -2024
rect 1855 -2058 1871 -2024
rect 1923 -2058 1939 -2024
rect 1973 -2058 1989 -2024
rect 2041 -2058 2057 -2024
rect 2091 -2058 2107 -2024
rect 2159 -2058 2175 -2024
rect 2209 -2058 2225 -2024
rect 2277 -2058 2293 -2024
rect 2327 -2058 2343 -2024
rect 2395 -2058 2411 -2024
rect 2445 -2058 2461 -2024
rect 2513 -2058 2529 -2024
rect 2563 -2058 2579 -2024
rect 2631 -2058 2647 -2024
rect 2681 -2058 2697 -2024
rect 2749 -2058 2765 -2024
rect 2799 -2058 2815 -2024
rect 2867 -2058 2883 -2024
rect 2917 -2058 2933 -2024
rect 2985 -2058 3001 -2024
rect 3035 -2058 3051 -2024
rect 3103 -2058 3119 -2024
rect 3153 -2058 3169 -2024
rect 3221 -2058 3237 -2024
rect 3271 -2058 3287 -2024
rect 3339 -2058 3355 -2024
rect 3389 -2058 3405 -2024
rect 3457 -2058 3473 -2024
rect 3507 -2058 3523 -2024
rect 3575 -2058 3591 -2024
rect 3625 -2058 3641 -2024
rect 3693 -2058 3709 -2024
rect 3743 -2058 3759 -2024
rect 3811 -2058 3827 -2024
rect 3861 -2058 3877 -2024
rect 3929 -2058 3945 -2024
rect 3979 -2058 3995 -2024
rect 4047 -2058 4063 -2024
rect 4097 -2058 4113 -2024
rect 4165 -2058 4181 -2024
rect 4215 -2058 4231 -2024
rect 4283 -2058 4299 -2024
rect 4333 -2058 4349 -2024
rect 4401 -2058 4417 -2024
rect 4451 -2058 4467 -2024
rect 4519 -2058 4535 -2024
rect 4569 -2058 4585 -2024
rect 4637 -2058 4653 -2024
rect 4687 -2058 4703 -2024
rect 4755 -2058 4771 -2024
rect 4805 -2058 4821 -2024
rect 4873 -2058 4889 -2024
rect 4923 -2058 4939 -2024
rect 4991 -2058 5007 -2024
rect 5041 -2058 5057 -2024
rect 5109 -2058 5125 -2024
rect 5159 -2058 5175 -2024
rect 5227 -2058 5243 -2024
rect 5277 -2058 5293 -2024
rect 5345 -2058 5361 -2024
rect 5395 -2058 5411 -2024
rect 5463 -2058 5479 -2024
rect 5513 -2058 5529 -2024
rect 5581 -2058 5597 -2024
rect 5631 -2058 5647 -2024
rect 5699 -2058 5715 -2024
rect 5749 -2058 5765 -2024
rect 5817 -2058 5833 -2024
rect 5867 -2058 5883 -2024
rect 5935 -2058 5951 -2024
rect 5985 -2058 6001 -2024
rect 6053 -2058 6069 -2024
rect 6103 -2058 6119 -2024
rect 6171 -2058 6187 -2024
rect 6221 -2058 6237 -2024
rect 6289 -2058 6305 -2024
rect 6339 -2058 6355 -2024
rect 6407 -2058 6423 -2024
rect 6457 -2058 6473 -2024
rect 6525 -2058 6541 -2024
rect 6575 -2058 6591 -2024
rect 6643 -2058 6659 -2024
rect 6693 -2058 6709 -2024
rect 6761 -2058 6777 -2024
rect 6811 -2058 6827 -2024
rect 6879 -2058 6895 -2024
rect 6929 -2058 6945 -2024
rect 6997 -2058 7013 -2024
rect 7047 -2058 7063 -2024
rect 7115 -2058 7131 -2024
rect 7165 -2058 7181 -2024
rect 1333 -3718 1349 -3684
rect 1383 -3718 1399 -3684
rect 1451 -3718 1467 -3684
rect 1501 -3718 1517 -3684
rect 1569 -3718 1585 -3684
rect 1619 -3718 1635 -3684
rect 1687 -3718 1703 -3684
rect 1737 -3718 1753 -3684
rect 1805 -3718 1821 -3684
rect 1855 -3718 1871 -3684
rect 1923 -3718 1939 -3684
rect 1973 -3718 1989 -3684
rect 2041 -3718 2057 -3684
rect 2091 -3718 2107 -3684
rect 2159 -3718 2175 -3684
rect 2209 -3718 2225 -3684
rect 2277 -3718 2293 -3684
rect 2327 -3718 2343 -3684
rect 2395 -3718 2411 -3684
rect 2445 -3718 2461 -3684
rect 2513 -3718 2529 -3684
rect 2563 -3718 2579 -3684
rect 2631 -3718 2647 -3684
rect 2681 -3718 2697 -3684
rect 2749 -3718 2765 -3684
rect 2799 -3718 2815 -3684
rect 2867 -3718 2883 -3684
rect 2917 -3718 2933 -3684
rect 2985 -3718 3001 -3684
rect 3035 -3718 3051 -3684
rect 3103 -3718 3119 -3684
rect 3153 -3718 3169 -3684
rect 3221 -3718 3237 -3684
rect 3271 -3718 3287 -3684
rect 3339 -3718 3355 -3684
rect 3389 -3718 3405 -3684
rect 3457 -3718 3473 -3684
rect 3507 -3718 3523 -3684
rect 3575 -3718 3591 -3684
rect 3625 -3718 3641 -3684
rect 3693 -3718 3709 -3684
rect 3743 -3718 3759 -3684
rect 3811 -3718 3827 -3684
rect 3861 -3718 3877 -3684
rect 3929 -3718 3945 -3684
rect 3979 -3718 3995 -3684
rect 4047 -3718 4063 -3684
rect 4097 -3718 4113 -3684
rect 4165 -3718 4181 -3684
rect 4215 -3718 4231 -3684
rect 4283 -3718 4299 -3684
rect 4333 -3718 4349 -3684
rect 4401 -3718 4417 -3684
rect 4451 -3718 4467 -3684
rect 4519 -3718 4535 -3684
rect 4569 -3718 4585 -3684
rect 4637 -3718 4653 -3684
rect 4687 -3718 4703 -3684
rect 4755 -3718 4771 -3684
rect 4805 -3718 4821 -3684
rect 4873 -3718 4889 -3684
rect 4923 -3718 4939 -3684
rect 4991 -3718 5007 -3684
rect 5041 -3718 5057 -3684
rect 5109 -3718 5125 -3684
rect 5159 -3718 5175 -3684
rect 5227 -3718 5243 -3684
rect 5277 -3718 5293 -3684
rect 5345 -3718 5361 -3684
rect 5395 -3718 5411 -3684
rect 5463 -3718 5479 -3684
rect 5513 -3718 5529 -3684
rect 5581 -3718 5597 -3684
rect 5631 -3718 5647 -3684
rect 5699 -3718 5715 -3684
rect 5749 -3718 5765 -3684
rect 5817 -3718 5833 -3684
rect 5867 -3718 5883 -3684
rect 5935 -3718 5951 -3684
rect 5985 -3718 6001 -3684
rect 6053 -3718 6069 -3684
rect 6103 -3718 6119 -3684
rect 6171 -3718 6187 -3684
rect 6221 -3718 6237 -3684
rect 6289 -3718 6305 -3684
rect 6339 -3718 6355 -3684
rect 6407 -3718 6423 -3684
rect 6457 -3718 6473 -3684
rect 6525 -3718 6541 -3684
rect 6575 -3718 6591 -3684
rect 6643 -3718 6659 -3684
rect 6693 -3718 6709 -3684
rect 6761 -3718 6777 -3684
rect 6811 -3718 6827 -3684
rect 6879 -3718 6895 -3684
rect 6929 -3718 6945 -3684
rect 6997 -3718 7013 -3684
rect 7047 -3718 7063 -3684
rect 7115 -3718 7131 -3684
rect 7165 -3718 7181 -3684
rect 1333 -3826 1349 -3792
rect 1383 -3826 1399 -3792
rect 1451 -3826 1467 -3792
rect 1501 -3826 1517 -3792
rect 1569 -3826 1585 -3792
rect 1619 -3826 1635 -3792
rect 1687 -3826 1703 -3792
rect 1737 -3826 1753 -3792
rect 1805 -3826 1821 -3792
rect 1855 -3826 1871 -3792
rect 1923 -3826 1939 -3792
rect 1973 -3826 1989 -3792
rect 2041 -3826 2057 -3792
rect 2091 -3826 2107 -3792
rect 2159 -3826 2175 -3792
rect 2209 -3826 2225 -3792
rect 2277 -3826 2293 -3792
rect 2327 -3826 2343 -3792
rect 2395 -3826 2411 -3792
rect 2445 -3826 2461 -3792
rect 2513 -3826 2529 -3792
rect 2563 -3826 2579 -3792
rect 2631 -3826 2647 -3792
rect 2681 -3826 2697 -3792
rect 2749 -3826 2765 -3792
rect 2799 -3826 2815 -3792
rect 2867 -3826 2883 -3792
rect 2917 -3826 2933 -3792
rect 2985 -3826 3001 -3792
rect 3035 -3826 3051 -3792
rect 3103 -3826 3119 -3792
rect 3153 -3826 3169 -3792
rect 3221 -3826 3237 -3792
rect 3271 -3826 3287 -3792
rect 3339 -3826 3355 -3792
rect 3389 -3826 3405 -3792
rect 3457 -3826 3473 -3792
rect 3507 -3826 3523 -3792
rect 3575 -3826 3591 -3792
rect 3625 -3826 3641 -3792
rect 3693 -3826 3709 -3792
rect 3743 -3826 3759 -3792
rect 3811 -3826 3827 -3792
rect 3861 -3826 3877 -3792
rect 3929 -3826 3945 -3792
rect 3979 -3826 3995 -3792
rect 4047 -3826 4063 -3792
rect 4097 -3826 4113 -3792
rect 4165 -3826 4181 -3792
rect 4215 -3826 4231 -3792
rect 4283 -3826 4299 -3792
rect 4333 -3826 4349 -3792
rect 4401 -3826 4417 -3792
rect 4451 -3826 4467 -3792
rect 4519 -3826 4535 -3792
rect 4569 -3826 4585 -3792
rect 4637 -3826 4653 -3792
rect 4687 -3826 4703 -3792
rect 4755 -3826 4771 -3792
rect 4805 -3826 4821 -3792
rect 4873 -3826 4889 -3792
rect 4923 -3826 4939 -3792
rect 4991 -3826 5007 -3792
rect 5041 -3826 5057 -3792
rect 5109 -3826 5125 -3792
rect 5159 -3826 5175 -3792
rect 5227 -3826 5243 -3792
rect 5277 -3826 5293 -3792
rect 5345 -3826 5361 -3792
rect 5395 -3826 5411 -3792
rect 5463 -3826 5479 -3792
rect 5513 -3826 5529 -3792
rect 5581 -3826 5597 -3792
rect 5631 -3826 5647 -3792
rect 5699 -3826 5715 -3792
rect 5749 -3826 5765 -3792
rect 5817 -3826 5833 -3792
rect 5867 -3826 5883 -3792
rect 5935 -3826 5951 -3792
rect 5985 -3826 6001 -3792
rect 6053 -3826 6069 -3792
rect 6103 -3826 6119 -3792
rect 6171 -3826 6187 -3792
rect 6221 -3826 6237 -3792
rect 6289 -3826 6305 -3792
rect 6339 -3826 6355 -3792
rect 6407 -3826 6423 -3792
rect 6457 -3826 6473 -3792
rect 6525 -3826 6541 -3792
rect 6575 -3826 6591 -3792
rect 6643 -3826 6659 -3792
rect 6693 -3826 6709 -3792
rect 6761 -3826 6777 -3792
rect 6811 -3826 6827 -3792
rect 6879 -3826 6895 -3792
rect 6929 -3826 6945 -3792
rect 6997 -3826 7013 -3792
rect 7047 -3826 7063 -3792
rect 7115 -3826 7131 -3792
rect 7165 -3826 7181 -3792
rect 1333 -5486 1349 -5452
rect 1383 -5486 1399 -5452
rect 1451 -5486 1467 -5452
rect 1501 -5486 1517 -5452
rect 1569 -5486 1585 -5452
rect 1619 -5486 1635 -5452
rect 1687 -5486 1703 -5452
rect 1737 -5486 1753 -5452
rect 1805 -5486 1821 -5452
rect 1855 -5486 1871 -5452
rect 1923 -5486 1939 -5452
rect 1973 -5486 1989 -5452
rect 2041 -5486 2057 -5452
rect 2091 -5486 2107 -5452
rect 2159 -5486 2175 -5452
rect 2209 -5486 2225 -5452
rect 2277 -5486 2293 -5452
rect 2327 -5486 2343 -5452
rect 2395 -5486 2411 -5452
rect 2445 -5486 2461 -5452
rect 2513 -5486 2529 -5452
rect 2563 -5486 2579 -5452
rect 2631 -5486 2647 -5452
rect 2681 -5486 2697 -5452
rect 2749 -5486 2765 -5452
rect 2799 -5486 2815 -5452
rect 2867 -5486 2883 -5452
rect 2917 -5486 2933 -5452
rect 2985 -5486 3001 -5452
rect 3035 -5486 3051 -5452
rect 3103 -5486 3119 -5452
rect 3153 -5486 3169 -5452
rect 3221 -5486 3237 -5452
rect 3271 -5486 3287 -5452
rect 3339 -5486 3355 -5452
rect 3389 -5486 3405 -5452
rect 3457 -5486 3473 -5452
rect 3507 -5486 3523 -5452
rect 3575 -5486 3591 -5452
rect 3625 -5486 3641 -5452
rect 3693 -5486 3709 -5452
rect 3743 -5486 3759 -5452
rect 3811 -5486 3827 -5452
rect 3861 -5486 3877 -5452
rect 3929 -5486 3945 -5452
rect 3979 -5486 3995 -5452
rect 4047 -5486 4063 -5452
rect 4097 -5486 4113 -5452
rect 4165 -5486 4181 -5452
rect 4215 -5486 4231 -5452
rect 4283 -5486 4299 -5452
rect 4333 -5486 4349 -5452
rect 4401 -5486 4417 -5452
rect 4451 -5486 4467 -5452
rect 4519 -5486 4535 -5452
rect 4569 -5486 4585 -5452
rect 4637 -5486 4653 -5452
rect 4687 -5486 4703 -5452
rect 4755 -5486 4771 -5452
rect 4805 -5486 4821 -5452
rect 4873 -5486 4889 -5452
rect 4923 -5486 4939 -5452
rect 4991 -5486 5007 -5452
rect 5041 -5486 5057 -5452
rect 5109 -5486 5125 -5452
rect 5159 -5486 5175 -5452
rect 5227 -5486 5243 -5452
rect 5277 -5486 5293 -5452
rect 5345 -5486 5361 -5452
rect 5395 -5486 5411 -5452
rect 5463 -5486 5479 -5452
rect 5513 -5486 5529 -5452
rect 5581 -5486 5597 -5452
rect 5631 -5486 5647 -5452
rect 5699 -5486 5715 -5452
rect 5749 -5486 5765 -5452
rect 5817 -5486 5833 -5452
rect 5867 -5486 5883 -5452
rect 5935 -5486 5951 -5452
rect 5985 -5486 6001 -5452
rect 6053 -5486 6069 -5452
rect 6103 -5486 6119 -5452
rect 6171 -5486 6187 -5452
rect 6221 -5486 6237 -5452
rect 6289 -5486 6305 -5452
rect 6339 -5486 6355 -5452
rect 6407 -5486 6423 -5452
rect 6457 -5486 6473 -5452
rect 6525 -5486 6541 -5452
rect 6575 -5486 6591 -5452
rect 6643 -5486 6659 -5452
rect 6693 -5486 6709 -5452
rect 6761 -5486 6777 -5452
rect 6811 -5486 6827 -5452
rect 6879 -5486 6895 -5452
rect 6929 -5486 6945 -5452
rect 6997 -5486 7013 -5452
rect 7047 -5486 7063 -5452
rect 7115 -5486 7131 -5452
rect 7165 -5486 7181 -5452
rect 1333 -5594 1349 -5560
rect 1383 -5594 1399 -5560
rect 1451 -5594 1467 -5560
rect 1501 -5594 1517 -5560
rect 1569 -5594 1585 -5560
rect 1619 -5594 1635 -5560
rect 1687 -5594 1703 -5560
rect 1737 -5594 1753 -5560
rect 1805 -5594 1821 -5560
rect 1855 -5594 1871 -5560
rect 1923 -5594 1939 -5560
rect 1973 -5594 1989 -5560
rect 2041 -5594 2057 -5560
rect 2091 -5594 2107 -5560
rect 2159 -5594 2175 -5560
rect 2209 -5594 2225 -5560
rect 2277 -5594 2293 -5560
rect 2327 -5594 2343 -5560
rect 2395 -5594 2411 -5560
rect 2445 -5594 2461 -5560
rect 2513 -5594 2529 -5560
rect 2563 -5594 2579 -5560
rect 2631 -5594 2647 -5560
rect 2681 -5594 2697 -5560
rect 2749 -5594 2765 -5560
rect 2799 -5594 2815 -5560
rect 2867 -5594 2883 -5560
rect 2917 -5594 2933 -5560
rect 2985 -5594 3001 -5560
rect 3035 -5594 3051 -5560
rect 3103 -5594 3119 -5560
rect 3153 -5594 3169 -5560
rect 3221 -5594 3237 -5560
rect 3271 -5594 3287 -5560
rect 3339 -5594 3355 -5560
rect 3389 -5594 3405 -5560
rect 3457 -5594 3473 -5560
rect 3507 -5594 3523 -5560
rect 3575 -5594 3591 -5560
rect 3625 -5594 3641 -5560
rect 3693 -5594 3709 -5560
rect 3743 -5594 3759 -5560
rect 3811 -5594 3827 -5560
rect 3861 -5594 3877 -5560
rect 3929 -5594 3945 -5560
rect 3979 -5594 3995 -5560
rect 4047 -5594 4063 -5560
rect 4097 -5594 4113 -5560
rect 4165 -5594 4181 -5560
rect 4215 -5594 4231 -5560
rect 4283 -5594 4299 -5560
rect 4333 -5594 4349 -5560
rect 4401 -5594 4417 -5560
rect 4451 -5594 4467 -5560
rect 4519 -5594 4535 -5560
rect 4569 -5594 4585 -5560
rect 4637 -5594 4653 -5560
rect 4687 -5594 4703 -5560
rect 4755 -5594 4771 -5560
rect 4805 -5594 4821 -5560
rect 4873 -5594 4889 -5560
rect 4923 -5594 4939 -5560
rect 4991 -5594 5007 -5560
rect 5041 -5594 5057 -5560
rect 5109 -5594 5125 -5560
rect 5159 -5594 5175 -5560
rect 5227 -5594 5243 -5560
rect 5277 -5594 5293 -5560
rect 5345 -5594 5361 -5560
rect 5395 -5594 5411 -5560
rect 5463 -5594 5479 -5560
rect 5513 -5594 5529 -5560
rect 5581 -5594 5597 -5560
rect 5631 -5594 5647 -5560
rect 5699 -5594 5715 -5560
rect 5749 -5594 5765 -5560
rect 5817 -5594 5833 -5560
rect 5867 -5594 5883 -5560
rect 5935 -5594 5951 -5560
rect 5985 -5594 6001 -5560
rect 6053 -5594 6069 -5560
rect 6103 -5594 6119 -5560
rect 6171 -5594 6187 -5560
rect 6221 -5594 6237 -5560
rect 6289 -5594 6305 -5560
rect 6339 -5594 6355 -5560
rect 6407 -5594 6423 -5560
rect 6457 -5594 6473 -5560
rect 6525 -5594 6541 -5560
rect 6575 -5594 6591 -5560
rect 6643 -5594 6659 -5560
rect 6693 -5594 6709 -5560
rect 6761 -5594 6777 -5560
rect 6811 -5594 6827 -5560
rect 6879 -5594 6895 -5560
rect 6929 -5594 6945 -5560
rect 6997 -5594 7013 -5560
rect 7047 -5594 7063 -5560
rect 7115 -5594 7131 -5560
rect 7165 -5594 7181 -5560
rect 11657 -7602 11673 -7568
rect 11731 -7602 11747 -7568
rect 11805 -7602 11821 -7568
rect 11879 -7602 11895 -7568
rect 11953 -7602 11969 -7568
rect 12027 -7602 12043 -7568
rect 12101 -7602 12117 -7568
rect 12175 -7602 12191 -7568
rect 12249 -7602 12265 -7568
rect 12323 -7602 12339 -7568
rect 12397 -7602 12413 -7568
rect 12471 -7602 12487 -7568
rect 12545 -7602 12561 -7568
rect 12619 -7602 12635 -7568
rect 12693 -7602 12709 -7568
rect 12767 -7602 12783 -7568
rect 12841 -7602 12857 -7568
rect 12915 -7602 12931 -7568
rect 12989 -7602 13005 -7568
rect 13063 -7602 13079 -7568
rect 13137 -7602 13153 -7568
rect 13211 -7602 13227 -7568
rect 13285 -7602 13301 -7568
rect 13359 -7602 13375 -7568
rect 13433 -7602 13449 -7568
rect 13507 -7602 13523 -7568
rect 13581 -7602 13597 -7568
rect 13655 -7602 13671 -7568
rect 13729 -7602 13745 -7568
rect 13803 -7602 13819 -7568
rect 13877 -7602 13893 -7568
rect 13951 -7602 13967 -7568
rect 14025 -7602 14041 -7568
rect 14099 -7602 14115 -7568
rect 14173 -7602 14189 -7568
rect 14247 -7602 14263 -7568
rect 14321 -7602 14337 -7568
rect 14395 -7602 14411 -7568
rect 14469 -7602 14485 -7568
rect 14543 -7602 14559 -7568
rect 14617 -7602 14633 -7568
rect 14691 -7602 14707 -7568
rect 14765 -7602 14781 -7568
rect 14839 -7602 14855 -7568
rect 14913 -7602 14929 -7568
rect 14987 -7602 15003 -7568
rect 15061 -7602 15077 -7568
rect 15135 -7602 15151 -7568
rect 15209 -7602 15225 -7568
rect 15283 -7602 15299 -7568
rect 15357 -7602 15373 -7568
rect 15431 -7602 15447 -7568
rect 15505 -7602 15521 -7568
rect 15579 -7602 15595 -7568
rect 15653 -7602 15669 -7568
rect 15727 -7602 15743 -7568
rect 15801 -7602 15817 -7568
rect 15875 -7602 15891 -7568
rect 15949 -7602 15965 -7568
rect 16023 -7602 16039 -7568
rect 16097 -7602 16113 -7568
rect 16171 -7602 16187 -7568
rect 16245 -7602 16261 -7568
rect 16319 -7602 16335 -7568
rect 16393 -7602 16409 -7568
rect 16467 -7602 16483 -7568
rect 16541 -7602 16557 -7568
rect 16615 -7602 16631 -7568
rect 16689 -7602 16705 -7568
rect 16763 -7602 16779 -7568
rect 16837 -7602 16853 -7568
rect 16911 -7602 16927 -7568
rect 16985 -7602 17001 -7568
rect 17059 -7602 17075 -7568
rect 17133 -7602 17149 -7568
rect 17207 -7602 17223 -7568
rect 17281 -7602 17297 -7568
rect 17355 -7602 17371 -7568
rect 17429 -7602 17445 -7568
rect 17503 -7602 17519 -7568
rect 17577 -7602 17593 -7568
rect 17651 -7602 17667 -7568
rect 17725 -7602 17741 -7568
rect 17799 -7602 17815 -7568
rect 17873 -7602 17889 -7568
rect 17947 -7602 17963 -7568
rect 18021 -7602 18037 -7568
rect 18095 -7602 18111 -7568
rect 18169 -7602 18185 -7568
rect 18243 -7602 18259 -7568
rect 18317 -7602 18333 -7568
rect 18391 -7602 18407 -7568
rect 18465 -7602 18481 -7568
rect 18539 -7602 18555 -7568
rect 18613 -7602 18629 -7568
rect 18687 -7602 18703 -7568
rect 18761 -7602 18777 -7568
rect 18835 -7602 18851 -7568
rect 18909 -7602 18925 -7568
rect 18983 -7602 18999 -7568
rect 19057 -7602 19073 -7568
rect 19131 -7602 19147 -7568
rect 19205 -7602 19221 -7568
rect 19279 -7602 19295 -7568
rect 19353 -7602 19369 -7568
rect 19427 -7602 19443 -7568
rect 19501 -7602 19517 -7568
rect 19575 -7602 19591 -7568
rect 19649 -7602 19665 -7568
rect 19723 -7602 19739 -7568
rect 19797 -7602 19813 -7568
rect 19871 -7602 19887 -7568
rect 19945 -7602 19961 -7568
rect 20019 -7602 20035 -7568
rect 20093 -7602 20109 -7568
rect 20167 -7602 20183 -7568
rect 20241 -7602 20257 -7568
rect 20315 -7602 20331 -7568
rect 20389 -7602 20405 -7568
rect 20463 -7602 20479 -7568
rect 20537 -7602 20553 -7568
rect 20611 -7602 20627 -7568
rect 20685 -7602 20701 -7568
rect 20759 -7602 20775 -7568
rect 20833 -7602 20849 -7568
rect 20907 -7602 20923 -7568
rect 20981 -7602 20997 -7568
rect 21055 -7602 21071 -7568
rect 21129 -7602 21145 -7568
rect 21203 -7602 21219 -7568
rect 21277 -7602 21293 -7568
rect 21351 -7602 21367 -7568
rect 21425 -7602 21441 -7568
rect 21499 -7602 21515 -7568
rect 21573 -7602 21589 -7568
rect 21647 -7602 21663 -7568
rect 21721 -7602 21737 -7568
rect 21795 -7602 21811 -7568
rect 21869 -7602 21885 -7568
rect 21943 -7602 21959 -7568
rect 22017 -7602 22033 -7568
rect 22091 -7602 22107 -7568
rect 22165 -7602 22181 -7568
rect 22239 -7602 22255 -7568
rect 22313 -7602 22329 -7568
rect 22387 -7602 22403 -7568
rect 22461 -7602 22477 -7568
rect 22535 -7602 22551 -7568
rect 11657 -7710 11673 -7676
rect 11731 -7710 11747 -7676
rect 11805 -7710 11821 -7676
rect 11879 -7710 11895 -7676
rect 11953 -7710 11969 -7676
rect 12027 -7710 12043 -7676
rect 12101 -7710 12117 -7676
rect 12175 -7710 12191 -7676
rect 12249 -7710 12265 -7676
rect 12323 -7710 12339 -7676
rect 12397 -7710 12413 -7676
rect 12471 -7710 12487 -7676
rect 12545 -7710 12561 -7676
rect 12619 -7710 12635 -7676
rect 12693 -7710 12709 -7676
rect 12767 -7710 12783 -7676
rect 12841 -7710 12857 -7676
rect 12915 -7710 12931 -7676
rect 12989 -7710 13005 -7676
rect 13063 -7710 13079 -7676
rect 13137 -7710 13153 -7676
rect 13211 -7710 13227 -7676
rect 13285 -7710 13301 -7676
rect 13359 -7710 13375 -7676
rect 13433 -7710 13449 -7676
rect 13507 -7710 13523 -7676
rect 13581 -7710 13597 -7676
rect 13655 -7710 13671 -7676
rect 13729 -7710 13745 -7676
rect 13803 -7710 13819 -7676
rect 13877 -7710 13893 -7676
rect 13951 -7710 13967 -7676
rect 14025 -7710 14041 -7676
rect 14099 -7710 14115 -7676
rect 14173 -7710 14189 -7676
rect 14247 -7710 14263 -7676
rect 14321 -7710 14337 -7676
rect 14395 -7710 14411 -7676
rect 14469 -7710 14485 -7676
rect 14543 -7710 14559 -7676
rect 14617 -7710 14633 -7676
rect 14691 -7710 14707 -7676
rect 14765 -7710 14781 -7676
rect 14839 -7710 14855 -7676
rect 14913 -7710 14929 -7676
rect 14987 -7710 15003 -7676
rect 15061 -7710 15077 -7676
rect 15135 -7710 15151 -7676
rect 15209 -7710 15225 -7676
rect 15283 -7710 15299 -7676
rect 15357 -7710 15373 -7676
rect 15431 -7710 15447 -7676
rect 15505 -7710 15521 -7676
rect 15579 -7710 15595 -7676
rect 15653 -7710 15669 -7676
rect 15727 -7710 15743 -7676
rect 15801 -7710 15817 -7676
rect 15875 -7710 15891 -7676
rect 15949 -7710 15965 -7676
rect 16023 -7710 16039 -7676
rect 16097 -7710 16113 -7676
rect 16171 -7710 16187 -7676
rect 16245 -7710 16261 -7676
rect 16319 -7710 16335 -7676
rect 16393 -7710 16409 -7676
rect 16467 -7710 16483 -7676
rect 16541 -7710 16557 -7676
rect 16615 -7710 16631 -7676
rect 16689 -7710 16705 -7676
rect 16763 -7710 16779 -7676
rect 16837 -7710 16853 -7676
rect 16911 -7710 16927 -7676
rect 16985 -7710 17001 -7676
rect 17059 -7710 17075 -7676
rect 17133 -7710 17149 -7676
rect 17207 -7710 17223 -7676
rect 17281 -7710 17297 -7676
rect 17355 -7710 17371 -7676
rect 17429 -7710 17445 -7676
rect 17503 -7710 17519 -7676
rect 17577 -7710 17593 -7676
rect 17651 -7710 17667 -7676
rect 17725 -7710 17741 -7676
rect 17799 -7710 17815 -7676
rect 17873 -7710 17889 -7676
rect 17947 -7710 17963 -7676
rect 18021 -7710 18037 -7676
rect 18095 -7710 18111 -7676
rect 18169 -7710 18185 -7676
rect 18243 -7710 18259 -7676
rect 18317 -7710 18333 -7676
rect 18391 -7710 18407 -7676
rect 18465 -7710 18481 -7676
rect 18539 -7710 18555 -7676
rect 18613 -7710 18629 -7676
rect 18687 -7710 18703 -7676
rect 18761 -7710 18777 -7676
rect 18835 -7710 18851 -7676
rect 18909 -7710 18925 -7676
rect 18983 -7710 18999 -7676
rect 19057 -7710 19073 -7676
rect 19131 -7710 19147 -7676
rect 19205 -7710 19221 -7676
rect 19279 -7710 19295 -7676
rect 19353 -7710 19369 -7676
rect 19427 -7710 19443 -7676
rect 19501 -7710 19517 -7676
rect 19575 -7710 19591 -7676
rect 19649 -7710 19665 -7676
rect 19723 -7710 19739 -7676
rect 19797 -7710 19813 -7676
rect 19871 -7710 19887 -7676
rect 19945 -7710 19961 -7676
rect 20019 -7710 20035 -7676
rect 20093 -7710 20109 -7676
rect 20167 -7710 20183 -7676
rect 20241 -7710 20257 -7676
rect 20315 -7710 20331 -7676
rect 20389 -7710 20405 -7676
rect 20463 -7710 20479 -7676
rect 20537 -7710 20553 -7676
rect 20611 -7710 20627 -7676
rect 20685 -7710 20701 -7676
rect 20759 -7710 20775 -7676
rect 20833 -7710 20849 -7676
rect 20907 -7710 20923 -7676
rect 20981 -7710 20997 -7676
rect 21055 -7710 21071 -7676
rect 21129 -7710 21145 -7676
rect 21203 -7710 21219 -7676
rect 21277 -7710 21293 -7676
rect 21351 -7710 21367 -7676
rect 21425 -7710 21441 -7676
rect 21499 -7710 21515 -7676
rect 21573 -7710 21589 -7676
rect 21647 -7710 21663 -7676
rect 21721 -7710 21737 -7676
rect 21795 -7710 21811 -7676
rect 21869 -7710 21885 -7676
rect 21943 -7710 21959 -7676
rect 22017 -7710 22033 -7676
rect 22091 -7710 22107 -7676
rect 22165 -7710 22181 -7676
rect 22239 -7710 22255 -7676
rect 22313 -7710 22329 -7676
rect 22387 -7710 22403 -7676
rect 22461 -7710 22477 -7676
rect 22535 -7710 22551 -7676
rect 3059 -7801 3075 -7767
rect 3109 -7801 3125 -7767
rect 3177 -7801 3193 -7767
rect 3227 -7801 3243 -7767
rect 3295 -7801 3311 -7767
rect 3345 -7801 3361 -7767
rect 3413 -7801 3429 -7767
rect 3463 -7801 3479 -7767
rect 3531 -7801 3547 -7767
rect 3581 -7801 3597 -7767
rect 3649 -7801 3665 -7767
rect 3699 -7801 3715 -7767
rect 3767 -7801 3783 -7767
rect 3817 -7801 3833 -7767
rect 3885 -7801 3901 -7767
rect 3935 -7801 3951 -7767
rect 4003 -7801 4019 -7767
rect 4053 -7801 4069 -7767
rect 4121 -7801 4137 -7767
rect 4171 -7801 4187 -7767
rect 4239 -7801 4255 -7767
rect 4289 -7801 4305 -7767
rect 4357 -7801 4373 -7767
rect 4407 -7801 4423 -7767
rect 4475 -7801 4491 -7767
rect 4525 -7801 4541 -7767
rect 4593 -7801 4609 -7767
rect 4643 -7801 4659 -7767
rect 4711 -7801 4727 -7767
rect 4761 -7801 4777 -7767
rect 5057 -7801 5073 -7767
rect 5107 -7801 5123 -7767
rect 5175 -7801 5191 -7767
rect 5225 -7801 5241 -7767
rect 5293 -7801 5309 -7767
rect 5343 -7801 5359 -7767
rect 5411 -7801 5427 -7767
rect 5461 -7801 5477 -7767
rect 5529 -7801 5545 -7767
rect 5579 -7801 5595 -7767
rect 5647 -7801 5663 -7767
rect 5697 -7801 5713 -7767
rect 5765 -7801 5781 -7767
rect 5815 -7801 5831 -7767
rect 5883 -7801 5899 -7767
rect 5933 -7801 5949 -7767
rect 6001 -7801 6017 -7767
rect 6051 -7801 6067 -7767
rect 6119 -7801 6135 -7767
rect 6169 -7801 6185 -7767
rect 6237 -7801 6253 -7767
rect 6287 -7801 6303 -7767
rect 6355 -7801 6371 -7767
rect 6405 -7801 6421 -7767
rect 6473 -7801 6489 -7767
rect 6523 -7801 6539 -7767
rect 6591 -7801 6607 -7767
rect 6641 -7801 6657 -7767
rect 6709 -7801 6725 -7767
rect 6759 -7801 6775 -7767
rect 3059 -7909 3075 -7875
rect 3109 -7909 3125 -7875
rect 3177 -7909 3193 -7875
rect 3227 -7909 3243 -7875
rect 3295 -7909 3311 -7875
rect 3345 -7909 3361 -7875
rect 3413 -7909 3429 -7875
rect 3463 -7909 3479 -7875
rect 3531 -7909 3547 -7875
rect 3581 -7909 3597 -7875
rect 3649 -7909 3665 -7875
rect 3699 -7909 3715 -7875
rect 3767 -7909 3783 -7875
rect 3817 -7909 3833 -7875
rect 3885 -7909 3901 -7875
rect 3935 -7909 3951 -7875
rect 4003 -7909 4019 -7875
rect 4053 -7909 4069 -7875
rect 4121 -7909 4137 -7875
rect 4171 -7909 4187 -7875
rect 4239 -7909 4255 -7875
rect 4289 -7909 4305 -7875
rect 4357 -7909 4373 -7875
rect 4407 -7909 4423 -7875
rect 4475 -7909 4491 -7875
rect 4525 -7909 4541 -7875
rect 4593 -7909 4609 -7875
rect 4643 -7909 4659 -7875
rect 4711 -7909 4727 -7875
rect 4761 -7909 4777 -7875
rect 5057 -7909 5073 -7875
rect 5107 -7909 5123 -7875
rect 5175 -7909 5191 -7875
rect 5225 -7909 5241 -7875
rect 5293 -7909 5309 -7875
rect 5343 -7909 5359 -7875
rect 5411 -7909 5427 -7875
rect 5461 -7909 5477 -7875
rect 5529 -7909 5545 -7875
rect 5579 -7909 5595 -7875
rect 5647 -7909 5663 -7875
rect 5697 -7909 5713 -7875
rect 5765 -7909 5781 -7875
rect 5815 -7909 5831 -7875
rect 5883 -7909 5899 -7875
rect 5933 -7909 5949 -7875
rect 6001 -7909 6017 -7875
rect 6051 -7909 6067 -7875
rect 6119 -7909 6135 -7875
rect 6169 -7909 6185 -7875
rect 6237 -7909 6253 -7875
rect 6287 -7909 6303 -7875
rect 6355 -7909 6371 -7875
rect 6405 -7909 6421 -7875
rect 6473 -7909 6489 -7875
rect 6523 -7909 6539 -7875
rect 6591 -7909 6607 -7875
rect 6641 -7909 6657 -7875
rect 6709 -7909 6725 -7875
rect 6759 -7909 6775 -7875
<< viali >>
rect 6788 2099 6822 2675
rect 4613 2006 4647 2040
rect 4731 2006 4765 2040
rect 4849 2006 4883 2040
rect 4967 2006 5001 2040
rect 5085 2006 5119 2040
rect 5203 2006 5237 2040
rect 5321 2006 5355 2040
rect 5439 2006 5473 2040
rect 5557 2006 5591 2040
rect 5675 2006 5709 2040
rect 5793 2006 5827 2040
rect 5911 2006 5945 2040
rect 6029 2006 6063 2040
rect 6147 2006 6181 2040
rect 6265 2006 6299 2040
rect 6847 2006 6881 2040
rect 6965 2006 6999 2040
rect 7083 2006 7117 2040
rect 7201 2006 7235 2040
rect 7319 2006 7353 2040
rect 7437 2006 7471 2040
rect 7555 2006 7589 2040
rect 7673 2006 7707 2040
rect 7791 2006 7825 2040
rect 7909 2006 7943 2040
rect 8027 2006 8061 2040
rect 8145 2006 8179 2040
rect 8263 2006 8297 2040
rect 8609 2006 8643 2040
rect 8727 2006 8761 2040
rect 8845 2006 8879 2040
rect 8963 2006 8997 2040
rect 9081 2006 9115 2040
rect 9199 2006 9233 2040
rect 9317 2006 9351 2040
rect 9435 2006 9469 2040
rect 9553 2006 9587 2040
rect 9671 2006 9705 2040
rect 9789 2006 9823 2040
rect 9907 2006 9941 2040
rect 10025 2006 10059 2040
rect 10143 2006 10177 2040
rect 10261 2006 10295 2040
rect 12677 2005 12711 2039
rect 12795 2005 12829 2039
rect 12913 2005 12947 2039
rect 13031 2005 13065 2039
rect 13149 2005 13183 2039
rect 13267 2005 13301 2039
rect 13385 2005 13419 2039
rect 13503 2005 13537 2039
rect 13621 2005 13655 2039
rect 13739 2005 13773 2039
rect 13857 2005 13891 2039
rect 13975 2005 14009 2039
rect 14093 2005 14127 2039
rect 14211 2005 14245 2039
rect 14329 2005 14363 2039
rect 14447 2005 14481 2039
rect 14565 2005 14599 2039
rect 14683 2005 14717 2039
rect 14801 2005 14835 2039
rect 14919 2005 14953 2039
rect 15037 2005 15071 2039
rect 15155 2005 15189 2039
rect 15273 2005 15307 2039
rect 15391 2005 15425 2039
rect 15509 2005 15543 2039
rect 15627 2005 15661 2039
rect 15745 2005 15779 2039
rect 15863 2005 15897 2039
rect 15981 2005 16015 2039
rect 16099 2005 16133 2039
rect 16217 2005 16251 2039
rect 16335 2005 16369 2039
rect 16453 2005 16487 2039
rect 16571 2005 16605 2039
rect 16689 2005 16723 2039
rect 16807 2005 16841 2039
rect 16925 2005 16959 2039
rect 17043 2005 17077 2039
rect 17161 2005 17195 2039
rect 17279 2005 17313 2039
rect 17397 2005 17431 2039
rect 17515 2005 17549 2039
rect 17633 2005 17667 2039
rect 17751 2005 17785 2039
rect 17869 2005 17903 2039
rect 17987 2005 18021 2039
rect 18105 2005 18139 2039
rect 18223 2005 18257 2039
rect 18341 2005 18375 2039
rect 18459 2005 18493 2039
rect 18577 2005 18611 2039
rect 18695 2005 18729 2039
rect 18813 2005 18847 2039
rect 18931 2005 18965 2039
rect 19049 2005 19083 2039
rect 19167 2005 19201 2039
rect 19285 2005 19319 2039
rect 19403 2005 19437 2039
rect 19521 2005 19555 2039
rect 19639 2005 19673 2039
rect 19757 2005 19791 2039
rect 19875 2005 19909 2039
rect 19993 2005 20027 2039
rect 20111 2005 20145 2039
rect 20229 2005 20263 2039
rect 20347 2005 20381 2039
rect 20465 2005 20499 2039
rect 20583 2005 20617 2039
rect 20701 2005 20735 2039
rect 20819 2005 20853 2039
rect 20937 2005 20971 2039
rect 21055 2005 21089 2039
rect 21173 2005 21207 2039
rect 21291 2005 21325 2039
rect 12677 1897 12711 1931
rect 12795 1897 12829 1931
rect 12913 1897 12947 1931
rect 13031 1897 13065 1931
rect 13149 1897 13183 1931
rect 13267 1897 13301 1931
rect 13385 1897 13419 1931
rect 13503 1897 13537 1931
rect 13621 1897 13655 1931
rect 13739 1897 13773 1931
rect 13857 1897 13891 1931
rect 13975 1897 14009 1931
rect 14093 1897 14127 1931
rect 14211 1897 14245 1931
rect 14329 1897 14363 1931
rect 14447 1897 14481 1931
rect 14565 1897 14599 1931
rect 14683 1897 14717 1931
rect 14801 1897 14835 1931
rect 14919 1897 14953 1931
rect 15037 1897 15071 1931
rect 15155 1897 15189 1931
rect 15273 1897 15307 1931
rect 15391 1897 15425 1931
rect 15509 1897 15543 1931
rect 15627 1897 15661 1931
rect 15745 1897 15779 1931
rect 15863 1897 15897 1931
rect 15981 1897 16015 1931
rect 16099 1897 16133 1931
rect 16217 1897 16251 1931
rect 16335 1897 16369 1931
rect 16453 1897 16487 1931
rect 16571 1897 16605 1931
rect 16689 1897 16723 1931
rect 16807 1897 16841 1931
rect 16925 1897 16959 1931
rect 17043 1897 17077 1931
rect 17161 1897 17195 1931
rect 17279 1897 17313 1931
rect 17397 1897 17431 1931
rect 17515 1897 17549 1931
rect 17633 1897 17667 1931
rect 17751 1897 17785 1931
rect 17869 1897 17903 1931
rect 17987 1897 18021 1931
rect 18105 1897 18139 1931
rect 18223 1897 18257 1931
rect 18341 1897 18375 1931
rect 18459 1897 18493 1931
rect 18577 1897 18611 1931
rect 18695 1897 18729 1931
rect 18813 1897 18847 1931
rect 18931 1897 18965 1931
rect 19049 1897 19083 1931
rect 19167 1897 19201 1931
rect 19285 1897 19319 1931
rect 19403 1897 19437 1931
rect 19521 1897 19555 1931
rect 19639 1897 19673 1931
rect 19757 1897 19791 1931
rect 19875 1897 19909 1931
rect 19993 1897 20027 1931
rect 20111 1897 20145 1931
rect 20229 1897 20263 1931
rect 20347 1897 20381 1931
rect 20465 1897 20499 1931
rect 20583 1897 20617 1931
rect 20701 1897 20735 1931
rect 20819 1897 20853 1931
rect 20937 1897 20971 1931
rect 21055 1897 21089 1931
rect 21173 1897 21207 1931
rect 21291 1897 21325 1931
rect 1467 -182 1501 -148
rect 1585 -182 1619 -148
rect 1703 -182 1737 -148
rect 1821 -182 1855 -148
rect 1939 -182 1973 -148
rect 2057 -182 2091 -148
rect 2175 -182 2209 -148
rect 2293 -182 2327 -148
rect 2411 -182 2445 -148
rect 2529 -182 2563 -148
rect 2647 -182 2681 -148
rect 2765 -182 2799 -148
rect 2883 -182 2917 -148
rect 3001 -182 3035 -148
rect 3119 -182 3153 -148
rect 3237 -182 3271 -148
rect 3355 -182 3389 -148
rect 3473 -182 3507 -148
rect 3591 -182 3625 -148
rect 3709 -182 3743 -148
rect 3827 -182 3861 -148
rect 3945 -182 3979 -148
rect 4063 -182 4097 -148
rect 4181 -182 4215 -148
rect 4299 -182 4333 -148
rect 4417 -182 4451 -148
rect 4535 -182 4569 -148
rect 4653 -182 4687 -148
rect 4771 -182 4805 -148
rect 4889 -182 4923 -148
rect 5007 -182 5041 -148
rect 5125 -182 5159 -148
rect 5243 -182 5277 -148
rect 5361 -182 5395 -148
rect 5479 -182 5513 -148
rect 5597 -182 5631 -148
rect 5715 -182 5749 -148
rect 5833 -182 5867 -148
rect 5951 -182 5985 -148
rect 6069 -182 6103 -148
rect 6187 -182 6221 -148
rect 6305 -182 6339 -148
rect 6423 -182 6457 -148
rect 6541 -182 6575 -148
rect 6659 -182 6693 -148
rect 6777 -182 6811 -148
rect 6895 -182 6929 -148
rect 7013 -182 7047 -148
rect 7131 -182 7165 -148
rect 1467 -290 1501 -256
rect 1585 -290 1619 -256
rect 1703 -290 1737 -256
rect 1821 -290 1855 -256
rect 1939 -290 1973 -256
rect 2057 -290 2091 -256
rect 2175 -290 2209 -256
rect 2293 -290 2327 -256
rect 2411 -290 2445 -256
rect 2529 -290 2563 -256
rect 2647 -290 2681 -256
rect 2765 -290 2799 -256
rect 2883 -290 2917 -256
rect 3001 -290 3035 -256
rect 3119 -290 3153 -256
rect 3237 -290 3271 -256
rect 3355 -290 3389 -256
rect 3473 -290 3507 -256
rect 3591 -290 3625 -256
rect 3709 -290 3743 -256
rect 3827 -290 3861 -256
rect 3945 -290 3979 -256
rect 4063 -290 4097 -256
rect 4181 -290 4215 -256
rect 4299 -290 4333 -256
rect 4417 -290 4451 -256
rect 4535 -290 4569 -256
rect 4653 -290 4687 -256
rect 4771 -290 4805 -256
rect 4889 -290 4923 -256
rect 5007 -290 5041 -256
rect 5125 -290 5159 -256
rect 5243 -290 5277 -256
rect 5361 -290 5395 -256
rect 5479 -290 5513 -256
rect 5597 -290 5631 -256
rect 5715 -290 5749 -256
rect 5833 -290 5867 -256
rect 5951 -290 5985 -256
rect 6069 -290 6103 -256
rect 6187 -290 6221 -256
rect 6305 -290 6339 -256
rect 6423 -290 6457 -256
rect 6541 -290 6575 -256
rect 6659 -290 6693 -256
rect 6777 -290 6811 -256
rect 6895 -290 6929 -256
rect 7013 -290 7047 -256
rect 7131 -290 7165 -256
rect 1349 -1950 1383 -1916
rect 1467 -1950 1501 -1916
rect 1585 -1950 1619 -1916
rect 1703 -1950 1737 -1916
rect 1821 -1950 1855 -1916
rect 1939 -1950 1973 -1916
rect 2057 -1950 2091 -1916
rect 2175 -1950 2209 -1916
rect 2293 -1950 2327 -1916
rect 2411 -1950 2445 -1916
rect 2529 -1950 2563 -1916
rect 2647 -1950 2681 -1916
rect 2765 -1950 2799 -1916
rect 2883 -1950 2917 -1916
rect 3001 -1950 3035 -1916
rect 3119 -1950 3153 -1916
rect 3237 -1950 3271 -1916
rect 3355 -1950 3389 -1916
rect 3473 -1950 3507 -1916
rect 3591 -1950 3625 -1916
rect 3709 -1950 3743 -1916
rect 3827 -1950 3861 -1916
rect 3945 -1950 3979 -1916
rect 4063 -1950 4097 -1916
rect 4181 -1950 4215 -1916
rect 4299 -1950 4333 -1916
rect 4417 -1950 4451 -1916
rect 4535 -1950 4569 -1916
rect 4653 -1950 4687 -1916
rect 4771 -1950 4805 -1916
rect 4889 -1950 4923 -1916
rect 5007 -1950 5041 -1916
rect 5125 -1950 5159 -1916
rect 5243 -1950 5277 -1916
rect 5361 -1950 5395 -1916
rect 5479 -1950 5513 -1916
rect 5597 -1950 5631 -1916
rect 5715 -1950 5749 -1916
rect 5833 -1950 5867 -1916
rect 5951 -1950 5985 -1916
rect 6069 -1950 6103 -1916
rect 6187 -1950 6221 -1916
rect 6305 -1950 6339 -1916
rect 6423 -1950 6457 -1916
rect 6541 -1950 6575 -1916
rect 6659 -1950 6693 -1916
rect 6777 -1950 6811 -1916
rect 6895 -1950 6929 -1916
rect 7013 -1950 7047 -1916
rect 7131 -1950 7165 -1916
rect 1349 -2058 1383 -2024
rect 1467 -2058 1501 -2024
rect 1585 -2058 1619 -2024
rect 1703 -2058 1737 -2024
rect 1821 -2058 1855 -2024
rect 1939 -2058 1973 -2024
rect 2057 -2058 2091 -2024
rect 2175 -2058 2209 -2024
rect 2293 -2058 2327 -2024
rect 2411 -2058 2445 -2024
rect 2529 -2058 2563 -2024
rect 2647 -2058 2681 -2024
rect 2765 -2058 2799 -2024
rect 2883 -2058 2917 -2024
rect 3001 -2058 3035 -2024
rect 3119 -2058 3153 -2024
rect 3237 -2058 3271 -2024
rect 3355 -2058 3389 -2024
rect 3473 -2058 3507 -2024
rect 3591 -2058 3625 -2024
rect 3709 -2058 3743 -2024
rect 3827 -2058 3861 -2024
rect 3945 -2058 3979 -2024
rect 4063 -2058 4097 -2024
rect 4181 -2058 4215 -2024
rect 4299 -2058 4333 -2024
rect 4417 -2058 4451 -2024
rect 4535 -2058 4569 -2024
rect 4653 -2058 4687 -2024
rect 4771 -2058 4805 -2024
rect 4889 -2058 4923 -2024
rect 5007 -2058 5041 -2024
rect 5125 -2058 5159 -2024
rect 5243 -2058 5277 -2024
rect 5361 -2058 5395 -2024
rect 5479 -2058 5513 -2024
rect 5597 -2058 5631 -2024
rect 5715 -2058 5749 -2024
rect 5833 -2058 5867 -2024
rect 5951 -2058 5985 -2024
rect 6069 -2058 6103 -2024
rect 6187 -2058 6221 -2024
rect 6305 -2058 6339 -2024
rect 6423 -2058 6457 -2024
rect 6541 -2058 6575 -2024
rect 6659 -2058 6693 -2024
rect 6777 -2058 6811 -2024
rect 6895 -2058 6929 -2024
rect 7013 -2058 7047 -2024
rect 7131 -2058 7165 -2024
rect 1349 -3718 1383 -3684
rect 1467 -3718 1501 -3684
rect 1585 -3718 1619 -3684
rect 1703 -3718 1737 -3684
rect 1821 -3718 1855 -3684
rect 1939 -3718 1973 -3684
rect 2057 -3718 2091 -3684
rect 2175 -3718 2209 -3684
rect 2293 -3718 2327 -3684
rect 2411 -3718 2445 -3684
rect 2529 -3718 2563 -3684
rect 2647 -3718 2681 -3684
rect 2765 -3718 2799 -3684
rect 2883 -3718 2917 -3684
rect 3001 -3718 3035 -3684
rect 3119 -3718 3153 -3684
rect 3237 -3718 3271 -3684
rect 3355 -3718 3389 -3684
rect 3473 -3718 3507 -3684
rect 3591 -3718 3625 -3684
rect 3709 -3718 3743 -3684
rect 3827 -3718 3861 -3684
rect 3945 -3718 3979 -3684
rect 4063 -3718 4097 -3684
rect 4181 -3718 4215 -3684
rect 4299 -3718 4333 -3684
rect 4417 -3718 4451 -3684
rect 4535 -3718 4569 -3684
rect 4653 -3718 4687 -3684
rect 4771 -3718 4805 -3684
rect 4889 -3718 4923 -3684
rect 5007 -3718 5041 -3684
rect 5125 -3718 5159 -3684
rect 5243 -3718 5277 -3684
rect 5361 -3718 5395 -3684
rect 5479 -3718 5513 -3684
rect 5597 -3718 5631 -3684
rect 5715 -3718 5749 -3684
rect 5833 -3718 5867 -3684
rect 5951 -3718 5985 -3684
rect 6069 -3718 6103 -3684
rect 6187 -3718 6221 -3684
rect 6305 -3718 6339 -3684
rect 6423 -3718 6457 -3684
rect 6541 -3718 6575 -3684
rect 6659 -3718 6693 -3684
rect 6777 -3718 6811 -3684
rect 6895 -3718 6929 -3684
rect 7013 -3718 7047 -3684
rect 7131 -3718 7165 -3684
rect 1349 -3826 1383 -3792
rect 1467 -3826 1501 -3792
rect 1585 -3826 1619 -3792
rect 1703 -3826 1737 -3792
rect 1821 -3826 1855 -3792
rect 1939 -3826 1973 -3792
rect 2057 -3826 2091 -3792
rect 2175 -3826 2209 -3792
rect 2293 -3826 2327 -3792
rect 2411 -3826 2445 -3792
rect 2529 -3826 2563 -3792
rect 2647 -3826 2681 -3792
rect 2765 -3826 2799 -3792
rect 2883 -3826 2917 -3792
rect 3001 -3826 3035 -3792
rect 3119 -3826 3153 -3792
rect 3237 -3826 3271 -3792
rect 3355 -3826 3389 -3792
rect 3473 -3826 3507 -3792
rect 3591 -3826 3625 -3792
rect 3709 -3826 3743 -3792
rect 3827 -3826 3861 -3792
rect 3945 -3826 3979 -3792
rect 4063 -3826 4097 -3792
rect 4181 -3826 4215 -3792
rect 4299 -3826 4333 -3792
rect 4417 -3826 4451 -3792
rect 4535 -3826 4569 -3792
rect 4653 -3826 4687 -3792
rect 4771 -3826 4805 -3792
rect 4889 -3826 4923 -3792
rect 5007 -3826 5041 -3792
rect 5125 -3826 5159 -3792
rect 5243 -3826 5277 -3792
rect 5361 -3826 5395 -3792
rect 5479 -3826 5513 -3792
rect 5597 -3826 5631 -3792
rect 5715 -3826 5749 -3792
rect 5833 -3826 5867 -3792
rect 5951 -3826 5985 -3792
rect 6069 -3826 6103 -3792
rect 6187 -3826 6221 -3792
rect 6305 -3826 6339 -3792
rect 6423 -3826 6457 -3792
rect 6541 -3826 6575 -3792
rect 6659 -3826 6693 -3792
rect 6777 -3826 6811 -3792
rect 6895 -3826 6929 -3792
rect 7013 -3826 7047 -3792
rect 7131 -3826 7165 -3792
rect 1349 -5486 1383 -5452
rect 1467 -5486 1501 -5452
rect 1585 -5486 1619 -5452
rect 1703 -5486 1737 -5452
rect 1821 -5486 1855 -5452
rect 1939 -5486 1973 -5452
rect 2057 -5486 2091 -5452
rect 2175 -5486 2209 -5452
rect 2293 -5486 2327 -5452
rect 2411 -5486 2445 -5452
rect 2529 -5486 2563 -5452
rect 2647 -5486 2681 -5452
rect 2765 -5486 2799 -5452
rect 2883 -5486 2917 -5452
rect 3001 -5486 3035 -5452
rect 3119 -5486 3153 -5452
rect 3237 -5486 3271 -5452
rect 3355 -5486 3389 -5452
rect 3473 -5486 3507 -5452
rect 3591 -5486 3625 -5452
rect 3709 -5486 3743 -5452
rect 3827 -5486 3861 -5452
rect 3945 -5486 3979 -5452
rect 4063 -5486 4097 -5452
rect 4181 -5486 4215 -5452
rect 4299 -5486 4333 -5452
rect 4417 -5486 4451 -5452
rect 4535 -5486 4569 -5452
rect 4653 -5486 4687 -5452
rect 4771 -5486 4805 -5452
rect 4889 -5486 4923 -5452
rect 5007 -5486 5041 -5452
rect 5125 -5486 5159 -5452
rect 5243 -5486 5277 -5452
rect 5361 -5486 5395 -5452
rect 5479 -5486 5513 -5452
rect 5597 -5486 5631 -5452
rect 5715 -5486 5749 -5452
rect 5833 -5486 5867 -5452
rect 5951 -5486 5985 -5452
rect 6069 -5486 6103 -5452
rect 6187 -5486 6221 -5452
rect 6305 -5486 6339 -5452
rect 6423 -5486 6457 -5452
rect 6541 -5486 6575 -5452
rect 6659 -5486 6693 -5452
rect 6777 -5486 6811 -5452
rect 6895 -5486 6929 -5452
rect 7013 -5486 7047 -5452
rect 7131 -5486 7165 -5452
rect 1349 -5594 1383 -5560
rect 1467 -5594 1501 -5560
rect 1585 -5594 1619 -5560
rect 1703 -5594 1737 -5560
rect 1821 -5594 1855 -5560
rect 1939 -5594 1973 -5560
rect 2057 -5594 2091 -5560
rect 2175 -5594 2209 -5560
rect 2293 -5594 2327 -5560
rect 2411 -5594 2445 -5560
rect 2529 -5594 2563 -5560
rect 2647 -5594 2681 -5560
rect 2765 -5594 2799 -5560
rect 2883 -5594 2917 -5560
rect 3001 -5594 3035 -5560
rect 3119 -5594 3153 -5560
rect 3237 -5594 3271 -5560
rect 3355 -5594 3389 -5560
rect 3473 -5594 3507 -5560
rect 3591 -5594 3625 -5560
rect 3709 -5594 3743 -5560
rect 3827 -5594 3861 -5560
rect 3945 -5594 3979 -5560
rect 4063 -5594 4097 -5560
rect 4181 -5594 4215 -5560
rect 4299 -5594 4333 -5560
rect 4417 -5594 4451 -5560
rect 4535 -5594 4569 -5560
rect 4653 -5594 4687 -5560
rect 4771 -5594 4805 -5560
rect 4889 -5594 4923 -5560
rect 5007 -5594 5041 -5560
rect 5125 -5594 5159 -5560
rect 5243 -5594 5277 -5560
rect 5361 -5594 5395 -5560
rect 5479 -5594 5513 -5560
rect 5597 -5594 5631 -5560
rect 5715 -5594 5749 -5560
rect 5833 -5594 5867 -5560
rect 5951 -5594 5985 -5560
rect 6069 -5594 6103 -5560
rect 6187 -5594 6221 -5560
rect 6305 -5594 6339 -5560
rect 6423 -5594 6457 -5560
rect 6541 -5594 6575 -5560
rect 6659 -5594 6693 -5560
rect 6777 -5594 6811 -5560
rect 6895 -5594 6929 -5560
rect 7013 -5594 7047 -5560
rect 7131 -5594 7165 -5560
rect 11463 -7518 11497 -6642
rect 11611 -7518 11645 -6642
rect 11759 -7518 11793 -6642
rect 11907 -7518 11941 -6642
rect 12055 -7518 12089 -6642
rect 12203 -7518 12237 -6642
rect 12351 -7518 12385 -6642
rect 12499 -7518 12533 -6642
rect 12647 -7518 12681 -6642
rect 12795 -7518 12829 -6642
rect 12943 -7518 12977 -6642
rect 13091 -7518 13125 -6642
rect 13239 -7518 13273 -6642
rect 13387 -7518 13421 -6642
rect 13535 -7518 13569 -6642
rect 13683 -7518 13717 -6642
rect 13831 -7518 13865 -6642
rect 13979 -7518 14013 -6642
rect 14127 -7518 14161 -6642
rect 14275 -7518 14309 -6642
rect 14423 -7518 14457 -6642
rect 14571 -7518 14605 -6642
rect 14719 -7518 14753 -6642
rect 14867 -7518 14901 -6642
rect 15015 -7518 15049 -6642
rect 15163 -7518 15197 -6642
rect 15311 -7518 15345 -6642
rect 15459 -7518 15493 -6642
rect 15607 -7518 15641 -6642
rect 15755 -7518 15789 -6642
rect 15903 -7518 15937 -6642
rect 16051 -7518 16085 -6642
rect 16199 -7518 16233 -6642
rect 16347 -7518 16381 -6642
rect 16495 -7518 16529 -6642
rect 16643 -7518 16677 -6642
rect 16791 -7518 16825 -6642
rect 16939 -7518 16973 -6642
rect 17087 -7518 17121 -6642
rect 17235 -7518 17269 -6642
rect 17383 -7518 17417 -6642
rect 17531 -7518 17565 -6642
rect 17679 -7518 17713 -6642
rect 17827 -7518 17861 -6642
rect 17975 -7518 18009 -6642
rect 18123 -7518 18157 -6642
rect 18271 -7518 18305 -6642
rect 18419 -7518 18453 -6642
rect 18567 -7518 18601 -6642
rect 18715 -7518 18749 -6642
rect 18863 -7518 18897 -6642
rect 19011 -7518 19045 -6642
rect 19159 -7518 19193 -6642
rect 19307 -7518 19341 -6642
rect 19455 -7518 19489 -6642
rect 19603 -7518 19637 -6642
rect 19751 -7518 19785 -6642
rect 19899 -7518 19933 -6642
rect 20047 -7518 20081 -6642
rect 20195 -7518 20229 -6642
rect 20343 -7518 20377 -6642
rect 20491 -7518 20525 -6642
rect 20639 -7518 20673 -6642
rect 20787 -7518 20821 -6642
rect 20935 -7518 20969 -6642
rect 21083 -7518 21117 -6642
rect 21231 -7518 21265 -6642
rect 21379 -7518 21413 -6642
rect 21527 -7518 21561 -6642
rect 21675 -7518 21709 -6642
rect 21823 -7518 21857 -6642
rect 21971 -7518 22005 -6642
rect 22119 -7518 22153 -6642
rect 22267 -7518 22301 -6642
rect 22563 -7518 22597 -6642
rect 11673 -7602 11731 -7568
rect 11821 -7602 11879 -7568
rect 11969 -7602 12027 -7568
rect 12117 -7602 12175 -7568
rect 12265 -7602 12323 -7568
rect 12413 -7602 12471 -7568
rect 12561 -7602 12619 -7568
rect 12709 -7602 12767 -7568
rect 12857 -7602 12915 -7568
rect 13005 -7602 13063 -7568
rect 13153 -7602 13211 -7568
rect 13301 -7602 13359 -7568
rect 13449 -7602 13507 -7568
rect 13597 -7602 13655 -7568
rect 13745 -7602 13803 -7568
rect 13893 -7602 13951 -7568
rect 14041 -7602 14099 -7568
rect 14189 -7602 14247 -7568
rect 14337 -7602 14395 -7568
rect 14485 -7602 14543 -7568
rect 14633 -7602 14691 -7568
rect 14781 -7602 14839 -7568
rect 14929 -7602 14987 -7568
rect 15077 -7602 15135 -7568
rect 15225 -7602 15283 -7568
rect 15373 -7602 15431 -7568
rect 15521 -7602 15579 -7568
rect 15669 -7602 15727 -7568
rect 15817 -7602 15875 -7568
rect 15965 -7602 16023 -7568
rect 16113 -7602 16171 -7568
rect 16261 -7602 16319 -7568
rect 16409 -7602 16467 -7568
rect 16557 -7602 16615 -7568
rect 16705 -7602 16763 -7568
rect 16853 -7602 16911 -7568
rect 17001 -7602 17059 -7568
rect 17149 -7602 17207 -7568
rect 17297 -7602 17355 -7568
rect 17445 -7602 17503 -7568
rect 17593 -7602 17651 -7568
rect 17741 -7602 17799 -7568
rect 17889 -7602 17947 -7568
rect 18037 -7602 18095 -7568
rect 18185 -7602 18243 -7568
rect 18333 -7602 18391 -7568
rect 18481 -7602 18539 -7568
rect 18629 -7602 18687 -7568
rect 18777 -7602 18835 -7568
rect 18925 -7602 18983 -7568
rect 19073 -7602 19131 -7568
rect 19221 -7602 19279 -7568
rect 19369 -7602 19427 -7568
rect 19517 -7602 19575 -7568
rect 19665 -7602 19723 -7568
rect 19813 -7602 19871 -7568
rect 19961 -7602 20019 -7568
rect 20109 -7602 20167 -7568
rect 20257 -7602 20315 -7568
rect 20405 -7602 20463 -7568
rect 20553 -7602 20611 -7568
rect 20701 -7602 20759 -7568
rect 20849 -7602 20907 -7568
rect 20997 -7602 21055 -7568
rect 21145 -7602 21203 -7568
rect 21293 -7602 21351 -7568
rect 21441 -7602 21499 -7568
rect 21589 -7602 21647 -7568
rect 21737 -7602 21795 -7568
rect 21885 -7602 21943 -7568
rect 22033 -7602 22091 -7568
rect 22181 -7602 22239 -7568
rect 22329 -7602 22387 -7568
rect 22477 -7602 22535 -7568
rect 11673 -7710 11731 -7676
rect 11821 -7710 11879 -7676
rect 11969 -7710 12027 -7676
rect 12117 -7710 12175 -7676
rect 12265 -7710 12323 -7676
rect 12413 -7710 12471 -7676
rect 12561 -7710 12619 -7676
rect 12709 -7710 12767 -7676
rect 12857 -7710 12915 -7676
rect 13005 -7710 13063 -7676
rect 13153 -7710 13211 -7676
rect 13301 -7710 13359 -7676
rect 13449 -7710 13507 -7676
rect 13597 -7710 13655 -7676
rect 13745 -7710 13803 -7676
rect 13893 -7710 13951 -7676
rect 14041 -7710 14099 -7676
rect 14189 -7710 14247 -7676
rect 14337 -7710 14395 -7676
rect 14485 -7710 14543 -7676
rect 14633 -7710 14691 -7676
rect 14781 -7710 14839 -7676
rect 14929 -7710 14987 -7676
rect 15077 -7710 15135 -7676
rect 15225 -7710 15283 -7676
rect 15373 -7710 15431 -7676
rect 15521 -7710 15579 -7676
rect 15669 -7710 15727 -7676
rect 15817 -7710 15875 -7676
rect 15965 -7710 16023 -7676
rect 16113 -7710 16171 -7676
rect 16261 -7710 16319 -7676
rect 16409 -7710 16467 -7676
rect 16557 -7710 16615 -7676
rect 16705 -7710 16763 -7676
rect 16853 -7710 16911 -7676
rect 17001 -7710 17059 -7676
rect 17149 -7710 17207 -7676
rect 17297 -7710 17355 -7676
rect 17445 -7710 17503 -7676
rect 17593 -7710 17651 -7676
rect 17741 -7710 17799 -7676
rect 17889 -7710 17947 -7676
rect 18037 -7710 18095 -7676
rect 18185 -7710 18243 -7676
rect 18333 -7710 18391 -7676
rect 18481 -7710 18539 -7676
rect 18629 -7710 18687 -7676
rect 18777 -7710 18835 -7676
rect 18925 -7710 18983 -7676
rect 19073 -7710 19131 -7676
rect 19221 -7710 19279 -7676
rect 19369 -7710 19427 -7676
rect 19517 -7710 19575 -7676
rect 19665 -7710 19723 -7676
rect 19813 -7710 19871 -7676
rect 19961 -7710 20019 -7676
rect 20109 -7710 20167 -7676
rect 20257 -7710 20315 -7676
rect 20405 -7710 20463 -7676
rect 20553 -7710 20611 -7676
rect 20701 -7710 20759 -7676
rect 20849 -7710 20907 -7676
rect 20997 -7710 21055 -7676
rect 21145 -7710 21203 -7676
rect 21293 -7710 21351 -7676
rect 21441 -7710 21499 -7676
rect 21589 -7710 21647 -7676
rect 21737 -7710 21795 -7676
rect 21885 -7710 21943 -7676
rect 22033 -7710 22091 -7676
rect 22181 -7710 22239 -7676
rect 22329 -7710 22387 -7676
rect 22477 -7710 22535 -7676
rect 3075 -7801 3109 -7767
rect 3193 -7801 3227 -7767
rect 3311 -7801 3345 -7767
rect 3429 -7801 3463 -7767
rect 3547 -7801 3581 -7767
rect 3665 -7801 3699 -7767
rect 3783 -7801 3817 -7767
rect 3901 -7801 3935 -7767
rect 4019 -7801 4053 -7767
rect 4137 -7801 4171 -7767
rect 4255 -7801 4289 -7767
rect 4373 -7801 4407 -7767
rect 4491 -7801 4525 -7767
rect 4609 -7801 4643 -7767
rect 4727 -7801 4761 -7767
rect 5073 -7801 5107 -7767
rect 5191 -7801 5225 -7767
rect 5309 -7801 5343 -7767
rect 5427 -7801 5461 -7767
rect 5545 -7801 5579 -7767
rect 5663 -7801 5697 -7767
rect 5781 -7801 5815 -7767
rect 5899 -7801 5933 -7767
rect 6017 -7801 6051 -7767
rect 6135 -7801 6169 -7767
rect 6253 -7801 6287 -7767
rect 6371 -7801 6405 -7767
rect 6489 -7801 6523 -7767
rect 6607 -7801 6641 -7767
rect 6725 -7801 6759 -7767
rect 3075 -7909 3109 -7875
rect 3193 -7909 3227 -7875
rect 3311 -7909 3345 -7875
rect 3429 -7909 3463 -7875
rect 3547 -7909 3581 -7875
rect 3665 -7909 3699 -7875
rect 3783 -7909 3817 -7875
rect 3901 -7909 3935 -7875
rect 4019 -7909 4053 -7875
rect 4137 -7909 4171 -7875
rect 4255 -7909 4289 -7875
rect 4373 -7909 4407 -7875
rect 4491 -7909 4525 -7875
rect 4609 -7909 4643 -7875
rect 4727 -7909 4761 -7875
rect 5073 -7909 5107 -7875
rect 5191 -7909 5225 -7875
rect 5309 -7909 5343 -7875
rect 5427 -7909 5461 -7875
rect 5545 -7909 5579 -7875
rect 5663 -7909 5697 -7875
rect 5781 -7909 5815 -7875
rect 5899 -7909 5933 -7875
rect 6017 -7909 6051 -7875
rect 6135 -7909 6169 -7875
rect 6253 -7909 6287 -7875
rect 6371 -7909 6405 -7875
rect 6489 -7909 6523 -7875
rect 6607 -7909 6641 -7875
rect 6725 -7909 6759 -7875
rect 11463 -8636 11497 -7760
rect 11611 -8636 11645 -7760
rect 11759 -8636 11793 -7760
rect 11907 -8636 11941 -7760
rect 12055 -8636 12089 -7760
rect 12203 -8636 12237 -7760
rect 12351 -8636 12385 -7760
rect 12499 -8636 12533 -7760
rect 12647 -8636 12681 -7760
rect 12795 -8636 12829 -7760
rect 12943 -8636 12977 -7760
rect 13091 -8636 13125 -7760
rect 13239 -8636 13273 -7760
rect 13387 -8636 13421 -7760
rect 13535 -8636 13569 -7760
rect 13683 -8636 13717 -7760
rect 13831 -8636 13865 -7760
rect 13979 -8636 14013 -7760
rect 14127 -8636 14161 -7760
rect 14275 -8636 14309 -7760
rect 14423 -8636 14457 -7760
rect 14571 -8636 14605 -7760
rect 14719 -8636 14753 -7760
rect 14867 -8636 14901 -7760
rect 15015 -8636 15049 -7760
rect 15163 -8636 15197 -7760
rect 15311 -8636 15345 -7760
rect 15459 -8636 15493 -7760
rect 15607 -8636 15641 -7760
rect 15755 -8636 15789 -7760
rect 15903 -8636 15937 -7760
rect 16051 -8636 16085 -7760
rect 16199 -8636 16233 -7760
rect 16347 -8636 16381 -7760
rect 16495 -8636 16529 -7760
rect 16643 -8636 16677 -7760
rect 16791 -8636 16825 -7760
rect 16939 -8636 16973 -7760
rect 17087 -8636 17121 -7760
rect 17235 -8636 17269 -7760
rect 17383 -8636 17417 -7760
rect 17531 -8636 17565 -7760
rect 17679 -8636 17713 -7760
rect 17827 -8636 17861 -7760
rect 17975 -8636 18009 -7760
rect 18123 -8636 18157 -7760
rect 18271 -8636 18305 -7760
rect 18419 -8636 18453 -7760
rect 18567 -8636 18601 -7760
rect 18715 -8636 18749 -7760
rect 18863 -8636 18897 -7760
rect 19011 -8636 19045 -7760
rect 19159 -8636 19193 -7760
rect 19307 -8636 19341 -7760
rect 19455 -8636 19489 -7760
rect 19603 -8636 19637 -7760
rect 19751 -8636 19785 -7760
rect 19899 -8636 19933 -7760
rect 20047 -8636 20081 -7760
rect 20195 -8636 20229 -7760
rect 20343 -8636 20377 -7760
rect 20491 -8636 20525 -7760
rect 20639 -8636 20673 -7760
rect 20787 -8636 20821 -7760
rect 20935 -8636 20969 -7760
rect 21083 -8636 21117 -7760
rect 21231 -8636 21265 -7760
rect 21379 -8636 21413 -7760
rect 21527 -8636 21561 -7760
rect 21675 -8636 21709 -7760
rect 21823 -8636 21857 -7760
rect 21971 -8636 22005 -7760
rect 22119 -8636 22153 -7760
rect 22267 -8636 22301 -7760
<< metal1 >>
rect 6520 2087 6530 2687
rect 6582 2087 6592 2687
rect 6664 2087 6700 2099
rect 6756 2087 6766 2687
rect 6818 2675 6828 2687
rect 6822 2099 6828 2675
rect 6818 2087 6828 2099
rect 4601 2044 4659 2046
rect 4719 2044 4777 2046
rect 4837 2044 4895 2046
rect 4955 2044 5013 2046
rect 5073 2044 5131 2046
rect 5191 2044 5249 2046
rect 5309 2044 5367 2046
rect 5427 2044 5485 2046
rect 5545 2044 5603 2046
rect 5663 2044 5721 2046
rect 5781 2044 5839 2046
rect 5899 2044 5957 2046
rect 6017 2044 6075 2046
rect 6135 2044 6193 2046
rect 6253 2044 6311 2046
rect 6835 2044 6893 2046
rect 6953 2044 7011 2046
rect 7071 2044 7129 2046
rect 7189 2044 7247 2046
rect 7307 2044 7365 2046
rect 7425 2044 7483 2046
rect 7543 2044 7601 2046
rect 7661 2044 7719 2046
rect 7779 2044 7837 2046
rect 7897 2044 7955 2046
rect 8015 2044 8073 2046
rect 8133 2044 8191 2046
rect 8251 2044 8309 2046
rect 8597 2044 8655 2046
rect 8715 2044 8773 2046
rect 8833 2044 8891 2046
rect 8951 2044 9009 2046
rect 9069 2044 9127 2046
rect 9187 2044 9245 2046
rect 9305 2044 9363 2046
rect 9423 2044 9481 2046
rect 9541 2044 9599 2046
rect 9659 2044 9717 2046
rect 9777 2044 9835 2046
rect 9895 2044 9953 2046
rect 10013 2044 10071 2046
rect 10131 2044 10189 2046
rect 10249 2044 10307 2046
rect 4591 1952 4601 2044
rect 4659 1952 4669 2044
rect 4709 1952 4719 2044
rect 4777 1952 4787 2044
rect 4827 1952 4837 2044
rect 4895 1952 4905 2044
rect 4945 1952 4955 2044
rect 5013 1952 5023 2044
rect 5063 1952 5073 2044
rect 5131 1952 5141 2044
rect 5181 1952 5191 2044
rect 5249 1952 5259 2044
rect 5299 1952 5309 2044
rect 5367 1952 5377 2044
rect 5417 1952 5427 2044
rect 5485 1952 5495 2044
rect 5535 1952 5545 2044
rect 5603 1952 5613 2044
rect 5653 1952 5663 2044
rect 5721 1952 5731 2044
rect 5771 1952 5781 2044
rect 5839 1952 5849 2044
rect 5889 1952 5899 2044
rect 5957 1952 5967 2044
rect 6007 1952 6017 2044
rect 6075 1952 6085 2044
rect 6125 1952 6135 2044
rect 6193 1952 6203 2044
rect 6243 1952 6253 2044
rect 6311 1952 6321 2044
rect 6589 1952 6599 2044
rect 6657 1952 6667 2044
rect 6707 1952 6717 2044
rect 6775 1952 6785 2044
rect 6825 1952 6835 2044
rect 6893 1952 6903 2044
rect 6943 1952 6953 2044
rect 7011 1952 7021 2044
rect 7061 1952 7071 2044
rect 7129 1952 7139 2044
rect 7179 1952 7189 2044
rect 7247 1952 7257 2044
rect 7297 1952 7307 2044
rect 7365 1952 7375 2044
rect 7415 1952 7425 2044
rect 7483 1952 7493 2044
rect 7533 1952 7543 2044
rect 7601 1952 7611 2044
rect 7651 1952 7661 2044
rect 7719 1952 7729 2044
rect 7769 1952 7779 2044
rect 7837 1952 7847 2044
rect 7887 1952 7897 2044
rect 7955 1952 7965 2044
rect 8005 1952 8015 2044
rect 8073 1952 8083 2044
rect 8123 1952 8133 2044
rect 8191 1952 8201 2044
rect 8241 1952 8251 2044
rect 8309 1952 8319 2044
rect 8587 1952 8597 2044
rect 8655 1952 8665 2044
rect 8705 1952 8715 2044
rect 8773 1952 8783 2044
rect 8823 1952 8833 2044
rect 8891 1952 8901 2044
rect 8941 1952 8951 2044
rect 9009 1952 9019 2044
rect 9059 1952 9069 2044
rect 9127 1952 9137 2044
rect 9177 1952 9187 2044
rect 9245 1952 9255 2044
rect 9295 1952 9305 2044
rect 9363 1952 9373 2044
rect 9413 1952 9423 2044
rect 9481 1952 9491 2044
rect 9531 1952 9541 2044
rect 9599 1952 9609 2044
rect 9649 1952 9659 2044
rect 9717 1952 9727 2044
rect 9767 1952 9777 2044
rect 9835 1952 9845 2044
rect 9885 1952 9895 2044
rect 9953 1952 9963 2044
rect 10003 1952 10013 2044
rect 10071 1952 10081 2044
rect 10121 1952 10131 2044
rect 10189 1952 10199 2044
rect 10239 1952 10249 2044
rect 10307 1952 10317 2044
rect 12537 1891 12547 2045
rect 12605 1891 12615 2045
rect 12655 1891 12665 2045
rect 12723 1891 12733 2045
rect 12773 1891 12783 2045
rect 12841 1891 12851 2045
rect 12891 1891 12901 2045
rect 12959 1891 12969 2045
rect 13009 1891 13019 2045
rect 13077 1891 13087 2045
rect 13127 1891 13137 2045
rect 13195 1891 13205 2045
rect 13245 1891 13255 2045
rect 13313 1891 13323 2045
rect 13363 1891 13373 2045
rect 13431 1891 13441 2045
rect 13481 1891 13491 2045
rect 13549 1891 13559 2045
rect 13599 1891 13609 2045
rect 13667 1891 13677 2045
rect 13717 1891 13727 2045
rect 13785 1891 13795 2045
rect 13835 1891 13845 2045
rect 13903 1891 13913 2045
rect 13953 1891 13963 2045
rect 14021 1891 14031 2045
rect 14071 1891 14081 2045
rect 14139 1891 14149 2045
rect 14189 1891 14199 2045
rect 14257 1891 14267 2045
rect 14307 1891 14317 2045
rect 14375 1891 14385 2045
rect 14425 1891 14435 2045
rect 14493 1891 14503 2045
rect 14543 1891 14553 2045
rect 14611 1891 14621 2045
rect 14661 1891 14671 2045
rect 14729 1891 14739 2045
rect 14779 1891 14789 2045
rect 14847 1891 14857 2045
rect 14897 1891 14907 2045
rect 14965 1891 14975 2045
rect 15015 1891 15025 2045
rect 15083 1891 15093 2045
rect 15133 1891 15143 2045
rect 15201 1891 15211 2045
rect 15251 1891 15261 2045
rect 15319 1891 15329 2045
rect 15369 1891 15379 2045
rect 15437 1891 15447 2045
rect 15487 1891 15497 2045
rect 15555 1891 15565 2045
rect 15605 1891 15615 2045
rect 15673 1891 15683 2045
rect 15723 1891 15733 2045
rect 15791 1891 15801 2045
rect 15841 1891 15851 2045
rect 15909 1891 15919 2045
rect 15959 1891 15969 2045
rect 16027 1891 16037 2045
rect 16077 1891 16087 2045
rect 16145 1891 16155 2045
rect 16195 1891 16205 2045
rect 16263 1891 16273 2045
rect 16313 1891 16323 2045
rect 16381 1891 16391 2045
rect 16431 1891 16441 2045
rect 16499 1891 16509 2045
rect 16549 1891 16559 2045
rect 16617 1891 16627 2045
rect 16667 1891 16677 2045
rect 16735 1891 16745 2045
rect 16785 1891 16795 2045
rect 16853 1891 16863 2045
rect 16903 1891 16913 2045
rect 16971 1891 16981 2045
rect 17021 1891 17031 2045
rect 17089 1891 17099 2045
rect 17139 1891 17149 2045
rect 17207 1891 17217 2045
rect 17257 1891 17267 2045
rect 17325 1891 17335 2045
rect 17375 1891 17385 2045
rect 17443 1891 17453 2045
rect 17493 1891 17503 2045
rect 17561 1891 17571 2045
rect 17611 1891 17621 2045
rect 17679 1891 17689 2045
rect 17729 1891 17739 2045
rect 17797 1891 17807 2045
rect 17847 1891 17857 2045
rect 17915 1891 17925 2045
rect 17965 1891 17975 2045
rect 18033 1891 18043 2045
rect 18083 1891 18093 2045
rect 18151 1891 18161 2045
rect 18201 1891 18211 2045
rect 18269 1891 18279 2045
rect 18319 1891 18329 2045
rect 18387 1891 18397 2045
rect 18437 1891 18447 2045
rect 18505 1891 18515 2045
rect 18555 1891 18565 2045
rect 18623 1891 18633 2045
rect 18673 1891 18683 2045
rect 18741 1891 18751 2045
rect 18791 1891 18801 2045
rect 18859 1891 18869 2045
rect 18909 1891 18919 2045
rect 18977 1891 18987 2045
rect 19027 1891 19037 2045
rect 19095 1891 19105 2045
rect 19145 1891 19155 2045
rect 19213 1891 19223 2045
rect 19263 1891 19273 2045
rect 19331 1891 19341 2045
rect 19381 1891 19391 2045
rect 19449 1891 19459 2045
rect 19499 1891 19509 2045
rect 19567 1891 19577 2045
rect 19617 1891 19627 2045
rect 19685 1891 19695 2045
rect 19735 1891 19745 2045
rect 19803 1891 19813 2045
rect 19853 1891 19863 2045
rect 19921 1891 19931 2045
rect 19971 1891 19981 2045
rect 20039 1891 20049 2045
rect 20089 1891 20099 2045
rect 20157 1891 20167 2045
rect 20207 1891 20217 2045
rect 20275 1891 20285 2045
rect 20325 1891 20335 2045
rect 20393 1891 20403 2045
rect 20443 1891 20453 2045
rect 20511 1891 20521 2045
rect 20561 1891 20571 2045
rect 20629 1891 20639 2045
rect 20679 1891 20689 2045
rect 20747 1891 20757 2045
rect 20797 1891 20807 2045
rect 20865 1891 20875 2045
rect 20915 1891 20925 2045
rect 20983 1891 20993 2045
rect 21033 1891 21043 2045
rect 21101 1891 21111 2045
rect 21151 1891 21161 2045
rect 21219 1891 21229 2045
rect 21269 1891 21279 2045
rect 21337 1891 21347 2045
rect 1327 -296 1337 -142
rect 1395 -296 1405 -142
rect 1445 -296 1455 -142
rect 1513 -296 1523 -142
rect 1563 -296 1573 -142
rect 1631 -296 1641 -142
rect 1681 -296 1691 -142
rect 1749 -296 1759 -142
rect 1799 -296 1809 -142
rect 1867 -296 1877 -142
rect 1917 -296 1927 -142
rect 1985 -296 1995 -142
rect 2035 -296 2045 -142
rect 2103 -296 2113 -142
rect 2153 -296 2163 -142
rect 2221 -296 2231 -142
rect 2271 -296 2281 -142
rect 2339 -296 2349 -142
rect 2389 -296 2399 -142
rect 2457 -296 2467 -142
rect 2507 -296 2517 -142
rect 2575 -296 2585 -142
rect 2625 -296 2635 -142
rect 2693 -296 2703 -142
rect 2743 -296 2753 -142
rect 2811 -296 2821 -142
rect 2861 -296 2871 -142
rect 2929 -296 2939 -142
rect 2979 -296 2989 -142
rect 3047 -296 3057 -142
rect 3097 -296 3107 -142
rect 3165 -296 3175 -142
rect 3215 -296 3225 -142
rect 3283 -296 3293 -142
rect 3333 -296 3343 -142
rect 3401 -296 3411 -142
rect 3451 -296 3461 -142
rect 3519 -296 3529 -142
rect 3569 -296 3579 -142
rect 3637 -296 3647 -142
rect 3687 -296 3697 -142
rect 3755 -296 3765 -142
rect 3805 -296 3815 -142
rect 3873 -296 3883 -142
rect 3923 -296 3933 -142
rect 3991 -296 4001 -142
rect 4041 -296 4051 -142
rect 4109 -296 4119 -142
rect 4159 -296 4169 -142
rect 4227 -296 4237 -142
rect 4277 -296 4287 -142
rect 4345 -296 4355 -142
rect 4395 -296 4405 -142
rect 4463 -296 4473 -142
rect 4513 -296 4523 -142
rect 4581 -296 4591 -142
rect 4631 -296 4641 -142
rect 4699 -296 4709 -142
rect 4749 -296 4759 -142
rect 4817 -296 4827 -142
rect 4867 -296 4877 -142
rect 4935 -296 4945 -142
rect 4985 -296 4995 -142
rect 5053 -296 5063 -142
rect 5103 -296 5113 -142
rect 5171 -296 5181 -142
rect 5221 -296 5231 -142
rect 5289 -296 5299 -142
rect 5339 -296 5349 -142
rect 5407 -296 5417 -142
rect 5457 -296 5467 -142
rect 5525 -296 5535 -142
rect 5575 -296 5585 -142
rect 5643 -296 5653 -142
rect 5693 -296 5703 -142
rect 5761 -296 5771 -142
rect 5811 -296 5821 -142
rect 5879 -296 5889 -142
rect 5929 -296 5939 -142
rect 5997 -296 6007 -142
rect 6047 -296 6057 -142
rect 6115 -296 6125 -142
rect 6165 -296 6175 -142
rect 6233 -296 6243 -142
rect 6283 -296 6293 -142
rect 6351 -296 6361 -142
rect 6401 -296 6411 -142
rect 6469 -296 6479 -142
rect 6519 -296 6529 -142
rect 6587 -296 6597 -142
rect 6637 -296 6647 -142
rect 6705 -296 6715 -142
rect 6755 -296 6765 -142
rect 6823 -296 6833 -142
rect 6873 -296 6883 -142
rect 6941 -296 6951 -142
rect 6991 -296 7001 -142
rect 7059 -296 7069 -142
rect 7109 -296 7119 -142
rect 7177 -296 7187 -142
rect 1327 -2064 1337 -1910
rect 1395 -2064 1405 -1910
rect 1445 -2064 1455 -1910
rect 1513 -2064 1523 -1910
rect 1563 -2064 1573 -1910
rect 1631 -2064 1641 -1910
rect 1681 -2064 1691 -1910
rect 1749 -2064 1759 -1910
rect 1799 -2064 1809 -1910
rect 1867 -2064 1877 -1910
rect 1917 -2064 1927 -1910
rect 1985 -2064 1995 -1910
rect 2035 -2064 2045 -1910
rect 2103 -2064 2113 -1910
rect 2153 -2064 2163 -1910
rect 2221 -2064 2231 -1910
rect 2271 -2064 2281 -1910
rect 2339 -2064 2349 -1910
rect 2389 -2064 2399 -1910
rect 2457 -2064 2467 -1910
rect 2507 -2064 2517 -1910
rect 2575 -2064 2585 -1910
rect 2625 -2064 2635 -1910
rect 2693 -2064 2703 -1910
rect 2743 -2064 2753 -1910
rect 2811 -2064 2821 -1910
rect 2861 -2064 2871 -1910
rect 2929 -2064 2939 -1910
rect 2979 -2064 2989 -1910
rect 3047 -2064 3057 -1910
rect 3097 -2064 3107 -1910
rect 3165 -2064 3175 -1910
rect 3215 -2064 3225 -1910
rect 3283 -2064 3293 -1910
rect 3333 -2064 3343 -1910
rect 3401 -2064 3411 -1910
rect 3451 -2064 3461 -1910
rect 3519 -2064 3529 -1910
rect 3569 -2064 3579 -1910
rect 3637 -2064 3647 -1910
rect 3687 -2064 3697 -1910
rect 3755 -2064 3765 -1910
rect 3805 -2064 3815 -1910
rect 3873 -2064 3883 -1910
rect 3923 -2064 3933 -1910
rect 3991 -2064 4001 -1910
rect 4041 -2064 4051 -1910
rect 4109 -2064 4119 -1910
rect 4159 -2064 4169 -1910
rect 4227 -2064 4237 -1910
rect 4277 -2064 4287 -1910
rect 4345 -2064 4355 -1910
rect 4395 -2064 4405 -1910
rect 4463 -2064 4473 -1910
rect 4513 -2064 4523 -1910
rect 4581 -2064 4591 -1910
rect 4631 -2064 4641 -1910
rect 4699 -2064 4709 -1910
rect 4749 -2064 4759 -1910
rect 4817 -2064 4827 -1910
rect 4867 -2064 4877 -1910
rect 4935 -2064 4945 -1910
rect 4985 -2064 4995 -1910
rect 5053 -2064 5063 -1910
rect 5103 -2064 5113 -1910
rect 5171 -2064 5181 -1910
rect 5221 -2064 5231 -1910
rect 5289 -2064 5299 -1910
rect 5339 -2064 5349 -1910
rect 5407 -2064 5417 -1910
rect 5457 -2064 5467 -1910
rect 5525 -2064 5535 -1910
rect 5575 -2064 5585 -1910
rect 5643 -2064 5653 -1910
rect 5693 -2064 5703 -1910
rect 5761 -2064 5771 -1910
rect 5811 -2064 5821 -1910
rect 5879 -2064 5889 -1910
rect 5929 -2064 5939 -1910
rect 5997 -2064 6007 -1910
rect 6047 -2064 6057 -1910
rect 6115 -2064 6125 -1910
rect 6165 -2064 6175 -1910
rect 6233 -2064 6243 -1910
rect 6283 -2064 6293 -1910
rect 6351 -2064 6361 -1910
rect 6401 -2064 6411 -1910
rect 6469 -2064 6479 -1910
rect 6519 -2064 6529 -1910
rect 6587 -2064 6597 -1910
rect 6637 -2064 6647 -1910
rect 6705 -2064 6715 -1910
rect 6755 -2064 6765 -1910
rect 6823 -2064 6833 -1910
rect 6873 -2064 6883 -1910
rect 6941 -2064 6951 -1910
rect 6991 -2064 7001 -1910
rect 7059 -2064 7069 -1910
rect 7109 -2064 7119 -1910
rect 7177 -2064 7187 -1910
rect 1327 -3832 1337 -3678
rect 1395 -3832 1405 -3678
rect 1445 -3832 1455 -3678
rect 1513 -3832 1523 -3678
rect 1563 -3832 1573 -3678
rect 1631 -3832 1641 -3678
rect 1681 -3832 1691 -3678
rect 1749 -3832 1759 -3678
rect 1799 -3832 1809 -3678
rect 1867 -3832 1877 -3678
rect 1917 -3832 1927 -3678
rect 1985 -3832 1995 -3678
rect 2035 -3832 2045 -3678
rect 2103 -3832 2113 -3678
rect 2153 -3832 2163 -3678
rect 2221 -3832 2231 -3678
rect 2271 -3832 2281 -3678
rect 2339 -3832 2349 -3678
rect 2389 -3832 2399 -3678
rect 2457 -3832 2467 -3678
rect 2507 -3832 2517 -3678
rect 2575 -3832 2585 -3678
rect 2625 -3832 2635 -3678
rect 2693 -3832 2703 -3678
rect 2743 -3832 2753 -3678
rect 2811 -3832 2821 -3678
rect 2861 -3832 2871 -3678
rect 2929 -3832 2939 -3678
rect 2979 -3832 2989 -3678
rect 3047 -3832 3057 -3678
rect 3097 -3832 3107 -3678
rect 3165 -3832 3175 -3678
rect 3215 -3832 3225 -3678
rect 3283 -3832 3293 -3678
rect 3333 -3832 3343 -3678
rect 3401 -3832 3411 -3678
rect 3451 -3832 3461 -3678
rect 3519 -3832 3529 -3678
rect 3569 -3832 3579 -3678
rect 3637 -3832 3647 -3678
rect 3687 -3832 3697 -3678
rect 3755 -3832 3765 -3678
rect 3805 -3832 3815 -3678
rect 3873 -3832 3883 -3678
rect 3923 -3832 3933 -3678
rect 3991 -3832 4001 -3678
rect 4041 -3832 4051 -3678
rect 4109 -3832 4119 -3678
rect 4159 -3832 4169 -3678
rect 4227 -3832 4237 -3678
rect 4277 -3832 4287 -3678
rect 4345 -3832 4355 -3678
rect 4395 -3832 4405 -3678
rect 4463 -3832 4473 -3678
rect 4513 -3832 4523 -3678
rect 4581 -3832 4591 -3678
rect 4631 -3832 4641 -3678
rect 4699 -3832 4709 -3678
rect 4749 -3832 4759 -3678
rect 4817 -3832 4827 -3678
rect 4867 -3832 4877 -3678
rect 4935 -3832 4945 -3678
rect 4985 -3832 4995 -3678
rect 5053 -3832 5063 -3678
rect 5103 -3832 5113 -3678
rect 5171 -3832 5181 -3678
rect 5221 -3832 5231 -3678
rect 5289 -3832 5299 -3678
rect 5339 -3832 5349 -3678
rect 5407 -3832 5417 -3678
rect 5457 -3832 5467 -3678
rect 5525 -3832 5535 -3678
rect 5575 -3832 5585 -3678
rect 5643 -3832 5653 -3678
rect 5693 -3832 5703 -3678
rect 5761 -3832 5771 -3678
rect 5811 -3832 5821 -3678
rect 5879 -3832 5889 -3678
rect 5929 -3832 5939 -3678
rect 5997 -3832 6007 -3678
rect 6047 -3832 6057 -3678
rect 6115 -3832 6125 -3678
rect 6165 -3832 6175 -3678
rect 6233 -3832 6243 -3678
rect 6283 -3832 6293 -3678
rect 6351 -3832 6361 -3678
rect 6401 -3832 6411 -3678
rect 6469 -3832 6479 -3678
rect 6519 -3832 6529 -3678
rect 6587 -3832 6597 -3678
rect 6637 -3832 6647 -3678
rect 6705 -3832 6715 -3678
rect 6755 -3832 6765 -3678
rect 6823 -3832 6833 -3678
rect 6873 -3832 6883 -3678
rect 6941 -3832 6951 -3678
rect 6991 -3832 7001 -3678
rect 7059 -3832 7069 -3678
rect 7109 -3832 7119 -3678
rect 7177 -3832 7187 -3678
rect 1327 -5600 1337 -5446
rect 1395 -5600 1405 -5446
rect 1445 -5600 1455 -5446
rect 1513 -5600 1523 -5446
rect 1563 -5600 1573 -5446
rect 1631 -5600 1641 -5446
rect 1681 -5600 1691 -5446
rect 1749 -5600 1759 -5446
rect 1799 -5600 1809 -5446
rect 1867 -5600 1877 -5446
rect 1917 -5600 1927 -5446
rect 1985 -5600 1995 -5446
rect 2035 -5600 2045 -5446
rect 2103 -5600 2113 -5446
rect 2153 -5600 2163 -5446
rect 2221 -5600 2231 -5446
rect 2271 -5600 2281 -5446
rect 2339 -5600 2349 -5446
rect 2389 -5600 2399 -5446
rect 2457 -5600 2467 -5446
rect 2507 -5600 2517 -5446
rect 2575 -5600 2585 -5446
rect 2625 -5600 2635 -5446
rect 2693 -5600 2703 -5446
rect 2743 -5600 2753 -5446
rect 2811 -5600 2821 -5446
rect 2861 -5600 2871 -5446
rect 2929 -5600 2939 -5446
rect 2979 -5600 2989 -5446
rect 3047 -5600 3057 -5446
rect 3097 -5600 3107 -5446
rect 3165 -5600 3175 -5446
rect 3215 -5600 3225 -5446
rect 3283 -5600 3293 -5446
rect 3333 -5600 3343 -5446
rect 3401 -5600 3411 -5446
rect 3451 -5600 3461 -5446
rect 3519 -5600 3529 -5446
rect 3569 -5600 3579 -5446
rect 3637 -5600 3647 -5446
rect 3687 -5600 3697 -5446
rect 3755 -5600 3765 -5446
rect 3805 -5600 3815 -5446
rect 3873 -5600 3883 -5446
rect 3923 -5600 3933 -5446
rect 3991 -5600 4001 -5446
rect 4041 -5600 4051 -5446
rect 4109 -5600 4119 -5446
rect 4159 -5600 4169 -5446
rect 4227 -5600 4237 -5446
rect 4277 -5600 4287 -5446
rect 4345 -5600 4355 -5446
rect 4395 -5600 4405 -5446
rect 4463 -5600 4473 -5446
rect 4513 -5600 4523 -5446
rect 4581 -5600 4591 -5446
rect 4631 -5600 4641 -5446
rect 4699 -5600 4709 -5446
rect 4749 -5600 4759 -5446
rect 4817 -5600 4827 -5446
rect 4867 -5600 4877 -5446
rect 4935 -5600 4945 -5446
rect 4985 -5600 4995 -5446
rect 5053 -5600 5063 -5446
rect 5103 -5600 5113 -5446
rect 5171 -5600 5181 -5446
rect 5221 -5600 5231 -5446
rect 5289 -5600 5299 -5446
rect 5339 -5600 5349 -5446
rect 5407 -5600 5417 -5446
rect 5457 -5600 5467 -5446
rect 5525 -5600 5535 -5446
rect 5575 -5600 5585 -5446
rect 5643 -5600 5653 -5446
rect 5693 -5600 5703 -5446
rect 5761 -5600 5771 -5446
rect 5811 -5600 5821 -5446
rect 5879 -5600 5889 -5446
rect 5929 -5600 5939 -5446
rect 5997 -5600 6007 -5446
rect 6047 -5600 6057 -5446
rect 6115 -5600 6125 -5446
rect 6165 -5600 6175 -5446
rect 6233 -5600 6243 -5446
rect 6283 -5600 6293 -5446
rect 6351 -5600 6361 -5446
rect 6401 -5600 6411 -5446
rect 6469 -5600 6479 -5446
rect 6519 -5600 6529 -5446
rect 6587 -5600 6597 -5446
rect 6637 -5600 6647 -5446
rect 6705 -5600 6715 -5446
rect 6755 -5600 6765 -5446
rect 6823 -5600 6833 -5446
rect 6873 -5600 6883 -5446
rect 6941 -5600 6951 -5446
rect 6991 -5600 7001 -5446
rect 7059 -5600 7069 -5446
rect 7109 -5600 7119 -5446
rect 7177 -5600 7187 -5446
rect 11457 -6642 11503 -6630
rect 11457 -6646 11463 -6642
rect 11497 -6646 11503 -6642
rect 11605 -6642 11651 -6630
rect 11605 -6646 11611 -6642
rect 11645 -6646 11651 -6642
rect 11753 -6642 11799 -6630
rect 11753 -6646 11759 -6642
rect 11793 -6646 11799 -6642
rect 11901 -6642 11947 -6630
rect 11901 -6646 11907 -6642
rect 11941 -6646 11947 -6642
rect 12049 -6642 12095 -6630
rect 12049 -6646 12055 -6642
rect 12089 -6646 12095 -6642
rect 12197 -6642 12243 -6630
rect 12197 -6646 12203 -6642
rect 12237 -6646 12243 -6642
rect 12345 -6642 12391 -6630
rect 12345 -6646 12351 -6642
rect 12385 -6646 12391 -6642
rect 12493 -6642 12539 -6630
rect 12493 -6646 12499 -6642
rect 12533 -6646 12539 -6642
rect 12641 -6642 12687 -6630
rect 12641 -6646 12647 -6642
rect 12681 -6646 12687 -6642
rect 12789 -6642 12835 -6630
rect 12789 -6646 12795 -6642
rect 12829 -6646 12835 -6642
rect 12937 -6642 12983 -6630
rect 12937 -6646 12943 -6642
rect 12977 -6646 12983 -6642
rect 13085 -6642 13131 -6630
rect 13085 -6646 13091 -6642
rect 13125 -6646 13131 -6642
rect 13233 -6642 13279 -6630
rect 13233 -6646 13239 -6642
rect 13273 -6646 13279 -6642
rect 13381 -6642 13427 -6630
rect 13381 -6646 13387 -6642
rect 13421 -6646 13427 -6642
rect 13529 -6642 13575 -6630
rect 13529 -6646 13535 -6642
rect 13569 -6646 13575 -6642
rect 13677 -6642 13723 -6630
rect 13677 -6646 13683 -6642
rect 13717 -6646 13723 -6642
rect 13825 -6642 13871 -6630
rect 13825 -6646 13831 -6642
rect 13865 -6646 13871 -6642
rect 13973 -6642 14019 -6630
rect 13973 -6646 13979 -6642
rect 14013 -6646 14019 -6642
rect 14121 -6642 14167 -6630
rect 14121 -6646 14127 -6642
rect 14161 -6646 14167 -6642
rect 14269 -6642 14315 -6630
rect 14269 -6646 14275 -6642
rect 14309 -6646 14315 -6642
rect 14417 -6642 14463 -6630
rect 14417 -6646 14423 -6642
rect 14457 -6646 14463 -6642
rect 14565 -6642 14611 -6630
rect 14565 -6646 14571 -6642
rect 14605 -6646 14611 -6642
rect 14713 -6642 14759 -6630
rect 14713 -6646 14719 -6642
rect 14753 -6646 14759 -6642
rect 14861 -6642 14907 -6630
rect 14861 -6646 14867 -6642
rect 14901 -6646 14907 -6642
rect 15009 -6642 15055 -6630
rect 15009 -6646 15015 -6642
rect 15049 -6646 15055 -6642
rect 15157 -6642 15203 -6630
rect 15157 -6646 15163 -6642
rect 15197 -6646 15203 -6642
rect 15305 -6642 15351 -6630
rect 15305 -6646 15311 -6642
rect 15345 -6646 15351 -6642
rect 15453 -6642 15499 -6630
rect 15453 -6646 15459 -6642
rect 15493 -6646 15499 -6642
rect 15601 -6642 15647 -6630
rect 15601 -6646 15607 -6642
rect 15641 -6646 15647 -6642
rect 15749 -6642 15795 -6630
rect 15749 -6646 15755 -6642
rect 15789 -6646 15795 -6642
rect 15897 -6642 15943 -6630
rect 15897 -6646 15903 -6642
rect 15937 -6646 15943 -6642
rect 16045 -6642 16091 -6630
rect 16045 -6646 16051 -6642
rect 16085 -6646 16091 -6642
rect 16193 -6642 16239 -6630
rect 16193 -6646 16199 -6642
rect 16233 -6646 16239 -6642
rect 16341 -6642 16387 -6630
rect 16341 -6646 16347 -6642
rect 16381 -6646 16387 -6642
rect 16489 -6642 16535 -6630
rect 16489 -6646 16495 -6642
rect 16529 -6646 16535 -6642
rect 16637 -6642 16683 -6630
rect 16637 -6646 16643 -6642
rect 16677 -6646 16683 -6642
rect 16785 -6642 16831 -6630
rect 16785 -6646 16791 -6642
rect 16825 -6646 16831 -6642
rect 16933 -6642 16979 -6630
rect 16933 -6646 16939 -6642
rect 16973 -6646 16979 -6642
rect 17081 -6642 17127 -6630
rect 17081 -6646 17087 -6642
rect 17121 -6646 17127 -6642
rect 17229 -6642 17275 -6630
rect 17229 -6646 17235 -6642
rect 17269 -6646 17275 -6642
rect 17377 -6642 17423 -6630
rect 17377 -6646 17383 -6642
rect 17417 -6646 17423 -6642
rect 17525 -6642 17571 -6630
rect 17525 -6646 17531 -6642
rect 17565 -6646 17571 -6642
rect 17673 -6642 17719 -6630
rect 17673 -6646 17679 -6642
rect 17713 -6646 17719 -6642
rect 17821 -6642 17867 -6630
rect 17821 -6646 17827 -6642
rect 17861 -6646 17867 -6642
rect 17969 -6642 18015 -6630
rect 17969 -6646 17975 -6642
rect 18009 -6646 18015 -6642
rect 18117 -6642 18163 -6630
rect 18117 -6646 18123 -6642
rect 18157 -6646 18163 -6642
rect 18265 -6642 18311 -6630
rect 18265 -6646 18271 -6642
rect 18305 -6646 18311 -6642
rect 18413 -6642 18459 -6630
rect 18413 -6646 18419 -6642
rect 18453 -6646 18459 -6642
rect 18561 -6642 18607 -6630
rect 18561 -6646 18567 -6642
rect 18601 -6646 18607 -6642
rect 18709 -6642 18755 -6630
rect 18709 -6646 18715 -6642
rect 18749 -6646 18755 -6642
rect 18857 -6642 18903 -6630
rect 18857 -6646 18863 -6642
rect 18897 -6646 18903 -6642
rect 19005 -6642 19051 -6630
rect 19005 -6646 19011 -6642
rect 19045 -6646 19051 -6642
rect 19153 -6642 19199 -6630
rect 19153 -6646 19159 -6642
rect 19193 -6646 19199 -6642
rect 19301 -6642 19347 -6630
rect 19301 -6646 19307 -6642
rect 19341 -6646 19347 -6642
rect 19449 -6642 19495 -6630
rect 19449 -6646 19455 -6642
rect 19489 -6646 19495 -6642
rect 19597 -6642 19643 -6630
rect 19597 -6646 19603 -6642
rect 19637 -6646 19643 -6642
rect 19745 -6642 19791 -6630
rect 19745 -6646 19751 -6642
rect 19785 -6646 19791 -6642
rect 19893 -6642 19939 -6630
rect 19893 -6646 19899 -6642
rect 19933 -6646 19939 -6642
rect 20041 -6642 20087 -6630
rect 20041 -6646 20047 -6642
rect 20081 -6646 20087 -6642
rect 20189 -6642 20235 -6630
rect 20189 -6646 20195 -6642
rect 20229 -6646 20235 -6642
rect 20337 -6642 20383 -6630
rect 20337 -6646 20343 -6642
rect 20377 -6646 20383 -6642
rect 20485 -6642 20531 -6630
rect 20485 -6646 20491 -6642
rect 20525 -6646 20531 -6642
rect 20633 -6642 20679 -6630
rect 20633 -6646 20639 -6642
rect 20673 -6646 20679 -6642
rect 20781 -6642 20827 -6630
rect 20781 -6646 20787 -6642
rect 20821 -6646 20827 -6642
rect 20929 -6642 20975 -6630
rect 20929 -6646 20935 -6642
rect 20969 -6646 20975 -6642
rect 21077 -6642 21123 -6630
rect 21077 -6646 21083 -6642
rect 21117 -6646 21123 -6642
rect 21225 -6642 21271 -6630
rect 21225 -6646 21231 -6642
rect 21265 -6646 21271 -6642
rect 21373 -6642 21419 -6630
rect 21373 -6646 21379 -6642
rect 21413 -6646 21419 -6642
rect 21521 -6642 21567 -6630
rect 21521 -6646 21527 -6642
rect 21561 -6646 21567 -6642
rect 21669 -6642 21715 -6630
rect 21669 -6646 21675 -6642
rect 21709 -6646 21715 -6642
rect 21817 -6642 21863 -6630
rect 21817 -6646 21823 -6642
rect 21857 -6646 21863 -6642
rect 21965 -6642 22011 -6630
rect 21965 -6646 21971 -6642
rect 22005 -6646 22011 -6642
rect 22113 -6642 22159 -6630
rect 22113 -6646 22119 -6642
rect 22153 -6646 22159 -6642
rect 22261 -6642 22307 -6630
rect 22261 -6646 22267 -6642
rect 22301 -6646 22307 -6642
rect 22557 -6642 22603 -6630
rect 22557 -6646 22563 -6642
rect 22597 -6646 22603 -6642
rect 11444 -7486 11454 -6646
rect 11506 -7486 11516 -6646
rect 11592 -7486 11602 -6646
rect 11654 -7486 11664 -6646
rect 11740 -7486 11750 -6646
rect 11802 -7486 11812 -6646
rect 11888 -7486 11898 -6646
rect 11950 -7486 11960 -6646
rect 12036 -7486 12046 -6646
rect 12098 -7486 12108 -6646
rect 12184 -7486 12194 -6646
rect 12246 -7486 12256 -6646
rect 12332 -7486 12342 -6646
rect 12394 -7486 12404 -6646
rect 12480 -7486 12490 -6646
rect 12542 -7486 12552 -6646
rect 12628 -7486 12638 -6646
rect 12690 -7486 12700 -6646
rect 12776 -7486 12786 -6646
rect 12838 -7486 12848 -6646
rect 12924 -7486 12934 -6646
rect 12986 -7486 12996 -6646
rect 13072 -7486 13082 -6646
rect 13134 -7486 13144 -6646
rect 13220 -7486 13230 -6646
rect 13282 -7486 13292 -6646
rect 13368 -7486 13378 -6646
rect 13430 -7486 13440 -6646
rect 13516 -7486 13526 -6646
rect 13578 -7486 13588 -6646
rect 13664 -7486 13674 -6646
rect 13726 -7486 13736 -6646
rect 13812 -7486 13822 -6646
rect 13874 -7486 13884 -6646
rect 13960 -7486 13970 -6646
rect 14022 -7486 14032 -6646
rect 14108 -7486 14118 -6646
rect 14170 -7486 14180 -6646
rect 14256 -7486 14266 -6646
rect 14318 -7486 14328 -6646
rect 14404 -7486 14414 -6646
rect 14466 -7486 14476 -6646
rect 14552 -7486 14562 -6646
rect 14614 -7486 14624 -6646
rect 14700 -7486 14710 -6646
rect 14762 -7486 14772 -6646
rect 14848 -7486 14858 -6646
rect 14910 -7486 14920 -6646
rect 14996 -7486 15006 -6646
rect 15058 -7486 15068 -6646
rect 15144 -7486 15154 -6646
rect 15206 -7486 15216 -6646
rect 15292 -7486 15302 -6646
rect 15354 -7486 15364 -6646
rect 15440 -7486 15450 -6646
rect 15502 -7486 15512 -6646
rect 15588 -7486 15598 -6646
rect 15650 -7486 15660 -6646
rect 15736 -7486 15746 -6646
rect 15798 -7486 15808 -6646
rect 15884 -7486 15894 -6646
rect 15946 -7486 15956 -6646
rect 16032 -7486 16042 -6646
rect 16094 -7486 16104 -6646
rect 16180 -7486 16190 -6646
rect 16242 -7486 16252 -6646
rect 16328 -7486 16338 -6646
rect 16390 -7486 16400 -6646
rect 16476 -7486 16486 -6646
rect 16538 -7486 16548 -6646
rect 16624 -7486 16634 -6646
rect 16686 -7486 16696 -6646
rect 16772 -7486 16782 -6646
rect 16834 -7486 16844 -6646
rect 16920 -7486 16930 -6646
rect 16982 -7486 16992 -6646
rect 17068 -7486 17078 -6646
rect 17130 -7486 17140 -6646
rect 17216 -7486 17226 -6646
rect 17278 -7486 17288 -6646
rect 17364 -7486 17374 -6646
rect 17426 -7486 17436 -6646
rect 17512 -7486 17522 -6646
rect 17574 -7486 17584 -6646
rect 17660 -7486 17670 -6646
rect 17722 -7486 17732 -6646
rect 17808 -7486 17818 -6646
rect 17870 -7486 17880 -6646
rect 17956 -7486 17966 -6646
rect 18018 -7486 18028 -6646
rect 18104 -7486 18114 -6646
rect 18166 -7486 18176 -6646
rect 18252 -7486 18262 -6646
rect 18314 -7486 18324 -6646
rect 18400 -7486 18410 -6646
rect 18462 -7486 18472 -6646
rect 18548 -7486 18558 -6646
rect 18610 -7486 18620 -6646
rect 18696 -7486 18706 -6646
rect 18758 -7486 18768 -6646
rect 18844 -7486 18854 -6646
rect 18906 -7486 18916 -6646
rect 18992 -7486 19002 -6646
rect 19054 -7486 19064 -6646
rect 19140 -7486 19150 -6646
rect 19202 -7486 19212 -6646
rect 19288 -7486 19298 -6646
rect 19350 -7486 19360 -6646
rect 19436 -7486 19446 -6646
rect 19498 -7486 19508 -6646
rect 19584 -7486 19594 -6646
rect 19646 -7486 19656 -6646
rect 19732 -7486 19742 -6646
rect 19794 -7486 19804 -6646
rect 19880 -7486 19890 -6646
rect 19942 -7486 19952 -6646
rect 20028 -7486 20038 -6646
rect 20090 -7486 20100 -6646
rect 20176 -7486 20186 -6646
rect 20238 -7486 20248 -6646
rect 20324 -7486 20334 -6646
rect 20386 -7486 20396 -6646
rect 20472 -7486 20482 -6646
rect 20534 -7486 20544 -6646
rect 20620 -7486 20630 -6646
rect 20682 -7486 20692 -6646
rect 20768 -7486 20778 -6646
rect 20830 -7486 20840 -6646
rect 20916 -7486 20926 -6646
rect 20978 -7486 20988 -6646
rect 21064 -7486 21074 -6646
rect 21126 -7486 21136 -6646
rect 21212 -7486 21222 -6646
rect 21274 -7486 21284 -6646
rect 21360 -7486 21370 -6646
rect 21422 -7486 21432 -6646
rect 21508 -7486 21518 -6646
rect 21570 -7486 21580 -6646
rect 21656 -7486 21666 -6646
rect 21718 -7486 21728 -6646
rect 21804 -7486 21814 -6646
rect 21866 -7486 21876 -6646
rect 21952 -7486 21962 -6646
rect 22014 -7486 22024 -6646
rect 22100 -7486 22110 -6646
rect 22162 -7486 22172 -6646
rect 22248 -7486 22258 -6646
rect 22310 -7486 22320 -6646
rect 22396 -7486 22406 -6646
rect 22458 -7486 22468 -6646
rect 22544 -7486 22554 -6646
rect 22606 -7486 22616 -6646
rect 11457 -7518 11463 -7486
rect 11497 -7518 11503 -7486
rect 11457 -7530 11503 -7518
rect 11605 -7518 11611 -7486
rect 11645 -7518 11651 -7486
rect 11605 -7530 11651 -7518
rect 11753 -7518 11759 -7486
rect 11793 -7518 11799 -7486
rect 11753 -7530 11799 -7518
rect 11901 -7518 11907 -7486
rect 11941 -7518 11947 -7486
rect 11901 -7530 11947 -7518
rect 12049 -7518 12055 -7486
rect 12089 -7518 12095 -7486
rect 12049 -7530 12095 -7518
rect 12197 -7518 12203 -7486
rect 12237 -7518 12243 -7486
rect 12197 -7530 12243 -7518
rect 12345 -7518 12351 -7486
rect 12385 -7518 12391 -7486
rect 12345 -7530 12391 -7518
rect 12493 -7518 12499 -7486
rect 12533 -7518 12539 -7486
rect 12493 -7530 12539 -7518
rect 12641 -7518 12647 -7486
rect 12681 -7518 12687 -7486
rect 12641 -7530 12687 -7518
rect 12789 -7518 12795 -7486
rect 12829 -7518 12835 -7486
rect 12789 -7530 12835 -7518
rect 12937 -7518 12943 -7486
rect 12977 -7518 12983 -7486
rect 12937 -7530 12983 -7518
rect 13085 -7518 13091 -7486
rect 13125 -7518 13131 -7486
rect 13085 -7530 13131 -7518
rect 13233 -7518 13239 -7486
rect 13273 -7518 13279 -7486
rect 13233 -7530 13279 -7518
rect 13381 -7518 13387 -7486
rect 13421 -7518 13427 -7486
rect 13381 -7530 13427 -7518
rect 13529 -7518 13535 -7486
rect 13569 -7518 13575 -7486
rect 13529 -7530 13575 -7518
rect 13677 -7518 13683 -7486
rect 13717 -7518 13723 -7486
rect 13677 -7530 13723 -7518
rect 13825 -7518 13831 -7486
rect 13865 -7518 13871 -7486
rect 13825 -7530 13871 -7518
rect 13973 -7518 13979 -7486
rect 14013 -7518 14019 -7486
rect 13973 -7530 14019 -7518
rect 14121 -7518 14127 -7486
rect 14161 -7518 14167 -7486
rect 14121 -7530 14167 -7518
rect 14269 -7518 14275 -7486
rect 14309 -7518 14315 -7486
rect 14269 -7530 14315 -7518
rect 14417 -7518 14423 -7486
rect 14457 -7518 14463 -7486
rect 14417 -7530 14463 -7518
rect 14565 -7518 14571 -7486
rect 14605 -7518 14611 -7486
rect 14565 -7530 14611 -7518
rect 14713 -7518 14719 -7486
rect 14753 -7518 14759 -7486
rect 14713 -7530 14759 -7518
rect 14861 -7518 14867 -7486
rect 14901 -7518 14907 -7486
rect 14861 -7530 14907 -7518
rect 15009 -7518 15015 -7486
rect 15049 -7518 15055 -7486
rect 15009 -7530 15055 -7518
rect 15157 -7518 15163 -7486
rect 15197 -7518 15203 -7486
rect 15157 -7530 15203 -7518
rect 15305 -7518 15311 -7486
rect 15345 -7518 15351 -7486
rect 15305 -7530 15351 -7518
rect 15453 -7518 15459 -7486
rect 15493 -7518 15499 -7486
rect 15453 -7530 15499 -7518
rect 15601 -7518 15607 -7486
rect 15641 -7518 15647 -7486
rect 15601 -7530 15647 -7518
rect 15749 -7518 15755 -7486
rect 15789 -7518 15795 -7486
rect 15749 -7530 15795 -7518
rect 15897 -7518 15903 -7486
rect 15937 -7518 15943 -7486
rect 15897 -7530 15943 -7518
rect 16045 -7518 16051 -7486
rect 16085 -7518 16091 -7486
rect 16045 -7530 16091 -7518
rect 16193 -7518 16199 -7486
rect 16233 -7518 16239 -7486
rect 16193 -7530 16239 -7518
rect 16341 -7518 16347 -7486
rect 16381 -7518 16387 -7486
rect 16341 -7530 16387 -7518
rect 16489 -7518 16495 -7486
rect 16529 -7518 16535 -7486
rect 16489 -7530 16535 -7518
rect 16637 -7518 16643 -7486
rect 16677 -7518 16683 -7486
rect 16637 -7530 16683 -7518
rect 16785 -7518 16791 -7486
rect 16825 -7518 16831 -7486
rect 16785 -7530 16831 -7518
rect 16933 -7518 16939 -7486
rect 16973 -7518 16979 -7486
rect 16933 -7530 16979 -7518
rect 17081 -7518 17087 -7486
rect 17121 -7518 17127 -7486
rect 17081 -7530 17127 -7518
rect 17229 -7518 17235 -7486
rect 17269 -7518 17275 -7486
rect 17229 -7530 17275 -7518
rect 17377 -7518 17383 -7486
rect 17417 -7518 17423 -7486
rect 17377 -7530 17423 -7518
rect 17525 -7518 17531 -7486
rect 17565 -7518 17571 -7486
rect 17525 -7530 17571 -7518
rect 17673 -7518 17679 -7486
rect 17713 -7518 17719 -7486
rect 17673 -7530 17719 -7518
rect 17821 -7518 17827 -7486
rect 17861 -7518 17867 -7486
rect 17821 -7530 17867 -7518
rect 17969 -7518 17975 -7486
rect 18009 -7518 18015 -7486
rect 17969 -7530 18015 -7518
rect 18117 -7518 18123 -7486
rect 18157 -7518 18163 -7486
rect 18117 -7530 18163 -7518
rect 18265 -7518 18271 -7486
rect 18305 -7518 18311 -7486
rect 18265 -7530 18311 -7518
rect 18413 -7518 18419 -7486
rect 18453 -7518 18459 -7486
rect 18413 -7530 18459 -7518
rect 18561 -7518 18567 -7486
rect 18601 -7518 18607 -7486
rect 18561 -7530 18607 -7518
rect 18709 -7518 18715 -7486
rect 18749 -7518 18755 -7486
rect 18709 -7530 18755 -7518
rect 18857 -7518 18863 -7486
rect 18897 -7518 18903 -7486
rect 18857 -7530 18903 -7518
rect 19005 -7518 19011 -7486
rect 19045 -7518 19051 -7486
rect 19005 -7530 19051 -7518
rect 19153 -7518 19159 -7486
rect 19193 -7518 19199 -7486
rect 19153 -7530 19199 -7518
rect 19301 -7518 19307 -7486
rect 19341 -7518 19347 -7486
rect 19301 -7530 19347 -7518
rect 19449 -7518 19455 -7486
rect 19489 -7518 19495 -7486
rect 19449 -7530 19495 -7518
rect 19597 -7518 19603 -7486
rect 19637 -7518 19643 -7486
rect 19597 -7530 19643 -7518
rect 19745 -7518 19751 -7486
rect 19785 -7518 19791 -7486
rect 19745 -7530 19791 -7518
rect 19893 -7518 19899 -7486
rect 19933 -7518 19939 -7486
rect 19893 -7530 19939 -7518
rect 20041 -7518 20047 -7486
rect 20081 -7518 20087 -7486
rect 20041 -7530 20087 -7518
rect 20189 -7518 20195 -7486
rect 20229 -7518 20235 -7486
rect 20189 -7530 20235 -7518
rect 20337 -7518 20343 -7486
rect 20377 -7518 20383 -7486
rect 20337 -7530 20383 -7518
rect 20485 -7518 20491 -7486
rect 20525 -7518 20531 -7486
rect 20485 -7530 20531 -7518
rect 20633 -7518 20639 -7486
rect 20673 -7518 20679 -7486
rect 20633 -7530 20679 -7518
rect 20781 -7518 20787 -7486
rect 20821 -7518 20827 -7486
rect 20781 -7530 20827 -7518
rect 20929 -7518 20935 -7486
rect 20969 -7518 20975 -7486
rect 20929 -7530 20975 -7518
rect 21077 -7518 21083 -7486
rect 21117 -7518 21123 -7486
rect 21077 -7530 21123 -7518
rect 21225 -7518 21231 -7486
rect 21265 -7518 21271 -7486
rect 21225 -7530 21271 -7518
rect 21373 -7518 21379 -7486
rect 21413 -7518 21419 -7486
rect 21373 -7530 21419 -7518
rect 21521 -7518 21527 -7486
rect 21561 -7518 21567 -7486
rect 21521 -7530 21567 -7518
rect 21669 -7518 21675 -7486
rect 21709 -7518 21715 -7486
rect 21669 -7530 21715 -7518
rect 21817 -7518 21823 -7486
rect 21857 -7518 21863 -7486
rect 21817 -7530 21863 -7518
rect 21965 -7518 21971 -7486
rect 22005 -7518 22011 -7486
rect 21965 -7530 22011 -7518
rect 22113 -7518 22119 -7486
rect 22153 -7518 22159 -7486
rect 22113 -7530 22159 -7518
rect 22261 -7518 22267 -7486
rect 22301 -7518 22307 -7486
rect 22261 -7530 22307 -7518
rect 22557 -7518 22563 -7486
rect 22597 -7518 22603 -7486
rect 22557 -7530 22603 -7518
rect 11499 -7716 11509 -7562
rect 11599 -7716 11609 -7562
rect 11647 -7716 11657 -7562
rect 11747 -7716 11757 -7562
rect 11795 -7716 11805 -7562
rect 11895 -7716 11905 -7562
rect 11943 -7716 11953 -7562
rect 12043 -7716 12053 -7562
rect 12091 -7716 12101 -7562
rect 12191 -7716 12201 -7562
rect 12239 -7716 12249 -7562
rect 12339 -7716 12349 -7562
rect 12387 -7716 12397 -7562
rect 12487 -7716 12497 -7562
rect 12535 -7716 12545 -7562
rect 12635 -7716 12645 -7562
rect 12683 -7716 12693 -7562
rect 12783 -7716 12793 -7562
rect 12831 -7716 12841 -7562
rect 12931 -7716 12941 -7562
rect 12979 -7716 12989 -7562
rect 13079 -7716 13089 -7562
rect 13127 -7716 13137 -7562
rect 13227 -7716 13237 -7562
rect 13275 -7716 13285 -7562
rect 13375 -7716 13385 -7562
rect 13423 -7716 13433 -7562
rect 13523 -7716 13533 -7562
rect 13571 -7716 13581 -7562
rect 13671 -7716 13681 -7562
rect 13719 -7716 13729 -7562
rect 13819 -7716 13829 -7562
rect 13867 -7716 13877 -7562
rect 13967 -7716 13977 -7562
rect 14015 -7716 14025 -7562
rect 14115 -7716 14125 -7562
rect 14163 -7716 14173 -7562
rect 14263 -7716 14273 -7562
rect 14311 -7716 14321 -7562
rect 14411 -7716 14421 -7562
rect 14459 -7716 14469 -7562
rect 14559 -7716 14569 -7562
rect 14607 -7716 14617 -7562
rect 14707 -7716 14717 -7562
rect 14755 -7716 14765 -7562
rect 14855 -7716 14865 -7562
rect 14903 -7716 14913 -7562
rect 15003 -7716 15013 -7562
rect 15051 -7716 15061 -7562
rect 15151 -7716 15161 -7562
rect 15199 -7716 15209 -7562
rect 15299 -7716 15309 -7562
rect 15347 -7716 15357 -7562
rect 15447 -7716 15457 -7562
rect 15495 -7716 15505 -7562
rect 15595 -7716 15605 -7562
rect 15643 -7716 15653 -7562
rect 15743 -7716 15753 -7562
rect 15791 -7716 15801 -7562
rect 15891 -7716 15901 -7562
rect 15939 -7716 15949 -7562
rect 16039 -7716 16049 -7562
rect 16087 -7716 16097 -7562
rect 16187 -7716 16197 -7562
rect 16235 -7716 16245 -7562
rect 16335 -7716 16345 -7562
rect 16383 -7716 16393 -7562
rect 16483 -7716 16493 -7562
rect 16531 -7716 16541 -7562
rect 16631 -7716 16641 -7562
rect 16679 -7716 16689 -7562
rect 16779 -7716 16789 -7562
rect 16827 -7716 16837 -7562
rect 16927 -7716 16937 -7562
rect 16975 -7716 16985 -7562
rect 17075 -7716 17085 -7562
rect 17123 -7716 17133 -7562
rect 17223 -7716 17233 -7562
rect 17271 -7716 17281 -7562
rect 17371 -7716 17381 -7562
rect 17419 -7716 17429 -7562
rect 17519 -7716 17529 -7562
rect 17567 -7716 17577 -7562
rect 17667 -7716 17677 -7562
rect 17715 -7716 17725 -7562
rect 17815 -7716 17825 -7562
rect 17863 -7716 17873 -7562
rect 17963 -7716 17973 -7562
rect 18011 -7716 18021 -7562
rect 18111 -7716 18121 -7562
rect 18159 -7716 18169 -7562
rect 18259 -7716 18269 -7562
rect 18307 -7716 18317 -7562
rect 18407 -7716 18417 -7562
rect 18455 -7716 18465 -7562
rect 18555 -7716 18565 -7562
rect 18603 -7716 18613 -7562
rect 18703 -7716 18713 -7562
rect 18751 -7716 18761 -7562
rect 18851 -7716 18861 -7562
rect 18899 -7716 18909 -7562
rect 18999 -7716 19009 -7562
rect 19047 -7716 19057 -7562
rect 19147 -7716 19157 -7562
rect 19195 -7716 19205 -7562
rect 19295 -7716 19305 -7562
rect 19343 -7716 19353 -7562
rect 19443 -7716 19453 -7562
rect 19491 -7716 19501 -7562
rect 19591 -7716 19601 -7562
rect 19639 -7716 19649 -7562
rect 19739 -7716 19749 -7562
rect 19787 -7716 19797 -7562
rect 19887 -7716 19897 -7562
rect 19935 -7716 19945 -7562
rect 20035 -7716 20045 -7562
rect 20083 -7716 20093 -7562
rect 20183 -7716 20193 -7562
rect 20231 -7716 20241 -7562
rect 20331 -7716 20341 -7562
rect 20379 -7716 20389 -7562
rect 20479 -7716 20489 -7562
rect 20527 -7716 20537 -7562
rect 20627 -7716 20637 -7562
rect 20675 -7716 20685 -7562
rect 20775 -7716 20785 -7562
rect 20823 -7716 20833 -7562
rect 20923 -7716 20933 -7562
rect 20971 -7716 20981 -7562
rect 21071 -7716 21081 -7562
rect 21119 -7716 21129 -7562
rect 21219 -7716 21229 -7562
rect 21267 -7716 21277 -7562
rect 21367 -7716 21377 -7562
rect 21415 -7716 21425 -7562
rect 21515 -7716 21525 -7562
rect 21563 -7716 21573 -7562
rect 21663 -7716 21673 -7562
rect 21711 -7716 21721 -7562
rect 21811 -7716 21821 -7562
rect 21859 -7716 21869 -7562
rect 21959 -7716 21969 -7562
rect 22007 -7716 22017 -7562
rect 22107 -7716 22117 -7562
rect 22155 -7716 22165 -7562
rect 22255 -7716 22265 -7562
rect 22303 -7716 22313 -7562
rect 22403 -7716 22413 -7562
rect 22451 -7716 22461 -7562
rect 22551 -7716 22561 -7562
rect 11457 -7760 11503 -7748
rect 3053 -7915 3063 -7761
rect 3121 -7915 3131 -7761
rect 3171 -7915 3181 -7761
rect 3239 -7915 3249 -7761
rect 3289 -7915 3299 -7761
rect 3357 -7915 3367 -7761
rect 3407 -7915 3417 -7761
rect 3475 -7915 3485 -7761
rect 3525 -7915 3535 -7761
rect 3593 -7915 3603 -7761
rect 3643 -7915 3653 -7761
rect 3711 -7915 3721 -7761
rect 3761 -7915 3771 -7761
rect 3829 -7915 3839 -7761
rect 3879 -7915 3889 -7761
rect 3947 -7915 3957 -7761
rect 3997 -7915 4007 -7761
rect 4065 -7915 4075 -7761
rect 4115 -7915 4125 -7761
rect 4183 -7915 4193 -7761
rect 4233 -7915 4243 -7761
rect 4301 -7915 4311 -7761
rect 4351 -7915 4361 -7761
rect 4419 -7915 4429 -7761
rect 4469 -7915 4479 -7761
rect 4537 -7915 4547 -7761
rect 4587 -7915 4597 -7761
rect 4655 -7915 4665 -7761
rect 4705 -7915 4715 -7761
rect 4773 -7915 4783 -7761
rect 5051 -7915 5061 -7761
rect 5119 -7915 5129 -7761
rect 5169 -7915 5179 -7761
rect 5237 -7915 5247 -7761
rect 5287 -7915 5297 -7761
rect 5355 -7915 5365 -7761
rect 5405 -7915 5415 -7761
rect 5473 -7915 5483 -7761
rect 5523 -7915 5533 -7761
rect 5591 -7915 5601 -7761
rect 5641 -7915 5651 -7761
rect 5709 -7915 5719 -7761
rect 5759 -7915 5769 -7761
rect 5827 -7915 5837 -7761
rect 5877 -7915 5887 -7761
rect 5945 -7915 5955 -7761
rect 5995 -7915 6005 -7761
rect 6063 -7915 6073 -7761
rect 6113 -7915 6123 -7761
rect 6181 -7915 6191 -7761
rect 6231 -7915 6241 -7761
rect 6299 -7915 6309 -7761
rect 6349 -7915 6359 -7761
rect 6417 -7915 6427 -7761
rect 6467 -7915 6477 -7761
rect 6535 -7915 6545 -7761
rect 6585 -7915 6595 -7761
rect 6653 -7915 6663 -7761
rect 6703 -7915 6713 -7761
rect 6771 -7915 6781 -7761
rect 11457 -7792 11463 -7760
rect 11497 -7792 11503 -7760
rect 11605 -7760 11651 -7748
rect 11605 -7792 11611 -7760
rect 11645 -7792 11651 -7760
rect 11753 -7760 11799 -7748
rect 11753 -7792 11759 -7760
rect 11793 -7792 11799 -7760
rect 11901 -7760 11947 -7748
rect 11901 -7792 11907 -7760
rect 11941 -7792 11947 -7760
rect 12049 -7760 12095 -7748
rect 12049 -7792 12055 -7760
rect 12089 -7792 12095 -7760
rect 12197 -7760 12243 -7748
rect 12197 -7792 12203 -7760
rect 12237 -7792 12243 -7760
rect 12345 -7760 12391 -7748
rect 12345 -7792 12351 -7760
rect 12385 -7792 12391 -7760
rect 12493 -7760 12539 -7748
rect 12493 -7792 12499 -7760
rect 12533 -7792 12539 -7760
rect 12641 -7760 12687 -7748
rect 12641 -7792 12647 -7760
rect 12681 -7792 12687 -7760
rect 12789 -7760 12835 -7748
rect 12789 -7792 12795 -7760
rect 12829 -7792 12835 -7760
rect 12937 -7760 12983 -7748
rect 12937 -7792 12943 -7760
rect 12977 -7792 12983 -7760
rect 13085 -7760 13131 -7748
rect 13085 -7792 13091 -7760
rect 13125 -7792 13131 -7760
rect 13233 -7760 13279 -7748
rect 13233 -7792 13239 -7760
rect 13273 -7792 13279 -7760
rect 13381 -7760 13427 -7748
rect 13381 -7792 13387 -7760
rect 13421 -7792 13427 -7760
rect 13529 -7760 13575 -7748
rect 13529 -7792 13535 -7760
rect 13569 -7792 13575 -7760
rect 13677 -7760 13723 -7748
rect 13677 -7792 13683 -7760
rect 13717 -7792 13723 -7760
rect 13825 -7760 13871 -7748
rect 13825 -7792 13831 -7760
rect 13865 -7792 13871 -7760
rect 13973 -7760 14019 -7748
rect 13973 -7792 13979 -7760
rect 14013 -7792 14019 -7760
rect 14121 -7760 14167 -7748
rect 14121 -7792 14127 -7760
rect 14161 -7792 14167 -7760
rect 14269 -7760 14315 -7748
rect 14269 -7792 14275 -7760
rect 14309 -7792 14315 -7760
rect 14417 -7760 14463 -7748
rect 14417 -7792 14423 -7760
rect 14457 -7792 14463 -7760
rect 14565 -7760 14611 -7748
rect 14565 -7792 14571 -7760
rect 14605 -7792 14611 -7760
rect 14713 -7760 14759 -7748
rect 14713 -7792 14719 -7760
rect 14753 -7792 14759 -7760
rect 14861 -7760 14907 -7748
rect 14861 -7792 14867 -7760
rect 14901 -7792 14907 -7760
rect 15009 -7760 15055 -7748
rect 15009 -7792 15015 -7760
rect 15049 -7792 15055 -7760
rect 15157 -7760 15203 -7748
rect 15157 -7792 15163 -7760
rect 15197 -7792 15203 -7760
rect 15305 -7760 15351 -7748
rect 15305 -7792 15311 -7760
rect 15345 -7792 15351 -7760
rect 15453 -7760 15499 -7748
rect 15453 -7792 15459 -7760
rect 15493 -7792 15499 -7760
rect 15601 -7760 15647 -7748
rect 15601 -7792 15607 -7760
rect 15641 -7792 15647 -7760
rect 15749 -7760 15795 -7748
rect 15749 -7792 15755 -7760
rect 15789 -7792 15795 -7760
rect 15897 -7760 15943 -7748
rect 15897 -7792 15903 -7760
rect 15937 -7792 15943 -7760
rect 16045 -7760 16091 -7748
rect 16045 -7792 16051 -7760
rect 16085 -7792 16091 -7760
rect 16193 -7760 16239 -7748
rect 16193 -7792 16199 -7760
rect 16233 -7792 16239 -7760
rect 16341 -7760 16387 -7748
rect 16341 -7792 16347 -7760
rect 16381 -7792 16387 -7760
rect 16489 -7760 16535 -7748
rect 16489 -7792 16495 -7760
rect 16529 -7792 16535 -7760
rect 16637 -7760 16683 -7748
rect 16637 -7792 16643 -7760
rect 16677 -7792 16683 -7760
rect 16785 -7760 16831 -7748
rect 16785 -7792 16791 -7760
rect 16825 -7792 16831 -7760
rect 16933 -7760 16979 -7748
rect 16933 -7792 16939 -7760
rect 16973 -7792 16979 -7760
rect 17081 -7760 17127 -7748
rect 17081 -7792 17087 -7760
rect 17121 -7792 17127 -7760
rect 17229 -7760 17275 -7748
rect 17229 -7792 17235 -7760
rect 17269 -7792 17275 -7760
rect 17377 -7760 17423 -7748
rect 17377 -7792 17383 -7760
rect 17417 -7792 17423 -7760
rect 17525 -7760 17571 -7748
rect 17525 -7792 17531 -7760
rect 17565 -7792 17571 -7760
rect 17673 -7760 17719 -7748
rect 17673 -7792 17679 -7760
rect 17713 -7792 17719 -7760
rect 17821 -7760 17867 -7748
rect 17821 -7792 17827 -7760
rect 17861 -7792 17867 -7760
rect 17969 -7760 18015 -7748
rect 17969 -7792 17975 -7760
rect 18009 -7792 18015 -7760
rect 18117 -7760 18163 -7748
rect 18117 -7792 18123 -7760
rect 18157 -7792 18163 -7760
rect 18265 -7760 18311 -7748
rect 18265 -7792 18271 -7760
rect 18305 -7792 18311 -7760
rect 18413 -7760 18459 -7748
rect 18413 -7792 18419 -7760
rect 18453 -7792 18459 -7760
rect 18561 -7760 18607 -7748
rect 18561 -7792 18567 -7760
rect 18601 -7792 18607 -7760
rect 18709 -7760 18755 -7748
rect 18709 -7792 18715 -7760
rect 18749 -7792 18755 -7760
rect 18857 -7760 18903 -7748
rect 18857 -7792 18863 -7760
rect 18897 -7792 18903 -7760
rect 19005 -7760 19051 -7748
rect 19005 -7792 19011 -7760
rect 19045 -7792 19051 -7760
rect 19153 -7760 19199 -7748
rect 19153 -7792 19159 -7760
rect 19193 -7792 19199 -7760
rect 19301 -7760 19347 -7748
rect 19301 -7792 19307 -7760
rect 19341 -7792 19347 -7760
rect 19449 -7760 19495 -7748
rect 19449 -7792 19455 -7760
rect 19489 -7792 19495 -7760
rect 19597 -7760 19643 -7748
rect 19597 -7792 19603 -7760
rect 19637 -7792 19643 -7760
rect 19745 -7760 19791 -7748
rect 19745 -7792 19751 -7760
rect 19785 -7792 19791 -7760
rect 19893 -7760 19939 -7748
rect 19893 -7792 19899 -7760
rect 19933 -7792 19939 -7760
rect 20041 -7760 20087 -7748
rect 20041 -7792 20047 -7760
rect 20081 -7792 20087 -7760
rect 20189 -7760 20235 -7748
rect 20189 -7792 20195 -7760
rect 20229 -7792 20235 -7760
rect 20337 -7760 20383 -7748
rect 20337 -7792 20343 -7760
rect 20377 -7792 20383 -7760
rect 20485 -7760 20531 -7748
rect 20485 -7792 20491 -7760
rect 20525 -7792 20531 -7760
rect 20633 -7760 20679 -7748
rect 20633 -7792 20639 -7760
rect 20673 -7792 20679 -7760
rect 20781 -7760 20827 -7748
rect 20781 -7792 20787 -7760
rect 20821 -7792 20827 -7760
rect 20929 -7760 20975 -7748
rect 20929 -7792 20935 -7760
rect 20969 -7792 20975 -7760
rect 21077 -7760 21123 -7748
rect 21077 -7792 21083 -7760
rect 21117 -7792 21123 -7760
rect 21225 -7760 21271 -7748
rect 21225 -7792 21231 -7760
rect 21265 -7792 21271 -7760
rect 21373 -7760 21419 -7748
rect 21373 -7792 21379 -7760
rect 21413 -7792 21419 -7760
rect 21521 -7760 21567 -7748
rect 21521 -7792 21527 -7760
rect 21561 -7792 21567 -7760
rect 21669 -7760 21715 -7748
rect 21669 -7792 21675 -7760
rect 21709 -7792 21715 -7760
rect 21817 -7760 21863 -7748
rect 21817 -7792 21823 -7760
rect 21857 -7792 21863 -7760
rect 21965 -7760 22011 -7748
rect 21965 -7792 21971 -7760
rect 22005 -7792 22011 -7760
rect 22113 -7760 22159 -7748
rect 22113 -7792 22119 -7760
rect 22153 -7792 22159 -7760
rect 22261 -7760 22307 -7748
rect 22261 -7792 22267 -7760
rect 22301 -7792 22307 -7760
rect 11444 -8632 11454 -7792
rect 11506 -8632 11516 -7792
rect 11592 -8632 11602 -7792
rect 11654 -8632 11664 -7792
rect 11740 -8632 11750 -7792
rect 11802 -8632 11812 -7792
rect 11888 -8632 11898 -7792
rect 11950 -8632 11960 -7792
rect 12036 -8632 12046 -7792
rect 12098 -8632 12108 -7792
rect 12184 -8632 12194 -7792
rect 12246 -8632 12256 -7792
rect 12332 -8632 12342 -7792
rect 12394 -8632 12404 -7792
rect 12480 -8632 12490 -7792
rect 12542 -8632 12552 -7792
rect 12628 -8632 12638 -7792
rect 12690 -8632 12700 -7792
rect 12776 -8632 12786 -7792
rect 12838 -8632 12848 -7792
rect 12924 -8632 12934 -7792
rect 12986 -8632 12996 -7792
rect 13072 -8632 13082 -7792
rect 13134 -8632 13144 -7792
rect 13220 -8632 13230 -7792
rect 13282 -8632 13292 -7792
rect 13368 -8632 13378 -7792
rect 13430 -8632 13440 -7792
rect 13516 -8632 13526 -7792
rect 13578 -8632 13588 -7792
rect 13664 -8632 13674 -7792
rect 13726 -8632 13736 -7792
rect 13812 -8632 13822 -7792
rect 13874 -8632 13884 -7792
rect 13960 -8632 13970 -7792
rect 14022 -8632 14032 -7792
rect 14108 -8632 14118 -7792
rect 14170 -8632 14180 -7792
rect 14256 -8632 14266 -7792
rect 14318 -8632 14328 -7792
rect 14404 -8632 14414 -7792
rect 14466 -8632 14476 -7792
rect 14552 -8632 14562 -7792
rect 14614 -8632 14624 -7792
rect 14700 -8632 14710 -7792
rect 14762 -8632 14772 -7792
rect 14848 -8632 14858 -7792
rect 14910 -8632 14920 -7792
rect 14996 -8632 15006 -7792
rect 15058 -8632 15068 -7792
rect 15144 -8632 15154 -7792
rect 15206 -8632 15216 -7792
rect 15292 -8632 15302 -7792
rect 15354 -8632 15364 -7792
rect 15440 -8632 15450 -7792
rect 15502 -8632 15512 -7792
rect 15588 -8632 15598 -7792
rect 15650 -8632 15660 -7792
rect 15736 -8632 15746 -7792
rect 15798 -8632 15808 -7792
rect 15884 -8632 15894 -7792
rect 15946 -8632 15956 -7792
rect 16032 -8632 16042 -7792
rect 16094 -8632 16104 -7792
rect 16180 -8632 16190 -7792
rect 16242 -8632 16252 -7792
rect 16328 -8632 16338 -7792
rect 16390 -8632 16400 -7792
rect 16476 -8632 16486 -7792
rect 16538 -8632 16548 -7792
rect 16624 -8632 16634 -7792
rect 16686 -8632 16696 -7792
rect 16772 -8632 16782 -7792
rect 16834 -8632 16844 -7792
rect 16920 -8632 16930 -7792
rect 16982 -8632 16992 -7792
rect 17068 -8632 17078 -7792
rect 17130 -8632 17140 -7792
rect 17216 -8632 17226 -7792
rect 17278 -8632 17288 -7792
rect 17364 -8632 17374 -7792
rect 17426 -8632 17436 -7792
rect 17512 -8632 17522 -7792
rect 17574 -8632 17584 -7792
rect 17660 -8632 17670 -7792
rect 17722 -8632 17732 -7792
rect 17808 -8632 17818 -7792
rect 17870 -8632 17880 -7792
rect 17956 -8632 17966 -7792
rect 18018 -8632 18028 -7792
rect 18104 -8632 18114 -7792
rect 18166 -8632 18176 -7792
rect 18252 -8632 18262 -7792
rect 18314 -8632 18324 -7792
rect 18400 -8632 18410 -7792
rect 18462 -8632 18472 -7792
rect 18548 -8632 18558 -7792
rect 18610 -8632 18620 -7792
rect 18696 -8632 18706 -7792
rect 18758 -8632 18768 -7792
rect 18844 -8632 18854 -7792
rect 18906 -8632 18916 -7792
rect 18992 -8632 19002 -7792
rect 19054 -8632 19064 -7792
rect 19140 -8632 19150 -7792
rect 19202 -8632 19212 -7792
rect 19288 -8632 19298 -7792
rect 19350 -8632 19360 -7792
rect 19436 -8632 19446 -7792
rect 19498 -8632 19508 -7792
rect 19584 -8632 19594 -7792
rect 19646 -8632 19656 -7792
rect 19732 -8632 19742 -7792
rect 19794 -8632 19804 -7792
rect 19880 -8632 19890 -7792
rect 19942 -8632 19952 -7792
rect 20028 -8632 20038 -7792
rect 20090 -8632 20100 -7792
rect 20176 -8632 20186 -7792
rect 20238 -8632 20248 -7792
rect 20324 -8632 20334 -7792
rect 20386 -8632 20396 -7792
rect 20472 -8632 20482 -7792
rect 20534 -8632 20544 -7792
rect 20620 -8632 20630 -7792
rect 20682 -8632 20692 -7792
rect 20768 -8632 20778 -7792
rect 20830 -8632 20840 -7792
rect 20916 -8632 20926 -7792
rect 20978 -8632 20988 -7792
rect 21064 -8632 21074 -7792
rect 21126 -8632 21136 -7792
rect 21212 -8632 21222 -7792
rect 21274 -8632 21284 -7792
rect 21360 -8632 21370 -7792
rect 21422 -8632 21432 -7792
rect 21508 -8632 21518 -7792
rect 21570 -8632 21580 -7792
rect 21656 -8632 21666 -7792
rect 21718 -8632 21728 -7792
rect 21804 -8632 21814 -7792
rect 21866 -8632 21876 -7792
rect 21952 -8632 21962 -7792
rect 22014 -8632 22024 -7792
rect 22100 -8632 22110 -7792
rect 22162 -8632 22172 -7792
rect 22248 -8632 22258 -7792
rect 22310 -8632 22320 -7792
rect 22396 -8632 22406 -7792
rect 22458 -8632 22468 -7792
rect 22544 -8632 22554 -7792
rect 22606 -8632 22616 -7792
rect 22820 -7926 22830 -7086
rect 22882 -7926 22892 -7086
rect 23045 -7926 23055 -7086
rect 23107 -7926 23117 -7086
rect 23223 -7939 23233 -7099
rect 23285 -7939 23295 -7099
rect 11457 -8636 11463 -8632
rect 11497 -8636 11503 -8632
rect 11457 -8648 11503 -8636
rect 11605 -8636 11611 -8632
rect 11645 -8636 11651 -8632
rect 11605 -8648 11651 -8636
rect 11753 -8636 11759 -8632
rect 11793 -8636 11799 -8632
rect 11753 -8648 11799 -8636
rect 11901 -8636 11907 -8632
rect 11941 -8636 11947 -8632
rect 11901 -8648 11947 -8636
rect 12049 -8636 12055 -8632
rect 12089 -8636 12095 -8632
rect 12049 -8648 12095 -8636
rect 12197 -8636 12203 -8632
rect 12237 -8636 12243 -8632
rect 12197 -8648 12243 -8636
rect 12345 -8636 12351 -8632
rect 12385 -8636 12391 -8632
rect 12345 -8648 12391 -8636
rect 12493 -8636 12499 -8632
rect 12533 -8636 12539 -8632
rect 12493 -8648 12539 -8636
rect 12641 -8636 12647 -8632
rect 12681 -8636 12687 -8632
rect 12641 -8648 12687 -8636
rect 12789 -8636 12795 -8632
rect 12829 -8636 12835 -8632
rect 12789 -8648 12835 -8636
rect 12937 -8636 12943 -8632
rect 12977 -8636 12983 -8632
rect 12937 -8648 12983 -8636
rect 13085 -8636 13091 -8632
rect 13125 -8636 13131 -8632
rect 13085 -8648 13131 -8636
rect 13233 -8636 13239 -8632
rect 13273 -8636 13279 -8632
rect 13233 -8648 13279 -8636
rect 13381 -8636 13387 -8632
rect 13421 -8636 13427 -8632
rect 13381 -8648 13427 -8636
rect 13529 -8636 13535 -8632
rect 13569 -8636 13575 -8632
rect 13529 -8648 13575 -8636
rect 13677 -8636 13683 -8632
rect 13717 -8636 13723 -8632
rect 13677 -8648 13723 -8636
rect 13825 -8636 13831 -8632
rect 13865 -8636 13871 -8632
rect 13825 -8648 13871 -8636
rect 13973 -8636 13979 -8632
rect 14013 -8636 14019 -8632
rect 13973 -8648 14019 -8636
rect 14121 -8636 14127 -8632
rect 14161 -8636 14167 -8632
rect 14121 -8648 14167 -8636
rect 14269 -8636 14275 -8632
rect 14309 -8636 14315 -8632
rect 14269 -8648 14315 -8636
rect 14417 -8636 14423 -8632
rect 14457 -8636 14463 -8632
rect 14417 -8648 14463 -8636
rect 14565 -8636 14571 -8632
rect 14605 -8636 14611 -8632
rect 14565 -8648 14611 -8636
rect 14713 -8636 14719 -8632
rect 14753 -8636 14759 -8632
rect 14713 -8648 14759 -8636
rect 14861 -8636 14867 -8632
rect 14901 -8636 14907 -8632
rect 14861 -8648 14907 -8636
rect 15009 -8636 15015 -8632
rect 15049 -8636 15055 -8632
rect 15009 -8648 15055 -8636
rect 15157 -8636 15163 -8632
rect 15197 -8636 15203 -8632
rect 15157 -8648 15203 -8636
rect 15305 -8636 15311 -8632
rect 15345 -8636 15351 -8632
rect 15305 -8648 15351 -8636
rect 15453 -8636 15459 -8632
rect 15493 -8636 15499 -8632
rect 15453 -8648 15499 -8636
rect 15601 -8636 15607 -8632
rect 15641 -8636 15647 -8632
rect 15601 -8648 15647 -8636
rect 15749 -8636 15755 -8632
rect 15789 -8636 15795 -8632
rect 15749 -8648 15795 -8636
rect 15897 -8636 15903 -8632
rect 15937 -8636 15943 -8632
rect 15897 -8648 15943 -8636
rect 16045 -8636 16051 -8632
rect 16085 -8636 16091 -8632
rect 16045 -8648 16091 -8636
rect 16193 -8636 16199 -8632
rect 16233 -8636 16239 -8632
rect 16193 -8648 16239 -8636
rect 16341 -8636 16347 -8632
rect 16381 -8636 16387 -8632
rect 16341 -8648 16387 -8636
rect 16489 -8636 16495 -8632
rect 16529 -8636 16535 -8632
rect 16489 -8648 16535 -8636
rect 16637 -8636 16643 -8632
rect 16677 -8636 16683 -8632
rect 16637 -8648 16683 -8636
rect 16785 -8636 16791 -8632
rect 16825 -8636 16831 -8632
rect 16785 -8648 16831 -8636
rect 16933 -8636 16939 -8632
rect 16973 -8636 16979 -8632
rect 16933 -8648 16979 -8636
rect 17081 -8636 17087 -8632
rect 17121 -8636 17127 -8632
rect 17081 -8648 17127 -8636
rect 17229 -8636 17235 -8632
rect 17269 -8636 17275 -8632
rect 17229 -8648 17275 -8636
rect 17377 -8636 17383 -8632
rect 17417 -8636 17423 -8632
rect 17377 -8648 17423 -8636
rect 17525 -8636 17531 -8632
rect 17565 -8636 17571 -8632
rect 17525 -8648 17571 -8636
rect 17673 -8636 17679 -8632
rect 17713 -8636 17719 -8632
rect 17673 -8648 17719 -8636
rect 17821 -8636 17827 -8632
rect 17861 -8636 17867 -8632
rect 17821 -8648 17867 -8636
rect 17969 -8636 17975 -8632
rect 18009 -8636 18015 -8632
rect 17969 -8648 18015 -8636
rect 18117 -8636 18123 -8632
rect 18157 -8636 18163 -8632
rect 18117 -8648 18163 -8636
rect 18265 -8636 18271 -8632
rect 18305 -8636 18311 -8632
rect 18265 -8648 18311 -8636
rect 18413 -8636 18419 -8632
rect 18453 -8636 18459 -8632
rect 18413 -8648 18459 -8636
rect 18561 -8636 18567 -8632
rect 18601 -8636 18607 -8632
rect 18561 -8648 18607 -8636
rect 18709 -8636 18715 -8632
rect 18749 -8636 18755 -8632
rect 18709 -8648 18755 -8636
rect 18857 -8636 18863 -8632
rect 18897 -8636 18903 -8632
rect 18857 -8648 18903 -8636
rect 19005 -8636 19011 -8632
rect 19045 -8636 19051 -8632
rect 19005 -8648 19051 -8636
rect 19153 -8636 19159 -8632
rect 19193 -8636 19199 -8632
rect 19153 -8648 19199 -8636
rect 19301 -8636 19307 -8632
rect 19341 -8636 19347 -8632
rect 19301 -8648 19347 -8636
rect 19449 -8636 19455 -8632
rect 19489 -8636 19495 -8632
rect 19449 -8648 19495 -8636
rect 19597 -8636 19603 -8632
rect 19637 -8636 19643 -8632
rect 19597 -8648 19643 -8636
rect 19745 -8636 19751 -8632
rect 19785 -8636 19791 -8632
rect 19745 -8648 19791 -8636
rect 19893 -8636 19899 -8632
rect 19933 -8636 19939 -8632
rect 19893 -8648 19939 -8636
rect 20041 -8636 20047 -8632
rect 20081 -8636 20087 -8632
rect 20041 -8648 20087 -8636
rect 20189 -8636 20195 -8632
rect 20229 -8636 20235 -8632
rect 20189 -8648 20235 -8636
rect 20337 -8636 20343 -8632
rect 20377 -8636 20383 -8632
rect 20337 -8648 20383 -8636
rect 20485 -8636 20491 -8632
rect 20525 -8636 20531 -8632
rect 20485 -8648 20531 -8636
rect 20633 -8636 20639 -8632
rect 20673 -8636 20679 -8632
rect 20633 -8648 20679 -8636
rect 20781 -8636 20787 -8632
rect 20821 -8636 20827 -8632
rect 20781 -8648 20827 -8636
rect 20929 -8636 20935 -8632
rect 20969 -8636 20975 -8632
rect 20929 -8648 20975 -8636
rect 21077 -8636 21083 -8632
rect 21117 -8636 21123 -8632
rect 21077 -8648 21123 -8636
rect 21225 -8636 21231 -8632
rect 21265 -8636 21271 -8632
rect 21225 -8648 21271 -8636
rect 21373 -8636 21379 -8632
rect 21413 -8636 21419 -8632
rect 21373 -8648 21419 -8636
rect 21521 -8636 21527 -8632
rect 21561 -8636 21567 -8632
rect 21521 -8648 21567 -8636
rect 21669 -8636 21675 -8632
rect 21709 -8636 21715 -8632
rect 21669 -8648 21715 -8636
rect 21817 -8636 21823 -8632
rect 21857 -8636 21863 -8632
rect 21817 -8648 21863 -8636
rect 21965 -8636 21971 -8632
rect 22005 -8636 22011 -8632
rect 21965 -8648 22011 -8636
rect 22113 -8636 22119 -8632
rect 22153 -8636 22159 -8632
rect 22113 -8648 22159 -8636
rect 22261 -8636 22267 -8632
rect 22301 -8636 22307 -8632
rect 22261 -8648 22307 -8636
<< via1 >>
rect 6530 2087 6582 2687
rect 6766 2675 6818 2687
rect 6766 2099 6788 2675
rect 6788 2099 6818 2675
rect 6766 2087 6818 2099
rect 4601 2040 4659 2044
rect 4601 2006 4613 2040
rect 4613 2006 4647 2040
rect 4647 2006 4659 2040
rect 4601 1952 4659 2006
rect 4719 2040 4777 2044
rect 4719 2006 4731 2040
rect 4731 2006 4765 2040
rect 4765 2006 4777 2040
rect 4719 1952 4777 2006
rect 4837 2040 4895 2044
rect 4837 2006 4849 2040
rect 4849 2006 4883 2040
rect 4883 2006 4895 2040
rect 4837 1952 4895 2006
rect 4955 2040 5013 2044
rect 4955 2006 4967 2040
rect 4967 2006 5001 2040
rect 5001 2006 5013 2040
rect 4955 1952 5013 2006
rect 5073 2040 5131 2044
rect 5073 2006 5085 2040
rect 5085 2006 5119 2040
rect 5119 2006 5131 2040
rect 5073 1952 5131 2006
rect 5191 2040 5249 2044
rect 5191 2006 5203 2040
rect 5203 2006 5237 2040
rect 5237 2006 5249 2040
rect 5191 1952 5249 2006
rect 5309 2040 5367 2044
rect 5309 2006 5321 2040
rect 5321 2006 5355 2040
rect 5355 2006 5367 2040
rect 5309 1952 5367 2006
rect 5427 2040 5485 2044
rect 5427 2006 5439 2040
rect 5439 2006 5473 2040
rect 5473 2006 5485 2040
rect 5427 1952 5485 2006
rect 5545 2040 5603 2044
rect 5545 2006 5557 2040
rect 5557 2006 5591 2040
rect 5591 2006 5603 2040
rect 5545 1952 5603 2006
rect 5663 2040 5721 2044
rect 5663 2006 5675 2040
rect 5675 2006 5709 2040
rect 5709 2006 5721 2040
rect 5663 1952 5721 2006
rect 5781 2040 5839 2044
rect 5781 2006 5793 2040
rect 5793 2006 5827 2040
rect 5827 2006 5839 2040
rect 5781 1952 5839 2006
rect 5899 2040 5957 2044
rect 5899 2006 5911 2040
rect 5911 2006 5945 2040
rect 5945 2006 5957 2040
rect 5899 1952 5957 2006
rect 6017 2040 6075 2044
rect 6017 2006 6029 2040
rect 6029 2006 6063 2040
rect 6063 2006 6075 2040
rect 6017 1952 6075 2006
rect 6135 2040 6193 2044
rect 6135 2006 6147 2040
rect 6147 2006 6181 2040
rect 6181 2006 6193 2040
rect 6135 1952 6193 2006
rect 6253 2040 6311 2044
rect 6253 2006 6265 2040
rect 6265 2006 6299 2040
rect 6299 2006 6311 2040
rect 6253 1952 6311 2006
rect 6599 1952 6657 2044
rect 6717 1952 6775 2044
rect 6835 2040 6893 2044
rect 6835 2006 6847 2040
rect 6847 2006 6881 2040
rect 6881 2006 6893 2040
rect 6835 1952 6893 2006
rect 6953 2040 7011 2044
rect 6953 2006 6965 2040
rect 6965 2006 6999 2040
rect 6999 2006 7011 2040
rect 6953 1952 7011 2006
rect 7071 2040 7129 2044
rect 7071 2006 7083 2040
rect 7083 2006 7117 2040
rect 7117 2006 7129 2040
rect 7071 1952 7129 2006
rect 7189 2040 7247 2044
rect 7189 2006 7201 2040
rect 7201 2006 7235 2040
rect 7235 2006 7247 2040
rect 7189 1952 7247 2006
rect 7307 2040 7365 2044
rect 7307 2006 7319 2040
rect 7319 2006 7353 2040
rect 7353 2006 7365 2040
rect 7307 1952 7365 2006
rect 7425 2040 7483 2044
rect 7425 2006 7437 2040
rect 7437 2006 7471 2040
rect 7471 2006 7483 2040
rect 7425 1952 7483 2006
rect 7543 2040 7601 2044
rect 7543 2006 7555 2040
rect 7555 2006 7589 2040
rect 7589 2006 7601 2040
rect 7543 1952 7601 2006
rect 7661 2040 7719 2044
rect 7661 2006 7673 2040
rect 7673 2006 7707 2040
rect 7707 2006 7719 2040
rect 7661 1952 7719 2006
rect 7779 2040 7837 2044
rect 7779 2006 7791 2040
rect 7791 2006 7825 2040
rect 7825 2006 7837 2040
rect 7779 1952 7837 2006
rect 7897 2040 7955 2044
rect 7897 2006 7909 2040
rect 7909 2006 7943 2040
rect 7943 2006 7955 2040
rect 7897 1952 7955 2006
rect 8015 2040 8073 2044
rect 8015 2006 8027 2040
rect 8027 2006 8061 2040
rect 8061 2006 8073 2040
rect 8015 1952 8073 2006
rect 8133 2040 8191 2044
rect 8133 2006 8145 2040
rect 8145 2006 8179 2040
rect 8179 2006 8191 2040
rect 8133 1952 8191 2006
rect 8251 2040 8309 2044
rect 8251 2006 8263 2040
rect 8263 2006 8297 2040
rect 8297 2006 8309 2040
rect 8251 1952 8309 2006
rect 8597 2040 8655 2044
rect 8597 2006 8609 2040
rect 8609 2006 8643 2040
rect 8643 2006 8655 2040
rect 8597 1952 8655 2006
rect 8715 2040 8773 2044
rect 8715 2006 8727 2040
rect 8727 2006 8761 2040
rect 8761 2006 8773 2040
rect 8715 1952 8773 2006
rect 8833 2040 8891 2044
rect 8833 2006 8845 2040
rect 8845 2006 8879 2040
rect 8879 2006 8891 2040
rect 8833 1952 8891 2006
rect 8951 2040 9009 2044
rect 8951 2006 8963 2040
rect 8963 2006 8997 2040
rect 8997 2006 9009 2040
rect 8951 1952 9009 2006
rect 9069 2040 9127 2044
rect 9069 2006 9081 2040
rect 9081 2006 9115 2040
rect 9115 2006 9127 2040
rect 9069 1952 9127 2006
rect 9187 2040 9245 2044
rect 9187 2006 9199 2040
rect 9199 2006 9233 2040
rect 9233 2006 9245 2040
rect 9187 1952 9245 2006
rect 9305 2040 9363 2044
rect 9305 2006 9317 2040
rect 9317 2006 9351 2040
rect 9351 2006 9363 2040
rect 9305 1952 9363 2006
rect 9423 2040 9481 2044
rect 9423 2006 9435 2040
rect 9435 2006 9469 2040
rect 9469 2006 9481 2040
rect 9423 1952 9481 2006
rect 9541 2040 9599 2044
rect 9541 2006 9553 2040
rect 9553 2006 9587 2040
rect 9587 2006 9599 2040
rect 9541 1952 9599 2006
rect 9659 2040 9717 2044
rect 9659 2006 9671 2040
rect 9671 2006 9705 2040
rect 9705 2006 9717 2040
rect 9659 1952 9717 2006
rect 9777 2040 9835 2044
rect 9777 2006 9789 2040
rect 9789 2006 9823 2040
rect 9823 2006 9835 2040
rect 9777 1952 9835 2006
rect 9895 2040 9953 2044
rect 9895 2006 9907 2040
rect 9907 2006 9941 2040
rect 9941 2006 9953 2040
rect 9895 1952 9953 2006
rect 10013 2040 10071 2044
rect 10013 2006 10025 2040
rect 10025 2006 10059 2040
rect 10059 2006 10071 2040
rect 10013 1952 10071 2006
rect 10131 2040 10189 2044
rect 10131 2006 10143 2040
rect 10143 2006 10177 2040
rect 10177 2006 10189 2040
rect 10131 1952 10189 2006
rect 10249 2040 10307 2044
rect 10249 2006 10261 2040
rect 10261 2006 10295 2040
rect 10295 2006 10307 2040
rect 10249 1952 10307 2006
rect 12547 1891 12605 2045
rect 12665 2039 12723 2045
rect 12665 2005 12677 2039
rect 12677 2005 12711 2039
rect 12711 2005 12723 2039
rect 12665 1931 12723 2005
rect 12665 1897 12677 1931
rect 12677 1897 12711 1931
rect 12711 1897 12723 1931
rect 12665 1891 12723 1897
rect 12783 2039 12841 2045
rect 12783 2005 12795 2039
rect 12795 2005 12829 2039
rect 12829 2005 12841 2039
rect 12783 1931 12841 2005
rect 12783 1897 12795 1931
rect 12795 1897 12829 1931
rect 12829 1897 12841 1931
rect 12783 1891 12841 1897
rect 12901 2039 12959 2045
rect 12901 2005 12913 2039
rect 12913 2005 12947 2039
rect 12947 2005 12959 2039
rect 12901 1931 12959 2005
rect 12901 1897 12913 1931
rect 12913 1897 12947 1931
rect 12947 1897 12959 1931
rect 12901 1891 12959 1897
rect 13019 2039 13077 2045
rect 13019 2005 13031 2039
rect 13031 2005 13065 2039
rect 13065 2005 13077 2039
rect 13019 1931 13077 2005
rect 13019 1897 13031 1931
rect 13031 1897 13065 1931
rect 13065 1897 13077 1931
rect 13019 1891 13077 1897
rect 13137 2039 13195 2045
rect 13137 2005 13149 2039
rect 13149 2005 13183 2039
rect 13183 2005 13195 2039
rect 13137 1931 13195 2005
rect 13137 1897 13149 1931
rect 13149 1897 13183 1931
rect 13183 1897 13195 1931
rect 13137 1891 13195 1897
rect 13255 2039 13313 2045
rect 13255 2005 13267 2039
rect 13267 2005 13301 2039
rect 13301 2005 13313 2039
rect 13255 1931 13313 2005
rect 13255 1897 13267 1931
rect 13267 1897 13301 1931
rect 13301 1897 13313 1931
rect 13255 1891 13313 1897
rect 13373 2039 13431 2045
rect 13373 2005 13385 2039
rect 13385 2005 13419 2039
rect 13419 2005 13431 2039
rect 13373 1931 13431 2005
rect 13373 1897 13385 1931
rect 13385 1897 13419 1931
rect 13419 1897 13431 1931
rect 13373 1891 13431 1897
rect 13491 2039 13549 2045
rect 13491 2005 13503 2039
rect 13503 2005 13537 2039
rect 13537 2005 13549 2039
rect 13491 1931 13549 2005
rect 13491 1897 13503 1931
rect 13503 1897 13537 1931
rect 13537 1897 13549 1931
rect 13491 1891 13549 1897
rect 13609 2039 13667 2045
rect 13609 2005 13621 2039
rect 13621 2005 13655 2039
rect 13655 2005 13667 2039
rect 13609 1931 13667 2005
rect 13609 1897 13621 1931
rect 13621 1897 13655 1931
rect 13655 1897 13667 1931
rect 13609 1891 13667 1897
rect 13727 2039 13785 2045
rect 13727 2005 13739 2039
rect 13739 2005 13773 2039
rect 13773 2005 13785 2039
rect 13727 1931 13785 2005
rect 13727 1897 13739 1931
rect 13739 1897 13773 1931
rect 13773 1897 13785 1931
rect 13727 1891 13785 1897
rect 13845 2039 13903 2045
rect 13845 2005 13857 2039
rect 13857 2005 13891 2039
rect 13891 2005 13903 2039
rect 13845 1931 13903 2005
rect 13845 1897 13857 1931
rect 13857 1897 13891 1931
rect 13891 1897 13903 1931
rect 13845 1891 13903 1897
rect 13963 2039 14021 2045
rect 13963 2005 13975 2039
rect 13975 2005 14009 2039
rect 14009 2005 14021 2039
rect 13963 1931 14021 2005
rect 13963 1897 13975 1931
rect 13975 1897 14009 1931
rect 14009 1897 14021 1931
rect 13963 1891 14021 1897
rect 14081 2039 14139 2045
rect 14081 2005 14093 2039
rect 14093 2005 14127 2039
rect 14127 2005 14139 2039
rect 14081 1931 14139 2005
rect 14081 1897 14093 1931
rect 14093 1897 14127 1931
rect 14127 1897 14139 1931
rect 14081 1891 14139 1897
rect 14199 2039 14257 2045
rect 14199 2005 14211 2039
rect 14211 2005 14245 2039
rect 14245 2005 14257 2039
rect 14199 1931 14257 2005
rect 14199 1897 14211 1931
rect 14211 1897 14245 1931
rect 14245 1897 14257 1931
rect 14199 1891 14257 1897
rect 14317 2039 14375 2045
rect 14317 2005 14329 2039
rect 14329 2005 14363 2039
rect 14363 2005 14375 2039
rect 14317 1931 14375 2005
rect 14317 1897 14329 1931
rect 14329 1897 14363 1931
rect 14363 1897 14375 1931
rect 14317 1891 14375 1897
rect 14435 2039 14493 2045
rect 14435 2005 14447 2039
rect 14447 2005 14481 2039
rect 14481 2005 14493 2039
rect 14435 1931 14493 2005
rect 14435 1897 14447 1931
rect 14447 1897 14481 1931
rect 14481 1897 14493 1931
rect 14435 1891 14493 1897
rect 14553 2039 14611 2045
rect 14553 2005 14565 2039
rect 14565 2005 14599 2039
rect 14599 2005 14611 2039
rect 14553 1931 14611 2005
rect 14553 1897 14565 1931
rect 14565 1897 14599 1931
rect 14599 1897 14611 1931
rect 14553 1891 14611 1897
rect 14671 2039 14729 2045
rect 14671 2005 14683 2039
rect 14683 2005 14717 2039
rect 14717 2005 14729 2039
rect 14671 1931 14729 2005
rect 14671 1897 14683 1931
rect 14683 1897 14717 1931
rect 14717 1897 14729 1931
rect 14671 1891 14729 1897
rect 14789 2039 14847 2045
rect 14789 2005 14801 2039
rect 14801 2005 14835 2039
rect 14835 2005 14847 2039
rect 14789 1931 14847 2005
rect 14789 1897 14801 1931
rect 14801 1897 14835 1931
rect 14835 1897 14847 1931
rect 14789 1891 14847 1897
rect 14907 2039 14965 2045
rect 14907 2005 14919 2039
rect 14919 2005 14953 2039
rect 14953 2005 14965 2039
rect 14907 1931 14965 2005
rect 14907 1897 14919 1931
rect 14919 1897 14953 1931
rect 14953 1897 14965 1931
rect 14907 1891 14965 1897
rect 15025 2039 15083 2045
rect 15025 2005 15037 2039
rect 15037 2005 15071 2039
rect 15071 2005 15083 2039
rect 15025 1931 15083 2005
rect 15025 1897 15037 1931
rect 15037 1897 15071 1931
rect 15071 1897 15083 1931
rect 15025 1891 15083 1897
rect 15143 2039 15201 2045
rect 15143 2005 15155 2039
rect 15155 2005 15189 2039
rect 15189 2005 15201 2039
rect 15143 1931 15201 2005
rect 15143 1897 15155 1931
rect 15155 1897 15189 1931
rect 15189 1897 15201 1931
rect 15143 1891 15201 1897
rect 15261 2039 15319 2045
rect 15261 2005 15273 2039
rect 15273 2005 15307 2039
rect 15307 2005 15319 2039
rect 15261 1931 15319 2005
rect 15261 1897 15273 1931
rect 15273 1897 15307 1931
rect 15307 1897 15319 1931
rect 15261 1891 15319 1897
rect 15379 2039 15437 2045
rect 15379 2005 15391 2039
rect 15391 2005 15425 2039
rect 15425 2005 15437 2039
rect 15379 1931 15437 2005
rect 15379 1897 15391 1931
rect 15391 1897 15425 1931
rect 15425 1897 15437 1931
rect 15379 1891 15437 1897
rect 15497 2039 15555 2045
rect 15497 2005 15509 2039
rect 15509 2005 15543 2039
rect 15543 2005 15555 2039
rect 15497 1931 15555 2005
rect 15497 1897 15509 1931
rect 15509 1897 15543 1931
rect 15543 1897 15555 1931
rect 15497 1891 15555 1897
rect 15615 2039 15673 2045
rect 15615 2005 15627 2039
rect 15627 2005 15661 2039
rect 15661 2005 15673 2039
rect 15615 1931 15673 2005
rect 15615 1897 15627 1931
rect 15627 1897 15661 1931
rect 15661 1897 15673 1931
rect 15615 1891 15673 1897
rect 15733 2039 15791 2045
rect 15733 2005 15745 2039
rect 15745 2005 15779 2039
rect 15779 2005 15791 2039
rect 15733 1931 15791 2005
rect 15733 1897 15745 1931
rect 15745 1897 15779 1931
rect 15779 1897 15791 1931
rect 15733 1891 15791 1897
rect 15851 2039 15909 2045
rect 15851 2005 15863 2039
rect 15863 2005 15897 2039
rect 15897 2005 15909 2039
rect 15851 1931 15909 2005
rect 15851 1897 15863 1931
rect 15863 1897 15897 1931
rect 15897 1897 15909 1931
rect 15851 1891 15909 1897
rect 15969 2039 16027 2045
rect 15969 2005 15981 2039
rect 15981 2005 16015 2039
rect 16015 2005 16027 2039
rect 15969 1931 16027 2005
rect 15969 1897 15981 1931
rect 15981 1897 16015 1931
rect 16015 1897 16027 1931
rect 15969 1891 16027 1897
rect 16087 2039 16145 2045
rect 16087 2005 16099 2039
rect 16099 2005 16133 2039
rect 16133 2005 16145 2039
rect 16087 1931 16145 2005
rect 16087 1897 16099 1931
rect 16099 1897 16133 1931
rect 16133 1897 16145 1931
rect 16087 1891 16145 1897
rect 16205 2039 16263 2045
rect 16205 2005 16217 2039
rect 16217 2005 16251 2039
rect 16251 2005 16263 2039
rect 16205 1931 16263 2005
rect 16205 1897 16217 1931
rect 16217 1897 16251 1931
rect 16251 1897 16263 1931
rect 16205 1891 16263 1897
rect 16323 2039 16381 2045
rect 16323 2005 16335 2039
rect 16335 2005 16369 2039
rect 16369 2005 16381 2039
rect 16323 1931 16381 2005
rect 16323 1897 16335 1931
rect 16335 1897 16369 1931
rect 16369 1897 16381 1931
rect 16323 1891 16381 1897
rect 16441 2039 16499 2045
rect 16441 2005 16453 2039
rect 16453 2005 16487 2039
rect 16487 2005 16499 2039
rect 16441 1931 16499 2005
rect 16441 1897 16453 1931
rect 16453 1897 16487 1931
rect 16487 1897 16499 1931
rect 16441 1891 16499 1897
rect 16559 2039 16617 2045
rect 16559 2005 16571 2039
rect 16571 2005 16605 2039
rect 16605 2005 16617 2039
rect 16559 1931 16617 2005
rect 16559 1897 16571 1931
rect 16571 1897 16605 1931
rect 16605 1897 16617 1931
rect 16559 1891 16617 1897
rect 16677 2039 16735 2045
rect 16677 2005 16689 2039
rect 16689 2005 16723 2039
rect 16723 2005 16735 2039
rect 16677 1931 16735 2005
rect 16677 1897 16689 1931
rect 16689 1897 16723 1931
rect 16723 1897 16735 1931
rect 16677 1891 16735 1897
rect 16795 2039 16853 2045
rect 16795 2005 16807 2039
rect 16807 2005 16841 2039
rect 16841 2005 16853 2039
rect 16795 1931 16853 2005
rect 16795 1897 16807 1931
rect 16807 1897 16841 1931
rect 16841 1897 16853 1931
rect 16795 1891 16853 1897
rect 16913 2039 16971 2045
rect 16913 2005 16925 2039
rect 16925 2005 16959 2039
rect 16959 2005 16971 2039
rect 16913 1931 16971 2005
rect 16913 1897 16925 1931
rect 16925 1897 16959 1931
rect 16959 1897 16971 1931
rect 16913 1891 16971 1897
rect 17031 2039 17089 2045
rect 17031 2005 17043 2039
rect 17043 2005 17077 2039
rect 17077 2005 17089 2039
rect 17031 1931 17089 2005
rect 17031 1897 17043 1931
rect 17043 1897 17077 1931
rect 17077 1897 17089 1931
rect 17031 1891 17089 1897
rect 17149 2039 17207 2045
rect 17149 2005 17161 2039
rect 17161 2005 17195 2039
rect 17195 2005 17207 2039
rect 17149 1931 17207 2005
rect 17149 1897 17161 1931
rect 17161 1897 17195 1931
rect 17195 1897 17207 1931
rect 17149 1891 17207 1897
rect 17267 2039 17325 2045
rect 17267 2005 17279 2039
rect 17279 2005 17313 2039
rect 17313 2005 17325 2039
rect 17267 1931 17325 2005
rect 17267 1897 17279 1931
rect 17279 1897 17313 1931
rect 17313 1897 17325 1931
rect 17267 1891 17325 1897
rect 17385 2039 17443 2045
rect 17385 2005 17397 2039
rect 17397 2005 17431 2039
rect 17431 2005 17443 2039
rect 17385 1931 17443 2005
rect 17385 1897 17397 1931
rect 17397 1897 17431 1931
rect 17431 1897 17443 1931
rect 17385 1891 17443 1897
rect 17503 2039 17561 2045
rect 17503 2005 17515 2039
rect 17515 2005 17549 2039
rect 17549 2005 17561 2039
rect 17503 1931 17561 2005
rect 17503 1897 17515 1931
rect 17515 1897 17549 1931
rect 17549 1897 17561 1931
rect 17503 1891 17561 1897
rect 17621 2039 17679 2045
rect 17621 2005 17633 2039
rect 17633 2005 17667 2039
rect 17667 2005 17679 2039
rect 17621 1931 17679 2005
rect 17621 1897 17633 1931
rect 17633 1897 17667 1931
rect 17667 1897 17679 1931
rect 17621 1891 17679 1897
rect 17739 2039 17797 2045
rect 17739 2005 17751 2039
rect 17751 2005 17785 2039
rect 17785 2005 17797 2039
rect 17739 1931 17797 2005
rect 17739 1897 17751 1931
rect 17751 1897 17785 1931
rect 17785 1897 17797 1931
rect 17739 1891 17797 1897
rect 17857 2039 17915 2045
rect 17857 2005 17869 2039
rect 17869 2005 17903 2039
rect 17903 2005 17915 2039
rect 17857 1931 17915 2005
rect 17857 1897 17869 1931
rect 17869 1897 17903 1931
rect 17903 1897 17915 1931
rect 17857 1891 17915 1897
rect 17975 2039 18033 2045
rect 17975 2005 17987 2039
rect 17987 2005 18021 2039
rect 18021 2005 18033 2039
rect 17975 1931 18033 2005
rect 17975 1897 17987 1931
rect 17987 1897 18021 1931
rect 18021 1897 18033 1931
rect 17975 1891 18033 1897
rect 18093 2039 18151 2045
rect 18093 2005 18105 2039
rect 18105 2005 18139 2039
rect 18139 2005 18151 2039
rect 18093 1931 18151 2005
rect 18093 1897 18105 1931
rect 18105 1897 18139 1931
rect 18139 1897 18151 1931
rect 18093 1891 18151 1897
rect 18211 2039 18269 2045
rect 18211 2005 18223 2039
rect 18223 2005 18257 2039
rect 18257 2005 18269 2039
rect 18211 1931 18269 2005
rect 18211 1897 18223 1931
rect 18223 1897 18257 1931
rect 18257 1897 18269 1931
rect 18211 1891 18269 1897
rect 18329 2039 18387 2045
rect 18329 2005 18341 2039
rect 18341 2005 18375 2039
rect 18375 2005 18387 2039
rect 18329 1931 18387 2005
rect 18329 1897 18341 1931
rect 18341 1897 18375 1931
rect 18375 1897 18387 1931
rect 18329 1891 18387 1897
rect 18447 2039 18505 2045
rect 18447 2005 18459 2039
rect 18459 2005 18493 2039
rect 18493 2005 18505 2039
rect 18447 1931 18505 2005
rect 18447 1897 18459 1931
rect 18459 1897 18493 1931
rect 18493 1897 18505 1931
rect 18447 1891 18505 1897
rect 18565 2039 18623 2045
rect 18565 2005 18577 2039
rect 18577 2005 18611 2039
rect 18611 2005 18623 2039
rect 18565 1931 18623 2005
rect 18565 1897 18577 1931
rect 18577 1897 18611 1931
rect 18611 1897 18623 1931
rect 18565 1891 18623 1897
rect 18683 2039 18741 2045
rect 18683 2005 18695 2039
rect 18695 2005 18729 2039
rect 18729 2005 18741 2039
rect 18683 1931 18741 2005
rect 18683 1897 18695 1931
rect 18695 1897 18729 1931
rect 18729 1897 18741 1931
rect 18683 1891 18741 1897
rect 18801 2039 18859 2045
rect 18801 2005 18813 2039
rect 18813 2005 18847 2039
rect 18847 2005 18859 2039
rect 18801 1931 18859 2005
rect 18801 1897 18813 1931
rect 18813 1897 18847 1931
rect 18847 1897 18859 1931
rect 18801 1891 18859 1897
rect 18919 2039 18977 2045
rect 18919 2005 18931 2039
rect 18931 2005 18965 2039
rect 18965 2005 18977 2039
rect 18919 1931 18977 2005
rect 18919 1897 18931 1931
rect 18931 1897 18965 1931
rect 18965 1897 18977 1931
rect 18919 1891 18977 1897
rect 19037 2039 19095 2045
rect 19037 2005 19049 2039
rect 19049 2005 19083 2039
rect 19083 2005 19095 2039
rect 19037 1931 19095 2005
rect 19037 1897 19049 1931
rect 19049 1897 19083 1931
rect 19083 1897 19095 1931
rect 19037 1891 19095 1897
rect 19155 2039 19213 2045
rect 19155 2005 19167 2039
rect 19167 2005 19201 2039
rect 19201 2005 19213 2039
rect 19155 1931 19213 2005
rect 19155 1897 19167 1931
rect 19167 1897 19201 1931
rect 19201 1897 19213 1931
rect 19155 1891 19213 1897
rect 19273 2039 19331 2045
rect 19273 2005 19285 2039
rect 19285 2005 19319 2039
rect 19319 2005 19331 2039
rect 19273 1931 19331 2005
rect 19273 1897 19285 1931
rect 19285 1897 19319 1931
rect 19319 1897 19331 1931
rect 19273 1891 19331 1897
rect 19391 2039 19449 2045
rect 19391 2005 19403 2039
rect 19403 2005 19437 2039
rect 19437 2005 19449 2039
rect 19391 1931 19449 2005
rect 19391 1897 19403 1931
rect 19403 1897 19437 1931
rect 19437 1897 19449 1931
rect 19391 1891 19449 1897
rect 19509 2039 19567 2045
rect 19509 2005 19521 2039
rect 19521 2005 19555 2039
rect 19555 2005 19567 2039
rect 19509 1931 19567 2005
rect 19509 1897 19521 1931
rect 19521 1897 19555 1931
rect 19555 1897 19567 1931
rect 19509 1891 19567 1897
rect 19627 2039 19685 2045
rect 19627 2005 19639 2039
rect 19639 2005 19673 2039
rect 19673 2005 19685 2039
rect 19627 1931 19685 2005
rect 19627 1897 19639 1931
rect 19639 1897 19673 1931
rect 19673 1897 19685 1931
rect 19627 1891 19685 1897
rect 19745 2039 19803 2045
rect 19745 2005 19757 2039
rect 19757 2005 19791 2039
rect 19791 2005 19803 2039
rect 19745 1931 19803 2005
rect 19745 1897 19757 1931
rect 19757 1897 19791 1931
rect 19791 1897 19803 1931
rect 19745 1891 19803 1897
rect 19863 2039 19921 2045
rect 19863 2005 19875 2039
rect 19875 2005 19909 2039
rect 19909 2005 19921 2039
rect 19863 1931 19921 2005
rect 19863 1897 19875 1931
rect 19875 1897 19909 1931
rect 19909 1897 19921 1931
rect 19863 1891 19921 1897
rect 19981 2039 20039 2045
rect 19981 2005 19993 2039
rect 19993 2005 20027 2039
rect 20027 2005 20039 2039
rect 19981 1931 20039 2005
rect 19981 1897 19993 1931
rect 19993 1897 20027 1931
rect 20027 1897 20039 1931
rect 19981 1891 20039 1897
rect 20099 2039 20157 2045
rect 20099 2005 20111 2039
rect 20111 2005 20145 2039
rect 20145 2005 20157 2039
rect 20099 1931 20157 2005
rect 20099 1897 20111 1931
rect 20111 1897 20145 1931
rect 20145 1897 20157 1931
rect 20099 1891 20157 1897
rect 20217 2039 20275 2045
rect 20217 2005 20229 2039
rect 20229 2005 20263 2039
rect 20263 2005 20275 2039
rect 20217 1931 20275 2005
rect 20217 1897 20229 1931
rect 20229 1897 20263 1931
rect 20263 1897 20275 1931
rect 20217 1891 20275 1897
rect 20335 2039 20393 2045
rect 20335 2005 20347 2039
rect 20347 2005 20381 2039
rect 20381 2005 20393 2039
rect 20335 1931 20393 2005
rect 20335 1897 20347 1931
rect 20347 1897 20381 1931
rect 20381 1897 20393 1931
rect 20335 1891 20393 1897
rect 20453 2039 20511 2045
rect 20453 2005 20465 2039
rect 20465 2005 20499 2039
rect 20499 2005 20511 2039
rect 20453 1931 20511 2005
rect 20453 1897 20465 1931
rect 20465 1897 20499 1931
rect 20499 1897 20511 1931
rect 20453 1891 20511 1897
rect 20571 2039 20629 2045
rect 20571 2005 20583 2039
rect 20583 2005 20617 2039
rect 20617 2005 20629 2039
rect 20571 1931 20629 2005
rect 20571 1897 20583 1931
rect 20583 1897 20617 1931
rect 20617 1897 20629 1931
rect 20571 1891 20629 1897
rect 20689 2039 20747 2045
rect 20689 2005 20701 2039
rect 20701 2005 20735 2039
rect 20735 2005 20747 2039
rect 20689 1931 20747 2005
rect 20689 1897 20701 1931
rect 20701 1897 20735 1931
rect 20735 1897 20747 1931
rect 20689 1891 20747 1897
rect 20807 2039 20865 2045
rect 20807 2005 20819 2039
rect 20819 2005 20853 2039
rect 20853 2005 20865 2039
rect 20807 1931 20865 2005
rect 20807 1897 20819 1931
rect 20819 1897 20853 1931
rect 20853 1897 20865 1931
rect 20807 1891 20865 1897
rect 20925 2039 20983 2045
rect 20925 2005 20937 2039
rect 20937 2005 20971 2039
rect 20971 2005 20983 2039
rect 20925 1931 20983 2005
rect 20925 1897 20937 1931
rect 20937 1897 20971 1931
rect 20971 1897 20983 1931
rect 20925 1891 20983 1897
rect 21043 2039 21101 2045
rect 21043 2005 21055 2039
rect 21055 2005 21089 2039
rect 21089 2005 21101 2039
rect 21043 1931 21101 2005
rect 21043 1897 21055 1931
rect 21055 1897 21089 1931
rect 21089 1897 21101 1931
rect 21043 1891 21101 1897
rect 21161 2039 21219 2045
rect 21161 2005 21173 2039
rect 21173 2005 21207 2039
rect 21207 2005 21219 2039
rect 21161 1931 21219 2005
rect 21161 1897 21173 1931
rect 21173 1897 21207 1931
rect 21207 1897 21219 1931
rect 21161 1891 21219 1897
rect 21279 2039 21337 2045
rect 21279 2005 21291 2039
rect 21291 2005 21325 2039
rect 21325 2005 21337 2039
rect 21279 1931 21337 2005
rect 21279 1897 21291 1931
rect 21291 1897 21325 1931
rect 21325 1897 21337 1931
rect 21279 1891 21337 1897
rect 1337 -296 1395 -142
rect 1455 -148 1513 -142
rect 1455 -182 1467 -148
rect 1467 -182 1501 -148
rect 1501 -182 1513 -148
rect 1455 -256 1513 -182
rect 1455 -290 1467 -256
rect 1467 -290 1501 -256
rect 1501 -290 1513 -256
rect 1455 -296 1513 -290
rect 1573 -148 1631 -142
rect 1573 -182 1585 -148
rect 1585 -182 1619 -148
rect 1619 -182 1631 -148
rect 1573 -256 1631 -182
rect 1573 -290 1585 -256
rect 1585 -290 1619 -256
rect 1619 -290 1631 -256
rect 1573 -296 1631 -290
rect 1691 -148 1749 -142
rect 1691 -182 1703 -148
rect 1703 -182 1737 -148
rect 1737 -182 1749 -148
rect 1691 -256 1749 -182
rect 1691 -290 1703 -256
rect 1703 -290 1737 -256
rect 1737 -290 1749 -256
rect 1691 -296 1749 -290
rect 1809 -148 1867 -142
rect 1809 -182 1821 -148
rect 1821 -182 1855 -148
rect 1855 -182 1867 -148
rect 1809 -256 1867 -182
rect 1809 -290 1821 -256
rect 1821 -290 1855 -256
rect 1855 -290 1867 -256
rect 1809 -296 1867 -290
rect 1927 -148 1985 -142
rect 1927 -182 1939 -148
rect 1939 -182 1973 -148
rect 1973 -182 1985 -148
rect 1927 -256 1985 -182
rect 1927 -290 1939 -256
rect 1939 -290 1973 -256
rect 1973 -290 1985 -256
rect 1927 -296 1985 -290
rect 2045 -148 2103 -142
rect 2045 -182 2057 -148
rect 2057 -182 2091 -148
rect 2091 -182 2103 -148
rect 2045 -256 2103 -182
rect 2045 -290 2057 -256
rect 2057 -290 2091 -256
rect 2091 -290 2103 -256
rect 2045 -296 2103 -290
rect 2163 -148 2221 -142
rect 2163 -182 2175 -148
rect 2175 -182 2209 -148
rect 2209 -182 2221 -148
rect 2163 -256 2221 -182
rect 2163 -290 2175 -256
rect 2175 -290 2209 -256
rect 2209 -290 2221 -256
rect 2163 -296 2221 -290
rect 2281 -148 2339 -142
rect 2281 -182 2293 -148
rect 2293 -182 2327 -148
rect 2327 -182 2339 -148
rect 2281 -256 2339 -182
rect 2281 -290 2293 -256
rect 2293 -290 2327 -256
rect 2327 -290 2339 -256
rect 2281 -296 2339 -290
rect 2399 -148 2457 -142
rect 2399 -182 2411 -148
rect 2411 -182 2445 -148
rect 2445 -182 2457 -148
rect 2399 -256 2457 -182
rect 2399 -290 2411 -256
rect 2411 -290 2445 -256
rect 2445 -290 2457 -256
rect 2399 -296 2457 -290
rect 2517 -148 2575 -142
rect 2517 -182 2529 -148
rect 2529 -182 2563 -148
rect 2563 -182 2575 -148
rect 2517 -256 2575 -182
rect 2517 -290 2529 -256
rect 2529 -290 2563 -256
rect 2563 -290 2575 -256
rect 2517 -296 2575 -290
rect 2635 -148 2693 -142
rect 2635 -182 2647 -148
rect 2647 -182 2681 -148
rect 2681 -182 2693 -148
rect 2635 -256 2693 -182
rect 2635 -290 2647 -256
rect 2647 -290 2681 -256
rect 2681 -290 2693 -256
rect 2635 -296 2693 -290
rect 2753 -148 2811 -142
rect 2753 -182 2765 -148
rect 2765 -182 2799 -148
rect 2799 -182 2811 -148
rect 2753 -256 2811 -182
rect 2753 -290 2765 -256
rect 2765 -290 2799 -256
rect 2799 -290 2811 -256
rect 2753 -296 2811 -290
rect 2871 -148 2929 -142
rect 2871 -182 2883 -148
rect 2883 -182 2917 -148
rect 2917 -182 2929 -148
rect 2871 -256 2929 -182
rect 2871 -290 2883 -256
rect 2883 -290 2917 -256
rect 2917 -290 2929 -256
rect 2871 -296 2929 -290
rect 2989 -148 3047 -142
rect 2989 -182 3001 -148
rect 3001 -182 3035 -148
rect 3035 -182 3047 -148
rect 2989 -256 3047 -182
rect 2989 -290 3001 -256
rect 3001 -290 3035 -256
rect 3035 -290 3047 -256
rect 2989 -296 3047 -290
rect 3107 -148 3165 -142
rect 3107 -182 3119 -148
rect 3119 -182 3153 -148
rect 3153 -182 3165 -148
rect 3107 -256 3165 -182
rect 3107 -290 3119 -256
rect 3119 -290 3153 -256
rect 3153 -290 3165 -256
rect 3107 -296 3165 -290
rect 3225 -148 3283 -142
rect 3225 -182 3237 -148
rect 3237 -182 3271 -148
rect 3271 -182 3283 -148
rect 3225 -256 3283 -182
rect 3225 -290 3237 -256
rect 3237 -290 3271 -256
rect 3271 -290 3283 -256
rect 3225 -296 3283 -290
rect 3343 -148 3401 -142
rect 3343 -182 3355 -148
rect 3355 -182 3389 -148
rect 3389 -182 3401 -148
rect 3343 -256 3401 -182
rect 3343 -290 3355 -256
rect 3355 -290 3389 -256
rect 3389 -290 3401 -256
rect 3343 -296 3401 -290
rect 3461 -148 3519 -142
rect 3461 -182 3473 -148
rect 3473 -182 3507 -148
rect 3507 -182 3519 -148
rect 3461 -256 3519 -182
rect 3461 -290 3473 -256
rect 3473 -290 3507 -256
rect 3507 -290 3519 -256
rect 3461 -296 3519 -290
rect 3579 -148 3637 -142
rect 3579 -182 3591 -148
rect 3591 -182 3625 -148
rect 3625 -182 3637 -148
rect 3579 -256 3637 -182
rect 3579 -290 3591 -256
rect 3591 -290 3625 -256
rect 3625 -290 3637 -256
rect 3579 -296 3637 -290
rect 3697 -148 3755 -142
rect 3697 -182 3709 -148
rect 3709 -182 3743 -148
rect 3743 -182 3755 -148
rect 3697 -256 3755 -182
rect 3697 -290 3709 -256
rect 3709 -290 3743 -256
rect 3743 -290 3755 -256
rect 3697 -296 3755 -290
rect 3815 -148 3873 -142
rect 3815 -182 3827 -148
rect 3827 -182 3861 -148
rect 3861 -182 3873 -148
rect 3815 -256 3873 -182
rect 3815 -290 3827 -256
rect 3827 -290 3861 -256
rect 3861 -290 3873 -256
rect 3815 -296 3873 -290
rect 3933 -148 3991 -142
rect 3933 -182 3945 -148
rect 3945 -182 3979 -148
rect 3979 -182 3991 -148
rect 3933 -256 3991 -182
rect 3933 -290 3945 -256
rect 3945 -290 3979 -256
rect 3979 -290 3991 -256
rect 3933 -296 3991 -290
rect 4051 -148 4109 -142
rect 4051 -182 4063 -148
rect 4063 -182 4097 -148
rect 4097 -182 4109 -148
rect 4051 -256 4109 -182
rect 4051 -290 4063 -256
rect 4063 -290 4097 -256
rect 4097 -290 4109 -256
rect 4051 -296 4109 -290
rect 4169 -148 4227 -142
rect 4169 -182 4181 -148
rect 4181 -182 4215 -148
rect 4215 -182 4227 -148
rect 4169 -256 4227 -182
rect 4169 -290 4181 -256
rect 4181 -290 4215 -256
rect 4215 -290 4227 -256
rect 4169 -296 4227 -290
rect 4287 -148 4345 -142
rect 4287 -182 4299 -148
rect 4299 -182 4333 -148
rect 4333 -182 4345 -148
rect 4287 -256 4345 -182
rect 4287 -290 4299 -256
rect 4299 -290 4333 -256
rect 4333 -290 4345 -256
rect 4287 -296 4345 -290
rect 4405 -148 4463 -142
rect 4405 -182 4417 -148
rect 4417 -182 4451 -148
rect 4451 -182 4463 -148
rect 4405 -256 4463 -182
rect 4405 -290 4417 -256
rect 4417 -290 4451 -256
rect 4451 -290 4463 -256
rect 4405 -296 4463 -290
rect 4523 -148 4581 -142
rect 4523 -182 4535 -148
rect 4535 -182 4569 -148
rect 4569 -182 4581 -148
rect 4523 -256 4581 -182
rect 4523 -290 4535 -256
rect 4535 -290 4569 -256
rect 4569 -290 4581 -256
rect 4523 -296 4581 -290
rect 4641 -148 4699 -142
rect 4641 -182 4653 -148
rect 4653 -182 4687 -148
rect 4687 -182 4699 -148
rect 4641 -256 4699 -182
rect 4641 -290 4653 -256
rect 4653 -290 4687 -256
rect 4687 -290 4699 -256
rect 4641 -296 4699 -290
rect 4759 -148 4817 -142
rect 4759 -182 4771 -148
rect 4771 -182 4805 -148
rect 4805 -182 4817 -148
rect 4759 -256 4817 -182
rect 4759 -290 4771 -256
rect 4771 -290 4805 -256
rect 4805 -290 4817 -256
rect 4759 -296 4817 -290
rect 4877 -148 4935 -142
rect 4877 -182 4889 -148
rect 4889 -182 4923 -148
rect 4923 -182 4935 -148
rect 4877 -256 4935 -182
rect 4877 -290 4889 -256
rect 4889 -290 4923 -256
rect 4923 -290 4935 -256
rect 4877 -296 4935 -290
rect 4995 -148 5053 -142
rect 4995 -182 5007 -148
rect 5007 -182 5041 -148
rect 5041 -182 5053 -148
rect 4995 -256 5053 -182
rect 4995 -290 5007 -256
rect 5007 -290 5041 -256
rect 5041 -290 5053 -256
rect 4995 -296 5053 -290
rect 5113 -148 5171 -142
rect 5113 -182 5125 -148
rect 5125 -182 5159 -148
rect 5159 -182 5171 -148
rect 5113 -256 5171 -182
rect 5113 -290 5125 -256
rect 5125 -290 5159 -256
rect 5159 -290 5171 -256
rect 5113 -296 5171 -290
rect 5231 -148 5289 -142
rect 5231 -182 5243 -148
rect 5243 -182 5277 -148
rect 5277 -182 5289 -148
rect 5231 -256 5289 -182
rect 5231 -290 5243 -256
rect 5243 -290 5277 -256
rect 5277 -290 5289 -256
rect 5231 -296 5289 -290
rect 5349 -148 5407 -142
rect 5349 -182 5361 -148
rect 5361 -182 5395 -148
rect 5395 -182 5407 -148
rect 5349 -256 5407 -182
rect 5349 -290 5361 -256
rect 5361 -290 5395 -256
rect 5395 -290 5407 -256
rect 5349 -296 5407 -290
rect 5467 -148 5525 -142
rect 5467 -182 5479 -148
rect 5479 -182 5513 -148
rect 5513 -182 5525 -148
rect 5467 -256 5525 -182
rect 5467 -290 5479 -256
rect 5479 -290 5513 -256
rect 5513 -290 5525 -256
rect 5467 -296 5525 -290
rect 5585 -148 5643 -142
rect 5585 -182 5597 -148
rect 5597 -182 5631 -148
rect 5631 -182 5643 -148
rect 5585 -256 5643 -182
rect 5585 -290 5597 -256
rect 5597 -290 5631 -256
rect 5631 -290 5643 -256
rect 5585 -296 5643 -290
rect 5703 -148 5761 -142
rect 5703 -182 5715 -148
rect 5715 -182 5749 -148
rect 5749 -182 5761 -148
rect 5703 -256 5761 -182
rect 5703 -290 5715 -256
rect 5715 -290 5749 -256
rect 5749 -290 5761 -256
rect 5703 -296 5761 -290
rect 5821 -148 5879 -142
rect 5821 -182 5833 -148
rect 5833 -182 5867 -148
rect 5867 -182 5879 -148
rect 5821 -256 5879 -182
rect 5821 -290 5833 -256
rect 5833 -290 5867 -256
rect 5867 -290 5879 -256
rect 5821 -296 5879 -290
rect 5939 -148 5997 -142
rect 5939 -182 5951 -148
rect 5951 -182 5985 -148
rect 5985 -182 5997 -148
rect 5939 -256 5997 -182
rect 5939 -290 5951 -256
rect 5951 -290 5985 -256
rect 5985 -290 5997 -256
rect 5939 -296 5997 -290
rect 6057 -148 6115 -142
rect 6057 -182 6069 -148
rect 6069 -182 6103 -148
rect 6103 -182 6115 -148
rect 6057 -256 6115 -182
rect 6057 -290 6069 -256
rect 6069 -290 6103 -256
rect 6103 -290 6115 -256
rect 6057 -296 6115 -290
rect 6175 -148 6233 -142
rect 6175 -182 6187 -148
rect 6187 -182 6221 -148
rect 6221 -182 6233 -148
rect 6175 -256 6233 -182
rect 6175 -290 6187 -256
rect 6187 -290 6221 -256
rect 6221 -290 6233 -256
rect 6175 -296 6233 -290
rect 6293 -148 6351 -142
rect 6293 -182 6305 -148
rect 6305 -182 6339 -148
rect 6339 -182 6351 -148
rect 6293 -256 6351 -182
rect 6293 -290 6305 -256
rect 6305 -290 6339 -256
rect 6339 -290 6351 -256
rect 6293 -296 6351 -290
rect 6411 -148 6469 -142
rect 6411 -182 6423 -148
rect 6423 -182 6457 -148
rect 6457 -182 6469 -148
rect 6411 -256 6469 -182
rect 6411 -290 6423 -256
rect 6423 -290 6457 -256
rect 6457 -290 6469 -256
rect 6411 -296 6469 -290
rect 6529 -148 6587 -142
rect 6529 -182 6541 -148
rect 6541 -182 6575 -148
rect 6575 -182 6587 -148
rect 6529 -256 6587 -182
rect 6529 -290 6541 -256
rect 6541 -290 6575 -256
rect 6575 -290 6587 -256
rect 6529 -296 6587 -290
rect 6647 -148 6705 -142
rect 6647 -182 6659 -148
rect 6659 -182 6693 -148
rect 6693 -182 6705 -148
rect 6647 -256 6705 -182
rect 6647 -290 6659 -256
rect 6659 -290 6693 -256
rect 6693 -290 6705 -256
rect 6647 -296 6705 -290
rect 6765 -148 6823 -142
rect 6765 -182 6777 -148
rect 6777 -182 6811 -148
rect 6811 -182 6823 -148
rect 6765 -256 6823 -182
rect 6765 -290 6777 -256
rect 6777 -290 6811 -256
rect 6811 -290 6823 -256
rect 6765 -296 6823 -290
rect 6883 -148 6941 -142
rect 6883 -182 6895 -148
rect 6895 -182 6929 -148
rect 6929 -182 6941 -148
rect 6883 -256 6941 -182
rect 6883 -290 6895 -256
rect 6895 -290 6929 -256
rect 6929 -290 6941 -256
rect 6883 -296 6941 -290
rect 7001 -148 7059 -142
rect 7001 -182 7013 -148
rect 7013 -182 7047 -148
rect 7047 -182 7059 -148
rect 7001 -256 7059 -182
rect 7001 -290 7013 -256
rect 7013 -290 7047 -256
rect 7047 -290 7059 -256
rect 7001 -296 7059 -290
rect 7119 -148 7177 -142
rect 7119 -182 7131 -148
rect 7131 -182 7165 -148
rect 7165 -182 7177 -148
rect 7119 -256 7177 -182
rect 7119 -290 7131 -256
rect 7131 -290 7165 -256
rect 7165 -290 7177 -256
rect 7119 -296 7177 -290
rect 1337 -1916 1395 -1910
rect 1337 -1950 1349 -1916
rect 1349 -1950 1383 -1916
rect 1383 -1950 1395 -1916
rect 1337 -2024 1395 -1950
rect 1337 -2058 1349 -2024
rect 1349 -2058 1383 -2024
rect 1383 -2058 1395 -2024
rect 1337 -2064 1395 -2058
rect 1455 -1916 1513 -1910
rect 1455 -1950 1467 -1916
rect 1467 -1950 1501 -1916
rect 1501 -1950 1513 -1916
rect 1455 -2024 1513 -1950
rect 1455 -2058 1467 -2024
rect 1467 -2058 1501 -2024
rect 1501 -2058 1513 -2024
rect 1455 -2064 1513 -2058
rect 1573 -1916 1631 -1910
rect 1573 -1950 1585 -1916
rect 1585 -1950 1619 -1916
rect 1619 -1950 1631 -1916
rect 1573 -2024 1631 -1950
rect 1573 -2058 1585 -2024
rect 1585 -2058 1619 -2024
rect 1619 -2058 1631 -2024
rect 1573 -2064 1631 -2058
rect 1691 -1916 1749 -1910
rect 1691 -1950 1703 -1916
rect 1703 -1950 1737 -1916
rect 1737 -1950 1749 -1916
rect 1691 -2024 1749 -1950
rect 1691 -2058 1703 -2024
rect 1703 -2058 1737 -2024
rect 1737 -2058 1749 -2024
rect 1691 -2064 1749 -2058
rect 1809 -1916 1867 -1910
rect 1809 -1950 1821 -1916
rect 1821 -1950 1855 -1916
rect 1855 -1950 1867 -1916
rect 1809 -2024 1867 -1950
rect 1809 -2058 1821 -2024
rect 1821 -2058 1855 -2024
rect 1855 -2058 1867 -2024
rect 1809 -2064 1867 -2058
rect 1927 -1916 1985 -1910
rect 1927 -1950 1939 -1916
rect 1939 -1950 1973 -1916
rect 1973 -1950 1985 -1916
rect 1927 -2024 1985 -1950
rect 1927 -2058 1939 -2024
rect 1939 -2058 1973 -2024
rect 1973 -2058 1985 -2024
rect 1927 -2064 1985 -2058
rect 2045 -1916 2103 -1910
rect 2045 -1950 2057 -1916
rect 2057 -1950 2091 -1916
rect 2091 -1950 2103 -1916
rect 2045 -2024 2103 -1950
rect 2045 -2058 2057 -2024
rect 2057 -2058 2091 -2024
rect 2091 -2058 2103 -2024
rect 2045 -2064 2103 -2058
rect 2163 -1916 2221 -1910
rect 2163 -1950 2175 -1916
rect 2175 -1950 2209 -1916
rect 2209 -1950 2221 -1916
rect 2163 -2024 2221 -1950
rect 2163 -2058 2175 -2024
rect 2175 -2058 2209 -2024
rect 2209 -2058 2221 -2024
rect 2163 -2064 2221 -2058
rect 2281 -1916 2339 -1910
rect 2281 -1950 2293 -1916
rect 2293 -1950 2327 -1916
rect 2327 -1950 2339 -1916
rect 2281 -2024 2339 -1950
rect 2281 -2058 2293 -2024
rect 2293 -2058 2327 -2024
rect 2327 -2058 2339 -2024
rect 2281 -2064 2339 -2058
rect 2399 -1916 2457 -1910
rect 2399 -1950 2411 -1916
rect 2411 -1950 2445 -1916
rect 2445 -1950 2457 -1916
rect 2399 -2024 2457 -1950
rect 2399 -2058 2411 -2024
rect 2411 -2058 2445 -2024
rect 2445 -2058 2457 -2024
rect 2399 -2064 2457 -2058
rect 2517 -1916 2575 -1910
rect 2517 -1950 2529 -1916
rect 2529 -1950 2563 -1916
rect 2563 -1950 2575 -1916
rect 2517 -2024 2575 -1950
rect 2517 -2058 2529 -2024
rect 2529 -2058 2563 -2024
rect 2563 -2058 2575 -2024
rect 2517 -2064 2575 -2058
rect 2635 -1916 2693 -1910
rect 2635 -1950 2647 -1916
rect 2647 -1950 2681 -1916
rect 2681 -1950 2693 -1916
rect 2635 -2024 2693 -1950
rect 2635 -2058 2647 -2024
rect 2647 -2058 2681 -2024
rect 2681 -2058 2693 -2024
rect 2635 -2064 2693 -2058
rect 2753 -1916 2811 -1910
rect 2753 -1950 2765 -1916
rect 2765 -1950 2799 -1916
rect 2799 -1950 2811 -1916
rect 2753 -2024 2811 -1950
rect 2753 -2058 2765 -2024
rect 2765 -2058 2799 -2024
rect 2799 -2058 2811 -2024
rect 2753 -2064 2811 -2058
rect 2871 -1916 2929 -1910
rect 2871 -1950 2883 -1916
rect 2883 -1950 2917 -1916
rect 2917 -1950 2929 -1916
rect 2871 -2024 2929 -1950
rect 2871 -2058 2883 -2024
rect 2883 -2058 2917 -2024
rect 2917 -2058 2929 -2024
rect 2871 -2064 2929 -2058
rect 2989 -1916 3047 -1910
rect 2989 -1950 3001 -1916
rect 3001 -1950 3035 -1916
rect 3035 -1950 3047 -1916
rect 2989 -2024 3047 -1950
rect 2989 -2058 3001 -2024
rect 3001 -2058 3035 -2024
rect 3035 -2058 3047 -2024
rect 2989 -2064 3047 -2058
rect 3107 -1916 3165 -1910
rect 3107 -1950 3119 -1916
rect 3119 -1950 3153 -1916
rect 3153 -1950 3165 -1916
rect 3107 -2024 3165 -1950
rect 3107 -2058 3119 -2024
rect 3119 -2058 3153 -2024
rect 3153 -2058 3165 -2024
rect 3107 -2064 3165 -2058
rect 3225 -1916 3283 -1910
rect 3225 -1950 3237 -1916
rect 3237 -1950 3271 -1916
rect 3271 -1950 3283 -1916
rect 3225 -2024 3283 -1950
rect 3225 -2058 3237 -2024
rect 3237 -2058 3271 -2024
rect 3271 -2058 3283 -2024
rect 3225 -2064 3283 -2058
rect 3343 -1916 3401 -1910
rect 3343 -1950 3355 -1916
rect 3355 -1950 3389 -1916
rect 3389 -1950 3401 -1916
rect 3343 -2024 3401 -1950
rect 3343 -2058 3355 -2024
rect 3355 -2058 3389 -2024
rect 3389 -2058 3401 -2024
rect 3343 -2064 3401 -2058
rect 3461 -1916 3519 -1910
rect 3461 -1950 3473 -1916
rect 3473 -1950 3507 -1916
rect 3507 -1950 3519 -1916
rect 3461 -2024 3519 -1950
rect 3461 -2058 3473 -2024
rect 3473 -2058 3507 -2024
rect 3507 -2058 3519 -2024
rect 3461 -2064 3519 -2058
rect 3579 -1916 3637 -1910
rect 3579 -1950 3591 -1916
rect 3591 -1950 3625 -1916
rect 3625 -1950 3637 -1916
rect 3579 -2024 3637 -1950
rect 3579 -2058 3591 -2024
rect 3591 -2058 3625 -2024
rect 3625 -2058 3637 -2024
rect 3579 -2064 3637 -2058
rect 3697 -1916 3755 -1910
rect 3697 -1950 3709 -1916
rect 3709 -1950 3743 -1916
rect 3743 -1950 3755 -1916
rect 3697 -2024 3755 -1950
rect 3697 -2058 3709 -2024
rect 3709 -2058 3743 -2024
rect 3743 -2058 3755 -2024
rect 3697 -2064 3755 -2058
rect 3815 -1916 3873 -1910
rect 3815 -1950 3827 -1916
rect 3827 -1950 3861 -1916
rect 3861 -1950 3873 -1916
rect 3815 -2024 3873 -1950
rect 3815 -2058 3827 -2024
rect 3827 -2058 3861 -2024
rect 3861 -2058 3873 -2024
rect 3815 -2064 3873 -2058
rect 3933 -1916 3991 -1910
rect 3933 -1950 3945 -1916
rect 3945 -1950 3979 -1916
rect 3979 -1950 3991 -1916
rect 3933 -2024 3991 -1950
rect 3933 -2058 3945 -2024
rect 3945 -2058 3979 -2024
rect 3979 -2058 3991 -2024
rect 3933 -2064 3991 -2058
rect 4051 -1916 4109 -1910
rect 4051 -1950 4063 -1916
rect 4063 -1950 4097 -1916
rect 4097 -1950 4109 -1916
rect 4051 -2024 4109 -1950
rect 4051 -2058 4063 -2024
rect 4063 -2058 4097 -2024
rect 4097 -2058 4109 -2024
rect 4051 -2064 4109 -2058
rect 4169 -1916 4227 -1910
rect 4169 -1950 4181 -1916
rect 4181 -1950 4215 -1916
rect 4215 -1950 4227 -1916
rect 4169 -2024 4227 -1950
rect 4169 -2058 4181 -2024
rect 4181 -2058 4215 -2024
rect 4215 -2058 4227 -2024
rect 4169 -2064 4227 -2058
rect 4287 -1916 4345 -1910
rect 4287 -1950 4299 -1916
rect 4299 -1950 4333 -1916
rect 4333 -1950 4345 -1916
rect 4287 -2024 4345 -1950
rect 4287 -2058 4299 -2024
rect 4299 -2058 4333 -2024
rect 4333 -2058 4345 -2024
rect 4287 -2064 4345 -2058
rect 4405 -1916 4463 -1910
rect 4405 -1950 4417 -1916
rect 4417 -1950 4451 -1916
rect 4451 -1950 4463 -1916
rect 4405 -2024 4463 -1950
rect 4405 -2058 4417 -2024
rect 4417 -2058 4451 -2024
rect 4451 -2058 4463 -2024
rect 4405 -2064 4463 -2058
rect 4523 -1916 4581 -1910
rect 4523 -1950 4535 -1916
rect 4535 -1950 4569 -1916
rect 4569 -1950 4581 -1916
rect 4523 -2024 4581 -1950
rect 4523 -2058 4535 -2024
rect 4535 -2058 4569 -2024
rect 4569 -2058 4581 -2024
rect 4523 -2064 4581 -2058
rect 4641 -1916 4699 -1910
rect 4641 -1950 4653 -1916
rect 4653 -1950 4687 -1916
rect 4687 -1950 4699 -1916
rect 4641 -2024 4699 -1950
rect 4641 -2058 4653 -2024
rect 4653 -2058 4687 -2024
rect 4687 -2058 4699 -2024
rect 4641 -2064 4699 -2058
rect 4759 -1916 4817 -1910
rect 4759 -1950 4771 -1916
rect 4771 -1950 4805 -1916
rect 4805 -1950 4817 -1916
rect 4759 -2024 4817 -1950
rect 4759 -2058 4771 -2024
rect 4771 -2058 4805 -2024
rect 4805 -2058 4817 -2024
rect 4759 -2064 4817 -2058
rect 4877 -1916 4935 -1910
rect 4877 -1950 4889 -1916
rect 4889 -1950 4923 -1916
rect 4923 -1950 4935 -1916
rect 4877 -2024 4935 -1950
rect 4877 -2058 4889 -2024
rect 4889 -2058 4923 -2024
rect 4923 -2058 4935 -2024
rect 4877 -2064 4935 -2058
rect 4995 -1916 5053 -1910
rect 4995 -1950 5007 -1916
rect 5007 -1950 5041 -1916
rect 5041 -1950 5053 -1916
rect 4995 -2024 5053 -1950
rect 4995 -2058 5007 -2024
rect 5007 -2058 5041 -2024
rect 5041 -2058 5053 -2024
rect 4995 -2064 5053 -2058
rect 5113 -1916 5171 -1910
rect 5113 -1950 5125 -1916
rect 5125 -1950 5159 -1916
rect 5159 -1950 5171 -1916
rect 5113 -2024 5171 -1950
rect 5113 -2058 5125 -2024
rect 5125 -2058 5159 -2024
rect 5159 -2058 5171 -2024
rect 5113 -2064 5171 -2058
rect 5231 -1916 5289 -1910
rect 5231 -1950 5243 -1916
rect 5243 -1950 5277 -1916
rect 5277 -1950 5289 -1916
rect 5231 -2024 5289 -1950
rect 5231 -2058 5243 -2024
rect 5243 -2058 5277 -2024
rect 5277 -2058 5289 -2024
rect 5231 -2064 5289 -2058
rect 5349 -1916 5407 -1910
rect 5349 -1950 5361 -1916
rect 5361 -1950 5395 -1916
rect 5395 -1950 5407 -1916
rect 5349 -2024 5407 -1950
rect 5349 -2058 5361 -2024
rect 5361 -2058 5395 -2024
rect 5395 -2058 5407 -2024
rect 5349 -2064 5407 -2058
rect 5467 -1916 5525 -1910
rect 5467 -1950 5479 -1916
rect 5479 -1950 5513 -1916
rect 5513 -1950 5525 -1916
rect 5467 -2024 5525 -1950
rect 5467 -2058 5479 -2024
rect 5479 -2058 5513 -2024
rect 5513 -2058 5525 -2024
rect 5467 -2064 5525 -2058
rect 5585 -1916 5643 -1910
rect 5585 -1950 5597 -1916
rect 5597 -1950 5631 -1916
rect 5631 -1950 5643 -1916
rect 5585 -2024 5643 -1950
rect 5585 -2058 5597 -2024
rect 5597 -2058 5631 -2024
rect 5631 -2058 5643 -2024
rect 5585 -2064 5643 -2058
rect 5703 -1916 5761 -1910
rect 5703 -1950 5715 -1916
rect 5715 -1950 5749 -1916
rect 5749 -1950 5761 -1916
rect 5703 -2024 5761 -1950
rect 5703 -2058 5715 -2024
rect 5715 -2058 5749 -2024
rect 5749 -2058 5761 -2024
rect 5703 -2064 5761 -2058
rect 5821 -1916 5879 -1910
rect 5821 -1950 5833 -1916
rect 5833 -1950 5867 -1916
rect 5867 -1950 5879 -1916
rect 5821 -2024 5879 -1950
rect 5821 -2058 5833 -2024
rect 5833 -2058 5867 -2024
rect 5867 -2058 5879 -2024
rect 5821 -2064 5879 -2058
rect 5939 -1916 5997 -1910
rect 5939 -1950 5951 -1916
rect 5951 -1950 5985 -1916
rect 5985 -1950 5997 -1916
rect 5939 -2024 5997 -1950
rect 5939 -2058 5951 -2024
rect 5951 -2058 5985 -2024
rect 5985 -2058 5997 -2024
rect 5939 -2064 5997 -2058
rect 6057 -1916 6115 -1910
rect 6057 -1950 6069 -1916
rect 6069 -1950 6103 -1916
rect 6103 -1950 6115 -1916
rect 6057 -2024 6115 -1950
rect 6057 -2058 6069 -2024
rect 6069 -2058 6103 -2024
rect 6103 -2058 6115 -2024
rect 6057 -2064 6115 -2058
rect 6175 -1916 6233 -1910
rect 6175 -1950 6187 -1916
rect 6187 -1950 6221 -1916
rect 6221 -1950 6233 -1916
rect 6175 -2024 6233 -1950
rect 6175 -2058 6187 -2024
rect 6187 -2058 6221 -2024
rect 6221 -2058 6233 -2024
rect 6175 -2064 6233 -2058
rect 6293 -1916 6351 -1910
rect 6293 -1950 6305 -1916
rect 6305 -1950 6339 -1916
rect 6339 -1950 6351 -1916
rect 6293 -2024 6351 -1950
rect 6293 -2058 6305 -2024
rect 6305 -2058 6339 -2024
rect 6339 -2058 6351 -2024
rect 6293 -2064 6351 -2058
rect 6411 -1916 6469 -1910
rect 6411 -1950 6423 -1916
rect 6423 -1950 6457 -1916
rect 6457 -1950 6469 -1916
rect 6411 -2024 6469 -1950
rect 6411 -2058 6423 -2024
rect 6423 -2058 6457 -2024
rect 6457 -2058 6469 -2024
rect 6411 -2064 6469 -2058
rect 6529 -1916 6587 -1910
rect 6529 -1950 6541 -1916
rect 6541 -1950 6575 -1916
rect 6575 -1950 6587 -1916
rect 6529 -2024 6587 -1950
rect 6529 -2058 6541 -2024
rect 6541 -2058 6575 -2024
rect 6575 -2058 6587 -2024
rect 6529 -2064 6587 -2058
rect 6647 -1916 6705 -1910
rect 6647 -1950 6659 -1916
rect 6659 -1950 6693 -1916
rect 6693 -1950 6705 -1916
rect 6647 -2024 6705 -1950
rect 6647 -2058 6659 -2024
rect 6659 -2058 6693 -2024
rect 6693 -2058 6705 -2024
rect 6647 -2064 6705 -2058
rect 6765 -1916 6823 -1910
rect 6765 -1950 6777 -1916
rect 6777 -1950 6811 -1916
rect 6811 -1950 6823 -1916
rect 6765 -2024 6823 -1950
rect 6765 -2058 6777 -2024
rect 6777 -2058 6811 -2024
rect 6811 -2058 6823 -2024
rect 6765 -2064 6823 -2058
rect 6883 -1916 6941 -1910
rect 6883 -1950 6895 -1916
rect 6895 -1950 6929 -1916
rect 6929 -1950 6941 -1916
rect 6883 -2024 6941 -1950
rect 6883 -2058 6895 -2024
rect 6895 -2058 6929 -2024
rect 6929 -2058 6941 -2024
rect 6883 -2064 6941 -2058
rect 7001 -1916 7059 -1910
rect 7001 -1950 7013 -1916
rect 7013 -1950 7047 -1916
rect 7047 -1950 7059 -1916
rect 7001 -2024 7059 -1950
rect 7001 -2058 7013 -2024
rect 7013 -2058 7047 -2024
rect 7047 -2058 7059 -2024
rect 7001 -2064 7059 -2058
rect 7119 -1916 7177 -1910
rect 7119 -1950 7131 -1916
rect 7131 -1950 7165 -1916
rect 7165 -1950 7177 -1916
rect 7119 -2024 7177 -1950
rect 7119 -2058 7131 -2024
rect 7131 -2058 7165 -2024
rect 7165 -2058 7177 -2024
rect 7119 -2064 7177 -2058
rect 1337 -3684 1395 -3678
rect 1337 -3718 1349 -3684
rect 1349 -3718 1383 -3684
rect 1383 -3718 1395 -3684
rect 1337 -3792 1395 -3718
rect 1337 -3826 1349 -3792
rect 1349 -3826 1383 -3792
rect 1383 -3826 1395 -3792
rect 1337 -3832 1395 -3826
rect 1455 -3684 1513 -3678
rect 1455 -3718 1467 -3684
rect 1467 -3718 1501 -3684
rect 1501 -3718 1513 -3684
rect 1455 -3792 1513 -3718
rect 1455 -3826 1467 -3792
rect 1467 -3826 1501 -3792
rect 1501 -3826 1513 -3792
rect 1455 -3832 1513 -3826
rect 1573 -3684 1631 -3678
rect 1573 -3718 1585 -3684
rect 1585 -3718 1619 -3684
rect 1619 -3718 1631 -3684
rect 1573 -3792 1631 -3718
rect 1573 -3826 1585 -3792
rect 1585 -3826 1619 -3792
rect 1619 -3826 1631 -3792
rect 1573 -3832 1631 -3826
rect 1691 -3684 1749 -3678
rect 1691 -3718 1703 -3684
rect 1703 -3718 1737 -3684
rect 1737 -3718 1749 -3684
rect 1691 -3792 1749 -3718
rect 1691 -3826 1703 -3792
rect 1703 -3826 1737 -3792
rect 1737 -3826 1749 -3792
rect 1691 -3832 1749 -3826
rect 1809 -3684 1867 -3678
rect 1809 -3718 1821 -3684
rect 1821 -3718 1855 -3684
rect 1855 -3718 1867 -3684
rect 1809 -3792 1867 -3718
rect 1809 -3826 1821 -3792
rect 1821 -3826 1855 -3792
rect 1855 -3826 1867 -3792
rect 1809 -3832 1867 -3826
rect 1927 -3684 1985 -3678
rect 1927 -3718 1939 -3684
rect 1939 -3718 1973 -3684
rect 1973 -3718 1985 -3684
rect 1927 -3792 1985 -3718
rect 1927 -3826 1939 -3792
rect 1939 -3826 1973 -3792
rect 1973 -3826 1985 -3792
rect 1927 -3832 1985 -3826
rect 2045 -3684 2103 -3678
rect 2045 -3718 2057 -3684
rect 2057 -3718 2091 -3684
rect 2091 -3718 2103 -3684
rect 2045 -3792 2103 -3718
rect 2045 -3826 2057 -3792
rect 2057 -3826 2091 -3792
rect 2091 -3826 2103 -3792
rect 2045 -3832 2103 -3826
rect 2163 -3684 2221 -3678
rect 2163 -3718 2175 -3684
rect 2175 -3718 2209 -3684
rect 2209 -3718 2221 -3684
rect 2163 -3792 2221 -3718
rect 2163 -3826 2175 -3792
rect 2175 -3826 2209 -3792
rect 2209 -3826 2221 -3792
rect 2163 -3832 2221 -3826
rect 2281 -3684 2339 -3678
rect 2281 -3718 2293 -3684
rect 2293 -3718 2327 -3684
rect 2327 -3718 2339 -3684
rect 2281 -3792 2339 -3718
rect 2281 -3826 2293 -3792
rect 2293 -3826 2327 -3792
rect 2327 -3826 2339 -3792
rect 2281 -3832 2339 -3826
rect 2399 -3684 2457 -3678
rect 2399 -3718 2411 -3684
rect 2411 -3718 2445 -3684
rect 2445 -3718 2457 -3684
rect 2399 -3792 2457 -3718
rect 2399 -3826 2411 -3792
rect 2411 -3826 2445 -3792
rect 2445 -3826 2457 -3792
rect 2399 -3832 2457 -3826
rect 2517 -3684 2575 -3678
rect 2517 -3718 2529 -3684
rect 2529 -3718 2563 -3684
rect 2563 -3718 2575 -3684
rect 2517 -3792 2575 -3718
rect 2517 -3826 2529 -3792
rect 2529 -3826 2563 -3792
rect 2563 -3826 2575 -3792
rect 2517 -3832 2575 -3826
rect 2635 -3684 2693 -3678
rect 2635 -3718 2647 -3684
rect 2647 -3718 2681 -3684
rect 2681 -3718 2693 -3684
rect 2635 -3792 2693 -3718
rect 2635 -3826 2647 -3792
rect 2647 -3826 2681 -3792
rect 2681 -3826 2693 -3792
rect 2635 -3832 2693 -3826
rect 2753 -3684 2811 -3678
rect 2753 -3718 2765 -3684
rect 2765 -3718 2799 -3684
rect 2799 -3718 2811 -3684
rect 2753 -3792 2811 -3718
rect 2753 -3826 2765 -3792
rect 2765 -3826 2799 -3792
rect 2799 -3826 2811 -3792
rect 2753 -3832 2811 -3826
rect 2871 -3684 2929 -3678
rect 2871 -3718 2883 -3684
rect 2883 -3718 2917 -3684
rect 2917 -3718 2929 -3684
rect 2871 -3792 2929 -3718
rect 2871 -3826 2883 -3792
rect 2883 -3826 2917 -3792
rect 2917 -3826 2929 -3792
rect 2871 -3832 2929 -3826
rect 2989 -3684 3047 -3678
rect 2989 -3718 3001 -3684
rect 3001 -3718 3035 -3684
rect 3035 -3718 3047 -3684
rect 2989 -3792 3047 -3718
rect 2989 -3826 3001 -3792
rect 3001 -3826 3035 -3792
rect 3035 -3826 3047 -3792
rect 2989 -3832 3047 -3826
rect 3107 -3684 3165 -3678
rect 3107 -3718 3119 -3684
rect 3119 -3718 3153 -3684
rect 3153 -3718 3165 -3684
rect 3107 -3792 3165 -3718
rect 3107 -3826 3119 -3792
rect 3119 -3826 3153 -3792
rect 3153 -3826 3165 -3792
rect 3107 -3832 3165 -3826
rect 3225 -3684 3283 -3678
rect 3225 -3718 3237 -3684
rect 3237 -3718 3271 -3684
rect 3271 -3718 3283 -3684
rect 3225 -3792 3283 -3718
rect 3225 -3826 3237 -3792
rect 3237 -3826 3271 -3792
rect 3271 -3826 3283 -3792
rect 3225 -3832 3283 -3826
rect 3343 -3684 3401 -3678
rect 3343 -3718 3355 -3684
rect 3355 -3718 3389 -3684
rect 3389 -3718 3401 -3684
rect 3343 -3792 3401 -3718
rect 3343 -3826 3355 -3792
rect 3355 -3826 3389 -3792
rect 3389 -3826 3401 -3792
rect 3343 -3832 3401 -3826
rect 3461 -3684 3519 -3678
rect 3461 -3718 3473 -3684
rect 3473 -3718 3507 -3684
rect 3507 -3718 3519 -3684
rect 3461 -3792 3519 -3718
rect 3461 -3826 3473 -3792
rect 3473 -3826 3507 -3792
rect 3507 -3826 3519 -3792
rect 3461 -3832 3519 -3826
rect 3579 -3684 3637 -3678
rect 3579 -3718 3591 -3684
rect 3591 -3718 3625 -3684
rect 3625 -3718 3637 -3684
rect 3579 -3792 3637 -3718
rect 3579 -3826 3591 -3792
rect 3591 -3826 3625 -3792
rect 3625 -3826 3637 -3792
rect 3579 -3832 3637 -3826
rect 3697 -3684 3755 -3678
rect 3697 -3718 3709 -3684
rect 3709 -3718 3743 -3684
rect 3743 -3718 3755 -3684
rect 3697 -3792 3755 -3718
rect 3697 -3826 3709 -3792
rect 3709 -3826 3743 -3792
rect 3743 -3826 3755 -3792
rect 3697 -3832 3755 -3826
rect 3815 -3684 3873 -3678
rect 3815 -3718 3827 -3684
rect 3827 -3718 3861 -3684
rect 3861 -3718 3873 -3684
rect 3815 -3792 3873 -3718
rect 3815 -3826 3827 -3792
rect 3827 -3826 3861 -3792
rect 3861 -3826 3873 -3792
rect 3815 -3832 3873 -3826
rect 3933 -3684 3991 -3678
rect 3933 -3718 3945 -3684
rect 3945 -3718 3979 -3684
rect 3979 -3718 3991 -3684
rect 3933 -3792 3991 -3718
rect 3933 -3826 3945 -3792
rect 3945 -3826 3979 -3792
rect 3979 -3826 3991 -3792
rect 3933 -3832 3991 -3826
rect 4051 -3684 4109 -3678
rect 4051 -3718 4063 -3684
rect 4063 -3718 4097 -3684
rect 4097 -3718 4109 -3684
rect 4051 -3792 4109 -3718
rect 4051 -3826 4063 -3792
rect 4063 -3826 4097 -3792
rect 4097 -3826 4109 -3792
rect 4051 -3832 4109 -3826
rect 4169 -3684 4227 -3678
rect 4169 -3718 4181 -3684
rect 4181 -3718 4215 -3684
rect 4215 -3718 4227 -3684
rect 4169 -3792 4227 -3718
rect 4169 -3826 4181 -3792
rect 4181 -3826 4215 -3792
rect 4215 -3826 4227 -3792
rect 4169 -3832 4227 -3826
rect 4287 -3684 4345 -3678
rect 4287 -3718 4299 -3684
rect 4299 -3718 4333 -3684
rect 4333 -3718 4345 -3684
rect 4287 -3792 4345 -3718
rect 4287 -3826 4299 -3792
rect 4299 -3826 4333 -3792
rect 4333 -3826 4345 -3792
rect 4287 -3832 4345 -3826
rect 4405 -3684 4463 -3678
rect 4405 -3718 4417 -3684
rect 4417 -3718 4451 -3684
rect 4451 -3718 4463 -3684
rect 4405 -3792 4463 -3718
rect 4405 -3826 4417 -3792
rect 4417 -3826 4451 -3792
rect 4451 -3826 4463 -3792
rect 4405 -3832 4463 -3826
rect 4523 -3684 4581 -3678
rect 4523 -3718 4535 -3684
rect 4535 -3718 4569 -3684
rect 4569 -3718 4581 -3684
rect 4523 -3792 4581 -3718
rect 4523 -3826 4535 -3792
rect 4535 -3826 4569 -3792
rect 4569 -3826 4581 -3792
rect 4523 -3832 4581 -3826
rect 4641 -3684 4699 -3678
rect 4641 -3718 4653 -3684
rect 4653 -3718 4687 -3684
rect 4687 -3718 4699 -3684
rect 4641 -3792 4699 -3718
rect 4641 -3826 4653 -3792
rect 4653 -3826 4687 -3792
rect 4687 -3826 4699 -3792
rect 4641 -3832 4699 -3826
rect 4759 -3684 4817 -3678
rect 4759 -3718 4771 -3684
rect 4771 -3718 4805 -3684
rect 4805 -3718 4817 -3684
rect 4759 -3792 4817 -3718
rect 4759 -3826 4771 -3792
rect 4771 -3826 4805 -3792
rect 4805 -3826 4817 -3792
rect 4759 -3832 4817 -3826
rect 4877 -3684 4935 -3678
rect 4877 -3718 4889 -3684
rect 4889 -3718 4923 -3684
rect 4923 -3718 4935 -3684
rect 4877 -3792 4935 -3718
rect 4877 -3826 4889 -3792
rect 4889 -3826 4923 -3792
rect 4923 -3826 4935 -3792
rect 4877 -3832 4935 -3826
rect 4995 -3684 5053 -3678
rect 4995 -3718 5007 -3684
rect 5007 -3718 5041 -3684
rect 5041 -3718 5053 -3684
rect 4995 -3792 5053 -3718
rect 4995 -3826 5007 -3792
rect 5007 -3826 5041 -3792
rect 5041 -3826 5053 -3792
rect 4995 -3832 5053 -3826
rect 5113 -3684 5171 -3678
rect 5113 -3718 5125 -3684
rect 5125 -3718 5159 -3684
rect 5159 -3718 5171 -3684
rect 5113 -3792 5171 -3718
rect 5113 -3826 5125 -3792
rect 5125 -3826 5159 -3792
rect 5159 -3826 5171 -3792
rect 5113 -3832 5171 -3826
rect 5231 -3684 5289 -3678
rect 5231 -3718 5243 -3684
rect 5243 -3718 5277 -3684
rect 5277 -3718 5289 -3684
rect 5231 -3792 5289 -3718
rect 5231 -3826 5243 -3792
rect 5243 -3826 5277 -3792
rect 5277 -3826 5289 -3792
rect 5231 -3832 5289 -3826
rect 5349 -3684 5407 -3678
rect 5349 -3718 5361 -3684
rect 5361 -3718 5395 -3684
rect 5395 -3718 5407 -3684
rect 5349 -3792 5407 -3718
rect 5349 -3826 5361 -3792
rect 5361 -3826 5395 -3792
rect 5395 -3826 5407 -3792
rect 5349 -3832 5407 -3826
rect 5467 -3684 5525 -3678
rect 5467 -3718 5479 -3684
rect 5479 -3718 5513 -3684
rect 5513 -3718 5525 -3684
rect 5467 -3792 5525 -3718
rect 5467 -3826 5479 -3792
rect 5479 -3826 5513 -3792
rect 5513 -3826 5525 -3792
rect 5467 -3832 5525 -3826
rect 5585 -3684 5643 -3678
rect 5585 -3718 5597 -3684
rect 5597 -3718 5631 -3684
rect 5631 -3718 5643 -3684
rect 5585 -3792 5643 -3718
rect 5585 -3826 5597 -3792
rect 5597 -3826 5631 -3792
rect 5631 -3826 5643 -3792
rect 5585 -3832 5643 -3826
rect 5703 -3684 5761 -3678
rect 5703 -3718 5715 -3684
rect 5715 -3718 5749 -3684
rect 5749 -3718 5761 -3684
rect 5703 -3792 5761 -3718
rect 5703 -3826 5715 -3792
rect 5715 -3826 5749 -3792
rect 5749 -3826 5761 -3792
rect 5703 -3832 5761 -3826
rect 5821 -3684 5879 -3678
rect 5821 -3718 5833 -3684
rect 5833 -3718 5867 -3684
rect 5867 -3718 5879 -3684
rect 5821 -3792 5879 -3718
rect 5821 -3826 5833 -3792
rect 5833 -3826 5867 -3792
rect 5867 -3826 5879 -3792
rect 5821 -3832 5879 -3826
rect 5939 -3684 5997 -3678
rect 5939 -3718 5951 -3684
rect 5951 -3718 5985 -3684
rect 5985 -3718 5997 -3684
rect 5939 -3792 5997 -3718
rect 5939 -3826 5951 -3792
rect 5951 -3826 5985 -3792
rect 5985 -3826 5997 -3792
rect 5939 -3832 5997 -3826
rect 6057 -3684 6115 -3678
rect 6057 -3718 6069 -3684
rect 6069 -3718 6103 -3684
rect 6103 -3718 6115 -3684
rect 6057 -3792 6115 -3718
rect 6057 -3826 6069 -3792
rect 6069 -3826 6103 -3792
rect 6103 -3826 6115 -3792
rect 6057 -3832 6115 -3826
rect 6175 -3684 6233 -3678
rect 6175 -3718 6187 -3684
rect 6187 -3718 6221 -3684
rect 6221 -3718 6233 -3684
rect 6175 -3792 6233 -3718
rect 6175 -3826 6187 -3792
rect 6187 -3826 6221 -3792
rect 6221 -3826 6233 -3792
rect 6175 -3832 6233 -3826
rect 6293 -3684 6351 -3678
rect 6293 -3718 6305 -3684
rect 6305 -3718 6339 -3684
rect 6339 -3718 6351 -3684
rect 6293 -3792 6351 -3718
rect 6293 -3826 6305 -3792
rect 6305 -3826 6339 -3792
rect 6339 -3826 6351 -3792
rect 6293 -3832 6351 -3826
rect 6411 -3684 6469 -3678
rect 6411 -3718 6423 -3684
rect 6423 -3718 6457 -3684
rect 6457 -3718 6469 -3684
rect 6411 -3792 6469 -3718
rect 6411 -3826 6423 -3792
rect 6423 -3826 6457 -3792
rect 6457 -3826 6469 -3792
rect 6411 -3832 6469 -3826
rect 6529 -3684 6587 -3678
rect 6529 -3718 6541 -3684
rect 6541 -3718 6575 -3684
rect 6575 -3718 6587 -3684
rect 6529 -3792 6587 -3718
rect 6529 -3826 6541 -3792
rect 6541 -3826 6575 -3792
rect 6575 -3826 6587 -3792
rect 6529 -3832 6587 -3826
rect 6647 -3684 6705 -3678
rect 6647 -3718 6659 -3684
rect 6659 -3718 6693 -3684
rect 6693 -3718 6705 -3684
rect 6647 -3792 6705 -3718
rect 6647 -3826 6659 -3792
rect 6659 -3826 6693 -3792
rect 6693 -3826 6705 -3792
rect 6647 -3832 6705 -3826
rect 6765 -3684 6823 -3678
rect 6765 -3718 6777 -3684
rect 6777 -3718 6811 -3684
rect 6811 -3718 6823 -3684
rect 6765 -3792 6823 -3718
rect 6765 -3826 6777 -3792
rect 6777 -3826 6811 -3792
rect 6811 -3826 6823 -3792
rect 6765 -3832 6823 -3826
rect 6883 -3684 6941 -3678
rect 6883 -3718 6895 -3684
rect 6895 -3718 6929 -3684
rect 6929 -3718 6941 -3684
rect 6883 -3792 6941 -3718
rect 6883 -3826 6895 -3792
rect 6895 -3826 6929 -3792
rect 6929 -3826 6941 -3792
rect 6883 -3832 6941 -3826
rect 7001 -3684 7059 -3678
rect 7001 -3718 7013 -3684
rect 7013 -3718 7047 -3684
rect 7047 -3718 7059 -3684
rect 7001 -3792 7059 -3718
rect 7001 -3826 7013 -3792
rect 7013 -3826 7047 -3792
rect 7047 -3826 7059 -3792
rect 7001 -3832 7059 -3826
rect 7119 -3684 7177 -3678
rect 7119 -3718 7131 -3684
rect 7131 -3718 7165 -3684
rect 7165 -3718 7177 -3684
rect 7119 -3792 7177 -3718
rect 7119 -3826 7131 -3792
rect 7131 -3826 7165 -3792
rect 7165 -3826 7177 -3792
rect 7119 -3832 7177 -3826
rect 1337 -5452 1395 -5446
rect 1337 -5486 1349 -5452
rect 1349 -5486 1383 -5452
rect 1383 -5486 1395 -5452
rect 1337 -5560 1395 -5486
rect 1337 -5594 1349 -5560
rect 1349 -5594 1383 -5560
rect 1383 -5594 1395 -5560
rect 1337 -5600 1395 -5594
rect 1455 -5452 1513 -5446
rect 1455 -5486 1467 -5452
rect 1467 -5486 1501 -5452
rect 1501 -5486 1513 -5452
rect 1455 -5560 1513 -5486
rect 1455 -5594 1467 -5560
rect 1467 -5594 1501 -5560
rect 1501 -5594 1513 -5560
rect 1455 -5600 1513 -5594
rect 1573 -5452 1631 -5446
rect 1573 -5486 1585 -5452
rect 1585 -5486 1619 -5452
rect 1619 -5486 1631 -5452
rect 1573 -5560 1631 -5486
rect 1573 -5594 1585 -5560
rect 1585 -5594 1619 -5560
rect 1619 -5594 1631 -5560
rect 1573 -5600 1631 -5594
rect 1691 -5452 1749 -5446
rect 1691 -5486 1703 -5452
rect 1703 -5486 1737 -5452
rect 1737 -5486 1749 -5452
rect 1691 -5560 1749 -5486
rect 1691 -5594 1703 -5560
rect 1703 -5594 1737 -5560
rect 1737 -5594 1749 -5560
rect 1691 -5600 1749 -5594
rect 1809 -5452 1867 -5446
rect 1809 -5486 1821 -5452
rect 1821 -5486 1855 -5452
rect 1855 -5486 1867 -5452
rect 1809 -5560 1867 -5486
rect 1809 -5594 1821 -5560
rect 1821 -5594 1855 -5560
rect 1855 -5594 1867 -5560
rect 1809 -5600 1867 -5594
rect 1927 -5452 1985 -5446
rect 1927 -5486 1939 -5452
rect 1939 -5486 1973 -5452
rect 1973 -5486 1985 -5452
rect 1927 -5560 1985 -5486
rect 1927 -5594 1939 -5560
rect 1939 -5594 1973 -5560
rect 1973 -5594 1985 -5560
rect 1927 -5600 1985 -5594
rect 2045 -5452 2103 -5446
rect 2045 -5486 2057 -5452
rect 2057 -5486 2091 -5452
rect 2091 -5486 2103 -5452
rect 2045 -5560 2103 -5486
rect 2045 -5594 2057 -5560
rect 2057 -5594 2091 -5560
rect 2091 -5594 2103 -5560
rect 2045 -5600 2103 -5594
rect 2163 -5452 2221 -5446
rect 2163 -5486 2175 -5452
rect 2175 -5486 2209 -5452
rect 2209 -5486 2221 -5452
rect 2163 -5560 2221 -5486
rect 2163 -5594 2175 -5560
rect 2175 -5594 2209 -5560
rect 2209 -5594 2221 -5560
rect 2163 -5600 2221 -5594
rect 2281 -5452 2339 -5446
rect 2281 -5486 2293 -5452
rect 2293 -5486 2327 -5452
rect 2327 -5486 2339 -5452
rect 2281 -5560 2339 -5486
rect 2281 -5594 2293 -5560
rect 2293 -5594 2327 -5560
rect 2327 -5594 2339 -5560
rect 2281 -5600 2339 -5594
rect 2399 -5452 2457 -5446
rect 2399 -5486 2411 -5452
rect 2411 -5486 2445 -5452
rect 2445 -5486 2457 -5452
rect 2399 -5560 2457 -5486
rect 2399 -5594 2411 -5560
rect 2411 -5594 2445 -5560
rect 2445 -5594 2457 -5560
rect 2399 -5600 2457 -5594
rect 2517 -5452 2575 -5446
rect 2517 -5486 2529 -5452
rect 2529 -5486 2563 -5452
rect 2563 -5486 2575 -5452
rect 2517 -5560 2575 -5486
rect 2517 -5594 2529 -5560
rect 2529 -5594 2563 -5560
rect 2563 -5594 2575 -5560
rect 2517 -5600 2575 -5594
rect 2635 -5452 2693 -5446
rect 2635 -5486 2647 -5452
rect 2647 -5486 2681 -5452
rect 2681 -5486 2693 -5452
rect 2635 -5560 2693 -5486
rect 2635 -5594 2647 -5560
rect 2647 -5594 2681 -5560
rect 2681 -5594 2693 -5560
rect 2635 -5600 2693 -5594
rect 2753 -5452 2811 -5446
rect 2753 -5486 2765 -5452
rect 2765 -5486 2799 -5452
rect 2799 -5486 2811 -5452
rect 2753 -5560 2811 -5486
rect 2753 -5594 2765 -5560
rect 2765 -5594 2799 -5560
rect 2799 -5594 2811 -5560
rect 2753 -5600 2811 -5594
rect 2871 -5452 2929 -5446
rect 2871 -5486 2883 -5452
rect 2883 -5486 2917 -5452
rect 2917 -5486 2929 -5452
rect 2871 -5560 2929 -5486
rect 2871 -5594 2883 -5560
rect 2883 -5594 2917 -5560
rect 2917 -5594 2929 -5560
rect 2871 -5600 2929 -5594
rect 2989 -5452 3047 -5446
rect 2989 -5486 3001 -5452
rect 3001 -5486 3035 -5452
rect 3035 -5486 3047 -5452
rect 2989 -5560 3047 -5486
rect 2989 -5594 3001 -5560
rect 3001 -5594 3035 -5560
rect 3035 -5594 3047 -5560
rect 2989 -5600 3047 -5594
rect 3107 -5452 3165 -5446
rect 3107 -5486 3119 -5452
rect 3119 -5486 3153 -5452
rect 3153 -5486 3165 -5452
rect 3107 -5560 3165 -5486
rect 3107 -5594 3119 -5560
rect 3119 -5594 3153 -5560
rect 3153 -5594 3165 -5560
rect 3107 -5600 3165 -5594
rect 3225 -5452 3283 -5446
rect 3225 -5486 3237 -5452
rect 3237 -5486 3271 -5452
rect 3271 -5486 3283 -5452
rect 3225 -5560 3283 -5486
rect 3225 -5594 3237 -5560
rect 3237 -5594 3271 -5560
rect 3271 -5594 3283 -5560
rect 3225 -5600 3283 -5594
rect 3343 -5452 3401 -5446
rect 3343 -5486 3355 -5452
rect 3355 -5486 3389 -5452
rect 3389 -5486 3401 -5452
rect 3343 -5560 3401 -5486
rect 3343 -5594 3355 -5560
rect 3355 -5594 3389 -5560
rect 3389 -5594 3401 -5560
rect 3343 -5600 3401 -5594
rect 3461 -5452 3519 -5446
rect 3461 -5486 3473 -5452
rect 3473 -5486 3507 -5452
rect 3507 -5486 3519 -5452
rect 3461 -5560 3519 -5486
rect 3461 -5594 3473 -5560
rect 3473 -5594 3507 -5560
rect 3507 -5594 3519 -5560
rect 3461 -5600 3519 -5594
rect 3579 -5452 3637 -5446
rect 3579 -5486 3591 -5452
rect 3591 -5486 3625 -5452
rect 3625 -5486 3637 -5452
rect 3579 -5560 3637 -5486
rect 3579 -5594 3591 -5560
rect 3591 -5594 3625 -5560
rect 3625 -5594 3637 -5560
rect 3579 -5600 3637 -5594
rect 3697 -5452 3755 -5446
rect 3697 -5486 3709 -5452
rect 3709 -5486 3743 -5452
rect 3743 -5486 3755 -5452
rect 3697 -5560 3755 -5486
rect 3697 -5594 3709 -5560
rect 3709 -5594 3743 -5560
rect 3743 -5594 3755 -5560
rect 3697 -5600 3755 -5594
rect 3815 -5452 3873 -5446
rect 3815 -5486 3827 -5452
rect 3827 -5486 3861 -5452
rect 3861 -5486 3873 -5452
rect 3815 -5560 3873 -5486
rect 3815 -5594 3827 -5560
rect 3827 -5594 3861 -5560
rect 3861 -5594 3873 -5560
rect 3815 -5600 3873 -5594
rect 3933 -5452 3991 -5446
rect 3933 -5486 3945 -5452
rect 3945 -5486 3979 -5452
rect 3979 -5486 3991 -5452
rect 3933 -5560 3991 -5486
rect 3933 -5594 3945 -5560
rect 3945 -5594 3979 -5560
rect 3979 -5594 3991 -5560
rect 3933 -5600 3991 -5594
rect 4051 -5452 4109 -5446
rect 4051 -5486 4063 -5452
rect 4063 -5486 4097 -5452
rect 4097 -5486 4109 -5452
rect 4051 -5560 4109 -5486
rect 4051 -5594 4063 -5560
rect 4063 -5594 4097 -5560
rect 4097 -5594 4109 -5560
rect 4051 -5600 4109 -5594
rect 4169 -5452 4227 -5446
rect 4169 -5486 4181 -5452
rect 4181 -5486 4215 -5452
rect 4215 -5486 4227 -5452
rect 4169 -5560 4227 -5486
rect 4169 -5594 4181 -5560
rect 4181 -5594 4215 -5560
rect 4215 -5594 4227 -5560
rect 4169 -5600 4227 -5594
rect 4287 -5452 4345 -5446
rect 4287 -5486 4299 -5452
rect 4299 -5486 4333 -5452
rect 4333 -5486 4345 -5452
rect 4287 -5560 4345 -5486
rect 4287 -5594 4299 -5560
rect 4299 -5594 4333 -5560
rect 4333 -5594 4345 -5560
rect 4287 -5600 4345 -5594
rect 4405 -5452 4463 -5446
rect 4405 -5486 4417 -5452
rect 4417 -5486 4451 -5452
rect 4451 -5486 4463 -5452
rect 4405 -5560 4463 -5486
rect 4405 -5594 4417 -5560
rect 4417 -5594 4451 -5560
rect 4451 -5594 4463 -5560
rect 4405 -5600 4463 -5594
rect 4523 -5452 4581 -5446
rect 4523 -5486 4535 -5452
rect 4535 -5486 4569 -5452
rect 4569 -5486 4581 -5452
rect 4523 -5560 4581 -5486
rect 4523 -5594 4535 -5560
rect 4535 -5594 4569 -5560
rect 4569 -5594 4581 -5560
rect 4523 -5600 4581 -5594
rect 4641 -5452 4699 -5446
rect 4641 -5486 4653 -5452
rect 4653 -5486 4687 -5452
rect 4687 -5486 4699 -5452
rect 4641 -5560 4699 -5486
rect 4641 -5594 4653 -5560
rect 4653 -5594 4687 -5560
rect 4687 -5594 4699 -5560
rect 4641 -5600 4699 -5594
rect 4759 -5452 4817 -5446
rect 4759 -5486 4771 -5452
rect 4771 -5486 4805 -5452
rect 4805 -5486 4817 -5452
rect 4759 -5560 4817 -5486
rect 4759 -5594 4771 -5560
rect 4771 -5594 4805 -5560
rect 4805 -5594 4817 -5560
rect 4759 -5600 4817 -5594
rect 4877 -5452 4935 -5446
rect 4877 -5486 4889 -5452
rect 4889 -5486 4923 -5452
rect 4923 -5486 4935 -5452
rect 4877 -5560 4935 -5486
rect 4877 -5594 4889 -5560
rect 4889 -5594 4923 -5560
rect 4923 -5594 4935 -5560
rect 4877 -5600 4935 -5594
rect 4995 -5452 5053 -5446
rect 4995 -5486 5007 -5452
rect 5007 -5486 5041 -5452
rect 5041 -5486 5053 -5452
rect 4995 -5560 5053 -5486
rect 4995 -5594 5007 -5560
rect 5007 -5594 5041 -5560
rect 5041 -5594 5053 -5560
rect 4995 -5600 5053 -5594
rect 5113 -5452 5171 -5446
rect 5113 -5486 5125 -5452
rect 5125 -5486 5159 -5452
rect 5159 -5486 5171 -5452
rect 5113 -5560 5171 -5486
rect 5113 -5594 5125 -5560
rect 5125 -5594 5159 -5560
rect 5159 -5594 5171 -5560
rect 5113 -5600 5171 -5594
rect 5231 -5452 5289 -5446
rect 5231 -5486 5243 -5452
rect 5243 -5486 5277 -5452
rect 5277 -5486 5289 -5452
rect 5231 -5560 5289 -5486
rect 5231 -5594 5243 -5560
rect 5243 -5594 5277 -5560
rect 5277 -5594 5289 -5560
rect 5231 -5600 5289 -5594
rect 5349 -5452 5407 -5446
rect 5349 -5486 5361 -5452
rect 5361 -5486 5395 -5452
rect 5395 -5486 5407 -5452
rect 5349 -5560 5407 -5486
rect 5349 -5594 5361 -5560
rect 5361 -5594 5395 -5560
rect 5395 -5594 5407 -5560
rect 5349 -5600 5407 -5594
rect 5467 -5452 5525 -5446
rect 5467 -5486 5479 -5452
rect 5479 -5486 5513 -5452
rect 5513 -5486 5525 -5452
rect 5467 -5560 5525 -5486
rect 5467 -5594 5479 -5560
rect 5479 -5594 5513 -5560
rect 5513 -5594 5525 -5560
rect 5467 -5600 5525 -5594
rect 5585 -5452 5643 -5446
rect 5585 -5486 5597 -5452
rect 5597 -5486 5631 -5452
rect 5631 -5486 5643 -5452
rect 5585 -5560 5643 -5486
rect 5585 -5594 5597 -5560
rect 5597 -5594 5631 -5560
rect 5631 -5594 5643 -5560
rect 5585 -5600 5643 -5594
rect 5703 -5452 5761 -5446
rect 5703 -5486 5715 -5452
rect 5715 -5486 5749 -5452
rect 5749 -5486 5761 -5452
rect 5703 -5560 5761 -5486
rect 5703 -5594 5715 -5560
rect 5715 -5594 5749 -5560
rect 5749 -5594 5761 -5560
rect 5703 -5600 5761 -5594
rect 5821 -5452 5879 -5446
rect 5821 -5486 5833 -5452
rect 5833 -5486 5867 -5452
rect 5867 -5486 5879 -5452
rect 5821 -5560 5879 -5486
rect 5821 -5594 5833 -5560
rect 5833 -5594 5867 -5560
rect 5867 -5594 5879 -5560
rect 5821 -5600 5879 -5594
rect 5939 -5452 5997 -5446
rect 5939 -5486 5951 -5452
rect 5951 -5486 5985 -5452
rect 5985 -5486 5997 -5452
rect 5939 -5560 5997 -5486
rect 5939 -5594 5951 -5560
rect 5951 -5594 5985 -5560
rect 5985 -5594 5997 -5560
rect 5939 -5600 5997 -5594
rect 6057 -5452 6115 -5446
rect 6057 -5486 6069 -5452
rect 6069 -5486 6103 -5452
rect 6103 -5486 6115 -5452
rect 6057 -5560 6115 -5486
rect 6057 -5594 6069 -5560
rect 6069 -5594 6103 -5560
rect 6103 -5594 6115 -5560
rect 6057 -5600 6115 -5594
rect 6175 -5452 6233 -5446
rect 6175 -5486 6187 -5452
rect 6187 -5486 6221 -5452
rect 6221 -5486 6233 -5452
rect 6175 -5560 6233 -5486
rect 6175 -5594 6187 -5560
rect 6187 -5594 6221 -5560
rect 6221 -5594 6233 -5560
rect 6175 -5600 6233 -5594
rect 6293 -5452 6351 -5446
rect 6293 -5486 6305 -5452
rect 6305 -5486 6339 -5452
rect 6339 -5486 6351 -5452
rect 6293 -5560 6351 -5486
rect 6293 -5594 6305 -5560
rect 6305 -5594 6339 -5560
rect 6339 -5594 6351 -5560
rect 6293 -5600 6351 -5594
rect 6411 -5452 6469 -5446
rect 6411 -5486 6423 -5452
rect 6423 -5486 6457 -5452
rect 6457 -5486 6469 -5452
rect 6411 -5560 6469 -5486
rect 6411 -5594 6423 -5560
rect 6423 -5594 6457 -5560
rect 6457 -5594 6469 -5560
rect 6411 -5600 6469 -5594
rect 6529 -5452 6587 -5446
rect 6529 -5486 6541 -5452
rect 6541 -5486 6575 -5452
rect 6575 -5486 6587 -5452
rect 6529 -5560 6587 -5486
rect 6529 -5594 6541 -5560
rect 6541 -5594 6575 -5560
rect 6575 -5594 6587 -5560
rect 6529 -5600 6587 -5594
rect 6647 -5452 6705 -5446
rect 6647 -5486 6659 -5452
rect 6659 -5486 6693 -5452
rect 6693 -5486 6705 -5452
rect 6647 -5560 6705 -5486
rect 6647 -5594 6659 -5560
rect 6659 -5594 6693 -5560
rect 6693 -5594 6705 -5560
rect 6647 -5600 6705 -5594
rect 6765 -5452 6823 -5446
rect 6765 -5486 6777 -5452
rect 6777 -5486 6811 -5452
rect 6811 -5486 6823 -5452
rect 6765 -5560 6823 -5486
rect 6765 -5594 6777 -5560
rect 6777 -5594 6811 -5560
rect 6811 -5594 6823 -5560
rect 6765 -5600 6823 -5594
rect 6883 -5452 6941 -5446
rect 6883 -5486 6895 -5452
rect 6895 -5486 6929 -5452
rect 6929 -5486 6941 -5452
rect 6883 -5560 6941 -5486
rect 6883 -5594 6895 -5560
rect 6895 -5594 6929 -5560
rect 6929 -5594 6941 -5560
rect 6883 -5600 6941 -5594
rect 7001 -5452 7059 -5446
rect 7001 -5486 7013 -5452
rect 7013 -5486 7047 -5452
rect 7047 -5486 7059 -5452
rect 7001 -5560 7059 -5486
rect 7001 -5594 7013 -5560
rect 7013 -5594 7047 -5560
rect 7047 -5594 7059 -5560
rect 7001 -5600 7059 -5594
rect 7119 -5452 7177 -5446
rect 7119 -5486 7131 -5452
rect 7131 -5486 7165 -5452
rect 7165 -5486 7177 -5452
rect 7119 -5560 7177 -5486
rect 7119 -5594 7131 -5560
rect 7131 -5594 7165 -5560
rect 7165 -5594 7177 -5560
rect 7119 -5600 7177 -5594
rect 11454 -7486 11463 -6646
rect 11463 -7486 11497 -6646
rect 11497 -7486 11506 -6646
rect 11602 -7486 11611 -6646
rect 11611 -7486 11645 -6646
rect 11645 -7486 11654 -6646
rect 11750 -7486 11759 -6646
rect 11759 -7486 11793 -6646
rect 11793 -7486 11802 -6646
rect 11898 -7486 11907 -6646
rect 11907 -7486 11941 -6646
rect 11941 -7486 11950 -6646
rect 12046 -7486 12055 -6646
rect 12055 -7486 12089 -6646
rect 12089 -7486 12098 -6646
rect 12194 -7486 12203 -6646
rect 12203 -7486 12237 -6646
rect 12237 -7486 12246 -6646
rect 12342 -7486 12351 -6646
rect 12351 -7486 12385 -6646
rect 12385 -7486 12394 -6646
rect 12490 -7486 12499 -6646
rect 12499 -7486 12533 -6646
rect 12533 -7486 12542 -6646
rect 12638 -7486 12647 -6646
rect 12647 -7486 12681 -6646
rect 12681 -7486 12690 -6646
rect 12786 -7486 12795 -6646
rect 12795 -7486 12829 -6646
rect 12829 -7486 12838 -6646
rect 12934 -7486 12943 -6646
rect 12943 -7486 12977 -6646
rect 12977 -7486 12986 -6646
rect 13082 -7486 13091 -6646
rect 13091 -7486 13125 -6646
rect 13125 -7486 13134 -6646
rect 13230 -7486 13239 -6646
rect 13239 -7486 13273 -6646
rect 13273 -7486 13282 -6646
rect 13378 -7486 13387 -6646
rect 13387 -7486 13421 -6646
rect 13421 -7486 13430 -6646
rect 13526 -7486 13535 -6646
rect 13535 -7486 13569 -6646
rect 13569 -7486 13578 -6646
rect 13674 -7486 13683 -6646
rect 13683 -7486 13717 -6646
rect 13717 -7486 13726 -6646
rect 13822 -7486 13831 -6646
rect 13831 -7486 13865 -6646
rect 13865 -7486 13874 -6646
rect 13970 -7486 13979 -6646
rect 13979 -7486 14013 -6646
rect 14013 -7486 14022 -6646
rect 14118 -7486 14127 -6646
rect 14127 -7486 14161 -6646
rect 14161 -7486 14170 -6646
rect 14266 -7486 14275 -6646
rect 14275 -7486 14309 -6646
rect 14309 -7486 14318 -6646
rect 14414 -7486 14423 -6646
rect 14423 -7486 14457 -6646
rect 14457 -7486 14466 -6646
rect 14562 -7486 14571 -6646
rect 14571 -7486 14605 -6646
rect 14605 -7486 14614 -6646
rect 14710 -7486 14719 -6646
rect 14719 -7486 14753 -6646
rect 14753 -7486 14762 -6646
rect 14858 -7486 14867 -6646
rect 14867 -7486 14901 -6646
rect 14901 -7486 14910 -6646
rect 15006 -7486 15015 -6646
rect 15015 -7486 15049 -6646
rect 15049 -7486 15058 -6646
rect 15154 -7486 15163 -6646
rect 15163 -7486 15197 -6646
rect 15197 -7486 15206 -6646
rect 15302 -7486 15311 -6646
rect 15311 -7486 15345 -6646
rect 15345 -7486 15354 -6646
rect 15450 -7486 15459 -6646
rect 15459 -7486 15493 -6646
rect 15493 -7486 15502 -6646
rect 15598 -7486 15607 -6646
rect 15607 -7486 15641 -6646
rect 15641 -7486 15650 -6646
rect 15746 -7486 15755 -6646
rect 15755 -7486 15789 -6646
rect 15789 -7486 15798 -6646
rect 15894 -7486 15903 -6646
rect 15903 -7486 15937 -6646
rect 15937 -7486 15946 -6646
rect 16042 -7486 16051 -6646
rect 16051 -7486 16085 -6646
rect 16085 -7486 16094 -6646
rect 16190 -7486 16199 -6646
rect 16199 -7486 16233 -6646
rect 16233 -7486 16242 -6646
rect 16338 -7486 16347 -6646
rect 16347 -7486 16381 -6646
rect 16381 -7486 16390 -6646
rect 16486 -7486 16495 -6646
rect 16495 -7486 16529 -6646
rect 16529 -7486 16538 -6646
rect 16634 -7486 16643 -6646
rect 16643 -7486 16677 -6646
rect 16677 -7486 16686 -6646
rect 16782 -7486 16791 -6646
rect 16791 -7486 16825 -6646
rect 16825 -7486 16834 -6646
rect 16930 -7486 16939 -6646
rect 16939 -7486 16973 -6646
rect 16973 -7486 16982 -6646
rect 17078 -7486 17087 -6646
rect 17087 -7486 17121 -6646
rect 17121 -7486 17130 -6646
rect 17226 -7486 17235 -6646
rect 17235 -7486 17269 -6646
rect 17269 -7486 17278 -6646
rect 17374 -7486 17383 -6646
rect 17383 -7486 17417 -6646
rect 17417 -7486 17426 -6646
rect 17522 -7486 17531 -6646
rect 17531 -7486 17565 -6646
rect 17565 -7486 17574 -6646
rect 17670 -7486 17679 -6646
rect 17679 -7486 17713 -6646
rect 17713 -7486 17722 -6646
rect 17818 -7486 17827 -6646
rect 17827 -7486 17861 -6646
rect 17861 -7486 17870 -6646
rect 17966 -7486 17975 -6646
rect 17975 -7486 18009 -6646
rect 18009 -7486 18018 -6646
rect 18114 -7486 18123 -6646
rect 18123 -7486 18157 -6646
rect 18157 -7486 18166 -6646
rect 18262 -7486 18271 -6646
rect 18271 -7486 18305 -6646
rect 18305 -7486 18314 -6646
rect 18410 -7486 18419 -6646
rect 18419 -7486 18453 -6646
rect 18453 -7486 18462 -6646
rect 18558 -7486 18567 -6646
rect 18567 -7486 18601 -6646
rect 18601 -7486 18610 -6646
rect 18706 -7486 18715 -6646
rect 18715 -7486 18749 -6646
rect 18749 -7486 18758 -6646
rect 18854 -7486 18863 -6646
rect 18863 -7486 18897 -6646
rect 18897 -7486 18906 -6646
rect 19002 -7486 19011 -6646
rect 19011 -7486 19045 -6646
rect 19045 -7486 19054 -6646
rect 19150 -7486 19159 -6646
rect 19159 -7486 19193 -6646
rect 19193 -7486 19202 -6646
rect 19298 -7486 19307 -6646
rect 19307 -7486 19341 -6646
rect 19341 -7486 19350 -6646
rect 19446 -7486 19455 -6646
rect 19455 -7486 19489 -6646
rect 19489 -7486 19498 -6646
rect 19594 -7486 19603 -6646
rect 19603 -7486 19637 -6646
rect 19637 -7486 19646 -6646
rect 19742 -7486 19751 -6646
rect 19751 -7486 19785 -6646
rect 19785 -7486 19794 -6646
rect 19890 -7486 19899 -6646
rect 19899 -7486 19933 -6646
rect 19933 -7486 19942 -6646
rect 20038 -7486 20047 -6646
rect 20047 -7486 20081 -6646
rect 20081 -7486 20090 -6646
rect 20186 -7486 20195 -6646
rect 20195 -7486 20229 -6646
rect 20229 -7486 20238 -6646
rect 20334 -7486 20343 -6646
rect 20343 -7486 20377 -6646
rect 20377 -7486 20386 -6646
rect 20482 -7486 20491 -6646
rect 20491 -7486 20525 -6646
rect 20525 -7486 20534 -6646
rect 20630 -7486 20639 -6646
rect 20639 -7486 20673 -6646
rect 20673 -7486 20682 -6646
rect 20778 -7486 20787 -6646
rect 20787 -7486 20821 -6646
rect 20821 -7486 20830 -6646
rect 20926 -7486 20935 -6646
rect 20935 -7486 20969 -6646
rect 20969 -7486 20978 -6646
rect 21074 -7486 21083 -6646
rect 21083 -7486 21117 -6646
rect 21117 -7486 21126 -6646
rect 21222 -7486 21231 -6646
rect 21231 -7486 21265 -6646
rect 21265 -7486 21274 -6646
rect 21370 -7486 21379 -6646
rect 21379 -7486 21413 -6646
rect 21413 -7486 21422 -6646
rect 21518 -7486 21527 -6646
rect 21527 -7486 21561 -6646
rect 21561 -7486 21570 -6646
rect 21666 -7486 21675 -6646
rect 21675 -7486 21709 -6646
rect 21709 -7486 21718 -6646
rect 21814 -7486 21823 -6646
rect 21823 -7486 21857 -6646
rect 21857 -7486 21866 -6646
rect 21962 -7486 21971 -6646
rect 21971 -7486 22005 -6646
rect 22005 -7486 22014 -6646
rect 22110 -7486 22162 -6646
rect 22258 -7486 22267 -6646
rect 22267 -7486 22301 -6646
rect 22301 -7486 22310 -6646
rect 22406 -7486 22458 -6646
rect 22554 -7486 22563 -6646
rect 22563 -7486 22597 -6646
rect 22597 -7486 22606 -6646
rect 11509 -7716 11599 -7562
rect 11657 -7568 11747 -7562
rect 11657 -7602 11673 -7568
rect 11673 -7602 11731 -7568
rect 11731 -7602 11747 -7568
rect 11657 -7676 11747 -7602
rect 11657 -7710 11673 -7676
rect 11673 -7710 11731 -7676
rect 11731 -7710 11747 -7676
rect 11657 -7716 11747 -7710
rect 11805 -7568 11895 -7562
rect 11805 -7602 11821 -7568
rect 11821 -7602 11879 -7568
rect 11879 -7602 11895 -7568
rect 11805 -7676 11895 -7602
rect 11805 -7710 11821 -7676
rect 11821 -7710 11879 -7676
rect 11879 -7710 11895 -7676
rect 11805 -7716 11895 -7710
rect 11953 -7568 12043 -7562
rect 11953 -7602 11969 -7568
rect 11969 -7602 12027 -7568
rect 12027 -7602 12043 -7568
rect 11953 -7676 12043 -7602
rect 11953 -7710 11969 -7676
rect 11969 -7710 12027 -7676
rect 12027 -7710 12043 -7676
rect 11953 -7716 12043 -7710
rect 12101 -7568 12191 -7562
rect 12101 -7602 12117 -7568
rect 12117 -7602 12175 -7568
rect 12175 -7602 12191 -7568
rect 12101 -7676 12191 -7602
rect 12101 -7710 12117 -7676
rect 12117 -7710 12175 -7676
rect 12175 -7710 12191 -7676
rect 12101 -7716 12191 -7710
rect 12249 -7568 12339 -7562
rect 12249 -7602 12265 -7568
rect 12265 -7602 12323 -7568
rect 12323 -7602 12339 -7568
rect 12249 -7676 12339 -7602
rect 12249 -7710 12265 -7676
rect 12265 -7710 12323 -7676
rect 12323 -7710 12339 -7676
rect 12249 -7716 12339 -7710
rect 12397 -7568 12487 -7562
rect 12397 -7602 12413 -7568
rect 12413 -7602 12471 -7568
rect 12471 -7602 12487 -7568
rect 12397 -7676 12487 -7602
rect 12397 -7710 12413 -7676
rect 12413 -7710 12471 -7676
rect 12471 -7710 12487 -7676
rect 12397 -7716 12487 -7710
rect 12545 -7568 12635 -7562
rect 12545 -7602 12561 -7568
rect 12561 -7602 12619 -7568
rect 12619 -7602 12635 -7568
rect 12545 -7676 12635 -7602
rect 12545 -7710 12561 -7676
rect 12561 -7710 12619 -7676
rect 12619 -7710 12635 -7676
rect 12545 -7716 12635 -7710
rect 12693 -7568 12783 -7562
rect 12693 -7602 12709 -7568
rect 12709 -7602 12767 -7568
rect 12767 -7602 12783 -7568
rect 12693 -7676 12783 -7602
rect 12693 -7710 12709 -7676
rect 12709 -7710 12767 -7676
rect 12767 -7710 12783 -7676
rect 12693 -7716 12783 -7710
rect 12841 -7568 12931 -7562
rect 12841 -7602 12857 -7568
rect 12857 -7602 12915 -7568
rect 12915 -7602 12931 -7568
rect 12841 -7676 12931 -7602
rect 12841 -7710 12857 -7676
rect 12857 -7710 12915 -7676
rect 12915 -7710 12931 -7676
rect 12841 -7716 12931 -7710
rect 12989 -7568 13079 -7562
rect 12989 -7602 13005 -7568
rect 13005 -7602 13063 -7568
rect 13063 -7602 13079 -7568
rect 12989 -7676 13079 -7602
rect 12989 -7710 13005 -7676
rect 13005 -7710 13063 -7676
rect 13063 -7710 13079 -7676
rect 12989 -7716 13079 -7710
rect 13137 -7568 13227 -7562
rect 13137 -7602 13153 -7568
rect 13153 -7602 13211 -7568
rect 13211 -7602 13227 -7568
rect 13137 -7676 13227 -7602
rect 13137 -7710 13153 -7676
rect 13153 -7710 13211 -7676
rect 13211 -7710 13227 -7676
rect 13137 -7716 13227 -7710
rect 13285 -7568 13375 -7562
rect 13285 -7602 13301 -7568
rect 13301 -7602 13359 -7568
rect 13359 -7602 13375 -7568
rect 13285 -7676 13375 -7602
rect 13285 -7710 13301 -7676
rect 13301 -7710 13359 -7676
rect 13359 -7710 13375 -7676
rect 13285 -7716 13375 -7710
rect 13433 -7568 13523 -7562
rect 13433 -7602 13449 -7568
rect 13449 -7602 13507 -7568
rect 13507 -7602 13523 -7568
rect 13433 -7676 13523 -7602
rect 13433 -7710 13449 -7676
rect 13449 -7710 13507 -7676
rect 13507 -7710 13523 -7676
rect 13433 -7716 13523 -7710
rect 13581 -7568 13671 -7562
rect 13581 -7602 13597 -7568
rect 13597 -7602 13655 -7568
rect 13655 -7602 13671 -7568
rect 13581 -7676 13671 -7602
rect 13581 -7710 13597 -7676
rect 13597 -7710 13655 -7676
rect 13655 -7710 13671 -7676
rect 13581 -7716 13671 -7710
rect 13729 -7568 13819 -7562
rect 13729 -7602 13745 -7568
rect 13745 -7602 13803 -7568
rect 13803 -7602 13819 -7568
rect 13729 -7676 13819 -7602
rect 13729 -7710 13745 -7676
rect 13745 -7710 13803 -7676
rect 13803 -7710 13819 -7676
rect 13729 -7716 13819 -7710
rect 13877 -7568 13967 -7562
rect 13877 -7602 13893 -7568
rect 13893 -7602 13951 -7568
rect 13951 -7602 13967 -7568
rect 13877 -7676 13967 -7602
rect 13877 -7710 13893 -7676
rect 13893 -7710 13951 -7676
rect 13951 -7710 13967 -7676
rect 13877 -7716 13967 -7710
rect 14025 -7568 14115 -7562
rect 14025 -7602 14041 -7568
rect 14041 -7602 14099 -7568
rect 14099 -7602 14115 -7568
rect 14025 -7676 14115 -7602
rect 14025 -7710 14041 -7676
rect 14041 -7710 14099 -7676
rect 14099 -7710 14115 -7676
rect 14025 -7716 14115 -7710
rect 14173 -7568 14263 -7562
rect 14173 -7602 14189 -7568
rect 14189 -7602 14247 -7568
rect 14247 -7602 14263 -7568
rect 14173 -7676 14263 -7602
rect 14173 -7710 14189 -7676
rect 14189 -7710 14247 -7676
rect 14247 -7710 14263 -7676
rect 14173 -7716 14263 -7710
rect 14321 -7568 14411 -7562
rect 14321 -7602 14337 -7568
rect 14337 -7602 14395 -7568
rect 14395 -7602 14411 -7568
rect 14321 -7676 14411 -7602
rect 14321 -7710 14337 -7676
rect 14337 -7710 14395 -7676
rect 14395 -7710 14411 -7676
rect 14321 -7716 14411 -7710
rect 14469 -7568 14559 -7562
rect 14469 -7602 14485 -7568
rect 14485 -7602 14543 -7568
rect 14543 -7602 14559 -7568
rect 14469 -7676 14559 -7602
rect 14469 -7710 14485 -7676
rect 14485 -7710 14543 -7676
rect 14543 -7710 14559 -7676
rect 14469 -7716 14559 -7710
rect 14617 -7568 14707 -7562
rect 14617 -7602 14633 -7568
rect 14633 -7602 14691 -7568
rect 14691 -7602 14707 -7568
rect 14617 -7676 14707 -7602
rect 14617 -7710 14633 -7676
rect 14633 -7710 14691 -7676
rect 14691 -7710 14707 -7676
rect 14617 -7716 14707 -7710
rect 14765 -7568 14855 -7562
rect 14765 -7602 14781 -7568
rect 14781 -7602 14839 -7568
rect 14839 -7602 14855 -7568
rect 14765 -7676 14855 -7602
rect 14765 -7710 14781 -7676
rect 14781 -7710 14839 -7676
rect 14839 -7710 14855 -7676
rect 14765 -7716 14855 -7710
rect 14913 -7568 15003 -7562
rect 14913 -7602 14929 -7568
rect 14929 -7602 14987 -7568
rect 14987 -7602 15003 -7568
rect 14913 -7676 15003 -7602
rect 14913 -7710 14929 -7676
rect 14929 -7710 14987 -7676
rect 14987 -7710 15003 -7676
rect 14913 -7716 15003 -7710
rect 15061 -7568 15151 -7562
rect 15061 -7602 15077 -7568
rect 15077 -7602 15135 -7568
rect 15135 -7602 15151 -7568
rect 15061 -7676 15151 -7602
rect 15061 -7710 15077 -7676
rect 15077 -7710 15135 -7676
rect 15135 -7710 15151 -7676
rect 15061 -7716 15151 -7710
rect 15209 -7568 15299 -7562
rect 15209 -7602 15225 -7568
rect 15225 -7602 15283 -7568
rect 15283 -7602 15299 -7568
rect 15209 -7676 15299 -7602
rect 15209 -7710 15225 -7676
rect 15225 -7710 15283 -7676
rect 15283 -7710 15299 -7676
rect 15209 -7716 15299 -7710
rect 15357 -7568 15447 -7562
rect 15357 -7602 15373 -7568
rect 15373 -7602 15431 -7568
rect 15431 -7602 15447 -7568
rect 15357 -7676 15447 -7602
rect 15357 -7710 15373 -7676
rect 15373 -7710 15431 -7676
rect 15431 -7710 15447 -7676
rect 15357 -7716 15447 -7710
rect 15505 -7568 15595 -7562
rect 15505 -7602 15521 -7568
rect 15521 -7602 15579 -7568
rect 15579 -7602 15595 -7568
rect 15505 -7676 15595 -7602
rect 15505 -7710 15521 -7676
rect 15521 -7710 15579 -7676
rect 15579 -7710 15595 -7676
rect 15505 -7716 15595 -7710
rect 15653 -7568 15743 -7562
rect 15653 -7602 15669 -7568
rect 15669 -7602 15727 -7568
rect 15727 -7602 15743 -7568
rect 15653 -7676 15743 -7602
rect 15653 -7710 15669 -7676
rect 15669 -7710 15727 -7676
rect 15727 -7710 15743 -7676
rect 15653 -7716 15743 -7710
rect 15801 -7568 15891 -7562
rect 15801 -7602 15817 -7568
rect 15817 -7602 15875 -7568
rect 15875 -7602 15891 -7568
rect 15801 -7676 15891 -7602
rect 15801 -7710 15817 -7676
rect 15817 -7710 15875 -7676
rect 15875 -7710 15891 -7676
rect 15801 -7716 15891 -7710
rect 15949 -7568 16039 -7562
rect 15949 -7602 15965 -7568
rect 15965 -7602 16023 -7568
rect 16023 -7602 16039 -7568
rect 15949 -7676 16039 -7602
rect 15949 -7710 15965 -7676
rect 15965 -7710 16023 -7676
rect 16023 -7710 16039 -7676
rect 15949 -7716 16039 -7710
rect 16097 -7568 16187 -7562
rect 16097 -7602 16113 -7568
rect 16113 -7602 16171 -7568
rect 16171 -7602 16187 -7568
rect 16097 -7676 16187 -7602
rect 16097 -7710 16113 -7676
rect 16113 -7710 16171 -7676
rect 16171 -7710 16187 -7676
rect 16097 -7716 16187 -7710
rect 16245 -7568 16335 -7562
rect 16245 -7602 16261 -7568
rect 16261 -7602 16319 -7568
rect 16319 -7602 16335 -7568
rect 16245 -7676 16335 -7602
rect 16245 -7710 16261 -7676
rect 16261 -7710 16319 -7676
rect 16319 -7710 16335 -7676
rect 16245 -7716 16335 -7710
rect 16393 -7568 16483 -7562
rect 16393 -7602 16409 -7568
rect 16409 -7602 16467 -7568
rect 16467 -7602 16483 -7568
rect 16393 -7676 16483 -7602
rect 16393 -7710 16409 -7676
rect 16409 -7710 16467 -7676
rect 16467 -7710 16483 -7676
rect 16393 -7716 16483 -7710
rect 16541 -7568 16631 -7562
rect 16541 -7602 16557 -7568
rect 16557 -7602 16615 -7568
rect 16615 -7602 16631 -7568
rect 16541 -7676 16631 -7602
rect 16541 -7710 16557 -7676
rect 16557 -7710 16615 -7676
rect 16615 -7710 16631 -7676
rect 16541 -7716 16631 -7710
rect 16689 -7568 16779 -7562
rect 16689 -7602 16705 -7568
rect 16705 -7602 16763 -7568
rect 16763 -7602 16779 -7568
rect 16689 -7676 16779 -7602
rect 16689 -7710 16705 -7676
rect 16705 -7710 16763 -7676
rect 16763 -7710 16779 -7676
rect 16689 -7716 16779 -7710
rect 16837 -7568 16927 -7562
rect 16837 -7602 16853 -7568
rect 16853 -7602 16911 -7568
rect 16911 -7602 16927 -7568
rect 16837 -7676 16927 -7602
rect 16837 -7710 16853 -7676
rect 16853 -7710 16911 -7676
rect 16911 -7710 16927 -7676
rect 16837 -7716 16927 -7710
rect 16985 -7568 17075 -7562
rect 16985 -7602 17001 -7568
rect 17001 -7602 17059 -7568
rect 17059 -7602 17075 -7568
rect 16985 -7676 17075 -7602
rect 16985 -7710 17001 -7676
rect 17001 -7710 17059 -7676
rect 17059 -7710 17075 -7676
rect 16985 -7716 17075 -7710
rect 17133 -7568 17223 -7562
rect 17133 -7602 17149 -7568
rect 17149 -7602 17207 -7568
rect 17207 -7602 17223 -7568
rect 17133 -7676 17223 -7602
rect 17133 -7710 17149 -7676
rect 17149 -7710 17207 -7676
rect 17207 -7710 17223 -7676
rect 17133 -7716 17223 -7710
rect 17281 -7568 17371 -7562
rect 17281 -7602 17297 -7568
rect 17297 -7602 17355 -7568
rect 17355 -7602 17371 -7568
rect 17281 -7676 17371 -7602
rect 17281 -7710 17297 -7676
rect 17297 -7710 17355 -7676
rect 17355 -7710 17371 -7676
rect 17281 -7716 17371 -7710
rect 17429 -7568 17519 -7562
rect 17429 -7602 17445 -7568
rect 17445 -7602 17503 -7568
rect 17503 -7602 17519 -7568
rect 17429 -7676 17519 -7602
rect 17429 -7710 17445 -7676
rect 17445 -7710 17503 -7676
rect 17503 -7710 17519 -7676
rect 17429 -7716 17519 -7710
rect 17577 -7568 17667 -7562
rect 17577 -7602 17593 -7568
rect 17593 -7602 17651 -7568
rect 17651 -7602 17667 -7568
rect 17577 -7676 17667 -7602
rect 17577 -7710 17593 -7676
rect 17593 -7710 17651 -7676
rect 17651 -7710 17667 -7676
rect 17577 -7716 17667 -7710
rect 17725 -7568 17815 -7562
rect 17725 -7602 17741 -7568
rect 17741 -7602 17799 -7568
rect 17799 -7602 17815 -7568
rect 17725 -7676 17815 -7602
rect 17725 -7710 17741 -7676
rect 17741 -7710 17799 -7676
rect 17799 -7710 17815 -7676
rect 17725 -7716 17815 -7710
rect 17873 -7568 17963 -7562
rect 17873 -7602 17889 -7568
rect 17889 -7602 17947 -7568
rect 17947 -7602 17963 -7568
rect 17873 -7676 17963 -7602
rect 17873 -7710 17889 -7676
rect 17889 -7710 17947 -7676
rect 17947 -7710 17963 -7676
rect 17873 -7716 17963 -7710
rect 18021 -7568 18111 -7562
rect 18021 -7602 18037 -7568
rect 18037 -7602 18095 -7568
rect 18095 -7602 18111 -7568
rect 18021 -7676 18111 -7602
rect 18021 -7710 18037 -7676
rect 18037 -7710 18095 -7676
rect 18095 -7710 18111 -7676
rect 18021 -7716 18111 -7710
rect 18169 -7568 18259 -7562
rect 18169 -7602 18185 -7568
rect 18185 -7602 18243 -7568
rect 18243 -7602 18259 -7568
rect 18169 -7676 18259 -7602
rect 18169 -7710 18185 -7676
rect 18185 -7710 18243 -7676
rect 18243 -7710 18259 -7676
rect 18169 -7716 18259 -7710
rect 18317 -7568 18407 -7562
rect 18317 -7602 18333 -7568
rect 18333 -7602 18391 -7568
rect 18391 -7602 18407 -7568
rect 18317 -7676 18407 -7602
rect 18317 -7710 18333 -7676
rect 18333 -7710 18391 -7676
rect 18391 -7710 18407 -7676
rect 18317 -7716 18407 -7710
rect 18465 -7568 18555 -7562
rect 18465 -7602 18481 -7568
rect 18481 -7602 18539 -7568
rect 18539 -7602 18555 -7568
rect 18465 -7676 18555 -7602
rect 18465 -7710 18481 -7676
rect 18481 -7710 18539 -7676
rect 18539 -7710 18555 -7676
rect 18465 -7716 18555 -7710
rect 18613 -7568 18703 -7562
rect 18613 -7602 18629 -7568
rect 18629 -7602 18687 -7568
rect 18687 -7602 18703 -7568
rect 18613 -7676 18703 -7602
rect 18613 -7710 18629 -7676
rect 18629 -7710 18687 -7676
rect 18687 -7710 18703 -7676
rect 18613 -7716 18703 -7710
rect 18761 -7568 18851 -7562
rect 18761 -7602 18777 -7568
rect 18777 -7602 18835 -7568
rect 18835 -7602 18851 -7568
rect 18761 -7676 18851 -7602
rect 18761 -7710 18777 -7676
rect 18777 -7710 18835 -7676
rect 18835 -7710 18851 -7676
rect 18761 -7716 18851 -7710
rect 18909 -7568 18999 -7562
rect 18909 -7602 18925 -7568
rect 18925 -7602 18983 -7568
rect 18983 -7602 18999 -7568
rect 18909 -7676 18999 -7602
rect 18909 -7710 18925 -7676
rect 18925 -7710 18983 -7676
rect 18983 -7710 18999 -7676
rect 18909 -7716 18999 -7710
rect 19057 -7568 19147 -7562
rect 19057 -7602 19073 -7568
rect 19073 -7602 19131 -7568
rect 19131 -7602 19147 -7568
rect 19057 -7676 19147 -7602
rect 19057 -7710 19073 -7676
rect 19073 -7710 19131 -7676
rect 19131 -7710 19147 -7676
rect 19057 -7716 19147 -7710
rect 19205 -7568 19295 -7562
rect 19205 -7602 19221 -7568
rect 19221 -7602 19279 -7568
rect 19279 -7602 19295 -7568
rect 19205 -7676 19295 -7602
rect 19205 -7710 19221 -7676
rect 19221 -7710 19279 -7676
rect 19279 -7710 19295 -7676
rect 19205 -7716 19295 -7710
rect 19353 -7568 19443 -7562
rect 19353 -7602 19369 -7568
rect 19369 -7602 19427 -7568
rect 19427 -7602 19443 -7568
rect 19353 -7676 19443 -7602
rect 19353 -7710 19369 -7676
rect 19369 -7710 19427 -7676
rect 19427 -7710 19443 -7676
rect 19353 -7716 19443 -7710
rect 19501 -7568 19591 -7562
rect 19501 -7602 19517 -7568
rect 19517 -7602 19575 -7568
rect 19575 -7602 19591 -7568
rect 19501 -7676 19591 -7602
rect 19501 -7710 19517 -7676
rect 19517 -7710 19575 -7676
rect 19575 -7710 19591 -7676
rect 19501 -7716 19591 -7710
rect 19649 -7568 19739 -7562
rect 19649 -7602 19665 -7568
rect 19665 -7602 19723 -7568
rect 19723 -7602 19739 -7568
rect 19649 -7676 19739 -7602
rect 19649 -7710 19665 -7676
rect 19665 -7710 19723 -7676
rect 19723 -7710 19739 -7676
rect 19649 -7716 19739 -7710
rect 19797 -7568 19887 -7562
rect 19797 -7602 19813 -7568
rect 19813 -7602 19871 -7568
rect 19871 -7602 19887 -7568
rect 19797 -7676 19887 -7602
rect 19797 -7710 19813 -7676
rect 19813 -7710 19871 -7676
rect 19871 -7710 19887 -7676
rect 19797 -7716 19887 -7710
rect 19945 -7568 20035 -7562
rect 19945 -7602 19961 -7568
rect 19961 -7602 20019 -7568
rect 20019 -7602 20035 -7568
rect 19945 -7676 20035 -7602
rect 19945 -7710 19961 -7676
rect 19961 -7710 20019 -7676
rect 20019 -7710 20035 -7676
rect 19945 -7716 20035 -7710
rect 20093 -7568 20183 -7562
rect 20093 -7602 20109 -7568
rect 20109 -7602 20167 -7568
rect 20167 -7602 20183 -7568
rect 20093 -7676 20183 -7602
rect 20093 -7710 20109 -7676
rect 20109 -7710 20167 -7676
rect 20167 -7710 20183 -7676
rect 20093 -7716 20183 -7710
rect 20241 -7568 20331 -7562
rect 20241 -7602 20257 -7568
rect 20257 -7602 20315 -7568
rect 20315 -7602 20331 -7568
rect 20241 -7676 20331 -7602
rect 20241 -7710 20257 -7676
rect 20257 -7710 20315 -7676
rect 20315 -7710 20331 -7676
rect 20241 -7716 20331 -7710
rect 20389 -7568 20479 -7562
rect 20389 -7602 20405 -7568
rect 20405 -7602 20463 -7568
rect 20463 -7602 20479 -7568
rect 20389 -7676 20479 -7602
rect 20389 -7710 20405 -7676
rect 20405 -7710 20463 -7676
rect 20463 -7710 20479 -7676
rect 20389 -7716 20479 -7710
rect 20537 -7568 20627 -7562
rect 20537 -7602 20553 -7568
rect 20553 -7602 20611 -7568
rect 20611 -7602 20627 -7568
rect 20537 -7676 20627 -7602
rect 20537 -7710 20553 -7676
rect 20553 -7710 20611 -7676
rect 20611 -7710 20627 -7676
rect 20537 -7716 20627 -7710
rect 20685 -7568 20775 -7562
rect 20685 -7602 20701 -7568
rect 20701 -7602 20759 -7568
rect 20759 -7602 20775 -7568
rect 20685 -7676 20775 -7602
rect 20685 -7710 20701 -7676
rect 20701 -7710 20759 -7676
rect 20759 -7710 20775 -7676
rect 20685 -7716 20775 -7710
rect 20833 -7568 20923 -7562
rect 20833 -7602 20849 -7568
rect 20849 -7602 20907 -7568
rect 20907 -7602 20923 -7568
rect 20833 -7676 20923 -7602
rect 20833 -7710 20849 -7676
rect 20849 -7710 20907 -7676
rect 20907 -7710 20923 -7676
rect 20833 -7716 20923 -7710
rect 20981 -7568 21071 -7562
rect 20981 -7602 20997 -7568
rect 20997 -7602 21055 -7568
rect 21055 -7602 21071 -7568
rect 20981 -7676 21071 -7602
rect 20981 -7710 20997 -7676
rect 20997 -7710 21055 -7676
rect 21055 -7710 21071 -7676
rect 20981 -7716 21071 -7710
rect 21129 -7568 21219 -7562
rect 21129 -7602 21145 -7568
rect 21145 -7602 21203 -7568
rect 21203 -7602 21219 -7568
rect 21129 -7676 21219 -7602
rect 21129 -7710 21145 -7676
rect 21145 -7710 21203 -7676
rect 21203 -7710 21219 -7676
rect 21129 -7716 21219 -7710
rect 21277 -7568 21367 -7562
rect 21277 -7602 21293 -7568
rect 21293 -7602 21351 -7568
rect 21351 -7602 21367 -7568
rect 21277 -7676 21367 -7602
rect 21277 -7710 21293 -7676
rect 21293 -7710 21351 -7676
rect 21351 -7710 21367 -7676
rect 21277 -7716 21367 -7710
rect 21425 -7568 21515 -7562
rect 21425 -7602 21441 -7568
rect 21441 -7602 21499 -7568
rect 21499 -7602 21515 -7568
rect 21425 -7676 21515 -7602
rect 21425 -7710 21441 -7676
rect 21441 -7710 21499 -7676
rect 21499 -7710 21515 -7676
rect 21425 -7716 21515 -7710
rect 21573 -7568 21663 -7562
rect 21573 -7602 21589 -7568
rect 21589 -7602 21647 -7568
rect 21647 -7602 21663 -7568
rect 21573 -7676 21663 -7602
rect 21573 -7710 21589 -7676
rect 21589 -7710 21647 -7676
rect 21647 -7710 21663 -7676
rect 21573 -7716 21663 -7710
rect 21721 -7568 21811 -7562
rect 21721 -7602 21737 -7568
rect 21737 -7602 21795 -7568
rect 21795 -7602 21811 -7568
rect 21721 -7676 21811 -7602
rect 21721 -7710 21737 -7676
rect 21737 -7710 21795 -7676
rect 21795 -7710 21811 -7676
rect 21721 -7716 21811 -7710
rect 21869 -7568 21959 -7562
rect 21869 -7602 21885 -7568
rect 21885 -7602 21943 -7568
rect 21943 -7602 21959 -7568
rect 21869 -7676 21959 -7602
rect 21869 -7710 21885 -7676
rect 21885 -7710 21943 -7676
rect 21943 -7710 21959 -7676
rect 21869 -7716 21959 -7710
rect 22017 -7568 22107 -7562
rect 22017 -7602 22033 -7568
rect 22033 -7602 22091 -7568
rect 22091 -7602 22107 -7568
rect 22017 -7676 22107 -7602
rect 22017 -7710 22033 -7676
rect 22033 -7710 22091 -7676
rect 22091 -7710 22107 -7676
rect 22017 -7716 22107 -7710
rect 22165 -7568 22255 -7562
rect 22165 -7602 22181 -7568
rect 22181 -7602 22239 -7568
rect 22239 -7602 22255 -7568
rect 22165 -7676 22255 -7602
rect 22165 -7710 22181 -7676
rect 22181 -7710 22239 -7676
rect 22239 -7710 22255 -7676
rect 22165 -7716 22255 -7710
rect 22313 -7568 22403 -7562
rect 22313 -7602 22329 -7568
rect 22329 -7602 22387 -7568
rect 22387 -7602 22403 -7568
rect 22313 -7676 22403 -7602
rect 22313 -7710 22329 -7676
rect 22329 -7710 22387 -7676
rect 22387 -7710 22403 -7676
rect 22313 -7716 22403 -7710
rect 22461 -7568 22551 -7562
rect 22461 -7602 22477 -7568
rect 22477 -7602 22535 -7568
rect 22535 -7602 22551 -7568
rect 22461 -7676 22551 -7602
rect 22461 -7710 22477 -7676
rect 22477 -7710 22535 -7676
rect 22535 -7710 22551 -7676
rect 22461 -7716 22551 -7710
rect 3063 -7767 3121 -7761
rect 3063 -7801 3075 -7767
rect 3075 -7801 3109 -7767
rect 3109 -7801 3121 -7767
rect 3063 -7875 3121 -7801
rect 3063 -7909 3075 -7875
rect 3075 -7909 3109 -7875
rect 3109 -7909 3121 -7875
rect 3063 -7915 3121 -7909
rect 3181 -7767 3239 -7761
rect 3181 -7801 3193 -7767
rect 3193 -7801 3227 -7767
rect 3227 -7801 3239 -7767
rect 3181 -7875 3239 -7801
rect 3181 -7909 3193 -7875
rect 3193 -7909 3227 -7875
rect 3227 -7909 3239 -7875
rect 3181 -7915 3239 -7909
rect 3299 -7767 3357 -7761
rect 3299 -7801 3311 -7767
rect 3311 -7801 3345 -7767
rect 3345 -7801 3357 -7767
rect 3299 -7875 3357 -7801
rect 3299 -7909 3311 -7875
rect 3311 -7909 3345 -7875
rect 3345 -7909 3357 -7875
rect 3299 -7915 3357 -7909
rect 3417 -7767 3475 -7761
rect 3417 -7801 3429 -7767
rect 3429 -7801 3463 -7767
rect 3463 -7801 3475 -7767
rect 3417 -7875 3475 -7801
rect 3417 -7909 3429 -7875
rect 3429 -7909 3463 -7875
rect 3463 -7909 3475 -7875
rect 3417 -7915 3475 -7909
rect 3535 -7767 3593 -7761
rect 3535 -7801 3547 -7767
rect 3547 -7801 3581 -7767
rect 3581 -7801 3593 -7767
rect 3535 -7875 3593 -7801
rect 3535 -7909 3547 -7875
rect 3547 -7909 3581 -7875
rect 3581 -7909 3593 -7875
rect 3535 -7915 3593 -7909
rect 3653 -7767 3711 -7761
rect 3653 -7801 3665 -7767
rect 3665 -7801 3699 -7767
rect 3699 -7801 3711 -7767
rect 3653 -7875 3711 -7801
rect 3653 -7909 3665 -7875
rect 3665 -7909 3699 -7875
rect 3699 -7909 3711 -7875
rect 3653 -7915 3711 -7909
rect 3771 -7767 3829 -7761
rect 3771 -7801 3783 -7767
rect 3783 -7801 3817 -7767
rect 3817 -7801 3829 -7767
rect 3771 -7875 3829 -7801
rect 3771 -7909 3783 -7875
rect 3783 -7909 3817 -7875
rect 3817 -7909 3829 -7875
rect 3771 -7915 3829 -7909
rect 3889 -7767 3947 -7761
rect 3889 -7801 3901 -7767
rect 3901 -7801 3935 -7767
rect 3935 -7801 3947 -7767
rect 3889 -7875 3947 -7801
rect 3889 -7909 3901 -7875
rect 3901 -7909 3935 -7875
rect 3935 -7909 3947 -7875
rect 3889 -7915 3947 -7909
rect 4007 -7767 4065 -7761
rect 4007 -7801 4019 -7767
rect 4019 -7801 4053 -7767
rect 4053 -7801 4065 -7767
rect 4007 -7875 4065 -7801
rect 4007 -7909 4019 -7875
rect 4019 -7909 4053 -7875
rect 4053 -7909 4065 -7875
rect 4007 -7915 4065 -7909
rect 4125 -7767 4183 -7761
rect 4125 -7801 4137 -7767
rect 4137 -7801 4171 -7767
rect 4171 -7801 4183 -7767
rect 4125 -7875 4183 -7801
rect 4125 -7909 4137 -7875
rect 4137 -7909 4171 -7875
rect 4171 -7909 4183 -7875
rect 4125 -7915 4183 -7909
rect 4243 -7767 4301 -7761
rect 4243 -7801 4255 -7767
rect 4255 -7801 4289 -7767
rect 4289 -7801 4301 -7767
rect 4243 -7875 4301 -7801
rect 4243 -7909 4255 -7875
rect 4255 -7909 4289 -7875
rect 4289 -7909 4301 -7875
rect 4243 -7915 4301 -7909
rect 4361 -7767 4419 -7761
rect 4361 -7801 4373 -7767
rect 4373 -7801 4407 -7767
rect 4407 -7801 4419 -7767
rect 4361 -7875 4419 -7801
rect 4361 -7909 4373 -7875
rect 4373 -7909 4407 -7875
rect 4407 -7909 4419 -7875
rect 4361 -7915 4419 -7909
rect 4479 -7767 4537 -7761
rect 4479 -7801 4491 -7767
rect 4491 -7801 4525 -7767
rect 4525 -7801 4537 -7767
rect 4479 -7875 4537 -7801
rect 4479 -7909 4491 -7875
rect 4491 -7909 4525 -7875
rect 4525 -7909 4537 -7875
rect 4479 -7915 4537 -7909
rect 4597 -7767 4655 -7761
rect 4597 -7801 4609 -7767
rect 4609 -7801 4643 -7767
rect 4643 -7801 4655 -7767
rect 4597 -7875 4655 -7801
rect 4597 -7909 4609 -7875
rect 4609 -7909 4643 -7875
rect 4643 -7909 4655 -7875
rect 4597 -7915 4655 -7909
rect 4715 -7767 4773 -7761
rect 4715 -7801 4727 -7767
rect 4727 -7801 4761 -7767
rect 4761 -7801 4773 -7767
rect 4715 -7875 4773 -7801
rect 4715 -7909 4727 -7875
rect 4727 -7909 4761 -7875
rect 4761 -7909 4773 -7875
rect 4715 -7915 4773 -7909
rect 5061 -7767 5119 -7761
rect 5061 -7801 5073 -7767
rect 5073 -7801 5107 -7767
rect 5107 -7801 5119 -7767
rect 5061 -7875 5119 -7801
rect 5061 -7909 5073 -7875
rect 5073 -7909 5107 -7875
rect 5107 -7909 5119 -7875
rect 5061 -7915 5119 -7909
rect 5179 -7767 5237 -7761
rect 5179 -7801 5191 -7767
rect 5191 -7801 5225 -7767
rect 5225 -7801 5237 -7767
rect 5179 -7875 5237 -7801
rect 5179 -7909 5191 -7875
rect 5191 -7909 5225 -7875
rect 5225 -7909 5237 -7875
rect 5179 -7915 5237 -7909
rect 5297 -7767 5355 -7761
rect 5297 -7801 5309 -7767
rect 5309 -7801 5343 -7767
rect 5343 -7801 5355 -7767
rect 5297 -7875 5355 -7801
rect 5297 -7909 5309 -7875
rect 5309 -7909 5343 -7875
rect 5343 -7909 5355 -7875
rect 5297 -7915 5355 -7909
rect 5415 -7767 5473 -7761
rect 5415 -7801 5427 -7767
rect 5427 -7801 5461 -7767
rect 5461 -7801 5473 -7767
rect 5415 -7875 5473 -7801
rect 5415 -7909 5427 -7875
rect 5427 -7909 5461 -7875
rect 5461 -7909 5473 -7875
rect 5415 -7915 5473 -7909
rect 5533 -7767 5591 -7761
rect 5533 -7801 5545 -7767
rect 5545 -7801 5579 -7767
rect 5579 -7801 5591 -7767
rect 5533 -7875 5591 -7801
rect 5533 -7909 5545 -7875
rect 5545 -7909 5579 -7875
rect 5579 -7909 5591 -7875
rect 5533 -7915 5591 -7909
rect 5651 -7767 5709 -7761
rect 5651 -7801 5663 -7767
rect 5663 -7801 5697 -7767
rect 5697 -7801 5709 -7767
rect 5651 -7875 5709 -7801
rect 5651 -7909 5663 -7875
rect 5663 -7909 5697 -7875
rect 5697 -7909 5709 -7875
rect 5651 -7915 5709 -7909
rect 5769 -7767 5827 -7761
rect 5769 -7801 5781 -7767
rect 5781 -7801 5815 -7767
rect 5815 -7801 5827 -7767
rect 5769 -7875 5827 -7801
rect 5769 -7909 5781 -7875
rect 5781 -7909 5815 -7875
rect 5815 -7909 5827 -7875
rect 5769 -7915 5827 -7909
rect 5887 -7767 5945 -7761
rect 5887 -7801 5899 -7767
rect 5899 -7801 5933 -7767
rect 5933 -7801 5945 -7767
rect 5887 -7875 5945 -7801
rect 5887 -7909 5899 -7875
rect 5899 -7909 5933 -7875
rect 5933 -7909 5945 -7875
rect 5887 -7915 5945 -7909
rect 6005 -7767 6063 -7761
rect 6005 -7801 6017 -7767
rect 6017 -7801 6051 -7767
rect 6051 -7801 6063 -7767
rect 6005 -7875 6063 -7801
rect 6005 -7909 6017 -7875
rect 6017 -7909 6051 -7875
rect 6051 -7909 6063 -7875
rect 6005 -7915 6063 -7909
rect 6123 -7767 6181 -7761
rect 6123 -7801 6135 -7767
rect 6135 -7801 6169 -7767
rect 6169 -7801 6181 -7767
rect 6123 -7875 6181 -7801
rect 6123 -7909 6135 -7875
rect 6135 -7909 6169 -7875
rect 6169 -7909 6181 -7875
rect 6123 -7915 6181 -7909
rect 6241 -7767 6299 -7761
rect 6241 -7801 6253 -7767
rect 6253 -7801 6287 -7767
rect 6287 -7801 6299 -7767
rect 6241 -7875 6299 -7801
rect 6241 -7909 6253 -7875
rect 6253 -7909 6287 -7875
rect 6287 -7909 6299 -7875
rect 6241 -7915 6299 -7909
rect 6359 -7767 6417 -7761
rect 6359 -7801 6371 -7767
rect 6371 -7801 6405 -7767
rect 6405 -7801 6417 -7767
rect 6359 -7875 6417 -7801
rect 6359 -7909 6371 -7875
rect 6371 -7909 6405 -7875
rect 6405 -7909 6417 -7875
rect 6359 -7915 6417 -7909
rect 6477 -7767 6535 -7761
rect 6477 -7801 6489 -7767
rect 6489 -7801 6523 -7767
rect 6523 -7801 6535 -7767
rect 6477 -7875 6535 -7801
rect 6477 -7909 6489 -7875
rect 6489 -7909 6523 -7875
rect 6523 -7909 6535 -7875
rect 6477 -7915 6535 -7909
rect 6595 -7767 6653 -7761
rect 6595 -7801 6607 -7767
rect 6607 -7801 6641 -7767
rect 6641 -7801 6653 -7767
rect 6595 -7875 6653 -7801
rect 6595 -7909 6607 -7875
rect 6607 -7909 6641 -7875
rect 6641 -7909 6653 -7875
rect 6595 -7915 6653 -7909
rect 6713 -7767 6771 -7761
rect 6713 -7801 6725 -7767
rect 6725 -7801 6759 -7767
rect 6759 -7801 6771 -7767
rect 6713 -7875 6771 -7801
rect 6713 -7909 6725 -7875
rect 6725 -7909 6759 -7875
rect 6759 -7909 6771 -7875
rect 6713 -7915 6771 -7909
rect 11454 -8632 11463 -7792
rect 11463 -8632 11497 -7792
rect 11497 -8632 11506 -7792
rect 11602 -8632 11611 -7792
rect 11611 -8632 11645 -7792
rect 11645 -8632 11654 -7792
rect 11750 -8632 11759 -7792
rect 11759 -8632 11793 -7792
rect 11793 -8632 11802 -7792
rect 11898 -8632 11907 -7792
rect 11907 -8632 11941 -7792
rect 11941 -8632 11950 -7792
rect 12046 -8632 12055 -7792
rect 12055 -8632 12089 -7792
rect 12089 -8632 12098 -7792
rect 12194 -8632 12203 -7792
rect 12203 -8632 12237 -7792
rect 12237 -8632 12246 -7792
rect 12342 -8632 12351 -7792
rect 12351 -8632 12385 -7792
rect 12385 -8632 12394 -7792
rect 12490 -8632 12499 -7792
rect 12499 -8632 12533 -7792
rect 12533 -8632 12542 -7792
rect 12638 -8632 12690 -7792
rect 12786 -8632 12838 -7792
rect 12934 -8632 12986 -7792
rect 13082 -8632 13134 -7792
rect 13230 -8632 13239 -7792
rect 13239 -8632 13273 -7792
rect 13273 -8632 13282 -7792
rect 13378 -8632 13387 -7792
rect 13387 -8632 13421 -7792
rect 13421 -8632 13430 -7792
rect 13526 -8632 13535 -7792
rect 13535 -8632 13569 -7792
rect 13569 -8632 13578 -7792
rect 13674 -8632 13683 -7792
rect 13683 -8632 13717 -7792
rect 13717 -8632 13726 -7792
rect 13822 -8632 13831 -7792
rect 13831 -8632 13865 -7792
rect 13865 -8632 13874 -7792
rect 13970 -8632 13979 -7792
rect 13979 -8632 14013 -7792
rect 14013 -8632 14022 -7792
rect 14118 -8632 14127 -7792
rect 14127 -8632 14161 -7792
rect 14161 -8632 14170 -7792
rect 14266 -8632 14275 -7792
rect 14275 -8632 14309 -7792
rect 14309 -8632 14318 -7792
rect 14414 -8632 14466 -7792
rect 14562 -8632 14614 -7792
rect 14710 -8632 14762 -7792
rect 14858 -8632 14910 -7792
rect 15006 -8632 15058 -7792
rect 15154 -8632 15206 -7792
rect 15302 -8632 15354 -7792
rect 15450 -8632 15502 -7792
rect 15598 -8632 15607 -7792
rect 15607 -8632 15641 -7792
rect 15641 -8632 15650 -7792
rect 15746 -8632 15755 -7792
rect 15755 -8632 15789 -7792
rect 15789 -8632 15798 -7792
rect 15894 -8632 15903 -7792
rect 15903 -8632 15937 -7792
rect 15937 -8632 15946 -7792
rect 16042 -8632 16051 -7792
rect 16051 -8632 16085 -7792
rect 16085 -8632 16094 -7792
rect 16190 -8632 16199 -7792
rect 16199 -8632 16233 -7792
rect 16233 -8632 16242 -7792
rect 16338 -8632 16347 -7792
rect 16347 -8632 16381 -7792
rect 16381 -8632 16390 -7792
rect 16486 -8632 16495 -7792
rect 16495 -8632 16529 -7792
rect 16529 -8632 16538 -7792
rect 16634 -8632 16643 -7792
rect 16643 -8632 16677 -7792
rect 16677 -8632 16686 -7792
rect 16782 -8632 16834 -7792
rect 16930 -8632 16982 -7792
rect 17078 -8632 17130 -7792
rect 17226 -8632 17278 -7792
rect 17374 -8632 17426 -7792
rect 17522 -8632 17574 -7792
rect 17670 -8632 17722 -7792
rect 17818 -8632 17870 -7792
rect 17966 -8632 17975 -7792
rect 17975 -8632 18009 -7792
rect 18009 -8632 18018 -7792
rect 18114 -8632 18123 -7792
rect 18123 -8632 18157 -7792
rect 18157 -8632 18166 -7792
rect 18262 -8632 18271 -7792
rect 18271 -8632 18305 -7792
rect 18305 -8632 18314 -7792
rect 18410 -8632 18419 -7792
rect 18419 -8632 18453 -7792
rect 18453 -8632 18462 -7792
rect 18558 -8632 18567 -7792
rect 18567 -8632 18601 -7792
rect 18601 -8632 18610 -7792
rect 18706 -8632 18715 -7792
rect 18715 -8632 18749 -7792
rect 18749 -8632 18758 -7792
rect 18854 -8632 18863 -7792
rect 18863 -8632 18897 -7792
rect 18897 -8632 18906 -7792
rect 19002 -8632 19011 -7792
rect 19011 -8632 19045 -7792
rect 19045 -8632 19054 -7792
rect 19150 -8632 19202 -7792
rect 19298 -8632 19350 -7792
rect 19446 -8632 19498 -7792
rect 19594 -8632 19646 -7792
rect 19742 -8632 19794 -7792
rect 19890 -8632 19942 -7792
rect 20038 -8632 20090 -7792
rect 20186 -8632 20238 -7792
rect 20334 -8632 20343 -7792
rect 20343 -8632 20377 -7792
rect 20377 -8632 20386 -7792
rect 20482 -8632 20491 -7792
rect 20491 -8632 20525 -7792
rect 20525 -8632 20534 -7792
rect 20630 -8632 20639 -7792
rect 20639 -8632 20673 -7792
rect 20673 -8632 20682 -7792
rect 20778 -8632 20787 -7792
rect 20787 -8632 20821 -7792
rect 20821 -8632 20830 -7792
rect 20926 -8632 20935 -7792
rect 20935 -8632 20969 -7792
rect 20969 -8632 20978 -7792
rect 21074 -8632 21083 -7792
rect 21083 -8632 21117 -7792
rect 21117 -8632 21126 -7792
rect 21222 -8632 21231 -7792
rect 21231 -8632 21265 -7792
rect 21265 -8632 21274 -7792
rect 21370 -8632 21379 -7792
rect 21379 -8632 21413 -7792
rect 21413 -8632 21422 -7792
rect 21518 -8632 21570 -7792
rect 21666 -8632 21718 -7792
rect 21814 -8632 21866 -7792
rect 21962 -8632 22014 -7792
rect 22110 -8632 22162 -7792
rect 22258 -8632 22310 -7792
rect 22406 -8632 22458 -7792
rect 22554 -8632 22606 -7792
rect 22830 -7926 22882 -7086
rect 23055 -7926 23107 -7086
rect 23233 -7939 23285 -7099
<< metal2 >>
rect 6530 2687 6582 2697
rect 6530 2077 6582 2087
rect 6766 2687 6818 2697
rect 6766 2077 6818 2087
rect 4482 2045 21337 2054
rect 4482 2044 12547 2045
rect 4482 1952 4601 2044
rect 4659 1952 4719 2044
rect 4777 1952 4837 2044
rect 4895 1952 4955 2044
rect 5013 1952 5073 2044
rect 5131 1952 5191 2044
rect 5249 1952 5309 2044
rect 5367 1952 5427 2044
rect 5485 1952 5545 2044
rect 5603 1952 5663 2044
rect 5721 1952 5781 2044
rect 5839 1952 5899 2044
rect 5957 1952 6017 2044
rect 6075 1952 6135 2044
rect 6193 1952 6253 2044
rect 6311 1952 6599 2044
rect 6657 1952 6717 2044
rect 6775 1952 6835 2044
rect 6893 1952 6953 2044
rect 7011 1952 7071 2044
rect 7129 1952 7189 2044
rect 7247 1952 7307 2044
rect 7365 1952 7425 2044
rect 7483 1952 7543 2044
rect 7601 1952 7661 2044
rect 7719 1952 7779 2044
rect 7837 1952 7897 2044
rect 7955 1952 8015 2044
rect 8073 1952 8133 2044
rect 8191 1952 8251 2044
rect 8309 1952 8597 2044
rect 8655 1952 8715 2044
rect 8773 1952 8833 2044
rect 8891 1952 8951 2044
rect 9009 1952 9069 2044
rect 9127 1952 9187 2044
rect 9245 1952 9305 2044
rect 9363 1952 9423 2044
rect 9481 1952 9541 2044
rect 9599 1952 9659 2044
rect 9717 1952 9777 2044
rect 9835 1952 9895 2044
rect 9953 1952 10013 2044
rect 10071 1952 10131 2044
rect 10189 1952 10249 2044
rect 10307 1952 12547 2044
rect 4482 1942 12547 1952
rect 12324 1891 12547 1942
rect 12605 1891 12665 2045
rect 12723 1891 12783 2045
rect 12841 1891 12901 2045
rect 12959 1891 13019 2045
rect 13077 1891 13137 2045
rect 13195 1891 13255 2045
rect 13313 1891 13373 2045
rect 13431 1891 13491 2045
rect 13549 1891 13609 2045
rect 13667 1891 13727 2045
rect 13785 1891 13845 2045
rect 13903 1891 13963 2045
rect 14021 1891 14081 2045
rect 14139 1891 14199 2045
rect 14257 1891 14317 2045
rect 14375 1891 14435 2045
rect 14493 1891 14553 2045
rect 14611 1891 14671 2045
rect 14729 1891 14789 2045
rect 14847 1891 14907 2045
rect 14965 1891 15025 2045
rect 15083 1891 15143 2045
rect 15201 1891 15261 2045
rect 15319 1891 15379 2045
rect 15437 1891 15497 2045
rect 15555 1891 15615 2045
rect 15673 1891 15733 2045
rect 15791 1891 15851 2045
rect 15909 1891 15969 2045
rect 16027 1891 16087 2045
rect 16145 1891 16205 2045
rect 16263 1891 16323 2045
rect 16381 1891 16441 2045
rect 16499 1891 16559 2045
rect 16617 1891 16677 2045
rect 16735 1891 16795 2045
rect 16853 1891 16913 2045
rect 16971 1891 17031 2045
rect 17089 1891 17149 2045
rect 17207 1891 17267 2045
rect 17325 1891 17385 2045
rect 17443 1891 17503 2045
rect 17561 1891 17621 2045
rect 17679 1891 17739 2045
rect 17797 1891 17857 2045
rect 17915 1891 17975 2045
rect 18033 1891 18093 2045
rect 18151 1891 18211 2045
rect 18269 1891 18329 2045
rect 18387 1891 18447 2045
rect 18505 1891 18565 2045
rect 18623 1891 18683 2045
rect 18741 1891 18801 2045
rect 18859 1891 18919 2045
rect 18977 1891 19037 2045
rect 19095 1891 19155 2045
rect 19213 1891 19273 2045
rect 19331 1891 19391 2045
rect 19449 1891 19509 2045
rect 19567 1891 19627 2045
rect 19685 1891 19745 2045
rect 19803 1891 19863 2045
rect 19921 1891 19981 2045
rect 20039 1891 20099 2045
rect 20157 1891 20217 2045
rect 20275 1891 20335 2045
rect 20393 1891 20453 2045
rect 20511 1891 20571 2045
rect 20629 1891 20689 2045
rect 20747 1891 20807 2045
rect 20865 1891 20925 2045
rect 20983 1891 21043 2045
rect 21101 1891 21161 2045
rect 21219 1891 21279 2045
rect 12324 1881 21337 1891
rect 1337 -142 7177 -132
rect 1395 -296 1455 -142
rect 1513 -296 1573 -142
rect 1631 -296 1691 -142
rect 1749 -296 1809 -142
rect 1867 -296 1927 -142
rect 1985 -296 2045 -142
rect 2103 -296 2163 -142
rect 2221 -296 2281 -142
rect 2339 -296 2399 -142
rect 2457 -296 2517 -142
rect 2575 -296 2635 -142
rect 2693 -296 2753 -142
rect 2811 -296 2871 -142
rect 2929 -296 2989 -142
rect 3047 -296 3107 -142
rect 3165 -296 3225 -142
rect 3283 -296 3343 -142
rect 3401 -296 3461 -142
rect 3519 -296 3579 -142
rect 3637 -296 3697 -142
rect 3755 -296 3815 -142
rect 3873 -296 3933 -142
rect 3991 -296 4051 -142
rect 4109 -296 4169 -142
rect 4227 -296 4287 -142
rect 4345 -296 4405 -142
rect 4463 -296 4523 -142
rect 4581 -296 4641 -142
rect 4699 -296 4759 -142
rect 4817 -296 4877 -142
rect 4935 -296 4995 -142
rect 5053 -296 5113 -142
rect 5171 -296 5231 -142
rect 5289 -296 5349 -142
rect 5407 -296 5467 -142
rect 5525 -296 5585 -142
rect 5643 -296 5703 -142
rect 5761 -296 5821 -142
rect 5879 -296 5939 -142
rect 5997 -296 6057 -142
rect 6115 -296 6175 -142
rect 6233 -296 6293 -142
rect 6351 -296 6411 -142
rect 6469 -296 6529 -142
rect 6587 -296 6647 -142
rect 6705 -296 6765 -142
rect 6823 -296 6883 -142
rect 6941 -296 7001 -142
rect 7059 -296 7119 -142
rect 1337 -306 7177 -296
rect 1337 -1910 7177 -1900
rect 1395 -2064 1455 -1910
rect 1513 -2064 1573 -1910
rect 1631 -2064 1691 -1910
rect 1749 -2064 1809 -1910
rect 1867 -2064 1927 -1910
rect 1985 -2064 2045 -1910
rect 2103 -2064 2163 -1910
rect 2221 -2064 2281 -1910
rect 2339 -2064 2399 -1910
rect 2457 -2064 2517 -1910
rect 2575 -2064 2635 -1910
rect 2693 -2064 2753 -1910
rect 2811 -2064 2871 -1910
rect 2929 -2064 2989 -1910
rect 3047 -2064 3107 -1910
rect 3165 -2064 3225 -1910
rect 3283 -2064 3343 -1910
rect 3401 -2064 3461 -1910
rect 3519 -2064 3579 -1910
rect 3637 -2064 3697 -1910
rect 3755 -2064 3815 -1910
rect 3873 -2064 3933 -1910
rect 3991 -2064 4051 -1910
rect 4109 -2064 4169 -1910
rect 4227 -2064 4287 -1910
rect 4345 -2064 4405 -1910
rect 4463 -2064 4523 -1910
rect 4581 -2064 4641 -1910
rect 4699 -2064 4759 -1910
rect 4817 -2064 4877 -1910
rect 4935 -2064 4995 -1910
rect 5053 -2064 5113 -1910
rect 5171 -2064 5231 -1910
rect 5289 -2064 5349 -1910
rect 5407 -2064 5467 -1910
rect 5525 -2064 5585 -1910
rect 5643 -2064 5703 -1910
rect 5761 -2064 5821 -1910
rect 5879 -2064 5939 -1910
rect 5997 -2064 6057 -1910
rect 6115 -2064 6175 -1910
rect 6233 -2064 6293 -1910
rect 6351 -2064 6411 -1910
rect 6469 -2064 6529 -1910
rect 6587 -2064 6647 -1910
rect 6705 -2064 6765 -1910
rect 6823 -2064 6883 -1910
rect 6941 -2064 7001 -1910
rect 7059 -2064 7119 -1910
rect 1337 -2074 7177 -2064
rect 1337 -3678 7177 -3668
rect 1395 -3832 1455 -3678
rect 1513 -3832 1573 -3678
rect 1631 -3832 1691 -3678
rect 1749 -3832 1809 -3678
rect 1867 -3832 1927 -3678
rect 1985 -3832 2045 -3678
rect 2103 -3832 2163 -3678
rect 2221 -3832 2281 -3678
rect 2339 -3832 2399 -3678
rect 2457 -3832 2517 -3678
rect 2575 -3832 2635 -3678
rect 2693 -3832 2753 -3678
rect 2811 -3832 2871 -3678
rect 2929 -3832 2989 -3678
rect 3047 -3832 3107 -3678
rect 3165 -3832 3225 -3678
rect 3283 -3832 3343 -3678
rect 3401 -3832 3461 -3678
rect 3519 -3832 3579 -3678
rect 3637 -3832 3697 -3678
rect 3755 -3832 3815 -3678
rect 3873 -3832 3933 -3678
rect 3991 -3832 4051 -3678
rect 4109 -3832 4169 -3678
rect 4227 -3832 4287 -3678
rect 4345 -3832 4405 -3678
rect 4463 -3832 4523 -3678
rect 4581 -3832 4641 -3678
rect 4699 -3832 4759 -3678
rect 4817 -3832 4877 -3678
rect 4935 -3832 4995 -3678
rect 5053 -3832 5113 -3678
rect 5171 -3832 5231 -3678
rect 5289 -3832 5349 -3678
rect 5407 -3832 5467 -3678
rect 5525 -3832 5585 -3678
rect 5643 -3832 5703 -3678
rect 5761 -3832 5821 -3678
rect 5879 -3832 5939 -3678
rect 5997 -3832 6057 -3678
rect 6115 -3832 6175 -3678
rect 6233 -3832 6293 -3678
rect 6351 -3832 6411 -3678
rect 6469 -3832 6529 -3678
rect 6587 -3832 6647 -3678
rect 6705 -3832 6765 -3678
rect 6823 -3832 6883 -3678
rect 6941 -3832 7001 -3678
rect 7059 -3832 7119 -3678
rect 1337 -3842 7177 -3832
rect 1337 -5446 7177 -5436
rect 1395 -5600 1455 -5446
rect 1513 -5600 1573 -5446
rect 1631 -5600 1691 -5446
rect 1749 -5600 1809 -5446
rect 1867 -5600 1927 -5446
rect 1985 -5600 2045 -5446
rect 2103 -5600 2163 -5446
rect 2221 -5600 2281 -5446
rect 2339 -5600 2399 -5446
rect 2457 -5600 2517 -5446
rect 2575 -5600 2635 -5446
rect 2693 -5600 2753 -5446
rect 2811 -5600 2871 -5446
rect 2929 -5600 2989 -5446
rect 3047 -5600 3107 -5446
rect 3165 -5600 3225 -5446
rect 3283 -5600 3343 -5446
rect 3401 -5600 3461 -5446
rect 3519 -5600 3579 -5446
rect 3637 -5600 3697 -5446
rect 3755 -5600 3815 -5446
rect 3873 -5600 3933 -5446
rect 3991 -5600 4051 -5446
rect 4109 -5600 4169 -5446
rect 4227 -5600 4287 -5446
rect 4345 -5600 4405 -5446
rect 4463 -5600 4523 -5446
rect 4581 -5600 4641 -5446
rect 4699 -5600 4759 -5446
rect 4817 -5600 4877 -5446
rect 4935 -5600 4995 -5446
rect 5053 -5600 5113 -5446
rect 5171 -5600 5231 -5446
rect 5289 -5600 5349 -5446
rect 5407 -5600 5467 -5446
rect 5525 -5600 5585 -5446
rect 5643 -5600 5703 -5446
rect 5761 -5600 5821 -5446
rect 5879 -5600 5939 -5446
rect 5997 -5600 6057 -5446
rect 6115 -5600 6175 -5446
rect 6233 -5600 6293 -5446
rect 6351 -5600 6411 -5446
rect 6469 -5600 6529 -5446
rect 6587 -5600 6647 -5446
rect 6705 -5600 6765 -5446
rect 6823 -5600 6883 -5446
rect 6941 -5600 7001 -5446
rect 7059 -5600 7119 -5446
rect 1337 -5610 7177 -5600
rect 11452 -6646 11508 -6636
rect 11452 -7496 11508 -7486
rect 11600 -6646 11656 -6636
rect 11600 -7496 11656 -7486
rect 11748 -6646 11804 -6636
rect 11748 -7496 11804 -7486
rect 11896 -6646 11952 -6636
rect 11896 -7496 11952 -7486
rect 12044 -6646 12100 -6636
rect 12044 -7496 12100 -7486
rect 12192 -6646 12248 -6636
rect 12192 -7496 12248 -7486
rect 12340 -6646 12396 -6636
rect 12340 -7496 12396 -7486
rect 12488 -6646 12544 -6636
rect 12488 -7496 12544 -7486
rect 12636 -6646 12692 -6636
rect 12636 -7496 12692 -7486
rect 12784 -6646 12840 -6636
rect 12784 -7496 12840 -7486
rect 12932 -6646 12988 -6636
rect 12932 -7496 12988 -7486
rect 13080 -6646 13136 -6636
rect 13080 -7496 13136 -7486
rect 13228 -6646 13284 -6636
rect 13228 -7496 13284 -7486
rect 13376 -6646 13432 -6636
rect 13376 -7496 13432 -7486
rect 13524 -6646 13580 -6636
rect 13524 -7496 13580 -7486
rect 13672 -6646 13728 -6636
rect 13672 -7496 13728 -7486
rect 13820 -6646 13876 -6636
rect 13820 -7496 13876 -7486
rect 13968 -6646 14024 -6636
rect 13968 -7496 14024 -7486
rect 14116 -6646 14172 -6636
rect 14116 -7496 14172 -7486
rect 14264 -6646 14320 -6636
rect 14264 -7496 14320 -7486
rect 14412 -6646 14468 -6636
rect 14412 -7496 14468 -7486
rect 14560 -6646 14616 -6636
rect 14560 -7496 14616 -7486
rect 14708 -6646 14764 -6636
rect 14708 -7496 14764 -7486
rect 14856 -6646 14912 -6636
rect 14856 -7496 14912 -7486
rect 15004 -6646 15060 -6636
rect 15004 -7496 15060 -7486
rect 15152 -6646 15208 -6636
rect 15152 -7496 15208 -7486
rect 15300 -6646 15356 -6636
rect 15300 -7496 15356 -7486
rect 15448 -6646 15504 -6636
rect 15448 -7496 15504 -7486
rect 15596 -6646 15652 -6636
rect 15596 -7496 15652 -7486
rect 15744 -6646 15800 -6636
rect 15744 -7496 15800 -7486
rect 15892 -6646 15948 -6636
rect 15892 -7496 15948 -7486
rect 16040 -6646 16096 -6636
rect 16040 -7496 16096 -7486
rect 16188 -6646 16244 -6636
rect 16188 -7496 16244 -7486
rect 16336 -6646 16392 -6636
rect 16336 -7496 16392 -7486
rect 16484 -6646 16540 -6636
rect 16484 -7496 16540 -7486
rect 16632 -6646 16688 -6636
rect 16632 -7496 16688 -7486
rect 16780 -6646 16836 -6636
rect 16780 -7496 16836 -7486
rect 16928 -6646 16984 -6636
rect 16928 -7496 16984 -7486
rect 17076 -6646 17132 -6636
rect 17076 -7496 17132 -7486
rect 17224 -6646 17280 -6636
rect 17224 -7496 17280 -7486
rect 17372 -6646 17428 -6636
rect 17372 -7496 17428 -7486
rect 17520 -6646 17576 -6636
rect 17520 -7496 17576 -7486
rect 17668 -6646 17724 -6636
rect 17668 -7496 17724 -7486
rect 17816 -6646 17872 -6636
rect 17816 -7496 17872 -7486
rect 17964 -6646 18020 -6636
rect 17964 -7496 18020 -7486
rect 18112 -6646 18168 -6636
rect 18112 -7496 18168 -7486
rect 18260 -6646 18316 -6636
rect 18260 -7496 18316 -7486
rect 18408 -6646 18464 -6636
rect 18408 -7496 18464 -7486
rect 18556 -6646 18612 -6636
rect 18556 -7496 18612 -7486
rect 18704 -6646 18760 -6636
rect 18704 -7496 18760 -7486
rect 18852 -6646 18908 -6636
rect 18852 -7496 18908 -7486
rect 19000 -6646 19056 -6636
rect 19000 -7496 19056 -7486
rect 19148 -6646 19204 -6636
rect 19148 -7496 19204 -7486
rect 19296 -6646 19352 -6636
rect 19296 -7496 19352 -7486
rect 19444 -6646 19500 -6636
rect 19444 -7496 19500 -7486
rect 19592 -6646 19648 -6636
rect 19592 -7496 19648 -7486
rect 19740 -6646 19796 -6636
rect 19740 -7496 19796 -7486
rect 19888 -6646 19944 -6636
rect 19888 -7496 19944 -7486
rect 20036 -6646 20092 -6636
rect 20036 -7496 20092 -7486
rect 20184 -6646 20240 -6636
rect 20184 -7496 20240 -7486
rect 20332 -6646 20388 -6636
rect 20332 -7496 20388 -7486
rect 20480 -6646 20536 -6636
rect 20480 -7496 20536 -7486
rect 20628 -6646 20684 -6636
rect 20628 -7496 20684 -7486
rect 20776 -6646 20832 -6636
rect 20776 -7496 20832 -7486
rect 20924 -6646 20980 -6636
rect 20924 -7496 20980 -7486
rect 21072 -6646 21128 -6636
rect 21072 -7496 21128 -7486
rect 21220 -6646 21276 -6636
rect 21220 -7496 21276 -7486
rect 21368 -6646 21424 -6636
rect 21368 -7496 21424 -7486
rect 21516 -6646 21572 -6636
rect 21516 -7496 21572 -7486
rect 21664 -6646 21720 -6636
rect 21664 -7496 21720 -7486
rect 21812 -6646 21868 -6636
rect 21812 -7496 21868 -7486
rect 21960 -6646 22016 -6636
rect 21960 -7496 22016 -7486
rect 22108 -6646 22164 -6636
rect 22108 -7496 22164 -7486
rect 22256 -6646 22312 -6636
rect 22256 -7496 22312 -7486
rect 22404 -6646 22460 -6636
rect 22404 -7496 22460 -7486
rect 22552 -6646 22608 -6636
rect 22552 -7496 22608 -7486
rect 22830 -7086 22882 -7076
rect 11509 -7562 22561 -7552
rect 11599 -7716 11657 -7562
rect 11747 -7716 11805 -7562
rect 11895 -7716 11953 -7562
rect 12043 -7716 12101 -7562
rect 12191 -7716 12249 -7562
rect 12339 -7716 12397 -7562
rect 12487 -7716 12545 -7562
rect 12635 -7716 12693 -7562
rect 12783 -7716 12841 -7562
rect 12931 -7716 12989 -7562
rect 13079 -7716 13137 -7562
rect 13227 -7716 13285 -7562
rect 13375 -7716 13433 -7562
rect 13523 -7716 13581 -7562
rect 13671 -7716 13729 -7562
rect 13819 -7716 13877 -7562
rect 13967 -7716 14025 -7562
rect 14115 -7716 14173 -7562
rect 14263 -7716 14321 -7562
rect 14411 -7716 14469 -7562
rect 14559 -7716 14617 -7562
rect 14707 -7716 14765 -7562
rect 14855 -7716 14913 -7562
rect 15003 -7716 15061 -7562
rect 15151 -7716 15209 -7562
rect 15299 -7716 15357 -7562
rect 15447 -7716 15505 -7562
rect 15595 -7716 15653 -7562
rect 15743 -7716 15801 -7562
rect 15891 -7716 15949 -7562
rect 16039 -7716 16097 -7562
rect 16187 -7716 16245 -7562
rect 16335 -7716 16393 -7562
rect 16483 -7716 16541 -7562
rect 16631 -7716 16689 -7562
rect 16779 -7716 16837 -7562
rect 16927 -7716 16985 -7562
rect 17075 -7716 17133 -7562
rect 17223 -7716 17281 -7562
rect 17371 -7716 17429 -7562
rect 17519 -7716 17577 -7562
rect 17667 -7716 17725 -7562
rect 17815 -7716 17873 -7562
rect 17963 -7716 18021 -7562
rect 18111 -7716 18169 -7562
rect 18259 -7716 18317 -7562
rect 18407 -7716 18465 -7562
rect 18555 -7716 18613 -7562
rect 18703 -7716 18761 -7562
rect 18851 -7716 18909 -7562
rect 18999 -7716 19057 -7562
rect 19147 -7716 19205 -7562
rect 19295 -7716 19353 -7562
rect 19443 -7716 19501 -7562
rect 19591 -7716 19649 -7562
rect 19739 -7716 19797 -7562
rect 19887 -7716 19945 -7562
rect 20035 -7716 20093 -7562
rect 20183 -7716 20241 -7562
rect 20331 -7716 20389 -7562
rect 20479 -7716 20537 -7562
rect 20627 -7716 20685 -7562
rect 20775 -7716 20833 -7562
rect 20923 -7716 20981 -7562
rect 21071 -7716 21129 -7562
rect 21219 -7716 21277 -7562
rect 21367 -7716 21425 -7562
rect 21515 -7716 21573 -7562
rect 21663 -7716 21721 -7562
rect 21811 -7716 21869 -7562
rect 21959 -7716 22017 -7562
rect 22107 -7716 22165 -7562
rect 22255 -7716 22313 -7562
rect 22403 -7716 22461 -7562
rect 22551 -7716 22561 -7562
rect 11509 -7726 22561 -7716
rect 3063 -7761 6818 -7751
rect 3121 -7915 3181 -7761
rect 3239 -7915 3299 -7761
rect 3357 -7915 3417 -7761
rect 3475 -7915 3535 -7761
rect 3593 -7915 3653 -7761
rect 3711 -7915 3771 -7761
rect 3829 -7915 3889 -7761
rect 3947 -7915 4007 -7761
rect 4065 -7915 4125 -7761
rect 4183 -7915 4243 -7761
rect 4301 -7915 4361 -7761
rect 4419 -7915 4479 -7761
rect 4537 -7915 4597 -7761
rect 4655 -7915 4715 -7761
rect 4773 -7915 5061 -7761
rect 5119 -7915 5179 -7761
rect 5237 -7915 5297 -7761
rect 5355 -7915 5415 -7761
rect 5473 -7915 5533 -7761
rect 5591 -7915 5651 -7761
rect 5709 -7915 5769 -7761
rect 5827 -7915 5887 -7761
rect 5945 -7915 6005 -7761
rect 6063 -7915 6123 -7761
rect 6181 -7915 6241 -7761
rect 6299 -7915 6359 -7761
rect 6417 -7915 6477 -7761
rect 6535 -7915 6595 -7761
rect 6653 -7915 6713 -7761
rect 6771 -7915 6818 -7761
rect 3063 -7925 6818 -7915
rect 11452 -7792 11508 -7782
rect 11452 -8642 11508 -8632
rect 11600 -7792 11656 -7782
rect 11600 -8642 11656 -8632
rect 11748 -7792 11804 -7782
rect 11748 -8642 11804 -8632
rect 11896 -7792 11952 -7782
rect 11896 -8642 11952 -8632
rect 12044 -7792 12100 -7782
rect 12044 -8642 12100 -8632
rect 12192 -7792 12248 -7782
rect 12192 -8642 12248 -8632
rect 12340 -7792 12396 -7782
rect 12340 -8642 12396 -8632
rect 12488 -7792 12544 -7782
rect 12488 -8642 12544 -8632
rect 12636 -7792 12692 -7782
rect 12636 -8642 12692 -8632
rect 12784 -7792 12840 -7782
rect 12784 -8642 12840 -8632
rect 12932 -7792 12988 -7782
rect 12932 -8642 12988 -8632
rect 13080 -7792 13136 -7782
rect 13080 -8642 13136 -8632
rect 13228 -7792 13284 -7782
rect 13228 -8642 13284 -8632
rect 13376 -7792 13432 -7782
rect 13376 -8642 13432 -8632
rect 13524 -7792 13580 -7782
rect 13524 -8642 13580 -8632
rect 13672 -7792 13728 -7782
rect 13672 -8642 13728 -8632
rect 13820 -7792 13876 -7782
rect 13820 -8642 13876 -8632
rect 13968 -7792 14024 -7782
rect 13968 -8642 14024 -8632
rect 14116 -7792 14172 -7782
rect 14116 -8642 14172 -8632
rect 14264 -7792 14320 -7782
rect 14264 -8642 14320 -8632
rect 14412 -7792 14468 -7782
rect 14412 -8642 14468 -8632
rect 14560 -7792 14616 -7782
rect 14560 -8642 14616 -8632
rect 14708 -7792 14764 -7782
rect 14708 -8642 14764 -8632
rect 14856 -7792 14912 -7782
rect 14856 -8642 14912 -8632
rect 15004 -7792 15060 -7782
rect 15004 -8642 15060 -8632
rect 15152 -7792 15208 -7782
rect 15152 -8642 15208 -8632
rect 15300 -7792 15356 -7782
rect 15300 -8642 15356 -8632
rect 15448 -7792 15504 -7782
rect 15448 -8642 15504 -8632
rect 15596 -7792 15652 -7782
rect 15596 -8642 15652 -8632
rect 15744 -7792 15800 -7782
rect 15744 -8642 15800 -8632
rect 15892 -7792 15948 -7782
rect 15892 -8642 15948 -8632
rect 16040 -7792 16096 -7782
rect 16040 -8642 16096 -8632
rect 16188 -7792 16244 -7782
rect 16188 -8642 16244 -8632
rect 16336 -7792 16392 -7782
rect 16336 -8642 16392 -8632
rect 16484 -7792 16540 -7782
rect 16484 -8642 16540 -8632
rect 16632 -7792 16688 -7782
rect 16632 -8642 16688 -8632
rect 16780 -7792 16836 -7782
rect 16780 -8642 16836 -8632
rect 16928 -7792 16984 -7782
rect 16928 -8642 16984 -8632
rect 17076 -7792 17132 -7782
rect 17076 -8642 17132 -8632
rect 17224 -7792 17280 -7782
rect 17224 -8642 17280 -8632
rect 17372 -7792 17428 -7782
rect 17372 -8642 17428 -8632
rect 17520 -7792 17576 -7782
rect 17520 -8642 17576 -8632
rect 17668 -7792 17724 -7782
rect 17668 -8642 17724 -8632
rect 17816 -7792 17872 -7782
rect 17816 -8642 17872 -8632
rect 17964 -7792 18020 -7782
rect 17964 -8642 18020 -8632
rect 18112 -7792 18168 -7782
rect 18112 -8642 18168 -8632
rect 18260 -7792 18316 -7782
rect 18260 -8642 18316 -8632
rect 18408 -7792 18464 -7782
rect 18408 -8642 18464 -8632
rect 18556 -7792 18612 -7782
rect 18556 -8642 18612 -8632
rect 18704 -7792 18760 -7782
rect 18704 -8642 18760 -8632
rect 18852 -7792 18908 -7782
rect 18852 -8642 18908 -8632
rect 19000 -7792 19056 -7782
rect 19000 -8642 19056 -8632
rect 19148 -7792 19204 -7782
rect 19148 -8642 19204 -8632
rect 19296 -7792 19352 -7782
rect 19296 -8642 19352 -8632
rect 19444 -7792 19500 -7782
rect 19444 -8642 19500 -8632
rect 19592 -7792 19648 -7782
rect 19592 -8642 19648 -8632
rect 19740 -7792 19796 -7782
rect 19740 -8642 19796 -8632
rect 19888 -7792 19944 -7782
rect 19888 -8642 19944 -8632
rect 20036 -7792 20092 -7782
rect 20036 -8642 20092 -8632
rect 20184 -7792 20240 -7782
rect 20184 -8642 20240 -8632
rect 20332 -7792 20388 -7782
rect 20332 -8642 20388 -8632
rect 20480 -7792 20536 -7782
rect 20480 -8642 20536 -8632
rect 20628 -7792 20684 -7782
rect 20628 -8642 20684 -8632
rect 20776 -7792 20832 -7782
rect 20776 -8642 20832 -8632
rect 20924 -7792 20980 -7782
rect 20924 -8642 20980 -8632
rect 21072 -7792 21128 -7782
rect 21072 -8642 21128 -8632
rect 21220 -7792 21276 -7782
rect 21220 -8642 21276 -8632
rect 21368 -7792 21424 -7782
rect 21368 -8642 21424 -8632
rect 21516 -7792 21572 -7782
rect 21516 -8642 21572 -8632
rect 21664 -7792 21720 -7782
rect 21664 -8642 21720 -8632
rect 21812 -7792 21868 -7782
rect 21812 -8642 21868 -8632
rect 21960 -7792 22016 -7782
rect 21960 -8642 22016 -8632
rect 22108 -7792 22164 -7782
rect 22108 -8642 22164 -8632
rect 22256 -7792 22312 -7782
rect 22256 -8642 22312 -8632
rect 22404 -7792 22460 -7782
rect 22404 -8642 22460 -8632
rect 22552 -7792 22608 -7782
rect 22830 -7936 22882 -7926
rect 23053 -7086 23109 -7076
rect 23053 -7936 23109 -7926
rect 23231 -7099 23287 -7089
rect 23231 -7949 23287 -7939
rect 22552 -8642 22608 -8632
<< via2 >>
rect 11452 -7486 11454 -6646
rect 11454 -7486 11506 -6646
rect 11506 -7486 11508 -6646
rect 11600 -7486 11602 -6646
rect 11602 -7486 11654 -6646
rect 11654 -7486 11656 -6646
rect 11748 -7486 11750 -6646
rect 11750 -7486 11802 -6646
rect 11802 -7486 11804 -6646
rect 11896 -7486 11898 -6646
rect 11898 -7486 11950 -6646
rect 11950 -7486 11952 -6646
rect 12044 -7486 12046 -6646
rect 12046 -7486 12098 -6646
rect 12098 -7486 12100 -6646
rect 12192 -7486 12194 -6646
rect 12194 -7486 12246 -6646
rect 12246 -7486 12248 -6646
rect 12340 -7486 12342 -6646
rect 12342 -7486 12394 -6646
rect 12394 -7486 12396 -6646
rect 12488 -7486 12490 -6646
rect 12490 -7486 12542 -6646
rect 12542 -7486 12544 -6646
rect 12636 -7486 12638 -6646
rect 12638 -7486 12690 -6646
rect 12690 -7486 12692 -6646
rect 12784 -7486 12786 -6646
rect 12786 -7486 12838 -6646
rect 12838 -7486 12840 -6646
rect 12932 -7486 12934 -6646
rect 12934 -7486 12986 -6646
rect 12986 -7486 12988 -6646
rect 13080 -7486 13082 -6646
rect 13082 -7486 13134 -6646
rect 13134 -7486 13136 -6646
rect 13228 -7486 13230 -6646
rect 13230 -7486 13282 -6646
rect 13282 -7486 13284 -6646
rect 13376 -7486 13378 -6646
rect 13378 -7486 13430 -6646
rect 13430 -7486 13432 -6646
rect 13524 -7486 13526 -6646
rect 13526 -7486 13578 -6646
rect 13578 -7486 13580 -6646
rect 13672 -7486 13674 -6646
rect 13674 -7486 13726 -6646
rect 13726 -7486 13728 -6646
rect 13820 -7486 13822 -6646
rect 13822 -7486 13874 -6646
rect 13874 -7486 13876 -6646
rect 13968 -7486 13970 -6646
rect 13970 -7486 14022 -6646
rect 14022 -7486 14024 -6646
rect 14116 -7486 14118 -6646
rect 14118 -7486 14170 -6646
rect 14170 -7486 14172 -6646
rect 14264 -7486 14266 -6646
rect 14266 -7486 14318 -6646
rect 14318 -7486 14320 -6646
rect 14412 -7486 14414 -6646
rect 14414 -7486 14466 -6646
rect 14466 -7486 14468 -6646
rect 14560 -7486 14562 -6646
rect 14562 -7486 14614 -6646
rect 14614 -7486 14616 -6646
rect 14708 -7486 14710 -6646
rect 14710 -7486 14762 -6646
rect 14762 -7486 14764 -6646
rect 14856 -7486 14858 -6646
rect 14858 -7486 14910 -6646
rect 14910 -7486 14912 -6646
rect 15004 -7486 15006 -6646
rect 15006 -7486 15058 -6646
rect 15058 -7486 15060 -6646
rect 15152 -7486 15154 -6646
rect 15154 -7486 15206 -6646
rect 15206 -7486 15208 -6646
rect 15300 -7486 15302 -6646
rect 15302 -7486 15354 -6646
rect 15354 -7486 15356 -6646
rect 15448 -7486 15450 -6646
rect 15450 -7486 15502 -6646
rect 15502 -7486 15504 -6646
rect 15596 -7486 15598 -6646
rect 15598 -7486 15650 -6646
rect 15650 -7486 15652 -6646
rect 15744 -7486 15746 -6646
rect 15746 -7486 15798 -6646
rect 15798 -7486 15800 -6646
rect 15892 -7486 15894 -6646
rect 15894 -7486 15946 -6646
rect 15946 -7486 15948 -6646
rect 16040 -7486 16042 -6646
rect 16042 -7486 16094 -6646
rect 16094 -7486 16096 -6646
rect 16188 -7486 16190 -6646
rect 16190 -7486 16242 -6646
rect 16242 -7486 16244 -6646
rect 16336 -7486 16338 -6646
rect 16338 -7486 16390 -6646
rect 16390 -7486 16392 -6646
rect 16484 -7486 16486 -6646
rect 16486 -7486 16538 -6646
rect 16538 -7486 16540 -6646
rect 16632 -7486 16634 -6646
rect 16634 -7486 16686 -6646
rect 16686 -7486 16688 -6646
rect 16780 -7486 16782 -6646
rect 16782 -7486 16834 -6646
rect 16834 -7486 16836 -6646
rect 16928 -7486 16930 -6646
rect 16930 -7486 16982 -6646
rect 16982 -7486 16984 -6646
rect 17076 -7486 17078 -6646
rect 17078 -7486 17130 -6646
rect 17130 -7486 17132 -6646
rect 17224 -7486 17226 -6646
rect 17226 -7486 17278 -6646
rect 17278 -7486 17280 -6646
rect 17372 -7486 17374 -6646
rect 17374 -7486 17426 -6646
rect 17426 -7486 17428 -6646
rect 17520 -7486 17522 -6646
rect 17522 -7486 17574 -6646
rect 17574 -7486 17576 -6646
rect 17668 -7486 17670 -6646
rect 17670 -7486 17722 -6646
rect 17722 -7486 17724 -6646
rect 17816 -7486 17818 -6646
rect 17818 -7486 17870 -6646
rect 17870 -7486 17872 -6646
rect 17964 -7486 17966 -6646
rect 17966 -7486 18018 -6646
rect 18018 -7486 18020 -6646
rect 18112 -7486 18114 -6646
rect 18114 -7486 18166 -6646
rect 18166 -7486 18168 -6646
rect 18260 -7486 18262 -6646
rect 18262 -7486 18314 -6646
rect 18314 -7486 18316 -6646
rect 18408 -7486 18410 -6646
rect 18410 -7486 18462 -6646
rect 18462 -7486 18464 -6646
rect 18556 -7486 18558 -6646
rect 18558 -7486 18610 -6646
rect 18610 -7486 18612 -6646
rect 18704 -7486 18706 -6646
rect 18706 -7486 18758 -6646
rect 18758 -7486 18760 -6646
rect 18852 -7486 18854 -6646
rect 18854 -7486 18906 -6646
rect 18906 -7486 18908 -6646
rect 19000 -7486 19002 -6646
rect 19002 -7486 19054 -6646
rect 19054 -7486 19056 -6646
rect 19148 -7486 19150 -6646
rect 19150 -7486 19202 -6646
rect 19202 -7486 19204 -6646
rect 19296 -7486 19298 -6646
rect 19298 -7486 19350 -6646
rect 19350 -7486 19352 -6646
rect 19444 -7486 19446 -6646
rect 19446 -7486 19498 -6646
rect 19498 -7486 19500 -6646
rect 19592 -7486 19594 -6646
rect 19594 -7486 19646 -6646
rect 19646 -7486 19648 -6646
rect 19740 -7486 19742 -6646
rect 19742 -7486 19794 -6646
rect 19794 -7486 19796 -6646
rect 19888 -7486 19890 -6646
rect 19890 -7486 19942 -6646
rect 19942 -7486 19944 -6646
rect 20036 -7486 20038 -6646
rect 20038 -7486 20090 -6646
rect 20090 -7486 20092 -6646
rect 20184 -7486 20186 -6646
rect 20186 -7486 20238 -6646
rect 20238 -7486 20240 -6646
rect 20332 -7486 20334 -6646
rect 20334 -7486 20386 -6646
rect 20386 -7486 20388 -6646
rect 20480 -7486 20482 -6646
rect 20482 -7486 20534 -6646
rect 20534 -7486 20536 -6646
rect 20628 -7486 20630 -6646
rect 20630 -7486 20682 -6646
rect 20682 -7486 20684 -6646
rect 20776 -7486 20778 -6646
rect 20778 -7486 20830 -6646
rect 20830 -7486 20832 -6646
rect 20924 -7486 20926 -6646
rect 20926 -7486 20978 -6646
rect 20978 -7486 20980 -6646
rect 21072 -7486 21074 -6646
rect 21074 -7486 21126 -6646
rect 21126 -7486 21128 -6646
rect 21220 -7486 21222 -6646
rect 21222 -7486 21274 -6646
rect 21274 -7486 21276 -6646
rect 21368 -7486 21370 -6646
rect 21370 -7486 21422 -6646
rect 21422 -7486 21424 -6646
rect 21516 -7486 21518 -6646
rect 21518 -7486 21570 -6646
rect 21570 -7486 21572 -6646
rect 21664 -7486 21666 -6646
rect 21666 -7486 21718 -6646
rect 21718 -7486 21720 -6646
rect 21812 -7486 21814 -6646
rect 21814 -7486 21866 -6646
rect 21866 -7486 21868 -6646
rect 21960 -7486 21962 -6646
rect 21962 -7486 22014 -6646
rect 22014 -7486 22016 -6646
rect 22108 -7486 22110 -6646
rect 22110 -7486 22162 -6646
rect 22162 -7486 22164 -6646
rect 22256 -7486 22258 -6646
rect 22258 -7486 22310 -6646
rect 22310 -7486 22312 -6646
rect 22404 -7486 22406 -6646
rect 22406 -7486 22458 -6646
rect 22458 -7486 22460 -6646
rect 22552 -7486 22554 -6646
rect 22554 -7486 22606 -6646
rect 22606 -7486 22608 -6646
rect 11452 -8632 11454 -7792
rect 11454 -8632 11506 -7792
rect 11506 -8632 11508 -7792
rect 11600 -8632 11602 -7792
rect 11602 -8632 11654 -7792
rect 11654 -8632 11656 -7792
rect 11748 -8632 11750 -7792
rect 11750 -8632 11802 -7792
rect 11802 -8632 11804 -7792
rect 11896 -8632 11898 -7792
rect 11898 -8632 11950 -7792
rect 11950 -8632 11952 -7792
rect 12044 -8632 12046 -7792
rect 12046 -8632 12098 -7792
rect 12098 -8632 12100 -7792
rect 12192 -8632 12194 -7792
rect 12194 -8632 12246 -7792
rect 12246 -8632 12248 -7792
rect 12340 -8632 12342 -7792
rect 12342 -8632 12394 -7792
rect 12394 -8632 12396 -7792
rect 12488 -8632 12490 -7792
rect 12490 -8632 12542 -7792
rect 12542 -8632 12544 -7792
rect 12636 -8632 12638 -7792
rect 12638 -8632 12690 -7792
rect 12690 -8632 12692 -7792
rect 12784 -8632 12786 -7792
rect 12786 -8632 12838 -7792
rect 12838 -8632 12840 -7792
rect 12932 -8632 12934 -7792
rect 12934 -8632 12986 -7792
rect 12986 -8632 12988 -7792
rect 13080 -8632 13082 -7792
rect 13082 -8632 13134 -7792
rect 13134 -8632 13136 -7792
rect 13228 -8632 13230 -7792
rect 13230 -8632 13282 -7792
rect 13282 -8632 13284 -7792
rect 13376 -8632 13378 -7792
rect 13378 -8632 13430 -7792
rect 13430 -8632 13432 -7792
rect 13524 -8632 13526 -7792
rect 13526 -8632 13578 -7792
rect 13578 -8632 13580 -7792
rect 13672 -8632 13674 -7792
rect 13674 -8632 13726 -7792
rect 13726 -8632 13728 -7792
rect 13820 -8632 13822 -7792
rect 13822 -8632 13874 -7792
rect 13874 -8632 13876 -7792
rect 13968 -8632 13970 -7792
rect 13970 -8632 14022 -7792
rect 14022 -8632 14024 -7792
rect 14116 -8632 14118 -7792
rect 14118 -8632 14170 -7792
rect 14170 -8632 14172 -7792
rect 14264 -8632 14266 -7792
rect 14266 -8632 14318 -7792
rect 14318 -8632 14320 -7792
rect 14412 -8632 14414 -7792
rect 14414 -8632 14466 -7792
rect 14466 -8632 14468 -7792
rect 14560 -8632 14562 -7792
rect 14562 -8632 14614 -7792
rect 14614 -8632 14616 -7792
rect 14708 -8632 14710 -7792
rect 14710 -8632 14762 -7792
rect 14762 -8632 14764 -7792
rect 14856 -8632 14858 -7792
rect 14858 -8632 14910 -7792
rect 14910 -8632 14912 -7792
rect 15004 -8632 15006 -7792
rect 15006 -8632 15058 -7792
rect 15058 -8632 15060 -7792
rect 15152 -8632 15154 -7792
rect 15154 -8632 15206 -7792
rect 15206 -8632 15208 -7792
rect 15300 -8632 15302 -7792
rect 15302 -8632 15354 -7792
rect 15354 -8632 15356 -7792
rect 15448 -8632 15450 -7792
rect 15450 -8632 15502 -7792
rect 15502 -8632 15504 -7792
rect 15596 -8632 15598 -7792
rect 15598 -8632 15650 -7792
rect 15650 -8632 15652 -7792
rect 15744 -8632 15746 -7792
rect 15746 -8632 15798 -7792
rect 15798 -8632 15800 -7792
rect 15892 -8632 15894 -7792
rect 15894 -8632 15946 -7792
rect 15946 -8632 15948 -7792
rect 16040 -8632 16042 -7792
rect 16042 -8632 16094 -7792
rect 16094 -8632 16096 -7792
rect 16188 -8632 16190 -7792
rect 16190 -8632 16242 -7792
rect 16242 -8632 16244 -7792
rect 16336 -8632 16338 -7792
rect 16338 -8632 16390 -7792
rect 16390 -8632 16392 -7792
rect 16484 -8632 16486 -7792
rect 16486 -8632 16538 -7792
rect 16538 -8632 16540 -7792
rect 16632 -8632 16634 -7792
rect 16634 -8632 16686 -7792
rect 16686 -8632 16688 -7792
rect 16780 -8632 16782 -7792
rect 16782 -8632 16834 -7792
rect 16834 -8632 16836 -7792
rect 16928 -8632 16930 -7792
rect 16930 -8632 16982 -7792
rect 16982 -8632 16984 -7792
rect 17076 -8632 17078 -7792
rect 17078 -8632 17130 -7792
rect 17130 -8632 17132 -7792
rect 17224 -8632 17226 -7792
rect 17226 -8632 17278 -7792
rect 17278 -8632 17280 -7792
rect 17372 -8632 17374 -7792
rect 17374 -8632 17426 -7792
rect 17426 -8632 17428 -7792
rect 17520 -8632 17522 -7792
rect 17522 -8632 17574 -7792
rect 17574 -8632 17576 -7792
rect 17668 -8632 17670 -7792
rect 17670 -8632 17722 -7792
rect 17722 -8632 17724 -7792
rect 17816 -8632 17818 -7792
rect 17818 -8632 17870 -7792
rect 17870 -8632 17872 -7792
rect 17964 -8632 17966 -7792
rect 17966 -8632 18018 -7792
rect 18018 -8632 18020 -7792
rect 18112 -8632 18114 -7792
rect 18114 -8632 18166 -7792
rect 18166 -8632 18168 -7792
rect 18260 -8632 18262 -7792
rect 18262 -8632 18314 -7792
rect 18314 -8632 18316 -7792
rect 18408 -8632 18410 -7792
rect 18410 -8632 18462 -7792
rect 18462 -8632 18464 -7792
rect 18556 -8632 18558 -7792
rect 18558 -8632 18610 -7792
rect 18610 -8632 18612 -7792
rect 18704 -8632 18706 -7792
rect 18706 -8632 18758 -7792
rect 18758 -8632 18760 -7792
rect 18852 -8632 18854 -7792
rect 18854 -8632 18906 -7792
rect 18906 -8632 18908 -7792
rect 19000 -8632 19002 -7792
rect 19002 -8632 19054 -7792
rect 19054 -8632 19056 -7792
rect 19148 -8632 19150 -7792
rect 19150 -8632 19202 -7792
rect 19202 -8632 19204 -7792
rect 19296 -8632 19298 -7792
rect 19298 -8632 19350 -7792
rect 19350 -8632 19352 -7792
rect 19444 -8632 19446 -7792
rect 19446 -8632 19498 -7792
rect 19498 -8632 19500 -7792
rect 19592 -8632 19594 -7792
rect 19594 -8632 19646 -7792
rect 19646 -8632 19648 -7792
rect 19740 -8632 19742 -7792
rect 19742 -8632 19794 -7792
rect 19794 -8632 19796 -7792
rect 19888 -8632 19890 -7792
rect 19890 -8632 19942 -7792
rect 19942 -8632 19944 -7792
rect 20036 -8632 20038 -7792
rect 20038 -8632 20090 -7792
rect 20090 -8632 20092 -7792
rect 20184 -8632 20186 -7792
rect 20186 -8632 20238 -7792
rect 20238 -8632 20240 -7792
rect 20332 -8632 20334 -7792
rect 20334 -8632 20386 -7792
rect 20386 -8632 20388 -7792
rect 20480 -8632 20482 -7792
rect 20482 -8632 20534 -7792
rect 20534 -8632 20536 -7792
rect 20628 -8632 20630 -7792
rect 20630 -8632 20682 -7792
rect 20682 -8632 20684 -7792
rect 20776 -8632 20778 -7792
rect 20778 -8632 20830 -7792
rect 20830 -8632 20832 -7792
rect 20924 -8632 20926 -7792
rect 20926 -8632 20978 -7792
rect 20978 -8632 20980 -7792
rect 21072 -8632 21074 -7792
rect 21074 -8632 21126 -7792
rect 21126 -8632 21128 -7792
rect 21220 -8632 21222 -7792
rect 21222 -8632 21274 -7792
rect 21274 -8632 21276 -7792
rect 21368 -8632 21370 -7792
rect 21370 -8632 21422 -7792
rect 21422 -8632 21424 -7792
rect 21516 -8632 21518 -7792
rect 21518 -8632 21570 -7792
rect 21570 -8632 21572 -7792
rect 21664 -8632 21666 -7792
rect 21666 -8632 21718 -7792
rect 21718 -8632 21720 -7792
rect 21812 -8632 21814 -7792
rect 21814 -8632 21866 -7792
rect 21866 -8632 21868 -7792
rect 21960 -8632 21962 -7792
rect 21962 -8632 22014 -7792
rect 22014 -8632 22016 -7792
rect 22108 -8632 22110 -7792
rect 22110 -8632 22162 -7792
rect 22162 -8632 22164 -7792
rect 22256 -8632 22258 -7792
rect 22258 -8632 22310 -7792
rect 22310 -8632 22312 -7792
rect 22404 -8632 22406 -7792
rect 22406 -8632 22458 -7792
rect 22458 -8632 22460 -7792
rect 22552 -8632 22554 -7792
rect 22554 -8632 22606 -7792
rect 22606 -8632 22608 -7792
rect 23053 -7926 23055 -7086
rect 23055 -7926 23107 -7086
rect 23107 -7926 23109 -7086
rect 23231 -7939 23233 -7099
rect 23233 -7939 23285 -7099
rect 23285 -7939 23287 -7099
<< metal3 >>
rect 11442 -6646 11518 -6641
rect 11442 -7486 11452 -6646
rect 11508 -7486 11518 -6646
rect 11442 -7792 11518 -7486
rect 11586 -7481 11596 -6641
rect 11660 -7481 11670 -6641
rect 11586 -7486 11600 -7481
rect 11656 -7486 11670 -7481
rect 11586 -7491 11670 -7486
rect 11738 -6646 11814 -6641
rect 11738 -7486 11748 -6646
rect 11804 -7486 11814 -6646
rect 11442 -8632 11452 -7792
rect 11508 -8632 11518 -7792
rect 11442 -8637 11518 -8632
rect 11586 -7792 11670 -7787
rect 11586 -7797 11600 -7792
rect 11656 -7797 11670 -7792
rect 11586 -8637 11596 -7797
rect 11660 -8637 11670 -7797
rect 11738 -7792 11814 -7486
rect 11882 -7481 11892 -6641
rect 11956 -7481 11966 -6641
rect 11882 -7486 11896 -7481
rect 11952 -7486 11966 -7481
rect 11882 -7491 11966 -7486
rect 12034 -6646 12110 -6641
rect 12034 -7486 12044 -6646
rect 12100 -7486 12110 -6646
rect 11738 -8632 11748 -7792
rect 11804 -8632 11814 -7792
rect 11738 -8637 11814 -8632
rect 11882 -7792 11966 -7787
rect 11882 -7797 11896 -7792
rect 11952 -7797 11966 -7792
rect 11882 -8637 11892 -7797
rect 11956 -8637 11966 -7797
rect 12034 -7792 12110 -7486
rect 12178 -7481 12188 -6641
rect 12252 -7481 12262 -6641
rect 12178 -7486 12192 -7481
rect 12248 -7486 12262 -7481
rect 12178 -7491 12262 -7486
rect 12330 -6646 12406 -6641
rect 12330 -7486 12340 -6646
rect 12396 -7486 12406 -6646
rect 12034 -8632 12044 -7792
rect 12100 -8632 12110 -7792
rect 12034 -8637 12110 -8632
rect 12178 -7792 12262 -7787
rect 12178 -7797 12192 -7792
rect 12248 -7797 12262 -7792
rect 12178 -8637 12188 -7797
rect 12252 -8637 12262 -7797
rect 12330 -7792 12406 -7486
rect 12474 -7481 12484 -6641
rect 12548 -7481 12558 -6641
rect 12474 -7486 12488 -7481
rect 12544 -7486 12558 -7481
rect 12474 -7491 12558 -7486
rect 12626 -6646 12702 -6641
rect 12626 -7486 12636 -6646
rect 12692 -7486 12702 -6646
rect 12330 -8632 12340 -7792
rect 12396 -8632 12406 -7792
rect 12330 -8637 12406 -8632
rect 12474 -7792 12558 -7787
rect 12474 -7797 12488 -7792
rect 12544 -7797 12558 -7792
rect 12474 -8637 12484 -7797
rect 12548 -8637 12558 -7797
rect 12626 -7792 12702 -7486
rect 12770 -7481 12780 -6641
rect 12844 -7481 12854 -6641
rect 12770 -7486 12784 -7481
rect 12840 -7486 12854 -7481
rect 12770 -7491 12854 -7486
rect 12922 -6646 12998 -6641
rect 12922 -7486 12932 -6646
rect 12988 -7486 12998 -6646
rect 12626 -8632 12636 -7792
rect 12692 -8632 12702 -7792
rect 12626 -8637 12702 -8632
rect 12770 -7792 12854 -7787
rect 12770 -7797 12784 -7792
rect 12840 -7797 12854 -7792
rect 12770 -8637 12780 -7797
rect 12844 -8637 12854 -7797
rect 12922 -7792 12998 -7486
rect 13066 -7481 13076 -6641
rect 13140 -7481 13150 -6641
rect 13066 -7486 13080 -7481
rect 13136 -7486 13150 -7481
rect 13066 -7491 13150 -7486
rect 13218 -6646 13294 -6641
rect 13218 -7486 13228 -6646
rect 13284 -7486 13294 -6646
rect 12922 -8632 12932 -7792
rect 12988 -8632 12998 -7792
rect 12922 -8637 12998 -8632
rect 13066 -7792 13150 -7787
rect 13066 -7797 13080 -7792
rect 13136 -7797 13150 -7792
rect 13066 -8637 13076 -7797
rect 13140 -8637 13150 -7797
rect 13218 -7792 13294 -7486
rect 13362 -7481 13372 -6641
rect 13436 -7481 13446 -6641
rect 13362 -7486 13376 -7481
rect 13432 -7486 13446 -7481
rect 13362 -7491 13446 -7486
rect 13514 -6646 13590 -6641
rect 13514 -7486 13524 -6646
rect 13580 -7486 13590 -6646
rect 13218 -8632 13228 -7792
rect 13284 -8632 13294 -7792
rect 13218 -8637 13294 -8632
rect 13362 -7792 13446 -7787
rect 13362 -7797 13376 -7792
rect 13432 -7797 13446 -7792
rect 13362 -8637 13372 -7797
rect 13436 -8637 13446 -7797
rect 13514 -7792 13590 -7486
rect 13658 -7481 13668 -6641
rect 13732 -7481 13742 -6641
rect 13658 -7486 13672 -7481
rect 13728 -7486 13742 -7481
rect 13658 -7491 13742 -7486
rect 13810 -6646 13886 -6641
rect 13810 -7486 13820 -6646
rect 13876 -7486 13886 -6646
rect 13514 -8632 13524 -7792
rect 13580 -8632 13590 -7792
rect 13514 -8637 13590 -8632
rect 13658 -7792 13742 -7787
rect 13658 -7797 13672 -7792
rect 13728 -7797 13742 -7792
rect 13658 -8637 13668 -7797
rect 13732 -8637 13742 -7797
rect 13810 -7792 13886 -7486
rect 13954 -7481 13964 -6641
rect 14028 -7481 14038 -6641
rect 13954 -7486 13968 -7481
rect 14024 -7486 14038 -7481
rect 13954 -7491 14038 -7486
rect 14106 -6646 14182 -6641
rect 14106 -7486 14116 -6646
rect 14172 -7486 14182 -6646
rect 13810 -8632 13820 -7792
rect 13876 -8632 13886 -7792
rect 13810 -8637 13886 -8632
rect 13954 -7792 14038 -7787
rect 13954 -7797 13968 -7792
rect 14024 -7797 14038 -7792
rect 13954 -8637 13964 -7797
rect 14028 -8637 14038 -7797
rect 14106 -7792 14182 -7486
rect 14250 -7481 14260 -6641
rect 14324 -7481 14334 -6641
rect 14250 -7486 14264 -7481
rect 14320 -7486 14334 -7481
rect 14250 -7491 14334 -7486
rect 14402 -6646 14478 -6641
rect 14402 -7486 14412 -6646
rect 14468 -7486 14478 -6646
rect 14106 -8632 14116 -7792
rect 14172 -8632 14182 -7792
rect 14106 -8637 14182 -8632
rect 14250 -7792 14334 -7787
rect 14250 -7797 14264 -7792
rect 14320 -7797 14334 -7792
rect 14250 -8637 14260 -7797
rect 14324 -8637 14334 -7797
rect 14402 -7792 14478 -7486
rect 14546 -7481 14556 -6641
rect 14620 -7481 14630 -6641
rect 14546 -7486 14560 -7481
rect 14616 -7486 14630 -7481
rect 14546 -7491 14630 -7486
rect 14698 -6646 14774 -6641
rect 14698 -7486 14708 -6646
rect 14764 -7486 14774 -6646
rect 14402 -8632 14412 -7792
rect 14468 -8632 14478 -7792
rect 14402 -8637 14478 -8632
rect 14546 -7792 14630 -7787
rect 14546 -7797 14560 -7792
rect 14616 -7797 14630 -7792
rect 14546 -8637 14556 -7797
rect 14620 -8637 14630 -7797
rect 14698 -7792 14774 -7486
rect 14842 -7481 14852 -6641
rect 14916 -7481 14926 -6641
rect 14842 -7486 14856 -7481
rect 14912 -7486 14926 -7481
rect 14842 -7491 14926 -7486
rect 14994 -6646 15070 -6641
rect 14994 -7486 15004 -6646
rect 15060 -7486 15070 -6646
rect 14698 -8632 14708 -7792
rect 14764 -8632 14774 -7792
rect 14698 -8637 14774 -8632
rect 14842 -7792 14926 -7787
rect 14842 -7797 14856 -7792
rect 14912 -7797 14926 -7792
rect 14842 -8637 14852 -7797
rect 14916 -8637 14926 -7797
rect 14994 -7792 15070 -7486
rect 15138 -7481 15148 -6641
rect 15212 -7481 15222 -6641
rect 15138 -7486 15152 -7481
rect 15208 -7486 15222 -7481
rect 15138 -7491 15222 -7486
rect 15290 -6646 15366 -6641
rect 15290 -7486 15300 -6646
rect 15356 -7486 15366 -6646
rect 14994 -8632 15004 -7792
rect 15060 -8632 15070 -7792
rect 14994 -8637 15070 -8632
rect 15138 -7792 15222 -7787
rect 15138 -7797 15152 -7792
rect 15208 -7797 15222 -7792
rect 15138 -8637 15148 -7797
rect 15212 -8637 15222 -7797
rect 15290 -7792 15366 -7486
rect 15434 -7481 15444 -6641
rect 15508 -7481 15518 -6641
rect 15434 -7486 15448 -7481
rect 15504 -7486 15518 -7481
rect 15434 -7491 15518 -7486
rect 15586 -6646 15662 -6641
rect 15586 -7486 15596 -6646
rect 15652 -7486 15662 -6646
rect 15290 -8632 15300 -7792
rect 15356 -8632 15366 -7792
rect 15290 -8637 15366 -8632
rect 15434 -7792 15518 -7787
rect 15434 -7797 15448 -7792
rect 15504 -7797 15518 -7792
rect 15434 -8637 15444 -7797
rect 15508 -8637 15518 -7797
rect 15586 -7792 15662 -7486
rect 15730 -7481 15740 -6641
rect 15804 -7481 15814 -6641
rect 15730 -7486 15744 -7481
rect 15800 -7486 15814 -7481
rect 15730 -7491 15814 -7486
rect 15882 -6646 15958 -6641
rect 15882 -7486 15892 -6646
rect 15948 -7486 15958 -6646
rect 15586 -8632 15596 -7792
rect 15652 -8632 15662 -7792
rect 15586 -8637 15662 -8632
rect 15730 -7792 15814 -7787
rect 15730 -7797 15744 -7792
rect 15800 -7797 15814 -7792
rect 15730 -8637 15740 -7797
rect 15804 -8637 15814 -7797
rect 15882 -7792 15958 -7486
rect 16026 -7481 16036 -6641
rect 16100 -7481 16110 -6641
rect 16026 -7486 16040 -7481
rect 16096 -7486 16110 -7481
rect 16026 -7491 16110 -7486
rect 16178 -6646 16254 -6641
rect 16178 -7486 16188 -6646
rect 16244 -7486 16254 -6646
rect 15882 -8632 15892 -7792
rect 15948 -8632 15958 -7792
rect 15882 -8637 15958 -8632
rect 16026 -7792 16110 -7787
rect 16026 -7797 16040 -7792
rect 16096 -7797 16110 -7792
rect 16026 -8637 16036 -7797
rect 16100 -8637 16110 -7797
rect 16178 -7792 16254 -7486
rect 16322 -7481 16332 -6641
rect 16396 -7481 16406 -6641
rect 16322 -7486 16336 -7481
rect 16392 -7486 16406 -7481
rect 16322 -7491 16406 -7486
rect 16474 -6646 16550 -6641
rect 16474 -7486 16484 -6646
rect 16540 -7486 16550 -6646
rect 16178 -8632 16188 -7792
rect 16244 -8632 16254 -7792
rect 16178 -8637 16254 -8632
rect 16322 -7792 16406 -7787
rect 16322 -7797 16336 -7792
rect 16392 -7797 16406 -7792
rect 16322 -8637 16332 -7797
rect 16396 -8637 16406 -7797
rect 16474 -7792 16550 -7486
rect 16618 -7481 16628 -6641
rect 16692 -7481 16702 -6641
rect 16618 -7486 16632 -7481
rect 16688 -7486 16702 -7481
rect 16618 -7491 16702 -7486
rect 16770 -6646 16846 -6641
rect 16770 -7486 16780 -6646
rect 16836 -7486 16846 -6646
rect 16474 -8632 16484 -7792
rect 16540 -8632 16550 -7792
rect 16474 -8637 16550 -8632
rect 16618 -7792 16702 -7787
rect 16618 -7797 16632 -7792
rect 16688 -7797 16702 -7792
rect 16618 -8637 16628 -7797
rect 16692 -8637 16702 -7797
rect 16770 -7792 16846 -7486
rect 16914 -7481 16924 -6641
rect 16988 -7481 16998 -6641
rect 16914 -7486 16928 -7481
rect 16984 -7486 16998 -7481
rect 16914 -7491 16998 -7486
rect 17066 -6646 17142 -6641
rect 17066 -7486 17076 -6646
rect 17132 -7486 17142 -6646
rect 16770 -8632 16780 -7792
rect 16836 -8632 16846 -7792
rect 16770 -8637 16846 -8632
rect 16914 -7792 16998 -7787
rect 16914 -7797 16928 -7792
rect 16984 -7797 16998 -7792
rect 16914 -8637 16924 -7797
rect 16988 -8637 16998 -7797
rect 17066 -7792 17142 -7486
rect 17210 -7481 17220 -6641
rect 17284 -7481 17294 -6641
rect 17210 -7486 17224 -7481
rect 17280 -7486 17294 -7481
rect 17210 -7491 17294 -7486
rect 17362 -6646 17438 -6641
rect 17362 -7486 17372 -6646
rect 17428 -7486 17438 -6646
rect 17066 -8632 17076 -7792
rect 17132 -8632 17142 -7792
rect 17066 -8637 17142 -8632
rect 17210 -7792 17294 -7787
rect 17210 -7797 17224 -7792
rect 17280 -7797 17294 -7792
rect 17210 -8637 17220 -7797
rect 17284 -8637 17294 -7797
rect 17362 -7792 17438 -7486
rect 17506 -7481 17516 -6641
rect 17580 -7481 17590 -6641
rect 17506 -7486 17520 -7481
rect 17576 -7486 17590 -7481
rect 17506 -7491 17590 -7486
rect 17658 -6646 17734 -6641
rect 17658 -7486 17668 -6646
rect 17724 -7486 17734 -6646
rect 17362 -8632 17372 -7792
rect 17428 -8632 17438 -7792
rect 17362 -8637 17438 -8632
rect 17506 -7792 17590 -7787
rect 17506 -7797 17520 -7792
rect 17576 -7797 17590 -7792
rect 17506 -8637 17516 -7797
rect 17580 -8637 17590 -7797
rect 17658 -7792 17734 -7486
rect 17802 -7481 17812 -6641
rect 17876 -7481 17886 -6641
rect 17802 -7486 17816 -7481
rect 17872 -7486 17886 -7481
rect 17802 -7491 17886 -7486
rect 17954 -6646 18030 -6641
rect 17954 -7486 17964 -6646
rect 18020 -7486 18030 -6646
rect 17658 -8632 17668 -7792
rect 17724 -8632 17734 -7792
rect 17658 -8637 17734 -8632
rect 17802 -7792 17886 -7787
rect 17802 -7797 17816 -7792
rect 17872 -7797 17886 -7792
rect 17802 -8637 17812 -7797
rect 17876 -8637 17886 -7797
rect 17954 -7792 18030 -7486
rect 18098 -7481 18108 -6641
rect 18172 -7481 18182 -6641
rect 18098 -7486 18112 -7481
rect 18168 -7486 18182 -7481
rect 18098 -7491 18182 -7486
rect 18250 -6646 18326 -6641
rect 18250 -7486 18260 -6646
rect 18316 -7486 18326 -6646
rect 17954 -8632 17964 -7792
rect 18020 -8632 18030 -7792
rect 17954 -8637 18030 -8632
rect 18098 -7792 18182 -7787
rect 18098 -7797 18112 -7792
rect 18168 -7797 18182 -7792
rect 18098 -8637 18108 -7797
rect 18172 -8637 18182 -7797
rect 18250 -7792 18326 -7486
rect 18394 -7481 18404 -6641
rect 18468 -7481 18478 -6641
rect 18394 -7486 18408 -7481
rect 18464 -7486 18478 -7481
rect 18394 -7491 18478 -7486
rect 18546 -6646 18622 -6641
rect 18546 -7486 18556 -6646
rect 18612 -7486 18622 -6646
rect 18250 -8632 18260 -7792
rect 18316 -8632 18326 -7792
rect 18250 -8637 18326 -8632
rect 18394 -7792 18478 -7787
rect 18394 -7797 18408 -7792
rect 18464 -7797 18478 -7792
rect 18394 -8637 18404 -7797
rect 18468 -8637 18478 -7797
rect 18546 -7792 18622 -7486
rect 18690 -7481 18700 -6641
rect 18764 -7481 18774 -6641
rect 18690 -7486 18704 -7481
rect 18760 -7486 18774 -7481
rect 18690 -7491 18774 -7486
rect 18842 -6646 18918 -6641
rect 18842 -7486 18852 -6646
rect 18908 -7486 18918 -6646
rect 18546 -8632 18556 -7792
rect 18612 -8632 18622 -7792
rect 18546 -8637 18622 -8632
rect 18690 -7792 18774 -7787
rect 18690 -7797 18704 -7792
rect 18760 -7797 18774 -7792
rect 18690 -8637 18700 -7797
rect 18764 -8637 18774 -7797
rect 18842 -7792 18918 -7486
rect 18986 -7481 18996 -6641
rect 19060 -7481 19070 -6641
rect 18986 -7486 19000 -7481
rect 19056 -7486 19070 -7481
rect 18986 -7491 19070 -7486
rect 19138 -6646 19214 -6641
rect 19138 -7486 19148 -6646
rect 19204 -7486 19214 -6646
rect 18842 -8632 18852 -7792
rect 18908 -8632 18918 -7792
rect 18842 -8637 18918 -8632
rect 18986 -7792 19070 -7787
rect 18986 -7797 19000 -7792
rect 19056 -7797 19070 -7792
rect 18986 -8637 18996 -7797
rect 19060 -8637 19070 -7797
rect 19138 -7792 19214 -7486
rect 19282 -7481 19292 -6641
rect 19356 -7481 19366 -6641
rect 19282 -7486 19296 -7481
rect 19352 -7486 19366 -7481
rect 19282 -7491 19366 -7486
rect 19434 -6646 19510 -6641
rect 19434 -7486 19444 -6646
rect 19500 -7486 19510 -6646
rect 19138 -8632 19148 -7792
rect 19204 -8632 19214 -7792
rect 19138 -8637 19214 -8632
rect 19282 -7792 19366 -7787
rect 19282 -7797 19296 -7792
rect 19352 -7797 19366 -7792
rect 19282 -8637 19292 -7797
rect 19356 -8637 19366 -7797
rect 19434 -7792 19510 -7486
rect 19578 -7481 19588 -6641
rect 19652 -7481 19662 -6641
rect 19578 -7486 19592 -7481
rect 19648 -7486 19662 -7481
rect 19578 -7491 19662 -7486
rect 19730 -6646 19806 -6641
rect 19730 -7486 19740 -6646
rect 19796 -7486 19806 -6646
rect 19434 -8632 19444 -7792
rect 19500 -8632 19510 -7792
rect 19434 -8637 19510 -8632
rect 19578 -7792 19662 -7787
rect 19578 -7797 19592 -7792
rect 19648 -7797 19662 -7792
rect 19578 -8637 19588 -7797
rect 19652 -8637 19662 -7797
rect 19730 -7792 19806 -7486
rect 19874 -7481 19884 -6641
rect 19948 -7481 19958 -6641
rect 19874 -7486 19888 -7481
rect 19944 -7486 19958 -7481
rect 19874 -7491 19958 -7486
rect 20026 -6646 20102 -6641
rect 20026 -7486 20036 -6646
rect 20092 -7486 20102 -6646
rect 19730 -8632 19740 -7792
rect 19796 -8632 19806 -7792
rect 19730 -8637 19806 -8632
rect 19874 -7792 19958 -7787
rect 19874 -7797 19888 -7792
rect 19944 -7797 19958 -7792
rect 19874 -8637 19884 -7797
rect 19948 -8637 19958 -7797
rect 20026 -7792 20102 -7486
rect 20170 -7481 20180 -6641
rect 20244 -7481 20254 -6641
rect 20170 -7486 20184 -7481
rect 20240 -7486 20254 -7481
rect 20170 -7491 20254 -7486
rect 20322 -6646 20398 -6641
rect 20322 -7486 20332 -6646
rect 20388 -7486 20398 -6646
rect 20026 -8632 20036 -7792
rect 20092 -8632 20102 -7792
rect 20026 -8637 20102 -8632
rect 20170 -7792 20254 -7787
rect 20170 -7797 20184 -7792
rect 20240 -7797 20254 -7792
rect 20170 -8637 20180 -7797
rect 20244 -8637 20254 -7797
rect 20322 -7792 20398 -7486
rect 20466 -7481 20476 -6641
rect 20540 -7481 20550 -6641
rect 20466 -7486 20480 -7481
rect 20536 -7486 20550 -7481
rect 20466 -7491 20550 -7486
rect 20618 -6646 20694 -6641
rect 20618 -7486 20628 -6646
rect 20684 -7486 20694 -6646
rect 20322 -8632 20332 -7792
rect 20388 -8632 20398 -7792
rect 20322 -8637 20398 -8632
rect 20466 -7792 20550 -7787
rect 20466 -7797 20480 -7792
rect 20536 -7797 20550 -7792
rect 20466 -8637 20476 -7797
rect 20540 -8637 20550 -7797
rect 20618 -7792 20694 -7486
rect 20762 -7481 20772 -6641
rect 20836 -7481 20846 -6641
rect 20762 -7486 20776 -7481
rect 20832 -7486 20846 -7481
rect 20762 -7491 20846 -7486
rect 20914 -6646 20990 -6641
rect 20914 -7486 20924 -6646
rect 20980 -7486 20990 -6646
rect 20618 -8632 20628 -7792
rect 20684 -8632 20694 -7792
rect 20618 -8637 20694 -8632
rect 20762 -7792 20846 -7787
rect 20762 -7797 20776 -7792
rect 20832 -7797 20846 -7792
rect 20762 -8637 20772 -7797
rect 20836 -8637 20846 -7797
rect 20914 -7792 20990 -7486
rect 21058 -7481 21068 -6641
rect 21132 -7481 21142 -6641
rect 21058 -7486 21072 -7481
rect 21128 -7486 21142 -7481
rect 21058 -7491 21142 -7486
rect 21210 -6646 21286 -6641
rect 21210 -7486 21220 -6646
rect 21276 -7486 21286 -6646
rect 20914 -8632 20924 -7792
rect 20980 -8632 20990 -7792
rect 20914 -8637 20990 -8632
rect 21058 -7792 21142 -7787
rect 21058 -7797 21072 -7792
rect 21128 -7797 21142 -7792
rect 21058 -8637 21068 -7797
rect 21132 -8637 21142 -7797
rect 21210 -7792 21286 -7486
rect 21354 -7481 21364 -6641
rect 21428 -7481 21438 -6641
rect 21354 -7486 21368 -7481
rect 21424 -7486 21438 -7481
rect 21354 -7491 21438 -7486
rect 21506 -6646 21582 -6641
rect 21506 -7486 21516 -6646
rect 21572 -7486 21582 -6646
rect 21210 -8632 21220 -7792
rect 21276 -8632 21286 -7792
rect 21210 -8637 21286 -8632
rect 21354 -7792 21438 -7787
rect 21354 -7797 21368 -7792
rect 21424 -7797 21438 -7792
rect 21354 -8637 21364 -7797
rect 21428 -8637 21438 -7797
rect 21506 -7792 21582 -7486
rect 21650 -7481 21660 -6641
rect 21724 -7481 21734 -6641
rect 21650 -7486 21664 -7481
rect 21720 -7486 21734 -7481
rect 21650 -7491 21734 -7486
rect 21802 -6646 21878 -6641
rect 21802 -7486 21812 -6646
rect 21868 -7486 21878 -6646
rect 21506 -8632 21516 -7792
rect 21572 -8632 21582 -7792
rect 21506 -8637 21582 -8632
rect 21650 -7792 21734 -7787
rect 21650 -7797 21664 -7792
rect 21720 -7797 21734 -7792
rect 21650 -8637 21660 -7797
rect 21724 -8637 21734 -7797
rect 21802 -7792 21878 -7486
rect 21946 -7481 21956 -6641
rect 22020 -7481 22030 -6641
rect 21946 -7486 21960 -7481
rect 22016 -7486 22030 -7481
rect 21946 -7491 22030 -7486
rect 22098 -6646 22174 -6641
rect 22098 -7486 22108 -6646
rect 22164 -7486 22174 -6646
rect 21802 -8632 21812 -7792
rect 21868 -8632 21878 -7792
rect 21802 -8637 21878 -8632
rect 21946 -7792 22030 -7787
rect 21946 -7797 21960 -7792
rect 22016 -7797 22030 -7792
rect 21946 -8637 21956 -7797
rect 22020 -8637 22030 -7797
rect 22098 -7792 22174 -7486
rect 22242 -7481 22252 -6641
rect 22316 -7481 22326 -6641
rect 22242 -7486 22256 -7481
rect 22312 -7486 22326 -7481
rect 22242 -7491 22326 -7486
rect 22394 -6646 22470 -6641
rect 22394 -7486 22404 -6646
rect 22460 -7486 22470 -6646
rect 22098 -8632 22108 -7792
rect 22164 -8632 22174 -7792
rect 22098 -8637 22174 -8632
rect 22242 -7792 22326 -7787
rect 22242 -7797 22256 -7792
rect 22312 -7797 22326 -7792
rect 22242 -8637 22252 -7797
rect 22316 -8637 22326 -7797
rect 22394 -7792 22470 -7486
rect 22538 -7481 22548 -6641
rect 22612 -7481 22622 -6641
rect 22538 -7486 22552 -7481
rect 22608 -7486 22622 -7481
rect 22538 -7491 22622 -7486
rect 23043 -7086 23119 -7081
rect 22394 -8632 22404 -7792
rect 22460 -8632 22470 -7792
rect 22394 -8637 22470 -8632
rect 22538 -7792 22622 -7787
rect 22538 -7797 22552 -7792
rect 22608 -7797 22622 -7792
rect 22538 -8637 22548 -7797
rect 22612 -8637 22622 -7797
rect 23043 -7926 23053 -7086
rect 23109 -7926 23119 -7086
rect 23043 -7931 23119 -7926
rect 23217 -7099 23301 -7094
rect 23217 -7104 23231 -7099
rect 23287 -7104 23301 -7099
rect 23217 -7944 23227 -7104
rect 23291 -7944 23301 -7104
<< via3 >>
rect 11596 -6646 11660 -6641
rect 11596 -7481 11600 -6646
rect 11600 -7481 11656 -6646
rect 11656 -7481 11660 -6646
rect 11596 -8632 11600 -7797
rect 11600 -8632 11656 -7797
rect 11656 -8632 11660 -7797
rect 11596 -8637 11660 -8632
rect 11892 -6646 11956 -6641
rect 11892 -7481 11896 -6646
rect 11896 -7481 11952 -6646
rect 11952 -7481 11956 -6646
rect 11892 -8632 11896 -7797
rect 11896 -8632 11952 -7797
rect 11952 -8632 11956 -7797
rect 11892 -8637 11956 -8632
rect 12188 -6646 12252 -6641
rect 12188 -7481 12192 -6646
rect 12192 -7481 12248 -6646
rect 12248 -7481 12252 -6646
rect 12188 -8632 12192 -7797
rect 12192 -8632 12248 -7797
rect 12248 -8632 12252 -7797
rect 12188 -8637 12252 -8632
rect 12484 -6646 12548 -6641
rect 12484 -7481 12488 -6646
rect 12488 -7481 12544 -6646
rect 12544 -7481 12548 -6646
rect 12484 -8632 12488 -7797
rect 12488 -8632 12544 -7797
rect 12544 -8632 12548 -7797
rect 12484 -8637 12548 -8632
rect 12780 -6646 12844 -6641
rect 12780 -7481 12784 -6646
rect 12784 -7481 12840 -6646
rect 12840 -7481 12844 -6646
rect 12780 -8632 12784 -7797
rect 12784 -8632 12840 -7797
rect 12840 -8632 12844 -7797
rect 12780 -8637 12844 -8632
rect 13076 -6646 13140 -6641
rect 13076 -7481 13080 -6646
rect 13080 -7481 13136 -6646
rect 13136 -7481 13140 -6646
rect 13076 -8632 13080 -7797
rect 13080 -8632 13136 -7797
rect 13136 -8632 13140 -7797
rect 13076 -8637 13140 -8632
rect 13372 -6646 13436 -6641
rect 13372 -7481 13376 -6646
rect 13376 -7481 13432 -6646
rect 13432 -7481 13436 -6646
rect 13372 -8632 13376 -7797
rect 13376 -8632 13432 -7797
rect 13432 -8632 13436 -7797
rect 13372 -8637 13436 -8632
rect 13668 -6646 13732 -6641
rect 13668 -7481 13672 -6646
rect 13672 -7481 13728 -6646
rect 13728 -7481 13732 -6646
rect 13668 -8632 13672 -7797
rect 13672 -8632 13728 -7797
rect 13728 -8632 13732 -7797
rect 13668 -8637 13732 -8632
rect 13964 -6646 14028 -6641
rect 13964 -7481 13968 -6646
rect 13968 -7481 14024 -6646
rect 14024 -7481 14028 -6646
rect 13964 -8632 13968 -7797
rect 13968 -8632 14024 -7797
rect 14024 -8632 14028 -7797
rect 13964 -8637 14028 -8632
rect 14260 -6646 14324 -6641
rect 14260 -7481 14264 -6646
rect 14264 -7481 14320 -6646
rect 14320 -7481 14324 -6646
rect 14260 -8632 14264 -7797
rect 14264 -8632 14320 -7797
rect 14320 -8632 14324 -7797
rect 14260 -8637 14324 -8632
rect 14556 -6646 14620 -6641
rect 14556 -7481 14560 -6646
rect 14560 -7481 14616 -6646
rect 14616 -7481 14620 -6646
rect 14556 -8632 14560 -7797
rect 14560 -8632 14616 -7797
rect 14616 -8632 14620 -7797
rect 14556 -8637 14620 -8632
rect 14852 -6646 14916 -6641
rect 14852 -7481 14856 -6646
rect 14856 -7481 14912 -6646
rect 14912 -7481 14916 -6646
rect 14852 -8632 14856 -7797
rect 14856 -8632 14912 -7797
rect 14912 -8632 14916 -7797
rect 14852 -8637 14916 -8632
rect 15148 -6646 15212 -6641
rect 15148 -7481 15152 -6646
rect 15152 -7481 15208 -6646
rect 15208 -7481 15212 -6646
rect 15148 -8632 15152 -7797
rect 15152 -8632 15208 -7797
rect 15208 -8632 15212 -7797
rect 15148 -8637 15212 -8632
rect 15444 -6646 15508 -6641
rect 15444 -7481 15448 -6646
rect 15448 -7481 15504 -6646
rect 15504 -7481 15508 -6646
rect 15444 -8632 15448 -7797
rect 15448 -8632 15504 -7797
rect 15504 -8632 15508 -7797
rect 15444 -8637 15508 -8632
rect 15740 -6646 15804 -6641
rect 15740 -7481 15744 -6646
rect 15744 -7481 15800 -6646
rect 15800 -7481 15804 -6646
rect 15740 -8632 15744 -7797
rect 15744 -8632 15800 -7797
rect 15800 -8632 15804 -7797
rect 15740 -8637 15804 -8632
rect 16036 -6646 16100 -6641
rect 16036 -7481 16040 -6646
rect 16040 -7481 16096 -6646
rect 16096 -7481 16100 -6646
rect 16036 -8632 16040 -7797
rect 16040 -8632 16096 -7797
rect 16096 -8632 16100 -7797
rect 16036 -8637 16100 -8632
rect 16332 -6646 16396 -6641
rect 16332 -7481 16336 -6646
rect 16336 -7481 16392 -6646
rect 16392 -7481 16396 -6646
rect 16332 -8632 16336 -7797
rect 16336 -8632 16392 -7797
rect 16392 -8632 16396 -7797
rect 16332 -8637 16396 -8632
rect 16628 -6646 16692 -6641
rect 16628 -7481 16632 -6646
rect 16632 -7481 16688 -6646
rect 16688 -7481 16692 -6646
rect 16628 -8632 16632 -7797
rect 16632 -8632 16688 -7797
rect 16688 -8632 16692 -7797
rect 16628 -8637 16692 -8632
rect 16924 -6646 16988 -6641
rect 16924 -7481 16928 -6646
rect 16928 -7481 16984 -6646
rect 16984 -7481 16988 -6646
rect 16924 -8632 16928 -7797
rect 16928 -8632 16984 -7797
rect 16984 -8632 16988 -7797
rect 16924 -8637 16988 -8632
rect 17220 -6646 17284 -6641
rect 17220 -7481 17224 -6646
rect 17224 -7481 17280 -6646
rect 17280 -7481 17284 -6646
rect 17220 -8632 17224 -7797
rect 17224 -8632 17280 -7797
rect 17280 -8632 17284 -7797
rect 17220 -8637 17284 -8632
rect 17516 -6646 17580 -6641
rect 17516 -7481 17520 -6646
rect 17520 -7481 17576 -6646
rect 17576 -7481 17580 -6646
rect 17516 -8632 17520 -7797
rect 17520 -8632 17576 -7797
rect 17576 -8632 17580 -7797
rect 17516 -8637 17580 -8632
rect 17812 -6646 17876 -6641
rect 17812 -7481 17816 -6646
rect 17816 -7481 17872 -6646
rect 17872 -7481 17876 -6646
rect 17812 -8632 17816 -7797
rect 17816 -8632 17872 -7797
rect 17872 -8632 17876 -7797
rect 17812 -8637 17876 -8632
rect 18108 -6646 18172 -6641
rect 18108 -7481 18112 -6646
rect 18112 -7481 18168 -6646
rect 18168 -7481 18172 -6646
rect 18108 -8632 18112 -7797
rect 18112 -8632 18168 -7797
rect 18168 -8632 18172 -7797
rect 18108 -8637 18172 -8632
rect 18404 -6646 18468 -6641
rect 18404 -7481 18408 -6646
rect 18408 -7481 18464 -6646
rect 18464 -7481 18468 -6646
rect 18404 -8632 18408 -7797
rect 18408 -8632 18464 -7797
rect 18464 -8632 18468 -7797
rect 18404 -8637 18468 -8632
rect 18700 -6646 18764 -6641
rect 18700 -7481 18704 -6646
rect 18704 -7481 18760 -6646
rect 18760 -7481 18764 -6646
rect 18700 -8632 18704 -7797
rect 18704 -8632 18760 -7797
rect 18760 -8632 18764 -7797
rect 18700 -8637 18764 -8632
rect 18996 -6646 19060 -6641
rect 18996 -7481 19000 -6646
rect 19000 -7481 19056 -6646
rect 19056 -7481 19060 -6646
rect 18996 -8632 19000 -7797
rect 19000 -8632 19056 -7797
rect 19056 -8632 19060 -7797
rect 18996 -8637 19060 -8632
rect 19292 -6646 19356 -6641
rect 19292 -7481 19296 -6646
rect 19296 -7481 19352 -6646
rect 19352 -7481 19356 -6646
rect 19292 -8632 19296 -7797
rect 19296 -8632 19352 -7797
rect 19352 -8632 19356 -7797
rect 19292 -8637 19356 -8632
rect 19588 -6646 19652 -6641
rect 19588 -7481 19592 -6646
rect 19592 -7481 19648 -6646
rect 19648 -7481 19652 -6646
rect 19588 -8632 19592 -7797
rect 19592 -8632 19648 -7797
rect 19648 -8632 19652 -7797
rect 19588 -8637 19652 -8632
rect 19884 -6646 19948 -6641
rect 19884 -7481 19888 -6646
rect 19888 -7481 19944 -6646
rect 19944 -7481 19948 -6646
rect 19884 -8632 19888 -7797
rect 19888 -8632 19944 -7797
rect 19944 -8632 19948 -7797
rect 19884 -8637 19948 -8632
rect 20180 -6646 20244 -6641
rect 20180 -7481 20184 -6646
rect 20184 -7481 20240 -6646
rect 20240 -7481 20244 -6646
rect 20180 -8632 20184 -7797
rect 20184 -8632 20240 -7797
rect 20240 -8632 20244 -7797
rect 20180 -8637 20244 -8632
rect 20476 -6646 20540 -6641
rect 20476 -7481 20480 -6646
rect 20480 -7481 20536 -6646
rect 20536 -7481 20540 -6646
rect 20476 -8632 20480 -7797
rect 20480 -8632 20536 -7797
rect 20536 -8632 20540 -7797
rect 20476 -8637 20540 -8632
rect 20772 -6646 20836 -6641
rect 20772 -7481 20776 -6646
rect 20776 -7481 20832 -6646
rect 20832 -7481 20836 -6646
rect 20772 -8632 20776 -7797
rect 20776 -8632 20832 -7797
rect 20832 -8632 20836 -7797
rect 20772 -8637 20836 -8632
rect 21068 -6646 21132 -6641
rect 21068 -7481 21072 -6646
rect 21072 -7481 21128 -6646
rect 21128 -7481 21132 -6646
rect 21068 -8632 21072 -7797
rect 21072 -8632 21128 -7797
rect 21128 -8632 21132 -7797
rect 21068 -8637 21132 -8632
rect 21364 -6646 21428 -6641
rect 21364 -7481 21368 -6646
rect 21368 -7481 21424 -6646
rect 21424 -7481 21428 -6646
rect 21364 -8632 21368 -7797
rect 21368 -8632 21424 -7797
rect 21424 -8632 21428 -7797
rect 21364 -8637 21428 -8632
rect 21660 -6646 21724 -6641
rect 21660 -7481 21664 -6646
rect 21664 -7481 21720 -6646
rect 21720 -7481 21724 -6646
rect 21660 -8632 21664 -7797
rect 21664 -8632 21720 -7797
rect 21720 -8632 21724 -7797
rect 21660 -8637 21724 -8632
rect 21956 -6646 22020 -6641
rect 21956 -7481 21960 -6646
rect 21960 -7481 22016 -6646
rect 22016 -7481 22020 -6646
rect 21956 -8632 21960 -7797
rect 21960 -8632 22016 -7797
rect 22016 -8632 22020 -7797
rect 21956 -8637 22020 -8632
rect 22252 -6646 22316 -6641
rect 22252 -7481 22256 -6646
rect 22256 -7481 22312 -6646
rect 22312 -7481 22316 -6646
rect 22252 -8632 22256 -7797
rect 22256 -8632 22312 -7797
rect 22312 -8632 22316 -7797
rect 22252 -8637 22316 -8632
rect 22548 -6646 22612 -6641
rect 22548 -7481 22552 -6646
rect 22552 -7481 22608 -6646
rect 22608 -7481 22612 -6646
rect 22548 -8632 22552 -7797
rect 22552 -8632 22608 -7797
rect 22608 -8632 22612 -7797
rect 22548 -8637 22612 -8632
rect 23227 -7939 23231 -7104
rect 23231 -7939 23287 -7104
rect 23287 -7939 23291 -7104
rect 23227 -7944 23291 -7939
<< metal4 >>
rect 11590 -6641 11666 -5394
rect 11590 -7481 11596 -6641
rect 11660 -7481 11666 -6641
rect 11590 -7797 11666 -7481
rect 11590 -8637 11596 -7797
rect 11660 -8637 11666 -7797
rect 11590 -8639 11666 -8637
rect 11886 -6641 11962 -5595
rect 11886 -7481 11892 -6641
rect 11956 -7481 11962 -6641
rect 11886 -7797 11962 -7481
rect 11886 -8637 11892 -7797
rect 11956 -8637 11962 -7797
rect 11886 -8639 11962 -8637
rect 12182 -6641 12258 -5608
rect 12182 -7481 12188 -6641
rect 12252 -7481 12258 -6641
rect 12182 -7797 12258 -7481
rect 12182 -8637 12188 -7797
rect 12252 -8637 12258 -7797
rect 12182 -8639 12258 -8637
rect 12478 -6641 12554 -5394
rect 12478 -7481 12484 -6641
rect 12548 -7481 12554 -6641
rect 12478 -7797 12554 -7481
rect 12478 -8637 12484 -7797
rect 12548 -8637 12554 -7797
rect 12478 -8639 12554 -8637
rect 12774 -6641 12850 -5595
rect 12774 -7481 12780 -6641
rect 12844 -7481 12850 -6641
rect 12774 -7797 12850 -7481
rect 12774 -8637 12780 -7797
rect 12844 -8637 12850 -7797
rect 12774 -8639 12850 -8637
rect 13070 -6641 13146 -5608
rect 13070 -7481 13076 -6641
rect 13140 -7481 13146 -6641
rect 13070 -7797 13146 -7481
rect 13070 -8637 13076 -7797
rect 13140 -8637 13146 -7797
rect 13070 -8639 13146 -8637
rect 13366 -6641 13442 -5394
rect 13366 -7481 13372 -6641
rect 13436 -7481 13442 -6641
rect 13366 -7797 13442 -7481
rect 13366 -8637 13372 -7797
rect 13436 -8637 13442 -7797
rect 13366 -8639 13442 -8637
rect 13662 -6641 13738 -5595
rect 13662 -7481 13668 -6641
rect 13732 -7481 13738 -6641
rect 13662 -7797 13738 -7481
rect 13662 -8637 13668 -7797
rect 13732 -8637 13738 -7797
rect 13662 -8639 13738 -8637
rect 13958 -6641 14034 -5608
rect 13958 -7481 13964 -6641
rect 14028 -7481 14034 -6641
rect 13958 -7797 14034 -7481
rect 13958 -8637 13964 -7797
rect 14028 -8637 14034 -7797
rect 13958 -8639 14034 -8637
rect 14254 -6641 14330 -5394
rect 14254 -7481 14260 -6641
rect 14324 -7481 14330 -6641
rect 14254 -7797 14330 -7481
rect 14254 -8637 14260 -7797
rect 14324 -8637 14330 -7797
rect 14254 -8639 14330 -8637
rect 14550 -6641 14626 -5394
rect 14550 -7481 14556 -6641
rect 14620 -7481 14626 -6641
rect 14550 -7797 14626 -7481
rect 14550 -8637 14556 -7797
rect 14620 -8637 14626 -7797
rect 14550 -8639 14626 -8637
rect 14846 -6641 14922 -5998
rect 14846 -7481 14852 -6641
rect 14916 -7481 14922 -6641
rect 14846 -7797 14922 -7481
rect 14846 -8637 14852 -7797
rect 14916 -8637 14922 -7797
rect 14846 -8639 14922 -8637
rect 15142 -6641 15218 -5910
rect 15142 -7481 15148 -6641
rect 15212 -7481 15218 -6641
rect 15142 -7797 15218 -7481
rect 15142 -8637 15148 -7797
rect 15212 -8637 15218 -7797
rect 15142 -8639 15218 -8637
rect 15438 -6641 15514 -5394
rect 15438 -7481 15444 -6641
rect 15508 -7481 15514 -6641
rect 15438 -7797 15514 -7481
rect 15438 -8637 15444 -7797
rect 15508 -8637 15514 -7797
rect 15438 -8639 15514 -8637
rect 15734 -6641 15810 -5595
rect 15734 -7481 15740 -6641
rect 15804 -7481 15810 -6641
rect 15734 -7797 15810 -7481
rect 15734 -8637 15740 -7797
rect 15804 -8637 15810 -7797
rect 15734 -8639 15810 -8637
rect 16030 -6641 16106 -5608
rect 16030 -7481 16036 -6641
rect 16100 -7481 16106 -6641
rect 16030 -7797 16106 -7481
rect 16030 -8637 16036 -7797
rect 16100 -8637 16106 -7797
rect 16030 -8639 16106 -8637
rect 16326 -6641 16402 -5394
rect 16326 -7481 16332 -6641
rect 16396 -7481 16402 -6641
rect 16326 -7797 16402 -7481
rect 16326 -8637 16332 -7797
rect 16396 -8637 16402 -7797
rect 16326 -8639 16402 -8637
rect 16622 -6641 16698 -5595
rect 16622 -7481 16628 -6641
rect 16692 -7481 16698 -6641
rect 16622 -7797 16698 -7481
rect 16622 -8637 16628 -7797
rect 16692 -8637 16698 -7797
rect 16622 -8639 16698 -8637
rect 16918 -6641 16994 -5608
rect 16918 -7481 16924 -6641
rect 16988 -7481 16994 -6641
rect 16918 -7797 16994 -7481
rect 16918 -8637 16924 -7797
rect 16988 -8637 16994 -7797
rect 16918 -8639 16994 -8637
rect 17214 -6641 17290 -5394
rect 17214 -7481 17220 -6641
rect 17284 -7481 17290 -6641
rect 17214 -7797 17290 -7481
rect 17214 -8637 17220 -7797
rect 17284 -8637 17290 -7797
rect 17214 -8639 17290 -8637
rect 17510 -6641 17586 -5394
rect 17510 -7481 17516 -6641
rect 17580 -7481 17586 -6641
rect 17510 -7797 17586 -7481
rect 17510 -8637 17516 -7797
rect 17580 -8637 17586 -7797
rect 17510 -8639 17586 -8637
rect 17806 -6641 17882 -5595
rect 17806 -7481 17812 -6641
rect 17876 -7481 17882 -6641
rect 17806 -7797 17882 -7481
rect 17806 -8637 17812 -7797
rect 17876 -8637 17882 -7797
rect 17806 -8639 17882 -8637
rect 18102 -6641 18178 -5608
rect 18102 -7481 18108 -6641
rect 18172 -7481 18178 -6641
rect 18102 -7797 18178 -7481
rect 18102 -8637 18108 -7797
rect 18172 -8637 18178 -7797
rect 18102 -8639 18178 -8637
rect 18398 -6641 18474 -5394
rect 18398 -7481 18404 -6641
rect 18468 -7481 18474 -6641
rect 18398 -7797 18474 -7481
rect 18398 -8637 18404 -7797
rect 18468 -8637 18474 -7797
rect 18398 -8639 18474 -8637
rect 18694 -6641 18770 -6019
rect 18694 -7481 18700 -6641
rect 18764 -7481 18770 -6641
rect 18694 -7797 18770 -7481
rect 18694 -8637 18700 -7797
rect 18764 -8637 18770 -7797
rect 18694 -8639 18770 -8637
rect 18990 -6641 19066 -5896
rect 18990 -7481 18996 -6641
rect 19060 -7481 19066 -6641
rect 18990 -7797 19066 -7481
rect 18990 -8637 18996 -7797
rect 19060 -8637 19066 -7797
rect 18990 -8639 19066 -8637
rect 19286 -6641 19362 -5394
rect 19286 -7481 19292 -6641
rect 19356 -7481 19362 -6641
rect 19286 -7797 19362 -7481
rect 19286 -8637 19292 -7797
rect 19356 -8637 19362 -7797
rect 19286 -8639 19362 -8637
rect 19582 -6641 19658 -5394
rect 19582 -7481 19588 -6641
rect 19652 -7481 19658 -6641
rect 19582 -7797 19658 -7481
rect 19582 -8637 19588 -7797
rect 19652 -8637 19658 -7797
rect 19582 -8639 19658 -8637
rect 19878 -6641 19954 -5595
rect 19878 -7481 19884 -6641
rect 19948 -7481 19954 -6641
rect 19878 -7797 19954 -7481
rect 19878 -8637 19884 -7797
rect 19948 -8637 19954 -7797
rect 19878 -8639 19954 -8637
rect 20174 -6641 20250 -5394
rect 20174 -7481 20180 -6641
rect 20244 -7481 20250 -6641
rect 20174 -7797 20250 -7481
rect 20174 -8637 20180 -7797
rect 20244 -8637 20250 -7797
rect 20174 -8639 20250 -8637
rect 20470 -6641 20546 -5394
rect 20470 -7481 20476 -6641
rect 20540 -7481 20546 -6641
rect 20470 -7797 20546 -7481
rect 20470 -8637 20476 -7797
rect 20540 -8637 20546 -7797
rect 20470 -8639 20546 -8637
rect 20766 -6641 20842 -5595
rect 20766 -7481 20772 -6641
rect 20836 -7481 20842 -6641
rect 20766 -7797 20842 -7481
rect 20766 -8637 20772 -7797
rect 20836 -8637 20842 -7797
rect 20766 -8639 20842 -8637
rect 21062 -6641 21138 -5608
rect 21062 -7481 21068 -6641
rect 21132 -7481 21138 -6641
rect 21062 -7797 21138 -7481
rect 21062 -8637 21068 -7797
rect 21132 -8637 21138 -7797
rect 21062 -8639 21138 -8637
rect 21358 -6641 21434 -5394
rect 21358 -7481 21364 -6641
rect 21428 -7481 21434 -6641
rect 21358 -7797 21434 -7481
rect 21358 -8637 21364 -7797
rect 21428 -8637 21434 -7797
rect 21358 -8639 21434 -8637
rect 21654 -6641 21730 -5595
rect 21654 -7481 21660 -6641
rect 21724 -7481 21730 -6641
rect 21654 -7797 21730 -7481
rect 21654 -8637 21660 -7797
rect 21724 -8637 21730 -7797
rect 21654 -8639 21730 -8637
rect 21950 -6641 22026 -5608
rect 21950 -7481 21956 -6641
rect 22020 -7481 22026 -6641
rect 21950 -7797 22026 -7481
rect 21950 -8637 21956 -7797
rect 22020 -8637 22026 -7797
rect 21950 -8639 22026 -8637
rect 22246 -6641 22322 -5394
rect 22246 -7481 22252 -6641
rect 22316 -7481 22322 -6641
rect 22246 -7797 22322 -7481
rect 22246 -8637 22252 -7797
rect 22316 -8637 22322 -7797
rect 22246 -8639 22322 -8637
rect 22542 -6641 22618 -5595
rect 22542 -7481 22548 -6641
rect 22612 -7481 22618 -6641
rect 22542 -7797 22618 -7481
rect 22542 -8637 22548 -7797
rect 22612 -8637 22618 -7797
rect 23226 -7104 23292 -7103
rect 23226 -7944 23227 -7104
rect 23291 -7944 23292 -7104
rect 23226 -7945 23292 -7944
rect 22542 -8639 22618 -8637
use sky130_fd_pr__nfet_01v8_M4T2ST  sky130_fd_pr__nfet_01v8_M4T2ST_0
timestamp 1606612150
transform 1 0 9823 0 1 -6885
box -285 -510 285 510
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_2
timestamp 1606520558
transform -1 0 16890 0 1 -4228
box -1941 -1600 1941 1600
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_3
timestamp 1606520558
transform -1 0 12851 0 1 -4228
box -1941 -1600 1941 1600
use sky130_fd_pr__nfet_01v8_8JUMX6  sky130_fd_pr__nfet_01v8_8JUMX6_0
timestamp 1606595467
transform 1 0 17030 0 1 -7639
box -5717 -1219 5717 1219
use sky130_fd_pr__nfet_01v8_8HUREQ  sky130_fd_pr__nfet_01v8_8HUREQ_1
timestamp 1606416512
transform 1 0 5916 0 1 -7838
box -1052 -919 1052 919
use sky130_fd_pr__pfet_01v8_YCMRKB  sky130_fd_pr__pfet_01v8_YCMRKB_3
timestamp 1606513430
transform 1 0 4257 0 1 -5523
box -3117 -937 3117 937
use sky130_fd_pr__nfet_01v8_8HUREQ  sky130_fd_pr__nfet_01v8_8HUREQ_0
timestamp 1606416512
transform 1 0 3918 0 1 -7838
box -1052 -919 1052 919
use sky130_fd_pr__pfet_01v8_YCMRKB  sky130_fd_pr__pfet_01v8_YCMRKB_2
timestamp 1606513430
transform 1 0 4257 0 1 -3755
box -3117 -937 3117 937
use sky130_fd_pr__pfet_01v8_YCMRKB  sky130_fd_pr__pfet_01v8_YCMRKB_0
timestamp 1606513430
transform 1 0 4257 0 1 -1987
box -3117 -937 3117 937
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_1
timestamp 1606520558
transform -1 0 16890 0 1 -820
box -1941 -1600 1941 1600
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_0
timestamp 1606520558
transform -1 0 12851 0 1 -820
box -1941 -1600 1941 1600
use sky130_fd_pr__pfet_01v8_YCMRKB  sky130_fd_pr__pfet_01v8_YCMRKB_1
timestamp 1606513430
transform 1 0 4257 0 1 -219
box -3117 -937 3117 937
use sky130_fd_pr__pfet_01v8_YC99EG  sky130_fd_pr__pfet_01v8_YC99EG_0
timestamp 1606509736
transform 1 0 16942 0 1 1968
box -4592 -937 4592 937
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_5
timestamp 1606520558
transform -1 0 20941 0 1 -820
box -1941 -1600 1941 1600
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_4
timestamp 1606520558
transform -1 0 20941 0 1 -4228
box -1941 -1600 1941 1600
use sky130_fd_pr__pfet_01v8_YC9MKB  sky130_fd_pr__pfet_01v8_YC9MKB_2
timestamp 1606509736
transform 1 0 9452 0 1 2387
box -1052 -519 1052 519
use sky130_fd_pr__pfet_01v8_YC9MKB  sky130_fd_pr__pfet_01v8_YC9MKB_1
timestamp 1606509736
transform 1 0 7454 0 1 2387
box -1052 -519 1052 519
use sky130_fd_pr__pfet_01v8_YC9MKB  sky130_fd_pr__pfet_01v8_YC9MKB_0
timestamp 1606509736
transform 1 0 5456 0 1 2387
box -1052 -519 1052 519
<< labels >>
rlabel metal2 12325 1931 12372 1992 1 iref
<< end >>
