magic
tech sky130A
magscale 1 2
timestamp 1605064714
<< viali >>
rect 3433 19593 3467 19627
rect 1409 19525 1443 19559
rect 1685 19457 1719 19491
rect 2145 19049 2179 19083
rect 4077 18981 4111 19015
rect 4353 18981 4387 19015
rect 6101 18981 6135 19015
rect 2329 18845 2363 18879
rect 5549 18641 5583 18675
rect 1685 18505 1719 18539
rect 1409 18437 1443 18471
rect 3433 18437 3467 18471
rect 4261 18437 4295 18471
rect 5365 18437 5399 18471
rect 4445 18301 4479 18335
rect 1961 18097 1995 18131
rect 4353 18029 4387 18063
rect 1777 17961 1811 17995
rect 2881 17961 2915 17995
rect 4077 17893 4111 17927
rect 6101 17893 6135 17927
rect 3065 17757 3099 17791
rect 1685 17417 1719 17451
rect 3433 17417 3467 17451
rect 1409 17349 1443 17383
rect 4169 16873 4203 16907
rect 4537 16805 4571 16839
rect 7113 16805 7147 16839
rect 6285 16669 6319 16703
rect 3433 16329 3467 16363
rect 3157 16261 3191 16295
rect 5181 16193 5215 16227
rect 5273 15921 5307 15955
rect 5089 15785 5123 15819
rect 6193 15785 6227 15819
rect 7389 15785 7423 15819
rect 7205 15717 7239 15751
rect 1409 15241 1443 15275
rect 4445 15241 4479 15275
rect 5825 15241 5859 15275
rect 4997 15173 5031 15207
rect 5181 15173 5215 15207
rect 5365 15173 5399 15207
rect 5733 15173 5767 15207
rect 7573 15173 7607 15207
rect 1685 15105 1719 15139
rect 3433 15105 3467 15139
rect 7665 15037 7699 15071
rect 4353 14765 4387 14799
rect 2145 14697 2179 14731
rect 4077 14697 4111 14731
rect 7021 14697 7055 14731
rect 7389 14697 7423 14731
rect 7665 14697 7699 14731
rect 6101 14629 6135 14663
rect 2329 14493 2363 14527
rect 6929 14289 6963 14323
rect 3433 14153 3467 14187
rect 5825 14153 5859 14187
rect 1409 14085 1443 14119
rect 4445 14085 4479 14119
rect 4997 14085 5031 14119
rect 5181 14085 5215 14119
rect 5365 14085 5399 14119
rect 5733 14085 5767 14119
rect 7113 14085 7147 14119
rect 7389 14085 7423 14119
rect 1685 14017 1719 14051
rect 7481 13745 7515 13779
rect 4537 13677 4571 13711
rect 3249 13609 3283 13643
rect 7205 13609 7239 13643
rect 7389 13609 7423 13643
rect 4261 13541 4295 13575
rect 6285 13541 6319 13575
rect 3065 13405 3099 13439
rect 7297 13201 7331 13235
rect 2237 13065 2271 13099
rect 3985 13065 4019 13099
rect 1961 12997 1995 13031
rect 4813 12997 4847 13031
rect 6929 12997 6963 13031
rect 7113 12997 7147 13031
rect 7021 12929 7055 12963
rect 4997 12861 5031 12895
rect 3065 12657 3099 12691
rect 4261 12657 4295 12691
rect 2881 12521 2915 12555
rect 4077 12521 4111 12555
rect 5181 12453 5215 12487
rect 5549 12453 5583 12487
rect 6929 12453 6963 12487
rect 2973 12113 3007 12147
rect 6929 12113 6963 12147
rect 3893 11977 3927 12011
rect 4169 11977 4203 12011
rect 2789 11909 2823 11943
rect 5917 11909 5951 11943
rect 6837 11909 6871 11943
rect 2329 11569 2363 11603
rect 5273 11569 5307 11603
rect 6377 11569 6411 11603
rect 2145 11433 2179 11467
rect 5089 11433 5123 11467
rect 6193 11433 6227 11467
rect 1409 10889 1443 10923
rect 3433 10889 3467 10923
rect 1685 10753 1719 10787
rect 4261 10753 4295 10787
rect 5549 10685 5583 10719
rect 2237 10345 2271 10379
rect 2421 10209 2455 10243
rect 1409 9801 1443 9835
rect 3433 9801 3467 9835
rect 7205 9733 7239 9767
rect 7297 9733 7331 9767
rect 1685 9665 1719 9699
rect 7757 9665 7791 9699
rect 1961 9393 1995 9427
rect 1777 9257 1811 9291
rect 2881 9257 2915 9291
rect 5457 9257 5491 9291
rect 5089 9189 5123 9223
rect 6837 9189 6871 9223
rect 3065 9053 3099 9087
rect 7021 8849 7055 8883
rect 4537 8713 4571 8747
rect 2513 8645 2547 8679
rect 5365 8645 5399 8679
rect 6837 8645 6871 8679
rect 2789 8577 2823 8611
rect 5549 8509 5583 8543
rect 3065 8305 3099 8339
rect 7481 8305 7515 8339
rect 6469 8237 6503 8271
rect 2789 8169 2823 8203
rect 2881 8169 2915 8203
rect 7303 8169 7337 8203
rect 4445 8101 4479 8135
rect 4721 8101 4755 8135
rect 2605 8033 2639 8067
rect 5733 7761 5767 7795
rect 4629 7693 4663 7727
rect 3341 7557 3375 7591
rect 4445 7557 4479 7591
rect 5549 7557 5583 7591
rect 3525 7421 3559 7455
rect 6377 7149 6411 7183
rect 4353 7013 4387 7047
rect 4629 7013 4663 7047
rect 5549 6673 5583 6707
rect 1409 6469 1443 6503
rect 4261 6469 4295 6503
rect 5365 6469 5399 6503
rect 1685 6401 1719 6435
rect 3433 6401 3467 6435
rect 4445 6333 4479 6367
rect 2145 5993 2179 6027
rect 2329 5789 2363 5823
rect 1409 5449 1443 5483
rect 1685 5449 1719 5483
rect 3433 5313 3467 5347
rect 2421 5041 2455 5075
rect 4353 4973 4387 5007
rect 2237 4905 2271 4939
rect 4077 4905 4111 4939
rect 6101 4837 6135 4871
rect 4629 4361 4663 4395
rect 2605 4293 2639 4327
rect 2881 4225 2915 4259
rect 3065 3953 3099 3987
rect 4353 3885 4387 3919
rect 2881 3817 2915 3851
rect 4077 3749 4111 3783
rect 6101 3749 6135 3783
rect 1672 3409 1706 3443
rect 5273 3409 5307 3443
rect 1409 3273 1443 3307
rect 5181 3205 5215 3239
rect 6837 3205 6871 3239
rect 3433 3137 3467 3171
rect 4997 3137 5031 3171
rect 6929 3069 6963 3103
rect 3065 2865 3099 2899
rect 2881 2729 2915 2763
rect 4997 2729 5031 2763
rect 5089 2729 5123 2763
rect 5273 2525 5307 2559
rect 4537 2321 4571 2355
rect 4353 2117 4387 2151
<< metal1 >>
rect 4062 22644 4068 22696
rect 4120 22684 4126 22696
rect 5166 22684 5172 22696
rect 4120 22656 5172 22684
rect 4120 22644 4126 22656
rect 5166 22644 5172 22656
rect 5224 22644 5230 22696
rect 1104 21506 8832 21528
rect 1104 21454 3579 21506
rect 3631 21454 3643 21506
rect 3695 21454 3707 21506
rect 3759 21454 3771 21506
rect 3823 21454 6176 21506
rect 6228 21454 6240 21506
rect 6292 21454 6304 21506
rect 6356 21454 6368 21506
rect 6420 21454 8832 21506
rect 1104 21432 8832 21454
rect 1104 20962 8832 20984
rect 1104 20910 2280 20962
rect 2332 20910 2344 20962
rect 2396 20910 2408 20962
rect 2460 20910 2472 20962
rect 2524 20910 4878 20962
rect 4930 20910 4942 20962
rect 4994 20910 5006 20962
rect 5058 20910 5070 20962
rect 5122 20910 7475 20962
rect 7527 20910 7539 20962
rect 7591 20910 7603 20962
rect 7655 20910 7667 20962
rect 7719 20910 8832 20962
rect 1104 20888 8832 20910
rect 1104 20418 8832 20440
rect 1104 20366 3579 20418
rect 3631 20366 3643 20418
rect 3695 20366 3707 20418
rect 3759 20366 3771 20418
rect 3823 20366 6176 20418
rect 6228 20366 6240 20418
rect 6292 20366 6304 20418
rect 6356 20366 6368 20418
rect 6420 20366 8832 20418
rect 1104 20344 8832 20366
rect 1104 19874 8832 19896
rect 1104 19822 2280 19874
rect 2332 19822 2344 19874
rect 2396 19822 2408 19874
rect 2460 19822 2472 19874
rect 2524 19822 4878 19874
rect 4930 19822 4942 19874
rect 4994 19822 5006 19874
rect 5058 19822 5070 19874
rect 5122 19822 7475 19874
rect 7527 19822 7539 19874
rect 7591 19822 7603 19874
rect 7655 19822 7667 19874
rect 7719 19822 8832 19874
rect 1104 19800 8832 19822
rect 3418 19624 3424 19636
rect 3379 19596 3424 19624
rect 3418 19584 3424 19596
rect 3476 19584 3482 19636
rect 1394 19556 1400 19568
rect 1355 19528 1400 19556
rect 1394 19516 1400 19528
rect 1452 19516 1458 19568
rect 1673 19491 1731 19497
rect 1673 19457 1685 19491
rect 1719 19457 1731 19491
rect 1673 19451 1731 19457
rect 1688 19420 1716 19451
rect 1946 19448 1952 19500
rect 2004 19488 2010 19500
rect 2004 19460 2162 19488
rect 2004 19448 2010 19460
rect 3326 19420 3332 19432
rect 1688 19392 3332 19420
rect 3326 19380 3332 19392
rect 3384 19380 3390 19432
rect 1104 19330 8832 19352
rect 1104 19278 3579 19330
rect 3631 19278 3643 19330
rect 3695 19278 3707 19330
rect 3759 19278 3771 19330
rect 3823 19278 6176 19330
rect 6228 19278 6240 19330
rect 6292 19278 6304 19330
rect 6356 19278 6368 19330
rect 6420 19278 8832 19330
rect 1104 19256 8832 19278
rect 1762 19040 1768 19092
rect 1820 19080 1826 19092
rect 2133 19083 2191 19089
rect 2133 19080 2145 19083
rect 1820 19052 2145 19080
rect 1820 19040 1826 19052
rect 2133 19049 2145 19052
rect 2179 19049 2191 19083
rect 5474 19052 5580 19080
rect 2133 19043 2191 19049
rect 5552 19024 5580 19052
rect 4062 19012 4068 19024
rect 4023 18984 4068 19012
rect 4062 18972 4068 18984
rect 4120 18972 4126 19024
rect 4341 19015 4399 19021
rect 4341 18981 4353 19015
rect 4387 19012 4399 19015
rect 5350 19012 5356 19024
rect 4387 18984 5356 19012
rect 4387 18981 4399 18984
rect 4341 18975 4399 18981
rect 5350 18972 5356 18984
rect 5408 18972 5414 19024
rect 5534 18972 5540 19024
rect 5592 18972 5598 19024
rect 6089 19015 6147 19021
rect 6089 18981 6101 19015
rect 6135 18981 6147 19015
rect 6089 18975 6147 18981
rect 2130 18836 2136 18888
rect 2188 18876 2194 18888
rect 2317 18879 2375 18885
rect 2317 18876 2329 18879
rect 2188 18848 2329 18876
rect 2188 18836 2194 18848
rect 2317 18845 2329 18848
rect 2363 18845 2375 18879
rect 2317 18839 2375 18845
rect 2682 18836 2688 18888
rect 2740 18876 2746 18888
rect 6104 18876 6132 18975
rect 2740 18848 6132 18876
rect 2740 18836 2746 18848
rect 1104 18786 8832 18808
rect 1104 18734 2280 18786
rect 2332 18734 2344 18786
rect 2396 18734 2408 18786
rect 2460 18734 2472 18786
rect 2524 18734 4878 18786
rect 4930 18734 4942 18786
rect 4994 18734 5006 18786
rect 5058 18734 5070 18786
rect 5122 18734 7475 18786
rect 7527 18734 7539 18786
rect 7591 18734 7603 18786
rect 7655 18734 7667 18786
rect 7719 18734 8832 18786
rect 1104 18712 8832 18734
rect 5534 18672 5540 18684
rect 5495 18644 5540 18672
rect 5534 18632 5540 18644
rect 5592 18632 5598 18684
rect 1670 18536 1676 18548
rect 1583 18508 1676 18536
rect 1670 18496 1676 18508
rect 1728 18536 1734 18548
rect 2682 18536 2688 18548
rect 1728 18508 2688 18536
rect 1728 18496 1734 18508
rect 2682 18496 2688 18508
rect 2740 18496 2746 18548
rect 1394 18468 1400 18480
rect 1355 18440 1400 18468
rect 1394 18428 1400 18440
rect 1452 18428 1458 18480
rect 3050 18428 3056 18480
rect 3108 18468 3114 18480
rect 3421 18471 3479 18477
rect 3421 18468 3433 18471
rect 3108 18440 3433 18468
rect 3108 18428 3114 18440
rect 3421 18437 3433 18440
rect 3467 18437 3479 18471
rect 3421 18431 3479 18437
rect 4249 18471 4307 18477
rect 4249 18437 4261 18471
rect 4295 18468 4307 18471
rect 4522 18468 4528 18480
rect 4295 18440 4528 18468
rect 4295 18437 4307 18440
rect 4249 18431 4307 18437
rect 4522 18428 4528 18440
rect 4580 18468 4586 18480
rect 5353 18471 5411 18477
rect 5353 18468 5365 18471
rect 4580 18440 5365 18468
rect 4580 18428 4586 18440
rect 5353 18437 5365 18440
rect 5399 18437 5411 18471
rect 5353 18431 5411 18437
rect 2130 18360 2136 18412
rect 2188 18360 2194 18412
rect 4430 18332 4436 18344
rect 4391 18304 4436 18332
rect 4430 18292 4436 18304
rect 4488 18292 4494 18344
rect 1104 18242 8832 18264
rect 1104 18190 3579 18242
rect 3631 18190 3643 18242
rect 3695 18190 3707 18242
rect 3759 18190 3771 18242
rect 3823 18190 6176 18242
rect 6228 18190 6240 18242
rect 6292 18190 6304 18242
rect 6356 18190 6368 18242
rect 6420 18190 8832 18242
rect 1104 18168 8832 18190
rect 1946 18128 1952 18140
rect 1907 18100 1952 18128
rect 1946 18088 1952 18100
rect 2004 18088 2010 18140
rect 4522 18128 4528 18140
rect 2884 18100 4528 18128
rect 1762 17992 1768 18004
rect 1723 17964 1768 17992
rect 1762 17952 1768 17964
rect 1820 17952 1826 18004
rect 2884 18001 2912 18100
rect 4522 18088 4528 18100
rect 4580 18088 4586 18140
rect 3326 18020 3332 18072
rect 3384 18060 3390 18072
rect 4341 18063 4399 18069
rect 4341 18060 4353 18063
rect 3384 18032 4353 18060
rect 3384 18020 3390 18032
rect 4341 18029 4353 18032
rect 4387 18029 4399 18063
rect 4341 18023 4399 18029
rect 4430 18020 4436 18072
rect 4488 18060 4494 18072
rect 4488 18032 4830 18060
rect 4488 18020 4494 18032
rect 2869 17995 2927 18001
rect 2869 17961 2881 17995
rect 2915 17961 2927 17995
rect 2869 17955 2927 17961
rect 2958 17884 2964 17936
rect 3016 17924 3022 17936
rect 4062 17924 4068 17936
rect 3016 17896 4068 17924
rect 3016 17884 3022 17896
rect 4062 17884 4068 17896
rect 4120 17884 4126 17936
rect 4706 17884 4712 17936
rect 4764 17924 4770 17936
rect 6089 17927 6147 17933
rect 6089 17924 6101 17927
rect 4764 17896 6101 17924
rect 4764 17884 4770 17896
rect 6089 17893 6101 17896
rect 6135 17893 6147 17927
rect 6089 17887 6147 17893
rect 3050 17788 3056 17800
rect 3011 17760 3056 17788
rect 3050 17748 3056 17760
rect 3108 17748 3114 17800
rect 1104 17698 8832 17720
rect 1104 17646 2280 17698
rect 2332 17646 2344 17698
rect 2396 17646 2408 17698
rect 2460 17646 2472 17698
rect 2524 17646 4878 17698
rect 4930 17646 4942 17698
rect 4994 17646 5006 17698
rect 5058 17646 5070 17698
rect 5122 17646 7475 17698
rect 7527 17646 7539 17698
rect 7591 17646 7603 17698
rect 7655 17646 7667 17698
rect 7719 17646 8832 17698
rect 1104 17624 8832 17646
rect 1394 17544 1400 17596
rect 1452 17584 1458 17596
rect 3418 17584 3424 17596
rect 1452 17556 3424 17584
rect 1452 17544 1458 17556
rect 3418 17544 3424 17556
rect 3476 17544 3482 17596
rect 1670 17448 1676 17460
rect 1631 17420 1676 17448
rect 1670 17408 1676 17420
rect 1728 17408 1734 17460
rect 3326 17408 3332 17460
rect 3384 17448 3390 17460
rect 3421 17451 3479 17457
rect 3421 17448 3433 17451
rect 3384 17420 3433 17448
rect 3384 17408 3390 17420
rect 3421 17417 3433 17420
rect 3467 17417 3479 17451
rect 3421 17411 3479 17417
rect 1397 17383 1455 17389
rect 1397 17349 1409 17383
rect 1443 17349 1455 17383
rect 3050 17380 3056 17392
rect 2806 17352 3056 17380
rect 1397 17343 1455 17349
rect 1412 17244 1440 17343
rect 3050 17340 3056 17352
rect 3108 17340 3114 17392
rect 2958 17244 2964 17256
rect 1412 17216 2964 17244
rect 2958 17204 2964 17216
rect 3016 17204 3022 17256
rect 1104 17154 8832 17176
rect 1104 17102 3579 17154
rect 3631 17102 3643 17154
rect 3695 17102 3707 17154
rect 3759 17102 3771 17154
rect 3823 17102 6176 17154
rect 6228 17102 6240 17154
rect 6292 17102 6304 17154
rect 6356 17102 6368 17154
rect 6420 17102 8832 17154
rect 1104 17080 8832 17102
rect 5258 16932 5264 16984
rect 5316 16932 5322 16984
rect 3418 16864 3424 16916
rect 3476 16904 3482 16916
rect 4157 16907 4215 16913
rect 4157 16904 4169 16907
rect 3476 16876 4169 16904
rect 3476 16864 3482 16876
rect 4157 16873 4169 16876
rect 4203 16873 4215 16907
rect 4157 16867 4215 16873
rect 4525 16839 4583 16845
rect 4525 16805 4537 16839
rect 4571 16836 4583 16839
rect 4706 16836 4712 16848
rect 4571 16808 4712 16836
rect 4571 16805 4583 16808
rect 4525 16799 4583 16805
rect 4706 16796 4712 16808
rect 4764 16796 4770 16848
rect 7098 16836 7104 16848
rect 7059 16808 7104 16836
rect 7098 16796 7104 16808
rect 7156 16796 7162 16848
rect 6273 16703 6331 16709
rect 6273 16669 6285 16703
rect 6319 16700 6331 16703
rect 6638 16700 6644 16712
rect 6319 16672 6644 16700
rect 6319 16669 6331 16672
rect 6273 16663 6331 16669
rect 6638 16660 6644 16672
rect 6696 16660 6702 16712
rect 1104 16610 8832 16632
rect 1104 16558 2280 16610
rect 2332 16558 2344 16610
rect 2396 16558 2408 16610
rect 2460 16558 2472 16610
rect 2524 16558 4878 16610
rect 4930 16558 4942 16610
rect 4994 16558 5006 16610
rect 5058 16558 5070 16610
rect 5122 16558 7475 16610
rect 7527 16558 7539 16610
rect 7591 16558 7603 16610
rect 7655 16558 7667 16610
rect 7719 16558 8832 16610
rect 1104 16536 8832 16558
rect 3421 16363 3479 16369
rect 3421 16329 3433 16363
rect 3467 16360 3479 16363
rect 4706 16360 4712 16372
rect 3467 16332 4712 16360
rect 3467 16329 3479 16332
rect 3421 16323 3479 16329
rect 4706 16320 4712 16332
rect 4764 16320 4770 16372
rect 2866 16252 2872 16304
rect 2924 16292 2930 16304
rect 3145 16295 3203 16301
rect 3145 16292 3157 16295
rect 2924 16264 3157 16292
rect 2924 16252 2930 16264
rect 3145 16261 3157 16264
rect 3191 16261 3203 16295
rect 3145 16255 3203 16261
rect 4522 16252 4528 16304
rect 4580 16252 4586 16304
rect 5166 16224 5172 16236
rect 5127 16196 5172 16224
rect 5166 16184 5172 16196
rect 5224 16184 5230 16236
rect 1104 16066 8832 16088
rect 1104 16014 3579 16066
rect 3631 16014 3643 16066
rect 3695 16014 3707 16066
rect 3759 16014 3771 16066
rect 3823 16014 6176 16066
rect 6228 16014 6240 16066
rect 6292 16014 6304 16066
rect 6356 16014 6368 16066
rect 6420 16014 8832 16066
rect 1104 15992 8832 16014
rect 5258 15952 5264 15964
rect 5219 15924 5264 15952
rect 5258 15912 5264 15924
rect 5316 15912 5322 15964
rect 4706 15776 4712 15828
rect 4764 15816 4770 15828
rect 5077 15819 5135 15825
rect 5077 15816 5089 15819
rect 4764 15788 5089 15816
rect 4764 15776 4770 15788
rect 5077 15785 5089 15788
rect 5123 15785 5135 15819
rect 5077 15779 5135 15785
rect 6181 15819 6239 15825
rect 6181 15785 6193 15819
rect 6227 15816 6239 15819
rect 7098 15816 7104 15828
rect 6227 15788 7104 15816
rect 6227 15785 6239 15788
rect 6181 15779 6239 15785
rect 7098 15776 7104 15788
rect 7156 15776 7162 15828
rect 7374 15816 7380 15828
rect 7335 15788 7380 15816
rect 7374 15776 7380 15788
rect 7432 15776 7438 15828
rect 6822 15708 6828 15760
rect 6880 15748 6886 15760
rect 7193 15751 7251 15757
rect 7193 15748 7205 15751
rect 6880 15720 7205 15748
rect 6880 15708 6886 15720
rect 7193 15717 7205 15720
rect 7239 15717 7251 15751
rect 7193 15711 7251 15717
rect 1104 15522 8832 15544
rect 1104 15470 2280 15522
rect 2332 15470 2344 15522
rect 2396 15470 2408 15522
rect 2460 15470 2472 15522
rect 2524 15470 4878 15522
rect 4930 15470 4942 15522
rect 4994 15470 5006 15522
rect 5058 15470 5070 15522
rect 5122 15470 7475 15522
rect 7527 15470 7539 15522
rect 7591 15470 7603 15522
rect 7655 15470 7667 15522
rect 7719 15470 8832 15522
rect 1104 15448 8832 15470
rect 5902 15340 5908 15352
rect 5644 15312 5908 15340
rect 1397 15275 1455 15281
rect 1397 15241 1409 15275
rect 1443 15272 1455 15275
rect 2866 15272 2872 15284
rect 1443 15244 2872 15272
rect 1443 15241 1455 15244
rect 1397 15235 1455 15241
rect 2866 15232 2872 15244
rect 2924 15232 2930 15284
rect 4154 15232 4160 15284
rect 4212 15272 4218 15284
rect 4433 15275 4491 15281
rect 4433 15272 4445 15275
rect 4212 15244 4445 15272
rect 4212 15232 4218 15244
rect 4433 15241 4445 15244
rect 4479 15241 4491 15275
rect 5534 15272 5540 15284
rect 4433 15235 4491 15241
rect 5184 15244 5540 15272
rect 5184 15213 5212 15244
rect 5534 15232 5540 15244
rect 5592 15232 5598 15284
rect 4985 15207 5043 15213
rect 4985 15173 4997 15207
rect 5031 15173 5043 15207
rect 4985 15167 5043 15173
rect 5169 15207 5227 15213
rect 5169 15173 5181 15207
rect 5215 15173 5227 15207
rect 5169 15167 5227 15173
rect 5353 15207 5411 15213
rect 5353 15173 5365 15207
rect 5399 15204 5411 15207
rect 5644 15204 5672 15312
rect 5902 15300 5908 15312
rect 5960 15300 5966 15352
rect 5810 15272 5816 15284
rect 5771 15244 5816 15272
rect 5810 15232 5816 15244
rect 5868 15232 5874 15284
rect 5399 15176 5672 15204
rect 5721 15207 5779 15213
rect 5399 15173 5411 15176
rect 5353 15167 5411 15173
rect 5721 15173 5733 15207
rect 5767 15173 5779 15207
rect 5721 15167 5779 15173
rect 1670 15136 1676 15148
rect 1631 15108 1676 15136
rect 1670 15096 1676 15108
rect 1728 15096 1734 15148
rect 2682 15096 2688 15148
rect 2740 15096 2746 15148
rect 3418 15136 3424 15148
rect 3379 15108 3424 15136
rect 3418 15096 3424 15108
rect 3476 15096 3482 15148
rect 5000 15136 5028 15167
rect 5626 15136 5632 15148
rect 5000 15108 5632 15136
rect 5626 15096 5632 15108
rect 5684 15096 5690 15148
rect 5736 15136 5764 15167
rect 5902 15164 5908 15216
rect 5960 15204 5966 15216
rect 7561 15207 7619 15213
rect 7561 15204 7573 15207
rect 5960 15176 7573 15204
rect 5960 15164 5966 15176
rect 7561 15173 7573 15176
rect 7607 15173 7619 15207
rect 7561 15167 7619 15173
rect 5810 15136 5816 15148
rect 5723 15108 5816 15136
rect 5810 15096 5816 15108
rect 5868 15136 5874 15148
rect 5868 15108 7696 15136
rect 5868 15096 5874 15108
rect 7668 15080 7696 15108
rect 7650 15068 7656 15080
rect 7611 15040 7656 15068
rect 7650 15028 7656 15040
rect 7708 15028 7714 15080
rect 1104 14978 8832 15000
rect 1104 14926 3579 14978
rect 3631 14926 3643 14978
rect 3695 14926 3707 14978
rect 3759 14926 3771 14978
rect 3823 14926 6176 14978
rect 6228 14926 6240 14978
rect 6292 14926 6304 14978
rect 6356 14926 6368 14978
rect 6420 14926 8832 14978
rect 1104 14904 8832 14926
rect 4522 14864 4528 14876
rect 4356 14836 4528 14864
rect 4356 14805 4384 14836
rect 4522 14824 4528 14836
rect 4580 14864 4586 14876
rect 5166 14864 5172 14876
rect 4580 14836 5172 14864
rect 4580 14824 4586 14836
rect 5166 14824 5172 14836
rect 5224 14824 5230 14876
rect 4341 14799 4399 14805
rect 4341 14765 4353 14799
rect 4387 14765 4399 14799
rect 4341 14759 4399 14765
rect 1762 14688 1768 14740
rect 1820 14728 1826 14740
rect 2133 14731 2191 14737
rect 2133 14728 2145 14731
rect 1820 14700 2145 14728
rect 1820 14688 1826 14700
rect 2133 14697 2145 14700
rect 2179 14697 2191 14731
rect 2133 14691 2191 14697
rect 2866 14688 2872 14740
rect 2924 14728 2930 14740
rect 4065 14731 4123 14737
rect 4065 14728 4077 14731
rect 2924 14700 4077 14728
rect 2924 14688 2930 14700
rect 4065 14697 4077 14700
rect 4111 14697 4123 14731
rect 7006 14728 7012 14740
rect 4065 14691 4123 14697
rect 5460 14660 5488 14714
rect 6967 14700 7012 14728
rect 7006 14688 7012 14700
rect 7064 14688 7070 14740
rect 7374 14728 7380 14740
rect 7335 14700 7380 14728
rect 7374 14688 7380 14700
rect 7432 14688 7438 14740
rect 7650 14728 7656 14740
rect 7611 14700 7656 14728
rect 7650 14688 7656 14700
rect 7708 14688 7714 14740
rect 4172 14632 5488 14660
rect 6089 14663 6147 14669
rect 3142 14552 3148 14604
rect 3200 14592 3206 14604
rect 4172 14592 4200 14632
rect 6089 14629 6101 14663
rect 6135 14629 6147 14663
rect 6089 14623 6147 14629
rect 3200 14564 4200 14592
rect 3200 14552 3206 14564
rect 5442 14552 5448 14604
rect 5500 14592 5506 14604
rect 6104 14592 6132 14623
rect 5500 14564 6132 14592
rect 5500 14552 5506 14564
rect 2130 14484 2136 14536
rect 2188 14524 2194 14536
rect 2317 14527 2375 14533
rect 2317 14524 2329 14527
rect 2188 14496 2329 14524
rect 2188 14484 2194 14496
rect 2317 14493 2329 14496
rect 2363 14493 2375 14527
rect 2317 14487 2375 14493
rect 1104 14434 8832 14456
rect 1104 14382 2280 14434
rect 2332 14382 2344 14434
rect 2396 14382 2408 14434
rect 2460 14382 2472 14434
rect 2524 14382 4878 14434
rect 4930 14382 4942 14434
rect 4994 14382 5006 14434
rect 5058 14382 5070 14434
rect 5122 14382 7475 14434
rect 7527 14382 7539 14434
rect 7591 14382 7603 14434
rect 7655 14382 7667 14434
rect 7719 14382 8832 14434
rect 1104 14360 8832 14382
rect 5626 14280 5632 14332
rect 5684 14320 5690 14332
rect 6917 14323 6975 14329
rect 6917 14320 6929 14323
rect 5684 14292 6929 14320
rect 5684 14280 5690 14292
rect 6917 14289 6929 14292
rect 6963 14289 6975 14323
rect 6917 14283 6975 14289
rect 5902 14252 5908 14264
rect 5092 14224 5908 14252
rect 3050 14144 3056 14196
rect 3108 14184 3114 14196
rect 3421 14187 3479 14193
rect 3421 14184 3433 14187
rect 3108 14156 3433 14184
rect 3108 14144 3114 14156
rect 3421 14153 3433 14156
rect 3467 14153 3479 14187
rect 3421 14147 3479 14153
rect 1394 14116 1400 14128
rect 1307 14088 1400 14116
rect 1394 14076 1400 14088
rect 1452 14076 1458 14128
rect 3234 14076 3240 14128
rect 3292 14116 3298 14128
rect 4433 14119 4491 14125
rect 4433 14116 4445 14119
rect 3292 14088 4445 14116
rect 3292 14076 3298 14088
rect 4433 14085 4445 14088
rect 4479 14085 4491 14119
rect 4433 14079 4491 14085
rect 4985 14119 5043 14125
rect 4985 14085 4997 14119
rect 5031 14116 5043 14119
rect 5092 14116 5120 14224
rect 5902 14212 5908 14224
rect 5960 14252 5966 14264
rect 6730 14252 6736 14264
rect 5960 14224 6736 14252
rect 5960 14212 5966 14224
rect 6730 14212 6736 14224
rect 6788 14212 6794 14264
rect 5810 14184 5816 14196
rect 5771 14156 5816 14184
rect 5810 14144 5816 14156
rect 5868 14144 5874 14196
rect 6638 14144 6644 14196
rect 6696 14184 6702 14196
rect 6696 14156 7420 14184
rect 6696 14144 6702 14156
rect 5031 14088 5120 14116
rect 5169 14119 5227 14125
rect 5031 14085 5043 14088
rect 4985 14079 5043 14085
rect 5169 14085 5181 14119
rect 5215 14116 5227 14119
rect 5353 14119 5411 14125
rect 5215 14088 5304 14116
rect 5215 14085 5227 14088
rect 5169 14079 5227 14085
rect 1412 13980 1440 14076
rect 1670 14048 1676 14060
rect 1631 14020 1676 14048
rect 1670 14008 1676 14020
rect 1728 14008 1734 14060
rect 2130 14008 2136 14060
rect 2188 14008 2194 14060
rect 3050 13980 3056 13992
rect 1412 13952 3056 13980
rect 3050 13940 3056 13952
rect 3108 13940 3114 13992
rect 5276 13980 5304 14088
rect 5353 14085 5365 14119
rect 5399 14085 5411 14119
rect 5718 14116 5724 14128
rect 5679 14088 5724 14116
rect 5353 14079 5411 14085
rect 5368 14048 5396 14079
rect 5718 14076 5724 14088
rect 5776 14076 5782 14128
rect 7098 14116 7104 14128
rect 7059 14088 7104 14116
rect 7098 14076 7104 14088
rect 7156 14076 7162 14128
rect 7392 14125 7420 14156
rect 7377 14119 7435 14125
rect 7377 14085 7389 14119
rect 7423 14085 7435 14119
rect 7377 14079 7435 14085
rect 5994 14048 6000 14060
rect 5368 14020 6000 14048
rect 5994 14008 6000 14020
rect 6052 14008 6058 14060
rect 6822 13980 6828 13992
rect 5276 13952 6828 13980
rect 6822 13940 6828 13952
rect 6880 13940 6886 13992
rect 1104 13890 8832 13912
rect 1104 13838 3579 13890
rect 3631 13838 3643 13890
rect 3695 13838 3707 13890
rect 3759 13838 3771 13890
rect 3823 13838 6176 13890
rect 6228 13838 6240 13890
rect 6292 13838 6304 13890
rect 6356 13838 6368 13890
rect 6420 13838 8832 13890
rect 1104 13816 8832 13838
rect 5534 13736 5540 13788
rect 5592 13776 5598 13788
rect 7469 13779 7527 13785
rect 7469 13776 7481 13779
rect 5592 13748 7481 13776
rect 5592 13736 5598 13748
rect 7469 13745 7481 13748
rect 7515 13745 7527 13779
rect 7469 13739 7527 13745
rect 4522 13708 4528 13720
rect 4483 13680 4528 13708
rect 4522 13668 4528 13680
rect 4580 13668 4586 13720
rect 5258 13668 5264 13720
rect 5316 13668 5322 13720
rect 3237 13643 3295 13649
rect 3237 13609 3249 13643
rect 3283 13640 3295 13643
rect 3970 13640 3976 13652
rect 3283 13612 3976 13640
rect 3283 13609 3295 13612
rect 3237 13603 3295 13609
rect 3970 13600 3976 13612
rect 4028 13600 4034 13652
rect 7190 13640 7196 13652
rect 7151 13612 7196 13640
rect 7190 13600 7196 13612
rect 7248 13600 7254 13652
rect 7377 13643 7435 13649
rect 7377 13609 7389 13643
rect 7423 13640 7435 13643
rect 7834 13640 7840 13652
rect 7423 13612 7840 13640
rect 7423 13609 7435 13612
rect 7377 13603 7435 13609
rect 7834 13600 7840 13612
rect 7892 13600 7898 13652
rect 3050 13532 3056 13584
rect 3108 13572 3114 13584
rect 3878 13572 3884 13584
rect 3108 13544 3884 13572
rect 3108 13532 3114 13544
rect 3878 13532 3884 13544
rect 3936 13572 3942 13584
rect 4249 13575 4307 13581
rect 4249 13572 4261 13575
rect 3936 13544 4261 13572
rect 3936 13532 3942 13544
rect 4249 13541 4261 13544
rect 4295 13541 4307 13575
rect 4249 13535 4307 13541
rect 6273 13575 6331 13581
rect 6273 13541 6285 13575
rect 6319 13541 6331 13575
rect 6273 13535 6331 13541
rect 5626 13464 5632 13516
rect 5684 13504 5690 13516
rect 6288 13504 6316 13535
rect 5684 13476 6316 13504
rect 5684 13464 5690 13476
rect 2866 13396 2872 13448
rect 2924 13436 2930 13448
rect 3053 13439 3111 13445
rect 3053 13436 3065 13439
rect 2924 13408 3065 13436
rect 2924 13396 2930 13408
rect 3053 13405 3065 13408
rect 3099 13405 3111 13439
rect 3053 13399 3111 13405
rect 4062 13396 4068 13448
rect 4120 13436 4126 13448
rect 7006 13436 7012 13448
rect 4120 13408 7012 13436
rect 4120 13396 4126 13408
rect 7006 13396 7012 13408
rect 7064 13436 7070 13448
rect 7282 13436 7288 13448
rect 7064 13408 7288 13436
rect 7064 13396 7070 13408
rect 7282 13396 7288 13408
rect 7340 13396 7346 13448
rect 1104 13346 8832 13368
rect 1104 13294 2280 13346
rect 2332 13294 2344 13346
rect 2396 13294 2408 13346
rect 2460 13294 2472 13346
rect 2524 13294 4878 13346
rect 4930 13294 4942 13346
rect 4994 13294 5006 13346
rect 5058 13294 5070 13346
rect 5122 13294 7475 13346
rect 7527 13294 7539 13346
rect 7591 13294 7603 13346
rect 7655 13294 7667 13346
rect 7719 13294 8832 13346
rect 1104 13272 8832 13294
rect 3418 13232 3424 13244
rect 2056 13204 3424 13232
rect 1762 13056 1768 13108
rect 1820 13096 1826 13108
rect 2056 13096 2084 13204
rect 3418 13192 3424 13204
rect 3476 13192 3482 13244
rect 7190 13192 7196 13244
rect 7248 13232 7254 13244
rect 7285 13235 7343 13241
rect 7285 13232 7297 13235
rect 7248 13204 7297 13232
rect 7248 13192 7254 13204
rect 7285 13201 7297 13204
rect 7331 13201 7343 13235
rect 7285 13195 7343 13201
rect 2225 13099 2283 13105
rect 2225 13096 2237 13099
rect 1820 13068 2237 13096
rect 1820 13056 1826 13068
rect 2225 13065 2237 13068
rect 2271 13065 2283 13099
rect 2225 13059 2283 13065
rect 3234 13056 3240 13108
rect 3292 13096 3298 13108
rect 3973 13099 4031 13105
rect 3973 13096 3985 13099
rect 3292 13068 3985 13096
rect 3292 13056 3298 13068
rect 3973 13065 3985 13068
rect 4019 13065 4031 13099
rect 3973 13059 4031 13065
rect 5626 13056 5632 13108
rect 5684 13096 5690 13108
rect 5684 13068 7144 13096
rect 5684 13056 5690 13068
rect 1949 13031 2007 13037
rect 1949 12997 1961 13031
rect 1995 12997 2007 13031
rect 1949 12991 2007 12997
rect 1964 12892 1992 12991
rect 4706 12988 4712 13040
rect 4764 13028 4770 13040
rect 4801 13031 4859 13037
rect 4801 13028 4813 13031
rect 4764 13000 4813 13028
rect 4764 12988 4770 13000
rect 4801 12997 4813 13000
rect 4847 12997 4859 13031
rect 4801 12991 4859 12997
rect 6822 12988 6828 13040
rect 6880 13028 6886 13040
rect 7116 13037 7144 13068
rect 6917 13031 6975 13037
rect 6917 13028 6929 13031
rect 6880 13000 6929 13028
rect 6880 12988 6886 13000
rect 6917 12997 6929 13000
rect 6963 12997 6975 13031
rect 6917 12991 6975 12997
rect 7101 13031 7159 13037
rect 7101 12997 7113 13031
rect 7147 12997 7159 13031
rect 7101 12991 7159 12997
rect 2958 12920 2964 12972
rect 3016 12920 3022 12972
rect 7006 12960 7012 12972
rect 6967 12932 7012 12960
rect 7006 12920 7012 12932
rect 7064 12920 7070 12972
rect 3050 12892 3056 12904
rect 1964 12864 3056 12892
rect 3050 12852 3056 12864
rect 3108 12852 3114 12904
rect 4985 12895 5043 12901
rect 4985 12861 4997 12895
rect 5031 12892 5043 12895
rect 5166 12892 5172 12904
rect 5031 12864 5172 12892
rect 5031 12861 5043 12864
rect 4985 12855 5043 12861
rect 5166 12852 5172 12864
rect 5224 12852 5230 12904
rect 1104 12802 8832 12824
rect 1104 12750 3579 12802
rect 3631 12750 3643 12802
rect 3695 12750 3707 12802
rect 3759 12750 3771 12802
rect 3823 12750 6176 12802
rect 6228 12750 6240 12802
rect 6292 12750 6304 12802
rect 6356 12750 6368 12802
rect 6420 12750 8832 12802
rect 1104 12728 8832 12750
rect 2958 12648 2964 12700
rect 3016 12688 3022 12700
rect 3053 12691 3111 12697
rect 3053 12688 3065 12691
rect 3016 12660 3065 12688
rect 3016 12648 3022 12660
rect 3053 12657 3065 12660
rect 3099 12657 3111 12691
rect 3053 12651 3111 12657
rect 4249 12691 4307 12697
rect 4249 12657 4261 12691
rect 4295 12688 4307 12691
rect 4706 12688 4712 12700
rect 4295 12660 4712 12688
rect 4295 12657 4307 12660
rect 4249 12651 4307 12657
rect 4264 12620 4292 12651
rect 4706 12648 4712 12660
rect 4764 12648 4770 12700
rect 2884 12592 4292 12620
rect 2884 12561 2912 12592
rect 6546 12580 6552 12632
rect 6604 12580 6610 12632
rect 2869 12555 2927 12561
rect 2869 12521 2881 12555
rect 2915 12521 2927 12555
rect 2869 12515 2927 12521
rect 2958 12512 2964 12564
rect 3016 12552 3022 12564
rect 4065 12555 4123 12561
rect 4065 12552 4077 12555
rect 3016 12524 4077 12552
rect 3016 12512 3022 12524
rect 4065 12521 4077 12524
rect 4111 12521 4123 12555
rect 4065 12515 4123 12521
rect 3878 12444 3884 12496
rect 3936 12484 3942 12496
rect 5169 12487 5227 12493
rect 5169 12484 5181 12487
rect 3936 12456 5181 12484
rect 3936 12444 3942 12456
rect 5169 12453 5181 12456
rect 5215 12453 5227 12487
rect 5534 12484 5540 12496
rect 5495 12456 5540 12484
rect 5169 12447 5227 12453
rect 5534 12444 5540 12456
rect 5592 12444 5598 12496
rect 5994 12444 6000 12496
rect 6052 12484 6058 12496
rect 6917 12487 6975 12493
rect 6917 12484 6929 12487
rect 6052 12456 6929 12484
rect 6052 12444 6058 12456
rect 6917 12453 6929 12456
rect 6963 12453 6975 12487
rect 6917 12447 6975 12453
rect 1104 12258 8832 12280
rect 1104 12206 2280 12258
rect 2332 12206 2344 12258
rect 2396 12206 2408 12258
rect 2460 12206 2472 12258
rect 2524 12206 4878 12258
rect 4930 12206 4942 12258
rect 4994 12206 5006 12258
rect 5058 12206 5070 12258
rect 5122 12206 7475 12258
rect 7527 12206 7539 12258
rect 7591 12206 7603 12258
rect 7655 12206 7667 12258
rect 7719 12206 8832 12258
rect 1104 12184 8832 12206
rect 2961 12147 3019 12153
rect 2961 12113 2973 12147
rect 3007 12144 3019 12147
rect 3142 12144 3148 12156
rect 3007 12116 3148 12144
rect 3007 12113 3019 12116
rect 2961 12107 3019 12113
rect 3142 12104 3148 12116
rect 3200 12104 3206 12156
rect 6917 12147 6975 12153
rect 6917 12113 6929 12147
rect 6963 12144 6975 12147
rect 7006 12144 7012 12156
rect 6963 12116 7012 12144
rect 6963 12113 6975 12116
rect 6917 12107 6975 12113
rect 7006 12104 7012 12116
rect 7064 12104 7070 12156
rect 3878 12008 3884 12020
rect 3839 11980 3884 12008
rect 3878 11968 3884 11980
rect 3936 11968 3942 12020
rect 4157 12011 4215 12017
rect 4157 11977 4169 12011
rect 4203 12008 4215 12011
rect 5442 12008 5448 12020
rect 4203 11980 5448 12008
rect 4203 11977 4215 11980
rect 4157 11971 4215 11977
rect 5442 11968 5448 11980
rect 5500 11968 5506 12020
rect 2777 11943 2835 11949
rect 2777 11909 2789 11943
rect 2823 11940 2835 11943
rect 2958 11940 2964 11952
rect 2823 11912 2964 11940
rect 2823 11909 2835 11912
rect 2777 11903 2835 11909
rect 2958 11900 2964 11912
rect 3016 11900 3022 11952
rect 5902 11940 5908 11952
rect 5815 11912 5908 11940
rect 5902 11900 5908 11912
rect 5960 11940 5966 11952
rect 6825 11943 6883 11949
rect 6825 11940 6837 11943
rect 5960 11912 6837 11940
rect 5960 11900 5966 11912
rect 6825 11909 6837 11912
rect 6871 11909 6883 11943
rect 6825 11903 6883 11909
rect 5166 11832 5172 11884
rect 5224 11832 5230 11884
rect 1104 11714 8832 11736
rect 1104 11662 3579 11714
rect 3631 11662 3643 11714
rect 3695 11662 3707 11714
rect 3759 11662 3771 11714
rect 3823 11662 6176 11714
rect 6228 11662 6240 11714
rect 6292 11662 6304 11714
rect 6356 11662 6368 11714
rect 6420 11662 8832 11714
rect 1104 11640 8832 11662
rect 2317 11603 2375 11609
rect 2317 11569 2329 11603
rect 2363 11600 2375 11603
rect 2682 11600 2688 11612
rect 2363 11572 2688 11600
rect 2363 11569 2375 11572
rect 2317 11563 2375 11569
rect 2682 11560 2688 11572
rect 2740 11560 2746 11612
rect 5258 11600 5264 11612
rect 5219 11572 5264 11600
rect 5258 11560 5264 11572
rect 5316 11560 5322 11612
rect 6365 11603 6423 11609
rect 6365 11569 6377 11603
rect 6411 11600 6423 11603
rect 6546 11600 6552 11612
rect 6411 11572 6552 11600
rect 6411 11569 6423 11572
rect 6365 11563 6423 11569
rect 6546 11560 6552 11572
rect 6604 11560 6610 11612
rect 2038 11424 2044 11476
rect 2096 11464 2102 11476
rect 2133 11467 2191 11473
rect 2133 11464 2145 11467
rect 2096 11436 2145 11464
rect 2096 11424 2102 11436
rect 2133 11433 2145 11436
rect 2179 11433 2191 11467
rect 2133 11427 2191 11433
rect 4706 11424 4712 11476
rect 4764 11464 4770 11476
rect 5077 11467 5135 11473
rect 5077 11464 5089 11467
rect 4764 11436 5089 11464
rect 4764 11424 4770 11436
rect 5077 11433 5089 11436
rect 5123 11464 5135 11467
rect 6181 11467 6239 11473
rect 6181 11464 6193 11467
rect 5123 11436 6193 11464
rect 5123 11433 5135 11436
rect 5077 11427 5135 11433
rect 6181 11433 6193 11436
rect 6227 11433 6239 11467
rect 6181 11427 6239 11433
rect 1104 11170 8832 11192
rect 1104 11118 2280 11170
rect 2332 11118 2344 11170
rect 2396 11118 2408 11170
rect 2460 11118 2472 11170
rect 2524 11118 4878 11170
rect 4930 11118 4942 11170
rect 4994 11118 5006 11170
rect 5058 11118 5070 11170
rect 5122 11118 7475 11170
rect 7527 11118 7539 11170
rect 7591 11118 7603 11170
rect 7655 11118 7667 11170
rect 7719 11118 8832 11170
rect 1104 11096 8832 11118
rect 2866 11056 2872 11068
rect 1412 11028 2872 11056
rect 1412 10929 1440 11028
rect 2866 11016 2872 11028
rect 2924 11016 2930 11068
rect 1397 10923 1455 10929
rect 1397 10889 1409 10923
rect 1443 10889 1455 10923
rect 1397 10883 1455 10889
rect 1670 10880 1676 10932
rect 1728 10920 1734 10932
rect 3421 10923 3479 10929
rect 3421 10920 3433 10923
rect 1728 10892 3433 10920
rect 1728 10880 1734 10892
rect 3421 10889 3433 10892
rect 3467 10889 3479 10923
rect 3421 10883 3479 10889
rect 1670 10784 1676 10796
rect 1631 10756 1676 10784
rect 1670 10744 1676 10756
rect 1728 10744 1734 10796
rect 1946 10744 1952 10796
rect 2004 10784 2010 10796
rect 4249 10787 4307 10793
rect 2004 10756 2162 10784
rect 2004 10744 2010 10756
rect 4249 10753 4261 10787
rect 4295 10784 4307 10787
rect 6638 10784 6644 10796
rect 4295 10756 6644 10784
rect 4295 10753 4307 10756
rect 4249 10747 4307 10753
rect 6638 10744 6644 10756
rect 6696 10744 6702 10796
rect 3970 10676 3976 10728
rect 4028 10716 4034 10728
rect 5537 10719 5595 10725
rect 5537 10716 5549 10719
rect 4028 10688 5549 10716
rect 4028 10676 4034 10688
rect 5537 10685 5549 10688
rect 5583 10685 5595 10719
rect 5537 10679 5595 10685
rect 1104 10626 8832 10648
rect 1104 10574 3579 10626
rect 3631 10574 3643 10626
rect 3695 10574 3707 10626
rect 3759 10574 3771 10626
rect 3823 10574 6176 10626
rect 6228 10574 6240 10626
rect 6292 10574 6304 10626
rect 6356 10574 6368 10626
rect 6420 10574 8832 10626
rect 1104 10552 8832 10574
rect 1854 10336 1860 10388
rect 1912 10376 1918 10388
rect 2225 10379 2283 10385
rect 2225 10376 2237 10379
rect 1912 10348 2237 10376
rect 1912 10336 1918 10348
rect 2225 10345 2237 10348
rect 2271 10345 2283 10379
rect 2225 10339 2283 10345
rect 2130 10200 2136 10252
rect 2188 10240 2194 10252
rect 2409 10243 2467 10249
rect 2409 10240 2421 10243
rect 2188 10212 2421 10240
rect 2188 10200 2194 10212
rect 2409 10209 2421 10212
rect 2455 10209 2467 10243
rect 2409 10203 2467 10209
rect 1104 10082 8832 10104
rect 1104 10030 2280 10082
rect 2332 10030 2344 10082
rect 2396 10030 2408 10082
rect 2460 10030 2472 10082
rect 2524 10030 4878 10082
rect 4930 10030 4942 10082
rect 4994 10030 5006 10082
rect 5058 10030 5070 10082
rect 5122 10030 7475 10082
rect 7527 10030 7539 10082
rect 7591 10030 7603 10082
rect 7655 10030 7667 10082
rect 7719 10030 8832 10082
rect 1104 10008 8832 10030
rect 1397 9835 1455 9841
rect 1397 9801 1409 9835
rect 1443 9832 1455 9835
rect 3418 9832 3424 9844
rect 1443 9804 3188 9832
rect 3379 9804 3424 9832
rect 1443 9801 1455 9804
rect 1397 9795 1455 9801
rect 3160 9764 3188 9804
rect 3418 9792 3424 9804
rect 3476 9792 3482 9844
rect 3878 9764 3884 9776
rect 3160 9736 3884 9764
rect 3878 9724 3884 9736
rect 3936 9724 3942 9776
rect 6822 9724 6828 9776
rect 6880 9764 6886 9776
rect 7193 9767 7251 9773
rect 7193 9764 7205 9767
rect 6880 9736 7205 9764
rect 6880 9724 6886 9736
rect 7193 9733 7205 9736
rect 7239 9733 7251 9767
rect 7193 9727 7251 9733
rect 7282 9724 7288 9776
rect 7340 9764 7346 9776
rect 7340 9736 7385 9764
rect 7340 9724 7346 9736
rect 1670 9696 1676 9708
rect 1631 9668 1676 9696
rect 1670 9656 1676 9668
rect 1728 9656 1734 9708
rect 2130 9656 2136 9708
rect 2188 9656 2194 9708
rect 7745 9699 7803 9705
rect 7745 9665 7757 9699
rect 7791 9696 7803 9699
rect 8202 9696 8208 9708
rect 7791 9668 8208 9696
rect 7791 9665 7803 9668
rect 7745 9659 7803 9665
rect 8202 9656 8208 9668
rect 8260 9656 8266 9708
rect 1104 9538 8832 9560
rect 1104 9486 3579 9538
rect 3631 9486 3643 9538
rect 3695 9486 3707 9538
rect 3759 9486 3771 9538
rect 3823 9486 6176 9538
rect 6228 9486 6240 9538
rect 6292 9486 6304 9538
rect 6356 9486 6368 9538
rect 6420 9486 8832 9538
rect 1104 9464 8832 9486
rect 1946 9424 1952 9436
rect 1907 9396 1952 9424
rect 1946 9384 1952 9396
rect 2004 9384 2010 9436
rect 7006 9356 7012 9368
rect 6486 9328 7012 9356
rect 7006 9316 7012 9328
rect 7064 9316 7070 9368
rect 1765 9291 1823 9297
rect 1765 9257 1777 9291
rect 1811 9288 1823 9291
rect 2038 9288 2044 9300
rect 1811 9260 2044 9288
rect 1811 9257 1823 9260
rect 1765 9251 1823 9257
rect 2038 9248 2044 9260
rect 2096 9288 2102 9300
rect 2682 9288 2688 9300
rect 2096 9260 2688 9288
rect 2096 9248 2102 9260
rect 2682 9248 2688 9260
rect 2740 9248 2746 9300
rect 2869 9291 2927 9297
rect 2869 9257 2881 9291
rect 2915 9288 2927 9291
rect 2958 9288 2964 9300
rect 2915 9260 2964 9288
rect 2915 9257 2927 9260
rect 2869 9251 2927 9257
rect 2958 9248 2964 9260
rect 3016 9248 3022 9300
rect 4706 9248 4712 9300
rect 4764 9288 4770 9300
rect 5445 9291 5503 9297
rect 5445 9288 5457 9291
rect 4764 9260 5457 9288
rect 4764 9248 4770 9260
rect 5445 9257 5457 9260
rect 5491 9257 5503 9291
rect 5445 9251 5503 9257
rect 3878 9180 3884 9232
rect 3936 9220 3942 9232
rect 5077 9223 5135 9229
rect 5077 9220 5089 9223
rect 3936 9192 5089 9220
rect 3936 9180 3942 9192
rect 5077 9189 5089 9192
rect 5123 9189 5135 9223
rect 6822 9220 6828 9232
rect 6783 9192 6828 9220
rect 5077 9183 5135 9189
rect 6822 9180 6828 9192
rect 6880 9180 6886 9232
rect 2682 9044 2688 9096
rect 2740 9084 2746 9096
rect 3053 9087 3111 9093
rect 3053 9084 3065 9087
rect 2740 9056 3065 9084
rect 2740 9044 2746 9056
rect 3053 9053 3065 9056
rect 3099 9053 3111 9087
rect 3053 9047 3111 9053
rect 1104 8994 8832 9016
rect 1104 8942 2280 8994
rect 2332 8942 2344 8994
rect 2396 8942 2408 8994
rect 2460 8942 2472 8994
rect 2524 8942 4878 8994
rect 4930 8942 4942 8994
rect 4994 8942 5006 8994
rect 5058 8942 5070 8994
rect 5122 8942 7475 8994
rect 7527 8942 7539 8994
rect 7591 8942 7603 8994
rect 7655 8942 7667 8994
rect 7719 8942 8832 8994
rect 1104 8920 8832 8942
rect 7006 8880 7012 8892
rect 2608 8852 4660 8880
rect 6967 8852 7012 8880
rect 1854 8772 1860 8824
rect 1912 8812 1918 8824
rect 2608 8812 2636 8852
rect 1912 8784 2636 8812
rect 1912 8772 1918 8784
rect 1670 8704 1676 8756
rect 1728 8744 1734 8756
rect 4525 8747 4583 8753
rect 4525 8744 4537 8747
rect 1728 8716 4537 8744
rect 1728 8704 1734 8716
rect 4525 8713 4537 8716
rect 4571 8713 4583 8747
rect 4632 8744 4660 8852
rect 7006 8840 7012 8852
rect 7064 8840 7070 8892
rect 4632 8716 6868 8744
rect 4525 8707 4583 8713
rect 2498 8676 2504 8688
rect 2459 8648 2504 8676
rect 2498 8636 2504 8648
rect 2556 8636 2562 8688
rect 4062 8636 4068 8688
rect 4120 8676 4126 8688
rect 6840 8685 6868 8716
rect 5353 8679 5411 8685
rect 5353 8676 5365 8679
rect 4120 8648 5365 8676
rect 4120 8636 4126 8648
rect 5353 8645 5365 8648
rect 5399 8645 5411 8679
rect 5353 8639 5411 8645
rect 6825 8679 6883 8685
rect 6825 8645 6837 8679
rect 6871 8676 6883 8679
rect 7466 8676 7472 8688
rect 6871 8648 7472 8676
rect 6871 8645 6883 8648
rect 6825 8639 6883 8645
rect 7466 8636 7472 8648
rect 7524 8636 7530 8688
rect 2777 8611 2835 8617
rect 2777 8577 2789 8611
rect 2823 8577 2835 8611
rect 2777 8571 2835 8577
rect 2792 8540 2820 8571
rect 3050 8568 3056 8620
rect 3108 8608 3114 8620
rect 3108 8580 3266 8608
rect 3108 8568 3114 8580
rect 4614 8568 4620 8620
rect 4672 8608 4678 8620
rect 4672 8580 5580 8608
rect 4672 8568 4678 8580
rect 5442 8540 5448 8552
rect 2792 8512 5448 8540
rect 5442 8500 5448 8512
rect 5500 8500 5506 8552
rect 5552 8549 5580 8580
rect 5537 8543 5595 8549
rect 5537 8509 5549 8543
rect 5583 8509 5595 8543
rect 5537 8503 5595 8509
rect 1104 8450 8832 8472
rect 1104 8398 3579 8450
rect 3631 8398 3643 8450
rect 3695 8398 3707 8450
rect 3759 8398 3771 8450
rect 3823 8398 6176 8450
rect 6228 8398 6240 8450
rect 6292 8398 6304 8450
rect 6356 8398 6368 8450
rect 6420 8398 8832 8450
rect 1104 8376 8832 8398
rect 3050 8336 3056 8348
rect 3011 8308 3056 8336
rect 3050 8296 3056 8308
rect 3108 8296 3114 8348
rect 5534 8296 5540 8348
rect 5592 8336 5598 8348
rect 7466 8336 7472 8348
rect 5592 8308 6500 8336
rect 7427 8308 7472 8336
rect 5592 8296 5598 8308
rect 3970 8268 3976 8280
rect 2792 8240 3976 8268
rect 2792 8209 2820 8240
rect 3970 8228 3976 8240
rect 4028 8228 4034 8280
rect 5718 8228 5724 8280
rect 5776 8228 5782 8280
rect 6472 8277 6500 8308
rect 7466 8296 7472 8308
rect 7524 8296 7530 8348
rect 6457 8271 6515 8277
rect 6457 8237 6469 8271
rect 6503 8237 6515 8271
rect 6457 8231 6515 8237
rect 2777 8203 2835 8209
rect 2777 8169 2789 8203
rect 2823 8169 2835 8203
rect 2777 8163 2835 8169
rect 2869 8203 2927 8209
rect 2869 8169 2881 8203
rect 2915 8169 2927 8203
rect 2869 8163 2927 8169
rect 7291 8203 7349 8209
rect 7291 8169 7303 8203
rect 7337 8169 7349 8203
rect 7291 8163 7349 8169
rect 2130 8092 2136 8144
rect 2188 8132 2194 8144
rect 2682 8132 2688 8144
rect 2188 8104 2688 8132
rect 2188 8092 2194 8104
rect 2682 8092 2688 8104
rect 2740 8132 2746 8144
rect 2884 8132 2912 8163
rect 2740 8104 2912 8132
rect 2740 8092 2746 8104
rect 4154 8092 4160 8144
rect 4212 8132 4218 8144
rect 4433 8135 4491 8141
rect 4433 8132 4445 8135
rect 4212 8104 4445 8132
rect 4212 8092 4218 8104
rect 4433 8101 4445 8104
rect 4479 8101 4491 8135
rect 4706 8132 4712 8144
rect 4667 8104 4712 8132
rect 4433 8095 4491 8101
rect 4706 8092 4712 8104
rect 4764 8092 4770 8144
rect 2498 8024 2504 8076
rect 2556 8064 2562 8076
rect 2593 8067 2651 8073
rect 2593 8064 2605 8067
rect 2556 8036 2605 8064
rect 2556 8024 2562 8036
rect 2593 8033 2605 8036
rect 2639 8064 2651 8067
rect 4172 8064 4200 8092
rect 2639 8036 4200 8064
rect 2639 8033 2651 8036
rect 2593 8027 2651 8033
rect 4430 7956 4436 8008
rect 4488 7996 4494 8008
rect 5258 7996 5264 8008
rect 4488 7968 5264 7996
rect 4488 7956 4494 7968
rect 5258 7956 5264 7968
rect 5316 7996 5322 8008
rect 7300 7996 7328 8163
rect 5316 7968 7328 7996
rect 5316 7956 5322 7968
rect 1104 7906 8832 7928
rect 1104 7854 2280 7906
rect 2332 7854 2344 7906
rect 2396 7854 2408 7906
rect 2460 7854 2472 7906
rect 2524 7854 4878 7906
rect 4930 7854 4942 7906
rect 4994 7854 5006 7906
rect 5058 7854 5070 7906
rect 5122 7854 7475 7906
rect 7527 7854 7539 7906
rect 7591 7854 7603 7906
rect 7655 7854 7667 7906
rect 7719 7854 8832 7906
rect 1104 7832 8832 7854
rect 3326 7752 3332 7804
rect 3384 7792 3390 7804
rect 5718 7792 5724 7804
rect 3384 7764 5580 7792
rect 5679 7764 5724 7792
rect 3384 7752 3390 7764
rect 4062 7724 4068 7736
rect 3344 7696 4068 7724
rect 2958 7548 2964 7600
rect 3016 7588 3022 7600
rect 3344 7597 3372 7696
rect 4062 7684 4068 7696
rect 4120 7724 4126 7736
rect 4617 7727 4675 7733
rect 4617 7724 4629 7727
rect 4120 7696 4629 7724
rect 4120 7684 4126 7696
rect 4617 7693 4629 7696
rect 4663 7693 4675 7727
rect 5552 7724 5580 7764
rect 5718 7752 5724 7764
rect 5776 7752 5782 7804
rect 5902 7724 5908 7736
rect 5552 7696 5908 7724
rect 4617 7687 4675 7693
rect 5902 7684 5908 7696
rect 5960 7684 5966 7736
rect 3329 7591 3387 7597
rect 3329 7588 3341 7591
rect 3016 7560 3341 7588
rect 3016 7548 3022 7560
rect 3329 7557 3341 7560
rect 3375 7557 3387 7591
rect 4430 7588 4436 7600
rect 4391 7560 4436 7588
rect 3329 7551 3387 7557
rect 4430 7548 4436 7560
rect 4488 7548 4494 7600
rect 5537 7591 5595 7597
rect 5537 7557 5549 7591
rect 5583 7557 5595 7591
rect 5537 7551 5595 7557
rect 5552 7520 5580 7551
rect 3528 7492 5580 7520
rect 3142 7412 3148 7464
rect 3200 7452 3206 7464
rect 3528 7461 3556 7492
rect 3513 7455 3571 7461
rect 3513 7452 3525 7455
rect 3200 7424 3525 7452
rect 3200 7412 3206 7424
rect 3513 7421 3525 7424
rect 3559 7421 3571 7455
rect 3513 7415 3571 7421
rect 4062 7412 4068 7464
rect 4120 7452 4126 7464
rect 5626 7452 5632 7464
rect 4120 7424 5632 7452
rect 4120 7412 4126 7424
rect 5626 7412 5632 7424
rect 5684 7412 5690 7464
rect 1104 7362 8832 7384
rect 1104 7310 3579 7362
rect 3631 7310 3643 7362
rect 3695 7310 3707 7362
rect 3759 7310 3771 7362
rect 3823 7310 6176 7362
rect 6228 7310 6240 7362
rect 6292 7310 6304 7362
rect 6356 7310 6368 7362
rect 6420 7310 8832 7362
rect 1104 7288 8832 7310
rect 4706 7208 4712 7260
rect 4764 7248 4770 7260
rect 4764 7220 6408 7248
rect 4764 7208 4770 7220
rect 6380 7189 6408 7220
rect 6365 7183 6423 7189
rect 6365 7149 6377 7183
rect 6411 7149 6423 7183
rect 6365 7143 6423 7149
rect 5718 7072 5724 7124
rect 5776 7072 5782 7124
rect 4154 7004 4160 7056
rect 4212 7044 4218 7056
rect 4341 7047 4399 7053
rect 4341 7044 4353 7047
rect 4212 7016 4353 7044
rect 4212 7004 4218 7016
rect 4341 7013 4353 7016
rect 4387 7013 4399 7047
rect 4341 7007 4399 7013
rect 4617 7047 4675 7053
rect 4617 7013 4629 7047
rect 4663 7044 4675 7047
rect 5626 7044 5632 7056
rect 4663 7016 5632 7044
rect 4663 7013 4675 7016
rect 4617 7007 4675 7013
rect 5626 7004 5632 7016
rect 5684 7004 5690 7056
rect 1104 6818 8832 6840
rect 1104 6766 2280 6818
rect 2332 6766 2344 6818
rect 2396 6766 2408 6818
rect 2460 6766 2472 6818
rect 2524 6766 4878 6818
rect 4930 6766 4942 6818
rect 4994 6766 5006 6818
rect 5058 6766 5070 6818
rect 5122 6766 7475 6818
rect 7527 6766 7539 6818
rect 7591 6766 7603 6818
rect 7655 6766 7667 6818
rect 7719 6766 8832 6818
rect 1104 6744 8832 6766
rect 5537 6707 5595 6713
rect 5537 6673 5549 6707
rect 5583 6704 5595 6707
rect 5718 6704 5724 6716
rect 5583 6676 5724 6704
rect 5583 6673 5595 6676
rect 5537 6667 5595 6673
rect 5718 6664 5724 6676
rect 5776 6664 5782 6716
rect 3142 6528 3148 6580
rect 3200 6568 3206 6580
rect 3200 6540 5396 6568
rect 3200 6528 3206 6540
rect 1394 6500 1400 6512
rect 1355 6472 1400 6500
rect 1394 6460 1400 6472
rect 1452 6460 1458 6512
rect 4249 6503 4307 6509
rect 4249 6469 4261 6503
rect 4295 6500 4307 6503
rect 4614 6500 4620 6512
rect 4295 6472 4620 6500
rect 4295 6469 4307 6472
rect 4249 6463 4307 6469
rect 4614 6460 4620 6472
rect 4672 6460 4678 6512
rect 5368 6509 5396 6540
rect 5353 6503 5411 6509
rect 5353 6469 5365 6503
rect 5399 6469 5411 6503
rect 5353 6463 5411 6469
rect 1670 6432 1676 6444
rect 1631 6404 1676 6432
rect 1670 6392 1676 6404
rect 1728 6392 1734 6444
rect 2682 6392 2688 6444
rect 2740 6392 2746 6444
rect 3418 6432 3424 6444
rect 3379 6404 3424 6432
rect 3418 6392 3424 6404
rect 3476 6392 3482 6444
rect 4430 6364 4436 6376
rect 4391 6336 4436 6364
rect 4430 6324 4436 6336
rect 4488 6324 4494 6376
rect 1104 6274 8832 6296
rect 1104 6222 3579 6274
rect 3631 6222 3643 6274
rect 3695 6222 3707 6274
rect 3759 6222 3771 6274
rect 3823 6222 6176 6274
rect 6228 6222 6240 6274
rect 6292 6222 6304 6274
rect 6356 6222 6368 6274
rect 6420 6222 8832 6274
rect 1104 6200 8832 6222
rect 1946 5984 1952 6036
rect 2004 6024 2010 6036
rect 2130 6024 2136 6036
rect 2004 5996 2136 6024
rect 2004 5984 2010 5996
rect 2130 5984 2136 5996
rect 2188 5984 2194 6036
rect 1394 5916 1400 5968
rect 1452 5956 1458 5968
rect 4154 5956 4160 5968
rect 1452 5928 4160 5956
rect 1452 5916 1458 5928
rect 4154 5916 4160 5928
rect 4212 5916 4218 5968
rect 2130 5780 2136 5832
rect 2188 5820 2194 5832
rect 2317 5823 2375 5829
rect 2317 5820 2329 5823
rect 2188 5792 2329 5820
rect 2188 5780 2194 5792
rect 2317 5789 2329 5792
rect 2363 5789 2375 5823
rect 2317 5783 2375 5789
rect 1104 5730 8832 5752
rect 1104 5678 2280 5730
rect 2332 5678 2344 5730
rect 2396 5678 2408 5730
rect 2460 5678 2472 5730
rect 2524 5678 4878 5730
rect 4930 5678 4942 5730
rect 4994 5678 5006 5730
rect 5058 5678 5070 5730
rect 5122 5678 7475 5730
rect 7527 5678 7539 5730
rect 7591 5678 7603 5730
rect 7655 5678 7667 5730
rect 7719 5678 8832 5730
rect 1104 5656 8832 5678
rect 1394 5480 1400 5492
rect 1355 5452 1400 5480
rect 1394 5440 1400 5452
rect 1452 5440 1458 5492
rect 1673 5483 1731 5489
rect 1673 5449 1685 5483
rect 1719 5480 1731 5483
rect 1762 5480 1768 5492
rect 1719 5452 1768 5480
rect 1719 5449 1731 5452
rect 1673 5443 1731 5449
rect 1762 5440 1768 5452
rect 1820 5440 1826 5492
rect 2130 5304 2136 5356
rect 2188 5304 2194 5356
rect 3421 5347 3479 5353
rect 3421 5313 3433 5347
rect 3467 5313 3479 5347
rect 3421 5307 3479 5313
rect 1670 5236 1676 5288
rect 1728 5276 1734 5288
rect 3436 5276 3464 5307
rect 1728 5248 3464 5276
rect 1728 5236 1734 5248
rect 1104 5186 8832 5208
rect 1104 5134 3579 5186
rect 3631 5134 3643 5186
rect 3695 5134 3707 5186
rect 3759 5134 3771 5186
rect 3823 5134 6176 5186
rect 6228 5134 6240 5186
rect 6292 5134 6304 5186
rect 6356 5134 6368 5186
rect 6420 5134 8832 5186
rect 1104 5112 8832 5134
rect 2409 5075 2467 5081
rect 2409 5041 2421 5075
rect 2455 5072 2467 5075
rect 2682 5072 2688 5084
rect 2455 5044 2688 5072
rect 2455 5041 2467 5044
rect 2409 5035 2467 5041
rect 2682 5032 2688 5044
rect 2740 5032 2746 5084
rect 3326 5032 3332 5084
rect 3384 5072 3390 5084
rect 6546 5072 6552 5084
rect 3384 5044 6552 5072
rect 3384 5032 3390 5044
rect 6546 5032 6552 5044
rect 6604 5032 6610 5084
rect 3142 4964 3148 5016
rect 3200 5004 3206 5016
rect 3418 5004 3424 5016
rect 3200 4976 3424 5004
rect 3200 4964 3206 4976
rect 3418 4964 3424 4976
rect 3476 5004 3482 5016
rect 4341 5007 4399 5013
rect 4341 5004 4353 5007
rect 3476 4976 4353 5004
rect 3476 4964 3482 4976
rect 4341 4973 4353 4976
rect 4387 4973 4399 5007
rect 4341 4967 4399 4973
rect 4430 4964 4436 5016
rect 4488 5004 4494 5016
rect 4488 4976 4830 5004
rect 4488 4964 4494 4976
rect 1946 4896 1952 4948
rect 2004 4936 2010 4948
rect 2225 4939 2283 4945
rect 2225 4936 2237 4939
rect 2004 4908 2237 4936
rect 2004 4896 2010 4908
rect 2225 4905 2237 4908
rect 2271 4905 2283 4939
rect 4062 4936 4068 4948
rect 4023 4908 4068 4936
rect 2225 4899 2283 4905
rect 4062 4896 4068 4908
rect 4120 4896 4126 4948
rect 4338 4828 4344 4880
rect 4396 4868 4402 4880
rect 5350 4868 5356 4880
rect 4396 4840 5356 4868
rect 4396 4828 4402 4840
rect 5350 4828 5356 4840
rect 5408 4868 5414 4880
rect 6089 4871 6147 4877
rect 6089 4868 6101 4871
rect 5408 4840 6101 4868
rect 5408 4828 5414 4840
rect 6089 4837 6101 4840
rect 6135 4837 6147 4871
rect 6089 4831 6147 4837
rect 1104 4642 8832 4664
rect 1104 4590 2280 4642
rect 2332 4590 2344 4642
rect 2396 4590 2408 4642
rect 2460 4590 2472 4642
rect 2524 4590 4878 4642
rect 4930 4590 4942 4642
rect 4994 4590 5006 4642
rect 5058 4590 5070 4642
rect 5122 4590 7475 4642
rect 7527 4590 7539 4642
rect 7591 4590 7603 4642
rect 7655 4590 7667 4642
rect 7719 4590 8832 4642
rect 1104 4568 8832 4590
rect 2866 4352 2872 4404
rect 2924 4392 2930 4404
rect 4617 4395 4675 4401
rect 4617 4392 4629 4395
rect 2924 4364 4629 4392
rect 2924 4352 2930 4364
rect 4617 4361 4629 4364
rect 4663 4361 4675 4395
rect 4617 4355 4675 4361
rect 2593 4327 2651 4333
rect 2593 4293 2605 4327
rect 2639 4293 2651 4327
rect 2593 4287 2651 4293
rect 2608 4256 2636 4287
rect 2774 4256 2780 4268
rect 2608 4228 2780 4256
rect 2774 4216 2780 4228
rect 2832 4216 2838 4268
rect 2869 4259 2927 4265
rect 2869 4225 2881 4259
rect 2915 4256 2927 4259
rect 3142 4256 3148 4268
rect 2915 4228 3148 4256
rect 2915 4225 2927 4228
rect 2869 4219 2927 4225
rect 3142 4216 3148 4228
rect 3200 4216 3206 4268
rect 3326 4216 3332 4268
rect 3384 4216 3390 4268
rect 1104 4098 8832 4120
rect 1104 4046 3579 4098
rect 3631 4046 3643 4098
rect 3695 4046 3707 4098
rect 3759 4046 3771 4098
rect 3823 4046 6176 4098
rect 6228 4046 6240 4098
rect 6292 4046 6304 4098
rect 6356 4046 6368 4098
rect 6420 4046 8832 4098
rect 1104 4024 8832 4046
rect 3053 3987 3111 3993
rect 3053 3953 3065 3987
rect 3099 3984 3111 3987
rect 3326 3984 3332 3996
rect 3099 3956 3332 3984
rect 3099 3953 3111 3956
rect 3053 3947 3111 3953
rect 3326 3944 3332 3956
rect 3384 3944 3390 3996
rect 4338 3916 4344 3928
rect 4299 3888 4344 3916
rect 4338 3876 4344 3888
rect 4396 3876 4402 3928
rect 4614 3876 4620 3928
rect 4672 3916 4678 3928
rect 4672 3888 4830 3916
rect 4672 3876 4678 3888
rect 2869 3851 2927 3857
rect 2869 3817 2881 3851
rect 2915 3848 2927 3851
rect 2958 3848 2964 3860
rect 2915 3820 2964 3848
rect 2915 3817 2927 3820
rect 2869 3811 2927 3817
rect 2958 3808 2964 3820
rect 3016 3808 3022 3860
rect 2774 3740 2780 3792
rect 2832 3780 2838 3792
rect 4062 3780 4068 3792
rect 2832 3752 4068 3780
rect 2832 3740 2838 3752
rect 4062 3740 4068 3752
rect 4120 3740 4126 3792
rect 6089 3783 6147 3789
rect 6089 3749 6101 3783
rect 6135 3749 6147 3783
rect 6089 3743 6147 3749
rect 4154 3604 4160 3656
rect 4212 3644 4218 3656
rect 6104 3644 6132 3743
rect 4212 3616 6132 3644
rect 4212 3604 4218 3616
rect 1104 3554 8832 3576
rect 1104 3502 2280 3554
rect 2332 3502 2344 3554
rect 2396 3502 2408 3554
rect 2460 3502 2472 3554
rect 2524 3502 4878 3554
rect 4930 3502 4942 3554
rect 4994 3502 5006 3554
rect 5058 3502 5070 3554
rect 5122 3502 7475 3554
rect 7527 3502 7539 3554
rect 7591 3502 7603 3554
rect 7655 3502 7667 3554
rect 7719 3502 8832 3554
rect 1104 3480 8832 3502
rect 1670 3449 1676 3452
rect 1660 3443 1676 3449
rect 1660 3409 1672 3443
rect 1660 3403 1676 3409
rect 1670 3400 1676 3403
rect 1728 3400 1734 3452
rect 5258 3440 5264 3452
rect 5219 3412 5264 3440
rect 5258 3400 5264 3412
rect 5316 3400 5322 3452
rect 2774 3332 2780 3384
rect 2832 3332 2838 3384
rect 1397 3307 1455 3313
rect 1397 3273 1409 3307
rect 1443 3304 1455 3307
rect 2792 3304 2820 3332
rect 1443 3276 2820 3304
rect 1443 3273 1455 3276
rect 1397 3267 1455 3273
rect 4246 3196 4252 3248
rect 4304 3236 4310 3248
rect 4890 3236 4896 3248
rect 4304 3208 4896 3236
rect 4304 3196 4310 3208
rect 4890 3196 4896 3208
rect 4948 3236 4954 3248
rect 5169 3239 5227 3245
rect 5169 3236 5181 3239
rect 4948 3208 5181 3236
rect 4948 3196 4954 3208
rect 5169 3205 5181 3208
rect 5215 3205 5227 3239
rect 6822 3236 6828 3248
rect 6783 3208 6828 3236
rect 5169 3199 5227 3205
rect 6822 3196 6828 3208
rect 6880 3196 6886 3248
rect 3050 3168 3056 3180
rect 2898 3140 3056 3168
rect 3050 3128 3056 3140
rect 3108 3128 3114 3180
rect 3418 3168 3424 3180
rect 3379 3140 3424 3168
rect 3418 3128 3424 3140
rect 3476 3128 3482 3180
rect 4985 3171 5043 3177
rect 4985 3137 4997 3171
rect 5031 3168 5043 3171
rect 6840 3168 6868 3196
rect 5031 3140 6868 3168
rect 5031 3137 5043 3140
rect 4985 3131 5043 3137
rect 6914 3060 6920 3112
rect 6972 3100 6978 3112
rect 6972 3072 7017 3100
rect 6972 3060 6978 3072
rect 1104 3010 8832 3032
rect 1104 2958 3579 3010
rect 3631 2958 3643 3010
rect 3695 2958 3707 3010
rect 3759 2958 3771 3010
rect 3823 2958 6176 3010
rect 6228 2958 6240 3010
rect 6292 2958 6304 3010
rect 6356 2958 6368 3010
rect 6420 2958 8832 3010
rect 1104 2936 8832 2958
rect 3050 2896 3056 2908
rect 3011 2868 3056 2896
rect 3050 2856 3056 2868
rect 3108 2856 3114 2908
rect 2869 2763 2927 2769
rect 2869 2729 2881 2763
rect 2915 2760 2927 2763
rect 2958 2760 2964 2772
rect 2915 2732 2964 2760
rect 2915 2729 2927 2732
rect 2869 2723 2927 2729
rect 2958 2720 2964 2732
rect 3016 2720 3022 2772
rect 4890 2720 4896 2772
rect 4948 2760 4954 2772
rect 4985 2763 5043 2769
rect 4985 2760 4997 2763
rect 4948 2732 4997 2760
rect 4948 2720 4954 2732
rect 4985 2729 4997 2732
rect 5031 2729 5043 2763
rect 4985 2723 5043 2729
rect 5077 2763 5135 2769
rect 5077 2729 5089 2763
rect 5123 2760 5135 2763
rect 6914 2760 6920 2772
rect 5123 2732 6920 2760
rect 5123 2729 5135 2732
rect 5077 2723 5135 2729
rect 6914 2720 6920 2732
rect 6972 2720 6978 2772
rect 4062 2516 4068 2568
rect 4120 2556 4126 2568
rect 5261 2559 5319 2565
rect 5261 2556 5273 2559
rect 4120 2528 5273 2556
rect 4120 2516 4126 2528
rect 5261 2525 5273 2528
rect 5307 2525 5319 2559
rect 5261 2519 5319 2525
rect 1104 2466 8832 2488
rect 1104 2414 2280 2466
rect 2332 2414 2344 2466
rect 2396 2414 2408 2466
rect 2460 2414 2472 2466
rect 2524 2414 4878 2466
rect 4930 2414 4942 2466
rect 4994 2414 5006 2466
rect 5058 2414 5070 2466
rect 5122 2414 7475 2466
rect 7527 2414 7539 2466
rect 7591 2414 7603 2466
rect 7655 2414 7667 2466
rect 7719 2414 8832 2466
rect 1104 2392 8832 2414
rect 4525 2355 4583 2361
rect 4525 2321 4537 2355
rect 4571 2352 4583 2355
rect 4614 2352 4620 2364
rect 4571 2324 4620 2352
rect 4571 2321 4583 2324
rect 4525 2315 4583 2321
rect 4614 2312 4620 2324
rect 4672 2312 4678 2364
rect 2958 2108 2964 2160
rect 3016 2148 3022 2160
rect 4341 2151 4399 2157
rect 4341 2148 4353 2151
rect 3016 2120 4353 2148
rect 3016 2108 3022 2120
rect 4341 2117 4353 2120
rect 4387 2117 4399 2151
rect 4341 2111 4399 2117
rect 1104 1922 8832 1944
rect 1104 1870 3579 1922
rect 3631 1870 3643 1922
rect 3695 1870 3707 1922
rect 3759 1870 3771 1922
rect 3823 1870 6176 1922
rect 6228 1870 6240 1922
rect 6292 1870 6304 1922
rect 6356 1870 6368 1922
rect 6420 1870 8832 1922
rect 1104 1848 8832 1870
rect 1104 1378 8832 1400
rect 1104 1326 2280 1378
rect 2332 1326 2344 1378
rect 2396 1326 2408 1378
rect 2460 1326 2472 1378
rect 2524 1326 4878 1378
rect 4930 1326 4942 1378
rect 4994 1326 5006 1378
rect 5058 1326 5070 1378
rect 5122 1326 7475 1378
rect 7527 1326 7539 1378
rect 7591 1326 7603 1378
rect 7655 1326 7667 1378
rect 7719 1326 8832 1378
rect 1104 1304 8832 1326
<< via1 >>
rect 4068 22644 4120 22696
rect 5172 22644 5224 22696
rect 3579 21454 3631 21506
rect 3643 21454 3695 21506
rect 3707 21454 3759 21506
rect 3771 21454 3823 21506
rect 6176 21454 6228 21506
rect 6240 21454 6292 21506
rect 6304 21454 6356 21506
rect 6368 21454 6420 21506
rect 2280 20910 2332 20962
rect 2344 20910 2396 20962
rect 2408 20910 2460 20962
rect 2472 20910 2524 20962
rect 4878 20910 4930 20962
rect 4942 20910 4994 20962
rect 5006 20910 5058 20962
rect 5070 20910 5122 20962
rect 7475 20910 7527 20962
rect 7539 20910 7591 20962
rect 7603 20910 7655 20962
rect 7667 20910 7719 20962
rect 3579 20366 3631 20418
rect 3643 20366 3695 20418
rect 3707 20366 3759 20418
rect 3771 20366 3823 20418
rect 6176 20366 6228 20418
rect 6240 20366 6292 20418
rect 6304 20366 6356 20418
rect 6368 20366 6420 20418
rect 2280 19822 2332 19874
rect 2344 19822 2396 19874
rect 2408 19822 2460 19874
rect 2472 19822 2524 19874
rect 4878 19822 4930 19874
rect 4942 19822 4994 19874
rect 5006 19822 5058 19874
rect 5070 19822 5122 19874
rect 7475 19822 7527 19874
rect 7539 19822 7591 19874
rect 7603 19822 7655 19874
rect 7667 19822 7719 19874
rect 3424 19627 3476 19636
rect 3424 19593 3433 19627
rect 3433 19593 3467 19627
rect 3467 19593 3476 19627
rect 3424 19584 3476 19593
rect 1400 19559 1452 19568
rect 1400 19525 1409 19559
rect 1409 19525 1443 19559
rect 1443 19525 1452 19559
rect 1400 19516 1452 19525
rect 1952 19448 2004 19500
rect 3332 19380 3384 19432
rect 3579 19278 3631 19330
rect 3643 19278 3695 19330
rect 3707 19278 3759 19330
rect 3771 19278 3823 19330
rect 6176 19278 6228 19330
rect 6240 19278 6292 19330
rect 6304 19278 6356 19330
rect 6368 19278 6420 19330
rect 1768 19040 1820 19092
rect 4068 19015 4120 19024
rect 4068 18981 4077 19015
rect 4077 18981 4111 19015
rect 4111 18981 4120 19015
rect 4068 18972 4120 18981
rect 5356 18972 5408 19024
rect 5540 18972 5592 19024
rect 2136 18836 2188 18888
rect 2688 18836 2740 18888
rect 2280 18734 2332 18786
rect 2344 18734 2396 18786
rect 2408 18734 2460 18786
rect 2472 18734 2524 18786
rect 4878 18734 4930 18786
rect 4942 18734 4994 18786
rect 5006 18734 5058 18786
rect 5070 18734 5122 18786
rect 7475 18734 7527 18786
rect 7539 18734 7591 18786
rect 7603 18734 7655 18786
rect 7667 18734 7719 18786
rect 5540 18675 5592 18684
rect 5540 18641 5549 18675
rect 5549 18641 5583 18675
rect 5583 18641 5592 18675
rect 5540 18632 5592 18641
rect 1676 18539 1728 18548
rect 1676 18505 1685 18539
rect 1685 18505 1719 18539
rect 1719 18505 1728 18539
rect 1676 18496 1728 18505
rect 2688 18496 2740 18548
rect 1400 18471 1452 18480
rect 1400 18437 1409 18471
rect 1409 18437 1443 18471
rect 1443 18437 1452 18471
rect 1400 18428 1452 18437
rect 3056 18428 3108 18480
rect 4528 18428 4580 18480
rect 2136 18360 2188 18412
rect 4436 18335 4488 18344
rect 4436 18301 4445 18335
rect 4445 18301 4479 18335
rect 4479 18301 4488 18335
rect 4436 18292 4488 18301
rect 3579 18190 3631 18242
rect 3643 18190 3695 18242
rect 3707 18190 3759 18242
rect 3771 18190 3823 18242
rect 6176 18190 6228 18242
rect 6240 18190 6292 18242
rect 6304 18190 6356 18242
rect 6368 18190 6420 18242
rect 1952 18131 2004 18140
rect 1952 18097 1961 18131
rect 1961 18097 1995 18131
rect 1995 18097 2004 18131
rect 1952 18088 2004 18097
rect 1768 17995 1820 18004
rect 1768 17961 1777 17995
rect 1777 17961 1811 17995
rect 1811 17961 1820 17995
rect 1768 17952 1820 17961
rect 4528 18088 4580 18140
rect 3332 18020 3384 18072
rect 4436 18020 4488 18072
rect 2964 17884 3016 17936
rect 4068 17927 4120 17936
rect 4068 17893 4077 17927
rect 4077 17893 4111 17927
rect 4111 17893 4120 17927
rect 4068 17884 4120 17893
rect 4712 17884 4764 17936
rect 3056 17791 3108 17800
rect 3056 17757 3065 17791
rect 3065 17757 3099 17791
rect 3099 17757 3108 17791
rect 3056 17748 3108 17757
rect 2280 17646 2332 17698
rect 2344 17646 2396 17698
rect 2408 17646 2460 17698
rect 2472 17646 2524 17698
rect 4878 17646 4930 17698
rect 4942 17646 4994 17698
rect 5006 17646 5058 17698
rect 5070 17646 5122 17698
rect 7475 17646 7527 17698
rect 7539 17646 7591 17698
rect 7603 17646 7655 17698
rect 7667 17646 7719 17698
rect 1400 17544 1452 17596
rect 3424 17544 3476 17596
rect 1676 17451 1728 17460
rect 1676 17417 1685 17451
rect 1685 17417 1719 17451
rect 1719 17417 1728 17451
rect 1676 17408 1728 17417
rect 3332 17408 3384 17460
rect 3056 17340 3108 17392
rect 2964 17204 3016 17256
rect 3579 17102 3631 17154
rect 3643 17102 3695 17154
rect 3707 17102 3759 17154
rect 3771 17102 3823 17154
rect 6176 17102 6228 17154
rect 6240 17102 6292 17154
rect 6304 17102 6356 17154
rect 6368 17102 6420 17154
rect 5264 16932 5316 16984
rect 3424 16864 3476 16916
rect 4712 16796 4764 16848
rect 7104 16839 7156 16848
rect 7104 16805 7113 16839
rect 7113 16805 7147 16839
rect 7147 16805 7156 16839
rect 7104 16796 7156 16805
rect 6644 16660 6696 16712
rect 2280 16558 2332 16610
rect 2344 16558 2396 16610
rect 2408 16558 2460 16610
rect 2472 16558 2524 16610
rect 4878 16558 4930 16610
rect 4942 16558 4994 16610
rect 5006 16558 5058 16610
rect 5070 16558 5122 16610
rect 7475 16558 7527 16610
rect 7539 16558 7591 16610
rect 7603 16558 7655 16610
rect 7667 16558 7719 16610
rect 4712 16320 4764 16372
rect 2872 16252 2924 16304
rect 4528 16252 4580 16304
rect 5172 16227 5224 16236
rect 5172 16193 5181 16227
rect 5181 16193 5215 16227
rect 5215 16193 5224 16227
rect 5172 16184 5224 16193
rect 3579 16014 3631 16066
rect 3643 16014 3695 16066
rect 3707 16014 3759 16066
rect 3771 16014 3823 16066
rect 6176 16014 6228 16066
rect 6240 16014 6292 16066
rect 6304 16014 6356 16066
rect 6368 16014 6420 16066
rect 5264 15955 5316 15964
rect 5264 15921 5273 15955
rect 5273 15921 5307 15955
rect 5307 15921 5316 15955
rect 5264 15912 5316 15921
rect 4712 15776 4764 15828
rect 7104 15776 7156 15828
rect 7380 15819 7432 15828
rect 7380 15785 7389 15819
rect 7389 15785 7423 15819
rect 7423 15785 7432 15819
rect 7380 15776 7432 15785
rect 6828 15708 6880 15760
rect 2280 15470 2332 15522
rect 2344 15470 2396 15522
rect 2408 15470 2460 15522
rect 2472 15470 2524 15522
rect 4878 15470 4930 15522
rect 4942 15470 4994 15522
rect 5006 15470 5058 15522
rect 5070 15470 5122 15522
rect 7475 15470 7527 15522
rect 7539 15470 7591 15522
rect 7603 15470 7655 15522
rect 7667 15470 7719 15522
rect 2872 15232 2924 15284
rect 4160 15232 4212 15284
rect 5540 15232 5592 15284
rect 5908 15300 5960 15352
rect 5816 15275 5868 15284
rect 5816 15241 5825 15275
rect 5825 15241 5859 15275
rect 5859 15241 5868 15275
rect 5816 15232 5868 15241
rect 1676 15139 1728 15148
rect 1676 15105 1685 15139
rect 1685 15105 1719 15139
rect 1719 15105 1728 15139
rect 1676 15096 1728 15105
rect 2688 15096 2740 15148
rect 3424 15139 3476 15148
rect 3424 15105 3433 15139
rect 3433 15105 3467 15139
rect 3467 15105 3476 15139
rect 3424 15096 3476 15105
rect 5632 15096 5684 15148
rect 5908 15164 5960 15216
rect 5816 15096 5868 15148
rect 7656 15071 7708 15080
rect 7656 15037 7665 15071
rect 7665 15037 7699 15071
rect 7699 15037 7708 15071
rect 7656 15028 7708 15037
rect 3579 14926 3631 14978
rect 3643 14926 3695 14978
rect 3707 14926 3759 14978
rect 3771 14926 3823 14978
rect 6176 14926 6228 14978
rect 6240 14926 6292 14978
rect 6304 14926 6356 14978
rect 6368 14926 6420 14978
rect 4528 14824 4580 14876
rect 5172 14824 5224 14876
rect 1768 14688 1820 14740
rect 2872 14688 2924 14740
rect 7012 14731 7064 14740
rect 7012 14697 7021 14731
rect 7021 14697 7055 14731
rect 7055 14697 7064 14731
rect 7012 14688 7064 14697
rect 7380 14731 7432 14740
rect 7380 14697 7389 14731
rect 7389 14697 7423 14731
rect 7423 14697 7432 14731
rect 7380 14688 7432 14697
rect 7656 14731 7708 14740
rect 7656 14697 7665 14731
rect 7665 14697 7699 14731
rect 7699 14697 7708 14731
rect 7656 14688 7708 14697
rect 3148 14552 3200 14604
rect 5448 14552 5500 14604
rect 2136 14484 2188 14536
rect 2280 14382 2332 14434
rect 2344 14382 2396 14434
rect 2408 14382 2460 14434
rect 2472 14382 2524 14434
rect 4878 14382 4930 14434
rect 4942 14382 4994 14434
rect 5006 14382 5058 14434
rect 5070 14382 5122 14434
rect 7475 14382 7527 14434
rect 7539 14382 7591 14434
rect 7603 14382 7655 14434
rect 7667 14382 7719 14434
rect 5632 14280 5684 14332
rect 3056 14144 3108 14196
rect 1400 14119 1452 14128
rect 1400 14085 1409 14119
rect 1409 14085 1443 14119
rect 1443 14085 1452 14119
rect 1400 14076 1452 14085
rect 3240 14076 3292 14128
rect 5908 14212 5960 14264
rect 6736 14212 6788 14264
rect 5816 14187 5868 14196
rect 5816 14153 5825 14187
rect 5825 14153 5859 14187
rect 5859 14153 5868 14187
rect 5816 14144 5868 14153
rect 6644 14144 6696 14196
rect 1676 14051 1728 14060
rect 1676 14017 1685 14051
rect 1685 14017 1719 14051
rect 1719 14017 1728 14051
rect 1676 14008 1728 14017
rect 2136 14008 2188 14060
rect 3056 13940 3108 13992
rect 5724 14119 5776 14128
rect 5724 14085 5733 14119
rect 5733 14085 5767 14119
rect 5767 14085 5776 14119
rect 5724 14076 5776 14085
rect 7104 14119 7156 14128
rect 7104 14085 7113 14119
rect 7113 14085 7147 14119
rect 7147 14085 7156 14119
rect 7104 14076 7156 14085
rect 6000 14008 6052 14060
rect 6828 13940 6880 13992
rect 3579 13838 3631 13890
rect 3643 13838 3695 13890
rect 3707 13838 3759 13890
rect 3771 13838 3823 13890
rect 6176 13838 6228 13890
rect 6240 13838 6292 13890
rect 6304 13838 6356 13890
rect 6368 13838 6420 13890
rect 5540 13736 5592 13788
rect 4528 13711 4580 13720
rect 4528 13677 4537 13711
rect 4537 13677 4571 13711
rect 4571 13677 4580 13711
rect 4528 13668 4580 13677
rect 5264 13668 5316 13720
rect 3976 13600 4028 13652
rect 7196 13643 7248 13652
rect 7196 13609 7205 13643
rect 7205 13609 7239 13643
rect 7239 13609 7248 13643
rect 7196 13600 7248 13609
rect 7840 13600 7892 13652
rect 3056 13532 3108 13584
rect 3884 13532 3936 13584
rect 5632 13464 5684 13516
rect 2872 13396 2924 13448
rect 4068 13396 4120 13448
rect 7012 13396 7064 13448
rect 7288 13396 7340 13448
rect 2280 13294 2332 13346
rect 2344 13294 2396 13346
rect 2408 13294 2460 13346
rect 2472 13294 2524 13346
rect 4878 13294 4930 13346
rect 4942 13294 4994 13346
rect 5006 13294 5058 13346
rect 5070 13294 5122 13346
rect 7475 13294 7527 13346
rect 7539 13294 7591 13346
rect 7603 13294 7655 13346
rect 7667 13294 7719 13346
rect 1768 13056 1820 13108
rect 3424 13192 3476 13244
rect 7196 13192 7248 13244
rect 3240 13056 3292 13108
rect 5632 13056 5684 13108
rect 4712 12988 4764 13040
rect 6828 12988 6880 13040
rect 2964 12920 3016 12972
rect 7012 12963 7064 12972
rect 7012 12929 7021 12963
rect 7021 12929 7055 12963
rect 7055 12929 7064 12963
rect 7012 12920 7064 12929
rect 3056 12852 3108 12904
rect 5172 12852 5224 12904
rect 3579 12750 3631 12802
rect 3643 12750 3695 12802
rect 3707 12750 3759 12802
rect 3771 12750 3823 12802
rect 6176 12750 6228 12802
rect 6240 12750 6292 12802
rect 6304 12750 6356 12802
rect 6368 12750 6420 12802
rect 2964 12648 3016 12700
rect 4712 12648 4764 12700
rect 6552 12580 6604 12632
rect 2964 12512 3016 12564
rect 3884 12444 3936 12496
rect 5540 12487 5592 12496
rect 5540 12453 5549 12487
rect 5549 12453 5583 12487
rect 5583 12453 5592 12487
rect 5540 12444 5592 12453
rect 6000 12444 6052 12496
rect 2280 12206 2332 12258
rect 2344 12206 2396 12258
rect 2408 12206 2460 12258
rect 2472 12206 2524 12258
rect 4878 12206 4930 12258
rect 4942 12206 4994 12258
rect 5006 12206 5058 12258
rect 5070 12206 5122 12258
rect 7475 12206 7527 12258
rect 7539 12206 7591 12258
rect 7603 12206 7655 12258
rect 7667 12206 7719 12258
rect 3148 12104 3200 12156
rect 7012 12104 7064 12156
rect 3884 12011 3936 12020
rect 3884 11977 3893 12011
rect 3893 11977 3927 12011
rect 3927 11977 3936 12011
rect 3884 11968 3936 11977
rect 5448 11968 5500 12020
rect 2964 11900 3016 11952
rect 5908 11943 5960 11952
rect 5908 11909 5917 11943
rect 5917 11909 5951 11943
rect 5951 11909 5960 11943
rect 5908 11900 5960 11909
rect 5172 11832 5224 11884
rect 3579 11662 3631 11714
rect 3643 11662 3695 11714
rect 3707 11662 3759 11714
rect 3771 11662 3823 11714
rect 6176 11662 6228 11714
rect 6240 11662 6292 11714
rect 6304 11662 6356 11714
rect 6368 11662 6420 11714
rect 2688 11560 2740 11612
rect 5264 11603 5316 11612
rect 5264 11569 5273 11603
rect 5273 11569 5307 11603
rect 5307 11569 5316 11603
rect 5264 11560 5316 11569
rect 6552 11560 6604 11612
rect 2044 11424 2096 11476
rect 4712 11424 4764 11476
rect 2280 11118 2332 11170
rect 2344 11118 2396 11170
rect 2408 11118 2460 11170
rect 2472 11118 2524 11170
rect 4878 11118 4930 11170
rect 4942 11118 4994 11170
rect 5006 11118 5058 11170
rect 5070 11118 5122 11170
rect 7475 11118 7527 11170
rect 7539 11118 7591 11170
rect 7603 11118 7655 11170
rect 7667 11118 7719 11170
rect 2872 11016 2924 11068
rect 1676 10880 1728 10932
rect 1676 10787 1728 10796
rect 1676 10753 1685 10787
rect 1685 10753 1719 10787
rect 1719 10753 1728 10787
rect 1676 10744 1728 10753
rect 1952 10744 2004 10796
rect 6644 10744 6696 10796
rect 3976 10676 4028 10728
rect 3579 10574 3631 10626
rect 3643 10574 3695 10626
rect 3707 10574 3759 10626
rect 3771 10574 3823 10626
rect 6176 10574 6228 10626
rect 6240 10574 6292 10626
rect 6304 10574 6356 10626
rect 6368 10574 6420 10626
rect 1860 10336 1912 10388
rect 2136 10200 2188 10252
rect 2280 10030 2332 10082
rect 2344 10030 2396 10082
rect 2408 10030 2460 10082
rect 2472 10030 2524 10082
rect 4878 10030 4930 10082
rect 4942 10030 4994 10082
rect 5006 10030 5058 10082
rect 5070 10030 5122 10082
rect 7475 10030 7527 10082
rect 7539 10030 7591 10082
rect 7603 10030 7655 10082
rect 7667 10030 7719 10082
rect 3424 9835 3476 9844
rect 3424 9801 3433 9835
rect 3433 9801 3467 9835
rect 3467 9801 3476 9835
rect 3424 9792 3476 9801
rect 3884 9724 3936 9776
rect 6828 9724 6880 9776
rect 7288 9767 7340 9776
rect 7288 9733 7297 9767
rect 7297 9733 7331 9767
rect 7331 9733 7340 9767
rect 7288 9724 7340 9733
rect 1676 9699 1728 9708
rect 1676 9665 1685 9699
rect 1685 9665 1719 9699
rect 1719 9665 1728 9699
rect 1676 9656 1728 9665
rect 2136 9656 2188 9708
rect 8208 9656 8260 9708
rect 3579 9486 3631 9538
rect 3643 9486 3695 9538
rect 3707 9486 3759 9538
rect 3771 9486 3823 9538
rect 6176 9486 6228 9538
rect 6240 9486 6292 9538
rect 6304 9486 6356 9538
rect 6368 9486 6420 9538
rect 1952 9427 2004 9436
rect 1952 9393 1961 9427
rect 1961 9393 1995 9427
rect 1995 9393 2004 9427
rect 1952 9384 2004 9393
rect 7012 9316 7064 9368
rect 2044 9248 2096 9300
rect 2688 9248 2740 9300
rect 2964 9248 3016 9300
rect 4712 9248 4764 9300
rect 3884 9180 3936 9232
rect 6828 9223 6880 9232
rect 6828 9189 6837 9223
rect 6837 9189 6871 9223
rect 6871 9189 6880 9223
rect 6828 9180 6880 9189
rect 2688 9044 2740 9096
rect 2280 8942 2332 8994
rect 2344 8942 2396 8994
rect 2408 8942 2460 8994
rect 2472 8942 2524 8994
rect 4878 8942 4930 8994
rect 4942 8942 4994 8994
rect 5006 8942 5058 8994
rect 5070 8942 5122 8994
rect 7475 8942 7527 8994
rect 7539 8942 7591 8994
rect 7603 8942 7655 8994
rect 7667 8942 7719 8994
rect 7012 8883 7064 8892
rect 1860 8772 1912 8824
rect 1676 8704 1728 8756
rect 7012 8849 7021 8883
rect 7021 8849 7055 8883
rect 7055 8849 7064 8883
rect 7012 8840 7064 8849
rect 2504 8679 2556 8688
rect 2504 8645 2513 8679
rect 2513 8645 2547 8679
rect 2547 8645 2556 8679
rect 2504 8636 2556 8645
rect 4068 8636 4120 8688
rect 7472 8636 7524 8688
rect 3056 8568 3108 8620
rect 4620 8568 4672 8620
rect 5448 8500 5500 8552
rect 3579 8398 3631 8450
rect 3643 8398 3695 8450
rect 3707 8398 3759 8450
rect 3771 8398 3823 8450
rect 6176 8398 6228 8450
rect 6240 8398 6292 8450
rect 6304 8398 6356 8450
rect 6368 8398 6420 8450
rect 3056 8339 3108 8348
rect 3056 8305 3065 8339
rect 3065 8305 3099 8339
rect 3099 8305 3108 8339
rect 3056 8296 3108 8305
rect 5540 8296 5592 8348
rect 7472 8339 7524 8348
rect 3976 8228 4028 8280
rect 5724 8228 5776 8280
rect 7472 8305 7481 8339
rect 7481 8305 7515 8339
rect 7515 8305 7524 8339
rect 7472 8296 7524 8305
rect 2136 8092 2188 8144
rect 2688 8092 2740 8144
rect 4160 8092 4212 8144
rect 4712 8135 4764 8144
rect 4712 8101 4721 8135
rect 4721 8101 4755 8135
rect 4755 8101 4764 8135
rect 4712 8092 4764 8101
rect 2504 8024 2556 8076
rect 4436 7956 4488 8008
rect 5264 7956 5316 8008
rect 2280 7854 2332 7906
rect 2344 7854 2396 7906
rect 2408 7854 2460 7906
rect 2472 7854 2524 7906
rect 4878 7854 4930 7906
rect 4942 7854 4994 7906
rect 5006 7854 5058 7906
rect 5070 7854 5122 7906
rect 7475 7854 7527 7906
rect 7539 7854 7591 7906
rect 7603 7854 7655 7906
rect 7667 7854 7719 7906
rect 3332 7752 3384 7804
rect 5724 7795 5776 7804
rect 2964 7548 3016 7600
rect 4068 7684 4120 7736
rect 5724 7761 5733 7795
rect 5733 7761 5767 7795
rect 5767 7761 5776 7795
rect 5724 7752 5776 7761
rect 5908 7684 5960 7736
rect 4436 7591 4488 7600
rect 4436 7557 4445 7591
rect 4445 7557 4479 7591
rect 4479 7557 4488 7591
rect 4436 7548 4488 7557
rect 3148 7412 3200 7464
rect 4068 7412 4120 7464
rect 5632 7412 5684 7464
rect 3579 7310 3631 7362
rect 3643 7310 3695 7362
rect 3707 7310 3759 7362
rect 3771 7310 3823 7362
rect 6176 7310 6228 7362
rect 6240 7310 6292 7362
rect 6304 7310 6356 7362
rect 6368 7310 6420 7362
rect 4712 7208 4764 7260
rect 5724 7072 5776 7124
rect 4160 7004 4212 7056
rect 5632 7004 5684 7056
rect 2280 6766 2332 6818
rect 2344 6766 2396 6818
rect 2408 6766 2460 6818
rect 2472 6766 2524 6818
rect 4878 6766 4930 6818
rect 4942 6766 4994 6818
rect 5006 6766 5058 6818
rect 5070 6766 5122 6818
rect 7475 6766 7527 6818
rect 7539 6766 7591 6818
rect 7603 6766 7655 6818
rect 7667 6766 7719 6818
rect 5724 6664 5776 6716
rect 3148 6528 3200 6580
rect 1400 6503 1452 6512
rect 1400 6469 1409 6503
rect 1409 6469 1443 6503
rect 1443 6469 1452 6503
rect 1400 6460 1452 6469
rect 4620 6460 4672 6512
rect 1676 6435 1728 6444
rect 1676 6401 1685 6435
rect 1685 6401 1719 6435
rect 1719 6401 1728 6435
rect 1676 6392 1728 6401
rect 2688 6392 2740 6444
rect 3424 6435 3476 6444
rect 3424 6401 3433 6435
rect 3433 6401 3467 6435
rect 3467 6401 3476 6435
rect 3424 6392 3476 6401
rect 4436 6367 4488 6376
rect 4436 6333 4445 6367
rect 4445 6333 4479 6367
rect 4479 6333 4488 6367
rect 4436 6324 4488 6333
rect 3579 6222 3631 6274
rect 3643 6222 3695 6274
rect 3707 6222 3759 6274
rect 3771 6222 3823 6274
rect 6176 6222 6228 6274
rect 6240 6222 6292 6274
rect 6304 6222 6356 6274
rect 6368 6222 6420 6274
rect 1952 5984 2004 6036
rect 2136 6027 2188 6036
rect 2136 5993 2145 6027
rect 2145 5993 2179 6027
rect 2179 5993 2188 6027
rect 2136 5984 2188 5993
rect 1400 5916 1452 5968
rect 4160 5916 4212 5968
rect 2136 5780 2188 5832
rect 2280 5678 2332 5730
rect 2344 5678 2396 5730
rect 2408 5678 2460 5730
rect 2472 5678 2524 5730
rect 4878 5678 4930 5730
rect 4942 5678 4994 5730
rect 5006 5678 5058 5730
rect 5070 5678 5122 5730
rect 7475 5678 7527 5730
rect 7539 5678 7591 5730
rect 7603 5678 7655 5730
rect 7667 5678 7719 5730
rect 1400 5483 1452 5492
rect 1400 5449 1409 5483
rect 1409 5449 1443 5483
rect 1443 5449 1452 5483
rect 1400 5440 1452 5449
rect 1768 5440 1820 5492
rect 2136 5304 2188 5356
rect 1676 5236 1728 5288
rect 3579 5134 3631 5186
rect 3643 5134 3695 5186
rect 3707 5134 3759 5186
rect 3771 5134 3823 5186
rect 6176 5134 6228 5186
rect 6240 5134 6292 5186
rect 6304 5134 6356 5186
rect 6368 5134 6420 5186
rect 2688 5032 2740 5084
rect 3332 5032 3384 5084
rect 6552 5032 6604 5084
rect 3148 4964 3200 5016
rect 3424 4964 3476 5016
rect 4436 4964 4488 5016
rect 1952 4896 2004 4948
rect 4068 4939 4120 4948
rect 4068 4905 4077 4939
rect 4077 4905 4111 4939
rect 4111 4905 4120 4939
rect 4068 4896 4120 4905
rect 4344 4828 4396 4880
rect 5356 4828 5408 4880
rect 2280 4590 2332 4642
rect 2344 4590 2396 4642
rect 2408 4590 2460 4642
rect 2472 4590 2524 4642
rect 4878 4590 4930 4642
rect 4942 4590 4994 4642
rect 5006 4590 5058 4642
rect 5070 4590 5122 4642
rect 7475 4590 7527 4642
rect 7539 4590 7591 4642
rect 7603 4590 7655 4642
rect 7667 4590 7719 4642
rect 2872 4352 2924 4404
rect 2780 4216 2832 4268
rect 3148 4216 3200 4268
rect 3332 4216 3384 4268
rect 3579 4046 3631 4098
rect 3643 4046 3695 4098
rect 3707 4046 3759 4098
rect 3771 4046 3823 4098
rect 6176 4046 6228 4098
rect 6240 4046 6292 4098
rect 6304 4046 6356 4098
rect 6368 4046 6420 4098
rect 3332 3944 3384 3996
rect 4344 3919 4396 3928
rect 4344 3885 4353 3919
rect 4353 3885 4387 3919
rect 4387 3885 4396 3919
rect 4344 3876 4396 3885
rect 4620 3876 4672 3928
rect 2964 3808 3016 3860
rect 2780 3740 2832 3792
rect 4068 3783 4120 3792
rect 4068 3749 4077 3783
rect 4077 3749 4111 3783
rect 4111 3749 4120 3783
rect 4068 3740 4120 3749
rect 4160 3604 4212 3656
rect 2280 3502 2332 3554
rect 2344 3502 2396 3554
rect 2408 3502 2460 3554
rect 2472 3502 2524 3554
rect 4878 3502 4930 3554
rect 4942 3502 4994 3554
rect 5006 3502 5058 3554
rect 5070 3502 5122 3554
rect 7475 3502 7527 3554
rect 7539 3502 7591 3554
rect 7603 3502 7655 3554
rect 7667 3502 7719 3554
rect 1676 3443 1728 3452
rect 1676 3409 1706 3443
rect 1706 3409 1728 3443
rect 1676 3400 1728 3409
rect 5264 3443 5316 3452
rect 5264 3409 5273 3443
rect 5273 3409 5307 3443
rect 5307 3409 5316 3443
rect 5264 3400 5316 3409
rect 2780 3332 2832 3384
rect 4252 3196 4304 3248
rect 4896 3196 4948 3248
rect 6828 3239 6880 3248
rect 6828 3205 6837 3239
rect 6837 3205 6871 3239
rect 6871 3205 6880 3239
rect 6828 3196 6880 3205
rect 3056 3128 3108 3180
rect 3424 3171 3476 3180
rect 3424 3137 3433 3171
rect 3433 3137 3467 3171
rect 3467 3137 3476 3171
rect 3424 3128 3476 3137
rect 6920 3103 6972 3112
rect 6920 3069 6929 3103
rect 6929 3069 6963 3103
rect 6963 3069 6972 3103
rect 6920 3060 6972 3069
rect 3579 2958 3631 3010
rect 3643 2958 3695 3010
rect 3707 2958 3759 3010
rect 3771 2958 3823 3010
rect 6176 2958 6228 3010
rect 6240 2958 6292 3010
rect 6304 2958 6356 3010
rect 6368 2958 6420 3010
rect 3056 2899 3108 2908
rect 3056 2865 3065 2899
rect 3065 2865 3099 2899
rect 3099 2865 3108 2899
rect 3056 2856 3108 2865
rect 2964 2720 3016 2772
rect 4896 2720 4948 2772
rect 6920 2720 6972 2772
rect 4068 2516 4120 2568
rect 2280 2414 2332 2466
rect 2344 2414 2396 2466
rect 2408 2414 2460 2466
rect 2472 2414 2524 2466
rect 4878 2414 4930 2466
rect 4942 2414 4994 2466
rect 5006 2414 5058 2466
rect 5070 2414 5122 2466
rect 7475 2414 7527 2466
rect 7539 2414 7591 2466
rect 7603 2414 7655 2466
rect 7667 2414 7719 2466
rect 4620 2312 4672 2364
rect 2964 2108 3016 2160
rect 3579 1870 3631 1922
rect 3643 1870 3695 1922
rect 3707 1870 3759 1922
rect 3771 1870 3823 1922
rect 6176 1870 6228 1922
rect 6240 1870 6292 1922
rect 6304 1870 6356 1922
rect 6368 1870 6420 1922
rect 2280 1326 2332 1378
rect 2344 1326 2396 1378
rect 2408 1326 2460 1378
rect 2472 1326 2524 1378
rect 4878 1326 4930 1378
rect 4942 1326 4994 1378
rect 5006 1326 5058 1378
rect 5070 1326 5122 1378
rect 7475 1326 7527 1378
rect 7539 1326 7591 1378
rect 7603 1326 7655 1378
rect 7667 1326 7719 1378
<< metal2 >>
rect 4066 23344 4122 23353
rect 4066 23279 4122 23288
rect 4080 22702 4108 23279
rect 5814 22800 5870 22809
rect 5814 22735 5870 22744
rect 4068 22696 4120 22702
rect 4068 22638 4120 22644
rect 5172 22696 5224 22702
rect 5172 22638 5224 22644
rect 3422 21712 3478 21721
rect 3422 21647 3478 21656
rect 2254 20964 2550 20984
rect 2310 20962 2334 20964
rect 2390 20962 2414 20964
rect 2470 20962 2494 20964
rect 2332 20910 2334 20962
rect 2396 20910 2408 20962
rect 2470 20910 2472 20962
rect 2310 20908 2334 20910
rect 2390 20908 2414 20910
rect 2470 20908 2494 20910
rect 2254 20888 2550 20908
rect 3054 20080 3110 20089
rect 3054 20015 3110 20024
rect 2254 19876 2550 19896
rect 2310 19874 2334 19876
rect 2390 19874 2414 19876
rect 2470 19874 2494 19876
rect 2332 19822 2334 19874
rect 2396 19822 2408 19874
rect 2470 19822 2472 19874
rect 2310 19820 2334 19822
rect 2390 19820 2414 19822
rect 2470 19820 2494 19822
rect 2254 19800 2550 19820
rect 1400 19568 1452 19574
rect 1400 19510 1452 19516
rect 1412 18486 1440 19510
rect 1952 19500 2004 19506
rect 1952 19442 2004 19448
rect 1768 19092 1820 19098
rect 1768 19034 1820 19040
rect 1676 18548 1728 18554
rect 1676 18490 1728 18496
rect 1400 18480 1452 18486
rect 1400 18422 1452 18428
rect 1412 17602 1440 18422
rect 1400 17596 1452 17602
rect 1400 17538 1452 17544
rect 1412 14134 1440 17538
rect 1688 17466 1716 18490
rect 1780 18010 1808 19034
rect 1964 18146 1992 19442
rect 2136 18888 2188 18894
rect 2136 18830 2188 18836
rect 2688 18888 2740 18894
rect 2688 18830 2740 18836
rect 2148 18418 2176 18830
rect 2254 18788 2550 18808
rect 2310 18786 2334 18788
rect 2390 18786 2414 18788
rect 2470 18786 2494 18788
rect 2332 18734 2334 18786
rect 2396 18734 2408 18786
rect 2470 18734 2472 18786
rect 2310 18732 2334 18734
rect 2390 18732 2414 18734
rect 2470 18732 2494 18734
rect 2254 18712 2550 18732
rect 2700 18554 2728 18830
rect 2688 18548 2740 18554
rect 2688 18490 2740 18496
rect 3068 18486 3096 20015
rect 3436 19642 3464 21647
rect 3553 21508 3849 21528
rect 3609 21506 3633 21508
rect 3689 21506 3713 21508
rect 3769 21506 3793 21508
rect 3631 21454 3633 21506
rect 3695 21454 3707 21506
rect 3769 21454 3771 21506
rect 3609 21452 3633 21454
rect 3689 21452 3713 21454
rect 3769 21452 3793 21454
rect 3553 21432 3849 21452
rect 4852 20964 5148 20984
rect 4908 20962 4932 20964
rect 4988 20962 5012 20964
rect 5068 20962 5092 20964
rect 4930 20910 4932 20962
rect 4994 20910 5006 20962
rect 5068 20910 5070 20962
rect 4908 20908 4932 20910
rect 4988 20908 5012 20910
rect 5068 20908 5092 20910
rect 4852 20888 5148 20908
rect 3553 20420 3849 20440
rect 3609 20418 3633 20420
rect 3689 20418 3713 20420
rect 3769 20418 3793 20420
rect 3631 20366 3633 20418
rect 3695 20366 3707 20418
rect 3769 20366 3771 20418
rect 3609 20364 3633 20366
rect 3689 20364 3713 20366
rect 3769 20364 3793 20366
rect 3553 20344 3849 20364
rect 4852 19876 5148 19896
rect 4908 19874 4932 19876
rect 4988 19874 5012 19876
rect 5068 19874 5092 19876
rect 4930 19822 4932 19874
rect 4994 19822 5006 19874
rect 5068 19822 5070 19874
rect 4908 19820 4932 19822
rect 4988 19820 5012 19822
rect 5068 19820 5092 19822
rect 4852 19800 5148 19820
rect 3424 19636 3476 19642
rect 3424 19578 3476 19584
rect 3332 19432 3384 19438
rect 3332 19374 3384 19380
rect 3056 18480 3108 18486
rect 3056 18422 3108 18428
rect 2136 18412 2188 18418
rect 2136 18354 2188 18360
rect 3238 18312 3294 18321
rect 3238 18247 3294 18256
rect 1952 18140 2004 18146
rect 1952 18082 2004 18088
rect 1768 18004 1820 18010
rect 1768 17946 1820 17952
rect 1676 17460 1728 17466
rect 1676 17402 1728 17408
rect 1676 15148 1728 15154
rect 1676 15090 1728 15096
rect 1400 14128 1452 14134
rect 1400 14070 1452 14076
rect 1688 14066 1716 15090
rect 1780 14746 1808 17946
rect 2964 17936 3016 17942
rect 2964 17878 3016 17884
rect 2254 17700 2550 17720
rect 2310 17698 2334 17700
rect 2390 17698 2414 17700
rect 2470 17698 2494 17700
rect 2332 17646 2334 17698
rect 2396 17646 2408 17698
rect 2470 17646 2472 17698
rect 2310 17644 2334 17646
rect 2390 17644 2414 17646
rect 2470 17644 2494 17646
rect 2254 17624 2550 17644
rect 2976 17262 3004 17878
rect 3056 17800 3108 17806
rect 3056 17742 3108 17748
rect 3068 17398 3096 17742
rect 3056 17392 3108 17398
rect 3056 17334 3108 17340
rect 2964 17256 3016 17262
rect 2884 17204 2964 17210
rect 2884 17198 3016 17204
rect 2884 17182 3004 17198
rect 2254 16612 2550 16632
rect 2310 16610 2334 16612
rect 2390 16610 2414 16612
rect 2470 16610 2494 16612
rect 2332 16558 2334 16610
rect 2396 16558 2408 16610
rect 2470 16558 2472 16610
rect 2310 16556 2334 16558
rect 2390 16556 2414 16558
rect 2470 16556 2494 16558
rect 2254 16536 2550 16556
rect 2884 16310 2912 17182
rect 2872 16304 2924 16310
rect 2872 16246 2924 16252
rect 2254 15524 2550 15544
rect 2310 15522 2334 15524
rect 2390 15522 2414 15524
rect 2470 15522 2494 15524
rect 2332 15470 2334 15522
rect 2396 15470 2408 15522
rect 2470 15470 2472 15522
rect 2310 15468 2334 15470
rect 2390 15468 2414 15470
rect 2470 15468 2494 15470
rect 2254 15448 2550 15468
rect 2884 15290 2912 16246
rect 2872 15284 2924 15290
rect 2872 15226 2924 15232
rect 2688 15148 2740 15154
rect 2688 15090 2740 15096
rect 1768 14740 1820 14746
rect 1820 14700 1900 14728
rect 1768 14682 1820 14688
rect 1676 14060 1728 14066
rect 1676 14002 1728 14008
rect 1688 10938 1716 14002
rect 1768 13108 1820 13114
rect 1768 13050 1820 13056
rect 1676 10932 1728 10938
rect 1676 10874 1728 10880
rect 1676 10796 1728 10802
rect 1676 10738 1728 10744
rect 1688 9714 1716 10738
rect 1676 9708 1728 9714
rect 1676 9650 1728 9656
rect 1688 8762 1716 9650
rect 1676 8756 1728 8762
rect 1676 8698 1728 8704
rect 1400 6512 1452 6518
rect 1400 6454 1452 6460
rect 1412 5974 1440 6454
rect 1676 6444 1728 6450
rect 1676 6386 1728 6392
rect 1400 5968 1452 5974
rect 1400 5910 1452 5916
rect 1412 5498 1440 5910
rect 1400 5492 1452 5498
rect 1400 5434 1452 5440
rect 1688 5294 1716 6386
rect 1780 5498 1808 13050
rect 1872 10394 1900 14700
rect 2136 14536 2188 14542
rect 2136 14478 2188 14484
rect 2148 14066 2176 14478
rect 2254 14436 2550 14456
rect 2310 14434 2334 14436
rect 2390 14434 2414 14436
rect 2470 14434 2494 14436
rect 2332 14382 2334 14434
rect 2396 14382 2408 14434
rect 2470 14382 2472 14434
rect 2310 14380 2334 14382
rect 2390 14380 2414 14382
rect 2470 14380 2494 14382
rect 2254 14360 2550 14380
rect 2136 14060 2188 14066
rect 2136 14002 2188 14008
rect 2254 13348 2550 13368
rect 2310 13346 2334 13348
rect 2390 13346 2414 13348
rect 2470 13346 2494 13348
rect 2332 13294 2334 13346
rect 2396 13294 2408 13346
rect 2470 13294 2472 13346
rect 2310 13292 2334 13294
rect 2390 13292 2414 13294
rect 2470 13292 2494 13294
rect 2254 13272 2550 13292
rect 2254 12260 2550 12280
rect 2310 12258 2334 12260
rect 2390 12258 2414 12260
rect 2470 12258 2494 12260
rect 2332 12206 2334 12258
rect 2396 12206 2408 12258
rect 2470 12206 2472 12258
rect 2310 12204 2334 12206
rect 2390 12204 2414 12206
rect 2470 12204 2494 12206
rect 2254 12184 2550 12204
rect 2700 11618 2728 15090
rect 2884 14746 2912 15226
rect 3054 15048 3110 15057
rect 3054 14983 3110 14992
rect 2872 14740 2924 14746
rect 2872 14682 2924 14688
rect 2884 13454 2912 14682
rect 3068 14202 3096 14983
rect 3148 14604 3200 14610
rect 3148 14546 3200 14552
rect 3056 14196 3108 14202
rect 3056 14138 3108 14144
rect 3056 13992 3108 13998
rect 3056 13934 3108 13940
rect 3068 13590 3096 13934
rect 3056 13584 3108 13590
rect 3056 13526 3108 13532
rect 2872 13448 2924 13454
rect 2872 13390 2924 13396
rect 2688 11612 2740 11618
rect 2688 11554 2740 11560
rect 2044 11476 2096 11482
rect 2044 11418 2096 11424
rect 1952 10796 2004 10802
rect 1952 10738 2004 10744
rect 1860 10388 1912 10394
rect 1860 10330 1912 10336
rect 1872 8830 1900 10330
rect 1964 9442 1992 10738
rect 1952 9436 2004 9442
rect 1952 9378 2004 9384
rect 2056 9306 2084 11418
rect 2254 11172 2550 11192
rect 2310 11170 2334 11172
rect 2390 11170 2414 11172
rect 2470 11170 2494 11172
rect 2332 11118 2334 11170
rect 2396 11118 2408 11170
rect 2470 11118 2472 11170
rect 2310 11116 2334 11118
rect 2390 11116 2414 11118
rect 2470 11116 2494 11118
rect 2254 11096 2550 11116
rect 2884 11074 2912 13390
rect 2964 12972 3016 12978
rect 2964 12914 3016 12920
rect 2976 12706 3004 12914
rect 3068 12910 3096 13526
rect 3056 12904 3108 12910
rect 3056 12846 3108 12852
rect 2964 12700 3016 12706
rect 2964 12642 3016 12648
rect 2964 12564 3016 12570
rect 2964 12506 3016 12512
rect 2976 11958 3004 12506
rect 3160 12162 3188 14546
rect 3252 14134 3280 18247
rect 3344 18078 3372 19374
rect 3553 19332 3849 19352
rect 3609 19330 3633 19332
rect 3689 19330 3713 19332
rect 3769 19330 3793 19332
rect 3631 19278 3633 19330
rect 3695 19278 3707 19330
rect 3769 19278 3771 19330
rect 3609 19276 3633 19278
rect 3689 19276 3713 19278
rect 3769 19276 3793 19278
rect 3553 19256 3849 19276
rect 5184 19114 5212 22638
rect 5722 20080 5778 20089
rect 5722 20015 5778 20024
rect 5184 19086 5488 19114
rect 4068 19024 4120 19030
rect 4068 18966 4120 18972
rect 5356 19024 5408 19030
rect 5356 18966 5408 18972
rect 3553 18244 3849 18264
rect 3609 18242 3633 18244
rect 3689 18242 3713 18244
rect 3769 18242 3793 18244
rect 3631 18190 3633 18242
rect 3695 18190 3707 18242
rect 3769 18190 3771 18242
rect 3609 18188 3633 18190
rect 3689 18188 3713 18190
rect 3769 18188 3793 18190
rect 3553 18168 3849 18188
rect 3332 18072 3384 18078
rect 3332 18014 3384 18020
rect 3344 17466 3372 18014
rect 4080 17942 4108 18966
rect 4852 18788 5148 18808
rect 4908 18786 4932 18788
rect 4988 18786 5012 18788
rect 5068 18786 5092 18788
rect 4930 18734 4932 18786
rect 4994 18734 5006 18786
rect 5068 18734 5070 18786
rect 4908 18732 4932 18734
rect 4988 18732 5012 18734
rect 5068 18732 5092 18734
rect 4852 18712 5148 18732
rect 4528 18480 4580 18486
rect 4528 18422 4580 18428
rect 4436 18344 4488 18350
rect 4436 18286 4488 18292
rect 4448 18078 4476 18286
rect 4540 18146 4568 18422
rect 4528 18140 4580 18146
rect 4528 18082 4580 18088
rect 4436 18072 4488 18078
rect 4436 18014 4488 18020
rect 4068 17936 4120 17942
rect 4068 17878 4120 17884
rect 3424 17596 3476 17602
rect 3424 17538 3476 17544
rect 3332 17460 3384 17466
rect 3332 17402 3384 17408
rect 3436 16922 3464 17538
rect 3553 17156 3849 17176
rect 3609 17154 3633 17156
rect 3689 17154 3713 17156
rect 3769 17154 3793 17156
rect 3631 17102 3633 17154
rect 3695 17102 3707 17154
rect 3769 17102 3771 17154
rect 3609 17100 3633 17102
rect 3689 17100 3713 17102
rect 3769 17100 3793 17102
rect 3553 17080 3849 17100
rect 3424 16916 3476 16922
rect 3424 16858 3476 16864
rect 4066 16408 4122 16417
rect 4122 16366 4200 16394
rect 4066 16343 4122 16352
rect 3553 16068 3849 16088
rect 3609 16066 3633 16068
rect 3689 16066 3713 16068
rect 3769 16066 3793 16068
rect 3631 16014 3633 16066
rect 3695 16014 3707 16066
rect 3769 16014 3771 16066
rect 3609 16012 3633 16014
rect 3689 16012 3713 16014
rect 3769 16012 3793 16014
rect 3553 15992 3849 16012
rect 4172 15290 4200 16366
rect 4540 16310 4568 18082
rect 4712 17936 4764 17942
rect 4712 17878 4764 17884
rect 4724 16854 4752 17878
rect 4852 17700 5148 17720
rect 4908 17698 4932 17700
rect 4988 17698 5012 17700
rect 5068 17698 5092 17700
rect 4930 17646 4932 17698
rect 4994 17646 5006 17698
rect 5068 17646 5070 17698
rect 4908 17644 4932 17646
rect 4988 17644 5012 17646
rect 5068 17644 5092 17646
rect 4852 17624 5148 17644
rect 5264 16984 5316 16990
rect 5264 16926 5316 16932
rect 4712 16848 4764 16854
rect 4712 16790 4764 16796
rect 4724 16378 4752 16790
rect 4852 16612 5148 16632
rect 4908 16610 4932 16612
rect 4988 16610 5012 16612
rect 5068 16610 5092 16612
rect 4930 16558 4932 16610
rect 4994 16558 5006 16610
rect 5068 16558 5070 16610
rect 4908 16556 4932 16558
rect 4988 16556 5012 16558
rect 5068 16556 5092 16558
rect 4852 16536 5148 16556
rect 4712 16372 4764 16378
rect 4712 16314 4764 16320
rect 4528 16304 4580 16310
rect 4528 16246 4580 16252
rect 4540 16122 4568 16246
rect 5172 16236 5224 16242
rect 5172 16178 5224 16184
rect 4540 16094 4660 16122
rect 4160 15284 4212 15290
rect 4160 15226 4212 15232
rect 3424 15148 3476 15154
rect 3424 15090 3476 15096
rect 3240 14128 3292 14134
rect 3240 14070 3292 14076
rect 3436 13250 3464 15090
rect 3553 14980 3849 15000
rect 3609 14978 3633 14980
rect 3689 14978 3713 14980
rect 3769 14978 3793 14980
rect 3631 14926 3633 14978
rect 3695 14926 3707 14978
rect 3769 14926 3771 14978
rect 3609 14924 3633 14926
rect 3689 14924 3713 14926
rect 3769 14924 3793 14926
rect 3553 14904 3849 14924
rect 4528 14876 4580 14882
rect 4528 14818 4580 14824
rect 3553 13892 3849 13912
rect 3609 13890 3633 13892
rect 3689 13890 3713 13892
rect 3769 13890 3793 13892
rect 3631 13838 3633 13890
rect 3695 13838 3707 13890
rect 3769 13838 3771 13890
rect 3609 13836 3633 13838
rect 3689 13836 3713 13838
rect 3769 13836 3793 13838
rect 3553 13816 3849 13836
rect 4540 13726 4568 14818
rect 4528 13720 4580 13726
rect 4528 13662 4580 13668
rect 3976 13652 4028 13658
rect 3976 13594 4028 13600
rect 3884 13584 3936 13590
rect 3884 13526 3936 13532
rect 3424 13244 3476 13250
rect 3424 13186 3476 13192
rect 3240 13108 3292 13114
rect 3240 13050 3292 13056
rect 3148 12156 3200 12162
rect 3148 12098 3200 12104
rect 2964 11952 3016 11958
rect 2964 11894 3016 11900
rect 2872 11068 2924 11074
rect 2872 11010 2924 11016
rect 2136 10252 2188 10258
rect 2136 10194 2188 10200
rect 2148 9714 2176 10194
rect 2254 10084 2550 10104
rect 2310 10082 2334 10084
rect 2390 10082 2414 10084
rect 2470 10082 2494 10084
rect 2332 10030 2334 10082
rect 2396 10030 2408 10082
rect 2470 10030 2472 10082
rect 2310 10028 2334 10030
rect 2390 10028 2414 10030
rect 2470 10028 2494 10030
rect 2254 10008 2550 10028
rect 2136 9708 2188 9714
rect 2136 9650 2188 9656
rect 2976 9306 3004 11894
rect 3252 11657 3280 13050
rect 3553 12804 3849 12824
rect 3609 12802 3633 12804
rect 3689 12802 3713 12804
rect 3769 12802 3793 12804
rect 3631 12750 3633 12802
rect 3695 12750 3707 12802
rect 3769 12750 3771 12802
rect 3609 12748 3633 12750
rect 3689 12748 3713 12750
rect 3769 12748 3793 12750
rect 3553 12728 3849 12748
rect 3896 12502 3924 13526
rect 3884 12496 3936 12502
rect 3884 12438 3936 12444
rect 3896 12026 3924 12438
rect 3884 12020 3936 12026
rect 3884 11962 3936 11968
rect 3553 11716 3849 11736
rect 3609 11714 3633 11716
rect 3689 11714 3713 11716
rect 3769 11714 3793 11716
rect 3631 11662 3633 11714
rect 3695 11662 3707 11714
rect 3769 11662 3771 11714
rect 3609 11660 3633 11662
rect 3689 11660 3713 11662
rect 3769 11660 3793 11662
rect 3238 11648 3294 11657
rect 3553 11640 3849 11660
rect 3238 11583 3294 11592
rect 3553 10628 3849 10648
rect 3609 10626 3633 10628
rect 3689 10626 3713 10628
rect 3769 10626 3793 10628
rect 3631 10574 3633 10626
rect 3695 10574 3707 10626
rect 3769 10574 3771 10626
rect 3609 10572 3633 10574
rect 3689 10572 3713 10574
rect 3769 10572 3793 10574
rect 3553 10552 3849 10572
rect 3422 9880 3478 9889
rect 3422 9815 3424 9824
rect 3476 9815 3478 9824
rect 3424 9786 3476 9792
rect 3896 9782 3924 11962
rect 3988 10734 4016 13594
rect 4066 13552 4122 13561
rect 4066 13487 4122 13496
rect 4080 13454 4108 13487
rect 4068 13448 4120 13454
rect 4068 13390 4120 13396
rect 3976 10728 4028 10734
rect 3976 10670 4028 10676
rect 3884 9776 3936 9782
rect 3884 9718 3936 9724
rect 3553 9540 3849 9560
rect 3609 9538 3633 9540
rect 3689 9538 3713 9540
rect 3769 9538 3793 9540
rect 3631 9486 3633 9538
rect 3695 9486 3707 9538
rect 3769 9486 3771 9538
rect 3609 9484 3633 9486
rect 3689 9484 3713 9486
rect 3769 9484 3793 9486
rect 3553 9464 3849 9484
rect 2044 9300 2096 9306
rect 2044 9242 2096 9248
rect 2688 9300 2740 9306
rect 2688 9242 2740 9248
rect 2964 9300 3016 9306
rect 2964 9242 3016 9248
rect 2700 9102 2728 9242
rect 2688 9096 2740 9102
rect 2688 9038 2740 9044
rect 2254 8996 2550 9016
rect 2310 8994 2334 8996
rect 2390 8994 2414 8996
rect 2470 8994 2494 8996
rect 2332 8942 2334 8994
rect 2396 8942 2408 8994
rect 2470 8942 2472 8994
rect 2310 8940 2334 8942
rect 2390 8940 2414 8942
rect 2470 8940 2494 8942
rect 2254 8920 2550 8940
rect 1860 8824 1912 8830
rect 1860 8766 1912 8772
rect 2504 8688 2556 8694
rect 2504 8630 2556 8636
rect 2136 8144 2188 8150
rect 2136 8086 2188 8092
rect 2148 6042 2176 8086
rect 2516 8082 2544 8630
rect 2700 8150 2728 9038
rect 2688 8144 2740 8150
rect 2688 8086 2740 8092
rect 2504 8076 2556 8082
rect 2504 8018 2556 8024
rect 2254 7908 2550 7928
rect 2310 7906 2334 7908
rect 2390 7906 2414 7908
rect 2470 7906 2494 7908
rect 2332 7854 2334 7906
rect 2396 7854 2408 7906
rect 2470 7854 2472 7906
rect 2310 7852 2334 7854
rect 2390 7852 2414 7854
rect 2470 7852 2494 7854
rect 2254 7832 2550 7852
rect 2976 7606 3004 9242
rect 3896 9238 3924 9718
rect 3884 9232 3936 9238
rect 3884 9174 3936 9180
rect 3056 8620 3108 8626
rect 3056 8562 3108 8568
rect 3068 8354 3096 8562
rect 3553 8452 3849 8472
rect 3609 8450 3633 8452
rect 3689 8450 3713 8452
rect 3769 8450 3793 8452
rect 3631 8398 3633 8450
rect 3695 8398 3707 8450
rect 3769 8398 3771 8450
rect 3609 8396 3633 8398
rect 3689 8396 3713 8398
rect 3769 8396 3793 8398
rect 3330 8384 3386 8393
rect 3056 8348 3108 8354
rect 3553 8376 3849 8396
rect 3330 8319 3386 8328
rect 3056 8290 3108 8296
rect 3344 7810 3372 8319
rect 3896 8098 3924 9174
rect 3988 8286 4016 10670
rect 4068 8688 4120 8694
rect 4068 8630 4120 8636
rect 3976 8280 4028 8286
rect 3976 8222 4028 8228
rect 3896 8070 4016 8098
rect 3332 7804 3384 7810
rect 3332 7746 3384 7752
rect 2964 7600 3016 7606
rect 2964 7542 3016 7548
rect 3148 7464 3200 7470
rect 3148 7406 3200 7412
rect 2254 6820 2550 6840
rect 2310 6818 2334 6820
rect 2390 6818 2414 6820
rect 2470 6818 2494 6820
rect 2332 6766 2334 6818
rect 2396 6766 2408 6818
rect 2470 6766 2472 6818
rect 2310 6764 2334 6766
rect 2390 6764 2414 6766
rect 2470 6764 2494 6766
rect 2254 6744 2550 6764
rect 3160 6586 3188 7406
rect 3553 7364 3849 7384
rect 3609 7362 3633 7364
rect 3689 7362 3713 7364
rect 3769 7362 3793 7364
rect 3631 7310 3633 7362
rect 3695 7310 3707 7362
rect 3769 7310 3771 7362
rect 3609 7308 3633 7310
rect 3689 7308 3713 7310
rect 3769 7308 3793 7310
rect 3553 7288 3849 7308
rect 3148 6580 3200 6586
rect 3148 6522 3200 6528
rect 2688 6444 2740 6450
rect 2688 6386 2740 6392
rect 1952 6036 2004 6042
rect 1952 5978 2004 5984
rect 2136 6036 2188 6042
rect 2136 5978 2188 5984
rect 1768 5492 1820 5498
rect 1768 5434 1820 5440
rect 1676 5288 1728 5294
rect 1676 5230 1728 5236
rect 1688 3458 1716 5230
rect 1964 4954 1992 5978
rect 2136 5832 2188 5838
rect 2136 5774 2188 5780
rect 2148 5362 2176 5774
rect 2254 5732 2550 5752
rect 2310 5730 2334 5732
rect 2390 5730 2414 5732
rect 2470 5730 2494 5732
rect 2332 5678 2334 5730
rect 2396 5678 2408 5730
rect 2470 5678 2472 5730
rect 2310 5676 2334 5678
rect 2390 5676 2414 5678
rect 2470 5676 2494 5678
rect 2254 5656 2550 5676
rect 2136 5356 2188 5362
rect 2136 5298 2188 5304
rect 2700 5090 2728 6386
rect 3160 5106 3188 6522
rect 3424 6444 3476 6450
rect 3424 6386 3476 6392
rect 2688 5084 2740 5090
rect 2688 5026 2740 5032
rect 2976 5078 3188 5106
rect 3332 5084 3384 5090
rect 1952 4948 2004 4954
rect 1952 4890 2004 4896
rect 2254 4644 2550 4664
rect 2310 4642 2334 4644
rect 2390 4642 2414 4644
rect 2470 4642 2494 4644
rect 2332 4590 2334 4642
rect 2396 4590 2408 4642
rect 2470 4590 2472 4642
rect 2310 4588 2334 4590
rect 2390 4588 2414 4590
rect 2470 4588 2494 4590
rect 2254 4568 2550 4588
rect 2872 4404 2924 4410
rect 2872 4346 2924 4352
rect 2780 4268 2832 4274
rect 2780 4210 2832 4216
rect 2792 3798 2820 4210
rect 2780 3792 2832 3798
rect 2780 3734 2832 3740
rect 2254 3556 2550 3576
rect 2310 3554 2334 3556
rect 2390 3554 2414 3556
rect 2470 3554 2494 3556
rect 2332 3502 2334 3554
rect 2396 3502 2408 3554
rect 2470 3502 2472 3554
rect 2310 3500 2334 3502
rect 2390 3500 2414 3502
rect 2470 3500 2494 3502
rect 2254 3480 2550 3500
rect 1676 3452 1728 3458
rect 1676 3394 1728 3400
rect 2792 3390 2820 3734
rect 2780 3384 2832 3390
rect 2884 3361 2912 4346
rect 2976 3866 3004 5078
rect 3332 5026 3384 5032
rect 3148 5016 3200 5022
rect 3344 4993 3372 5026
rect 3436 5022 3464 6386
rect 3553 6276 3849 6296
rect 3609 6274 3633 6276
rect 3689 6274 3713 6276
rect 3769 6274 3793 6276
rect 3631 6222 3633 6274
rect 3695 6222 3707 6274
rect 3769 6222 3771 6274
rect 3609 6220 3633 6222
rect 3689 6220 3713 6222
rect 3769 6220 3793 6222
rect 3553 6200 3849 6220
rect 3553 5188 3849 5208
rect 3609 5186 3633 5188
rect 3689 5186 3713 5188
rect 3769 5186 3793 5188
rect 3631 5134 3633 5186
rect 3695 5134 3707 5186
rect 3769 5134 3771 5186
rect 3609 5132 3633 5134
rect 3689 5132 3713 5134
rect 3769 5132 3793 5134
rect 3553 5112 3849 5132
rect 3424 5016 3476 5022
rect 3148 4958 3200 4964
rect 3330 4984 3386 4993
rect 3160 4274 3188 4958
rect 3424 4958 3476 4964
rect 3330 4919 3386 4928
rect 3148 4268 3200 4274
rect 3148 4210 3200 4216
rect 3332 4268 3384 4274
rect 3332 4210 3384 4216
rect 3344 4002 3372 4210
rect 3553 4100 3849 4120
rect 3609 4098 3633 4100
rect 3689 4098 3713 4100
rect 3769 4098 3793 4100
rect 3631 4046 3633 4098
rect 3695 4046 3707 4098
rect 3769 4046 3771 4098
rect 3609 4044 3633 4046
rect 3689 4044 3713 4046
rect 3769 4044 3793 4046
rect 3553 4024 3849 4044
rect 3988 4018 4016 8070
rect 4080 7742 4108 8630
rect 4632 8626 4660 16094
rect 4712 15828 4764 15834
rect 4712 15770 4764 15776
rect 4724 13046 4752 15770
rect 4852 15524 5148 15544
rect 4908 15522 4932 15524
rect 4988 15522 5012 15524
rect 5068 15522 5092 15524
rect 4930 15470 4932 15522
rect 4994 15470 5006 15522
rect 5068 15470 5070 15522
rect 4908 15468 4932 15470
rect 4988 15468 5012 15470
rect 5068 15468 5092 15470
rect 4852 15448 5148 15468
rect 5184 14882 5212 16178
rect 5276 15970 5304 16926
rect 5264 15964 5316 15970
rect 5264 15906 5316 15912
rect 5172 14876 5224 14882
rect 5172 14818 5224 14824
rect 4852 14436 5148 14456
rect 4908 14434 4932 14436
rect 4988 14434 5012 14436
rect 5068 14434 5092 14436
rect 4930 14382 4932 14434
rect 4994 14382 5006 14434
rect 5068 14382 5070 14434
rect 4908 14380 4932 14382
rect 4988 14380 5012 14382
rect 5068 14380 5092 14382
rect 4852 14360 5148 14380
rect 5264 13720 5316 13726
rect 5264 13662 5316 13668
rect 4852 13348 5148 13368
rect 4908 13346 4932 13348
rect 4988 13346 5012 13348
rect 5068 13346 5092 13348
rect 4930 13294 4932 13346
rect 4994 13294 5006 13346
rect 5068 13294 5070 13346
rect 4908 13292 4932 13294
rect 4988 13292 5012 13294
rect 5068 13292 5092 13294
rect 4852 13272 5148 13292
rect 4712 13040 4764 13046
rect 4712 12982 4764 12988
rect 4724 12706 4752 12982
rect 5172 12904 5224 12910
rect 5172 12846 5224 12852
rect 4712 12700 4764 12706
rect 4712 12642 4764 12648
rect 4724 11482 4752 12642
rect 4852 12260 5148 12280
rect 4908 12258 4932 12260
rect 4988 12258 5012 12260
rect 5068 12258 5092 12260
rect 4930 12206 4932 12258
rect 4994 12206 5006 12258
rect 5068 12206 5070 12258
rect 4908 12204 4932 12206
rect 4988 12204 5012 12206
rect 5068 12204 5092 12206
rect 4852 12184 5148 12204
rect 5184 11890 5212 12846
rect 5172 11884 5224 11890
rect 5172 11826 5224 11832
rect 5276 11618 5304 13662
rect 5264 11612 5316 11618
rect 5264 11554 5316 11560
rect 4712 11476 4764 11482
rect 4712 11418 4764 11424
rect 4852 11172 5148 11192
rect 4908 11170 4932 11172
rect 4988 11170 5012 11172
rect 5068 11170 5092 11172
rect 4930 11118 4932 11170
rect 4994 11118 5006 11170
rect 5068 11118 5070 11170
rect 4908 11116 4932 11118
rect 4988 11116 5012 11118
rect 5068 11116 5092 11118
rect 4852 11096 5148 11116
rect 4852 10084 5148 10104
rect 4908 10082 4932 10084
rect 4988 10082 5012 10084
rect 5068 10082 5092 10084
rect 4930 10030 4932 10082
rect 4994 10030 5006 10082
rect 5068 10030 5070 10082
rect 4908 10028 4932 10030
rect 4988 10028 5012 10030
rect 5068 10028 5092 10030
rect 4852 10008 5148 10028
rect 4712 9300 4764 9306
rect 4712 9242 4764 9248
rect 4620 8620 4672 8626
rect 4620 8562 4672 8568
rect 4160 8144 4212 8150
rect 4160 8086 4212 8092
rect 4068 7736 4120 7742
rect 4068 7678 4120 7684
rect 4068 7464 4120 7470
rect 4068 7406 4120 7412
rect 4080 7033 4108 7406
rect 4172 7062 4200 8086
rect 4436 8008 4488 8014
rect 4436 7950 4488 7956
rect 4448 7606 4476 7950
rect 4436 7600 4488 7606
rect 4436 7542 4488 7548
rect 4160 7056 4212 7062
rect 4066 7024 4122 7033
rect 4160 6998 4212 7004
rect 4066 6959 4122 6968
rect 4172 5974 4200 6998
rect 4632 6518 4660 8562
rect 4724 8150 4752 9242
rect 4852 8996 5148 9016
rect 4908 8994 4932 8996
rect 4988 8994 5012 8996
rect 5068 8994 5092 8996
rect 4930 8942 4932 8994
rect 4994 8942 5006 8994
rect 5068 8942 5070 8994
rect 4908 8940 4932 8942
rect 4988 8940 5012 8942
rect 5068 8940 5092 8942
rect 4852 8920 5148 8940
rect 4712 8144 4764 8150
rect 4712 8086 4764 8092
rect 4724 7266 4752 8086
rect 5264 8008 5316 8014
rect 5264 7950 5316 7956
rect 4852 7908 5148 7928
rect 4908 7906 4932 7908
rect 4988 7906 5012 7908
rect 5068 7906 5092 7908
rect 4930 7854 4932 7906
rect 4994 7854 5006 7906
rect 5068 7854 5070 7906
rect 4908 7852 4932 7854
rect 4988 7852 5012 7854
rect 5068 7852 5092 7854
rect 4852 7832 5148 7852
rect 4712 7260 4764 7266
rect 4712 7202 4764 7208
rect 4852 6820 5148 6840
rect 4908 6818 4932 6820
rect 4988 6818 5012 6820
rect 5068 6818 5092 6820
rect 4930 6766 4932 6818
rect 4994 6766 5006 6818
rect 5068 6766 5070 6818
rect 4908 6764 4932 6766
rect 4988 6764 5012 6766
rect 5068 6764 5092 6766
rect 4852 6744 5148 6764
rect 4620 6512 4672 6518
rect 4620 6454 4672 6460
rect 4436 6376 4488 6382
rect 4436 6318 4488 6324
rect 4160 5968 4212 5974
rect 4160 5910 4212 5916
rect 4172 4970 4200 5910
rect 4448 5022 4476 6318
rect 4852 5732 5148 5752
rect 4908 5730 4932 5732
rect 4988 5730 5012 5732
rect 5068 5730 5092 5732
rect 4930 5678 4932 5730
rect 4994 5678 5006 5730
rect 5068 5678 5070 5730
rect 4908 5676 4932 5678
rect 4988 5676 5012 5678
rect 5068 5676 5092 5678
rect 4852 5656 5148 5676
rect 4436 5016 4488 5022
rect 4080 4954 4292 4970
rect 4436 4958 4488 4964
rect 4068 4948 4292 4954
rect 4120 4942 4292 4948
rect 4068 4890 4120 4896
rect 3332 3996 3384 4002
rect 3988 3990 4108 4018
rect 3332 3938 3384 3944
rect 2964 3860 3016 3866
rect 2964 3802 3016 3808
rect 2780 3326 2832 3332
rect 2870 3352 2926 3361
rect 2870 3287 2926 3296
rect 2976 2778 3004 3802
rect 4080 3798 4108 3990
rect 4068 3792 4120 3798
rect 4068 3734 4120 3740
rect 3056 3180 3108 3186
rect 3056 3122 3108 3128
rect 3424 3180 3476 3186
rect 3424 3122 3476 3128
rect 3068 2914 3096 3122
rect 3056 2908 3108 2914
rect 3056 2850 3108 2856
rect 2964 2772 3016 2778
rect 2964 2714 3016 2720
rect 2254 2468 2550 2488
rect 2310 2466 2334 2468
rect 2390 2466 2414 2468
rect 2470 2466 2494 2468
rect 2332 2414 2334 2466
rect 2396 2414 2408 2466
rect 2470 2414 2472 2466
rect 2310 2412 2334 2414
rect 2390 2412 2414 2414
rect 2470 2412 2494 2414
rect 2254 2392 2550 2412
rect 2976 2166 3004 2714
rect 2964 2160 3016 2166
rect 2964 2102 3016 2108
rect 2254 1380 2550 1400
rect 2310 1378 2334 1380
rect 2390 1378 2414 1380
rect 2470 1378 2494 1380
rect 2332 1326 2334 1378
rect 2396 1326 2408 1378
rect 2470 1326 2472 1378
rect 2310 1324 2334 1326
rect 2390 1324 2414 1326
rect 2470 1324 2494 1326
rect 2254 1304 2550 1324
rect 3436 97 3464 3122
rect 3553 3012 3849 3032
rect 3609 3010 3633 3012
rect 3689 3010 3713 3012
rect 3769 3010 3793 3012
rect 3631 2958 3633 3010
rect 3695 2958 3707 3010
rect 3769 2958 3771 3010
rect 3609 2956 3633 2958
rect 3689 2956 3713 2958
rect 3769 2956 3793 2958
rect 3553 2936 3849 2956
rect 4080 2574 4108 3734
rect 4160 3656 4212 3662
rect 4160 3598 4212 3604
rect 4068 2568 4120 2574
rect 4068 2510 4120 2516
rect 3553 1924 3849 1944
rect 3609 1922 3633 1924
rect 3689 1922 3713 1924
rect 3769 1922 3793 1924
rect 3631 1870 3633 1922
rect 3695 1870 3707 1922
rect 3769 1870 3771 1922
rect 3609 1868 3633 1870
rect 3689 1868 3713 1870
rect 3769 1868 3793 1870
rect 3553 1848 3849 1868
rect 4066 1720 4122 1729
rect 4172 1706 4200 3598
rect 4264 3254 4292 4942
rect 4344 4880 4396 4886
rect 4344 4822 4396 4828
rect 4356 3934 4384 4822
rect 4852 4644 5148 4664
rect 4908 4642 4932 4644
rect 4988 4642 5012 4644
rect 5068 4642 5092 4644
rect 4930 4590 4932 4642
rect 4994 4590 5006 4642
rect 5068 4590 5070 4642
rect 4908 4588 4932 4590
rect 4988 4588 5012 4590
rect 5068 4588 5092 4590
rect 4852 4568 5148 4588
rect 4344 3928 4396 3934
rect 4344 3870 4396 3876
rect 4620 3928 4672 3934
rect 4620 3870 4672 3876
rect 4252 3248 4304 3254
rect 4252 3190 4304 3196
rect 4632 2370 4660 3870
rect 4852 3556 5148 3576
rect 4908 3554 4932 3556
rect 4988 3554 5012 3556
rect 5068 3554 5092 3556
rect 4930 3502 4932 3554
rect 4994 3502 5006 3554
rect 5068 3502 5070 3554
rect 4908 3500 4932 3502
rect 4988 3500 5012 3502
rect 5068 3500 5092 3502
rect 4852 3480 5148 3500
rect 5276 3458 5304 7950
rect 5368 4886 5396 18966
rect 5460 14610 5488 19086
rect 5540 19024 5592 19030
rect 5540 18966 5592 18972
rect 5552 18690 5580 18966
rect 5540 18684 5592 18690
rect 5540 18626 5592 18632
rect 5540 15284 5592 15290
rect 5540 15226 5592 15232
rect 5448 14604 5500 14610
rect 5448 14546 5500 14552
rect 5460 12026 5488 14546
rect 5552 13794 5580 15226
rect 5632 15148 5684 15154
rect 5632 15090 5684 15096
rect 5644 14338 5672 15090
rect 5632 14332 5684 14338
rect 5632 14274 5684 14280
rect 5736 14134 5764 20015
rect 5828 15290 5856 22735
rect 6150 21508 6446 21528
rect 6206 21506 6230 21508
rect 6286 21506 6310 21508
rect 6366 21506 6390 21508
rect 6228 21454 6230 21506
rect 6292 21454 6304 21506
rect 6366 21454 6368 21506
rect 6206 21452 6230 21454
rect 6286 21452 6310 21454
rect 6366 21452 6390 21454
rect 6150 21432 6446 21452
rect 7449 20964 7745 20984
rect 7505 20962 7529 20964
rect 7585 20962 7609 20964
rect 7665 20962 7689 20964
rect 7527 20910 7529 20962
rect 7591 20910 7603 20962
rect 7665 20910 7667 20962
rect 7505 20908 7529 20910
rect 7585 20908 7609 20910
rect 7665 20908 7689 20910
rect 7449 20888 7745 20908
rect 6150 20420 6446 20440
rect 6206 20418 6230 20420
rect 6286 20418 6310 20420
rect 6366 20418 6390 20420
rect 6228 20366 6230 20418
rect 6292 20366 6304 20418
rect 6366 20366 6368 20418
rect 6206 20364 6230 20366
rect 6286 20364 6310 20366
rect 6366 20364 6390 20366
rect 6150 20344 6446 20364
rect 7449 19876 7745 19896
rect 7505 19874 7529 19876
rect 7585 19874 7609 19876
rect 7665 19874 7689 19876
rect 7527 19822 7529 19874
rect 7591 19822 7603 19874
rect 7665 19822 7667 19874
rect 7505 19820 7529 19822
rect 7585 19820 7609 19822
rect 7665 19820 7689 19822
rect 7449 19800 7745 19820
rect 6150 19332 6446 19352
rect 6206 19330 6230 19332
rect 6286 19330 6310 19332
rect 6366 19330 6390 19332
rect 6228 19278 6230 19330
rect 6292 19278 6304 19330
rect 6366 19278 6368 19330
rect 6206 19276 6230 19278
rect 6286 19276 6310 19278
rect 6366 19276 6390 19278
rect 6150 19256 6446 19276
rect 7449 18788 7745 18808
rect 7505 18786 7529 18788
rect 7585 18786 7609 18788
rect 7665 18786 7689 18788
rect 7527 18734 7529 18786
rect 7591 18734 7603 18786
rect 7665 18734 7667 18786
rect 7505 18732 7529 18734
rect 7585 18732 7609 18734
rect 7665 18732 7689 18734
rect 7449 18712 7745 18732
rect 6150 18244 6446 18264
rect 6206 18242 6230 18244
rect 6286 18242 6310 18244
rect 6366 18242 6390 18244
rect 6228 18190 6230 18242
rect 6292 18190 6304 18242
rect 6366 18190 6368 18242
rect 6206 18188 6230 18190
rect 6286 18188 6310 18190
rect 6366 18188 6390 18190
rect 6150 18168 6446 18188
rect 7449 17700 7745 17720
rect 7505 17698 7529 17700
rect 7585 17698 7609 17700
rect 7665 17698 7689 17700
rect 7527 17646 7529 17698
rect 7591 17646 7603 17698
rect 7665 17646 7667 17698
rect 7505 17644 7529 17646
rect 7585 17644 7609 17646
rect 7665 17644 7689 17646
rect 7449 17624 7745 17644
rect 6826 17224 6882 17233
rect 6150 17156 6446 17176
rect 6826 17159 6882 17168
rect 6206 17154 6230 17156
rect 6286 17154 6310 17156
rect 6366 17154 6390 17156
rect 6228 17102 6230 17154
rect 6292 17102 6304 17154
rect 6366 17102 6368 17154
rect 6206 17100 6230 17102
rect 6286 17100 6310 17102
rect 6366 17100 6390 17102
rect 6150 17080 6446 17100
rect 6644 16712 6696 16718
rect 6644 16654 6696 16660
rect 6150 16068 6446 16088
rect 6206 16066 6230 16068
rect 6286 16066 6310 16068
rect 6366 16066 6390 16068
rect 6228 16014 6230 16066
rect 6292 16014 6304 16066
rect 6366 16014 6368 16066
rect 6206 16012 6230 16014
rect 6286 16012 6310 16014
rect 6366 16012 6390 16014
rect 6150 15992 6446 16012
rect 5908 15352 5960 15358
rect 5908 15294 5960 15300
rect 5816 15284 5868 15290
rect 5816 15226 5868 15232
rect 5920 15222 5948 15294
rect 5908 15216 5960 15222
rect 5908 15158 5960 15164
rect 5816 15148 5868 15154
rect 5816 15090 5868 15096
rect 5828 14202 5856 15090
rect 5920 14270 5948 15158
rect 6150 14980 6446 15000
rect 6206 14978 6230 14980
rect 6286 14978 6310 14980
rect 6366 14978 6390 14980
rect 6228 14926 6230 14978
rect 6292 14926 6304 14978
rect 6366 14926 6368 14978
rect 6206 14924 6230 14926
rect 6286 14924 6310 14926
rect 6366 14924 6390 14926
rect 6150 14904 6446 14924
rect 5908 14264 5960 14270
rect 5908 14206 5960 14212
rect 6656 14202 6684 16654
rect 6840 15766 6868 17159
rect 7104 16848 7156 16854
rect 7104 16790 7156 16796
rect 7116 15834 7144 16790
rect 7449 16612 7745 16632
rect 7505 16610 7529 16612
rect 7585 16610 7609 16612
rect 7665 16610 7689 16612
rect 7527 16558 7529 16610
rect 7591 16558 7603 16610
rect 7665 16558 7667 16610
rect 7505 16556 7529 16558
rect 7585 16556 7609 16558
rect 7665 16556 7689 16558
rect 7449 16536 7745 16556
rect 7104 15828 7156 15834
rect 7104 15770 7156 15776
rect 7380 15828 7432 15834
rect 7380 15770 7432 15776
rect 6828 15760 6880 15766
rect 6828 15702 6880 15708
rect 7392 14746 7420 15770
rect 7449 15524 7745 15544
rect 7505 15522 7529 15524
rect 7585 15522 7609 15524
rect 7665 15522 7689 15524
rect 7527 15470 7529 15522
rect 7591 15470 7603 15522
rect 7665 15470 7667 15522
rect 7505 15468 7529 15470
rect 7585 15468 7609 15470
rect 7665 15468 7689 15470
rect 7449 15448 7745 15468
rect 7656 15080 7708 15086
rect 7656 15022 7708 15028
rect 7668 14746 7696 15022
rect 7012 14740 7064 14746
rect 7012 14682 7064 14688
rect 7380 14740 7432 14746
rect 7380 14682 7432 14688
rect 7656 14740 7708 14746
rect 7656 14682 7708 14688
rect 6736 14264 6788 14270
rect 6736 14206 6788 14212
rect 5816 14196 5868 14202
rect 5816 14138 5868 14144
rect 6644 14196 6696 14202
rect 6644 14138 6696 14144
rect 5724 14128 5776 14134
rect 5724 14070 5776 14076
rect 6000 14060 6052 14066
rect 6000 14002 6052 14008
rect 5540 13788 5592 13794
rect 5540 13730 5592 13736
rect 5632 13516 5684 13522
rect 5632 13458 5684 13464
rect 5644 13114 5672 13458
rect 5632 13108 5684 13114
rect 5632 13050 5684 13056
rect 5540 12496 5592 12502
rect 5540 12438 5592 12444
rect 5448 12020 5500 12026
rect 5448 11962 5500 11968
rect 5448 8552 5500 8558
rect 5552 8506 5580 12438
rect 5500 8500 5580 8506
rect 5448 8494 5580 8500
rect 5460 8478 5580 8494
rect 5552 8354 5580 8478
rect 5540 8348 5592 8354
rect 5540 8290 5592 8296
rect 5644 7470 5672 13050
rect 6012 12502 6040 14002
rect 6150 13892 6446 13912
rect 6206 13890 6230 13892
rect 6286 13890 6310 13892
rect 6366 13890 6390 13892
rect 6228 13838 6230 13890
rect 6292 13838 6304 13890
rect 6366 13838 6368 13890
rect 6206 13836 6230 13838
rect 6286 13836 6310 13838
rect 6366 13836 6390 13838
rect 6150 13816 6446 13836
rect 6150 12804 6446 12824
rect 6206 12802 6230 12804
rect 6286 12802 6310 12804
rect 6366 12802 6390 12804
rect 6228 12750 6230 12802
rect 6292 12750 6304 12802
rect 6366 12750 6368 12802
rect 6206 12748 6230 12750
rect 6286 12748 6310 12750
rect 6366 12748 6390 12750
rect 6150 12728 6446 12748
rect 6552 12632 6604 12638
rect 6552 12574 6604 12580
rect 6000 12496 6052 12502
rect 6000 12438 6052 12444
rect 5908 11952 5960 11958
rect 5908 11894 5960 11900
rect 5724 8280 5776 8286
rect 5724 8222 5776 8228
rect 5736 7810 5764 8222
rect 5724 7804 5776 7810
rect 5724 7746 5776 7752
rect 5920 7742 5948 11894
rect 6150 11716 6446 11736
rect 6206 11714 6230 11716
rect 6286 11714 6310 11716
rect 6366 11714 6390 11716
rect 6228 11662 6230 11714
rect 6292 11662 6304 11714
rect 6366 11662 6368 11714
rect 6206 11660 6230 11662
rect 6286 11660 6310 11662
rect 6366 11660 6390 11662
rect 6150 11640 6446 11660
rect 6564 11618 6592 12574
rect 6552 11612 6604 11618
rect 6552 11554 6604 11560
rect 6656 11498 6684 14138
rect 6564 11470 6684 11498
rect 6748 11498 6776 14206
rect 6828 13992 6880 13998
rect 6828 13934 6880 13940
rect 6840 13046 6868 13934
rect 7024 13454 7052 14682
rect 7838 14504 7894 14513
rect 7449 14436 7745 14456
rect 7838 14439 7894 14448
rect 7505 14434 7529 14436
rect 7585 14434 7609 14436
rect 7665 14434 7689 14436
rect 7527 14382 7529 14434
rect 7591 14382 7603 14434
rect 7665 14382 7667 14434
rect 7505 14380 7529 14382
rect 7585 14380 7609 14382
rect 7665 14380 7689 14382
rect 7449 14360 7745 14380
rect 7104 14128 7156 14134
rect 7104 14070 7156 14076
rect 7116 13946 7144 14070
rect 7116 13918 7236 13946
rect 7208 13658 7236 13918
rect 7852 13658 7880 14439
rect 7196 13652 7248 13658
rect 7196 13594 7248 13600
rect 7840 13652 7892 13658
rect 7840 13594 7892 13600
rect 7012 13448 7064 13454
rect 7012 13390 7064 13396
rect 7208 13250 7236 13594
rect 7288 13448 7340 13454
rect 7288 13390 7340 13396
rect 7196 13244 7248 13250
rect 7196 13186 7248 13192
rect 6828 13040 6880 13046
rect 6828 12982 6880 12988
rect 6840 11657 6868 12982
rect 7012 12972 7064 12978
rect 7012 12914 7064 12920
rect 7024 12162 7052 12914
rect 7012 12156 7064 12162
rect 7012 12098 7064 12104
rect 6826 11648 6882 11657
rect 6826 11583 6882 11592
rect 6748 11470 6868 11498
rect 6150 10628 6446 10648
rect 6206 10626 6230 10628
rect 6286 10626 6310 10628
rect 6366 10626 6390 10628
rect 6228 10574 6230 10626
rect 6292 10574 6304 10626
rect 6366 10574 6368 10626
rect 6206 10572 6230 10574
rect 6286 10572 6310 10574
rect 6366 10572 6390 10574
rect 6150 10552 6446 10572
rect 6150 9540 6446 9560
rect 6206 9538 6230 9540
rect 6286 9538 6310 9540
rect 6366 9538 6390 9540
rect 6228 9486 6230 9538
rect 6292 9486 6304 9538
rect 6366 9486 6368 9538
rect 6206 9484 6230 9486
rect 6286 9484 6310 9486
rect 6366 9484 6390 9486
rect 6150 9464 6446 9484
rect 6150 8452 6446 8472
rect 6206 8450 6230 8452
rect 6286 8450 6310 8452
rect 6366 8450 6390 8452
rect 6228 8398 6230 8450
rect 6292 8398 6304 8450
rect 6366 8398 6368 8450
rect 6206 8396 6230 8398
rect 6286 8396 6310 8398
rect 6366 8396 6390 8398
rect 6150 8376 6446 8396
rect 5908 7736 5960 7742
rect 5908 7678 5960 7684
rect 5632 7464 5684 7470
rect 5632 7406 5684 7412
rect 6150 7364 6446 7384
rect 6206 7362 6230 7364
rect 6286 7362 6310 7364
rect 6366 7362 6390 7364
rect 6228 7310 6230 7362
rect 6292 7310 6304 7362
rect 6366 7310 6368 7362
rect 6206 7308 6230 7310
rect 6286 7308 6310 7310
rect 6366 7308 6390 7310
rect 6150 7288 6446 7308
rect 5724 7124 5776 7130
rect 5724 7066 5776 7072
rect 5632 7056 5684 7062
rect 5632 6998 5684 7004
rect 5644 6081 5672 6998
rect 5736 6722 5764 7066
rect 5724 6716 5776 6722
rect 5724 6658 5776 6664
rect 6150 6276 6446 6296
rect 6206 6274 6230 6276
rect 6286 6274 6310 6276
rect 6366 6274 6390 6276
rect 6228 6222 6230 6274
rect 6292 6222 6304 6274
rect 6366 6222 6368 6274
rect 6206 6220 6230 6222
rect 6286 6220 6310 6222
rect 6366 6220 6390 6222
rect 6150 6200 6446 6220
rect 5630 6072 5686 6081
rect 5630 6007 5686 6016
rect 6150 5188 6446 5208
rect 6206 5186 6230 5188
rect 6286 5186 6310 5188
rect 6366 5186 6390 5188
rect 6228 5134 6230 5186
rect 6292 5134 6304 5186
rect 6366 5134 6368 5186
rect 6206 5132 6230 5134
rect 6286 5132 6310 5134
rect 6366 5132 6390 5134
rect 6150 5112 6446 5132
rect 6564 5090 6592 11470
rect 6644 10796 6696 10802
rect 6644 10738 6696 10744
rect 6552 5084 6604 5090
rect 6552 5026 6604 5032
rect 5356 4880 5408 4886
rect 5356 4822 5408 4828
rect 6150 4100 6446 4120
rect 6206 4098 6230 4100
rect 6286 4098 6310 4100
rect 6366 4098 6390 4100
rect 6228 4046 6230 4098
rect 6292 4046 6304 4098
rect 6366 4046 6368 4098
rect 6206 4044 6230 4046
rect 6286 4044 6310 4046
rect 6366 4044 6390 4046
rect 6150 4024 6446 4044
rect 5264 3452 5316 3458
rect 5264 3394 5316 3400
rect 6656 3361 6684 10738
rect 6840 9782 6868 11470
rect 7300 9782 7328 13390
rect 7449 13348 7745 13368
rect 7505 13346 7529 13348
rect 7585 13346 7609 13348
rect 7665 13346 7689 13348
rect 7527 13294 7529 13346
rect 7591 13294 7603 13346
rect 7665 13294 7667 13346
rect 7505 13292 7529 13294
rect 7585 13292 7609 13294
rect 7665 13292 7689 13294
rect 7449 13272 7745 13292
rect 7449 12260 7745 12280
rect 7505 12258 7529 12260
rect 7585 12258 7609 12260
rect 7665 12258 7689 12260
rect 7527 12206 7529 12258
rect 7591 12206 7603 12258
rect 7665 12206 7667 12258
rect 7505 12204 7529 12206
rect 7585 12204 7609 12206
rect 7665 12204 7689 12206
rect 7449 12184 7745 12204
rect 7449 11172 7745 11192
rect 7505 11170 7529 11172
rect 7585 11170 7609 11172
rect 7665 11170 7689 11172
rect 7527 11118 7529 11170
rect 7591 11118 7603 11170
rect 7665 11118 7667 11170
rect 7505 11116 7529 11118
rect 7585 11116 7609 11118
rect 7665 11116 7689 11118
rect 7449 11096 7745 11116
rect 7449 10084 7745 10104
rect 7505 10082 7529 10084
rect 7585 10082 7609 10084
rect 7665 10082 7689 10084
rect 7527 10030 7529 10082
rect 7591 10030 7603 10082
rect 7665 10030 7667 10082
rect 7505 10028 7529 10030
rect 7585 10028 7609 10030
rect 7665 10028 7689 10030
rect 7449 10008 7745 10028
rect 6828 9776 6880 9782
rect 6828 9718 6880 9724
rect 7288 9776 7340 9782
rect 7288 9718 7340 9724
rect 6840 9238 6868 9718
rect 8208 9708 8260 9714
rect 8208 9650 8260 9656
rect 7012 9368 7064 9374
rect 7012 9310 7064 9316
rect 6828 9232 6880 9238
rect 6828 9174 6880 9180
rect 7024 8898 7052 9310
rect 7449 8996 7745 9016
rect 7505 8994 7529 8996
rect 7585 8994 7609 8996
rect 7665 8994 7689 8996
rect 7527 8942 7529 8994
rect 7591 8942 7603 8994
rect 7665 8942 7667 8994
rect 7505 8940 7529 8942
rect 7585 8940 7609 8942
rect 7665 8940 7689 8942
rect 7449 8920 7745 8940
rect 8220 8937 8248 9650
rect 8206 8928 8262 8937
rect 7012 8892 7064 8898
rect 8206 8863 8262 8872
rect 7012 8834 7064 8840
rect 7472 8688 7524 8694
rect 7472 8630 7524 8636
rect 7484 8354 7512 8630
rect 7472 8348 7524 8354
rect 7472 8290 7524 8296
rect 7449 7908 7745 7928
rect 7505 7906 7529 7908
rect 7585 7906 7609 7908
rect 7665 7906 7689 7908
rect 7527 7854 7529 7906
rect 7591 7854 7603 7906
rect 7665 7854 7667 7906
rect 7505 7852 7529 7854
rect 7585 7852 7609 7854
rect 7665 7852 7689 7854
rect 7449 7832 7745 7852
rect 7449 6820 7745 6840
rect 7505 6818 7529 6820
rect 7585 6818 7609 6820
rect 7665 6818 7689 6820
rect 7527 6766 7529 6818
rect 7591 6766 7603 6818
rect 7665 6766 7667 6818
rect 7505 6764 7529 6766
rect 7585 6764 7609 6766
rect 7665 6764 7689 6766
rect 7449 6744 7745 6764
rect 7449 5732 7745 5752
rect 7505 5730 7529 5732
rect 7585 5730 7609 5732
rect 7665 5730 7689 5732
rect 7527 5678 7529 5730
rect 7591 5678 7603 5730
rect 7665 5678 7667 5730
rect 7505 5676 7529 5678
rect 7585 5676 7609 5678
rect 7665 5676 7689 5678
rect 7449 5656 7745 5676
rect 7449 4644 7745 4664
rect 7505 4642 7529 4644
rect 7585 4642 7609 4644
rect 7665 4642 7689 4644
rect 7527 4590 7529 4642
rect 7591 4590 7603 4642
rect 7665 4590 7667 4642
rect 7505 4588 7529 4590
rect 7585 4588 7609 4590
rect 7665 4588 7689 4590
rect 7449 4568 7745 4588
rect 7449 3556 7745 3576
rect 7505 3554 7529 3556
rect 7585 3554 7609 3556
rect 7665 3554 7689 3556
rect 7527 3502 7529 3554
rect 7591 3502 7603 3554
rect 7665 3502 7667 3554
rect 7505 3500 7529 3502
rect 7585 3500 7609 3502
rect 7665 3500 7689 3502
rect 7449 3480 7745 3500
rect 6642 3352 6698 3361
rect 6642 3287 6698 3296
rect 4896 3248 4948 3254
rect 4896 3190 4948 3196
rect 6828 3248 6880 3254
rect 6828 3190 6880 3196
rect 4908 2778 4936 3190
rect 6150 3012 6446 3032
rect 6206 3010 6230 3012
rect 6286 3010 6310 3012
rect 6366 3010 6390 3012
rect 6228 2958 6230 3010
rect 6292 2958 6304 3010
rect 6366 2958 6368 3010
rect 6206 2956 6230 2958
rect 6286 2956 6310 2958
rect 6366 2956 6390 2958
rect 6150 2936 6446 2956
rect 4896 2772 4948 2778
rect 4896 2714 4948 2720
rect 4852 2468 5148 2488
rect 4908 2466 4932 2468
rect 4988 2466 5012 2468
rect 5068 2466 5092 2468
rect 4930 2414 4932 2466
rect 4994 2414 5006 2466
rect 5068 2414 5070 2466
rect 4908 2412 4932 2414
rect 4988 2412 5012 2414
rect 5068 2412 5092 2414
rect 4852 2392 5148 2412
rect 4620 2364 4672 2370
rect 4620 2306 4672 2312
rect 6150 1924 6446 1944
rect 6206 1922 6230 1924
rect 6286 1922 6310 1924
rect 6366 1922 6390 1924
rect 6228 1870 6230 1922
rect 6292 1870 6304 1922
rect 6366 1870 6368 1922
rect 6206 1868 6230 1870
rect 6286 1868 6310 1870
rect 6366 1868 6390 1870
rect 6150 1848 6446 1868
rect 4122 1678 4200 1706
rect 4066 1655 4122 1664
rect 4852 1380 5148 1400
rect 4908 1378 4932 1380
rect 4988 1378 5012 1380
rect 5068 1378 5092 1380
rect 4930 1326 4932 1378
rect 4994 1326 5006 1378
rect 5068 1326 5070 1378
rect 4908 1324 4932 1326
rect 4988 1324 5012 1326
rect 5068 1324 5092 1326
rect 4852 1304 5148 1324
rect 6840 641 6868 3190
rect 6920 3112 6972 3118
rect 6920 3054 6972 3060
rect 6932 2778 6960 3054
rect 6920 2772 6972 2778
rect 6920 2714 6972 2720
rect 7449 2468 7745 2488
rect 7505 2466 7529 2468
rect 7585 2466 7609 2468
rect 7665 2466 7689 2468
rect 7527 2414 7529 2466
rect 7591 2414 7603 2466
rect 7665 2414 7667 2466
rect 7505 2412 7529 2414
rect 7585 2412 7609 2414
rect 7665 2412 7689 2414
rect 7449 2392 7745 2412
rect 7449 1380 7745 1400
rect 7505 1378 7529 1380
rect 7585 1378 7609 1380
rect 7665 1378 7689 1380
rect 7527 1326 7529 1378
rect 7591 1326 7603 1378
rect 7665 1326 7667 1378
rect 7505 1324 7529 1326
rect 7585 1324 7609 1326
rect 7665 1324 7689 1326
rect 7449 1304 7745 1324
rect 6826 632 6882 641
rect 6826 567 6882 576
rect 3422 88 3478 97
rect 3422 23 3478 32
<< via2 >>
rect 4066 23288 4122 23344
rect 5814 22744 5870 22800
rect 3422 21656 3478 21712
rect 2254 20962 2310 20964
rect 2334 20962 2390 20964
rect 2414 20962 2470 20964
rect 2494 20962 2550 20964
rect 2254 20910 2280 20962
rect 2280 20910 2310 20962
rect 2334 20910 2344 20962
rect 2344 20910 2390 20962
rect 2414 20910 2460 20962
rect 2460 20910 2470 20962
rect 2494 20910 2524 20962
rect 2524 20910 2550 20962
rect 2254 20908 2310 20910
rect 2334 20908 2390 20910
rect 2414 20908 2470 20910
rect 2494 20908 2550 20910
rect 3054 20024 3110 20080
rect 2254 19874 2310 19876
rect 2334 19874 2390 19876
rect 2414 19874 2470 19876
rect 2494 19874 2550 19876
rect 2254 19822 2280 19874
rect 2280 19822 2310 19874
rect 2334 19822 2344 19874
rect 2344 19822 2390 19874
rect 2414 19822 2460 19874
rect 2460 19822 2470 19874
rect 2494 19822 2524 19874
rect 2524 19822 2550 19874
rect 2254 19820 2310 19822
rect 2334 19820 2390 19822
rect 2414 19820 2470 19822
rect 2494 19820 2550 19822
rect 2254 18786 2310 18788
rect 2334 18786 2390 18788
rect 2414 18786 2470 18788
rect 2494 18786 2550 18788
rect 2254 18734 2280 18786
rect 2280 18734 2310 18786
rect 2334 18734 2344 18786
rect 2344 18734 2390 18786
rect 2414 18734 2460 18786
rect 2460 18734 2470 18786
rect 2494 18734 2524 18786
rect 2524 18734 2550 18786
rect 2254 18732 2310 18734
rect 2334 18732 2390 18734
rect 2414 18732 2470 18734
rect 2494 18732 2550 18734
rect 3553 21506 3609 21508
rect 3633 21506 3689 21508
rect 3713 21506 3769 21508
rect 3793 21506 3849 21508
rect 3553 21454 3579 21506
rect 3579 21454 3609 21506
rect 3633 21454 3643 21506
rect 3643 21454 3689 21506
rect 3713 21454 3759 21506
rect 3759 21454 3769 21506
rect 3793 21454 3823 21506
rect 3823 21454 3849 21506
rect 3553 21452 3609 21454
rect 3633 21452 3689 21454
rect 3713 21452 3769 21454
rect 3793 21452 3849 21454
rect 4852 20962 4908 20964
rect 4932 20962 4988 20964
rect 5012 20962 5068 20964
rect 5092 20962 5148 20964
rect 4852 20910 4878 20962
rect 4878 20910 4908 20962
rect 4932 20910 4942 20962
rect 4942 20910 4988 20962
rect 5012 20910 5058 20962
rect 5058 20910 5068 20962
rect 5092 20910 5122 20962
rect 5122 20910 5148 20962
rect 4852 20908 4908 20910
rect 4932 20908 4988 20910
rect 5012 20908 5068 20910
rect 5092 20908 5148 20910
rect 3553 20418 3609 20420
rect 3633 20418 3689 20420
rect 3713 20418 3769 20420
rect 3793 20418 3849 20420
rect 3553 20366 3579 20418
rect 3579 20366 3609 20418
rect 3633 20366 3643 20418
rect 3643 20366 3689 20418
rect 3713 20366 3759 20418
rect 3759 20366 3769 20418
rect 3793 20366 3823 20418
rect 3823 20366 3849 20418
rect 3553 20364 3609 20366
rect 3633 20364 3689 20366
rect 3713 20364 3769 20366
rect 3793 20364 3849 20366
rect 4852 19874 4908 19876
rect 4932 19874 4988 19876
rect 5012 19874 5068 19876
rect 5092 19874 5148 19876
rect 4852 19822 4878 19874
rect 4878 19822 4908 19874
rect 4932 19822 4942 19874
rect 4942 19822 4988 19874
rect 5012 19822 5058 19874
rect 5058 19822 5068 19874
rect 5092 19822 5122 19874
rect 5122 19822 5148 19874
rect 4852 19820 4908 19822
rect 4932 19820 4988 19822
rect 5012 19820 5068 19822
rect 5092 19820 5148 19822
rect 3238 18256 3294 18312
rect 2254 17698 2310 17700
rect 2334 17698 2390 17700
rect 2414 17698 2470 17700
rect 2494 17698 2550 17700
rect 2254 17646 2280 17698
rect 2280 17646 2310 17698
rect 2334 17646 2344 17698
rect 2344 17646 2390 17698
rect 2414 17646 2460 17698
rect 2460 17646 2470 17698
rect 2494 17646 2524 17698
rect 2524 17646 2550 17698
rect 2254 17644 2310 17646
rect 2334 17644 2390 17646
rect 2414 17644 2470 17646
rect 2494 17644 2550 17646
rect 2254 16610 2310 16612
rect 2334 16610 2390 16612
rect 2414 16610 2470 16612
rect 2494 16610 2550 16612
rect 2254 16558 2280 16610
rect 2280 16558 2310 16610
rect 2334 16558 2344 16610
rect 2344 16558 2390 16610
rect 2414 16558 2460 16610
rect 2460 16558 2470 16610
rect 2494 16558 2524 16610
rect 2524 16558 2550 16610
rect 2254 16556 2310 16558
rect 2334 16556 2390 16558
rect 2414 16556 2470 16558
rect 2494 16556 2550 16558
rect 2254 15522 2310 15524
rect 2334 15522 2390 15524
rect 2414 15522 2470 15524
rect 2494 15522 2550 15524
rect 2254 15470 2280 15522
rect 2280 15470 2310 15522
rect 2334 15470 2344 15522
rect 2344 15470 2390 15522
rect 2414 15470 2460 15522
rect 2460 15470 2470 15522
rect 2494 15470 2524 15522
rect 2524 15470 2550 15522
rect 2254 15468 2310 15470
rect 2334 15468 2390 15470
rect 2414 15468 2470 15470
rect 2494 15468 2550 15470
rect 2254 14434 2310 14436
rect 2334 14434 2390 14436
rect 2414 14434 2470 14436
rect 2494 14434 2550 14436
rect 2254 14382 2280 14434
rect 2280 14382 2310 14434
rect 2334 14382 2344 14434
rect 2344 14382 2390 14434
rect 2414 14382 2460 14434
rect 2460 14382 2470 14434
rect 2494 14382 2524 14434
rect 2524 14382 2550 14434
rect 2254 14380 2310 14382
rect 2334 14380 2390 14382
rect 2414 14380 2470 14382
rect 2494 14380 2550 14382
rect 2254 13346 2310 13348
rect 2334 13346 2390 13348
rect 2414 13346 2470 13348
rect 2494 13346 2550 13348
rect 2254 13294 2280 13346
rect 2280 13294 2310 13346
rect 2334 13294 2344 13346
rect 2344 13294 2390 13346
rect 2414 13294 2460 13346
rect 2460 13294 2470 13346
rect 2494 13294 2524 13346
rect 2524 13294 2550 13346
rect 2254 13292 2310 13294
rect 2334 13292 2390 13294
rect 2414 13292 2470 13294
rect 2494 13292 2550 13294
rect 2254 12258 2310 12260
rect 2334 12258 2390 12260
rect 2414 12258 2470 12260
rect 2494 12258 2550 12260
rect 2254 12206 2280 12258
rect 2280 12206 2310 12258
rect 2334 12206 2344 12258
rect 2344 12206 2390 12258
rect 2414 12206 2460 12258
rect 2460 12206 2470 12258
rect 2494 12206 2524 12258
rect 2524 12206 2550 12258
rect 2254 12204 2310 12206
rect 2334 12204 2390 12206
rect 2414 12204 2470 12206
rect 2494 12204 2550 12206
rect 3054 14992 3110 15048
rect 2254 11170 2310 11172
rect 2334 11170 2390 11172
rect 2414 11170 2470 11172
rect 2494 11170 2550 11172
rect 2254 11118 2280 11170
rect 2280 11118 2310 11170
rect 2334 11118 2344 11170
rect 2344 11118 2390 11170
rect 2414 11118 2460 11170
rect 2460 11118 2470 11170
rect 2494 11118 2524 11170
rect 2524 11118 2550 11170
rect 2254 11116 2310 11118
rect 2334 11116 2390 11118
rect 2414 11116 2470 11118
rect 2494 11116 2550 11118
rect 3553 19330 3609 19332
rect 3633 19330 3689 19332
rect 3713 19330 3769 19332
rect 3793 19330 3849 19332
rect 3553 19278 3579 19330
rect 3579 19278 3609 19330
rect 3633 19278 3643 19330
rect 3643 19278 3689 19330
rect 3713 19278 3759 19330
rect 3759 19278 3769 19330
rect 3793 19278 3823 19330
rect 3823 19278 3849 19330
rect 3553 19276 3609 19278
rect 3633 19276 3689 19278
rect 3713 19276 3769 19278
rect 3793 19276 3849 19278
rect 5722 20024 5778 20080
rect 3553 18242 3609 18244
rect 3633 18242 3689 18244
rect 3713 18242 3769 18244
rect 3793 18242 3849 18244
rect 3553 18190 3579 18242
rect 3579 18190 3609 18242
rect 3633 18190 3643 18242
rect 3643 18190 3689 18242
rect 3713 18190 3759 18242
rect 3759 18190 3769 18242
rect 3793 18190 3823 18242
rect 3823 18190 3849 18242
rect 3553 18188 3609 18190
rect 3633 18188 3689 18190
rect 3713 18188 3769 18190
rect 3793 18188 3849 18190
rect 4852 18786 4908 18788
rect 4932 18786 4988 18788
rect 5012 18786 5068 18788
rect 5092 18786 5148 18788
rect 4852 18734 4878 18786
rect 4878 18734 4908 18786
rect 4932 18734 4942 18786
rect 4942 18734 4988 18786
rect 5012 18734 5058 18786
rect 5058 18734 5068 18786
rect 5092 18734 5122 18786
rect 5122 18734 5148 18786
rect 4852 18732 4908 18734
rect 4932 18732 4988 18734
rect 5012 18732 5068 18734
rect 5092 18732 5148 18734
rect 3553 17154 3609 17156
rect 3633 17154 3689 17156
rect 3713 17154 3769 17156
rect 3793 17154 3849 17156
rect 3553 17102 3579 17154
rect 3579 17102 3609 17154
rect 3633 17102 3643 17154
rect 3643 17102 3689 17154
rect 3713 17102 3759 17154
rect 3759 17102 3769 17154
rect 3793 17102 3823 17154
rect 3823 17102 3849 17154
rect 3553 17100 3609 17102
rect 3633 17100 3689 17102
rect 3713 17100 3769 17102
rect 3793 17100 3849 17102
rect 4066 16352 4122 16408
rect 3553 16066 3609 16068
rect 3633 16066 3689 16068
rect 3713 16066 3769 16068
rect 3793 16066 3849 16068
rect 3553 16014 3579 16066
rect 3579 16014 3609 16066
rect 3633 16014 3643 16066
rect 3643 16014 3689 16066
rect 3713 16014 3759 16066
rect 3759 16014 3769 16066
rect 3793 16014 3823 16066
rect 3823 16014 3849 16066
rect 3553 16012 3609 16014
rect 3633 16012 3689 16014
rect 3713 16012 3769 16014
rect 3793 16012 3849 16014
rect 4852 17698 4908 17700
rect 4932 17698 4988 17700
rect 5012 17698 5068 17700
rect 5092 17698 5148 17700
rect 4852 17646 4878 17698
rect 4878 17646 4908 17698
rect 4932 17646 4942 17698
rect 4942 17646 4988 17698
rect 5012 17646 5058 17698
rect 5058 17646 5068 17698
rect 5092 17646 5122 17698
rect 5122 17646 5148 17698
rect 4852 17644 4908 17646
rect 4932 17644 4988 17646
rect 5012 17644 5068 17646
rect 5092 17644 5148 17646
rect 4852 16610 4908 16612
rect 4932 16610 4988 16612
rect 5012 16610 5068 16612
rect 5092 16610 5148 16612
rect 4852 16558 4878 16610
rect 4878 16558 4908 16610
rect 4932 16558 4942 16610
rect 4942 16558 4988 16610
rect 5012 16558 5058 16610
rect 5058 16558 5068 16610
rect 5092 16558 5122 16610
rect 5122 16558 5148 16610
rect 4852 16556 4908 16558
rect 4932 16556 4988 16558
rect 5012 16556 5068 16558
rect 5092 16556 5148 16558
rect 3553 14978 3609 14980
rect 3633 14978 3689 14980
rect 3713 14978 3769 14980
rect 3793 14978 3849 14980
rect 3553 14926 3579 14978
rect 3579 14926 3609 14978
rect 3633 14926 3643 14978
rect 3643 14926 3689 14978
rect 3713 14926 3759 14978
rect 3759 14926 3769 14978
rect 3793 14926 3823 14978
rect 3823 14926 3849 14978
rect 3553 14924 3609 14926
rect 3633 14924 3689 14926
rect 3713 14924 3769 14926
rect 3793 14924 3849 14926
rect 3553 13890 3609 13892
rect 3633 13890 3689 13892
rect 3713 13890 3769 13892
rect 3793 13890 3849 13892
rect 3553 13838 3579 13890
rect 3579 13838 3609 13890
rect 3633 13838 3643 13890
rect 3643 13838 3689 13890
rect 3713 13838 3759 13890
rect 3759 13838 3769 13890
rect 3793 13838 3823 13890
rect 3823 13838 3849 13890
rect 3553 13836 3609 13838
rect 3633 13836 3689 13838
rect 3713 13836 3769 13838
rect 3793 13836 3849 13838
rect 2254 10082 2310 10084
rect 2334 10082 2390 10084
rect 2414 10082 2470 10084
rect 2494 10082 2550 10084
rect 2254 10030 2280 10082
rect 2280 10030 2310 10082
rect 2334 10030 2344 10082
rect 2344 10030 2390 10082
rect 2414 10030 2460 10082
rect 2460 10030 2470 10082
rect 2494 10030 2524 10082
rect 2524 10030 2550 10082
rect 2254 10028 2310 10030
rect 2334 10028 2390 10030
rect 2414 10028 2470 10030
rect 2494 10028 2550 10030
rect 3553 12802 3609 12804
rect 3633 12802 3689 12804
rect 3713 12802 3769 12804
rect 3793 12802 3849 12804
rect 3553 12750 3579 12802
rect 3579 12750 3609 12802
rect 3633 12750 3643 12802
rect 3643 12750 3689 12802
rect 3713 12750 3759 12802
rect 3759 12750 3769 12802
rect 3793 12750 3823 12802
rect 3823 12750 3849 12802
rect 3553 12748 3609 12750
rect 3633 12748 3689 12750
rect 3713 12748 3769 12750
rect 3793 12748 3849 12750
rect 3553 11714 3609 11716
rect 3633 11714 3689 11716
rect 3713 11714 3769 11716
rect 3793 11714 3849 11716
rect 3553 11662 3579 11714
rect 3579 11662 3609 11714
rect 3633 11662 3643 11714
rect 3643 11662 3689 11714
rect 3713 11662 3759 11714
rect 3759 11662 3769 11714
rect 3793 11662 3823 11714
rect 3823 11662 3849 11714
rect 3553 11660 3609 11662
rect 3633 11660 3689 11662
rect 3713 11660 3769 11662
rect 3793 11660 3849 11662
rect 3238 11592 3294 11648
rect 3553 10626 3609 10628
rect 3633 10626 3689 10628
rect 3713 10626 3769 10628
rect 3793 10626 3849 10628
rect 3553 10574 3579 10626
rect 3579 10574 3609 10626
rect 3633 10574 3643 10626
rect 3643 10574 3689 10626
rect 3713 10574 3759 10626
rect 3759 10574 3769 10626
rect 3793 10574 3823 10626
rect 3823 10574 3849 10626
rect 3553 10572 3609 10574
rect 3633 10572 3689 10574
rect 3713 10572 3769 10574
rect 3793 10572 3849 10574
rect 3422 9844 3478 9880
rect 3422 9824 3424 9844
rect 3424 9824 3476 9844
rect 3476 9824 3478 9844
rect 4066 13496 4122 13552
rect 3553 9538 3609 9540
rect 3633 9538 3689 9540
rect 3713 9538 3769 9540
rect 3793 9538 3849 9540
rect 3553 9486 3579 9538
rect 3579 9486 3609 9538
rect 3633 9486 3643 9538
rect 3643 9486 3689 9538
rect 3713 9486 3759 9538
rect 3759 9486 3769 9538
rect 3793 9486 3823 9538
rect 3823 9486 3849 9538
rect 3553 9484 3609 9486
rect 3633 9484 3689 9486
rect 3713 9484 3769 9486
rect 3793 9484 3849 9486
rect 2254 8994 2310 8996
rect 2334 8994 2390 8996
rect 2414 8994 2470 8996
rect 2494 8994 2550 8996
rect 2254 8942 2280 8994
rect 2280 8942 2310 8994
rect 2334 8942 2344 8994
rect 2344 8942 2390 8994
rect 2414 8942 2460 8994
rect 2460 8942 2470 8994
rect 2494 8942 2524 8994
rect 2524 8942 2550 8994
rect 2254 8940 2310 8942
rect 2334 8940 2390 8942
rect 2414 8940 2470 8942
rect 2494 8940 2550 8942
rect 2254 7906 2310 7908
rect 2334 7906 2390 7908
rect 2414 7906 2470 7908
rect 2494 7906 2550 7908
rect 2254 7854 2280 7906
rect 2280 7854 2310 7906
rect 2334 7854 2344 7906
rect 2344 7854 2390 7906
rect 2414 7854 2460 7906
rect 2460 7854 2470 7906
rect 2494 7854 2524 7906
rect 2524 7854 2550 7906
rect 2254 7852 2310 7854
rect 2334 7852 2390 7854
rect 2414 7852 2470 7854
rect 2494 7852 2550 7854
rect 3553 8450 3609 8452
rect 3633 8450 3689 8452
rect 3713 8450 3769 8452
rect 3793 8450 3849 8452
rect 3553 8398 3579 8450
rect 3579 8398 3609 8450
rect 3633 8398 3643 8450
rect 3643 8398 3689 8450
rect 3713 8398 3759 8450
rect 3759 8398 3769 8450
rect 3793 8398 3823 8450
rect 3823 8398 3849 8450
rect 3553 8396 3609 8398
rect 3633 8396 3689 8398
rect 3713 8396 3769 8398
rect 3793 8396 3849 8398
rect 3330 8328 3386 8384
rect 2254 6818 2310 6820
rect 2334 6818 2390 6820
rect 2414 6818 2470 6820
rect 2494 6818 2550 6820
rect 2254 6766 2280 6818
rect 2280 6766 2310 6818
rect 2334 6766 2344 6818
rect 2344 6766 2390 6818
rect 2414 6766 2460 6818
rect 2460 6766 2470 6818
rect 2494 6766 2524 6818
rect 2524 6766 2550 6818
rect 2254 6764 2310 6766
rect 2334 6764 2390 6766
rect 2414 6764 2470 6766
rect 2494 6764 2550 6766
rect 3553 7362 3609 7364
rect 3633 7362 3689 7364
rect 3713 7362 3769 7364
rect 3793 7362 3849 7364
rect 3553 7310 3579 7362
rect 3579 7310 3609 7362
rect 3633 7310 3643 7362
rect 3643 7310 3689 7362
rect 3713 7310 3759 7362
rect 3759 7310 3769 7362
rect 3793 7310 3823 7362
rect 3823 7310 3849 7362
rect 3553 7308 3609 7310
rect 3633 7308 3689 7310
rect 3713 7308 3769 7310
rect 3793 7308 3849 7310
rect 2254 5730 2310 5732
rect 2334 5730 2390 5732
rect 2414 5730 2470 5732
rect 2494 5730 2550 5732
rect 2254 5678 2280 5730
rect 2280 5678 2310 5730
rect 2334 5678 2344 5730
rect 2344 5678 2390 5730
rect 2414 5678 2460 5730
rect 2460 5678 2470 5730
rect 2494 5678 2524 5730
rect 2524 5678 2550 5730
rect 2254 5676 2310 5678
rect 2334 5676 2390 5678
rect 2414 5676 2470 5678
rect 2494 5676 2550 5678
rect 2254 4642 2310 4644
rect 2334 4642 2390 4644
rect 2414 4642 2470 4644
rect 2494 4642 2550 4644
rect 2254 4590 2280 4642
rect 2280 4590 2310 4642
rect 2334 4590 2344 4642
rect 2344 4590 2390 4642
rect 2414 4590 2460 4642
rect 2460 4590 2470 4642
rect 2494 4590 2524 4642
rect 2524 4590 2550 4642
rect 2254 4588 2310 4590
rect 2334 4588 2390 4590
rect 2414 4588 2470 4590
rect 2494 4588 2550 4590
rect 2254 3554 2310 3556
rect 2334 3554 2390 3556
rect 2414 3554 2470 3556
rect 2494 3554 2550 3556
rect 2254 3502 2280 3554
rect 2280 3502 2310 3554
rect 2334 3502 2344 3554
rect 2344 3502 2390 3554
rect 2414 3502 2460 3554
rect 2460 3502 2470 3554
rect 2494 3502 2524 3554
rect 2524 3502 2550 3554
rect 2254 3500 2310 3502
rect 2334 3500 2390 3502
rect 2414 3500 2470 3502
rect 2494 3500 2550 3502
rect 3553 6274 3609 6276
rect 3633 6274 3689 6276
rect 3713 6274 3769 6276
rect 3793 6274 3849 6276
rect 3553 6222 3579 6274
rect 3579 6222 3609 6274
rect 3633 6222 3643 6274
rect 3643 6222 3689 6274
rect 3713 6222 3759 6274
rect 3759 6222 3769 6274
rect 3793 6222 3823 6274
rect 3823 6222 3849 6274
rect 3553 6220 3609 6222
rect 3633 6220 3689 6222
rect 3713 6220 3769 6222
rect 3793 6220 3849 6222
rect 3553 5186 3609 5188
rect 3633 5186 3689 5188
rect 3713 5186 3769 5188
rect 3793 5186 3849 5188
rect 3553 5134 3579 5186
rect 3579 5134 3609 5186
rect 3633 5134 3643 5186
rect 3643 5134 3689 5186
rect 3713 5134 3759 5186
rect 3759 5134 3769 5186
rect 3793 5134 3823 5186
rect 3823 5134 3849 5186
rect 3553 5132 3609 5134
rect 3633 5132 3689 5134
rect 3713 5132 3769 5134
rect 3793 5132 3849 5134
rect 3330 4928 3386 4984
rect 3553 4098 3609 4100
rect 3633 4098 3689 4100
rect 3713 4098 3769 4100
rect 3793 4098 3849 4100
rect 3553 4046 3579 4098
rect 3579 4046 3609 4098
rect 3633 4046 3643 4098
rect 3643 4046 3689 4098
rect 3713 4046 3759 4098
rect 3759 4046 3769 4098
rect 3793 4046 3823 4098
rect 3823 4046 3849 4098
rect 3553 4044 3609 4046
rect 3633 4044 3689 4046
rect 3713 4044 3769 4046
rect 3793 4044 3849 4046
rect 4852 15522 4908 15524
rect 4932 15522 4988 15524
rect 5012 15522 5068 15524
rect 5092 15522 5148 15524
rect 4852 15470 4878 15522
rect 4878 15470 4908 15522
rect 4932 15470 4942 15522
rect 4942 15470 4988 15522
rect 5012 15470 5058 15522
rect 5058 15470 5068 15522
rect 5092 15470 5122 15522
rect 5122 15470 5148 15522
rect 4852 15468 4908 15470
rect 4932 15468 4988 15470
rect 5012 15468 5068 15470
rect 5092 15468 5148 15470
rect 4852 14434 4908 14436
rect 4932 14434 4988 14436
rect 5012 14434 5068 14436
rect 5092 14434 5148 14436
rect 4852 14382 4878 14434
rect 4878 14382 4908 14434
rect 4932 14382 4942 14434
rect 4942 14382 4988 14434
rect 5012 14382 5058 14434
rect 5058 14382 5068 14434
rect 5092 14382 5122 14434
rect 5122 14382 5148 14434
rect 4852 14380 4908 14382
rect 4932 14380 4988 14382
rect 5012 14380 5068 14382
rect 5092 14380 5148 14382
rect 4852 13346 4908 13348
rect 4932 13346 4988 13348
rect 5012 13346 5068 13348
rect 5092 13346 5148 13348
rect 4852 13294 4878 13346
rect 4878 13294 4908 13346
rect 4932 13294 4942 13346
rect 4942 13294 4988 13346
rect 5012 13294 5058 13346
rect 5058 13294 5068 13346
rect 5092 13294 5122 13346
rect 5122 13294 5148 13346
rect 4852 13292 4908 13294
rect 4932 13292 4988 13294
rect 5012 13292 5068 13294
rect 5092 13292 5148 13294
rect 4852 12258 4908 12260
rect 4932 12258 4988 12260
rect 5012 12258 5068 12260
rect 5092 12258 5148 12260
rect 4852 12206 4878 12258
rect 4878 12206 4908 12258
rect 4932 12206 4942 12258
rect 4942 12206 4988 12258
rect 5012 12206 5058 12258
rect 5058 12206 5068 12258
rect 5092 12206 5122 12258
rect 5122 12206 5148 12258
rect 4852 12204 4908 12206
rect 4932 12204 4988 12206
rect 5012 12204 5068 12206
rect 5092 12204 5148 12206
rect 4852 11170 4908 11172
rect 4932 11170 4988 11172
rect 5012 11170 5068 11172
rect 5092 11170 5148 11172
rect 4852 11118 4878 11170
rect 4878 11118 4908 11170
rect 4932 11118 4942 11170
rect 4942 11118 4988 11170
rect 5012 11118 5058 11170
rect 5058 11118 5068 11170
rect 5092 11118 5122 11170
rect 5122 11118 5148 11170
rect 4852 11116 4908 11118
rect 4932 11116 4988 11118
rect 5012 11116 5068 11118
rect 5092 11116 5148 11118
rect 4852 10082 4908 10084
rect 4932 10082 4988 10084
rect 5012 10082 5068 10084
rect 5092 10082 5148 10084
rect 4852 10030 4878 10082
rect 4878 10030 4908 10082
rect 4932 10030 4942 10082
rect 4942 10030 4988 10082
rect 5012 10030 5058 10082
rect 5058 10030 5068 10082
rect 5092 10030 5122 10082
rect 5122 10030 5148 10082
rect 4852 10028 4908 10030
rect 4932 10028 4988 10030
rect 5012 10028 5068 10030
rect 5092 10028 5148 10030
rect 4066 6968 4122 7024
rect 4852 8994 4908 8996
rect 4932 8994 4988 8996
rect 5012 8994 5068 8996
rect 5092 8994 5148 8996
rect 4852 8942 4878 8994
rect 4878 8942 4908 8994
rect 4932 8942 4942 8994
rect 4942 8942 4988 8994
rect 5012 8942 5058 8994
rect 5058 8942 5068 8994
rect 5092 8942 5122 8994
rect 5122 8942 5148 8994
rect 4852 8940 4908 8942
rect 4932 8940 4988 8942
rect 5012 8940 5068 8942
rect 5092 8940 5148 8942
rect 4852 7906 4908 7908
rect 4932 7906 4988 7908
rect 5012 7906 5068 7908
rect 5092 7906 5148 7908
rect 4852 7854 4878 7906
rect 4878 7854 4908 7906
rect 4932 7854 4942 7906
rect 4942 7854 4988 7906
rect 5012 7854 5058 7906
rect 5058 7854 5068 7906
rect 5092 7854 5122 7906
rect 5122 7854 5148 7906
rect 4852 7852 4908 7854
rect 4932 7852 4988 7854
rect 5012 7852 5068 7854
rect 5092 7852 5148 7854
rect 4852 6818 4908 6820
rect 4932 6818 4988 6820
rect 5012 6818 5068 6820
rect 5092 6818 5148 6820
rect 4852 6766 4878 6818
rect 4878 6766 4908 6818
rect 4932 6766 4942 6818
rect 4942 6766 4988 6818
rect 5012 6766 5058 6818
rect 5058 6766 5068 6818
rect 5092 6766 5122 6818
rect 5122 6766 5148 6818
rect 4852 6764 4908 6766
rect 4932 6764 4988 6766
rect 5012 6764 5068 6766
rect 5092 6764 5148 6766
rect 4852 5730 4908 5732
rect 4932 5730 4988 5732
rect 5012 5730 5068 5732
rect 5092 5730 5148 5732
rect 4852 5678 4878 5730
rect 4878 5678 4908 5730
rect 4932 5678 4942 5730
rect 4942 5678 4988 5730
rect 5012 5678 5058 5730
rect 5058 5678 5068 5730
rect 5092 5678 5122 5730
rect 5122 5678 5148 5730
rect 4852 5676 4908 5678
rect 4932 5676 4988 5678
rect 5012 5676 5068 5678
rect 5092 5676 5148 5678
rect 2870 3296 2926 3352
rect 2254 2466 2310 2468
rect 2334 2466 2390 2468
rect 2414 2466 2470 2468
rect 2494 2466 2550 2468
rect 2254 2414 2280 2466
rect 2280 2414 2310 2466
rect 2334 2414 2344 2466
rect 2344 2414 2390 2466
rect 2414 2414 2460 2466
rect 2460 2414 2470 2466
rect 2494 2414 2524 2466
rect 2524 2414 2550 2466
rect 2254 2412 2310 2414
rect 2334 2412 2390 2414
rect 2414 2412 2470 2414
rect 2494 2412 2550 2414
rect 2254 1378 2310 1380
rect 2334 1378 2390 1380
rect 2414 1378 2470 1380
rect 2494 1378 2550 1380
rect 2254 1326 2280 1378
rect 2280 1326 2310 1378
rect 2334 1326 2344 1378
rect 2344 1326 2390 1378
rect 2414 1326 2460 1378
rect 2460 1326 2470 1378
rect 2494 1326 2524 1378
rect 2524 1326 2550 1378
rect 2254 1324 2310 1326
rect 2334 1324 2390 1326
rect 2414 1324 2470 1326
rect 2494 1324 2550 1326
rect 3553 3010 3609 3012
rect 3633 3010 3689 3012
rect 3713 3010 3769 3012
rect 3793 3010 3849 3012
rect 3553 2958 3579 3010
rect 3579 2958 3609 3010
rect 3633 2958 3643 3010
rect 3643 2958 3689 3010
rect 3713 2958 3759 3010
rect 3759 2958 3769 3010
rect 3793 2958 3823 3010
rect 3823 2958 3849 3010
rect 3553 2956 3609 2958
rect 3633 2956 3689 2958
rect 3713 2956 3769 2958
rect 3793 2956 3849 2958
rect 3553 1922 3609 1924
rect 3633 1922 3689 1924
rect 3713 1922 3769 1924
rect 3793 1922 3849 1924
rect 3553 1870 3579 1922
rect 3579 1870 3609 1922
rect 3633 1870 3643 1922
rect 3643 1870 3689 1922
rect 3713 1870 3759 1922
rect 3759 1870 3769 1922
rect 3793 1870 3823 1922
rect 3823 1870 3849 1922
rect 3553 1868 3609 1870
rect 3633 1868 3689 1870
rect 3713 1868 3769 1870
rect 3793 1868 3849 1870
rect 4066 1664 4122 1720
rect 4852 4642 4908 4644
rect 4932 4642 4988 4644
rect 5012 4642 5068 4644
rect 5092 4642 5148 4644
rect 4852 4590 4878 4642
rect 4878 4590 4908 4642
rect 4932 4590 4942 4642
rect 4942 4590 4988 4642
rect 5012 4590 5058 4642
rect 5058 4590 5068 4642
rect 5092 4590 5122 4642
rect 5122 4590 5148 4642
rect 4852 4588 4908 4590
rect 4932 4588 4988 4590
rect 5012 4588 5068 4590
rect 5092 4588 5148 4590
rect 4852 3554 4908 3556
rect 4932 3554 4988 3556
rect 5012 3554 5068 3556
rect 5092 3554 5148 3556
rect 4852 3502 4878 3554
rect 4878 3502 4908 3554
rect 4932 3502 4942 3554
rect 4942 3502 4988 3554
rect 5012 3502 5058 3554
rect 5058 3502 5068 3554
rect 5092 3502 5122 3554
rect 5122 3502 5148 3554
rect 4852 3500 4908 3502
rect 4932 3500 4988 3502
rect 5012 3500 5068 3502
rect 5092 3500 5148 3502
rect 6150 21506 6206 21508
rect 6230 21506 6286 21508
rect 6310 21506 6366 21508
rect 6390 21506 6446 21508
rect 6150 21454 6176 21506
rect 6176 21454 6206 21506
rect 6230 21454 6240 21506
rect 6240 21454 6286 21506
rect 6310 21454 6356 21506
rect 6356 21454 6366 21506
rect 6390 21454 6420 21506
rect 6420 21454 6446 21506
rect 6150 21452 6206 21454
rect 6230 21452 6286 21454
rect 6310 21452 6366 21454
rect 6390 21452 6446 21454
rect 7449 20962 7505 20964
rect 7529 20962 7585 20964
rect 7609 20962 7665 20964
rect 7689 20962 7745 20964
rect 7449 20910 7475 20962
rect 7475 20910 7505 20962
rect 7529 20910 7539 20962
rect 7539 20910 7585 20962
rect 7609 20910 7655 20962
rect 7655 20910 7665 20962
rect 7689 20910 7719 20962
rect 7719 20910 7745 20962
rect 7449 20908 7505 20910
rect 7529 20908 7585 20910
rect 7609 20908 7665 20910
rect 7689 20908 7745 20910
rect 6150 20418 6206 20420
rect 6230 20418 6286 20420
rect 6310 20418 6366 20420
rect 6390 20418 6446 20420
rect 6150 20366 6176 20418
rect 6176 20366 6206 20418
rect 6230 20366 6240 20418
rect 6240 20366 6286 20418
rect 6310 20366 6356 20418
rect 6356 20366 6366 20418
rect 6390 20366 6420 20418
rect 6420 20366 6446 20418
rect 6150 20364 6206 20366
rect 6230 20364 6286 20366
rect 6310 20364 6366 20366
rect 6390 20364 6446 20366
rect 7449 19874 7505 19876
rect 7529 19874 7585 19876
rect 7609 19874 7665 19876
rect 7689 19874 7745 19876
rect 7449 19822 7475 19874
rect 7475 19822 7505 19874
rect 7529 19822 7539 19874
rect 7539 19822 7585 19874
rect 7609 19822 7655 19874
rect 7655 19822 7665 19874
rect 7689 19822 7719 19874
rect 7719 19822 7745 19874
rect 7449 19820 7505 19822
rect 7529 19820 7585 19822
rect 7609 19820 7665 19822
rect 7689 19820 7745 19822
rect 6150 19330 6206 19332
rect 6230 19330 6286 19332
rect 6310 19330 6366 19332
rect 6390 19330 6446 19332
rect 6150 19278 6176 19330
rect 6176 19278 6206 19330
rect 6230 19278 6240 19330
rect 6240 19278 6286 19330
rect 6310 19278 6356 19330
rect 6356 19278 6366 19330
rect 6390 19278 6420 19330
rect 6420 19278 6446 19330
rect 6150 19276 6206 19278
rect 6230 19276 6286 19278
rect 6310 19276 6366 19278
rect 6390 19276 6446 19278
rect 7449 18786 7505 18788
rect 7529 18786 7585 18788
rect 7609 18786 7665 18788
rect 7689 18786 7745 18788
rect 7449 18734 7475 18786
rect 7475 18734 7505 18786
rect 7529 18734 7539 18786
rect 7539 18734 7585 18786
rect 7609 18734 7655 18786
rect 7655 18734 7665 18786
rect 7689 18734 7719 18786
rect 7719 18734 7745 18786
rect 7449 18732 7505 18734
rect 7529 18732 7585 18734
rect 7609 18732 7665 18734
rect 7689 18732 7745 18734
rect 6150 18242 6206 18244
rect 6230 18242 6286 18244
rect 6310 18242 6366 18244
rect 6390 18242 6446 18244
rect 6150 18190 6176 18242
rect 6176 18190 6206 18242
rect 6230 18190 6240 18242
rect 6240 18190 6286 18242
rect 6310 18190 6356 18242
rect 6356 18190 6366 18242
rect 6390 18190 6420 18242
rect 6420 18190 6446 18242
rect 6150 18188 6206 18190
rect 6230 18188 6286 18190
rect 6310 18188 6366 18190
rect 6390 18188 6446 18190
rect 7449 17698 7505 17700
rect 7529 17698 7585 17700
rect 7609 17698 7665 17700
rect 7689 17698 7745 17700
rect 7449 17646 7475 17698
rect 7475 17646 7505 17698
rect 7529 17646 7539 17698
rect 7539 17646 7585 17698
rect 7609 17646 7655 17698
rect 7655 17646 7665 17698
rect 7689 17646 7719 17698
rect 7719 17646 7745 17698
rect 7449 17644 7505 17646
rect 7529 17644 7585 17646
rect 7609 17644 7665 17646
rect 7689 17644 7745 17646
rect 6826 17168 6882 17224
rect 6150 17154 6206 17156
rect 6230 17154 6286 17156
rect 6310 17154 6366 17156
rect 6390 17154 6446 17156
rect 6150 17102 6176 17154
rect 6176 17102 6206 17154
rect 6230 17102 6240 17154
rect 6240 17102 6286 17154
rect 6310 17102 6356 17154
rect 6356 17102 6366 17154
rect 6390 17102 6420 17154
rect 6420 17102 6446 17154
rect 6150 17100 6206 17102
rect 6230 17100 6286 17102
rect 6310 17100 6366 17102
rect 6390 17100 6446 17102
rect 6150 16066 6206 16068
rect 6230 16066 6286 16068
rect 6310 16066 6366 16068
rect 6390 16066 6446 16068
rect 6150 16014 6176 16066
rect 6176 16014 6206 16066
rect 6230 16014 6240 16066
rect 6240 16014 6286 16066
rect 6310 16014 6356 16066
rect 6356 16014 6366 16066
rect 6390 16014 6420 16066
rect 6420 16014 6446 16066
rect 6150 16012 6206 16014
rect 6230 16012 6286 16014
rect 6310 16012 6366 16014
rect 6390 16012 6446 16014
rect 6150 14978 6206 14980
rect 6230 14978 6286 14980
rect 6310 14978 6366 14980
rect 6390 14978 6446 14980
rect 6150 14926 6176 14978
rect 6176 14926 6206 14978
rect 6230 14926 6240 14978
rect 6240 14926 6286 14978
rect 6310 14926 6356 14978
rect 6356 14926 6366 14978
rect 6390 14926 6420 14978
rect 6420 14926 6446 14978
rect 6150 14924 6206 14926
rect 6230 14924 6286 14926
rect 6310 14924 6366 14926
rect 6390 14924 6446 14926
rect 7449 16610 7505 16612
rect 7529 16610 7585 16612
rect 7609 16610 7665 16612
rect 7689 16610 7745 16612
rect 7449 16558 7475 16610
rect 7475 16558 7505 16610
rect 7529 16558 7539 16610
rect 7539 16558 7585 16610
rect 7609 16558 7655 16610
rect 7655 16558 7665 16610
rect 7689 16558 7719 16610
rect 7719 16558 7745 16610
rect 7449 16556 7505 16558
rect 7529 16556 7585 16558
rect 7609 16556 7665 16558
rect 7689 16556 7745 16558
rect 7449 15522 7505 15524
rect 7529 15522 7585 15524
rect 7609 15522 7665 15524
rect 7689 15522 7745 15524
rect 7449 15470 7475 15522
rect 7475 15470 7505 15522
rect 7529 15470 7539 15522
rect 7539 15470 7585 15522
rect 7609 15470 7655 15522
rect 7655 15470 7665 15522
rect 7689 15470 7719 15522
rect 7719 15470 7745 15522
rect 7449 15468 7505 15470
rect 7529 15468 7585 15470
rect 7609 15468 7665 15470
rect 7689 15468 7745 15470
rect 6150 13890 6206 13892
rect 6230 13890 6286 13892
rect 6310 13890 6366 13892
rect 6390 13890 6446 13892
rect 6150 13838 6176 13890
rect 6176 13838 6206 13890
rect 6230 13838 6240 13890
rect 6240 13838 6286 13890
rect 6310 13838 6356 13890
rect 6356 13838 6366 13890
rect 6390 13838 6420 13890
rect 6420 13838 6446 13890
rect 6150 13836 6206 13838
rect 6230 13836 6286 13838
rect 6310 13836 6366 13838
rect 6390 13836 6446 13838
rect 6150 12802 6206 12804
rect 6230 12802 6286 12804
rect 6310 12802 6366 12804
rect 6390 12802 6446 12804
rect 6150 12750 6176 12802
rect 6176 12750 6206 12802
rect 6230 12750 6240 12802
rect 6240 12750 6286 12802
rect 6310 12750 6356 12802
rect 6356 12750 6366 12802
rect 6390 12750 6420 12802
rect 6420 12750 6446 12802
rect 6150 12748 6206 12750
rect 6230 12748 6286 12750
rect 6310 12748 6366 12750
rect 6390 12748 6446 12750
rect 6150 11714 6206 11716
rect 6230 11714 6286 11716
rect 6310 11714 6366 11716
rect 6390 11714 6446 11716
rect 6150 11662 6176 11714
rect 6176 11662 6206 11714
rect 6230 11662 6240 11714
rect 6240 11662 6286 11714
rect 6310 11662 6356 11714
rect 6356 11662 6366 11714
rect 6390 11662 6420 11714
rect 6420 11662 6446 11714
rect 6150 11660 6206 11662
rect 6230 11660 6286 11662
rect 6310 11660 6366 11662
rect 6390 11660 6446 11662
rect 7838 14448 7894 14504
rect 7449 14434 7505 14436
rect 7529 14434 7585 14436
rect 7609 14434 7665 14436
rect 7689 14434 7745 14436
rect 7449 14382 7475 14434
rect 7475 14382 7505 14434
rect 7529 14382 7539 14434
rect 7539 14382 7585 14434
rect 7609 14382 7655 14434
rect 7655 14382 7665 14434
rect 7689 14382 7719 14434
rect 7719 14382 7745 14434
rect 7449 14380 7505 14382
rect 7529 14380 7585 14382
rect 7609 14380 7665 14382
rect 7689 14380 7745 14382
rect 6826 11592 6882 11648
rect 6150 10626 6206 10628
rect 6230 10626 6286 10628
rect 6310 10626 6366 10628
rect 6390 10626 6446 10628
rect 6150 10574 6176 10626
rect 6176 10574 6206 10626
rect 6230 10574 6240 10626
rect 6240 10574 6286 10626
rect 6310 10574 6356 10626
rect 6356 10574 6366 10626
rect 6390 10574 6420 10626
rect 6420 10574 6446 10626
rect 6150 10572 6206 10574
rect 6230 10572 6286 10574
rect 6310 10572 6366 10574
rect 6390 10572 6446 10574
rect 6150 9538 6206 9540
rect 6230 9538 6286 9540
rect 6310 9538 6366 9540
rect 6390 9538 6446 9540
rect 6150 9486 6176 9538
rect 6176 9486 6206 9538
rect 6230 9486 6240 9538
rect 6240 9486 6286 9538
rect 6310 9486 6356 9538
rect 6356 9486 6366 9538
rect 6390 9486 6420 9538
rect 6420 9486 6446 9538
rect 6150 9484 6206 9486
rect 6230 9484 6286 9486
rect 6310 9484 6366 9486
rect 6390 9484 6446 9486
rect 6150 8450 6206 8452
rect 6230 8450 6286 8452
rect 6310 8450 6366 8452
rect 6390 8450 6446 8452
rect 6150 8398 6176 8450
rect 6176 8398 6206 8450
rect 6230 8398 6240 8450
rect 6240 8398 6286 8450
rect 6310 8398 6356 8450
rect 6356 8398 6366 8450
rect 6390 8398 6420 8450
rect 6420 8398 6446 8450
rect 6150 8396 6206 8398
rect 6230 8396 6286 8398
rect 6310 8396 6366 8398
rect 6390 8396 6446 8398
rect 6150 7362 6206 7364
rect 6230 7362 6286 7364
rect 6310 7362 6366 7364
rect 6390 7362 6446 7364
rect 6150 7310 6176 7362
rect 6176 7310 6206 7362
rect 6230 7310 6240 7362
rect 6240 7310 6286 7362
rect 6310 7310 6356 7362
rect 6356 7310 6366 7362
rect 6390 7310 6420 7362
rect 6420 7310 6446 7362
rect 6150 7308 6206 7310
rect 6230 7308 6286 7310
rect 6310 7308 6366 7310
rect 6390 7308 6446 7310
rect 6150 6274 6206 6276
rect 6230 6274 6286 6276
rect 6310 6274 6366 6276
rect 6390 6274 6446 6276
rect 6150 6222 6176 6274
rect 6176 6222 6206 6274
rect 6230 6222 6240 6274
rect 6240 6222 6286 6274
rect 6310 6222 6356 6274
rect 6356 6222 6366 6274
rect 6390 6222 6420 6274
rect 6420 6222 6446 6274
rect 6150 6220 6206 6222
rect 6230 6220 6286 6222
rect 6310 6220 6366 6222
rect 6390 6220 6446 6222
rect 5630 6016 5686 6072
rect 6150 5186 6206 5188
rect 6230 5186 6286 5188
rect 6310 5186 6366 5188
rect 6390 5186 6446 5188
rect 6150 5134 6176 5186
rect 6176 5134 6206 5186
rect 6230 5134 6240 5186
rect 6240 5134 6286 5186
rect 6310 5134 6356 5186
rect 6356 5134 6366 5186
rect 6390 5134 6420 5186
rect 6420 5134 6446 5186
rect 6150 5132 6206 5134
rect 6230 5132 6286 5134
rect 6310 5132 6366 5134
rect 6390 5132 6446 5134
rect 6150 4098 6206 4100
rect 6230 4098 6286 4100
rect 6310 4098 6366 4100
rect 6390 4098 6446 4100
rect 6150 4046 6176 4098
rect 6176 4046 6206 4098
rect 6230 4046 6240 4098
rect 6240 4046 6286 4098
rect 6310 4046 6356 4098
rect 6356 4046 6366 4098
rect 6390 4046 6420 4098
rect 6420 4046 6446 4098
rect 6150 4044 6206 4046
rect 6230 4044 6286 4046
rect 6310 4044 6366 4046
rect 6390 4044 6446 4046
rect 7449 13346 7505 13348
rect 7529 13346 7585 13348
rect 7609 13346 7665 13348
rect 7689 13346 7745 13348
rect 7449 13294 7475 13346
rect 7475 13294 7505 13346
rect 7529 13294 7539 13346
rect 7539 13294 7585 13346
rect 7609 13294 7655 13346
rect 7655 13294 7665 13346
rect 7689 13294 7719 13346
rect 7719 13294 7745 13346
rect 7449 13292 7505 13294
rect 7529 13292 7585 13294
rect 7609 13292 7665 13294
rect 7689 13292 7745 13294
rect 7449 12258 7505 12260
rect 7529 12258 7585 12260
rect 7609 12258 7665 12260
rect 7689 12258 7745 12260
rect 7449 12206 7475 12258
rect 7475 12206 7505 12258
rect 7529 12206 7539 12258
rect 7539 12206 7585 12258
rect 7609 12206 7655 12258
rect 7655 12206 7665 12258
rect 7689 12206 7719 12258
rect 7719 12206 7745 12258
rect 7449 12204 7505 12206
rect 7529 12204 7585 12206
rect 7609 12204 7665 12206
rect 7689 12204 7745 12206
rect 7449 11170 7505 11172
rect 7529 11170 7585 11172
rect 7609 11170 7665 11172
rect 7689 11170 7745 11172
rect 7449 11118 7475 11170
rect 7475 11118 7505 11170
rect 7529 11118 7539 11170
rect 7539 11118 7585 11170
rect 7609 11118 7655 11170
rect 7655 11118 7665 11170
rect 7689 11118 7719 11170
rect 7719 11118 7745 11170
rect 7449 11116 7505 11118
rect 7529 11116 7585 11118
rect 7609 11116 7665 11118
rect 7689 11116 7745 11118
rect 7449 10082 7505 10084
rect 7529 10082 7585 10084
rect 7609 10082 7665 10084
rect 7689 10082 7745 10084
rect 7449 10030 7475 10082
rect 7475 10030 7505 10082
rect 7529 10030 7539 10082
rect 7539 10030 7585 10082
rect 7609 10030 7655 10082
rect 7655 10030 7665 10082
rect 7689 10030 7719 10082
rect 7719 10030 7745 10082
rect 7449 10028 7505 10030
rect 7529 10028 7585 10030
rect 7609 10028 7665 10030
rect 7689 10028 7745 10030
rect 7449 8994 7505 8996
rect 7529 8994 7585 8996
rect 7609 8994 7665 8996
rect 7689 8994 7745 8996
rect 7449 8942 7475 8994
rect 7475 8942 7505 8994
rect 7529 8942 7539 8994
rect 7539 8942 7585 8994
rect 7609 8942 7655 8994
rect 7655 8942 7665 8994
rect 7689 8942 7719 8994
rect 7719 8942 7745 8994
rect 7449 8940 7505 8942
rect 7529 8940 7585 8942
rect 7609 8940 7665 8942
rect 7689 8940 7745 8942
rect 8206 8872 8262 8928
rect 7449 7906 7505 7908
rect 7529 7906 7585 7908
rect 7609 7906 7665 7908
rect 7689 7906 7745 7908
rect 7449 7854 7475 7906
rect 7475 7854 7505 7906
rect 7529 7854 7539 7906
rect 7539 7854 7585 7906
rect 7609 7854 7655 7906
rect 7655 7854 7665 7906
rect 7689 7854 7719 7906
rect 7719 7854 7745 7906
rect 7449 7852 7505 7854
rect 7529 7852 7585 7854
rect 7609 7852 7665 7854
rect 7689 7852 7745 7854
rect 7449 6818 7505 6820
rect 7529 6818 7585 6820
rect 7609 6818 7665 6820
rect 7689 6818 7745 6820
rect 7449 6766 7475 6818
rect 7475 6766 7505 6818
rect 7529 6766 7539 6818
rect 7539 6766 7585 6818
rect 7609 6766 7655 6818
rect 7655 6766 7665 6818
rect 7689 6766 7719 6818
rect 7719 6766 7745 6818
rect 7449 6764 7505 6766
rect 7529 6764 7585 6766
rect 7609 6764 7665 6766
rect 7689 6764 7745 6766
rect 7449 5730 7505 5732
rect 7529 5730 7585 5732
rect 7609 5730 7665 5732
rect 7689 5730 7745 5732
rect 7449 5678 7475 5730
rect 7475 5678 7505 5730
rect 7529 5678 7539 5730
rect 7539 5678 7585 5730
rect 7609 5678 7655 5730
rect 7655 5678 7665 5730
rect 7689 5678 7719 5730
rect 7719 5678 7745 5730
rect 7449 5676 7505 5678
rect 7529 5676 7585 5678
rect 7609 5676 7665 5678
rect 7689 5676 7745 5678
rect 7449 4642 7505 4644
rect 7529 4642 7585 4644
rect 7609 4642 7665 4644
rect 7689 4642 7745 4644
rect 7449 4590 7475 4642
rect 7475 4590 7505 4642
rect 7529 4590 7539 4642
rect 7539 4590 7585 4642
rect 7609 4590 7655 4642
rect 7655 4590 7665 4642
rect 7689 4590 7719 4642
rect 7719 4590 7745 4642
rect 7449 4588 7505 4590
rect 7529 4588 7585 4590
rect 7609 4588 7665 4590
rect 7689 4588 7745 4590
rect 7449 3554 7505 3556
rect 7529 3554 7585 3556
rect 7609 3554 7665 3556
rect 7689 3554 7745 3556
rect 7449 3502 7475 3554
rect 7475 3502 7505 3554
rect 7529 3502 7539 3554
rect 7539 3502 7585 3554
rect 7609 3502 7655 3554
rect 7655 3502 7665 3554
rect 7689 3502 7719 3554
rect 7719 3502 7745 3554
rect 7449 3500 7505 3502
rect 7529 3500 7585 3502
rect 7609 3500 7665 3502
rect 7689 3500 7745 3502
rect 6642 3296 6698 3352
rect 6150 3010 6206 3012
rect 6230 3010 6286 3012
rect 6310 3010 6366 3012
rect 6390 3010 6446 3012
rect 6150 2958 6176 3010
rect 6176 2958 6206 3010
rect 6230 2958 6240 3010
rect 6240 2958 6286 3010
rect 6310 2958 6356 3010
rect 6356 2958 6366 3010
rect 6390 2958 6420 3010
rect 6420 2958 6446 3010
rect 6150 2956 6206 2958
rect 6230 2956 6286 2958
rect 6310 2956 6366 2958
rect 6390 2956 6446 2958
rect 4852 2466 4908 2468
rect 4932 2466 4988 2468
rect 5012 2466 5068 2468
rect 5092 2466 5148 2468
rect 4852 2414 4878 2466
rect 4878 2414 4908 2466
rect 4932 2414 4942 2466
rect 4942 2414 4988 2466
rect 5012 2414 5058 2466
rect 5058 2414 5068 2466
rect 5092 2414 5122 2466
rect 5122 2414 5148 2466
rect 4852 2412 4908 2414
rect 4932 2412 4988 2414
rect 5012 2412 5068 2414
rect 5092 2412 5148 2414
rect 6150 1922 6206 1924
rect 6230 1922 6286 1924
rect 6310 1922 6366 1924
rect 6390 1922 6446 1924
rect 6150 1870 6176 1922
rect 6176 1870 6206 1922
rect 6230 1870 6240 1922
rect 6240 1870 6286 1922
rect 6310 1870 6356 1922
rect 6356 1870 6366 1922
rect 6390 1870 6420 1922
rect 6420 1870 6446 1922
rect 6150 1868 6206 1870
rect 6230 1868 6286 1870
rect 6310 1868 6366 1870
rect 6390 1868 6446 1870
rect 4852 1378 4908 1380
rect 4932 1378 4988 1380
rect 5012 1378 5068 1380
rect 5092 1378 5148 1380
rect 4852 1326 4878 1378
rect 4878 1326 4908 1378
rect 4932 1326 4942 1378
rect 4942 1326 4988 1378
rect 5012 1326 5058 1378
rect 5058 1326 5068 1378
rect 5092 1326 5122 1378
rect 5122 1326 5148 1378
rect 4852 1324 4908 1326
rect 4932 1324 4988 1326
rect 5012 1324 5068 1326
rect 5092 1324 5148 1326
rect 7449 2466 7505 2468
rect 7529 2466 7585 2468
rect 7609 2466 7665 2468
rect 7689 2466 7745 2468
rect 7449 2414 7475 2466
rect 7475 2414 7505 2466
rect 7529 2414 7539 2466
rect 7539 2414 7585 2466
rect 7609 2414 7655 2466
rect 7655 2414 7665 2466
rect 7689 2414 7719 2466
rect 7719 2414 7745 2466
rect 7449 2412 7505 2414
rect 7529 2412 7585 2414
rect 7609 2412 7665 2414
rect 7689 2412 7745 2414
rect 7449 1378 7505 1380
rect 7529 1378 7585 1380
rect 7609 1378 7665 1380
rect 7689 1378 7745 1380
rect 7449 1326 7475 1378
rect 7475 1326 7505 1378
rect 7529 1326 7539 1378
rect 7539 1326 7585 1378
rect 7609 1326 7655 1378
rect 7655 1326 7665 1378
rect 7689 1326 7719 1378
rect 7719 1326 7745 1378
rect 7449 1324 7505 1326
rect 7529 1324 7585 1326
rect 7609 1324 7665 1326
rect 7689 1324 7745 1326
rect 6826 576 6882 632
rect 3422 32 3478 88
<< metal3 >>
rect 0 23346 480 23376
rect 4061 23346 4127 23349
rect 0 23344 4127 23346
rect 0 23288 4066 23344
rect 4122 23288 4127 23344
rect 0 23286 4127 23288
rect 0 23256 480 23286
rect 4061 23283 4127 23286
rect 5809 22802 5875 22805
rect 9520 22802 10000 22832
rect 5809 22800 10000 22802
rect 5809 22744 5814 22800
rect 5870 22744 10000 22800
rect 5809 22742 10000 22744
rect 5809 22739 5875 22742
rect 9520 22712 10000 22742
rect 0 21714 480 21744
rect 3417 21714 3483 21717
rect 0 21712 3483 21714
rect 0 21656 3422 21712
rect 3478 21656 3483 21712
rect 0 21654 3483 21656
rect 0 21624 480 21654
rect 3417 21651 3483 21654
rect 3541 21512 3861 21513
rect 3541 21448 3549 21512
rect 3613 21448 3629 21512
rect 3693 21448 3709 21512
rect 3773 21448 3789 21512
rect 3853 21448 3861 21512
rect 3541 21447 3861 21448
rect 6138 21512 6458 21513
rect 6138 21448 6146 21512
rect 6210 21448 6226 21512
rect 6290 21448 6306 21512
rect 6370 21448 6386 21512
rect 6450 21448 6458 21512
rect 6138 21447 6458 21448
rect 2242 20968 2562 20969
rect 2242 20904 2250 20968
rect 2314 20904 2330 20968
rect 2394 20904 2410 20968
rect 2474 20904 2490 20968
rect 2554 20904 2562 20968
rect 2242 20903 2562 20904
rect 4840 20968 5160 20969
rect 4840 20904 4848 20968
rect 4912 20904 4928 20968
rect 4992 20904 5008 20968
rect 5072 20904 5088 20968
rect 5152 20904 5160 20968
rect 4840 20903 5160 20904
rect 7437 20968 7757 20969
rect 7437 20904 7445 20968
rect 7509 20904 7525 20968
rect 7589 20904 7605 20968
rect 7669 20904 7685 20968
rect 7749 20904 7757 20968
rect 7437 20903 7757 20904
rect 3541 20424 3861 20425
rect 3541 20360 3549 20424
rect 3613 20360 3629 20424
rect 3693 20360 3709 20424
rect 3773 20360 3789 20424
rect 3853 20360 3861 20424
rect 3541 20359 3861 20360
rect 6138 20424 6458 20425
rect 6138 20360 6146 20424
rect 6210 20360 6226 20424
rect 6290 20360 6306 20424
rect 6370 20360 6386 20424
rect 6450 20360 6458 20424
rect 6138 20359 6458 20360
rect 0 20082 480 20112
rect 3049 20082 3115 20085
rect 0 20080 3115 20082
rect 0 20024 3054 20080
rect 3110 20024 3115 20080
rect 0 20022 3115 20024
rect 0 19992 480 20022
rect 3049 20019 3115 20022
rect 5717 20082 5783 20085
rect 9520 20082 10000 20112
rect 5717 20080 10000 20082
rect 5717 20024 5722 20080
rect 5778 20024 10000 20080
rect 5717 20022 10000 20024
rect 5717 20019 5783 20022
rect 9520 19992 10000 20022
rect 2242 19880 2562 19881
rect 2242 19816 2250 19880
rect 2314 19816 2330 19880
rect 2394 19816 2410 19880
rect 2474 19816 2490 19880
rect 2554 19816 2562 19880
rect 2242 19815 2562 19816
rect 4840 19880 5160 19881
rect 4840 19816 4848 19880
rect 4912 19816 4928 19880
rect 4992 19816 5008 19880
rect 5072 19816 5088 19880
rect 5152 19816 5160 19880
rect 4840 19815 5160 19816
rect 7437 19880 7757 19881
rect 7437 19816 7445 19880
rect 7509 19816 7525 19880
rect 7589 19816 7605 19880
rect 7669 19816 7685 19880
rect 7749 19816 7757 19880
rect 7437 19815 7757 19816
rect 3541 19336 3861 19337
rect 3541 19272 3549 19336
rect 3613 19272 3629 19336
rect 3693 19272 3709 19336
rect 3773 19272 3789 19336
rect 3853 19272 3861 19336
rect 3541 19271 3861 19272
rect 6138 19336 6458 19337
rect 6138 19272 6146 19336
rect 6210 19272 6226 19336
rect 6290 19272 6306 19336
rect 6370 19272 6386 19336
rect 6450 19272 6458 19336
rect 6138 19271 6458 19272
rect 2242 18792 2562 18793
rect 2242 18728 2250 18792
rect 2314 18728 2330 18792
rect 2394 18728 2410 18792
rect 2474 18728 2490 18792
rect 2554 18728 2562 18792
rect 2242 18727 2562 18728
rect 4840 18792 5160 18793
rect 4840 18728 4848 18792
rect 4912 18728 4928 18792
rect 4992 18728 5008 18792
rect 5072 18728 5088 18792
rect 5152 18728 5160 18792
rect 4840 18727 5160 18728
rect 7437 18792 7757 18793
rect 7437 18728 7445 18792
rect 7509 18728 7525 18792
rect 7589 18728 7605 18792
rect 7669 18728 7685 18792
rect 7749 18728 7757 18792
rect 7437 18727 7757 18728
rect 0 18314 480 18344
rect 3233 18314 3299 18317
rect 0 18312 3299 18314
rect 0 18256 3238 18312
rect 3294 18256 3299 18312
rect 0 18254 3299 18256
rect 0 18224 480 18254
rect 3233 18251 3299 18254
rect 3541 18248 3861 18249
rect 3541 18184 3549 18248
rect 3613 18184 3629 18248
rect 3693 18184 3709 18248
rect 3773 18184 3789 18248
rect 3853 18184 3861 18248
rect 3541 18183 3861 18184
rect 6138 18248 6458 18249
rect 6138 18184 6146 18248
rect 6210 18184 6226 18248
rect 6290 18184 6306 18248
rect 6370 18184 6386 18248
rect 6450 18184 6458 18248
rect 6138 18183 6458 18184
rect 2242 17704 2562 17705
rect 2242 17640 2250 17704
rect 2314 17640 2330 17704
rect 2394 17640 2410 17704
rect 2474 17640 2490 17704
rect 2554 17640 2562 17704
rect 2242 17639 2562 17640
rect 4840 17704 5160 17705
rect 4840 17640 4848 17704
rect 4912 17640 4928 17704
rect 4992 17640 5008 17704
rect 5072 17640 5088 17704
rect 5152 17640 5160 17704
rect 4840 17639 5160 17640
rect 7437 17704 7757 17705
rect 7437 17640 7445 17704
rect 7509 17640 7525 17704
rect 7589 17640 7605 17704
rect 7669 17640 7685 17704
rect 7749 17640 7757 17704
rect 7437 17639 7757 17640
rect 6821 17226 6887 17229
rect 9520 17226 10000 17256
rect 6821 17224 10000 17226
rect 6821 17168 6826 17224
rect 6882 17168 10000 17224
rect 6821 17166 10000 17168
rect 6821 17163 6887 17166
rect 3541 17160 3861 17161
rect 3541 17096 3549 17160
rect 3613 17096 3629 17160
rect 3693 17096 3709 17160
rect 3773 17096 3789 17160
rect 3853 17096 3861 17160
rect 3541 17095 3861 17096
rect 6138 17160 6458 17161
rect 6138 17096 6146 17160
rect 6210 17096 6226 17160
rect 6290 17096 6306 17160
rect 6370 17096 6386 17160
rect 6450 17096 6458 17160
rect 9520 17136 10000 17166
rect 6138 17095 6458 17096
rect 0 16682 480 16712
rect 0 16622 2146 16682
rect 0 16592 480 16622
rect 2086 16410 2146 16622
rect 2242 16616 2562 16617
rect 2242 16552 2250 16616
rect 2314 16552 2330 16616
rect 2394 16552 2410 16616
rect 2474 16552 2490 16616
rect 2554 16552 2562 16616
rect 2242 16551 2562 16552
rect 4840 16616 5160 16617
rect 4840 16552 4848 16616
rect 4912 16552 4928 16616
rect 4992 16552 5008 16616
rect 5072 16552 5088 16616
rect 5152 16552 5160 16616
rect 4840 16551 5160 16552
rect 7437 16616 7757 16617
rect 7437 16552 7445 16616
rect 7509 16552 7525 16616
rect 7589 16552 7605 16616
rect 7669 16552 7685 16616
rect 7749 16552 7757 16616
rect 7437 16551 7757 16552
rect 4061 16410 4127 16413
rect 2086 16408 4127 16410
rect 2086 16352 4066 16408
rect 4122 16352 4127 16408
rect 2086 16350 4127 16352
rect 4061 16347 4127 16350
rect 3541 16072 3861 16073
rect 3541 16008 3549 16072
rect 3613 16008 3629 16072
rect 3693 16008 3709 16072
rect 3773 16008 3789 16072
rect 3853 16008 3861 16072
rect 3541 16007 3861 16008
rect 6138 16072 6458 16073
rect 6138 16008 6146 16072
rect 6210 16008 6226 16072
rect 6290 16008 6306 16072
rect 6370 16008 6386 16072
rect 6450 16008 6458 16072
rect 6138 16007 6458 16008
rect 2242 15528 2562 15529
rect 2242 15464 2250 15528
rect 2314 15464 2330 15528
rect 2394 15464 2410 15528
rect 2474 15464 2490 15528
rect 2554 15464 2562 15528
rect 2242 15463 2562 15464
rect 4840 15528 5160 15529
rect 4840 15464 4848 15528
rect 4912 15464 4928 15528
rect 4992 15464 5008 15528
rect 5072 15464 5088 15528
rect 5152 15464 5160 15528
rect 4840 15463 5160 15464
rect 7437 15528 7757 15529
rect 7437 15464 7445 15528
rect 7509 15464 7525 15528
rect 7589 15464 7605 15528
rect 7669 15464 7685 15528
rect 7749 15464 7757 15528
rect 7437 15463 7757 15464
rect 0 15050 480 15080
rect 3049 15050 3115 15053
rect 0 15048 3115 15050
rect 0 14992 3054 15048
rect 3110 14992 3115 15048
rect 0 14990 3115 14992
rect 0 14960 480 14990
rect 3049 14987 3115 14990
rect 3541 14984 3861 14985
rect 3541 14920 3549 14984
rect 3613 14920 3629 14984
rect 3693 14920 3709 14984
rect 3773 14920 3789 14984
rect 3853 14920 3861 14984
rect 3541 14919 3861 14920
rect 6138 14984 6458 14985
rect 6138 14920 6146 14984
rect 6210 14920 6226 14984
rect 6290 14920 6306 14984
rect 6370 14920 6386 14984
rect 6450 14920 6458 14984
rect 6138 14919 6458 14920
rect 7833 14506 7899 14509
rect 9520 14506 10000 14536
rect 7833 14504 10000 14506
rect 7833 14448 7838 14504
rect 7894 14448 10000 14504
rect 7833 14446 10000 14448
rect 7833 14443 7899 14446
rect 2242 14440 2562 14441
rect 2242 14376 2250 14440
rect 2314 14376 2330 14440
rect 2394 14376 2410 14440
rect 2474 14376 2490 14440
rect 2554 14376 2562 14440
rect 2242 14375 2562 14376
rect 4840 14440 5160 14441
rect 4840 14376 4848 14440
rect 4912 14376 4928 14440
rect 4992 14376 5008 14440
rect 5072 14376 5088 14440
rect 5152 14376 5160 14440
rect 4840 14375 5160 14376
rect 7437 14440 7757 14441
rect 7437 14376 7445 14440
rect 7509 14376 7525 14440
rect 7589 14376 7605 14440
rect 7669 14376 7685 14440
rect 7749 14376 7757 14440
rect 9520 14416 10000 14446
rect 7437 14375 7757 14376
rect 3541 13896 3861 13897
rect 3541 13832 3549 13896
rect 3613 13832 3629 13896
rect 3693 13832 3709 13896
rect 3773 13832 3789 13896
rect 3853 13832 3861 13896
rect 3541 13831 3861 13832
rect 6138 13896 6458 13897
rect 6138 13832 6146 13896
rect 6210 13832 6226 13896
rect 6290 13832 6306 13896
rect 6370 13832 6386 13896
rect 6450 13832 6458 13896
rect 6138 13831 6458 13832
rect 4061 13554 4127 13557
rect 2086 13552 4127 13554
rect 2086 13496 4066 13552
rect 4122 13496 4127 13552
rect 2086 13494 4127 13496
rect 0 13418 480 13448
rect 2086 13418 2146 13494
rect 4061 13491 4127 13494
rect 0 13358 2146 13418
rect 0 13328 480 13358
rect 2242 13352 2562 13353
rect 2242 13288 2250 13352
rect 2314 13288 2330 13352
rect 2394 13288 2410 13352
rect 2474 13288 2490 13352
rect 2554 13288 2562 13352
rect 2242 13287 2562 13288
rect 4840 13352 5160 13353
rect 4840 13288 4848 13352
rect 4912 13288 4928 13352
rect 4992 13288 5008 13352
rect 5072 13288 5088 13352
rect 5152 13288 5160 13352
rect 4840 13287 5160 13288
rect 7437 13352 7757 13353
rect 7437 13288 7445 13352
rect 7509 13288 7525 13352
rect 7589 13288 7605 13352
rect 7669 13288 7685 13352
rect 7749 13288 7757 13352
rect 7437 13287 7757 13288
rect 3541 12808 3861 12809
rect 3541 12744 3549 12808
rect 3613 12744 3629 12808
rect 3693 12744 3709 12808
rect 3773 12744 3789 12808
rect 3853 12744 3861 12808
rect 3541 12743 3861 12744
rect 6138 12808 6458 12809
rect 6138 12744 6146 12808
rect 6210 12744 6226 12808
rect 6290 12744 6306 12808
rect 6370 12744 6386 12808
rect 6450 12744 6458 12808
rect 6138 12743 6458 12744
rect 2242 12264 2562 12265
rect 2242 12200 2250 12264
rect 2314 12200 2330 12264
rect 2394 12200 2410 12264
rect 2474 12200 2490 12264
rect 2554 12200 2562 12264
rect 2242 12199 2562 12200
rect 4840 12264 5160 12265
rect 4840 12200 4848 12264
rect 4912 12200 4928 12264
rect 4992 12200 5008 12264
rect 5072 12200 5088 12264
rect 5152 12200 5160 12264
rect 4840 12199 5160 12200
rect 7437 12264 7757 12265
rect 7437 12200 7445 12264
rect 7509 12200 7525 12264
rect 7589 12200 7605 12264
rect 7669 12200 7685 12264
rect 7749 12200 7757 12264
rect 7437 12199 7757 12200
rect 3541 11720 3861 11721
rect 0 11650 480 11680
rect 3541 11656 3549 11720
rect 3613 11656 3629 11720
rect 3693 11656 3709 11720
rect 3773 11656 3789 11720
rect 3853 11656 3861 11720
rect 3541 11655 3861 11656
rect 6138 11720 6458 11721
rect 6138 11656 6146 11720
rect 6210 11656 6226 11720
rect 6290 11656 6306 11720
rect 6370 11656 6386 11720
rect 6450 11656 6458 11720
rect 6138 11655 6458 11656
rect 3233 11650 3299 11653
rect 0 11648 3299 11650
rect 0 11592 3238 11648
rect 3294 11592 3299 11648
rect 0 11590 3299 11592
rect 0 11560 480 11590
rect 3233 11587 3299 11590
rect 6821 11650 6887 11653
rect 9520 11650 10000 11680
rect 6821 11648 10000 11650
rect 6821 11592 6826 11648
rect 6882 11592 10000 11648
rect 6821 11590 10000 11592
rect 6821 11587 6887 11590
rect 9520 11560 10000 11590
rect 2242 11176 2562 11177
rect 2242 11112 2250 11176
rect 2314 11112 2330 11176
rect 2394 11112 2410 11176
rect 2474 11112 2490 11176
rect 2554 11112 2562 11176
rect 2242 11111 2562 11112
rect 4840 11176 5160 11177
rect 4840 11112 4848 11176
rect 4912 11112 4928 11176
rect 4992 11112 5008 11176
rect 5072 11112 5088 11176
rect 5152 11112 5160 11176
rect 4840 11111 5160 11112
rect 7437 11176 7757 11177
rect 7437 11112 7445 11176
rect 7509 11112 7525 11176
rect 7589 11112 7605 11176
rect 7669 11112 7685 11176
rect 7749 11112 7757 11176
rect 7437 11111 7757 11112
rect 3541 10632 3861 10633
rect 3541 10568 3549 10632
rect 3613 10568 3629 10632
rect 3693 10568 3709 10632
rect 3773 10568 3789 10632
rect 3853 10568 3861 10632
rect 3541 10567 3861 10568
rect 6138 10632 6458 10633
rect 6138 10568 6146 10632
rect 6210 10568 6226 10632
rect 6290 10568 6306 10632
rect 6370 10568 6386 10632
rect 6450 10568 6458 10632
rect 6138 10567 6458 10568
rect 2242 10088 2562 10089
rect 0 10018 480 10048
rect 2242 10024 2250 10088
rect 2314 10024 2330 10088
rect 2394 10024 2410 10088
rect 2474 10024 2490 10088
rect 2554 10024 2562 10088
rect 2242 10023 2562 10024
rect 4840 10088 5160 10089
rect 4840 10024 4848 10088
rect 4912 10024 4928 10088
rect 4992 10024 5008 10088
rect 5072 10024 5088 10088
rect 5152 10024 5160 10088
rect 4840 10023 5160 10024
rect 7437 10088 7757 10089
rect 7437 10024 7445 10088
rect 7509 10024 7525 10088
rect 7589 10024 7605 10088
rect 7669 10024 7685 10088
rect 7749 10024 7757 10088
rect 7437 10023 7757 10024
rect 0 9958 2146 10018
rect 0 9928 480 9958
rect 2086 9882 2146 9958
rect 3417 9882 3483 9885
rect 2086 9880 3483 9882
rect 2086 9824 3422 9880
rect 3478 9824 3483 9880
rect 2086 9822 3483 9824
rect 3417 9819 3483 9822
rect 3541 9544 3861 9545
rect 3541 9480 3549 9544
rect 3613 9480 3629 9544
rect 3693 9480 3709 9544
rect 3773 9480 3789 9544
rect 3853 9480 3861 9544
rect 3541 9479 3861 9480
rect 6138 9544 6458 9545
rect 6138 9480 6146 9544
rect 6210 9480 6226 9544
rect 6290 9480 6306 9544
rect 6370 9480 6386 9544
rect 6450 9480 6458 9544
rect 6138 9479 6458 9480
rect 2242 9000 2562 9001
rect 2242 8936 2250 9000
rect 2314 8936 2330 9000
rect 2394 8936 2410 9000
rect 2474 8936 2490 9000
rect 2554 8936 2562 9000
rect 2242 8935 2562 8936
rect 4840 9000 5160 9001
rect 4840 8936 4848 9000
rect 4912 8936 4928 9000
rect 4992 8936 5008 9000
rect 5072 8936 5088 9000
rect 5152 8936 5160 9000
rect 4840 8935 5160 8936
rect 7437 9000 7757 9001
rect 7437 8936 7445 9000
rect 7509 8936 7525 9000
rect 7589 8936 7605 9000
rect 7669 8936 7685 9000
rect 7749 8936 7757 9000
rect 7437 8935 7757 8936
rect 8201 8930 8267 8933
rect 9520 8930 10000 8960
rect 8201 8928 10000 8930
rect 8201 8872 8206 8928
rect 8262 8872 10000 8928
rect 8201 8870 10000 8872
rect 8201 8867 8267 8870
rect 9520 8840 10000 8870
rect 3541 8456 3861 8457
rect 0 8386 480 8416
rect 3541 8392 3549 8456
rect 3613 8392 3629 8456
rect 3693 8392 3709 8456
rect 3773 8392 3789 8456
rect 3853 8392 3861 8456
rect 3541 8391 3861 8392
rect 6138 8456 6458 8457
rect 6138 8392 6146 8456
rect 6210 8392 6226 8456
rect 6290 8392 6306 8456
rect 6370 8392 6386 8456
rect 6450 8392 6458 8456
rect 6138 8391 6458 8392
rect 3325 8386 3391 8389
rect 0 8384 3391 8386
rect 0 8328 3330 8384
rect 3386 8328 3391 8384
rect 0 8326 3391 8328
rect 0 8296 480 8326
rect 3325 8323 3391 8326
rect 2242 7912 2562 7913
rect 2242 7848 2250 7912
rect 2314 7848 2330 7912
rect 2394 7848 2410 7912
rect 2474 7848 2490 7912
rect 2554 7848 2562 7912
rect 2242 7847 2562 7848
rect 4840 7912 5160 7913
rect 4840 7848 4848 7912
rect 4912 7848 4928 7912
rect 4992 7848 5008 7912
rect 5072 7848 5088 7912
rect 5152 7848 5160 7912
rect 4840 7847 5160 7848
rect 7437 7912 7757 7913
rect 7437 7848 7445 7912
rect 7509 7848 7525 7912
rect 7589 7848 7605 7912
rect 7669 7848 7685 7912
rect 7749 7848 7757 7912
rect 7437 7847 7757 7848
rect 3541 7368 3861 7369
rect 3541 7304 3549 7368
rect 3613 7304 3629 7368
rect 3693 7304 3709 7368
rect 3773 7304 3789 7368
rect 3853 7304 3861 7368
rect 3541 7303 3861 7304
rect 6138 7368 6458 7369
rect 6138 7304 6146 7368
rect 6210 7304 6226 7368
rect 6290 7304 6306 7368
rect 6370 7304 6386 7368
rect 6450 7304 6458 7368
rect 6138 7303 6458 7304
rect 4061 7026 4127 7029
rect 2086 7024 4127 7026
rect 2086 6968 4066 7024
rect 4122 6968 4127 7024
rect 2086 6966 4127 6968
rect 0 6754 480 6784
rect 2086 6754 2146 6966
rect 4061 6963 4127 6966
rect 2242 6824 2562 6825
rect 2242 6760 2250 6824
rect 2314 6760 2330 6824
rect 2394 6760 2410 6824
rect 2474 6760 2490 6824
rect 2554 6760 2562 6824
rect 2242 6759 2562 6760
rect 4840 6824 5160 6825
rect 4840 6760 4848 6824
rect 4912 6760 4928 6824
rect 4992 6760 5008 6824
rect 5072 6760 5088 6824
rect 5152 6760 5160 6824
rect 4840 6759 5160 6760
rect 7437 6824 7757 6825
rect 7437 6760 7445 6824
rect 7509 6760 7525 6824
rect 7589 6760 7605 6824
rect 7669 6760 7685 6824
rect 7749 6760 7757 6824
rect 7437 6759 7757 6760
rect 0 6694 2146 6754
rect 0 6664 480 6694
rect 3541 6280 3861 6281
rect 3541 6216 3549 6280
rect 3613 6216 3629 6280
rect 3693 6216 3709 6280
rect 3773 6216 3789 6280
rect 3853 6216 3861 6280
rect 3541 6215 3861 6216
rect 6138 6280 6458 6281
rect 6138 6216 6146 6280
rect 6210 6216 6226 6280
rect 6290 6216 6306 6280
rect 6370 6216 6386 6280
rect 6450 6216 6458 6280
rect 6138 6215 6458 6216
rect 5625 6074 5691 6077
rect 9520 6074 10000 6104
rect 5625 6072 10000 6074
rect 5625 6016 5630 6072
rect 5686 6016 10000 6072
rect 5625 6014 10000 6016
rect 5625 6011 5691 6014
rect 9520 5984 10000 6014
rect 2242 5736 2562 5737
rect 2242 5672 2250 5736
rect 2314 5672 2330 5736
rect 2394 5672 2410 5736
rect 2474 5672 2490 5736
rect 2554 5672 2562 5736
rect 2242 5671 2562 5672
rect 4840 5736 5160 5737
rect 4840 5672 4848 5736
rect 4912 5672 4928 5736
rect 4992 5672 5008 5736
rect 5072 5672 5088 5736
rect 5152 5672 5160 5736
rect 4840 5671 5160 5672
rect 7437 5736 7757 5737
rect 7437 5672 7445 5736
rect 7509 5672 7525 5736
rect 7589 5672 7605 5736
rect 7669 5672 7685 5736
rect 7749 5672 7757 5736
rect 7437 5671 7757 5672
rect 3541 5192 3861 5193
rect 3541 5128 3549 5192
rect 3613 5128 3629 5192
rect 3693 5128 3709 5192
rect 3773 5128 3789 5192
rect 3853 5128 3861 5192
rect 3541 5127 3861 5128
rect 6138 5192 6458 5193
rect 6138 5128 6146 5192
rect 6210 5128 6226 5192
rect 6290 5128 6306 5192
rect 6370 5128 6386 5192
rect 6450 5128 6458 5192
rect 6138 5127 6458 5128
rect 0 4986 480 5016
rect 3325 4986 3391 4989
rect 0 4984 3391 4986
rect 0 4928 3330 4984
rect 3386 4928 3391 4984
rect 0 4926 3391 4928
rect 0 4896 480 4926
rect 3325 4923 3391 4926
rect 2242 4648 2562 4649
rect 2242 4584 2250 4648
rect 2314 4584 2330 4648
rect 2394 4584 2410 4648
rect 2474 4584 2490 4648
rect 2554 4584 2562 4648
rect 2242 4583 2562 4584
rect 4840 4648 5160 4649
rect 4840 4584 4848 4648
rect 4912 4584 4928 4648
rect 4992 4584 5008 4648
rect 5072 4584 5088 4648
rect 5152 4584 5160 4648
rect 4840 4583 5160 4584
rect 7437 4648 7757 4649
rect 7437 4584 7445 4648
rect 7509 4584 7525 4648
rect 7589 4584 7605 4648
rect 7669 4584 7685 4648
rect 7749 4584 7757 4648
rect 7437 4583 7757 4584
rect 3541 4104 3861 4105
rect 3541 4040 3549 4104
rect 3613 4040 3629 4104
rect 3693 4040 3709 4104
rect 3773 4040 3789 4104
rect 3853 4040 3861 4104
rect 3541 4039 3861 4040
rect 6138 4104 6458 4105
rect 6138 4040 6146 4104
rect 6210 4040 6226 4104
rect 6290 4040 6306 4104
rect 6370 4040 6386 4104
rect 6450 4040 6458 4104
rect 6138 4039 6458 4040
rect 2242 3560 2562 3561
rect 2242 3496 2250 3560
rect 2314 3496 2330 3560
rect 2394 3496 2410 3560
rect 2474 3496 2490 3560
rect 2554 3496 2562 3560
rect 2242 3495 2562 3496
rect 4840 3560 5160 3561
rect 4840 3496 4848 3560
rect 4912 3496 4928 3560
rect 4992 3496 5008 3560
rect 5072 3496 5088 3560
rect 5152 3496 5160 3560
rect 4840 3495 5160 3496
rect 7437 3560 7757 3561
rect 7437 3496 7445 3560
rect 7509 3496 7525 3560
rect 7589 3496 7605 3560
rect 7669 3496 7685 3560
rect 7749 3496 7757 3560
rect 7437 3495 7757 3496
rect 0 3354 480 3384
rect 2865 3354 2931 3357
rect 0 3352 2931 3354
rect 0 3296 2870 3352
rect 2926 3296 2931 3352
rect 0 3294 2931 3296
rect 0 3264 480 3294
rect 2865 3291 2931 3294
rect 6637 3354 6703 3357
rect 9520 3354 10000 3384
rect 6637 3352 10000 3354
rect 6637 3296 6642 3352
rect 6698 3296 10000 3352
rect 6637 3294 10000 3296
rect 6637 3291 6703 3294
rect 9520 3264 10000 3294
rect 3541 3016 3861 3017
rect 3541 2952 3549 3016
rect 3613 2952 3629 3016
rect 3693 2952 3709 3016
rect 3773 2952 3789 3016
rect 3853 2952 3861 3016
rect 3541 2951 3861 2952
rect 6138 3016 6458 3017
rect 6138 2952 6146 3016
rect 6210 2952 6226 3016
rect 6290 2952 6306 3016
rect 6370 2952 6386 3016
rect 6450 2952 6458 3016
rect 6138 2951 6458 2952
rect 2242 2472 2562 2473
rect 2242 2408 2250 2472
rect 2314 2408 2330 2472
rect 2394 2408 2410 2472
rect 2474 2408 2490 2472
rect 2554 2408 2562 2472
rect 2242 2407 2562 2408
rect 4840 2472 5160 2473
rect 4840 2408 4848 2472
rect 4912 2408 4928 2472
rect 4992 2408 5008 2472
rect 5072 2408 5088 2472
rect 5152 2408 5160 2472
rect 4840 2407 5160 2408
rect 7437 2472 7757 2473
rect 7437 2408 7445 2472
rect 7509 2408 7525 2472
rect 7589 2408 7605 2472
rect 7669 2408 7685 2472
rect 7749 2408 7757 2472
rect 7437 2407 7757 2408
rect 3541 1928 3861 1929
rect 3541 1864 3549 1928
rect 3613 1864 3629 1928
rect 3693 1864 3709 1928
rect 3773 1864 3789 1928
rect 3853 1864 3861 1928
rect 3541 1863 3861 1864
rect 6138 1928 6458 1929
rect 6138 1864 6146 1928
rect 6210 1864 6226 1928
rect 6290 1864 6306 1928
rect 6370 1864 6386 1928
rect 6450 1864 6458 1928
rect 6138 1863 6458 1864
rect 0 1722 480 1752
rect 4061 1722 4127 1725
rect 0 1720 4127 1722
rect 0 1664 4066 1720
rect 4122 1664 4127 1720
rect 0 1662 4127 1664
rect 0 1632 480 1662
rect 4061 1659 4127 1662
rect 2242 1384 2562 1385
rect 2242 1320 2250 1384
rect 2314 1320 2330 1384
rect 2394 1320 2410 1384
rect 2474 1320 2490 1384
rect 2554 1320 2562 1384
rect 2242 1319 2562 1320
rect 4840 1384 5160 1385
rect 4840 1320 4848 1384
rect 4912 1320 4928 1384
rect 4992 1320 5008 1384
rect 5072 1320 5088 1384
rect 5152 1320 5160 1384
rect 4840 1319 5160 1320
rect 7437 1384 7757 1385
rect 7437 1320 7445 1384
rect 7509 1320 7525 1384
rect 7589 1320 7605 1384
rect 7669 1320 7685 1384
rect 7749 1320 7757 1384
rect 7437 1319 7757 1320
rect 6821 634 6887 637
rect 9520 634 10000 664
rect 6821 632 10000 634
rect 6821 576 6826 632
rect 6882 576 10000 632
rect 6821 574 10000 576
rect 6821 571 6887 574
rect 9520 544 10000 574
rect 0 90 480 120
rect 3417 90 3483 93
rect 0 88 3483 90
rect 0 32 3422 88
rect 3478 32 3483 88
rect 0 30 3483 32
rect 0 0 480 30
rect 3417 27 3483 30
<< via3 >>
rect 3549 21508 3613 21512
rect 3549 21452 3553 21508
rect 3553 21452 3609 21508
rect 3609 21452 3613 21508
rect 3549 21448 3613 21452
rect 3629 21508 3693 21512
rect 3629 21452 3633 21508
rect 3633 21452 3689 21508
rect 3689 21452 3693 21508
rect 3629 21448 3693 21452
rect 3709 21508 3773 21512
rect 3709 21452 3713 21508
rect 3713 21452 3769 21508
rect 3769 21452 3773 21508
rect 3709 21448 3773 21452
rect 3789 21508 3853 21512
rect 3789 21452 3793 21508
rect 3793 21452 3849 21508
rect 3849 21452 3853 21508
rect 3789 21448 3853 21452
rect 6146 21508 6210 21512
rect 6146 21452 6150 21508
rect 6150 21452 6206 21508
rect 6206 21452 6210 21508
rect 6146 21448 6210 21452
rect 6226 21508 6290 21512
rect 6226 21452 6230 21508
rect 6230 21452 6286 21508
rect 6286 21452 6290 21508
rect 6226 21448 6290 21452
rect 6306 21508 6370 21512
rect 6306 21452 6310 21508
rect 6310 21452 6366 21508
rect 6366 21452 6370 21508
rect 6306 21448 6370 21452
rect 6386 21508 6450 21512
rect 6386 21452 6390 21508
rect 6390 21452 6446 21508
rect 6446 21452 6450 21508
rect 6386 21448 6450 21452
rect 2250 20964 2314 20968
rect 2250 20908 2254 20964
rect 2254 20908 2310 20964
rect 2310 20908 2314 20964
rect 2250 20904 2314 20908
rect 2330 20964 2394 20968
rect 2330 20908 2334 20964
rect 2334 20908 2390 20964
rect 2390 20908 2394 20964
rect 2330 20904 2394 20908
rect 2410 20964 2474 20968
rect 2410 20908 2414 20964
rect 2414 20908 2470 20964
rect 2470 20908 2474 20964
rect 2410 20904 2474 20908
rect 2490 20964 2554 20968
rect 2490 20908 2494 20964
rect 2494 20908 2550 20964
rect 2550 20908 2554 20964
rect 2490 20904 2554 20908
rect 4848 20964 4912 20968
rect 4848 20908 4852 20964
rect 4852 20908 4908 20964
rect 4908 20908 4912 20964
rect 4848 20904 4912 20908
rect 4928 20964 4992 20968
rect 4928 20908 4932 20964
rect 4932 20908 4988 20964
rect 4988 20908 4992 20964
rect 4928 20904 4992 20908
rect 5008 20964 5072 20968
rect 5008 20908 5012 20964
rect 5012 20908 5068 20964
rect 5068 20908 5072 20964
rect 5008 20904 5072 20908
rect 5088 20964 5152 20968
rect 5088 20908 5092 20964
rect 5092 20908 5148 20964
rect 5148 20908 5152 20964
rect 5088 20904 5152 20908
rect 7445 20964 7509 20968
rect 7445 20908 7449 20964
rect 7449 20908 7505 20964
rect 7505 20908 7509 20964
rect 7445 20904 7509 20908
rect 7525 20964 7589 20968
rect 7525 20908 7529 20964
rect 7529 20908 7585 20964
rect 7585 20908 7589 20964
rect 7525 20904 7589 20908
rect 7605 20964 7669 20968
rect 7605 20908 7609 20964
rect 7609 20908 7665 20964
rect 7665 20908 7669 20964
rect 7605 20904 7669 20908
rect 7685 20964 7749 20968
rect 7685 20908 7689 20964
rect 7689 20908 7745 20964
rect 7745 20908 7749 20964
rect 7685 20904 7749 20908
rect 3549 20420 3613 20424
rect 3549 20364 3553 20420
rect 3553 20364 3609 20420
rect 3609 20364 3613 20420
rect 3549 20360 3613 20364
rect 3629 20420 3693 20424
rect 3629 20364 3633 20420
rect 3633 20364 3689 20420
rect 3689 20364 3693 20420
rect 3629 20360 3693 20364
rect 3709 20420 3773 20424
rect 3709 20364 3713 20420
rect 3713 20364 3769 20420
rect 3769 20364 3773 20420
rect 3709 20360 3773 20364
rect 3789 20420 3853 20424
rect 3789 20364 3793 20420
rect 3793 20364 3849 20420
rect 3849 20364 3853 20420
rect 3789 20360 3853 20364
rect 6146 20420 6210 20424
rect 6146 20364 6150 20420
rect 6150 20364 6206 20420
rect 6206 20364 6210 20420
rect 6146 20360 6210 20364
rect 6226 20420 6290 20424
rect 6226 20364 6230 20420
rect 6230 20364 6286 20420
rect 6286 20364 6290 20420
rect 6226 20360 6290 20364
rect 6306 20420 6370 20424
rect 6306 20364 6310 20420
rect 6310 20364 6366 20420
rect 6366 20364 6370 20420
rect 6306 20360 6370 20364
rect 6386 20420 6450 20424
rect 6386 20364 6390 20420
rect 6390 20364 6446 20420
rect 6446 20364 6450 20420
rect 6386 20360 6450 20364
rect 2250 19876 2314 19880
rect 2250 19820 2254 19876
rect 2254 19820 2310 19876
rect 2310 19820 2314 19876
rect 2250 19816 2314 19820
rect 2330 19876 2394 19880
rect 2330 19820 2334 19876
rect 2334 19820 2390 19876
rect 2390 19820 2394 19876
rect 2330 19816 2394 19820
rect 2410 19876 2474 19880
rect 2410 19820 2414 19876
rect 2414 19820 2470 19876
rect 2470 19820 2474 19876
rect 2410 19816 2474 19820
rect 2490 19876 2554 19880
rect 2490 19820 2494 19876
rect 2494 19820 2550 19876
rect 2550 19820 2554 19876
rect 2490 19816 2554 19820
rect 4848 19876 4912 19880
rect 4848 19820 4852 19876
rect 4852 19820 4908 19876
rect 4908 19820 4912 19876
rect 4848 19816 4912 19820
rect 4928 19876 4992 19880
rect 4928 19820 4932 19876
rect 4932 19820 4988 19876
rect 4988 19820 4992 19876
rect 4928 19816 4992 19820
rect 5008 19876 5072 19880
rect 5008 19820 5012 19876
rect 5012 19820 5068 19876
rect 5068 19820 5072 19876
rect 5008 19816 5072 19820
rect 5088 19876 5152 19880
rect 5088 19820 5092 19876
rect 5092 19820 5148 19876
rect 5148 19820 5152 19876
rect 5088 19816 5152 19820
rect 7445 19876 7509 19880
rect 7445 19820 7449 19876
rect 7449 19820 7505 19876
rect 7505 19820 7509 19876
rect 7445 19816 7509 19820
rect 7525 19876 7589 19880
rect 7525 19820 7529 19876
rect 7529 19820 7585 19876
rect 7585 19820 7589 19876
rect 7525 19816 7589 19820
rect 7605 19876 7669 19880
rect 7605 19820 7609 19876
rect 7609 19820 7665 19876
rect 7665 19820 7669 19876
rect 7605 19816 7669 19820
rect 7685 19876 7749 19880
rect 7685 19820 7689 19876
rect 7689 19820 7745 19876
rect 7745 19820 7749 19876
rect 7685 19816 7749 19820
rect 3549 19332 3613 19336
rect 3549 19276 3553 19332
rect 3553 19276 3609 19332
rect 3609 19276 3613 19332
rect 3549 19272 3613 19276
rect 3629 19332 3693 19336
rect 3629 19276 3633 19332
rect 3633 19276 3689 19332
rect 3689 19276 3693 19332
rect 3629 19272 3693 19276
rect 3709 19332 3773 19336
rect 3709 19276 3713 19332
rect 3713 19276 3769 19332
rect 3769 19276 3773 19332
rect 3709 19272 3773 19276
rect 3789 19332 3853 19336
rect 3789 19276 3793 19332
rect 3793 19276 3849 19332
rect 3849 19276 3853 19332
rect 3789 19272 3853 19276
rect 6146 19332 6210 19336
rect 6146 19276 6150 19332
rect 6150 19276 6206 19332
rect 6206 19276 6210 19332
rect 6146 19272 6210 19276
rect 6226 19332 6290 19336
rect 6226 19276 6230 19332
rect 6230 19276 6286 19332
rect 6286 19276 6290 19332
rect 6226 19272 6290 19276
rect 6306 19332 6370 19336
rect 6306 19276 6310 19332
rect 6310 19276 6366 19332
rect 6366 19276 6370 19332
rect 6306 19272 6370 19276
rect 6386 19332 6450 19336
rect 6386 19276 6390 19332
rect 6390 19276 6446 19332
rect 6446 19276 6450 19332
rect 6386 19272 6450 19276
rect 2250 18788 2314 18792
rect 2250 18732 2254 18788
rect 2254 18732 2310 18788
rect 2310 18732 2314 18788
rect 2250 18728 2314 18732
rect 2330 18788 2394 18792
rect 2330 18732 2334 18788
rect 2334 18732 2390 18788
rect 2390 18732 2394 18788
rect 2330 18728 2394 18732
rect 2410 18788 2474 18792
rect 2410 18732 2414 18788
rect 2414 18732 2470 18788
rect 2470 18732 2474 18788
rect 2410 18728 2474 18732
rect 2490 18788 2554 18792
rect 2490 18732 2494 18788
rect 2494 18732 2550 18788
rect 2550 18732 2554 18788
rect 2490 18728 2554 18732
rect 4848 18788 4912 18792
rect 4848 18732 4852 18788
rect 4852 18732 4908 18788
rect 4908 18732 4912 18788
rect 4848 18728 4912 18732
rect 4928 18788 4992 18792
rect 4928 18732 4932 18788
rect 4932 18732 4988 18788
rect 4988 18732 4992 18788
rect 4928 18728 4992 18732
rect 5008 18788 5072 18792
rect 5008 18732 5012 18788
rect 5012 18732 5068 18788
rect 5068 18732 5072 18788
rect 5008 18728 5072 18732
rect 5088 18788 5152 18792
rect 5088 18732 5092 18788
rect 5092 18732 5148 18788
rect 5148 18732 5152 18788
rect 5088 18728 5152 18732
rect 7445 18788 7509 18792
rect 7445 18732 7449 18788
rect 7449 18732 7505 18788
rect 7505 18732 7509 18788
rect 7445 18728 7509 18732
rect 7525 18788 7589 18792
rect 7525 18732 7529 18788
rect 7529 18732 7585 18788
rect 7585 18732 7589 18788
rect 7525 18728 7589 18732
rect 7605 18788 7669 18792
rect 7605 18732 7609 18788
rect 7609 18732 7665 18788
rect 7665 18732 7669 18788
rect 7605 18728 7669 18732
rect 7685 18788 7749 18792
rect 7685 18732 7689 18788
rect 7689 18732 7745 18788
rect 7745 18732 7749 18788
rect 7685 18728 7749 18732
rect 3549 18244 3613 18248
rect 3549 18188 3553 18244
rect 3553 18188 3609 18244
rect 3609 18188 3613 18244
rect 3549 18184 3613 18188
rect 3629 18244 3693 18248
rect 3629 18188 3633 18244
rect 3633 18188 3689 18244
rect 3689 18188 3693 18244
rect 3629 18184 3693 18188
rect 3709 18244 3773 18248
rect 3709 18188 3713 18244
rect 3713 18188 3769 18244
rect 3769 18188 3773 18244
rect 3709 18184 3773 18188
rect 3789 18244 3853 18248
rect 3789 18188 3793 18244
rect 3793 18188 3849 18244
rect 3849 18188 3853 18244
rect 3789 18184 3853 18188
rect 6146 18244 6210 18248
rect 6146 18188 6150 18244
rect 6150 18188 6206 18244
rect 6206 18188 6210 18244
rect 6146 18184 6210 18188
rect 6226 18244 6290 18248
rect 6226 18188 6230 18244
rect 6230 18188 6286 18244
rect 6286 18188 6290 18244
rect 6226 18184 6290 18188
rect 6306 18244 6370 18248
rect 6306 18188 6310 18244
rect 6310 18188 6366 18244
rect 6366 18188 6370 18244
rect 6306 18184 6370 18188
rect 6386 18244 6450 18248
rect 6386 18188 6390 18244
rect 6390 18188 6446 18244
rect 6446 18188 6450 18244
rect 6386 18184 6450 18188
rect 2250 17700 2314 17704
rect 2250 17644 2254 17700
rect 2254 17644 2310 17700
rect 2310 17644 2314 17700
rect 2250 17640 2314 17644
rect 2330 17700 2394 17704
rect 2330 17644 2334 17700
rect 2334 17644 2390 17700
rect 2390 17644 2394 17700
rect 2330 17640 2394 17644
rect 2410 17700 2474 17704
rect 2410 17644 2414 17700
rect 2414 17644 2470 17700
rect 2470 17644 2474 17700
rect 2410 17640 2474 17644
rect 2490 17700 2554 17704
rect 2490 17644 2494 17700
rect 2494 17644 2550 17700
rect 2550 17644 2554 17700
rect 2490 17640 2554 17644
rect 4848 17700 4912 17704
rect 4848 17644 4852 17700
rect 4852 17644 4908 17700
rect 4908 17644 4912 17700
rect 4848 17640 4912 17644
rect 4928 17700 4992 17704
rect 4928 17644 4932 17700
rect 4932 17644 4988 17700
rect 4988 17644 4992 17700
rect 4928 17640 4992 17644
rect 5008 17700 5072 17704
rect 5008 17644 5012 17700
rect 5012 17644 5068 17700
rect 5068 17644 5072 17700
rect 5008 17640 5072 17644
rect 5088 17700 5152 17704
rect 5088 17644 5092 17700
rect 5092 17644 5148 17700
rect 5148 17644 5152 17700
rect 5088 17640 5152 17644
rect 7445 17700 7509 17704
rect 7445 17644 7449 17700
rect 7449 17644 7505 17700
rect 7505 17644 7509 17700
rect 7445 17640 7509 17644
rect 7525 17700 7589 17704
rect 7525 17644 7529 17700
rect 7529 17644 7585 17700
rect 7585 17644 7589 17700
rect 7525 17640 7589 17644
rect 7605 17700 7669 17704
rect 7605 17644 7609 17700
rect 7609 17644 7665 17700
rect 7665 17644 7669 17700
rect 7605 17640 7669 17644
rect 7685 17700 7749 17704
rect 7685 17644 7689 17700
rect 7689 17644 7745 17700
rect 7745 17644 7749 17700
rect 7685 17640 7749 17644
rect 3549 17156 3613 17160
rect 3549 17100 3553 17156
rect 3553 17100 3609 17156
rect 3609 17100 3613 17156
rect 3549 17096 3613 17100
rect 3629 17156 3693 17160
rect 3629 17100 3633 17156
rect 3633 17100 3689 17156
rect 3689 17100 3693 17156
rect 3629 17096 3693 17100
rect 3709 17156 3773 17160
rect 3709 17100 3713 17156
rect 3713 17100 3769 17156
rect 3769 17100 3773 17156
rect 3709 17096 3773 17100
rect 3789 17156 3853 17160
rect 3789 17100 3793 17156
rect 3793 17100 3849 17156
rect 3849 17100 3853 17156
rect 3789 17096 3853 17100
rect 6146 17156 6210 17160
rect 6146 17100 6150 17156
rect 6150 17100 6206 17156
rect 6206 17100 6210 17156
rect 6146 17096 6210 17100
rect 6226 17156 6290 17160
rect 6226 17100 6230 17156
rect 6230 17100 6286 17156
rect 6286 17100 6290 17156
rect 6226 17096 6290 17100
rect 6306 17156 6370 17160
rect 6306 17100 6310 17156
rect 6310 17100 6366 17156
rect 6366 17100 6370 17156
rect 6306 17096 6370 17100
rect 6386 17156 6450 17160
rect 6386 17100 6390 17156
rect 6390 17100 6446 17156
rect 6446 17100 6450 17156
rect 6386 17096 6450 17100
rect 2250 16612 2314 16616
rect 2250 16556 2254 16612
rect 2254 16556 2310 16612
rect 2310 16556 2314 16612
rect 2250 16552 2314 16556
rect 2330 16612 2394 16616
rect 2330 16556 2334 16612
rect 2334 16556 2390 16612
rect 2390 16556 2394 16612
rect 2330 16552 2394 16556
rect 2410 16612 2474 16616
rect 2410 16556 2414 16612
rect 2414 16556 2470 16612
rect 2470 16556 2474 16612
rect 2410 16552 2474 16556
rect 2490 16612 2554 16616
rect 2490 16556 2494 16612
rect 2494 16556 2550 16612
rect 2550 16556 2554 16612
rect 2490 16552 2554 16556
rect 4848 16612 4912 16616
rect 4848 16556 4852 16612
rect 4852 16556 4908 16612
rect 4908 16556 4912 16612
rect 4848 16552 4912 16556
rect 4928 16612 4992 16616
rect 4928 16556 4932 16612
rect 4932 16556 4988 16612
rect 4988 16556 4992 16612
rect 4928 16552 4992 16556
rect 5008 16612 5072 16616
rect 5008 16556 5012 16612
rect 5012 16556 5068 16612
rect 5068 16556 5072 16612
rect 5008 16552 5072 16556
rect 5088 16612 5152 16616
rect 5088 16556 5092 16612
rect 5092 16556 5148 16612
rect 5148 16556 5152 16612
rect 5088 16552 5152 16556
rect 7445 16612 7509 16616
rect 7445 16556 7449 16612
rect 7449 16556 7505 16612
rect 7505 16556 7509 16612
rect 7445 16552 7509 16556
rect 7525 16612 7589 16616
rect 7525 16556 7529 16612
rect 7529 16556 7585 16612
rect 7585 16556 7589 16612
rect 7525 16552 7589 16556
rect 7605 16612 7669 16616
rect 7605 16556 7609 16612
rect 7609 16556 7665 16612
rect 7665 16556 7669 16612
rect 7605 16552 7669 16556
rect 7685 16612 7749 16616
rect 7685 16556 7689 16612
rect 7689 16556 7745 16612
rect 7745 16556 7749 16612
rect 7685 16552 7749 16556
rect 3549 16068 3613 16072
rect 3549 16012 3553 16068
rect 3553 16012 3609 16068
rect 3609 16012 3613 16068
rect 3549 16008 3613 16012
rect 3629 16068 3693 16072
rect 3629 16012 3633 16068
rect 3633 16012 3689 16068
rect 3689 16012 3693 16068
rect 3629 16008 3693 16012
rect 3709 16068 3773 16072
rect 3709 16012 3713 16068
rect 3713 16012 3769 16068
rect 3769 16012 3773 16068
rect 3709 16008 3773 16012
rect 3789 16068 3853 16072
rect 3789 16012 3793 16068
rect 3793 16012 3849 16068
rect 3849 16012 3853 16068
rect 3789 16008 3853 16012
rect 6146 16068 6210 16072
rect 6146 16012 6150 16068
rect 6150 16012 6206 16068
rect 6206 16012 6210 16068
rect 6146 16008 6210 16012
rect 6226 16068 6290 16072
rect 6226 16012 6230 16068
rect 6230 16012 6286 16068
rect 6286 16012 6290 16068
rect 6226 16008 6290 16012
rect 6306 16068 6370 16072
rect 6306 16012 6310 16068
rect 6310 16012 6366 16068
rect 6366 16012 6370 16068
rect 6306 16008 6370 16012
rect 6386 16068 6450 16072
rect 6386 16012 6390 16068
rect 6390 16012 6446 16068
rect 6446 16012 6450 16068
rect 6386 16008 6450 16012
rect 2250 15524 2314 15528
rect 2250 15468 2254 15524
rect 2254 15468 2310 15524
rect 2310 15468 2314 15524
rect 2250 15464 2314 15468
rect 2330 15524 2394 15528
rect 2330 15468 2334 15524
rect 2334 15468 2390 15524
rect 2390 15468 2394 15524
rect 2330 15464 2394 15468
rect 2410 15524 2474 15528
rect 2410 15468 2414 15524
rect 2414 15468 2470 15524
rect 2470 15468 2474 15524
rect 2410 15464 2474 15468
rect 2490 15524 2554 15528
rect 2490 15468 2494 15524
rect 2494 15468 2550 15524
rect 2550 15468 2554 15524
rect 2490 15464 2554 15468
rect 4848 15524 4912 15528
rect 4848 15468 4852 15524
rect 4852 15468 4908 15524
rect 4908 15468 4912 15524
rect 4848 15464 4912 15468
rect 4928 15524 4992 15528
rect 4928 15468 4932 15524
rect 4932 15468 4988 15524
rect 4988 15468 4992 15524
rect 4928 15464 4992 15468
rect 5008 15524 5072 15528
rect 5008 15468 5012 15524
rect 5012 15468 5068 15524
rect 5068 15468 5072 15524
rect 5008 15464 5072 15468
rect 5088 15524 5152 15528
rect 5088 15468 5092 15524
rect 5092 15468 5148 15524
rect 5148 15468 5152 15524
rect 5088 15464 5152 15468
rect 7445 15524 7509 15528
rect 7445 15468 7449 15524
rect 7449 15468 7505 15524
rect 7505 15468 7509 15524
rect 7445 15464 7509 15468
rect 7525 15524 7589 15528
rect 7525 15468 7529 15524
rect 7529 15468 7585 15524
rect 7585 15468 7589 15524
rect 7525 15464 7589 15468
rect 7605 15524 7669 15528
rect 7605 15468 7609 15524
rect 7609 15468 7665 15524
rect 7665 15468 7669 15524
rect 7605 15464 7669 15468
rect 7685 15524 7749 15528
rect 7685 15468 7689 15524
rect 7689 15468 7745 15524
rect 7745 15468 7749 15524
rect 7685 15464 7749 15468
rect 3549 14980 3613 14984
rect 3549 14924 3553 14980
rect 3553 14924 3609 14980
rect 3609 14924 3613 14980
rect 3549 14920 3613 14924
rect 3629 14980 3693 14984
rect 3629 14924 3633 14980
rect 3633 14924 3689 14980
rect 3689 14924 3693 14980
rect 3629 14920 3693 14924
rect 3709 14980 3773 14984
rect 3709 14924 3713 14980
rect 3713 14924 3769 14980
rect 3769 14924 3773 14980
rect 3709 14920 3773 14924
rect 3789 14980 3853 14984
rect 3789 14924 3793 14980
rect 3793 14924 3849 14980
rect 3849 14924 3853 14980
rect 3789 14920 3853 14924
rect 6146 14980 6210 14984
rect 6146 14924 6150 14980
rect 6150 14924 6206 14980
rect 6206 14924 6210 14980
rect 6146 14920 6210 14924
rect 6226 14980 6290 14984
rect 6226 14924 6230 14980
rect 6230 14924 6286 14980
rect 6286 14924 6290 14980
rect 6226 14920 6290 14924
rect 6306 14980 6370 14984
rect 6306 14924 6310 14980
rect 6310 14924 6366 14980
rect 6366 14924 6370 14980
rect 6306 14920 6370 14924
rect 6386 14980 6450 14984
rect 6386 14924 6390 14980
rect 6390 14924 6446 14980
rect 6446 14924 6450 14980
rect 6386 14920 6450 14924
rect 2250 14436 2314 14440
rect 2250 14380 2254 14436
rect 2254 14380 2310 14436
rect 2310 14380 2314 14436
rect 2250 14376 2314 14380
rect 2330 14436 2394 14440
rect 2330 14380 2334 14436
rect 2334 14380 2390 14436
rect 2390 14380 2394 14436
rect 2330 14376 2394 14380
rect 2410 14436 2474 14440
rect 2410 14380 2414 14436
rect 2414 14380 2470 14436
rect 2470 14380 2474 14436
rect 2410 14376 2474 14380
rect 2490 14436 2554 14440
rect 2490 14380 2494 14436
rect 2494 14380 2550 14436
rect 2550 14380 2554 14436
rect 2490 14376 2554 14380
rect 4848 14436 4912 14440
rect 4848 14380 4852 14436
rect 4852 14380 4908 14436
rect 4908 14380 4912 14436
rect 4848 14376 4912 14380
rect 4928 14436 4992 14440
rect 4928 14380 4932 14436
rect 4932 14380 4988 14436
rect 4988 14380 4992 14436
rect 4928 14376 4992 14380
rect 5008 14436 5072 14440
rect 5008 14380 5012 14436
rect 5012 14380 5068 14436
rect 5068 14380 5072 14436
rect 5008 14376 5072 14380
rect 5088 14436 5152 14440
rect 5088 14380 5092 14436
rect 5092 14380 5148 14436
rect 5148 14380 5152 14436
rect 5088 14376 5152 14380
rect 7445 14436 7509 14440
rect 7445 14380 7449 14436
rect 7449 14380 7505 14436
rect 7505 14380 7509 14436
rect 7445 14376 7509 14380
rect 7525 14436 7589 14440
rect 7525 14380 7529 14436
rect 7529 14380 7585 14436
rect 7585 14380 7589 14436
rect 7525 14376 7589 14380
rect 7605 14436 7669 14440
rect 7605 14380 7609 14436
rect 7609 14380 7665 14436
rect 7665 14380 7669 14436
rect 7605 14376 7669 14380
rect 7685 14436 7749 14440
rect 7685 14380 7689 14436
rect 7689 14380 7745 14436
rect 7745 14380 7749 14436
rect 7685 14376 7749 14380
rect 3549 13892 3613 13896
rect 3549 13836 3553 13892
rect 3553 13836 3609 13892
rect 3609 13836 3613 13892
rect 3549 13832 3613 13836
rect 3629 13892 3693 13896
rect 3629 13836 3633 13892
rect 3633 13836 3689 13892
rect 3689 13836 3693 13892
rect 3629 13832 3693 13836
rect 3709 13892 3773 13896
rect 3709 13836 3713 13892
rect 3713 13836 3769 13892
rect 3769 13836 3773 13892
rect 3709 13832 3773 13836
rect 3789 13892 3853 13896
rect 3789 13836 3793 13892
rect 3793 13836 3849 13892
rect 3849 13836 3853 13892
rect 3789 13832 3853 13836
rect 6146 13892 6210 13896
rect 6146 13836 6150 13892
rect 6150 13836 6206 13892
rect 6206 13836 6210 13892
rect 6146 13832 6210 13836
rect 6226 13892 6290 13896
rect 6226 13836 6230 13892
rect 6230 13836 6286 13892
rect 6286 13836 6290 13892
rect 6226 13832 6290 13836
rect 6306 13892 6370 13896
rect 6306 13836 6310 13892
rect 6310 13836 6366 13892
rect 6366 13836 6370 13892
rect 6306 13832 6370 13836
rect 6386 13892 6450 13896
rect 6386 13836 6390 13892
rect 6390 13836 6446 13892
rect 6446 13836 6450 13892
rect 6386 13832 6450 13836
rect 2250 13348 2314 13352
rect 2250 13292 2254 13348
rect 2254 13292 2310 13348
rect 2310 13292 2314 13348
rect 2250 13288 2314 13292
rect 2330 13348 2394 13352
rect 2330 13292 2334 13348
rect 2334 13292 2390 13348
rect 2390 13292 2394 13348
rect 2330 13288 2394 13292
rect 2410 13348 2474 13352
rect 2410 13292 2414 13348
rect 2414 13292 2470 13348
rect 2470 13292 2474 13348
rect 2410 13288 2474 13292
rect 2490 13348 2554 13352
rect 2490 13292 2494 13348
rect 2494 13292 2550 13348
rect 2550 13292 2554 13348
rect 2490 13288 2554 13292
rect 4848 13348 4912 13352
rect 4848 13292 4852 13348
rect 4852 13292 4908 13348
rect 4908 13292 4912 13348
rect 4848 13288 4912 13292
rect 4928 13348 4992 13352
rect 4928 13292 4932 13348
rect 4932 13292 4988 13348
rect 4988 13292 4992 13348
rect 4928 13288 4992 13292
rect 5008 13348 5072 13352
rect 5008 13292 5012 13348
rect 5012 13292 5068 13348
rect 5068 13292 5072 13348
rect 5008 13288 5072 13292
rect 5088 13348 5152 13352
rect 5088 13292 5092 13348
rect 5092 13292 5148 13348
rect 5148 13292 5152 13348
rect 5088 13288 5152 13292
rect 7445 13348 7509 13352
rect 7445 13292 7449 13348
rect 7449 13292 7505 13348
rect 7505 13292 7509 13348
rect 7445 13288 7509 13292
rect 7525 13348 7589 13352
rect 7525 13292 7529 13348
rect 7529 13292 7585 13348
rect 7585 13292 7589 13348
rect 7525 13288 7589 13292
rect 7605 13348 7669 13352
rect 7605 13292 7609 13348
rect 7609 13292 7665 13348
rect 7665 13292 7669 13348
rect 7605 13288 7669 13292
rect 7685 13348 7749 13352
rect 7685 13292 7689 13348
rect 7689 13292 7745 13348
rect 7745 13292 7749 13348
rect 7685 13288 7749 13292
rect 3549 12804 3613 12808
rect 3549 12748 3553 12804
rect 3553 12748 3609 12804
rect 3609 12748 3613 12804
rect 3549 12744 3613 12748
rect 3629 12804 3693 12808
rect 3629 12748 3633 12804
rect 3633 12748 3689 12804
rect 3689 12748 3693 12804
rect 3629 12744 3693 12748
rect 3709 12804 3773 12808
rect 3709 12748 3713 12804
rect 3713 12748 3769 12804
rect 3769 12748 3773 12804
rect 3709 12744 3773 12748
rect 3789 12804 3853 12808
rect 3789 12748 3793 12804
rect 3793 12748 3849 12804
rect 3849 12748 3853 12804
rect 3789 12744 3853 12748
rect 6146 12804 6210 12808
rect 6146 12748 6150 12804
rect 6150 12748 6206 12804
rect 6206 12748 6210 12804
rect 6146 12744 6210 12748
rect 6226 12804 6290 12808
rect 6226 12748 6230 12804
rect 6230 12748 6286 12804
rect 6286 12748 6290 12804
rect 6226 12744 6290 12748
rect 6306 12804 6370 12808
rect 6306 12748 6310 12804
rect 6310 12748 6366 12804
rect 6366 12748 6370 12804
rect 6306 12744 6370 12748
rect 6386 12804 6450 12808
rect 6386 12748 6390 12804
rect 6390 12748 6446 12804
rect 6446 12748 6450 12804
rect 6386 12744 6450 12748
rect 2250 12260 2314 12264
rect 2250 12204 2254 12260
rect 2254 12204 2310 12260
rect 2310 12204 2314 12260
rect 2250 12200 2314 12204
rect 2330 12260 2394 12264
rect 2330 12204 2334 12260
rect 2334 12204 2390 12260
rect 2390 12204 2394 12260
rect 2330 12200 2394 12204
rect 2410 12260 2474 12264
rect 2410 12204 2414 12260
rect 2414 12204 2470 12260
rect 2470 12204 2474 12260
rect 2410 12200 2474 12204
rect 2490 12260 2554 12264
rect 2490 12204 2494 12260
rect 2494 12204 2550 12260
rect 2550 12204 2554 12260
rect 2490 12200 2554 12204
rect 4848 12260 4912 12264
rect 4848 12204 4852 12260
rect 4852 12204 4908 12260
rect 4908 12204 4912 12260
rect 4848 12200 4912 12204
rect 4928 12260 4992 12264
rect 4928 12204 4932 12260
rect 4932 12204 4988 12260
rect 4988 12204 4992 12260
rect 4928 12200 4992 12204
rect 5008 12260 5072 12264
rect 5008 12204 5012 12260
rect 5012 12204 5068 12260
rect 5068 12204 5072 12260
rect 5008 12200 5072 12204
rect 5088 12260 5152 12264
rect 5088 12204 5092 12260
rect 5092 12204 5148 12260
rect 5148 12204 5152 12260
rect 5088 12200 5152 12204
rect 7445 12260 7509 12264
rect 7445 12204 7449 12260
rect 7449 12204 7505 12260
rect 7505 12204 7509 12260
rect 7445 12200 7509 12204
rect 7525 12260 7589 12264
rect 7525 12204 7529 12260
rect 7529 12204 7585 12260
rect 7585 12204 7589 12260
rect 7525 12200 7589 12204
rect 7605 12260 7669 12264
rect 7605 12204 7609 12260
rect 7609 12204 7665 12260
rect 7665 12204 7669 12260
rect 7605 12200 7669 12204
rect 7685 12260 7749 12264
rect 7685 12204 7689 12260
rect 7689 12204 7745 12260
rect 7745 12204 7749 12260
rect 7685 12200 7749 12204
rect 3549 11716 3613 11720
rect 3549 11660 3553 11716
rect 3553 11660 3609 11716
rect 3609 11660 3613 11716
rect 3549 11656 3613 11660
rect 3629 11716 3693 11720
rect 3629 11660 3633 11716
rect 3633 11660 3689 11716
rect 3689 11660 3693 11716
rect 3629 11656 3693 11660
rect 3709 11716 3773 11720
rect 3709 11660 3713 11716
rect 3713 11660 3769 11716
rect 3769 11660 3773 11716
rect 3709 11656 3773 11660
rect 3789 11716 3853 11720
rect 3789 11660 3793 11716
rect 3793 11660 3849 11716
rect 3849 11660 3853 11716
rect 3789 11656 3853 11660
rect 6146 11716 6210 11720
rect 6146 11660 6150 11716
rect 6150 11660 6206 11716
rect 6206 11660 6210 11716
rect 6146 11656 6210 11660
rect 6226 11716 6290 11720
rect 6226 11660 6230 11716
rect 6230 11660 6286 11716
rect 6286 11660 6290 11716
rect 6226 11656 6290 11660
rect 6306 11716 6370 11720
rect 6306 11660 6310 11716
rect 6310 11660 6366 11716
rect 6366 11660 6370 11716
rect 6306 11656 6370 11660
rect 6386 11716 6450 11720
rect 6386 11660 6390 11716
rect 6390 11660 6446 11716
rect 6446 11660 6450 11716
rect 6386 11656 6450 11660
rect 2250 11172 2314 11176
rect 2250 11116 2254 11172
rect 2254 11116 2310 11172
rect 2310 11116 2314 11172
rect 2250 11112 2314 11116
rect 2330 11172 2394 11176
rect 2330 11116 2334 11172
rect 2334 11116 2390 11172
rect 2390 11116 2394 11172
rect 2330 11112 2394 11116
rect 2410 11172 2474 11176
rect 2410 11116 2414 11172
rect 2414 11116 2470 11172
rect 2470 11116 2474 11172
rect 2410 11112 2474 11116
rect 2490 11172 2554 11176
rect 2490 11116 2494 11172
rect 2494 11116 2550 11172
rect 2550 11116 2554 11172
rect 2490 11112 2554 11116
rect 4848 11172 4912 11176
rect 4848 11116 4852 11172
rect 4852 11116 4908 11172
rect 4908 11116 4912 11172
rect 4848 11112 4912 11116
rect 4928 11172 4992 11176
rect 4928 11116 4932 11172
rect 4932 11116 4988 11172
rect 4988 11116 4992 11172
rect 4928 11112 4992 11116
rect 5008 11172 5072 11176
rect 5008 11116 5012 11172
rect 5012 11116 5068 11172
rect 5068 11116 5072 11172
rect 5008 11112 5072 11116
rect 5088 11172 5152 11176
rect 5088 11116 5092 11172
rect 5092 11116 5148 11172
rect 5148 11116 5152 11172
rect 5088 11112 5152 11116
rect 7445 11172 7509 11176
rect 7445 11116 7449 11172
rect 7449 11116 7505 11172
rect 7505 11116 7509 11172
rect 7445 11112 7509 11116
rect 7525 11172 7589 11176
rect 7525 11116 7529 11172
rect 7529 11116 7585 11172
rect 7585 11116 7589 11172
rect 7525 11112 7589 11116
rect 7605 11172 7669 11176
rect 7605 11116 7609 11172
rect 7609 11116 7665 11172
rect 7665 11116 7669 11172
rect 7605 11112 7669 11116
rect 7685 11172 7749 11176
rect 7685 11116 7689 11172
rect 7689 11116 7745 11172
rect 7745 11116 7749 11172
rect 7685 11112 7749 11116
rect 3549 10628 3613 10632
rect 3549 10572 3553 10628
rect 3553 10572 3609 10628
rect 3609 10572 3613 10628
rect 3549 10568 3613 10572
rect 3629 10628 3693 10632
rect 3629 10572 3633 10628
rect 3633 10572 3689 10628
rect 3689 10572 3693 10628
rect 3629 10568 3693 10572
rect 3709 10628 3773 10632
rect 3709 10572 3713 10628
rect 3713 10572 3769 10628
rect 3769 10572 3773 10628
rect 3709 10568 3773 10572
rect 3789 10628 3853 10632
rect 3789 10572 3793 10628
rect 3793 10572 3849 10628
rect 3849 10572 3853 10628
rect 3789 10568 3853 10572
rect 6146 10628 6210 10632
rect 6146 10572 6150 10628
rect 6150 10572 6206 10628
rect 6206 10572 6210 10628
rect 6146 10568 6210 10572
rect 6226 10628 6290 10632
rect 6226 10572 6230 10628
rect 6230 10572 6286 10628
rect 6286 10572 6290 10628
rect 6226 10568 6290 10572
rect 6306 10628 6370 10632
rect 6306 10572 6310 10628
rect 6310 10572 6366 10628
rect 6366 10572 6370 10628
rect 6306 10568 6370 10572
rect 6386 10628 6450 10632
rect 6386 10572 6390 10628
rect 6390 10572 6446 10628
rect 6446 10572 6450 10628
rect 6386 10568 6450 10572
rect 2250 10084 2314 10088
rect 2250 10028 2254 10084
rect 2254 10028 2310 10084
rect 2310 10028 2314 10084
rect 2250 10024 2314 10028
rect 2330 10084 2394 10088
rect 2330 10028 2334 10084
rect 2334 10028 2390 10084
rect 2390 10028 2394 10084
rect 2330 10024 2394 10028
rect 2410 10084 2474 10088
rect 2410 10028 2414 10084
rect 2414 10028 2470 10084
rect 2470 10028 2474 10084
rect 2410 10024 2474 10028
rect 2490 10084 2554 10088
rect 2490 10028 2494 10084
rect 2494 10028 2550 10084
rect 2550 10028 2554 10084
rect 2490 10024 2554 10028
rect 4848 10084 4912 10088
rect 4848 10028 4852 10084
rect 4852 10028 4908 10084
rect 4908 10028 4912 10084
rect 4848 10024 4912 10028
rect 4928 10084 4992 10088
rect 4928 10028 4932 10084
rect 4932 10028 4988 10084
rect 4988 10028 4992 10084
rect 4928 10024 4992 10028
rect 5008 10084 5072 10088
rect 5008 10028 5012 10084
rect 5012 10028 5068 10084
rect 5068 10028 5072 10084
rect 5008 10024 5072 10028
rect 5088 10084 5152 10088
rect 5088 10028 5092 10084
rect 5092 10028 5148 10084
rect 5148 10028 5152 10084
rect 5088 10024 5152 10028
rect 7445 10084 7509 10088
rect 7445 10028 7449 10084
rect 7449 10028 7505 10084
rect 7505 10028 7509 10084
rect 7445 10024 7509 10028
rect 7525 10084 7589 10088
rect 7525 10028 7529 10084
rect 7529 10028 7585 10084
rect 7585 10028 7589 10084
rect 7525 10024 7589 10028
rect 7605 10084 7669 10088
rect 7605 10028 7609 10084
rect 7609 10028 7665 10084
rect 7665 10028 7669 10084
rect 7605 10024 7669 10028
rect 7685 10084 7749 10088
rect 7685 10028 7689 10084
rect 7689 10028 7745 10084
rect 7745 10028 7749 10084
rect 7685 10024 7749 10028
rect 3549 9540 3613 9544
rect 3549 9484 3553 9540
rect 3553 9484 3609 9540
rect 3609 9484 3613 9540
rect 3549 9480 3613 9484
rect 3629 9540 3693 9544
rect 3629 9484 3633 9540
rect 3633 9484 3689 9540
rect 3689 9484 3693 9540
rect 3629 9480 3693 9484
rect 3709 9540 3773 9544
rect 3709 9484 3713 9540
rect 3713 9484 3769 9540
rect 3769 9484 3773 9540
rect 3709 9480 3773 9484
rect 3789 9540 3853 9544
rect 3789 9484 3793 9540
rect 3793 9484 3849 9540
rect 3849 9484 3853 9540
rect 3789 9480 3853 9484
rect 6146 9540 6210 9544
rect 6146 9484 6150 9540
rect 6150 9484 6206 9540
rect 6206 9484 6210 9540
rect 6146 9480 6210 9484
rect 6226 9540 6290 9544
rect 6226 9484 6230 9540
rect 6230 9484 6286 9540
rect 6286 9484 6290 9540
rect 6226 9480 6290 9484
rect 6306 9540 6370 9544
rect 6306 9484 6310 9540
rect 6310 9484 6366 9540
rect 6366 9484 6370 9540
rect 6306 9480 6370 9484
rect 6386 9540 6450 9544
rect 6386 9484 6390 9540
rect 6390 9484 6446 9540
rect 6446 9484 6450 9540
rect 6386 9480 6450 9484
rect 2250 8996 2314 9000
rect 2250 8940 2254 8996
rect 2254 8940 2310 8996
rect 2310 8940 2314 8996
rect 2250 8936 2314 8940
rect 2330 8996 2394 9000
rect 2330 8940 2334 8996
rect 2334 8940 2390 8996
rect 2390 8940 2394 8996
rect 2330 8936 2394 8940
rect 2410 8996 2474 9000
rect 2410 8940 2414 8996
rect 2414 8940 2470 8996
rect 2470 8940 2474 8996
rect 2410 8936 2474 8940
rect 2490 8996 2554 9000
rect 2490 8940 2494 8996
rect 2494 8940 2550 8996
rect 2550 8940 2554 8996
rect 2490 8936 2554 8940
rect 4848 8996 4912 9000
rect 4848 8940 4852 8996
rect 4852 8940 4908 8996
rect 4908 8940 4912 8996
rect 4848 8936 4912 8940
rect 4928 8996 4992 9000
rect 4928 8940 4932 8996
rect 4932 8940 4988 8996
rect 4988 8940 4992 8996
rect 4928 8936 4992 8940
rect 5008 8996 5072 9000
rect 5008 8940 5012 8996
rect 5012 8940 5068 8996
rect 5068 8940 5072 8996
rect 5008 8936 5072 8940
rect 5088 8996 5152 9000
rect 5088 8940 5092 8996
rect 5092 8940 5148 8996
rect 5148 8940 5152 8996
rect 5088 8936 5152 8940
rect 7445 8996 7509 9000
rect 7445 8940 7449 8996
rect 7449 8940 7505 8996
rect 7505 8940 7509 8996
rect 7445 8936 7509 8940
rect 7525 8996 7589 9000
rect 7525 8940 7529 8996
rect 7529 8940 7585 8996
rect 7585 8940 7589 8996
rect 7525 8936 7589 8940
rect 7605 8996 7669 9000
rect 7605 8940 7609 8996
rect 7609 8940 7665 8996
rect 7665 8940 7669 8996
rect 7605 8936 7669 8940
rect 7685 8996 7749 9000
rect 7685 8940 7689 8996
rect 7689 8940 7745 8996
rect 7745 8940 7749 8996
rect 7685 8936 7749 8940
rect 3549 8452 3613 8456
rect 3549 8396 3553 8452
rect 3553 8396 3609 8452
rect 3609 8396 3613 8452
rect 3549 8392 3613 8396
rect 3629 8452 3693 8456
rect 3629 8396 3633 8452
rect 3633 8396 3689 8452
rect 3689 8396 3693 8452
rect 3629 8392 3693 8396
rect 3709 8452 3773 8456
rect 3709 8396 3713 8452
rect 3713 8396 3769 8452
rect 3769 8396 3773 8452
rect 3709 8392 3773 8396
rect 3789 8452 3853 8456
rect 3789 8396 3793 8452
rect 3793 8396 3849 8452
rect 3849 8396 3853 8452
rect 3789 8392 3853 8396
rect 6146 8452 6210 8456
rect 6146 8396 6150 8452
rect 6150 8396 6206 8452
rect 6206 8396 6210 8452
rect 6146 8392 6210 8396
rect 6226 8452 6290 8456
rect 6226 8396 6230 8452
rect 6230 8396 6286 8452
rect 6286 8396 6290 8452
rect 6226 8392 6290 8396
rect 6306 8452 6370 8456
rect 6306 8396 6310 8452
rect 6310 8396 6366 8452
rect 6366 8396 6370 8452
rect 6306 8392 6370 8396
rect 6386 8452 6450 8456
rect 6386 8396 6390 8452
rect 6390 8396 6446 8452
rect 6446 8396 6450 8452
rect 6386 8392 6450 8396
rect 2250 7908 2314 7912
rect 2250 7852 2254 7908
rect 2254 7852 2310 7908
rect 2310 7852 2314 7908
rect 2250 7848 2314 7852
rect 2330 7908 2394 7912
rect 2330 7852 2334 7908
rect 2334 7852 2390 7908
rect 2390 7852 2394 7908
rect 2330 7848 2394 7852
rect 2410 7908 2474 7912
rect 2410 7852 2414 7908
rect 2414 7852 2470 7908
rect 2470 7852 2474 7908
rect 2410 7848 2474 7852
rect 2490 7908 2554 7912
rect 2490 7852 2494 7908
rect 2494 7852 2550 7908
rect 2550 7852 2554 7908
rect 2490 7848 2554 7852
rect 4848 7908 4912 7912
rect 4848 7852 4852 7908
rect 4852 7852 4908 7908
rect 4908 7852 4912 7908
rect 4848 7848 4912 7852
rect 4928 7908 4992 7912
rect 4928 7852 4932 7908
rect 4932 7852 4988 7908
rect 4988 7852 4992 7908
rect 4928 7848 4992 7852
rect 5008 7908 5072 7912
rect 5008 7852 5012 7908
rect 5012 7852 5068 7908
rect 5068 7852 5072 7908
rect 5008 7848 5072 7852
rect 5088 7908 5152 7912
rect 5088 7852 5092 7908
rect 5092 7852 5148 7908
rect 5148 7852 5152 7908
rect 5088 7848 5152 7852
rect 7445 7908 7509 7912
rect 7445 7852 7449 7908
rect 7449 7852 7505 7908
rect 7505 7852 7509 7908
rect 7445 7848 7509 7852
rect 7525 7908 7589 7912
rect 7525 7852 7529 7908
rect 7529 7852 7585 7908
rect 7585 7852 7589 7908
rect 7525 7848 7589 7852
rect 7605 7908 7669 7912
rect 7605 7852 7609 7908
rect 7609 7852 7665 7908
rect 7665 7852 7669 7908
rect 7605 7848 7669 7852
rect 7685 7908 7749 7912
rect 7685 7852 7689 7908
rect 7689 7852 7745 7908
rect 7745 7852 7749 7908
rect 7685 7848 7749 7852
rect 3549 7364 3613 7368
rect 3549 7308 3553 7364
rect 3553 7308 3609 7364
rect 3609 7308 3613 7364
rect 3549 7304 3613 7308
rect 3629 7364 3693 7368
rect 3629 7308 3633 7364
rect 3633 7308 3689 7364
rect 3689 7308 3693 7364
rect 3629 7304 3693 7308
rect 3709 7364 3773 7368
rect 3709 7308 3713 7364
rect 3713 7308 3769 7364
rect 3769 7308 3773 7364
rect 3709 7304 3773 7308
rect 3789 7364 3853 7368
rect 3789 7308 3793 7364
rect 3793 7308 3849 7364
rect 3849 7308 3853 7364
rect 3789 7304 3853 7308
rect 6146 7364 6210 7368
rect 6146 7308 6150 7364
rect 6150 7308 6206 7364
rect 6206 7308 6210 7364
rect 6146 7304 6210 7308
rect 6226 7364 6290 7368
rect 6226 7308 6230 7364
rect 6230 7308 6286 7364
rect 6286 7308 6290 7364
rect 6226 7304 6290 7308
rect 6306 7364 6370 7368
rect 6306 7308 6310 7364
rect 6310 7308 6366 7364
rect 6366 7308 6370 7364
rect 6306 7304 6370 7308
rect 6386 7364 6450 7368
rect 6386 7308 6390 7364
rect 6390 7308 6446 7364
rect 6446 7308 6450 7364
rect 6386 7304 6450 7308
rect 2250 6820 2314 6824
rect 2250 6764 2254 6820
rect 2254 6764 2310 6820
rect 2310 6764 2314 6820
rect 2250 6760 2314 6764
rect 2330 6820 2394 6824
rect 2330 6764 2334 6820
rect 2334 6764 2390 6820
rect 2390 6764 2394 6820
rect 2330 6760 2394 6764
rect 2410 6820 2474 6824
rect 2410 6764 2414 6820
rect 2414 6764 2470 6820
rect 2470 6764 2474 6820
rect 2410 6760 2474 6764
rect 2490 6820 2554 6824
rect 2490 6764 2494 6820
rect 2494 6764 2550 6820
rect 2550 6764 2554 6820
rect 2490 6760 2554 6764
rect 4848 6820 4912 6824
rect 4848 6764 4852 6820
rect 4852 6764 4908 6820
rect 4908 6764 4912 6820
rect 4848 6760 4912 6764
rect 4928 6820 4992 6824
rect 4928 6764 4932 6820
rect 4932 6764 4988 6820
rect 4988 6764 4992 6820
rect 4928 6760 4992 6764
rect 5008 6820 5072 6824
rect 5008 6764 5012 6820
rect 5012 6764 5068 6820
rect 5068 6764 5072 6820
rect 5008 6760 5072 6764
rect 5088 6820 5152 6824
rect 5088 6764 5092 6820
rect 5092 6764 5148 6820
rect 5148 6764 5152 6820
rect 5088 6760 5152 6764
rect 7445 6820 7509 6824
rect 7445 6764 7449 6820
rect 7449 6764 7505 6820
rect 7505 6764 7509 6820
rect 7445 6760 7509 6764
rect 7525 6820 7589 6824
rect 7525 6764 7529 6820
rect 7529 6764 7585 6820
rect 7585 6764 7589 6820
rect 7525 6760 7589 6764
rect 7605 6820 7669 6824
rect 7605 6764 7609 6820
rect 7609 6764 7665 6820
rect 7665 6764 7669 6820
rect 7605 6760 7669 6764
rect 7685 6820 7749 6824
rect 7685 6764 7689 6820
rect 7689 6764 7745 6820
rect 7745 6764 7749 6820
rect 7685 6760 7749 6764
rect 3549 6276 3613 6280
rect 3549 6220 3553 6276
rect 3553 6220 3609 6276
rect 3609 6220 3613 6276
rect 3549 6216 3613 6220
rect 3629 6276 3693 6280
rect 3629 6220 3633 6276
rect 3633 6220 3689 6276
rect 3689 6220 3693 6276
rect 3629 6216 3693 6220
rect 3709 6276 3773 6280
rect 3709 6220 3713 6276
rect 3713 6220 3769 6276
rect 3769 6220 3773 6276
rect 3709 6216 3773 6220
rect 3789 6276 3853 6280
rect 3789 6220 3793 6276
rect 3793 6220 3849 6276
rect 3849 6220 3853 6276
rect 3789 6216 3853 6220
rect 6146 6276 6210 6280
rect 6146 6220 6150 6276
rect 6150 6220 6206 6276
rect 6206 6220 6210 6276
rect 6146 6216 6210 6220
rect 6226 6276 6290 6280
rect 6226 6220 6230 6276
rect 6230 6220 6286 6276
rect 6286 6220 6290 6276
rect 6226 6216 6290 6220
rect 6306 6276 6370 6280
rect 6306 6220 6310 6276
rect 6310 6220 6366 6276
rect 6366 6220 6370 6276
rect 6306 6216 6370 6220
rect 6386 6276 6450 6280
rect 6386 6220 6390 6276
rect 6390 6220 6446 6276
rect 6446 6220 6450 6276
rect 6386 6216 6450 6220
rect 2250 5732 2314 5736
rect 2250 5676 2254 5732
rect 2254 5676 2310 5732
rect 2310 5676 2314 5732
rect 2250 5672 2314 5676
rect 2330 5732 2394 5736
rect 2330 5676 2334 5732
rect 2334 5676 2390 5732
rect 2390 5676 2394 5732
rect 2330 5672 2394 5676
rect 2410 5732 2474 5736
rect 2410 5676 2414 5732
rect 2414 5676 2470 5732
rect 2470 5676 2474 5732
rect 2410 5672 2474 5676
rect 2490 5732 2554 5736
rect 2490 5676 2494 5732
rect 2494 5676 2550 5732
rect 2550 5676 2554 5732
rect 2490 5672 2554 5676
rect 4848 5732 4912 5736
rect 4848 5676 4852 5732
rect 4852 5676 4908 5732
rect 4908 5676 4912 5732
rect 4848 5672 4912 5676
rect 4928 5732 4992 5736
rect 4928 5676 4932 5732
rect 4932 5676 4988 5732
rect 4988 5676 4992 5732
rect 4928 5672 4992 5676
rect 5008 5732 5072 5736
rect 5008 5676 5012 5732
rect 5012 5676 5068 5732
rect 5068 5676 5072 5732
rect 5008 5672 5072 5676
rect 5088 5732 5152 5736
rect 5088 5676 5092 5732
rect 5092 5676 5148 5732
rect 5148 5676 5152 5732
rect 5088 5672 5152 5676
rect 7445 5732 7509 5736
rect 7445 5676 7449 5732
rect 7449 5676 7505 5732
rect 7505 5676 7509 5732
rect 7445 5672 7509 5676
rect 7525 5732 7589 5736
rect 7525 5676 7529 5732
rect 7529 5676 7585 5732
rect 7585 5676 7589 5732
rect 7525 5672 7589 5676
rect 7605 5732 7669 5736
rect 7605 5676 7609 5732
rect 7609 5676 7665 5732
rect 7665 5676 7669 5732
rect 7605 5672 7669 5676
rect 7685 5732 7749 5736
rect 7685 5676 7689 5732
rect 7689 5676 7745 5732
rect 7745 5676 7749 5732
rect 7685 5672 7749 5676
rect 3549 5188 3613 5192
rect 3549 5132 3553 5188
rect 3553 5132 3609 5188
rect 3609 5132 3613 5188
rect 3549 5128 3613 5132
rect 3629 5188 3693 5192
rect 3629 5132 3633 5188
rect 3633 5132 3689 5188
rect 3689 5132 3693 5188
rect 3629 5128 3693 5132
rect 3709 5188 3773 5192
rect 3709 5132 3713 5188
rect 3713 5132 3769 5188
rect 3769 5132 3773 5188
rect 3709 5128 3773 5132
rect 3789 5188 3853 5192
rect 3789 5132 3793 5188
rect 3793 5132 3849 5188
rect 3849 5132 3853 5188
rect 3789 5128 3853 5132
rect 6146 5188 6210 5192
rect 6146 5132 6150 5188
rect 6150 5132 6206 5188
rect 6206 5132 6210 5188
rect 6146 5128 6210 5132
rect 6226 5188 6290 5192
rect 6226 5132 6230 5188
rect 6230 5132 6286 5188
rect 6286 5132 6290 5188
rect 6226 5128 6290 5132
rect 6306 5188 6370 5192
rect 6306 5132 6310 5188
rect 6310 5132 6366 5188
rect 6366 5132 6370 5188
rect 6306 5128 6370 5132
rect 6386 5188 6450 5192
rect 6386 5132 6390 5188
rect 6390 5132 6446 5188
rect 6446 5132 6450 5188
rect 6386 5128 6450 5132
rect 2250 4644 2314 4648
rect 2250 4588 2254 4644
rect 2254 4588 2310 4644
rect 2310 4588 2314 4644
rect 2250 4584 2314 4588
rect 2330 4644 2394 4648
rect 2330 4588 2334 4644
rect 2334 4588 2390 4644
rect 2390 4588 2394 4644
rect 2330 4584 2394 4588
rect 2410 4644 2474 4648
rect 2410 4588 2414 4644
rect 2414 4588 2470 4644
rect 2470 4588 2474 4644
rect 2410 4584 2474 4588
rect 2490 4644 2554 4648
rect 2490 4588 2494 4644
rect 2494 4588 2550 4644
rect 2550 4588 2554 4644
rect 2490 4584 2554 4588
rect 4848 4644 4912 4648
rect 4848 4588 4852 4644
rect 4852 4588 4908 4644
rect 4908 4588 4912 4644
rect 4848 4584 4912 4588
rect 4928 4644 4992 4648
rect 4928 4588 4932 4644
rect 4932 4588 4988 4644
rect 4988 4588 4992 4644
rect 4928 4584 4992 4588
rect 5008 4644 5072 4648
rect 5008 4588 5012 4644
rect 5012 4588 5068 4644
rect 5068 4588 5072 4644
rect 5008 4584 5072 4588
rect 5088 4644 5152 4648
rect 5088 4588 5092 4644
rect 5092 4588 5148 4644
rect 5148 4588 5152 4644
rect 5088 4584 5152 4588
rect 7445 4644 7509 4648
rect 7445 4588 7449 4644
rect 7449 4588 7505 4644
rect 7505 4588 7509 4644
rect 7445 4584 7509 4588
rect 7525 4644 7589 4648
rect 7525 4588 7529 4644
rect 7529 4588 7585 4644
rect 7585 4588 7589 4644
rect 7525 4584 7589 4588
rect 7605 4644 7669 4648
rect 7605 4588 7609 4644
rect 7609 4588 7665 4644
rect 7665 4588 7669 4644
rect 7605 4584 7669 4588
rect 7685 4644 7749 4648
rect 7685 4588 7689 4644
rect 7689 4588 7745 4644
rect 7745 4588 7749 4644
rect 7685 4584 7749 4588
rect 3549 4100 3613 4104
rect 3549 4044 3553 4100
rect 3553 4044 3609 4100
rect 3609 4044 3613 4100
rect 3549 4040 3613 4044
rect 3629 4100 3693 4104
rect 3629 4044 3633 4100
rect 3633 4044 3689 4100
rect 3689 4044 3693 4100
rect 3629 4040 3693 4044
rect 3709 4100 3773 4104
rect 3709 4044 3713 4100
rect 3713 4044 3769 4100
rect 3769 4044 3773 4100
rect 3709 4040 3773 4044
rect 3789 4100 3853 4104
rect 3789 4044 3793 4100
rect 3793 4044 3849 4100
rect 3849 4044 3853 4100
rect 3789 4040 3853 4044
rect 6146 4100 6210 4104
rect 6146 4044 6150 4100
rect 6150 4044 6206 4100
rect 6206 4044 6210 4100
rect 6146 4040 6210 4044
rect 6226 4100 6290 4104
rect 6226 4044 6230 4100
rect 6230 4044 6286 4100
rect 6286 4044 6290 4100
rect 6226 4040 6290 4044
rect 6306 4100 6370 4104
rect 6306 4044 6310 4100
rect 6310 4044 6366 4100
rect 6366 4044 6370 4100
rect 6306 4040 6370 4044
rect 6386 4100 6450 4104
rect 6386 4044 6390 4100
rect 6390 4044 6446 4100
rect 6446 4044 6450 4100
rect 6386 4040 6450 4044
rect 2250 3556 2314 3560
rect 2250 3500 2254 3556
rect 2254 3500 2310 3556
rect 2310 3500 2314 3556
rect 2250 3496 2314 3500
rect 2330 3556 2394 3560
rect 2330 3500 2334 3556
rect 2334 3500 2390 3556
rect 2390 3500 2394 3556
rect 2330 3496 2394 3500
rect 2410 3556 2474 3560
rect 2410 3500 2414 3556
rect 2414 3500 2470 3556
rect 2470 3500 2474 3556
rect 2410 3496 2474 3500
rect 2490 3556 2554 3560
rect 2490 3500 2494 3556
rect 2494 3500 2550 3556
rect 2550 3500 2554 3556
rect 2490 3496 2554 3500
rect 4848 3556 4912 3560
rect 4848 3500 4852 3556
rect 4852 3500 4908 3556
rect 4908 3500 4912 3556
rect 4848 3496 4912 3500
rect 4928 3556 4992 3560
rect 4928 3500 4932 3556
rect 4932 3500 4988 3556
rect 4988 3500 4992 3556
rect 4928 3496 4992 3500
rect 5008 3556 5072 3560
rect 5008 3500 5012 3556
rect 5012 3500 5068 3556
rect 5068 3500 5072 3556
rect 5008 3496 5072 3500
rect 5088 3556 5152 3560
rect 5088 3500 5092 3556
rect 5092 3500 5148 3556
rect 5148 3500 5152 3556
rect 5088 3496 5152 3500
rect 7445 3556 7509 3560
rect 7445 3500 7449 3556
rect 7449 3500 7505 3556
rect 7505 3500 7509 3556
rect 7445 3496 7509 3500
rect 7525 3556 7589 3560
rect 7525 3500 7529 3556
rect 7529 3500 7585 3556
rect 7585 3500 7589 3556
rect 7525 3496 7589 3500
rect 7605 3556 7669 3560
rect 7605 3500 7609 3556
rect 7609 3500 7665 3556
rect 7665 3500 7669 3556
rect 7605 3496 7669 3500
rect 7685 3556 7749 3560
rect 7685 3500 7689 3556
rect 7689 3500 7745 3556
rect 7745 3500 7749 3556
rect 7685 3496 7749 3500
rect 3549 3012 3613 3016
rect 3549 2956 3553 3012
rect 3553 2956 3609 3012
rect 3609 2956 3613 3012
rect 3549 2952 3613 2956
rect 3629 3012 3693 3016
rect 3629 2956 3633 3012
rect 3633 2956 3689 3012
rect 3689 2956 3693 3012
rect 3629 2952 3693 2956
rect 3709 3012 3773 3016
rect 3709 2956 3713 3012
rect 3713 2956 3769 3012
rect 3769 2956 3773 3012
rect 3709 2952 3773 2956
rect 3789 3012 3853 3016
rect 3789 2956 3793 3012
rect 3793 2956 3849 3012
rect 3849 2956 3853 3012
rect 3789 2952 3853 2956
rect 6146 3012 6210 3016
rect 6146 2956 6150 3012
rect 6150 2956 6206 3012
rect 6206 2956 6210 3012
rect 6146 2952 6210 2956
rect 6226 3012 6290 3016
rect 6226 2956 6230 3012
rect 6230 2956 6286 3012
rect 6286 2956 6290 3012
rect 6226 2952 6290 2956
rect 6306 3012 6370 3016
rect 6306 2956 6310 3012
rect 6310 2956 6366 3012
rect 6366 2956 6370 3012
rect 6306 2952 6370 2956
rect 6386 3012 6450 3016
rect 6386 2956 6390 3012
rect 6390 2956 6446 3012
rect 6446 2956 6450 3012
rect 6386 2952 6450 2956
rect 2250 2468 2314 2472
rect 2250 2412 2254 2468
rect 2254 2412 2310 2468
rect 2310 2412 2314 2468
rect 2250 2408 2314 2412
rect 2330 2468 2394 2472
rect 2330 2412 2334 2468
rect 2334 2412 2390 2468
rect 2390 2412 2394 2468
rect 2330 2408 2394 2412
rect 2410 2468 2474 2472
rect 2410 2412 2414 2468
rect 2414 2412 2470 2468
rect 2470 2412 2474 2468
rect 2410 2408 2474 2412
rect 2490 2468 2554 2472
rect 2490 2412 2494 2468
rect 2494 2412 2550 2468
rect 2550 2412 2554 2468
rect 2490 2408 2554 2412
rect 4848 2468 4912 2472
rect 4848 2412 4852 2468
rect 4852 2412 4908 2468
rect 4908 2412 4912 2468
rect 4848 2408 4912 2412
rect 4928 2468 4992 2472
rect 4928 2412 4932 2468
rect 4932 2412 4988 2468
rect 4988 2412 4992 2468
rect 4928 2408 4992 2412
rect 5008 2468 5072 2472
rect 5008 2412 5012 2468
rect 5012 2412 5068 2468
rect 5068 2412 5072 2468
rect 5008 2408 5072 2412
rect 5088 2468 5152 2472
rect 5088 2412 5092 2468
rect 5092 2412 5148 2468
rect 5148 2412 5152 2468
rect 5088 2408 5152 2412
rect 7445 2468 7509 2472
rect 7445 2412 7449 2468
rect 7449 2412 7505 2468
rect 7505 2412 7509 2468
rect 7445 2408 7509 2412
rect 7525 2468 7589 2472
rect 7525 2412 7529 2468
rect 7529 2412 7585 2468
rect 7585 2412 7589 2468
rect 7525 2408 7589 2412
rect 7605 2468 7669 2472
rect 7605 2412 7609 2468
rect 7609 2412 7665 2468
rect 7665 2412 7669 2468
rect 7605 2408 7669 2412
rect 7685 2468 7749 2472
rect 7685 2412 7689 2468
rect 7689 2412 7745 2468
rect 7745 2412 7749 2468
rect 7685 2408 7749 2412
rect 3549 1924 3613 1928
rect 3549 1868 3553 1924
rect 3553 1868 3609 1924
rect 3609 1868 3613 1924
rect 3549 1864 3613 1868
rect 3629 1924 3693 1928
rect 3629 1868 3633 1924
rect 3633 1868 3689 1924
rect 3689 1868 3693 1924
rect 3629 1864 3693 1868
rect 3709 1924 3773 1928
rect 3709 1868 3713 1924
rect 3713 1868 3769 1924
rect 3769 1868 3773 1924
rect 3709 1864 3773 1868
rect 3789 1924 3853 1928
rect 3789 1868 3793 1924
rect 3793 1868 3849 1924
rect 3849 1868 3853 1924
rect 3789 1864 3853 1868
rect 6146 1924 6210 1928
rect 6146 1868 6150 1924
rect 6150 1868 6206 1924
rect 6206 1868 6210 1924
rect 6146 1864 6210 1868
rect 6226 1924 6290 1928
rect 6226 1868 6230 1924
rect 6230 1868 6286 1924
rect 6286 1868 6290 1924
rect 6226 1864 6290 1868
rect 6306 1924 6370 1928
rect 6306 1868 6310 1924
rect 6310 1868 6366 1924
rect 6366 1868 6370 1924
rect 6306 1864 6370 1868
rect 6386 1924 6450 1928
rect 6386 1868 6390 1924
rect 6390 1868 6446 1924
rect 6446 1868 6450 1924
rect 6386 1864 6450 1868
rect 2250 1380 2314 1384
rect 2250 1324 2254 1380
rect 2254 1324 2310 1380
rect 2310 1324 2314 1380
rect 2250 1320 2314 1324
rect 2330 1380 2394 1384
rect 2330 1324 2334 1380
rect 2334 1324 2390 1380
rect 2390 1324 2394 1380
rect 2330 1320 2394 1324
rect 2410 1380 2474 1384
rect 2410 1324 2414 1380
rect 2414 1324 2470 1380
rect 2470 1324 2474 1380
rect 2410 1320 2474 1324
rect 2490 1380 2554 1384
rect 2490 1324 2494 1380
rect 2494 1324 2550 1380
rect 2550 1324 2554 1380
rect 2490 1320 2554 1324
rect 4848 1380 4912 1384
rect 4848 1324 4852 1380
rect 4852 1324 4908 1380
rect 4908 1324 4912 1380
rect 4848 1320 4912 1324
rect 4928 1380 4992 1384
rect 4928 1324 4932 1380
rect 4932 1324 4988 1380
rect 4988 1324 4992 1380
rect 4928 1320 4992 1324
rect 5008 1380 5072 1384
rect 5008 1324 5012 1380
rect 5012 1324 5068 1380
rect 5068 1324 5072 1380
rect 5008 1320 5072 1324
rect 5088 1380 5152 1384
rect 5088 1324 5092 1380
rect 5092 1324 5148 1380
rect 5148 1324 5152 1380
rect 5088 1320 5152 1324
rect 7445 1380 7509 1384
rect 7445 1324 7449 1380
rect 7449 1324 7505 1380
rect 7505 1324 7509 1380
rect 7445 1320 7509 1324
rect 7525 1380 7589 1384
rect 7525 1324 7529 1380
rect 7529 1324 7585 1380
rect 7585 1324 7589 1380
rect 7525 1320 7589 1324
rect 7605 1380 7669 1384
rect 7605 1324 7609 1380
rect 7609 1324 7665 1380
rect 7665 1324 7669 1380
rect 7605 1320 7669 1324
rect 7685 1380 7749 1384
rect 7685 1324 7689 1380
rect 7689 1324 7745 1380
rect 7745 1324 7749 1380
rect 7685 1320 7749 1324
<< metal4 >>
rect 2242 20968 2562 21528
rect 2242 20904 2250 20968
rect 2314 20904 2330 20968
rect 2394 20904 2410 20968
rect 2474 20904 2490 20968
rect 2554 20904 2562 20968
rect 2242 19880 2562 20904
rect 2242 19816 2250 19880
rect 2314 19816 2330 19880
rect 2394 19816 2410 19880
rect 2474 19816 2490 19880
rect 2554 19816 2562 19880
rect 2242 18792 2562 19816
rect 2242 18728 2250 18792
rect 2314 18728 2330 18792
rect 2394 18728 2410 18792
rect 2474 18728 2490 18792
rect 2554 18728 2562 18792
rect 2242 18628 2562 18728
rect 2242 18392 2284 18628
rect 2520 18392 2562 18628
rect 2242 17704 2562 18392
rect 2242 17640 2250 17704
rect 2314 17640 2330 17704
rect 2394 17640 2410 17704
rect 2474 17640 2490 17704
rect 2554 17640 2562 17704
rect 2242 16616 2562 17640
rect 2242 16552 2250 16616
rect 2314 16552 2330 16616
rect 2394 16552 2410 16616
rect 2474 16552 2490 16616
rect 2554 16552 2562 16616
rect 2242 15528 2562 16552
rect 2242 15464 2250 15528
rect 2314 15464 2330 15528
rect 2394 15464 2410 15528
rect 2474 15464 2490 15528
rect 2554 15464 2562 15528
rect 2242 14440 2562 15464
rect 2242 14376 2250 14440
rect 2314 14376 2330 14440
rect 2394 14376 2410 14440
rect 2474 14376 2490 14440
rect 2554 14376 2562 14440
rect 2242 13352 2562 14376
rect 2242 13288 2250 13352
rect 2314 13288 2330 13352
rect 2394 13288 2410 13352
rect 2474 13288 2490 13352
rect 2554 13288 2562 13352
rect 2242 12264 2562 13288
rect 2242 12200 2250 12264
rect 2314 12200 2330 12264
rect 2394 12200 2410 12264
rect 2474 12200 2490 12264
rect 2554 12200 2562 12264
rect 2242 11746 2562 12200
rect 2242 11510 2284 11746
rect 2520 11510 2562 11746
rect 2242 11176 2562 11510
rect 2242 11112 2250 11176
rect 2314 11112 2330 11176
rect 2394 11112 2410 11176
rect 2474 11112 2490 11176
rect 2554 11112 2562 11176
rect 2242 10088 2562 11112
rect 2242 10024 2250 10088
rect 2314 10024 2330 10088
rect 2394 10024 2410 10088
rect 2474 10024 2490 10088
rect 2554 10024 2562 10088
rect 2242 9000 2562 10024
rect 2242 8936 2250 9000
rect 2314 8936 2330 9000
rect 2394 8936 2410 9000
rect 2474 8936 2490 9000
rect 2554 8936 2562 9000
rect 2242 7912 2562 8936
rect 2242 7848 2250 7912
rect 2314 7848 2330 7912
rect 2394 7848 2410 7912
rect 2474 7848 2490 7912
rect 2554 7848 2562 7912
rect 2242 6824 2562 7848
rect 2242 6760 2250 6824
rect 2314 6760 2330 6824
rect 2394 6760 2410 6824
rect 2474 6760 2490 6824
rect 2554 6760 2562 6824
rect 2242 5736 2562 6760
rect 2242 5672 2250 5736
rect 2314 5672 2330 5736
rect 2394 5672 2410 5736
rect 2474 5672 2490 5736
rect 2554 5672 2562 5736
rect 2242 4863 2562 5672
rect 2242 4648 2284 4863
rect 2520 4648 2562 4863
rect 2242 4584 2250 4648
rect 2314 4584 2330 4627
rect 2394 4584 2410 4627
rect 2474 4584 2490 4627
rect 2554 4584 2562 4648
rect 2242 3560 2562 4584
rect 2242 3496 2250 3560
rect 2314 3496 2330 3560
rect 2394 3496 2410 3560
rect 2474 3496 2490 3560
rect 2554 3496 2562 3560
rect 2242 2472 2562 3496
rect 2242 2408 2250 2472
rect 2314 2408 2330 2472
rect 2394 2408 2410 2472
rect 2474 2408 2490 2472
rect 2554 2408 2562 2472
rect 2242 1384 2562 2408
rect 2242 1320 2250 1384
rect 2314 1320 2330 1384
rect 2394 1320 2410 1384
rect 2474 1320 2490 1384
rect 2554 1320 2562 1384
rect 2242 1304 2562 1320
rect 3541 21512 3861 21528
rect 3541 21448 3549 21512
rect 3613 21448 3629 21512
rect 3693 21448 3709 21512
rect 3773 21448 3789 21512
rect 3853 21448 3861 21512
rect 3541 20424 3861 21448
rect 3541 20360 3549 20424
rect 3613 20360 3629 20424
rect 3693 20360 3709 20424
rect 3773 20360 3789 20424
rect 3853 20360 3861 20424
rect 3541 19336 3861 20360
rect 3541 19272 3549 19336
rect 3613 19272 3629 19336
rect 3693 19272 3709 19336
rect 3773 19272 3789 19336
rect 3853 19272 3861 19336
rect 3541 18248 3861 19272
rect 3541 18184 3549 18248
rect 3613 18184 3629 18248
rect 3693 18184 3709 18248
rect 3773 18184 3789 18248
rect 3853 18184 3861 18248
rect 3541 17160 3861 18184
rect 3541 17096 3549 17160
rect 3613 17096 3629 17160
rect 3693 17096 3709 17160
rect 3773 17096 3789 17160
rect 3853 17096 3861 17160
rect 3541 16072 3861 17096
rect 3541 16008 3549 16072
rect 3613 16008 3629 16072
rect 3693 16008 3709 16072
rect 3773 16008 3789 16072
rect 3853 16008 3861 16072
rect 3541 15187 3861 16008
rect 3541 14984 3583 15187
rect 3819 14984 3861 15187
rect 3541 14920 3549 14984
rect 3613 14920 3629 14951
rect 3693 14920 3709 14951
rect 3773 14920 3789 14951
rect 3853 14920 3861 14984
rect 3541 13896 3861 14920
rect 3541 13832 3549 13896
rect 3613 13832 3629 13896
rect 3693 13832 3709 13896
rect 3773 13832 3789 13896
rect 3853 13832 3861 13896
rect 3541 12808 3861 13832
rect 3541 12744 3549 12808
rect 3613 12744 3629 12808
rect 3693 12744 3709 12808
rect 3773 12744 3789 12808
rect 3853 12744 3861 12808
rect 3541 11720 3861 12744
rect 3541 11656 3549 11720
rect 3613 11656 3629 11720
rect 3693 11656 3709 11720
rect 3773 11656 3789 11720
rect 3853 11656 3861 11720
rect 3541 10632 3861 11656
rect 3541 10568 3549 10632
rect 3613 10568 3629 10632
rect 3693 10568 3709 10632
rect 3773 10568 3789 10632
rect 3853 10568 3861 10632
rect 3541 9544 3861 10568
rect 3541 9480 3549 9544
rect 3613 9480 3629 9544
rect 3693 9480 3709 9544
rect 3773 9480 3789 9544
rect 3853 9480 3861 9544
rect 3541 8456 3861 9480
rect 3541 8392 3549 8456
rect 3613 8392 3629 8456
rect 3693 8392 3709 8456
rect 3773 8392 3789 8456
rect 3853 8392 3861 8456
rect 3541 8304 3861 8392
rect 3541 8068 3583 8304
rect 3819 8068 3861 8304
rect 3541 7368 3861 8068
rect 3541 7304 3549 7368
rect 3613 7304 3629 7368
rect 3693 7304 3709 7368
rect 3773 7304 3789 7368
rect 3853 7304 3861 7368
rect 3541 6280 3861 7304
rect 3541 6216 3549 6280
rect 3613 6216 3629 6280
rect 3693 6216 3709 6280
rect 3773 6216 3789 6280
rect 3853 6216 3861 6280
rect 3541 5192 3861 6216
rect 3541 5128 3549 5192
rect 3613 5128 3629 5192
rect 3693 5128 3709 5192
rect 3773 5128 3789 5192
rect 3853 5128 3861 5192
rect 3541 4104 3861 5128
rect 3541 4040 3549 4104
rect 3613 4040 3629 4104
rect 3693 4040 3709 4104
rect 3773 4040 3789 4104
rect 3853 4040 3861 4104
rect 3541 3016 3861 4040
rect 3541 2952 3549 3016
rect 3613 2952 3629 3016
rect 3693 2952 3709 3016
rect 3773 2952 3789 3016
rect 3853 2952 3861 3016
rect 3541 1928 3861 2952
rect 3541 1864 3549 1928
rect 3613 1864 3629 1928
rect 3693 1864 3709 1928
rect 3773 1864 3789 1928
rect 3853 1864 3861 1928
rect 3541 1304 3861 1864
rect 4840 20968 5160 21528
rect 4840 20904 4848 20968
rect 4912 20904 4928 20968
rect 4992 20904 5008 20968
rect 5072 20904 5088 20968
rect 5152 20904 5160 20968
rect 4840 19880 5160 20904
rect 4840 19816 4848 19880
rect 4912 19816 4928 19880
rect 4992 19816 5008 19880
rect 5072 19816 5088 19880
rect 5152 19816 5160 19880
rect 4840 18792 5160 19816
rect 4840 18728 4848 18792
rect 4912 18728 4928 18792
rect 4992 18728 5008 18792
rect 5072 18728 5088 18792
rect 5152 18728 5160 18792
rect 4840 18628 5160 18728
rect 4840 18392 4882 18628
rect 5118 18392 5160 18628
rect 4840 17704 5160 18392
rect 4840 17640 4848 17704
rect 4912 17640 4928 17704
rect 4992 17640 5008 17704
rect 5072 17640 5088 17704
rect 5152 17640 5160 17704
rect 4840 16616 5160 17640
rect 4840 16552 4848 16616
rect 4912 16552 4928 16616
rect 4992 16552 5008 16616
rect 5072 16552 5088 16616
rect 5152 16552 5160 16616
rect 4840 15528 5160 16552
rect 4840 15464 4848 15528
rect 4912 15464 4928 15528
rect 4992 15464 5008 15528
rect 5072 15464 5088 15528
rect 5152 15464 5160 15528
rect 4840 14440 5160 15464
rect 4840 14376 4848 14440
rect 4912 14376 4928 14440
rect 4992 14376 5008 14440
rect 5072 14376 5088 14440
rect 5152 14376 5160 14440
rect 4840 13352 5160 14376
rect 4840 13288 4848 13352
rect 4912 13288 4928 13352
rect 4992 13288 5008 13352
rect 5072 13288 5088 13352
rect 5152 13288 5160 13352
rect 4840 12264 5160 13288
rect 4840 12200 4848 12264
rect 4912 12200 4928 12264
rect 4992 12200 5008 12264
rect 5072 12200 5088 12264
rect 5152 12200 5160 12264
rect 4840 11746 5160 12200
rect 4840 11510 4882 11746
rect 5118 11510 5160 11746
rect 4840 11176 5160 11510
rect 4840 11112 4848 11176
rect 4912 11112 4928 11176
rect 4992 11112 5008 11176
rect 5072 11112 5088 11176
rect 5152 11112 5160 11176
rect 4840 10088 5160 11112
rect 4840 10024 4848 10088
rect 4912 10024 4928 10088
rect 4992 10024 5008 10088
rect 5072 10024 5088 10088
rect 5152 10024 5160 10088
rect 4840 9000 5160 10024
rect 4840 8936 4848 9000
rect 4912 8936 4928 9000
rect 4992 8936 5008 9000
rect 5072 8936 5088 9000
rect 5152 8936 5160 9000
rect 4840 7912 5160 8936
rect 4840 7848 4848 7912
rect 4912 7848 4928 7912
rect 4992 7848 5008 7912
rect 5072 7848 5088 7912
rect 5152 7848 5160 7912
rect 4840 6824 5160 7848
rect 4840 6760 4848 6824
rect 4912 6760 4928 6824
rect 4992 6760 5008 6824
rect 5072 6760 5088 6824
rect 5152 6760 5160 6824
rect 4840 5736 5160 6760
rect 4840 5672 4848 5736
rect 4912 5672 4928 5736
rect 4992 5672 5008 5736
rect 5072 5672 5088 5736
rect 5152 5672 5160 5736
rect 4840 4863 5160 5672
rect 4840 4648 4882 4863
rect 5118 4648 5160 4863
rect 4840 4584 4848 4648
rect 4912 4584 4928 4627
rect 4992 4584 5008 4627
rect 5072 4584 5088 4627
rect 5152 4584 5160 4648
rect 4840 3560 5160 4584
rect 4840 3496 4848 3560
rect 4912 3496 4928 3560
rect 4992 3496 5008 3560
rect 5072 3496 5088 3560
rect 5152 3496 5160 3560
rect 4840 2472 5160 3496
rect 4840 2408 4848 2472
rect 4912 2408 4928 2472
rect 4992 2408 5008 2472
rect 5072 2408 5088 2472
rect 5152 2408 5160 2472
rect 4840 1384 5160 2408
rect 4840 1320 4848 1384
rect 4912 1320 4928 1384
rect 4992 1320 5008 1384
rect 5072 1320 5088 1384
rect 5152 1320 5160 1384
rect 4840 1304 5160 1320
rect 6138 21512 6458 21528
rect 6138 21448 6146 21512
rect 6210 21448 6226 21512
rect 6290 21448 6306 21512
rect 6370 21448 6386 21512
rect 6450 21448 6458 21512
rect 6138 20424 6458 21448
rect 6138 20360 6146 20424
rect 6210 20360 6226 20424
rect 6290 20360 6306 20424
rect 6370 20360 6386 20424
rect 6450 20360 6458 20424
rect 6138 19336 6458 20360
rect 6138 19272 6146 19336
rect 6210 19272 6226 19336
rect 6290 19272 6306 19336
rect 6370 19272 6386 19336
rect 6450 19272 6458 19336
rect 6138 18248 6458 19272
rect 6138 18184 6146 18248
rect 6210 18184 6226 18248
rect 6290 18184 6306 18248
rect 6370 18184 6386 18248
rect 6450 18184 6458 18248
rect 6138 17160 6458 18184
rect 6138 17096 6146 17160
rect 6210 17096 6226 17160
rect 6290 17096 6306 17160
rect 6370 17096 6386 17160
rect 6450 17096 6458 17160
rect 6138 16072 6458 17096
rect 6138 16008 6146 16072
rect 6210 16008 6226 16072
rect 6290 16008 6306 16072
rect 6370 16008 6386 16072
rect 6450 16008 6458 16072
rect 6138 15187 6458 16008
rect 6138 14984 6180 15187
rect 6416 14984 6458 15187
rect 6138 14920 6146 14984
rect 6210 14920 6226 14951
rect 6290 14920 6306 14951
rect 6370 14920 6386 14951
rect 6450 14920 6458 14984
rect 6138 13896 6458 14920
rect 6138 13832 6146 13896
rect 6210 13832 6226 13896
rect 6290 13832 6306 13896
rect 6370 13832 6386 13896
rect 6450 13832 6458 13896
rect 6138 12808 6458 13832
rect 6138 12744 6146 12808
rect 6210 12744 6226 12808
rect 6290 12744 6306 12808
rect 6370 12744 6386 12808
rect 6450 12744 6458 12808
rect 6138 11720 6458 12744
rect 6138 11656 6146 11720
rect 6210 11656 6226 11720
rect 6290 11656 6306 11720
rect 6370 11656 6386 11720
rect 6450 11656 6458 11720
rect 6138 10632 6458 11656
rect 6138 10568 6146 10632
rect 6210 10568 6226 10632
rect 6290 10568 6306 10632
rect 6370 10568 6386 10632
rect 6450 10568 6458 10632
rect 6138 9544 6458 10568
rect 6138 9480 6146 9544
rect 6210 9480 6226 9544
rect 6290 9480 6306 9544
rect 6370 9480 6386 9544
rect 6450 9480 6458 9544
rect 6138 8456 6458 9480
rect 6138 8392 6146 8456
rect 6210 8392 6226 8456
rect 6290 8392 6306 8456
rect 6370 8392 6386 8456
rect 6450 8392 6458 8456
rect 6138 8304 6458 8392
rect 6138 8068 6180 8304
rect 6416 8068 6458 8304
rect 6138 7368 6458 8068
rect 6138 7304 6146 7368
rect 6210 7304 6226 7368
rect 6290 7304 6306 7368
rect 6370 7304 6386 7368
rect 6450 7304 6458 7368
rect 6138 6280 6458 7304
rect 6138 6216 6146 6280
rect 6210 6216 6226 6280
rect 6290 6216 6306 6280
rect 6370 6216 6386 6280
rect 6450 6216 6458 6280
rect 6138 5192 6458 6216
rect 6138 5128 6146 5192
rect 6210 5128 6226 5192
rect 6290 5128 6306 5192
rect 6370 5128 6386 5192
rect 6450 5128 6458 5192
rect 6138 4104 6458 5128
rect 6138 4040 6146 4104
rect 6210 4040 6226 4104
rect 6290 4040 6306 4104
rect 6370 4040 6386 4104
rect 6450 4040 6458 4104
rect 6138 3016 6458 4040
rect 6138 2952 6146 3016
rect 6210 2952 6226 3016
rect 6290 2952 6306 3016
rect 6370 2952 6386 3016
rect 6450 2952 6458 3016
rect 6138 1928 6458 2952
rect 6138 1864 6146 1928
rect 6210 1864 6226 1928
rect 6290 1864 6306 1928
rect 6370 1864 6386 1928
rect 6450 1864 6458 1928
rect 6138 1304 6458 1864
rect 7437 20968 7757 21528
rect 7437 20904 7445 20968
rect 7509 20904 7525 20968
rect 7589 20904 7605 20968
rect 7669 20904 7685 20968
rect 7749 20904 7757 20968
rect 7437 19880 7757 20904
rect 7437 19816 7445 19880
rect 7509 19816 7525 19880
rect 7589 19816 7605 19880
rect 7669 19816 7685 19880
rect 7749 19816 7757 19880
rect 7437 18792 7757 19816
rect 7437 18728 7445 18792
rect 7509 18728 7525 18792
rect 7589 18728 7605 18792
rect 7669 18728 7685 18792
rect 7749 18728 7757 18792
rect 7437 18628 7757 18728
rect 7437 18392 7479 18628
rect 7715 18392 7757 18628
rect 7437 17704 7757 18392
rect 7437 17640 7445 17704
rect 7509 17640 7525 17704
rect 7589 17640 7605 17704
rect 7669 17640 7685 17704
rect 7749 17640 7757 17704
rect 7437 16616 7757 17640
rect 7437 16552 7445 16616
rect 7509 16552 7525 16616
rect 7589 16552 7605 16616
rect 7669 16552 7685 16616
rect 7749 16552 7757 16616
rect 7437 15528 7757 16552
rect 7437 15464 7445 15528
rect 7509 15464 7525 15528
rect 7589 15464 7605 15528
rect 7669 15464 7685 15528
rect 7749 15464 7757 15528
rect 7437 14440 7757 15464
rect 7437 14376 7445 14440
rect 7509 14376 7525 14440
rect 7589 14376 7605 14440
rect 7669 14376 7685 14440
rect 7749 14376 7757 14440
rect 7437 13352 7757 14376
rect 7437 13288 7445 13352
rect 7509 13288 7525 13352
rect 7589 13288 7605 13352
rect 7669 13288 7685 13352
rect 7749 13288 7757 13352
rect 7437 12264 7757 13288
rect 7437 12200 7445 12264
rect 7509 12200 7525 12264
rect 7589 12200 7605 12264
rect 7669 12200 7685 12264
rect 7749 12200 7757 12264
rect 7437 11746 7757 12200
rect 7437 11510 7479 11746
rect 7715 11510 7757 11746
rect 7437 11176 7757 11510
rect 7437 11112 7445 11176
rect 7509 11112 7525 11176
rect 7589 11112 7605 11176
rect 7669 11112 7685 11176
rect 7749 11112 7757 11176
rect 7437 10088 7757 11112
rect 7437 10024 7445 10088
rect 7509 10024 7525 10088
rect 7589 10024 7605 10088
rect 7669 10024 7685 10088
rect 7749 10024 7757 10088
rect 7437 9000 7757 10024
rect 7437 8936 7445 9000
rect 7509 8936 7525 9000
rect 7589 8936 7605 9000
rect 7669 8936 7685 9000
rect 7749 8936 7757 9000
rect 7437 7912 7757 8936
rect 7437 7848 7445 7912
rect 7509 7848 7525 7912
rect 7589 7848 7605 7912
rect 7669 7848 7685 7912
rect 7749 7848 7757 7912
rect 7437 6824 7757 7848
rect 7437 6760 7445 6824
rect 7509 6760 7525 6824
rect 7589 6760 7605 6824
rect 7669 6760 7685 6824
rect 7749 6760 7757 6824
rect 7437 5736 7757 6760
rect 7437 5672 7445 5736
rect 7509 5672 7525 5736
rect 7589 5672 7605 5736
rect 7669 5672 7685 5736
rect 7749 5672 7757 5736
rect 7437 4863 7757 5672
rect 7437 4648 7479 4863
rect 7715 4648 7757 4863
rect 7437 4584 7445 4648
rect 7509 4584 7525 4627
rect 7589 4584 7605 4627
rect 7669 4584 7685 4627
rect 7749 4584 7757 4648
rect 7437 3560 7757 4584
rect 7437 3496 7445 3560
rect 7509 3496 7525 3560
rect 7589 3496 7605 3560
rect 7669 3496 7685 3560
rect 7749 3496 7757 3560
rect 7437 2472 7757 3496
rect 7437 2408 7445 2472
rect 7509 2408 7525 2472
rect 7589 2408 7605 2472
rect 7669 2408 7685 2472
rect 7749 2408 7757 2472
rect 7437 1384 7757 2408
rect 7437 1320 7445 1384
rect 7509 1320 7525 1384
rect 7589 1320 7605 1384
rect 7669 1320 7685 1384
rect 7749 1320 7757 1384
rect 7437 1304 7757 1320
<< via4 >>
rect 2284 18392 2520 18628
rect 2284 11510 2520 11746
rect 2284 4648 2520 4863
rect 2284 4627 2314 4648
rect 2314 4627 2330 4648
rect 2330 4627 2394 4648
rect 2394 4627 2410 4648
rect 2410 4627 2474 4648
rect 2474 4627 2490 4648
rect 2490 4627 2520 4648
rect 3583 14984 3819 15187
rect 3583 14951 3613 14984
rect 3613 14951 3629 14984
rect 3629 14951 3693 14984
rect 3693 14951 3709 14984
rect 3709 14951 3773 14984
rect 3773 14951 3789 14984
rect 3789 14951 3819 14984
rect 3583 8068 3819 8304
rect 4882 18392 5118 18628
rect 4882 11510 5118 11746
rect 4882 4648 5118 4863
rect 4882 4627 4912 4648
rect 4912 4627 4928 4648
rect 4928 4627 4992 4648
rect 4992 4627 5008 4648
rect 5008 4627 5072 4648
rect 5072 4627 5088 4648
rect 5088 4627 5118 4648
rect 6180 14984 6416 15187
rect 6180 14951 6210 14984
rect 6210 14951 6226 14984
rect 6226 14951 6290 14984
rect 6290 14951 6306 14984
rect 6306 14951 6370 14984
rect 6370 14951 6386 14984
rect 6386 14951 6416 14984
rect 6180 8068 6416 8304
rect 7479 18392 7715 18628
rect 7479 11510 7715 11746
rect 7479 4648 7715 4863
rect 7479 4627 7509 4648
rect 7509 4627 7525 4648
rect 7525 4627 7589 4648
rect 7589 4627 7605 4648
rect 7605 4627 7669 4648
rect 7669 4627 7685 4648
rect 7685 4627 7715 4648
<< metal5 >>
rect 1104 18628 8832 18670
rect 1104 18392 2284 18628
rect 2520 18392 4882 18628
rect 5118 18392 7479 18628
rect 7715 18392 8832 18628
rect 1104 18350 8832 18392
rect 1104 15187 8832 15229
rect 1104 14951 3583 15187
rect 3819 14951 6180 15187
rect 6416 14951 8832 15187
rect 1104 14909 8832 14951
rect 1104 11746 8832 11788
rect 1104 11510 2284 11746
rect 2520 11510 4882 11746
rect 5118 11510 7479 11746
rect 7715 11510 8832 11746
rect 1104 11468 8832 11510
rect 1104 8304 8832 8347
rect 1104 8068 3583 8304
rect 3819 8068 6180 8304
rect 6416 8068 8832 8304
rect 1104 8026 8832 8068
rect 1104 4863 8832 4905
rect 1104 4627 2284 4863
rect 2520 4627 4882 4863
rect 5118 4627 7479 4863
rect 7715 4627 8832 4863
rect 1104 4585 8832 4627
use sky130_fd_sc_hd__decap_3  PHY_0 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 1104 0 -1 1896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604489732
transform 1 0 1104 0 1 1896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 1380 0 -1 1896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604489732
transform 1 0 2484 0 -1 1896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604489732
transform 1 0 1380 0 1 1896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604489732
transform 1 0 2484 0 1 1896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _055_ /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 4324 0 1 1896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 3956 0 -1 1896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 3588 0 -1 1896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604489732
transform 1 0 4048 0 -1 1896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604489732
transform 1 0 5152 0 -1 1896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_27 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 3588 0 1 1896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604489732
transform 1 0 4692 0 1 1896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604489732
transform 1 0 6808 0 -1 1896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604489732
transform 1 0 6716 0 1 1896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 6256 0 -1 1896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604489732
transform 1 0 6900 0 -1 1896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51
timestamp 1604489732
transform 1 0 5796 0 1 1896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 6532 0 1 1896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604489732
transform 1 0 6808 0 1 1896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_74
timestamp 1604489732
transform 1 0 7912 0 1 1896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604489732
transform -1 0 8832 0 -1 1896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604489732
transform -1 0 8832 0 1 1896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75
timestamp 1604489732
transform 1 0 8004 0 -1 1896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_80 /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 8464 0 1 1896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1604489732
transform 1 0 2852 0 -1 2984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604489732
transform 1 0 1104 0 -1 2984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604489732
transform 1 0 1380 0 -1 2984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1604489732
transform 1 0 2484 0 -1 2984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_23
timestamp 1604489732
transform 1 0 3220 0 -1 2984
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _079_ /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 4968 0 -1 2984
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604489732
transform 1 0 3956 0 -1 2984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_32
timestamp 1604489732
transform 1 0 4048 0 -1 2984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_40
timestamp 1604489732
transform 1 0 4784 0 -1 2984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_49
timestamp 1604489732
transform 1 0 5612 0 -1 2984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_61
timestamp 1604489732
transform 1 0 6716 0 -1 2984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_73
timestamp 1604489732
transform 1 0 7820 0 -1 2984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604489732
transform -1 0 8832 0 -1 2984
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _092_ /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 1380 0 1 2984
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604489732
transform 1 0 1104 0 1 2984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _039_ /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 4968 0 1 2984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_3_26
timestamp 1604489732
transform 1 0 3496 0 1 2984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_38
timestamp 1604489732
transform 1 0 4600 0 1 2984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_49
timestamp 1604489732
transform 1 0 5612 0 1 2984
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _078_ /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 6808 0 1 2984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604489732
transform 1 0 6716 0 1 2984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_65
timestamp 1604489732
transform 1 0 7084 0 1 2984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604489732
transform -1 0 8832 0 1 2984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_77
timestamp 1604489732
transform 1 0 8188 0 1 2984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1604489732
transform 1 0 2852 0 -1 4072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604489732
transform 1 0 1104 0 -1 4072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604489732
transform 1 0 1380 0 -1 4072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1604489732
transform 1 0 2484 0 -1 4072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_23
timestamp 1604489732
transform 1 0 3220 0 -1 4072
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _094_
timestamp 1604489732
transform 1 0 4048 0 -1 4072
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604489732
transform 1 0 3956 0 -1 4072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_55
timestamp 1604489732
transform 1 0 6164 0 -1 4072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_67
timestamp 1604489732
transform 1 0 7268 0 -1 4072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604489732
transform -1 0 8832 0 -1 4072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_79
timestamp 1604489732
transform 1 0 8372 0 -1 4072
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _093_
timestamp 1604489732
transform 1 0 2576 0 1 4072
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604489732
transform 1 0 1104 0 1 4072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604489732
transform 1 0 1380 0 1 4072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_15
timestamp 1604489732
transform 1 0 2484 0 1 4072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604489732
transform 1 0 4692 0 1 4072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604489732
transform 1 0 6716 0 1 4072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604489732
transform 1 0 5796 0 1 4072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604489732
transform 1 0 6532 0 1 4072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604489732
transform 1 0 6808 0 1 4072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_74
timestamp 1604489732
transform 1 0 7912 0 1 4072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604489732
transform -1 0 8832 0 1 4072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_80
timestamp 1604489732
transform 1 0 8464 0 1 4072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _047_
timestamp 1604489732
transform 1 0 2208 0 -1 5160
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _100_
timestamp 1604489732
transform 1 0 1380 0 1 5160
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604489732
transform 1 0 1104 0 -1 5160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604489732
transform 1 0 1104 0 1 5160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1604489732
transform 1 0 1380 0 -1 5160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_11
timestamp 1604489732
transform 1 0 2116 0 -1 5160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_16
timestamp 1604489732
transform 1 0 2576 0 -1 5160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _102_
timestamp 1604489732
transform 1 0 4048 0 -1 5160
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604489732
transform 1 0 3956 0 -1 5160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_28
timestamp 1604489732
transform 1 0 3680 0 -1 5160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_26
timestamp 1604489732
transform 1 0 3496 0 1 5160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_38
timestamp 1604489732
transform 1 0 4600 0 1 5160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604489732
transform 1 0 6716 0 1 5160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_55
timestamp 1604489732
transform 1 0 6164 0 -1 5160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_67
timestamp 1604489732
transform 1 0 7268 0 -1 5160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_50
timestamp 1604489732
transform 1 0 5704 0 1 5160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_58
timestamp 1604489732
transform 1 0 6440 0 1 5160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604489732
transform 1 0 6808 0 1 5160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_74
timestamp 1604489732
transform 1 0 7912 0 1 5160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604489732
transform -1 0 8832 0 -1 5160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604489732
transform -1 0 8832 0 1 5160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_79
timestamp 1604489732
transform 1 0 8372 0 -1 5160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_80
timestamp 1604489732
transform 1 0 8464 0 1 5160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _048_
timestamp 1604489732
transform 1 0 2116 0 -1 6248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604489732
transform 1 0 1104 0 -1 6248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1604489732
transform 1 0 1380 0 -1 6248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604489732
transform 1 0 2484 0 -1 6248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604489732
transform 1 0 3956 0 -1 6248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604489732
transform 1 0 3588 0 -1 6248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604489732
transform 1 0 4048 0 -1 6248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604489732
transform 1 0 5152 0 -1 6248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604489732
transform 1 0 6256 0 -1 6248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604489732
transform 1 0 7360 0 -1 6248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604489732
transform -1 0 8832 0 -1 6248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_80
timestamp 1604489732
transform 1 0 8464 0 -1 6248
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _101_
timestamp 1604489732
transform 1 0 1380 0 1 6248
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604489732
transform 1 0 1104 0 1 6248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _045_
timestamp 1604489732
transform 1 0 4232 0 1 6248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _054_
timestamp 1604489732
transform 1 0 5336 0 1 6248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_26
timestamp 1604489732
transform 1 0 3496 0 1 6248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_38
timestamp 1604489732
transform 1 0 4600 0 1 6248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604489732
transform 1 0 6716 0 1 6248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_50
timestamp 1604489732
transform 1 0 5704 0 1 6248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1604489732
transform 1 0 6440 0 1 6248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604489732
transform 1 0 6808 0 1 6248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_74
timestamp 1604489732
transform 1 0 7912 0 1 6248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604489732
transform -1 0 8832 0 1 6248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_80
timestamp 1604489732
transform 1 0 8464 0 1 6248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604489732
transform 1 0 1104 0 -1 7336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604489732
transform 1 0 1380 0 -1 7336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604489732
transform 1 0 2484 0 -1 7336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _095_
timestamp 1604489732
transform 1 0 4324 0 -1 7336
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604489732
transform 1 0 3956 0 -1 7336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604489732
transform 1 0 3588 0 -1 7336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_32
timestamp 1604489732
transform 1 0 4048 0 -1 7336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_58
timestamp 1604489732
transform 1 0 6440 0 -1 7336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_70
timestamp 1604489732
transform 1 0 7544 0 -1 7336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604489732
transform -1 0 8832 0 -1 7336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_78
timestamp 1604489732
transform 1 0 8280 0 -1 7336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _052_
timestamp 1604489732
transform 1 0 3312 0 1 7336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604489732
transform 1 0 1104 0 1 7336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604489732
transform 1 0 1380 0 1 7336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_15
timestamp 1604489732
transform 1 0 2484 0 1 7336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_23
timestamp 1604489732
transform 1 0 3220 0 1 7336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _040_
timestamp 1604489732
transform 1 0 4416 0 1 7336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _053_
timestamp 1604489732
transform 1 0 5520 0 1 7336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_28
timestamp 1604489732
transform 1 0 3680 0 1 7336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_40
timestamp 1604489732
transform 1 0 4784 0 1 7336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604489732
transform 1 0 6716 0 1 7336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_52
timestamp 1604489732
transform 1 0 5888 0 1 7336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1604489732
transform 1 0 6624 0 1 7336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604489732
transform 1 0 6808 0 1 7336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_74
timestamp 1604489732
transform 1 0 7912 0 1 7336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604489732
transform -1 0 8832 0 1 7336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_80
timestamp 1604489732
transform 1 0 8464 0 1 7336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _051_
timestamp 1604489732
transform 1 0 2852 0 -1 8424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604489732
transform 1 0 1104 0 -1 8424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_serial_clock /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 2576 0 -1 8424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604489732
transform 1 0 1380 0 -1 8424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_15
timestamp 1604489732
transform 1 0 2484 0 -1 8424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_23
timestamp 1604489732
transform 1 0 3220 0 -1 8424
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _096_
timestamp 1604489732
transform 1 0 4416 0 -1 8424
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604489732
transform 1 0 3956 0 -1 8424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1604489732
transform 1 0 4048 0 -1 8424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1604489732
transform 1 0 7268 0 -1 8424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_59
timestamp 1604489732
transform 1 0 6532 0 -1 8424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_71
timestamp 1604489732
transform 1 0 7636 0 -1 8424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604489732
transform -1 0 8832 0 -1 8424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_79
timestamp 1604489732
transform 1 0 8372 0 -1 8424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _046_
timestamp 1604489732
transform 1 0 2852 0 -1 9512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _050_
timestamp 1604489732
transform 1 0 1748 0 -1 9512
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _097_
timestamp 1604489732
transform 1 0 2484 0 1 8424
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604489732
transform 1 0 1104 0 1 8424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604489732
transform 1 0 1104 0 -1 9512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604489732
transform 1 0 1380 0 1 8424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1604489732
transform 1 0 1380 0 -1 9512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_11
timestamp 1604489732
transform 1 0 2116 0 -1 9512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_23
timestamp 1604489732
transform 1 0 3220 0 -1 9512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _041_
timestamp 1604489732
transform 1 0 5336 0 1 8424
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_4  _082_ /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 5060 0 -1 9512
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604489732
transform 1 0 3956 0 -1 9512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_38
timestamp 1604489732
transform 1 0 4600 0 1 8424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_32
timestamp 1604489732
transform 1 0 4048 0 -1 9512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_40
timestamp 1604489732
transform 1 0 4784 0 -1 9512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604489732
transform 1 0 6808 0 1 8424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604489732
transform 1 0 6716 0 1 8424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_50
timestamp 1604489732
transform 1 0 5704 0 1 8424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_58
timestamp 1604489732
transform 1 0 6440 0 1 8424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_66
timestamp 1604489732
transform 1 0 7176 0 1 8424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_67
timestamp 1604489732
transform 1 0 7268 0 -1 9512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604489732
transform -1 0 8832 0 1 8424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604489732
transform -1 0 8832 0 -1 9512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_78
timestamp 1604489732
transform 1 0 8280 0 1 8424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_79
timestamp 1604489732
transform 1 0 8372 0 -1 9512
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _083_
timestamp 1604489732
transform 1 0 1380 0 1 9512
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604489732
transform 1 0 1104 0 1 9512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_26
timestamp 1604489732
transform 1 0 3496 0 1 9512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_38
timestamp 1604489732
transform 1 0 4600 0 1 9512
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _080_
timestamp 1604489732
transform 1 0 7176 0 1 9512
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604489732
transform 1 0 6716 0 1 9512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_50
timestamp 1604489732
transform 1 0 5704 0 1 9512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_58
timestamp 1604489732
transform 1 0 6440 0 1 9512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1604489732
transform 1 0 6808 0 1 9512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_73
timestamp 1604489732
transform 1 0 7820 0 1 9512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604489732
transform -1 0 8832 0 1 9512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604489732
transform 1 0 2208 0 -1 10600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604489732
transform 1 0 1104 0 -1 10600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1604489732
transform 1 0 1380 0 -1 10600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_11
timestamp 1604489732
transform 1 0 2116 0 -1 10600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_16
timestamp 1604489732
transform 1 0 2576 0 -1 10600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604489732
transform 1 0 3956 0 -1 10600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_28
timestamp 1604489732
transform 1 0 3680 0 -1 10600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604489732
transform 1 0 4048 0 -1 10600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604489732
transform 1 0 5152 0 -1 10600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1604489732
transform 1 0 6256 0 -1 10600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1604489732
transform 1 0 7360 0 -1 10600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604489732
transform -1 0 8832 0 -1 10600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_80
timestamp 1604489732
transform 1 0 8464 0 -1 10600
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _098_
timestamp 1604489732
transform 1 0 1380 0 1 10600
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604489732
transform 1 0 1104 0 1 10600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 4232 0 1 10600
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_17_26
timestamp 1604489732
transform 1 0 3496 0 1 10600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604489732
transform 1 0 6716 0 1 10600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_54
timestamp 1604489732
transform 1 0 6072 0 1 10600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1604489732
transform 1 0 6624 0 1 10600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1604489732
transform 1 0 6808 0 1 10600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_74
timestamp 1604489732
transform 1 0 7912 0 1 10600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604489732
transform -1 0 8832 0 1 10600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_80
timestamp 1604489732
transform 1 0 8464 0 1 10600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _049_
timestamp 1604489732
transform 1 0 2116 0 -1 11688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604489732
transform 1 0 1104 0 -1 11688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1604489732
transform 1 0 1380 0 -1 11688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1604489732
transform 1 0 2484 0 -1 11688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1604489732
transform 1 0 5060 0 -1 11688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604489732
transform 1 0 3956 0 -1 11688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1604489732
transform 1 0 3588 0 -1 11688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_32
timestamp 1604489732
transform 1 0 4048 0 -1 11688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_40
timestamp 1604489732
transform 1 0 4784 0 -1 11688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_47
timestamp 1604489732
transform 1 0 5428 0 -1 11688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1604489732
transform 1 0 6164 0 -1 11688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_59
timestamp 1604489732
transform 1 0 6532 0 -1 11688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_71
timestamp 1604489732
transform 1 0 7636 0 -1 11688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604489732
transform -1 0 8832 0 -1 11688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_79
timestamp 1604489732
transform 1 0 8372 0 -1 11688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604489732
transform 1 0 1104 0 -1 12776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604489732
transform 1 0 1104 0 1 11688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_23
timestamp 1604489732
transform 1 0 3220 0 -1 12776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_15
timestamp 1604489732
transform 1 0 2484 0 -1 12776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_22
timestamp 1604489732
transform 1 0 3128 0 1 11688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_15
timestamp 1604489732
transform 1 0 2484 0 1 11688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604489732
transform 1 0 2760 0 1 11688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1604489732
transform 1 0 2852 0 -1 12776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604489732
transform 1 0 1380 0 -1 12776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604489732
transform 1 0 1380 0 1 11688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1604489732
transform 1 0 4048 0 -1 12776
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_4  _088_
timestamp 1604489732
transform 1 0 5152 0 -1 12776
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrtp_4  _091_
timestamp 1604489732
transform 1 0 3864 0 1 11688
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604489732
transform 1 0 3956 0 -1 12776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_36
timestamp 1604489732
transform 1 0 4416 0 -1 12776
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _072_
timestamp 1604489732
transform 1 0 6808 0 1 11688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604489732
transform 1 0 6716 0 1 11688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_53
timestamp 1604489732
transform 1 0 5980 0 1 11688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_65
timestamp 1604489732
transform 1 0 7084 0 1 11688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1604489732
transform 1 0 7360 0 -1 12776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604489732
transform -1 0 8832 0 1 11688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604489732
transform -1 0 8832 0 -1 12776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_77
timestamp 1604489732
transform 1 0 8188 0 1 11688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_80
timestamp 1604489732
transform 1 0 8464 0 -1 12776
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _087_
timestamp 1604489732
transform 1 0 1932 0 1 12776
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604489732
transform 1 0 1104 0 1 12776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1604489732
transform 1 0 1380 0 1 12776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1604489732
transform 1 0 4784 0 1 12776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_32
timestamp 1604489732
transform 1 0 4048 0 1 12776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_44
timestamp 1604489732
transform 1 0 5152 0 1 12776
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _073_ /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 6808 0 1 12776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604489732
transform 1 0 6716 0 1 12776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_56
timestamp 1604489732
transform 1 0 6256 0 1 12776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1604489732
transform 1 0 6624 0 1 12776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_71
timestamp 1604489732
transform 1 0 7636 0 1 12776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604489732
transform -1 0 8832 0 1 12776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_79
timestamp 1604489732
transform 1 0 8372 0 1 12776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604489732
transform 1 0 1104 0 -1 13864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_serial_clock
timestamp 1604489732
transform 1 0 3036 0 -1 13864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604489732
transform 1 0 1380 0 -1 13864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_15
timestamp 1604489732
transform 1 0 2484 0 -1 13864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_24
timestamp 1604489732
transform 1 0 3312 0 -1 13864
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_4  _090_
timestamp 1604489732
transform 1 0 4232 0 -1 13864
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604489732
transform 1 0 3956 0 -1 13864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_30
timestamp 1604489732
transform 1 0 3864 0 -1 13864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1604489732
transform 1 0 4048 0 -1 13864
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _074_
timestamp 1604489732
transform 1 0 7176 0 -1 13864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_22_57
timestamp 1604489732
transform 1 0 6348 0 -1 13864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_65
timestamp 1604489732
transform 1 0 7084 0 -1 13864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_73
timestamp 1604489732
transform 1 0 7820 0 -1 13864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604489732
transform -1 0 8832 0 -1 13864
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _086_
timestamp 1604489732
transform 1 0 1380 0 1 13864
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604489732
transform 1 0 1104 0 1 13864
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_4  _071_ /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 4416 0 1 13864
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_23_26
timestamp 1604489732
transform 1 0 3496 0 1 13864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_34
timestamp 1604489732
transform 1 0 4232 0 1 13864
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _075_ /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 6808 0 1 13864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604489732
transform 1 0 6716 0 1 13864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_53
timestamp 1604489732
transform 1 0 5980 0 1 13864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_71
timestamp 1604489732
transform 1 0 7636 0 1 13864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604489732
transform -1 0 8832 0 1 13864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_79
timestamp 1604489732
transform 1 0 8372 0 1 13864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1604489732
transform 1 0 2116 0 -1 14952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604489732
transform 1 0 1104 0 -1 14952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1604489732
transform 1 0 1380 0 -1 14952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604489732
transform 1 0 2484 0 -1 14952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _107_
timestamp 1604489732
transform 1 0 4048 0 -1 14952
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604489732
transform 1 0 3956 0 -1 14952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604489732
transform 1 0 3588 0 -1 14952
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _077_
timestamp 1604489732
transform 1 0 6992 0 -1 14952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_55
timestamp 1604489732
transform 1 0 6164 0 -1 14952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_63
timestamp 1604489732
transform 1 0 6900 0 -1 14952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_73
timestamp 1604489732
transform 1 0 7820 0 -1 14952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604489732
transform -1 0 8832 0 -1 14952
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _099_
timestamp 1604489732
transform 1 0 1380 0 1 14952
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604489732
transform 1 0 1104 0 1 14952
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_4  _076_
timestamp 1604489732
transform 1 0 4416 0 1 14952
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_25_26
timestamp 1604489732
transform 1 0 3496 0 1 14952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_34
timestamp 1604489732
transform 1 0 4232 0 1 14952
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _070_
timestamp 1604489732
transform 1 0 7544 0 1 14952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604489732
transform 1 0 6716 0 1 14952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_53
timestamp 1604489732
transform 1 0 5980 0 1 14952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_62
timestamp 1604489732
transform 1 0 6808 0 1 14952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_73
timestamp 1604489732
transform 1 0 7820 0 1 14952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604489732
transform -1 0 8832 0 1 14952
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _106_
timestamp 1604489732
transform 1 0 3128 0 1 16040
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604489732
transform 1 0 1104 0 -1 16040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604489732
transform 1 0 1104 0 1 16040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604489732
transform 1 0 1380 0 -1 16040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604489732
transform 1 0 2484 0 -1 16040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604489732
transform 1 0 1380 0 1 16040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_15
timestamp 1604489732
transform 1 0 2484 0 1 16040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_21
timestamp 1604489732
transform 1 0 3036 0 1 16040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1604489732
transform 1 0 5060 0 -1 16040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604489732
transform 1 0 3956 0 -1 16040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604489732
transform 1 0 3588 0 -1 16040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_32
timestamp 1604489732
transform 1 0 4048 0 -1 16040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_40
timestamp 1604489732
transform 1 0 4784 0 -1 16040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_47
timestamp 1604489732
transform 1 0 5428 0 -1 16040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_45
timestamp 1604489732
transform 1 0 5244 0 1 16040
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  gpio_in_buf /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 6164 0 -1 16040
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604489732
transform 1 0 6716 0 1 16040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_73
timestamp 1604489732
transform 1 0 7820 0 -1 16040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1604489732
transform 1 0 6348 0 1 16040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604489732
transform 1 0 6808 0 1 16040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_74
timestamp 1604489732
transform 1 0 7912 0 1 16040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604489732
transform -1 0 8832 0 -1 16040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604489732
transform -1 0 8832 0 1 16040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_80
timestamp 1604489732
transform 1 0 8464 0 1 16040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604489732
transform 1 0 1104 0 -1 17128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604489732
transform 1 0 1380 0 -1 17128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604489732
transform 1 0 2484 0 -1 17128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfstp_4  _089_
timestamp 1604489732
transform 1 0 4140 0 -1 17128
box -38 -48 2246 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604489732
transform 1 0 3956 0 -1 17128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604489732
transform 1 0 3588 0 -1 17128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_32
timestamp 1604489732
transform 1 0 4048 0 -1 17128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  gpio_logic_high /home/xrex/usr/devel/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604489732
transform 1 0 7084 0 -1 17128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_57
timestamp 1604489732
transform 1 0 6348 0 -1 17128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604489732
transform 1 0 7360 0 -1 17128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604489732
transform -1 0 8832 0 -1 17128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_80
timestamp 1604489732
transform 1 0 8464 0 -1 17128
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _104_
timestamp 1604489732
transform 1 0 1380 0 1 17128
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604489732
transform 1 0 1104 0 1 17128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_26
timestamp 1604489732
transform 1 0 3496 0 1 17128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_38
timestamp 1604489732
transform 1 0 4600 0 1 17128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604489732
transform 1 0 6716 0 1 17128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_50
timestamp 1604489732
transform 1 0 5704 0 1 17128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_58
timestamp 1604489732
transform 1 0 6440 0 1 17128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604489732
transform 1 0 6808 0 1 17128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_74
timestamp 1604489732
transform 1 0 7912 0 1 17128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604489732
transform -1 0 8832 0 1 17128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_80
timestamp 1604489732
transform 1 0 8464 0 1 17128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _043_
timestamp 1604489732
transform 1 0 2852 0 -1 18216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604489732
transform 1 0 1748 0 -1 18216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604489732
transform 1 0 1104 0 -1 18216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1604489732
transform 1 0 1380 0 -1 18216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_11
timestamp 1604489732
transform 1 0 2116 0 -1 18216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_23
timestamp 1604489732
transform 1 0 3220 0 -1 18216
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _105_
timestamp 1604489732
transform 1 0 4048 0 -1 18216
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604489732
transform 1 0 3956 0 -1 18216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_55
timestamp 1604489732
transform 1 0 6164 0 -1 18216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_67
timestamp 1604489732
transform 1 0 7268 0 -1 18216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604489732
transform -1 0 8832 0 -1 18216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_79
timestamp 1604489732
transform 1 0 8372 0 -1 18216
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _084_
timestamp 1604489732
transform 1 0 1380 0 1 18216
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604489732
transform 1 0 1104 0 1 18216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _042_
timestamp 1604489732
transform 1 0 4232 0 1 18216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _044_
timestamp 1604489732
transform 1 0 5336 0 1 18216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_26
timestamp 1604489732
transform 1 0 3496 0 1 18216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_38
timestamp 1604489732
transform 1 0 4600 0 1 18216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604489732
transform 1 0 6716 0 1 18216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_50
timestamp 1604489732
transform 1 0 5704 0 1 18216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_58
timestamp 1604489732
transform 1 0 6440 0 1 18216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604489732
transform 1 0 6808 0 1 18216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_74
timestamp 1604489732
transform 1 0 7912 0 1 18216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604489732
transform -1 0 8832 0 1 18216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_80
timestamp 1604489732
transform 1 0 8464 0 1 18216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604489732
transform 1 0 2116 0 -1 19304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604489732
transform 1 0 1104 0 -1 19304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1604489732
transform 1 0 1380 0 -1 19304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604489732
transform 1 0 2484 0 -1 19304
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_4  _103_
timestamp 1604489732
transform 1 0 4048 0 -1 19304
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604489732
transform 1 0 3956 0 -1 19304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604489732
transform 1 0 3588 0 -1 19304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_55
timestamp 1604489732
transform 1 0 6164 0 -1 19304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_67
timestamp 1604489732
transform 1 0 7268 0 -1 19304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604489732
transform -1 0 8832 0 -1 19304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_79
timestamp 1604489732
transform 1 0 8372 0 -1 19304
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _085_
timestamp 1604489732
transform 1 0 1380 0 1 19304
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604489732
transform 1 0 1104 0 1 19304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604489732
transform 1 0 1104 0 -1 20392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604489732
transform 1 0 1380 0 -1 20392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604489732
transform 1 0 2484 0 -1 20392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604489732
transform 1 0 3956 0 -1 20392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_26
timestamp 1604489732
transform 1 0 3496 0 1 19304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_38
timestamp 1604489732
transform 1 0 4600 0 1 19304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604489732
transform 1 0 3588 0 -1 20392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604489732
transform 1 0 4048 0 -1 20392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604489732
transform 1 0 5152 0 -1 20392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604489732
transform 1 0 6716 0 1 19304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_50
timestamp 1604489732
transform 1 0 5704 0 1 19304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_58
timestamp 1604489732
transform 1 0 6440 0 1 19304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1604489732
transform 1 0 6808 0 1 19304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_74
timestamp 1604489732
transform 1 0 7912 0 1 19304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604489732
transform 1 0 6256 0 -1 20392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604489732
transform 1 0 7360 0 -1 20392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604489732
transform -1 0 8832 0 1 19304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604489732
transform -1 0 8832 0 -1 20392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_80
timestamp 1604489732
transform 1 0 8464 0 1 19304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_80
timestamp 1604489732
transform 1 0 8464 0 -1 20392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604489732
transform 1 0 1104 0 1 20392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604489732
transform 1 0 1380 0 1 20392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604489732
transform 1 0 2484 0 1 20392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1604489732
transform 1 0 3588 0 1 20392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1604489732
transform 1 0 4692 0 1 20392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604489732
transform 1 0 6716 0 1 20392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1604489732
transform 1 0 5796 0 1 20392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1604489732
transform 1 0 6532 0 1 20392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1604489732
transform 1 0 6808 0 1 20392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_74
timestamp 1604489732
transform 1 0 7912 0 1 20392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604489732
transform -1 0 8832 0 1 20392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_80
timestamp 1604489732
transform 1 0 8464 0 1 20392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604489732
transform 1 0 1104 0 -1 21480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604489732
transform 1 0 1380 0 -1 21480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604489732
transform 1 0 2484 0 -1 21480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604489732
transform 1 0 3956 0 -1 21480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1604489732
transform 1 0 3588 0 -1 21480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1604489732
transform 1 0 4048 0 -1 21480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1604489732
transform 1 0 5152 0 -1 21480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604489732
transform 1 0 6808 0 -1 21480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_56
timestamp 1604489732
transform 1 0 6256 0 -1 21480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_63
timestamp 1604489732
transform 1 0 6900 0 -1 21480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604489732
transform -1 0 8832 0 -1 21480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_75
timestamp 1604489732
transform 1 0 8004 0 -1 21480
box -38 -48 590 592
<< labels >>
rlabel metal3 s 9520 8840 10000 8960 6 mgmt_gpio_in
port 0 nsew default tristate
rlabel metal3 s 9520 11560 10000 11680 6 mgmt_gpio_oeb
port 1 nsew default input
rlabel metal3 s 9520 14416 10000 14536 6 mgmt_gpio_out
port 2 nsew default input
rlabel metal3 s 0 0 480 120 6 pad_gpio_ana_en
port 3 nsew default tristate
rlabel metal3 s 0 1632 480 1752 6 pad_gpio_ana_pol
port 4 nsew default tristate
rlabel metal3 s 0 3264 480 3384 6 pad_gpio_ana_sel
port 5 nsew default tristate
rlabel metal3 s 0 4896 480 5016 6 pad_gpio_dm[0]
port 6 nsew default tristate
rlabel metal3 s 0 6664 480 6784 6 pad_gpio_dm[1]
port 7 nsew default tristate
rlabel metal3 s 0 8296 480 8416 6 pad_gpio_dm[2]
port 8 nsew default tristate
rlabel metal3 s 0 9928 480 10048 6 pad_gpio_holdover
port 9 nsew default tristate
rlabel metal3 s 0 11560 480 11680 6 pad_gpio_ib_mode_sel
port 10 nsew default tristate
rlabel metal3 s 0 13328 480 13448 6 pad_gpio_in
port 11 nsew default input
rlabel metal3 s 0 14960 480 15080 6 pad_gpio_inenb
port 12 nsew default tristate
rlabel metal3 s 0 16592 480 16712 6 pad_gpio_out
port 13 nsew default tristate
rlabel metal3 s 0 18224 480 18344 6 pad_gpio_outenb
port 14 nsew default tristate
rlabel metal3 s 0 19992 480 20112 6 pad_gpio_slow_sel
port 15 nsew default tristate
rlabel metal3 s 0 21624 480 21744 6 pad_gpio_vtrip_sel
port 16 nsew default tristate
rlabel metal3 s 9520 544 10000 664 6 resetn
port 17 nsew default input
rlabel metal3 s 9520 3264 10000 3384 6 serial_clock
port 18 nsew default input
rlabel metal3 s 9520 5984 10000 6104 6 serial_data_in
port 19 nsew default input
rlabel metal3 s 0 23256 480 23376 6 serial_data_out
port 20 nsew default tristate
rlabel metal3 s 9520 17136 10000 17256 6 user_gpio_in
port 21 nsew default tristate
rlabel metal3 s 9520 19992 10000 20112 6 user_gpio_oeb
port 22 nsew default input
rlabel metal3 s 9520 22712 10000 22832 6 user_gpio_out
port 23 nsew default input
rlabel metal5 s 1104 4585 8832 4905 6 VPWR
port 24 nsew default input
rlabel metal5 s 1104 8027 8832 8347 6 VGND
port 25 nsew default input
<< properties >>
string FIXED_BBOX 0 0 10000 23376
<< end >>
