magic
tech sky130A
magscale 1 2
timestamp 1625003591
<< metal1 >>
rect 287920 993609 287926 993661
rect 287978 993649 287984 993661
rect 291280 993649 291286 993661
rect 287978 993621 291286 993649
rect 287978 993609 287984 993621
rect 291280 993609 291286 993621
rect 291338 993609 291344 993661
rect 175600 992795 175606 992847
rect 175658 992835 175664 992847
rect 178480 992835 178486 992847
rect 175658 992807 178486 992835
rect 175658 992795 175664 992807
rect 178480 992795 178486 992807
rect 178538 992795 178544 992847
rect 129520 984951 129526 985003
rect 129578 984991 129584 985003
rect 132400 984991 132406 985003
rect 129578 984963 132406 984991
rect 129578 984951 129584 984963
rect 132400 984951 132406 984963
rect 132458 984951 132464 985003
rect 399568 983471 399574 983523
rect 399626 983511 399632 983523
rect 432016 983511 432022 983523
rect 399626 983483 432022 983511
rect 399626 983471 399632 983483
rect 432016 983471 432022 983483
rect 432074 983471 432080 983523
rect 578866 983039 610574 983067
rect 178576 982953 178582 983005
rect 178634 982993 178640 983005
rect 184240 982993 184246 983005
rect 178634 982965 184246 982993
rect 178634 982953 178640 982965
rect 184240 982953 184246 982965
rect 184298 982953 184304 983005
rect 392464 982879 392470 982931
rect 392522 982919 392528 982931
rect 578866 982919 578894 983039
rect 392522 982891 578894 982919
rect 588994 982965 590414 982993
rect 392522 982879 392528 982891
rect 394576 982805 394582 982857
rect 394634 982845 394640 982857
rect 588994 982845 589022 982965
rect 394634 982817 589022 982845
rect 590386 982845 590414 982965
rect 610546 982919 610574 983039
rect 649456 982919 649462 982931
rect 610546 982891 649462 982919
rect 649456 982879 649462 982891
rect 649514 982879 649520 982931
rect 590386 982817 649406 982845
rect 394634 982805 394640 982817
rect 649378 982031 649406 982817
rect 652240 982031 652246 982043
rect 649378 982003 652246 982031
rect 652240 981991 652246 982003
rect 652298 981991 652304 982043
rect 649456 981917 649462 981969
rect 649514 981957 649520 981969
rect 656656 981957 656662 981969
rect 649514 981929 656662 981957
rect 649514 981917 649520 981929
rect 656656 981917 656662 981929
rect 656714 981917 656720 981969
rect 652240 979179 652246 979231
rect 652298 979219 652304 979231
rect 679696 979219 679702 979231
rect 652298 979191 679702 979219
rect 652298 979179 652304 979191
rect 679696 979179 679702 979191
rect 679754 979179 679760 979231
rect 656656 974887 656662 974939
rect 656714 974927 656720 974939
rect 671056 974927 671062 974939
rect 656714 974899 671062 974927
rect 656714 974887 656720 974899
rect 671056 974887 671062 974899
rect 671114 974887 671120 974939
rect 671056 963935 671062 963987
rect 671114 963975 671120 963987
rect 677584 963975 677590 963987
rect 671114 963947 677590 963975
rect 671114 963935 671120 963947
rect 677584 963935 677590 963947
rect 677642 963935 677648 963987
rect 40144 961863 40150 961915
rect 40202 961903 40208 961915
rect 60016 961903 60022 961915
rect 40202 961875 60022 961903
rect 40202 961863 40208 961875
rect 60016 961863 60022 961875
rect 60074 961863 60080 961915
rect 677488 959051 677494 959103
rect 677546 959091 677552 959103
rect 679696 959091 679702 959103
rect 677546 959063 679702 959091
rect 677546 959051 677552 959063
rect 679696 959051 679702 959063
rect 679754 959051 679760 959103
rect 653776 944325 653782 944377
rect 653834 944365 653840 944377
rect 676816 944365 676822 944377
rect 653834 944337 676822 944365
rect 653834 944325 653840 944337
rect 676816 944325 676822 944337
rect 676874 944325 676880 944377
rect 654256 878613 654262 878665
rect 654314 878653 654320 878665
rect 676240 878653 676246 878665
rect 654314 878625 676246 878653
rect 654314 878613 654320 878625
rect 676240 878613 676246 878625
rect 676298 878613 676304 878665
rect 654160 878539 654166 878591
rect 654218 878579 654224 878591
rect 676144 878579 676150 878591
rect 654218 878551 676150 878579
rect 654218 878539 654224 878551
rect 676144 878539 676150 878551
rect 676202 878539 676208 878591
rect 654064 878465 654070 878517
rect 654122 878505 654128 878517
rect 676336 878505 676342 878517
rect 654122 878477 676342 878505
rect 654122 878465 654128 878477
rect 676336 878465 676342 878477
rect 676394 878465 676400 878517
rect 673360 878391 673366 878443
rect 673418 878431 673424 878443
rect 676048 878431 676054 878443
rect 673418 878403 676054 878431
rect 673418 878391 673424 878403
rect 676048 878391 676054 878403
rect 676106 878391 676112 878443
rect 670864 877207 670870 877259
rect 670922 877247 670928 877259
rect 676240 877247 676246 877259
rect 670922 877219 676246 877247
rect 670922 877207 670928 877219
rect 676240 877207 676246 877219
rect 676298 877207 676304 877259
rect 670960 876171 670966 876223
rect 671018 876211 671024 876223
rect 676240 876211 676246 876223
rect 671018 876183 676246 876211
rect 671018 876171 671024 876183
rect 676240 876171 676246 876183
rect 676298 876171 676304 876223
rect 674032 872693 674038 872745
rect 674090 872733 674096 872745
rect 676240 872733 676246 872745
rect 674090 872705 676246 872733
rect 674090 872693 674096 872705
rect 676240 872693 676246 872705
rect 676298 872693 676304 872745
rect 674320 872619 674326 872671
rect 674378 872659 674384 872671
rect 676048 872659 676054 872671
rect 674378 872631 676054 872659
rect 674378 872619 674384 872631
rect 676048 872619 676054 872631
rect 676106 872619 676112 872671
rect 674128 870103 674134 870155
rect 674186 870143 674192 870155
rect 676048 870143 676054 870155
rect 674186 870115 676054 870143
rect 674186 870103 674192 870115
rect 676048 870103 676054 870115
rect 676106 870103 676112 870155
rect 674896 869881 674902 869933
rect 674954 869921 674960 869933
rect 676240 869921 676246 869933
rect 674954 869893 676246 869921
rect 674954 869881 674960 869893
rect 676240 869881 676246 869893
rect 676298 869881 676304 869933
rect 675088 869807 675094 869859
rect 675146 869847 675152 869859
rect 676048 869847 676054 869859
rect 675146 869819 676054 869847
rect 675146 869807 675152 869819
rect 676048 869807 676054 869819
rect 676106 869807 676112 869859
rect 674992 869733 674998 869785
rect 675050 869773 675056 869785
rect 679696 869773 679702 869785
rect 675050 869745 679702 869773
rect 675050 869733 675056 869745
rect 679696 869733 679702 869745
rect 679754 869733 679760 869785
rect 675184 869659 675190 869711
rect 675242 869699 675248 869711
rect 679792 869699 679798 869711
rect 675242 869671 679798 869699
rect 675242 869659 675248 869671
rect 679792 869659 679798 869671
rect 679850 869659 679856 869711
rect 674512 866995 674518 867047
rect 674570 867035 674576 867047
rect 676240 867035 676246 867047
rect 674570 867007 676246 867035
rect 674570 866995 674576 867007
rect 676240 866995 676246 867007
rect 676298 866995 676304 867047
rect 649456 866921 649462 866973
rect 649514 866961 649520 866973
rect 679792 866961 679798 866973
rect 649514 866933 679798 866961
rect 649514 866921 649520 866933
rect 679792 866921 679798 866933
rect 679850 866921 679856 866973
rect 674608 864257 674614 864309
rect 674666 864297 674672 864309
rect 679888 864297 679894 864309
rect 674666 864269 679894 864297
rect 674666 864257 674672 864269
rect 679888 864257 679894 864269
rect 679946 864257 679952 864309
rect 674992 864183 674998 864235
rect 675050 864223 675056 864235
rect 680176 864223 680182 864235
rect 675050 864195 680182 864223
rect 675050 864183 675056 864195
rect 680176 864183 680182 864195
rect 680234 864183 680240 864235
rect 675280 864109 675286 864161
rect 675338 864149 675344 864161
rect 680272 864149 680278 864161
rect 675338 864121 680278 864149
rect 675338 864109 675344 864121
rect 680272 864109 680278 864121
rect 680330 864109 680336 864161
rect 654256 864035 654262 864087
rect 654314 864075 654320 864087
rect 675472 864075 675478 864087
rect 654314 864047 675478 864075
rect 654314 864035 654320 864047
rect 675472 864035 675478 864047
rect 675530 864035 675536 864087
rect 674224 863147 674230 863199
rect 674282 863187 674288 863199
rect 680080 863187 680086 863199
rect 674282 863159 680086 863187
rect 674282 863147 674288 863159
rect 680080 863147 680086 863159
rect 680138 863147 680144 863199
rect 674416 863073 674422 863125
rect 674474 863113 674480 863125
rect 679984 863113 679990 863125
rect 674474 863085 679990 863113
rect 674474 863073 674480 863085
rect 679984 863073 679990 863085
rect 680042 863073 680048 863125
rect 675184 862407 675190 862459
rect 675242 862447 675248 862459
rect 675376 862447 675382 862459
rect 675242 862419 675382 862447
rect 675242 862407 675248 862419
rect 675376 862407 675382 862419
rect 675434 862407 675440 862459
rect 674896 861963 674902 862015
rect 674954 862003 674960 862015
rect 675376 862003 675382 862015
rect 674954 861975 675382 862003
rect 674954 861963 674960 861975
rect 675376 861963 675382 861975
rect 675434 861963 675440 862015
rect 674608 861815 674614 861867
rect 674666 861855 674672 861867
rect 674896 861855 674902 861867
rect 674666 861827 674902 861855
rect 674666 861815 674672 861827
rect 674896 861815 674902 861827
rect 674954 861815 674960 861867
rect 656368 861223 656374 861275
rect 656426 861263 656432 861275
rect 674608 861263 674614 861275
rect 656426 861235 674614 861263
rect 656426 861223 656432 861235
rect 674608 861223 674614 861235
rect 674666 861223 674672 861275
rect 654832 861149 654838 861201
rect 654890 861189 654896 861201
rect 675184 861189 675190 861201
rect 654890 861161 675190 861189
rect 654890 861149 654896 861161
rect 675184 861149 675190 861161
rect 675242 861149 675248 861201
rect 674992 859521 674998 859573
rect 675050 859561 675056 859573
rect 675472 859561 675478 859573
rect 675050 859533 675478 859561
rect 675050 859521 675056 859533
rect 675472 859521 675478 859533
rect 675530 859521 675536 859573
rect 674896 858707 674902 858759
rect 674954 858747 674960 858759
rect 675376 858747 675382 858759
rect 674954 858719 675382 858747
rect 674954 858707 674960 858719
rect 675376 858707 675382 858719
rect 675434 858707 675440 858759
rect 674032 858263 674038 858315
rect 674090 858303 674096 858315
rect 674992 858303 674998 858315
rect 674090 858275 674998 858303
rect 674090 858263 674096 858275
rect 674992 858263 674998 858275
rect 675050 858263 675056 858315
rect 674224 858115 674230 858167
rect 674282 858155 674288 858167
rect 675472 858155 675478 858167
rect 674282 858127 675478 858155
rect 674282 858115 674288 858127
rect 675472 858115 675478 858127
rect 675530 858115 675536 858167
rect 674416 857671 674422 857723
rect 674474 857711 674480 857723
rect 675376 857711 675382 857723
rect 674474 857683 675382 857711
rect 674474 857671 674480 857683
rect 675376 857671 675382 857683
rect 675434 857671 675440 857723
rect 674992 855155 674998 855207
rect 675050 855195 675056 855207
rect 675376 855195 675382 855207
rect 675050 855167 675382 855195
rect 675050 855155 675056 855167
rect 675376 855155 675382 855167
rect 675434 855155 675440 855207
rect 675088 854489 675094 854541
rect 675146 854529 675152 854541
rect 675376 854529 675382 854541
rect 675146 854501 675382 854529
rect 675146 854489 675152 854501
rect 675376 854489 675382 854501
rect 675434 854489 675440 854541
rect 674896 853971 674902 854023
rect 674954 854011 674960 854023
rect 675376 854011 675382 854023
rect 674954 853983 675382 854011
rect 674954 853971 674960 853983
rect 675376 853971 675382 853983
rect 675434 853971 675440 854023
rect 674512 853157 674518 853209
rect 674570 853197 674576 853209
rect 675472 853197 675478 853209
rect 674570 853169 675478 853197
rect 674570 853157 674576 853169
rect 675472 853157 675478 853169
rect 675530 853157 675536 853209
rect 675184 852713 675190 852765
rect 675242 852753 675248 852765
rect 675376 852753 675382 852765
rect 675242 852725 675382 852753
rect 675242 852713 675248 852725
rect 675376 852713 675382 852725
rect 675434 852713 675440 852765
rect 674128 852121 674134 852173
rect 674186 852161 674192 852173
rect 675376 852161 675382 852173
rect 674186 852133 675382 852161
rect 674186 852121 674192 852133
rect 675376 852121 675382 852133
rect 675434 852121 675440 852173
rect 674608 850863 674614 850915
rect 674666 850903 674672 850915
rect 675376 850903 675382 850915
rect 674666 850875 675382 850903
rect 674666 850863 674672 850875
rect 675376 850863 675382 850875
rect 675434 850863 675440 850915
rect 674320 850123 674326 850175
rect 674378 850163 674384 850175
rect 675472 850163 675478 850175
rect 674378 850135 675478 850163
rect 674378 850123 674384 850135
rect 675472 850123 675478 850135
rect 675530 850123 675536 850175
rect 675184 848421 675190 848473
rect 675242 848461 675248 848473
rect 675472 848461 675478 848473
rect 675242 848433 675478 848461
rect 675242 848421 675248 848433
rect 675472 848421 675478 848433
rect 675530 848421 675536 848473
rect 41776 817933 41782 817985
rect 41834 817973 41840 817985
rect 47536 817973 47542 817985
rect 41834 817945 47542 817973
rect 41834 817933 41840 817945
rect 47536 817933 47542 817945
rect 47594 817933 47600 817985
rect 41776 817267 41782 817319
rect 41834 817307 41840 817319
rect 44752 817307 44758 817319
rect 41834 817279 44758 817307
rect 41834 817267 41840 817279
rect 44752 817267 44758 817279
rect 44810 817267 44816 817319
rect 41584 816527 41590 816579
rect 41642 816567 41648 816579
rect 44848 816567 44854 816579
rect 41642 816539 44854 816567
rect 41642 816527 41648 816539
rect 44848 816527 44854 816539
rect 44906 816527 44912 816579
rect 41776 815787 41782 815839
rect 41834 815827 41840 815839
rect 43216 815827 43222 815839
rect 41834 815799 43222 815827
rect 41834 815787 41840 815799
rect 43216 815787 43222 815799
rect 43274 815787 43280 815839
rect 41776 814825 41782 814877
rect 41834 814865 41840 814877
rect 44656 814865 44662 814877
rect 41834 814837 44662 814865
rect 41834 814825 41840 814837
rect 44656 814825 44662 814837
rect 44714 814825 44720 814877
rect 41584 813567 41590 813619
rect 41642 813607 41648 813619
rect 44560 813607 44566 813619
rect 41642 813579 44566 813607
rect 41642 813567 41648 813579
rect 44560 813567 44566 813579
rect 44618 813567 44624 813619
rect 41872 808757 41878 808809
rect 41930 808797 41936 808809
rect 42736 808797 42742 808809
rect 41930 808769 42742 808797
rect 41930 808757 41936 808769
rect 42736 808757 42742 808769
rect 42794 808757 42800 808809
rect 41872 807055 41878 807107
rect 41930 807095 41936 807107
rect 43024 807095 43030 807107
rect 41930 807067 43030 807095
rect 41930 807055 41936 807067
rect 43024 807055 43030 807067
rect 43082 807055 43088 807107
rect 41392 806981 41398 807033
rect 41450 807021 41456 807033
rect 43120 807021 43126 807033
rect 41450 806993 43126 807021
rect 41450 806981 41456 806993
rect 43120 806981 43126 806993
rect 43178 806981 43184 807033
rect 41584 806759 41590 806811
rect 41642 806799 41648 806811
rect 42832 806799 42838 806811
rect 41642 806771 42838 806799
rect 41642 806759 41648 806771
rect 42832 806759 42838 806771
rect 42890 806759 42896 806811
rect 41584 806463 41590 806515
rect 41642 806503 41648 806515
rect 42928 806503 42934 806515
rect 41642 806475 42934 806503
rect 41642 806463 41648 806475
rect 42928 806463 42934 806475
rect 42986 806463 42992 806515
rect 37360 806315 37366 806367
rect 37418 806355 37424 806367
rect 42640 806355 42646 806367
rect 37418 806327 42646 806355
rect 37418 806315 37424 806327
rect 42640 806315 42646 806327
rect 42698 806315 42704 806367
rect 41584 805131 41590 805183
rect 41642 805171 41648 805183
rect 47440 805171 47446 805183
rect 41642 805143 47446 805171
rect 41642 805131 41648 805143
rect 47440 805131 47446 805143
rect 47498 805131 47504 805183
rect 34384 804909 34390 804961
rect 34442 804949 34448 804961
rect 41872 804949 41878 804961
rect 34442 804921 41878 804949
rect 34442 804909 34448 804921
rect 41872 804909 41878 804921
rect 41930 804909 41936 804961
rect 40144 801357 40150 801409
rect 40202 801397 40208 801409
rect 43408 801397 43414 801409
rect 40202 801369 43414 801397
rect 40202 801357 40208 801369
rect 43408 801357 43414 801369
rect 43466 801357 43472 801409
rect 40240 801283 40246 801335
rect 40298 801323 40304 801335
rect 43312 801323 43318 801335
rect 40298 801295 43318 801323
rect 40298 801283 40304 801295
rect 43312 801283 43318 801295
rect 43370 801283 43376 801335
rect 41968 801061 41974 801113
rect 42026 801101 42032 801113
rect 43504 801101 43510 801113
rect 42026 801073 43510 801101
rect 42026 801061 42032 801073
rect 43504 801061 43510 801073
rect 43562 801061 43568 801113
rect 41776 800987 41782 801039
rect 41834 800987 41840 801039
rect 42064 800987 42070 801039
rect 42122 801027 42128 801039
rect 42122 800999 42206 801027
rect 42122 800987 42128 800999
rect 41794 800817 41822 800987
rect 42178 800879 42206 800999
rect 42178 800851 42686 800879
rect 41776 800765 41782 800817
rect 41834 800765 41840 800817
rect 42658 800669 42686 800851
rect 43024 800765 43030 800817
rect 43082 800805 43088 800817
rect 43600 800805 43606 800817
rect 43082 800777 43606 800805
rect 43082 800765 43088 800777
rect 43600 800765 43606 800777
rect 43658 800765 43664 800817
rect 42640 800617 42646 800669
rect 42698 800617 42704 800669
rect 43024 800617 43030 800669
rect 43082 800657 43088 800669
rect 57616 800657 57622 800669
rect 43082 800629 57622 800657
rect 43082 800617 43088 800629
rect 57616 800617 57622 800629
rect 57674 800617 57680 800669
rect 43120 800543 43126 800595
rect 43178 800583 43184 800595
rect 43178 800555 43454 800583
rect 43178 800543 43184 800555
rect 43426 800521 43454 800555
rect 43408 800469 43414 800521
rect 43466 800469 43472 800521
rect 43312 799211 43318 799263
rect 43370 799251 43376 799263
rect 43600 799251 43606 799263
rect 43370 799223 43606 799251
rect 43370 799211 43376 799223
rect 43600 799211 43606 799223
rect 43658 799211 43664 799263
rect 42160 798915 42166 798967
rect 42218 798955 42224 798967
rect 42640 798955 42646 798967
rect 42218 798927 42646 798955
rect 42218 798915 42224 798927
rect 42640 798915 42646 798927
rect 42698 798915 42704 798967
rect 42160 797879 42166 797931
rect 42218 797919 42224 797931
rect 43312 797919 43318 797931
rect 42218 797891 43318 797919
rect 42218 797879 42224 797891
rect 43312 797879 43318 797891
rect 43370 797879 43376 797931
rect 42160 797065 42166 797117
rect 42218 797105 42224 797117
rect 42736 797105 42742 797117
rect 42218 797077 42742 797105
rect 42218 797065 42224 797077
rect 42736 797065 42742 797077
rect 42794 797065 42800 797117
rect 42736 796917 42742 796969
rect 42794 796957 42800 796969
rect 43504 796957 43510 796969
rect 42794 796929 43510 796957
rect 42794 796917 42800 796929
rect 43504 796917 43510 796929
rect 43562 796917 43568 796969
rect 42064 796251 42070 796303
rect 42122 796291 42128 796303
rect 43024 796291 43030 796303
rect 42122 796263 43030 796291
rect 42122 796251 42128 796263
rect 43024 796251 43030 796263
rect 43082 796251 43088 796303
rect 43024 796103 43030 796155
rect 43082 796143 43088 796155
rect 43408 796143 43414 796155
rect 43082 796115 43414 796143
rect 43082 796103 43088 796115
rect 43408 796103 43414 796115
rect 43466 796103 43472 796155
rect 42160 795659 42166 795711
rect 42218 795699 42224 795711
rect 42928 795699 42934 795711
rect 42218 795671 42934 795699
rect 42218 795659 42224 795671
rect 42928 795659 42934 795671
rect 42986 795659 42992 795711
rect 42640 795511 42646 795563
rect 42698 795551 42704 795563
rect 42928 795551 42934 795563
rect 42698 795523 42934 795551
rect 42698 795511 42704 795523
rect 42928 795511 42934 795523
rect 42986 795511 42992 795563
rect 42160 795215 42166 795267
rect 42218 795255 42224 795267
rect 42832 795255 42838 795267
rect 42218 795227 42838 795255
rect 42218 795215 42224 795227
rect 42832 795215 42838 795227
rect 42890 795215 42896 795267
rect 42832 795067 42838 795119
rect 42890 795107 42896 795119
rect 43600 795107 43606 795119
rect 42890 795079 43606 795107
rect 42890 795067 42896 795079
rect 43600 795067 43606 795079
rect 43658 795067 43664 795119
rect 42640 794919 42646 794971
rect 42698 794959 42704 794971
rect 43696 794959 43702 794971
rect 42698 794931 43702 794959
rect 42698 794919 42704 794931
rect 43696 794919 43702 794931
rect 43754 794919 43760 794971
rect 42064 794475 42070 794527
rect 42122 794515 42128 794527
rect 43024 794515 43030 794527
rect 42122 794487 43030 794515
rect 42122 794475 42128 794487
rect 43024 794475 43030 794487
rect 43082 794475 43088 794527
rect 42160 793735 42166 793787
rect 42218 793775 42224 793787
rect 42736 793775 42742 793787
rect 42218 793747 42742 793775
rect 42218 793735 42224 793747
rect 42736 793735 42742 793747
rect 42794 793735 42800 793787
rect 42640 792107 42646 792159
rect 42698 792107 42704 792159
rect 42832 792107 42838 792159
rect 42890 792107 42896 792159
rect 42544 791885 42550 791937
rect 42602 791925 42608 791937
rect 42658 791925 42686 792107
rect 42602 791897 42686 791925
rect 42602 791885 42608 791897
rect 42640 791811 42646 791863
rect 42698 791851 42704 791863
rect 42850 791851 42878 792107
rect 42698 791823 42878 791851
rect 42698 791811 42704 791823
rect 42064 791441 42070 791493
rect 42122 791481 42128 791493
rect 42544 791481 42550 791493
rect 42122 791453 42550 791481
rect 42122 791441 42128 791453
rect 42544 791441 42550 791453
rect 42602 791441 42608 791493
rect 42160 790775 42166 790827
rect 42218 790815 42224 790827
rect 42640 790815 42646 790827
rect 42218 790787 42646 790815
rect 42218 790775 42224 790787
rect 42640 790775 42646 790787
rect 42698 790775 42704 790827
rect 43312 789739 43318 789791
rect 43370 789779 43376 789791
rect 58000 789779 58006 789791
rect 43370 789751 58006 789779
rect 43370 789739 43376 789751
rect 58000 789739 58006 789751
rect 58058 789739 58064 789791
rect 42064 789591 42070 789643
rect 42122 789631 42128 789643
rect 43120 789631 43126 789643
rect 42122 789603 43126 789631
rect 42122 789591 42128 789603
rect 43120 789591 43126 789603
rect 43178 789591 43184 789643
rect 42640 789147 42646 789199
rect 42698 789187 42704 789199
rect 58192 789187 58198 789199
rect 42698 789159 58198 789187
rect 42698 789147 42704 789159
rect 58192 789147 58198 789159
rect 58250 789147 58256 789199
rect 44848 789073 44854 789125
rect 44906 789113 44912 789125
rect 58384 789113 58390 789125
rect 44906 789085 58390 789113
rect 44906 789073 44912 789085
rect 58384 789073 58390 789085
rect 58442 789073 58448 789125
rect 42256 787815 42262 787867
rect 42314 787855 42320 787867
rect 43024 787855 43030 787867
rect 42314 787827 43030 787855
rect 42314 787815 42320 787827
rect 43024 787815 43030 787827
rect 43082 787815 43088 787867
rect 42160 787223 42166 787275
rect 42218 787263 42224 787275
rect 42928 787263 42934 787275
rect 42218 787235 42934 787263
rect 42218 787223 42224 787235
rect 42928 787223 42934 787235
rect 42986 787223 42992 787275
rect 42160 785891 42166 785943
rect 42218 785931 42224 785943
rect 42640 785931 42646 785943
rect 42218 785903 42646 785931
rect 42218 785891 42224 785903
rect 42640 785891 42646 785903
rect 42698 785891 42704 785943
rect 44752 785595 44758 785647
rect 44810 785635 44816 785647
rect 58672 785635 58678 785647
rect 44810 785607 58678 785635
rect 44810 785595 44816 785607
rect 58672 785595 58678 785607
rect 58730 785595 58736 785647
rect 47536 785225 47542 785277
rect 47594 785265 47600 785277
rect 59632 785265 59638 785277
rect 47594 785237 59638 785265
rect 47594 785225 47600 785237
rect 59632 785225 59638 785237
rect 59690 785225 59696 785277
rect 675376 774831 675382 774843
rect 659506 774803 675382 774831
rect 654160 774717 654166 774769
rect 654218 774757 654224 774769
rect 659506 774757 659534 774803
rect 675376 774791 675382 774803
rect 675434 774791 675440 774843
rect 654218 774729 659534 774757
rect 654218 774717 654224 774729
rect 41776 774643 41782 774695
rect 41834 774683 41840 774695
rect 47632 774683 47638 774695
rect 41834 774655 47638 774683
rect 41834 774643 41840 774655
rect 47632 774643 47638 774655
rect 47690 774643 47696 774695
rect 41584 773903 41590 773955
rect 41642 773943 41648 773955
rect 44752 773943 44758 773955
rect 41642 773915 44758 773943
rect 41642 773903 41648 773915
rect 44752 773903 44758 773915
rect 44810 773903 44816 773955
rect 41776 773459 41782 773511
rect 41834 773499 41840 773511
rect 44944 773499 44950 773511
rect 41834 773471 44950 773499
rect 41834 773459 41840 773471
rect 44944 773459 44950 773471
rect 45002 773459 45008 773511
rect 41584 773385 41590 773437
rect 41642 773425 41648 773437
rect 43216 773425 43222 773437
rect 41642 773397 43222 773425
rect 41642 773385 41648 773397
rect 43216 773385 43222 773397
rect 43274 773385 43280 773437
rect 41776 772571 41782 772623
rect 41834 772611 41840 772623
rect 43216 772611 43222 772623
rect 41834 772583 43222 772611
rect 41834 772571 41840 772583
rect 43216 772571 43222 772583
rect 43274 772571 43280 772623
rect 41584 772127 41590 772179
rect 41642 772167 41648 772179
rect 62032 772167 62038 772179
rect 41642 772139 62038 772167
rect 41642 772127 41648 772139
rect 62032 772127 62038 772139
rect 62090 772127 62096 772179
rect 43120 771905 43126 771957
rect 43178 771945 43184 771957
rect 61840 771945 61846 771957
rect 43178 771917 61846 771945
rect 43178 771905 43184 771917
rect 61840 771905 61846 771917
rect 61898 771905 61904 771957
rect 654832 771905 654838 771957
rect 654890 771945 654896 771957
rect 674992 771945 674998 771957
rect 654890 771917 674998 771945
rect 654890 771905 654896 771917
rect 674992 771905 674998 771917
rect 675050 771905 675056 771957
rect 656176 771831 656182 771883
rect 656234 771871 656240 771883
rect 675088 771871 675094 771883
rect 656234 771843 675094 771871
rect 656234 771831 656240 771843
rect 675088 771831 675094 771843
rect 675146 771831 675152 771883
rect 674224 771313 674230 771365
rect 674282 771353 674288 771365
rect 675376 771353 675382 771365
rect 674282 771325 675382 771353
rect 674282 771313 674288 771325
rect 675376 771313 675382 771325
rect 675434 771313 675440 771365
rect 41776 769611 41782 769663
rect 41834 769651 41840 769663
rect 43120 769651 43126 769663
rect 41834 769623 43126 769651
rect 41834 769611 41840 769623
rect 43120 769611 43126 769623
rect 43178 769611 43184 769663
rect 674416 766799 674422 766851
rect 674474 766839 674480 766851
rect 675376 766839 675382 766851
rect 674474 766811 675382 766839
rect 674474 766799 674480 766811
rect 675376 766799 675382 766811
rect 675434 766799 675440 766851
rect 674128 766281 674134 766333
rect 674186 766321 674192 766333
rect 675472 766321 675478 766333
rect 674186 766293 675478 766321
rect 674186 766281 674192 766293
rect 675472 766281 675478 766293
rect 675530 766281 675536 766333
rect 674320 765689 674326 765741
rect 674378 765729 674384 765741
rect 675472 765729 675478 765741
rect 674378 765701 675478 765729
rect 674378 765689 674384 765701
rect 675472 765689 675478 765701
rect 675530 765689 675536 765741
rect 675088 765245 675094 765297
rect 675146 765285 675152 765297
rect 675376 765285 675382 765297
rect 675146 765257 675382 765285
rect 675146 765245 675152 765257
rect 675376 765245 675382 765257
rect 675434 765245 675440 765297
rect 41776 765097 41782 765149
rect 41834 765137 41840 765149
rect 42736 765137 42742 765149
rect 41834 765109 42742 765137
rect 41834 765097 41840 765109
rect 42736 765097 42742 765109
rect 42794 765097 42800 765149
rect 674512 765097 674518 765149
rect 674570 765137 674576 765149
rect 675472 765137 675478 765149
rect 674570 765109 675478 765137
rect 674570 765097 674576 765109
rect 675472 765097 675478 765109
rect 675530 765097 675536 765149
rect 674896 763691 674902 763743
rect 674954 763731 674960 763743
rect 675376 763731 675382 763743
rect 674954 763703 675382 763731
rect 674954 763691 674960 763703
rect 675376 763691 675382 763703
rect 675434 763691 675440 763743
rect 41584 763543 41590 763595
rect 41642 763583 41648 763595
rect 42928 763583 42934 763595
rect 41642 763555 42934 763583
rect 41642 763543 41648 763555
rect 42928 763543 42934 763555
rect 42986 763543 42992 763595
rect 674992 763469 674998 763521
rect 675050 763509 675056 763521
rect 675376 763509 675382 763521
rect 675050 763481 675382 763509
rect 675050 763469 675056 763481
rect 675376 763469 675382 763481
rect 675434 763469 675440 763521
rect 41584 763395 41590 763447
rect 41642 763435 41648 763447
rect 42832 763435 42838 763447
rect 41642 763407 42838 763435
rect 41642 763395 41648 763407
rect 42832 763395 42838 763407
rect 42890 763395 42896 763447
rect 41776 762063 41782 762115
rect 41834 762103 41840 762115
rect 47536 762103 47542 762115
rect 41834 762075 47542 762103
rect 41834 762063 41840 762075
rect 47536 762063 47542 762075
rect 47594 762063 47600 762115
rect 674992 761841 674998 761893
rect 675050 761881 675056 761893
rect 675376 761881 675382 761893
rect 675050 761853 675382 761881
rect 675050 761841 675056 761853
rect 675376 761841 675382 761853
rect 675434 761841 675440 761893
rect 40240 760287 40246 760339
rect 40298 760327 40304 760339
rect 41008 760327 41014 760339
rect 40298 760299 41014 760327
rect 40298 760287 40304 760299
rect 41008 760287 41014 760299
rect 41066 760287 41072 760339
rect 674896 760287 674902 760339
rect 674954 760327 674960 760339
rect 675376 760327 675382 760339
rect 674954 760299 675382 760327
rect 674954 760287 674960 760299
rect 675376 760287 675382 760299
rect 675434 760287 675440 760339
rect 37360 760213 37366 760265
rect 37418 760253 37424 760265
rect 41776 760253 41782 760265
rect 37418 760225 41782 760253
rect 37418 760213 37424 760225
rect 41776 760213 41782 760225
rect 41834 760213 41840 760265
rect 40144 758067 40150 758119
rect 40202 758107 40208 758119
rect 43600 758107 43606 758119
rect 40202 758079 43606 758107
rect 40202 758067 40208 758079
rect 43600 758067 43606 758079
rect 43658 758067 43664 758119
rect 42256 757919 42262 757971
rect 42314 757959 42320 757971
rect 43504 757959 43510 757971
rect 42314 757931 43510 757959
rect 42314 757919 42320 757931
rect 43504 757919 43510 757931
rect 43562 757919 43568 757971
rect 41968 757845 41974 757897
rect 42026 757885 42032 757897
rect 43408 757885 43414 757897
rect 42026 757857 43414 757885
rect 42026 757845 42032 757857
rect 43408 757845 43414 757857
rect 43466 757845 43472 757897
rect 41872 757771 41878 757823
rect 41930 757771 41936 757823
rect 42160 757771 42166 757823
rect 42218 757811 42224 757823
rect 43312 757811 43318 757823
rect 42218 757783 43318 757811
rect 42218 757771 42224 757783
rect 43312 757771 43318 757783
rect 43370 757771 43376 757823
rect 41890 757601 41918 757771
rect 41872 757549 41878 757601
rect 41930 757549 41936 757601
rect 42736 756365 42742 756417
rect 42794 756405 42800 756417
rect 42794 756377 42878 756405
rect 42794 756365 42800 756377
rect 42352 756143 42358 756195
rect 42410 756183 42416 756195
rect 42850 756183 42878 756377
rect 42410 756155 42878 756183
rect 42410 756143 42416 756155
rect 42160 755699 42166 755751
rect 42218 755739 42224 755751
rect 43120 755739 43126 755751
rect 42218 755711 43126 755739
rect 42218 755699 42224 755711
rect 43120 755699 43126 755711
rect 43178 755699 43184 755751
rect 43120 755551 43126 755603
rect 43178 755591 43184 755603
rect 43312 755591 43318 755603
rect 43178 755563 43318 755591
rect 43178 755551 43184 755563
rect 43312 755551 43318 755563
rect 43370 755551 43376 755603
rect 42064 754663 42070 754715
rect 42122 754703 42128 754715
rect 43312 754703 43318 754715
rect 42122 754675 43318 754703
rect 42122 754663 42128 754675
rect 43312 754663 43318 754675
rect 43370 754663 43376 754715
rect 42160 753849 42166 753901
rect 42218 753889 42224 753901
rect 42928 753889 42934 753901
rect 42218 753861 42934 753889
rect 42218 753849 42224 753861
rect 42928 753849 42934 753861
rect 42986 753849 42992 753901
rect 42928 753701 42934 753753
rect 42986 753741 42992 753753
rect 43408 753741 43414 753753
rect 42986 753713 43414 753741
rect 42986 753701 42992 753713
rect 43408 753701 43414 753713
rect 43466 753701 43472 753753
rect 42160 752591 42166 752643
rect 42218 752631 42224 752643
rect 42832 752631 42838 752643
rect 42218 752603 42838 752631
rect 42218 752591 42224 752603
rect 42832 752591 42838 752603
rect 42890 752591 42896 752643
rect 42064 752369 42070 752421
rect 42122 752409 42128 752421
rect 43408 752409 43414 752421
rect 42122 752381 43414 752409
rect 42122 752369 42128 752381
rect 43408 752369 43414 752381
rect 43466 752369 43472 752421
rect 42352 752039 42358 752051
rect 42274 752011 42358 752039
rect 42064 751851 42070 751903
rect 42122 751891 42128 751903
rect 42274 751891 42302 752011
rect 42352 751999 42358 752011
rect 42410 751999 42416 752051
rect 42122 751863 42302 751891
rect 42122 751851 42128 751863
rect 42352 751851 42358 751903
rect 42410 751891 42416 751903
rect 43120 751891 43126 751903
rect 42410 751863 43126 751891
rect 42410 751851 42416 751863
rect 43120 751851 43126 751863
rect 43178 751851 43184 751903
rect 43024 751777 43030 751829
rect 43082 751817 43088 751829
rect 43504 751817 43510 751829
rect 43082 751789 43510 751817
rect 43082 751777 43088 751789
rect 43504 751777 43510 751789
rect 43562 751777 43568 751829
rect 42832 751629 42838 751681
rect 42890 751669 42896 751681
rect 43120 751669 43126 751681
rect 42890 751641 43126 751669
rect 42890 751629 42896 751641
rect 43120 751629 43126 751641
rect 43178 751629 43184 751681
rect 42352 751555 42358 751607
rect 42410 751595 42416 751607
rect 42410 751567 42878 751595
rect 42410 751555 42416 751567
rect 42850 751533 42878 751567
rect 42832 751481 42838 751533
rect 42890 751481 42896 751533
rect 42160 751259 42166 751311
rect 42218 751299 42224 751311
rect 42928 751299 42934 751311
rect 42218 751271 42934 751299
rect 42218 751259 42224 751271
rect 42928 751259 42934 751271
rect 42986 751259 42992 751311
rect 42160 750519 42166 750571
rect 42218 750559 42224 750571
rect 43024 750559 43030 750571
rect 42218 750531 43030 750559
rect 42218 750519 42224 750531
rect 43024 750519 43030 750531
rect 43082 750519 43088 750571
rect 43312 748743 43318 748795
rect 43370 748783 43376 748795
rect 57904 748783 57910 748795
rect 43370 748755 57910 748783
rect 43370 748743 43376 748755
rect 57904 748743 57910 748755
rect 57962 748743 57968 748795
rect 42160 748151 42166 748203
rect 42218 748191 42224 748203
rect 42832 748191 42838 748203
rect 42218 748163 42838 748191
rect 42218 748151 42224 748163
rect 42832 748151 42838 748163
rect 42890 748151 42896 748203
rect 42160 747559 42166 747611
rect 42218 747599 42224 747611
rect 43600 747599 43606 747611
rect 42218 747571 43606 747599
rect 42218 747559 42224 747571
rect 43600 747559 43606 747571
rect 43658 747559 43664 747611
rect 42160 746227 42166 746279
rect 42218 746267 42224 746279
rect 42928 746267 42934 746279
rect 42218 746239 42934 746267
rect 42218 746227 42224 746239
rect 42928 746227 42934 746239
rect 42986 746227 42992 746279
rect 42352 746079 42358 746131
rect 42410 746119 42416 746131
rect 44848 746119 44854 746131
rect 42410 746091 44854 746119
rect 42410 746079 42416 746091
rect 44848 746079 44854 746091
rect 44906 746079 44912 746131
rect 42352 745931 42358 745983
rect 42410 745971 42416 745983
rect 54640 745971 54646 745983
rect 42410 745943 54646 745971
rect 42410 745931 42416 745943
rect 54640 745931 54646 745943
rect 54698 745931 54704 745983
rect 54736 745931 54742 745983
rect 54794 745971 54800 745983
rect 57616 745971 57622 745983
rect 54794 745943 57622 745971
rect 54794 745931 54800 745943
rect 57616 745931 57622 745943
rect 57674 745931 57680 745983
rect 44944 745339 44950 745391
rect 45002 745379 45008 745391
rect 59248 745379 59254 745391
rect 45002 745351 59254 745379
rect 45002 745339 45008 745351
rect 59248 745339 59254 745351
rect 59306 745339 59312 745391
rect 43408 745265 43414 745317
rect 43466 745305 43472 745317
rect 59632 745305 59638 745317
rect 43466 745277 59638 745305
rect 43466 745265 43472 745277
rect 59632 745265 59638 745277
rect 59690 745265 59696 745317
rect 42160 744599 42166 744651
rect 42218 744639 42224 744651
rect 43024 744639 43030 744651
rect 42218 744611 43030 744639
rect 42218 744599 42224 744611
rect 43024 744599 43030 744611
rect 43082 744599 43088 744651
rect 42160 744007 42166 744059
rect 42218 744047 42224 744059
rect 43120 744047 43126 744059
rect 42218 744019 43126 744047
rect 42218 744007 42224 744019
rect 43120 744007 43126 744019
rect 43178 744007 43184 744059
rect 42064 743341 42070 743393
rect 42122 743381 42128 743393
rect 42832 743381 42838 743393
rect 42122 743353 42838 743381
rect 42122 743341 42128 743353
rect 42832 743341 42838 743353
rect 42890 743341 42896 743393
rect 47632 742971 47638 743023
rect 47690 743011 47696 743023
rect 59632 743011 59638 743023
rect 47690 742983 59638 743011
rect 47690 742971 47696 742983
rect 59632 742971 59638 742983
rect 59690 742971 59696 743023
rect 44752 742897 44758 742949
rect 44810 742937 44816 742949
rect 59728 742937 59734 742949
rect 44810 742909 59734 742937
rect 44810 742897 44816 742909
rect 59728 742897 59734 742909
rect 59786 742897 59792 742949
rect 42160 742749 42166 742801
rect 42218 742789 42224 742801
rect 42352 742789 42358 742801
rect 42218 742761 42358 742789
rect 42218 742749 42224 742761
rect 42352 742749 42358 742761
rect 42410 742749 42416 742801
rect 41776 731427 41782 731479
rect 41834 731467 41840 731479
rect 50320 731467 50326 731479
rect 41834 731439 50326 731467
rect 41834 731427 41840 731439
rect 50320 731427 50326 731439
rect 50378 731427 50384 731479
rect 41584 730687 41590 730739
rect 41642 730727 41648 730739
rect 47728 730727 47734 730739
rect 41642 730699 47734 730727
rect 41642 730687 41648 730699
rect 47728 730687 47734 730699
rect 47786 730687 47792 730739
rect 41776 730317 41782 730369
rect 41834 730357 41840 730369
rect 44752 730357 44758 730369
rect 41834 730329 44758 730357
rect 41834 730317 41840 730329
rect 44752 730317 44758 730329
rect 44810 730317 44816 730369
rect 41584 730169 41590 730221
rect 41642 730209 41648 730221
rect 43216 730209 43222 730221
rect 41642 730181 43222 730209
rect 41642 730169 41648 730181
rect 43216 730169 43222 730181
rect 43274 730169 43280 730221
rect 41584 729207 41590 729259
rect 41642 729247 41648 729259
rect 43696 729247 43702 729259
rect 41642 729219 43702 729247
rect 41642 729207 41648 729219
rect 43696 729207 43702 729219
rect 43754 729207 43760 729259
rect 41200 728837 41206 728889
rect 41258 728877 41264 728889
rect 62224 728877 62230 728889
rect 41258 728849 62230 728877
rect 41258 728837 41264 728849
rect 62224 728837 62230 728849
rect 62282 728837 62288 728889
rect 40432 728763 40438 728815
rect 40490 728803 40496 728815
rect 62416 728803 62422 728815
rect 40490 728775 62422 728803
rect 40490 728763 40496 728775
rect 62416 728763 62422 728775
rect 62474 728763 62480 728815
rect 654160 728689 654166 728741
rect 654218 728729 654224 728741
rect 675280 728729 675286 728741
rect 654218 728701 675286 728729
rect 654218 728689 654224 728701
rect 675280 728689 675286 728701
rect 675338 728689 675344 728741
rect 41584 728615 41590 728667
rect 41642 728655 41648 728667
rect 43504 728655 43510 728667
rect 41642 728627 43510 728655
rect 41642 728615 41648 728627
rect 43504 728615 43510 728627
rect 43562 728615 43568 728667
rect 41776 727875 41782 727927
rect 41834 727915 41840 727927
rect 43408 727915 43414 727927
rect 41834 727887 43414 727915
rect 41834 727875 41840 727887
rect 43408 727875 43414 727887
rect 43466 727875 43472 727927
rect 654256 727135 654262 727187
rect 654314 727175 654320 727187
rect 674608 727175 674614 727187
rect 654314 727147 674614 727175
rect 654314 727135 654320 727147
rect 674608 727135 674614 727147
rect 674666 727135 674672 727187
rect 41776 726099 41782 726151
rect 41834 726139 41840 726151
rect 42928 726139 42934 726151
rect 41834 726111 42934 726139
rect 41834 726099 41840 726111
rect 42928 726099 42934 726111
rect 42986 726099 42992 726151
rect 673264 724915 673270 724967
rect 673322 724955 673328 724967
rect 675472 724955 675478 724967
rect 673322 724927 675478 724955
rect 673322 724915 673328 724927
rect 675472 724915 675478 724927
rect 675530 724915 675536 724967
rect 654160 724323 654166 724375
rect 654218 724363 654224 724375
rect 673936 724363 673942 724375
rect 654218 724335 673942 724363
rect 654218 724323 654224 724335
rect 673936 724323 673942 724335
rect 673994 724323 674000 724375
rect 673936 723361 673942 723413
rect 673994 723401 674000 723413
rect 675280 723401 675286 723413
rect 673994 723373 675286 723401
rect 673994 723361 674000 723373
rect 675280 723361 675286 723373
rect 675338 723361 675344 723413
rect 674512 722399 674518 722451
rect 674570 722439 674576 722451
rect 675376 722439 675382 722451
rect 674570 722411 675382 722439
rect 674570 722399 674576 722411
rect 675376 722399 675382 722411
rect 675434 722399 675440 722451
rect 41584 721363 41590 721415
rect 41642 721403 41648 721415
rect 43120 721403 43126 721415
rect 41642 721375 43126 721403
rect 41642 721363 41648 721375
rect 43120 721363 43126 721375
rect 43178 721363 43184 721415
rect 674032 721141 674038 721193
rect 674090 721181 674096 721193
rect 675472 721181 675478 721193
rect 674090 721153 675478 721181
rect 674090 721141 674096 721153
rect 675472 721141 675478 721153
rect 675530 721141 675536 721193
rect 674608 720845 674614 720897
rect 674666 720885 674672 720897
rect 675376 720885 675382 720897
rect 674666 720857 675382 720885
rect 674666 720845 674672 720857
rect 675376 720845 675382 720857
rect 675434 720845 675440 720897
rect 672880 720697 672886 720749
rect 672938 720737 672944 720749
rect 675472 720737 675478 720749
rect 672938 720709 675478 720737
rect 672938 720697 672944 720709
rect 675472 720697 675478 720709
rect 675530 720697 675536 720749
rect 41584 720401 41590 720453
rect 41642 720441 41648 720453
rect 42832 720441 42838 720453
rect 41642 720413 42838 720441
rect 41642 720401 41648 720413
rect 42832 720401 42838 720413
rect 42890 720401 42896 720453
rect 41584 720179 41590 720231
rect 41642 720219 41648 720231
rect 43024 720219 43030 720231
rect 41642 720191 43030 720219
rect 41642 720179 41648 720191
rect 43024 720179 43030 720191
rect 43082 720179 43088 720231
rect 674512 719291 674518 719343
rect 674570 719331 674576 719343
rect 675376 719331 675382 719343
rect 674570 719303 675382 719331
rect 674570 719291 674576 719303
rect 675376 719291 675382 719303
rect 675434 719291 675440 719343
rect 41584 718699 41590 718751
rect 41642 718739 41648 718751
rect 47632 718739 47638 718751
rect 41642 718711 47638 718739
rect 41642 718699 41648 718711
rect 47632 718699 47638 718711
rect 47690 718699 47696 718751
rect 675280 715591 675286 715643
rect 675338 715591 675344 715643
rect 675376 715591 675382 715643
rect 675434 715591 675440 715643
rect 675298 715335 675326 715591
rect 675394 715421 675422 715591
rect 675376 715369 675382 715421
rect 675434 715369 675440 715421
rect 675568 715335 675574 715347
rect 675298 715307 675574 715335
rect 675568 715295 675574 715307
rect 675626 715295 675632 715347
rect 41968 714629 41974 714681
rect 42026 714669 42032 714681
rect 43312 714669 43318 714681
rect 42026 714641 43318 714669
rect 42026 714629 42032 714641
rect 43312 714629 43318 714641
rect 43370 714629 43376 714681
rect 41776 714555 41782 714607
rect 41834 714555 41840 714607
rect 41872 714555 41878 714607
rect 41930 714595 41936 714607
rect 43600 714595 43606 714607
rect 41930 714567 43606 714595
rect 41930 714555 41936 714567
rect 43600 714555 43606 714567
rect 43658 714555 43664 714607
rect 41794 714385 41822 714555
rect 41776 714333 41782 714385
rect 41834 714333 41840 714385
rect 42256 714259 42262 714311
rect 42314 714299 42320 714311
rect 43216 714299 43222 714311
rect 42314 714271 43222 714299
rect 42314 714259 42320 714271
rect 43216 714259 43222 714271
rect 43274 714259 43280 714311
rect 673360 714185 673366 714237
rect 673418 714225 673424 714237
rect 679696 714225 679702 714237
rect 673418 714197 679702 714225
rect 673418 714185 673424 714197
rect 679696 714185 679702 714197
rect 679754 714185 679760 714237
rect 42832 712853 42838 712905
rect 42890 712893 42896 712905
rect 43120 712893 43126 712905
rect 42890 712865 43126 712893
rect 42890 712853 42896 712865
rect 43120 712853 43126 712865
rect 43178 712853 43184 712905
rect 43216 712557 43222 712609
rect 43274 712597 43280 712609
rect 43504 712597 43510 712609
rect 43274 712569 43510 712597
rect 43274 712557 43280 712569
rect 43504 712557 43510 712569
rect 43562 712557 43568 712609
rect 42064 712483 42070 712535
rect 42122 712523 42128 712535
rect 42928 712523 42934 712535
rect 42122 712495 42934 712523
rect 42122 712483 42128 712495
rect 42928 712483 42934 712495
rect 42986 712483 42992 712535
rect 42928 712335 42934 712387
rect 42986 712375 42992 712387
rect 43312 712375 43318 712387
rect 42986 712347 43318 712375
rect 42986 712335 42992 712347
rect 43312 712335 43318 712347
rect 43370 712335 43376 712387
rect 43312 712187 43318 712239
rect 43370 712227 43376 712239
rect 43696 712227 43702 712239
rect 43370 712199 43702 712227
rect 43370 712187 43376 712199
rect 43696 712187 43702 712199
rect 43754 712187 43760 712239
rect 42160 711225 42166 711277
rect 42218 711265 42224 711277
rect 43696 711265 43702 711277
rect 42218 711237 43702 711265
rect 42218 711225 42224 711237
rect 43696 711225 43702 711237
rect 43754 711225 43760 711277
rect 42064 710633 42070 710685
rect 42122 710673 42128 710685
rect 42832 710673 42838 710685
rect 42122 710645 42838 710673
rect 42122 710633 42128 710645
rect 42832 710633 42838 710645
rect 42890 710633 42896 710685
rect 42832 710485 42838 710537
rect 42890 710525 42896 710537
rect 43600 710525 43606 710537
rect 42890 710497 43606 710525
rect 42890 710485 42896 710497
rect 43600 710485 43606 710497
rect 43658 710485 43664 710537
rect 674032 709893 674038 709945
rect 674090 709933 674096 709945
rect 675664 709933 675670 709945
rect 674090 709905 675670 709933
rect 674090 709893 674096 709905
rect 675664 709893 675670 709905
rect 675722 709893 675728 709945
rect 42160 709597 42166 709649
rect 42218 709637 42224 709649
rect 43504 709637 43510 709649
rect 42218 709609 43510 709637
rect 42218 709597 42224 709609
rect 43504 709597 43510 709609
rect 43562 709597 43568 709649
rect 42064 709375 42070 709427
rect 42122 709415 42128 709427
rect 43024 709415 43030 709427
rect 42122 709387 43030 709415
rect 42122 709375 42128 709387
rect 43024 709375 43030 709387
rect 43082 709375 43088 709427
rect 43024 708783 43030 708835
rect 43082 708783 43088 708835
rect 42160 708635 42166 708687
rect 42218 708675 42224 708687
rect 42832 708675 42838 708687
rect 42218 708647 42838 708675
rect 42218 708635 42224 708647
rect 42832 708635 42838 708647
rect 42890 708635 42896 708687
rect 42160 708191 42166 708243
rect 42218 708231 42224 708243
rect 42736 708231 42742 708243
rect 42218 708203 42742 708231
rect 42218 708191 42224 708203
rect 42736 708191 42742 708203
rect 42794 708191 42800 708243
rect 42736 708043 42742 708095
rect 42794 708083 42800 708095
rect 43042 708083 43070 708783
rect 42794 708055 43070 708083
rect 42794 708043 42800 708055
rect 42064 707229 42070 707281
rect 42122 707269 42128 707281
rect 42928 707269 42934 707281
rect 42122 707241 42934 707269
rect 42122 707229 42128 707241
rect 42928 707229 42934 707241
rect 42986 707229 42992 707281
rect 42352 705527 42358 705579
rect 42410 705567 42416 705579
rect 42736 705567 42742 705579
rect 42410 705539 42742 705567
rect 42410 705527 42416 705539
rect 42736 705527 42742 705539
rect 42794 705527 42800 705579
rect 42160 705083 42166 705135
rect 42218 705123 42224 705135
rect 42352 705123 42358 705135
rect 42218 705095 42358 705123
rect 42218 705083 42224 705095
rect 42352 705083 42358 705095
rect 42410 705083 42416 705135
rect 43696 704861 43702 704913
rect 43754 704901 43760 704913
rect 58384 704901 58390 704913
rect 43754 704873 58390 704901
rect 43754 704861 43760 704873
rect 58384 704861 58390 704873
rect 58442 704861 58448 704913
rect 42160 704491 42166 704543
rect 42218 704531 42224 704543
rect 42832 704531 42838 704543
rect 42218 704503 42838 704531
rect 42218 704491 42224 704503
rect 42832 704491 42838 704503
rect 42890 704491 42896 704543
rect 42064 703751 42070 703803
rect 42122 703791 42128 703803
rect 43120 703791 43126 703803
rect 42122 703763 43126 703791
rect 42122 703751 42128 703763
rect 43120 703751 43126 703763
rect 43178 703751 43184 703803
rect 42160 703233 42166 703285
rect 42218 703273 42224 703285
rect 43024 703273 43030 703285
rect 42218 703245 43030 703273
rect 42218 703233 42224 703245
rect 43024 703233 43030 703245
rect 43082 703233 43088 703285
rect 655600 703011 655606 703063
rect 655658 703051 655664 703063
rect 676240 703051 676246 703063
rect 655658 703023 676246 703051
rect 655658 703011 655664 703023
rect 676240 703011 676246 703023
rect 676298 703011 676304 703063
rect 655216 702863 655222 702915
rect 655274 702903 655280 702915
rect 676240 702903 676246 702915
rect 655274 702875 676246 702903
rect 655274 702863 655280 702875
rect 676240 702863 676246 702875
rect 676298 702863 676304 702915
rect 43504 702641 43510 702693
rect 43562 702681 43568 702693
rect 58768 702681 58774 702693
rect 43562 702653 58774 702681
rect 43562 702641 43568 702653
rect 58768 702641 58774 702653
rect 58826 702641 58832 702693
rect 44752 702567 44758 702619
rect 44810 702607 44816 702619
rect 58672 702607 58678 702619
rect 44810 702579 58678 702607
rect 44810 702567 44816 702579
rect 58672 702567 58678 702579
rect 58730 702567 58736 702619
rect 42064 700791 42070 700843
rect 42122 700831 42128 700843
rect 42928 700831 42934 700843
rect 42122 700803 42934 700831
rect 42122 700791 42128 700803
rect 42928 700791 42934 700803
rect 42986 700791 42992 700843
rect 669520 700791 669526 700843
rect 669578 700831 669584 700843
rect 670864 700831 670870 700843
rect 669578 700803 670870 700831
rect 669578 700791 669584 700803
rect 670864 700791 670870 700803
rect 670922 700831 670928 700843
rect 676240 700831 676246 700843
rect 670922 700803 676246 700831
rect 670922 700791 670928 700803
rect 676240 700791 676246 700803
rect 676298 700791 676304 700843
rect 42160 700199 42166 700251
rect 42218 700239 42224 700251
rect 42736 700239 42742 700251
rect 42218 700211 42742 700239
rect 42218 700199 42224 700211
rect 42736 700199 42742 700211
rect 42794 700199 42800 700251
rect 670672 700051 670678 700103
rect 670730 700091 670736 700103
rect 676240 700091 676246 700103
rect 670730 700063 676246 700091
rect 670730 700051 670736 700063
rect 676240 700051 676246 700063
rect 676298 700051 676304 700103
rect 655408 699829 655414 699881
rect 655466 699869 655472 699881
rect 676048 699869 676054 699881
rect 655466 699841 676054 699869
rect 655466 699829 655472 699841
rect 676048 699829 676054 699841
rect 676106 699829 676112 699881
rect 50320 699755 50326 699807
rect 50378 699795 50384 699807
rect 59248 699795 59254 699807
rect 50378 699767 59254 699795
rect 50378 699755 50384 699767
rect 59248 699755 59254 699767
rect 59306 699755 59312 699807
rect 47728 699681 47734 699733
rect 47786 699721 47792 699733
rect 58864 699721 58870 699733
rect 47786 699693 58870 699721
rect 47786 699681 47792 699693
rect 58864 699681 58870 699693
rect 58922 699681 58928 699733
rect 670960 699681 670966 699733
rect 671018 699721 671024 699733
rect 676048 699721 676054 699733
rect 671018 699693 676054 699721
rect 671018 699681 671024 699693
rect 676048 699681 676054 699693
rect 676106 699681 676112 699733
rect 42064 699533 42070 699585
rect 42122 699573 42128 699585
rect 42832 699573 42838 699585
rect 42122 699545 42838 699573
rect 42122 699533 42128 699545
rect 42832 699533 42838 699545
rect 42890 699533 42896 699585
rect 674224 699163 674230 699215
rect 674282 699203 674288 699215
rect 676240 699203 676246 699215
rect 674282 699175 676246 699203
rect 674282 699163 674288 699175
rect 676240 699163 676246 699175
rect 676298 699163 676304 699215
rect 670864 699089 670870 699141
rect 670922 699129 670928 699141
rect 676048 699129 676054 699141
rect 670922 699101 676054 699129
rect 670922 699089 670928 699101
rect 676048 699089 676054 699101
rect 676106 699089 676112 699141
rect 674992 698941 674998 698993
rect 675050 698981 675056 698993
rect 676048 698981 676054 698993
rect 675050 698953 676054 698981
rect 675050 698941 675056 698953
rect 676048 698941 676054 698953
rect 676106 698941 676112 698993
rect 669712 696943 669718 696995
rect 669770 696983 669776 696995
rect 670960 696983 670966 696995
rect 669770 696955 670966 696983
rect 669770 696943 669776 696955
rect 670960 696943 670966 696955
rect 671018 696943 671024 696995
rect 674896 696869 674902 696921
rect 674954 696909 674960 696921
rect 676048 696909 676054 696921
rect 674954 696881 676054 696909
rect 674954 696869 674960 696881
rect 676048 696869 676054 696881
rect 676106 696869 676112 696921
rect 674416 696795 674422 696847
rect 674474 696835 674480 696847
rect 675952 696835 675958 696847
rect 674474 696807 675958 696835
rect 674474 696795 674480 696807
rect 675952 696795 675958 696807
rect 676010 696795 676016 696847
rect 674896 696647 674902 696699
rect 674954 696687 674960 696699
rect 676240 696687 676246 696699
rect 674954 696659 676246 696687
rect 674954 696647 674960 696659
rect 676240 696647 676246 696659
rect 676298 696647 676304 696699
rect 674320 693983 674326 694035
rect 674378 694023 674384 694035
rect 676048 694023 676054 694035
rect 674378 693995 676054 694023
rect 674378 693983 674384 693995
rect 676048 693983 676054 693995
rect 676106 693983 676112 694035
rect 674128 693613 674134 693665
rect 674186 693653 674192 693665
rect 676048 693653 676054 693665
rect 674186 693625 676054 693653
rect 674186 693613 674192 693625
rect 676048 693613 676054 693625
rect 676106 693613 676112 693665
rect 670768 691171 670774 691223
rect 670826 691211 670832 691223
rect 679696 691211 679702 691223
rect 670826 691183 679702 691211
rect 670826 691171 670832 691183
rect 679696 691171 679702 691183
rect 679754 691171 679760 691223
rect 674320 689765 674326 689817
rect 674378 689805 674384 689817
rect 675664 689805 675670 689817
rect 674378 689777 675670 689805
rect 674378 689765 674384 689777
rect 675664 689765 675670 689777
rect 675722 689765 675728 689817
rect 674992 689395 674998 689447
rect 675050 689435 675056 689447
rect 675568 689435 675574 689447
rect 675050 689407 675574 689435
rect 675050 689395 675056 689407
rect 675568 689395 675574 689407
rect 675626 689395 675632 689447
rect 649456 688359 649462 688411
rect 649514 688399 649520 688411
rect 679984 688399 679990 688411
rect 649514 688371 679990 688399
rect 649514 688359 649520 688371
rect 679984 688359 679990 688371
rect 680042 688359 680048 688411
rect 41776 688211 41782 688263
rect 41834 688251 41840 688263
rect 53200 688251 53206 688263
rect 41834 688223 53206 688251
rect 41834 688211 41840 688223
rect 53200 688211 53206 688223
rect 53258 688211 53264 688263
rect 41584 687471 41590 687523
rect 41642 687511 41648 687523
rect 50320 687511 50326 687523
rect 41642 687483 50326 687511
rect 41642 687471 41648 687483
rect 50320 687471 50326 687483
rect 50378 687471 50384 687523
rect 41776 687175 41782 687227
rect 41834 687215 41840 687227
rect 47824 687215 47830 687227
rect 41834 687187 47830 687215
rect 41834 687175 41840 687187
rect 47824 687175 47830 687187
rect 47882 687175 47888 687227
rect 41584 686953 41590 687005
rect 41642 686993 41648 687005
rect 43312 686993 43318 687005
rect 41642 686965 43318 686993
rect 41642 686953 41648 686965
rect 43312 686953 43318 686965
rect 43370 686953 43376 687005
rect 674032 686213 674038 686265
rect 674090 686253 674096 686265
rect 675376 686253 675382 686265
rect 674090 686225 675382 686253
rect 674090 686213 674096 686225
rect 675376 686213 675382 686225
rect 675434 686213 675440 686265
rect 41584 685991 41590 686043
rect 41642 686031 41648 686043
rect 43504 686031 43510 686043
rect 41642 686003 43510 686031
rect 41642 685991 41648 686003
rect 43504 685991 43510 686003
rect 43562 685991 43568 686043
rect 656368 685547 656374 685599
rect 656426 685587 656432 685599
rect 674032 685587 674038 685599
rect 656426 685559 674038 685587
rect 656426 685547 656432 685559
rect 674032 685547 674038 685559
rect 674090 685547 674096 685599
rect 41776 685325 41782 685377
rect 41834 685365 41840 685377
rect 43216 685365 43222 685377
rect 41834 685337 43222 685365
rect 41834 685325 41840 685337
rect 43216 685325 43222 685337
rect 43274 685365 43280 685377
rect 44752 685365 44758 685377
rect 43274 685337 44758 685365
rect 43274 685325 43280 685337
rect 44752 685325 44758 685337
rect 44810 685325 44816 685377
rect 672400 685325 672406 685377
rect 672458 685365 672464 685377
rect 675472 685365 675478 685377
rect 672458 685337 675478 685365
rect 672458 685325 672464 685337
rect 675472 685325 675478 685337
rect 675530 685325 675536 685377
rect 41584 684511 41590 684563
rect 41642 684551 41648 684563
rect 43312 684551 43318 684563
rect 41642 684523 43318 684551
rect 41642 684511 41648 684523
rect 43312 684511 43318 684523
rect 43370 684511 43376 684563
rect 41776 684141 41782 684193
rect 41834 684181 41840 684193
rect 43408 684181 43414 684193
rect 41834 684153 43414 684181
rect 41834 684141 41840 684153
rect 43408 684141 43414 684153
rect 43466 684181 43472 684193
rect 44944 684181 44950 684193
rect 43466 684153 44950 684181
rect 43466 684141 43472 684153
rect 44944 684141 44950 684153
rect 45002 684141 45008 684193
rect 41776 682735 41782 682787
rect 41834 682775 41840 682787
rect 43120 682775 43126 682787
rect 41834 682747 43126 682775
rect 41834 682735 41840 682747
rect 43120 682735 43126 682747
rect 43178 682735 43184 682787
rect 672688 682069 672694 682121
rect 672746 682109 672752 682121
rect 675472 682109 675478 682121
rect 672746 682081 675478 682109
rect 672746 682069 672752 682081
rect 675472 682069 675478 682081
rect 675530 682069 675536 682121
rect 672976 681255 672982 681307
rect 673034 681295 673040 681307
rect 675376 681295 675382 681307
rect 673034 681267 675382 681295
rect 673034 681255 673040 681267
rect 675376 681255 675382 681267
rect 675434 681255 675440 681307
rect 655984 681181 655990 681233
rect 656042 681221 656048 681233
rect 674896 681221 674902 681233
rect 656042 681193 674902 681221
rect 656042 681181 656048 681193
rect 674896 681181 674902 681193
rect 674954 681181 674960 681233
rect 654448 681107 654454 681159
rect 654506 681147 654512 681159
rect 674416 681147 674422 681159
rect 654506 681119 674422 681147
rect 654506 681107 654512 681119
rect 674416 681107 674422 681119
rect 674474 681107 674480 681159
rect 672208 680737 672214 680789
rect 672266 680777 672272 680789
rect 675376 680777 675382 680789
rect 672266 680749 675382 680777
rect 672266 680737 672272 680749
rect 675376 680737 675382 680749
rect 675434 680737 675440 680789
rect 674896 679627 674902 679679
rect 674954 679667 674960 679679
rect 675280 679667 675286 679679
rect 674954 679639 675286 679667
rect 674954 679627 674960 679639
rect 675280 679627 675286 679639
rect 675338 679627 675344 679679
rect 675184 679075 675190 679087
rect 675010 679047 675190 679075
rect 675010 678865 675038 679047
rect 675184 679035 675190 679047
rect 675242 679035 675248 679087
rect 674992 678813 674998 678865
rect 675050 678813 675056 678865
rect 673072 677555 673078 677607
rect 673130 677595 673136 677607
rect 675376 677595 675382 677607
rect 673130 677567 675382 677595
rect 673130 677555 673136 677567
rect 675376 677555 675382 677567
rect 675434 677555 675440 677607
rect 41584 677259 41590 677311
rect 41642 677299 41648 677311
rect 42928 677299 42934 677311
rect 41642 677271 42934 677299
rect 41642 677259 41648 677271
rect 42928 677259 42934 677271
rect 42986 677259 42992 677311
rect 41776 677185 41782 677237
rect 41834 677225 41840 677237
rect 42832 677225 42838 677237
rect 41834 677197 42838 677225
rect 41834 677185 41840 677197
rect 42832 677185 42838 677197
rect 42890 677185 42896 677237
rect 672496 677037 672502 677089
rect 672554 677077 672560 677089
rect 675472 677077 675478 677089
rect 672554 677049 675478 677077
rect 672554 677037 672560 677049
rect 675472 677037 675478 677049
rect 675530 677037 675536 677089
rect 673168 676667 673174 676719
rect 673226 676707 673232 676719
rect 675472 676707 675478 676719
rect 673226 676679 675478 676707
rect 673226 676667 673232 676679
rect 675472 676667 675478 676679
rect 675530 676667 675536 676719
rect 674416 676149 674422 676201
rect 674474 676189 674480 676201
rect 675280 676189 675286 676201
rect 674474 676161 675286 676189
rect 674474 676149 674480 676161
rect 675280 676149 675286 676161
rect 675338 676149 675344 676201
rect 41776 675705 41782 675757
rect 41834 675745 41840 675757
rect 47728 675745 47734 675757
rect 41834 675717 47734 675745
rect 41834 675705 41840 675717
rect 47728 675705 47734 675717
rect 47786 675705 47792 675757
rect 672304 675113 672310 675165
rect 672362 675153 672368 675165
rect 675472 675153 675478 675165
rect 672362 675125 675478 675153
rect 672362 675113 672368 675125
rect 675472 675113 675478 675125
rect 675530 675113 675536 675165
rect 42736 671043 42742 671095
rect 42794 671083 42800 671095
rect 59632 671083 59638 671095
rect 42794 671055 59638 671083
rect 42794 671043 42800 671055
rect 59632 671043 59638 671055
rect 59690 671043 59696 671095
rect 42256 670787 42262 670799
rect 42178 670759 42262 670787
rect 42178 670577 42206 670759
rect 42256 670747 42262 670759
rect 42314 670747 42320 670799
rect 42160 670525 42166 670577
rect 42218 670525 42224 670577
rect 674896 669637 674902 669689
rect 674954 669677 674960 669689
rect 675568 669677 675574 669689
rect 674954 669649 675574 669677
rect 674954 669637 674960 669649
rect 675568 669637 675574 669649
rect 675626 669637 675632 669689
rect 674992 669563 674998 669615
rect 675050 669603 675056 669615
rect 675472 669603 675478 669615
rect 675050 669575 675478 669603
rect 675050 669563 675056 669575
rect 675472 669563 675478 669575
rect 675530 669563 675536 669615
rect 42160 669119 42166 669171
rect 42218 669159 42224 669171
rect 43120 669159 43126 669171
rect 42218 669131 43126 669159
rect 42218 669119 42224 669131
rect 43120 669119 43126 669131
rect 43178 669119 43184 669171
rect 42832 668527 42838 668579
rect 42890 668567 42896 668579
rect 43120 668567 43126 668579
rect 42890 668539 43126 668567
rect 42890 668527 42896 668539
rect 43120 668527 43126 668539
rect 43178 668527 43184 668579
rect 42160 668453 42166 668505
rect 42218 668493 42224 668505
rect 42736 668493 42742 668505
rect 42218 668465 42742 668493
rect 42218 668453 42224 668465
rect 42736 668453 42742 668465
rect 42794 668453 42800 668505
rect 42160 667269 42166 667321
rect 42218 667309 42224 667321
rect 43024 667309 43030 667321
rect 42218 667281 43030 667309
rect 42218 667269 42224 667281
rect 43024 667269 43030 667281
rect 43082 667269 43088 667321
rect 42064 665863 42070 665915
rect 42122 665903 42128 665915
rect 43120 665903 43126 665915
rect 42122 665875 43126 665903
rect 42122 665863 42128 665875
rect 43120 665863 43126 665875
rect 43178 665863 43184 665915
rect 42160 665641 42166 665693
rect 42218 665681 42224 665693
rect 43216 665681 43222 665693
rect 42218 665653 43222 665681
rect 42218 665641 42224 665653
rect 43216 665641 43222 665653
rect 43274 665641 43280 665693
rect 42160 665419 42166 665471
rect 42218 665459 42224 665471
rect 42736 665459 42742 665471
rect 42218 665431 42742 665459
rect 42218 665419 42224 665431
rect 42736 665419 42742 665431
rect 42794 665419 42800 665471
rect 42064 664605 42070 664657
rect 42122 664645 42128 664657
rect 42928 664645 42934 664657
rect 42122 664617 42934 664645
rect 42122 664605 42128 664617
rect 42928 664605 42934 664617
rect 42986 664605 42992 664657
rect 42160 664161 42166 664213
rect 42218 664201 42224 664213
rect 42832 664201 42838 664213
rect 42218 664173 42838 664201
rect 42218 664161 42224 664173
rect 42832 664161 42838 664173
rect 42890 664161 42896 664213
rect 42064 661645 42070 661697
rect 42122 661685 42128 661697
rect 43024 661685 43030 661697
rect 42122 661657 43030 661685
rect 42122 661645 42128 661657
rect 43024 661645 43030 661657
rect 43082 661645 43088 661697
rect 42160 661127 42166 661179
rect 42218 661167 42224 661179
rect 42736 661167 42742 661179
rect 42218 661139 42742 661167
rect 42218 661127 42224 661139
rect 42736 661127 42742 661139
rect 42794 661127 42800 661179
rect 42160 660239 42166 660291
rect 42218 660279 42224 660291
rect 43120 660279 43126 660291
rect 42218 660251 43126 660279
rect 42218 660239 42224 660251
rect 43120 660239 43126 660251
rect 43178 660239 43184 660291
rect 42064 659647 42070 659699
rect 42122 659687 42128 659699
rect 42352 659687 42358 659699
rect 42122 659659 42358 659687
rect 42122 659647 42128 659659
rect 42352 659647 42358 659659
rect 42410 659647 42416 659699
rect 47824 659425 47830 659477
rect 47882 659465 47888 659477
rect 59152 659465 59158 659477
rect 47882 659437 59158 659465
rect 47882 659425 47888 659437
rect 59152 659425 59158 659437
rect 59210 659425 59216 659477
rect 43216 659351 43222 659403
rect 43274 659391 43280 659403
rect 58768 659391 58774 659403
rect 43274 659363 58774 659391
rect 43274 659351 43280 659363
rect 58768 659351 58774 659363
rect 58826 659351 58832 659403
rect 42160 657945 42166 657997
rect 42218 657985 42224 657997
rect 42928 657985 42934 657997
rect 42218 657957 42934 657985
rect 42218 657945 42224 657957
rect 42928 657945 42934 657957
rect 42986 657945 42992 657997
rect 670768 657575 670774 657627
rect 670826 657615 670832 657627
rect 676048 657615 676054 657627
rect 670826 657587 676054 657615
rect 670826 657575 670832 657587
rect 676048 657575 676054 657587
rect 676106 657575 676112 657627
rect 42160 657427 42166 657479
rect 42218 657467 42224 657479
rect 42832 657467 42838 657479
rect 42218 657439 42838 657467
rect 42218 657427 42224 657439
rect 42832 657427 42838 657439
rect 42890 657427 42896 657479
rect 655504 657131 655510 657183
rect 655562 657171 655568 657183
rect 676144 657171 676150 657183
rect 655562 657143 676150 657171
rect 655562 657131 655568 657143
rect 676144 657131 676150 657143
rect 676202 657131 676208 657183
rect 655312 656983 655318 657035
rect 655370 657023 655376 657035
rect 676240 657023 676246 657035
rect 655370 656995 676246 657023
rect 655370 656983 655376 656995
rect 676240 656983 676246 656995
rect 676298 656983 676304 657035
rect 673744 656909 673750 656961
rect 673802 656949 673808 656961
rect 676048 656949 676054 656961
rect 673802 656921 676054 656949
rect 673802 656909 673808 656921
rect 676048 656909 676054 656921
rect 676106 656909 676112 656961
rect 655120 656835 655126 656887
rect 655178 656875 655184 656887
rect 676336 656875 676342 656887
rect 655178 656847 676342 656875
rect 655178 656835 655184 656847
rect 676336 656835 676342 656847
rect 676394 656835 676400 656887
rect 42160 656761 42166 656813
rect 42218 656801 42224 656813
rect 43024 656801 43030 656813
rect 42218 656773 43030 656801
rect 42218 656761 42224 656773
rect 43024 656761 43030 656773
rect 43082 656761 43088 656813
rect 53200 656613 53206 656665
rect 53258 656653 53264 656665
rect 58192 656653 58198 656665
rect 53258 656625 58198 656653
rect 53258 656613 53264 656625
rect 58192 656613 58198 656625
rect 58250 656613 58256 656665
rect 50320 656539 50326 656591
rect 50378 656579 50384 656591
rect 58384 656579 58390 656591
rect 50378 656551 58390 656579
rect 50378 656539 50384 656551
rect 58384 656539 58390 656551
rect 58442 656539 58448 656591
rect 670672 656465 670678 656517
rect 670730 656505 670736 656517
rect 676048 656505 676054 656517
rect 670730 656477 676054 656505
rect 670730 656465 670736 656477
rect 676048 656465 676054 656477
rect 676106 656465 676112 656517
rect 42160 656095 42166 656147
rect 42218 656135 42224 656147
rect 45040 656135 45046 656147
rect 42218 656107 45046 656135
rect 42218 656095 42224 656107
rect 45040 656095 45046 656107
rect 45098 656095 45104 656147
rect 670864 656021 670870 656073
rect 670922 656061 670928 656073
rect 676048 656061 676054 656073
rect 670922 656033 676054 656061
rect 670922 656021 670928 656033
rect 676048 656021 676054 656033
rect 676106 656021 676112 656073
rect 670960 655725 670966 655777
rect 671018 655765 671024 655777
rect 676240 655765 676246 655777
rect 671018 655737 676246 655765
rect 671018 655725 671024 655737
rect 676240 655725 676246 655737
rect 676298 655725 676304 655777
rect 652240 655281 652246 655333
rect 652298 655321 652304 655333
rect 670960 655321 670966 655333
rect 652298 655293 670966 655321
rect 652298 655281 652304 655293
rect 670960 655281 670966 655293
rect 671018 655281 671024 655333
rect 649744 655207 649750 655259
rect 649802 655247 649808 655259
rect 670672 655247 670678 655259
rect 649802 655219 670678 655247
rect 649802 655207 649808 655219
rect 670672 655207 670678 655219
rect 670730 655207 670736 655259
rect 670768 654763 670774 654815
rect 670826 654803 670832 654815
rect 676240 654803 676246 654815
rect 670826 654775 676246 654803
rect 670826 654763 670832 654775
rect 676240 654763 676246 654775
rect 676298 654763 676304 654815
rect 674608 653727 674614 653779
rect 674666 653767 674672 653779
rect 676048 653767 676054 653779
rect 674666 653739 676054 653767
rect 674666 653727 674672 653739
rect 676048 653727 676054 653739
rect 676106 653727 676112 653779
rect 674512 650841 674518 650893
rect 674570 650881 674576 650893
rect 676048 650881 676054 650893
rect 674570 650853 676054 650881
rect 674570 650841 674576 650853
rect 676048 650841 676054 650853
rect 676106 650841 676112 650893
rect 673264 649213 673270 649265
rect 673322 649253 673328 649265
rect 676240 649253 676246 649265
rect 673322 649225 676246 649253
rect 673322 649213 673328 649225
rect 676240 649213 676246 649225
rect 676298 649213 676304 649265
rect 672880 648029 672886 648081
rect 672938 648069 672944 648081
rect 676048 648069 676054 648081
rect 672938 648041 676054 648069
rect 672938 648029 672944 648041
rect 676048 648029 676054 648041
rect 676106 648029 676112 648081
rect 649552 645143 649558 645195
rect 649610 645183 649616 645195
rect 679792 645183 679798 645195
rect 649610 645155 679798 645183
rect 649610 645143 649616 645155
rect 679792 645143 679798 645155
rect 679850 645143 679856 645195
rect 41584 644847 41590 644899
rect 41642 644887 41648 644899
rect 53200 644887 53206 644899
rect 41642 644859 53206 644887
rect 41642 644847 41648 644859
rect 53200 644847 53206 644859
rect 53258 644847 53264 644899
rect 41584 644255 41590 644307
rect 41642 644295 41648 644307
rect 50320 644295 50326 644307
rect 41642 644267 50326 644295
rect 41642 644255 41648 644267
rect 50320 644255 50326 644267
rect 50378 644255 50384 644307
rect 41776 643959 41782 644011
rect 41834 643999 41840 644011
rect 47920 643999 47926 644011
rect 41834 643971 47926 643999
rect 41834 643959 41840 643971
rect 47920 643959 47926 643971
rect 47978 643959 47984 644011
rect 41584 643737 41590 643789
rect 41642 643777 41648 643789
rect 43504 643777 43510 643789
rect 41642 643749 43510 643777
rect 41642 643737 41648 643749
rect 43504 643737 43510 643749
rect 43562 643737 43568 643789
rect 41584 642775 41590 642827
rect 41642 642815 41648 642827
rect 43216 642815 43222 642827
rect 41642 642787 43222 642815
rect 41642 642775 41648 642787
rect 43216 642775 43222 642787
rect 43274 642775 43280 642827
rect 43120 642479 43126 642531
rect 43178 642519 43184 642531
rect 61936 642519 61942 642531
rect 43178 642491 61942 642519
rect 43178 642479 43184 642491
rect 61936 642479 61942 642491
rect 61994 642479 62000 642531
rect 43408 642257 43414 642309
rect 43466 642297 43472 642309
rect 45136 642297 45142 642309
rect 43466 642269 45142 642297
rect 43466 642257 43472 642269
rect 45136 642257 45142 642269
rect 45194 642257 45200 642309
rect 654160 642183 654166 642235
rect 654218 642223 654224 642235
rect 675184 642223 675190 642235
rect 654218 642195 675190 642223
rect 654218 642183 654224 642195
rect 675184 642183 675190 642195
rect 675242 642183 675248 642235
rect 41584 641295 41590 641347
rect 41642 641335 41648 641347
rect 43312 641335 43318 641347
rect 41642 641307 43318 641335
rect 41642 641295 41648 641307
rect 43312 641295 43318 641307
rect 43370 641295 43376 641347
rect 41584 639667 41590 639719
rect 41642 639707 41648 639719
rect 43024 639707 43030 639719
rect 41642 639679 43030 639707
rect 41642 639667 41648 639679
rect 43024 639667 43030 639679
rect 43082 639667 43088 639719
rect 670960 637817 670966 637869
rect 671018 637857 671024 637869
rect 675376 637857 675382 637869
rect 671018 637829 675382 637857
rect 671018 637817 671024 637829
rect 675376 637817 675382 637829
rect 675434 637817 675440 637869
rect 673360 637077 673366 637129
rect 673418 637117 673424 637129
rect 675472 637117 675478 637129
rect 673418 637089 675478 637117
rect 673418 637077 673424 637089
rect 675472 637077 675478 637089
rect 675530 637077 675536 637129
rect 655792 636633 655798 636685
rect 655850 636673 655856 636685
rect 675184 636673 675190 636685
rect 655850 636645 675190 636673
rect 655850 636633 655856 636645
rect 675184 636633 675190 636645
rect 675242 636633 675248 636685
rect 673264 636485 673270 636537
rect 673322 636525 673328 636537
rect 675376 636525 675382 636537
rect 673322 636497 675382 636525
rect 673322 636485 673328 636497
rect 675376 636485 675382 636497
rect 675434 636485 675440 636537
rect 655888 635005 655894 635057
rect 655946 635045 655952 635057
rect 674992 635045 674998 635057
rect 655946 635017 674998 635045
rect 655946 635005 655952 635017
rect 674992 635005 674998 635017
rect 675050 635005 675056 635057
rect 41776 634191 41782 634243
rect 41834 634231 41840 634243
rect 43120 634231 43126 634243
rect 41834 634203 43126 634231
rect 41834 634191 41840 634203
rect 43120 634191 43126 634203
rect 43178 634191 43184 634243
rect 41776 633895 41782 633947
rect 41834 633935 41840 633947
rect 42928 633935 42934 633947
rect 41834 633907 42934 633935
rect 41834 633895 41840 633907
rect 42928 633895 42934 633907
rect 42986 633895 42992 633947
rect 672784 633599 672790 633651
rect 672842 633639 672848 633651
rect 675376 633639 675382 633651
rect 672842 633611 675382 633639
rect 672842 633599 672848 633611
rect 675376 633599 675382 633611
rect 675434 633599 675440 633651
rect 41776 632489 41782 632541
rect 41834 632529 41840 632541
rect 47824 632529 47830 632541
rect 41834 632501 47830 632529
rect 41834 632489 41840 632501
rect 47824 632489 47830 632501
rect 47882 632489 47888 632541
rect 672880 632341 672886 632393
rect 672938 632381 672944 632393
rect 675472 632381 675478 632393
rect 672938 632353 675478 632381
rect 672938 632341 672944 632353
rect 675472 632341 675478 632353
rect 675530 632341 675536 632393
rect 672592 630713 672598 630765
rect 672650 630753 672656 630765
rect 675280 630753 675286 630765
rect 672650 630725 675286 630753
rect 672650 630713 672656 630725
rect 675280 630713 675286 630725
rect 675338 630713 675344 630765
rect 674992 630639 674998 630691
rect 675050 630679 675056 630691
rect 675472 630679 675478 630691
rect 675050 630651 675478 630679
rect 675050 630639 675056 630651
rect 675472 630639 675478 630651
rect 675530 630639 675536 630691
rect 41872 627975 41878 628027
rect 41930 627975 41936 628027
rect 41890 627805 41918 627975
rect 42832 627827 42838 627879
rect 42890 627867 42896 627879
rect 54640 627867 54646 627879
rect 42890 627839 54646 627867
rect 42890 627827 42896 627839
rect 54640 627827 54646 627839
rect 54698 627827 54704 627879
rect 41872 627753 41878 627805
rect 41930 627753 41936 627805
rect 43120 626643 43126 626695
rect 43178 626683 43184 626695
rect 43178 626655 43262 626683
rect 43178 626643 43184 626655
rect 42928 626495 42934 626547
rect 42986 626535 42992 626547
rect 43120 626535 43126 626547
rect 42986 626507 43126 626535
rect 42986 626495 42992 626507
rect 43120 626495 43126 626507
rect 43178 626495 43184 626547
rect 42160 625903 42166 625955
rect 42218 625943 42224 625955
rect 43024 625943 43030 625955
rect 42218 625915 43030 625943
rect 42218 625903 42224 625915
rect 43024 625903 43030 625915
rect 43082 625903 43088 625955
rect 43024 625755 43030 625807
rect 43082 625795 43088 625807
rect 43234 625795 43262 626655
rect 43082 625767 43262 625795
rect 43082 625755 43088 625767
rect 42064 625237 42070 625289
rect 42122 625277 42128 625289
rect 42832 625277 42838 625289
rect 42122 625249 42838 625277
rect 42122 625237 42128 625249
rect 42832 625237 42838 625249
rect 42890 625237 42896 625289
rect 54640 624793 54646 624845
rect 54698 624833 54704 624845
rect 58960 624833 58966 624845
rect 54698 624805 58966 624833
rect 54698 624793 54704 624805
rect 58960 624793 58966 624805
rect 59018 624793 59024 624845
rect 42160 624053 42166 624105
rect 42218 624093 42224 624105
rect 43024 624093 43030 624105
rect 42218 624065 43030 624093
rect 42218 624053 42224 624065
rect 43024 624053 43030 624065
rect 43082 624053 43088 624105
rect 42064 622647 42070 622699
rect 42122 622687 42128 622699
rect 43120 622687 43126 622699
rect 42122 622659 43126 622687
rect 42122 622647 42128 622659
rect 43120 622647 43126 622659
rect 43178 622647 43184 622699
rect 42160 622499 42166 622551
rect 42218 622539 42224 622551
rect 43408 622539 43414 622551
rect 42218 622511 43414 622539
rect 42218 622499 42224 622511
rect 43408 622499 43414 622511
rect 43466 622499 43472 622551
rect 42064 622203 42070 622255
rect 42122 622243 42128 622255
rect 42832 622243 42838 622255
rect 42122 622215 42838 622243
rect 42122 622203 42128 622215
rect 42832 622203 42838 622215
rect 42890 622203 42896 622255
rect 42160 621463 42166 621515
rect 42218 621503 42224 621515
rect 42928 621503 42934 621515
rect 42218 621475 42934 621503
rect 42218 621463 42224 621475
rect 42928 621463 42934 621475
rect 42986 621463 42992 621515
rect 42160 618429 42166 618481
rect 42218 618469 42224 618481
rect 42832 618469 42838 618481
rect 42218 618441 42838 618469
rect 42218 618429 42224 618441
rect 42832 618429 42838 618441
rect 42890 618429 42896 618481
rect 42160 617763 42166 617815
rect 42218 617803 42224 617815
rect 43024 617803 43030 617815
rect 42218 617775 43030 617803
rect 42218 617763 42224 617775
rect 43024 617763 43030 617775
rect 43082 617763 43088 617815
rect 42832 616357 42838 616409
rect 42890 616397 42896 616409
rect 58192 616397 58198 616409
rect 42890 616369 58198 616397
rect 42890 616357 42896 616369
rect 58192 616357 58198 616369
rect 58250 616357 58256 616409
rect 47920 616283 47926 616335
rect 47978 616323 47984 616335
rect 58960 616323 58966 616335
rect 47978 616295 58966 616323
rect 47978 616283 47984 616295
rect 58960 616283 58966 616295
rect 59018 616283 59024 616335
rect 43408 616209 43414 616261
rect 43466 616249 43472 616261
rect 59632 616249 59638 616261
rect 43466 616221 59638 616249
rect 43466 616209 43472 616221
rect 59632 616209 59638 616221
rect 59690 616209 59696 616261
rect 42160 614803 42166 614855
rect 42218 614843 42224 614855
rect 42928 614843 42934 614855
rect 42218 614815 42934 614843
rect 42218 614803 42224 614815
rect 42928 614803 42934 614815
rect 42986 614803 42992 614855
rect 42160 614211 42166 614263
rect 42218 614251 42224 614263
rect 43120 614251 43126 614263
rect 42218 614223 43126 614251
rect 42218 614211 42224 614223
rect 43120 614211 43126 614223
rect 43178 614211 43184 614263
rect 655600 613915 655606 613967
rect 655658 613955 655664 613967
rect 676240 613955 676246 613967
rect 655658 613927 676246 613955
rect 655658 613915 655664 613927
rect 676240 613915 676246 613927
rect 676298 613915 676304 613967
rect 655408 613767 655414 613819
rect 655466 613807 655472 613819
rect 676144 613807 676150 613819
rect 655466 613779 676150 613807
rect 655466 613767 655472 613779
rect 676144 613767 676150 613779
rect 676202 613767 676208 613819
rect 655216 613619 655222 613671
rect 655274 613659 655280 613671
rect 676048 613659 676054 613671
rect 655274 613631 676054 613659
rect 655274 613619 655280 613631
rect 676048 613619 676054 613631
rect 676106 613619 676112 613671
rect 42064 613471 42070 613523
rect 42122 613511 42128 613523
rect 43024 613511 43030 613523
rect 42122 613483 43030 613511
rect 42122 613471 42128 613483
rect 43024 613471 43030 613483
rect 43082 613471 43088 613523
rect 53200 613397 53206 613449
rect 53258 613437 53264 613449
rect 59632 613437 59638 613449
rect 53258 613409 59638 613437
rect 53258 613397 53264 613409
rect 59632 613397 59638 613409
rect 59690 613397 59696 613449
rect 50320 613323 50326 613375
rect 50378 613363 50384 613375
rect 59536 613363 59542 613375
rect 50378 613335 59542 613363
rect 50378 613323 50384 613335
rect 59536 613323 59542 613335
rect 59594 613323 59600 613375
rect 673744 613175 673750 613227
rect 673802 613215 673808 613227
rect 676048 613215 676054 613227
rect 673802 613187 676054 613215
rect 673802 613175 673808 613187
rect 676048 613175 676054 613187
rect 676106 613175 676112 613227
rect 42160 612953 42166 613005
rect 42218 612993 42224 613005
rect 42832 612993 42838 613005
rect 42218 612965 42838 612993
rect 42218 612953 42224 612965
rect 42832 612953 42838 612965
rect 42890 612953 42896 613005
rect 672112 612583 672118 612635
rect 672170 612623 672176 612635
rect 676048 612623 676054 612635
rect 672170 612595 676054 612623
rect 672170 612583 672176 612595
rect 676048 612583 676054 612595
rect 676106 612583 676112 612635
rect 669808 611843 669814 611895
rect 669866 611883 669872 611895
rect 670864 611883 670870 611895
rect 669866 611855 670870 611883
rect 669866 611843 669872 611855
rect 670864 611843 670870 611855
rect 670922 611883 670928 611895
rect 676240 611883 676246 611895
rect 670922 611855 676246 611883
rect 670922 611843 670928 611855
rect 676240 611843 676246 611855
rect 676298 611843 676304 611895
rect 670576 611621 670582 611673
rect 670634 611661 670640 611673
rect 676048 611661 676054 611673
rect 670634 611633 676054 611661
rect 670634 611621 670640 611633
rect 676048 611621 676054 611633
rect 676106 611621 676112 611673
rect 669616 611103 669622 611155
rect 669674 611143 669680 611155
rect 670768 611143 670774 611155
rect 669674 611115 670774 611143
rect 669674 611103 669680 611115
rect 670768 611103 670774 611115
rect 670826 611143 670832 611155
rect 676048 611143 676054 611155
rect 670826 611115 676054 611143
rect 670826 611103 670832 611115
rect 676048 611103 676054 611115
rect 676106 611103 676112 611155
rect 670672 610585 670678 610637
rect 670730 610625 670736 610637
rect 676048 610625 676054 610637
rect 670730 610597 676054 610625
rect 670730 610585 670736 610597
rect 676048 610585 676054 610597
rect 676106 610585 676112 610637
rect 672400 607181 672406 607233
rect 672458 607221 672464 607233
rect 676048 607221 676054 607233
rect 672458 607193 676054 607221
rect 672458 607181 672464 607193
rect 676048 607181 676054 607193
rect 676106 607181 676112 607233
rect 672688 606663 672694 606715
rect 672746 606703 672752 606715
rect 676048 606703 676054 606715
rect 672746 606675 676054 606703
rect 672746 606663 672752 606675
rect 676048 606663 676054 606675
rect 676106 606663 676112 606715
rect 672976 606293 672982 606345
rect 673034 606333 673040 606345
rect 676240 606333 676246 606345
rect 673034 606305 676246 606333
rect 673034 606293 673040 606305
rect 676240 606293 676246 606305
rect 676298 606293 676304 606345
rect 672304 605701 672310 605753
rect 672362 605741 672368 605753
rect 676048 605741 676054 605753
rect 672362 605713 676054 605741
rect 672362 605701 672368 605713
rect 676048 605701 676054 605713
rect 676106 605701 676112 605753
rect 672496 605109 672502 605161
rect 672554 605149 672560 605161
rect 676048 605149 676054 605161
rect 672554 605121 676054 605149
rect 672554 605109 672560 605121
rect 676048 605109 676054 605121
rect 676106 605109 676112 605161
rect 672208 604665 672214 604717
rect 672266 604705 672272 604717
rect 676048 604705 676054 604717
rect 672266 604677 676054 604705
rect 672266 604665 672272 604677
rect 676048 604665 676054 604677
rect 676106 604665 676112 604717
rect 673072 604369 673078 604421
rect 673130 604409 673136 604421
rect 676240 604409 676246 604421
rect 673130 604381 676246 604409
rect 673130 604369 673136 604381
rect 676240 604369 676246 604381
rect 676298 604369 676304 604421
rect 673168 603629 673174 603681
rect 673226 603669 673232 603681
rect 676048 603669 676054 603681
rect 673226 603641 676054 603669
rect 673226 603629 673232 603641
rect 676048 603629 676054 603641
rect 676106 603629 676112 603681
rect 654544 602001 654550 602053
rect 654602 602041 654608 602053
rect 675376 602041 675382 602053
rect 654602 602013 675382 602041
rect 654602 602001 654608 602013
rect 675376 602001 675382 602013
rect 675434 602001 675440 602053
rect 649648 601927 649654 601979
rect 649706 601967 649712 601979
rect 679984 601967 679990 601979
rect 649706 601939 679990 601967
rect 649706 601927 649712 601939
rect 679984 601927 679990 601939
rect 680042 601927 680048 601979
rect 41776 601335 41782 601387
rect 41834 601375 41840 601387
rect 53200 601375 53206 601387
rect 41834 601347 53206 601375
rect 41834 601335 41840 601347
rect 53200 601335 53206 601347
rect 53258 601335 53264 601387
rect 41776 600743 41782 600795
rect 41834 600783 41840 600795
rect 50320 600783 50326 600795
rect 41834 600755 50326 600783
rect 41834 600743 41840 600755
rect 50320 600743 50326 600755
rect 50378 600743 50384 600795
rect 43312 600447 43318 600499
rect 43370 600487 43376 600499
rect 62320 600487 62326 600499
rect 43370 600459 62326 600487
rect 43370 600447 43376 600459
rect 62320 600447 62326 600459
rect 62378 600447 62384 600499
rect 41776 600373 41782 600425
rect 41834 600413 41840 600425
rect 43216 600413 43222 600425
rect 41834 600385 43222 600413
rect 41834 600373 41840 600385
rect 43216 600373 43222 600385
rect 43274 600373 43280 600425
rect 41776 599781 41782 599833
rect 41834 599821 41840 599833
rect 43216 599821 43222 599833
rect 41834 599793 43222 599821
rect 41834 599781 41840 599793
rect 43216 599781 43222 599793
rect 43274 599781 43280 599833
rect 39760 599411 39766 599463
rect 39818 599451 39824 599463
rect 43312 599451 43318 599463
rect 39818 599423 43318 599451
rect 39818 599411 39824 599423
rect 43312 599411 43318 599423
rect 43370 599411 43376 599463
rect 41776 599263 41782 599315
rect 41834 599303 41840 599315
rect 43312 599303 43318 599315
rect 41834 599275 43318 599303
rect 41834 599263 41840 599275
rect 43312 599263 43318 599275
rect 43370 599263 43376 599315
rect 40336 599189 40342 599241
rect 40394 599229 40400 599241
rect 62128 599229 62134 599241
rect 40394 599201 62134 599229
rect 40394 599189 40400 599201
rect 62128 599189 62134 599201
rect 62186 599189 62192 599241
rect 41584 599041 41590 599093
rect 41642 599081 41648 599093
rect 56176 599081 56182 599093
rect 41642 599053 56182 599081
rect 41642 599041 41648 599053
rect 56176 599041 56182 599053
rect 56234 599041 56240 599093
rect 41776 598301 41782 598353
rect 41834 598341 41840 598353
rect 46096 598341 46102 598353
rect 41834 598313 46102 598341
rect 41834 598301 41840 598313
rect 46096 598301 46102 598313
rect 46154 598301 46160 598353
rect 41584 596599 41590 596651
rect 41642 596639 41648 596651
rect 43120 596639 43126 596651
rect 41642 596611 43126 596639
rect 41642 596599 41648 596611
rect 43120 596599 43126 596611
rect 43178 596599 43184 596651
rect 674896 596303 674902 596355
rect 674954 596343 674960 596355
rect 675376 596343 675382 596355
rect 674954 596315 675382 596343
rect 674954 596303 674960 596315
rect 675376 596303 675382 596315
rect 675434 596303 675440 596355
rect 654160 593343 654166 593395
rect 654218 593383 654224 593395
rect 674896 593383 674902 593395
rect 654218 593355 674902 593383
rect 654218 593343 654224 593355
rect 674896 593343 674902 593355
rect 674954 593343 674960 593395
rect 673648 593269 673654 593321
rect 673706 593309 673712 593321
rect 675376 593309 675382 593321
rect 673706 593281 675382 593309
rect 673706 593269 673712 593281
rect 675376 593269 675382 593281
rect 675434 593269 675440 593321
rect 672976 592677 672982 592729
rect 673034 592717 673040 592729
rect 675472 592717 675478 592729
rect 673034 592689 675478 592717
rect 673034 592677 673040 592689
rect 675472 592677 675478 592689
rect 675530 592677 675536 592729
rect 672304 592085 672310 592137
rect 672362 592125 672368 592137
rect 675376 592125 675382 592137
rect 672362 592097 675382 592125
rect 672362 592085 672368 592097
rect 675376 592085 675382 592097
rect 675434 592085 675440 592137
rect 41776 590975 41782 591027
rect 41834 591015 41840 591027
rect 43024 591015 43030 591027
rect 41834 590987 43030 591015
rect 41834 590975 41840 590987
rect 43024 590975 43030 590987
rect 43082 590975 43088 591027
rect 41776 590827 41782 590879
rect 41834 590867 41840 590879
rect 42928 590867 42934 590879
rect 41834 590839 42934 590867
rect 41834 590827 41840 590839
rect 42928 590827 42934 590839
rect 42986 590827 42992 590879
rect 654352 590457 654358 590509
rect 654410 590497 654416 590509
rect 674992 590497 674998 590509
rect 654410 590469 674998 590497
rect 654410 590457 654416 590469
rect 674992 590457 674998 590469
rect 675050 590457 675056 590509
rect 673168 588977 673174 589029
rect 673226 589017 673232 589029
rect 675376 589017 675382 589029
rect 673226 588989 675382 589017
rect 673226 588977 673232 588989
rect 675376 588977 675382 588989
rect 675434 588977 675440 589029
rect 672208 588533 672214 588585
rect 672266 588573 672272 588585
rect 675376 588573 675382 588585
rect 672266 588545 675382 588573
rect 672266 588533 672272 588545
rect 675376 588533 675382 588545
rect 675434 588533 675440 588585
rect 674896 588089 674902 588141
rect 674954 588129 674960 588141
rect 675376 588129 675382 588141
rect 674954 588101 675382 588129
rect 674954 588089 674960 588101
rect 675376 588089 675382 588101
rect 675434 588089 675440 588141
rect 673072 587941 673078 587993
rect 673130 587981 673136 587993
rect 675472 587981 675478 587993
rect 673130 587953 675478 587981
rect 673130 587941 673136 587953
rect 675472 587941 675478 587953
rect 675530 587941 675536 587993
rect 41584 587497 41590 587549
rect 41642 587537 41648 587549
rect 56080 587537 56086 587549
rect 41642 587509 56086 587537
rect 41642 587497 41648 587509
rect 56080 587497 56086 587509
rect 56138 587497 56144 587549
rect 672688 586461 672694 586513
rect 672746 586501 672752 586513
rect 675376 586501 675382 586513
rect 672746 586473 675382 586501
rect 672746 586461 672752 586473
rect 675376 586461 675382 586473
rect 675434 586461 675440 586513
rect 674992 586239 674998 586291
rect 675050 586279 675056 586291
rect 675472 586279 675478 586291
rect 675050 586251 675478 586279
rect 675050 586239 675056 586251
rect 675472 586239 675478 586251
rect 675530 586239 675536 586291
rect 41872 584759 41878 584811
rect 41930 584759 41936 584811
rect 41890 584589 41918 584759
rect 42832 584685 42838 584737
rect 42890 584725 42896 584737
rect 58960 584725 58966 584737
rect 42890 584697 58966 584725
rect 42890 584685 42896 584697
rect 58960 584685 58966 584697
rect 59018 584685 59024 584737
rect 41872 584537 41878 584589
rect 41930 584537 41936 584589
rect 42064 582687 42070 582739
rect 42122 582727 42128 582739
rect 43120 582727 43126 582739
rect 42122 582699 43126 582727
rect 42122 582687 42128 582699
rect 43120 582687 43126 582699
rect 43178 582687 43184 582739
rect 42064 582021 42070 582073
rect 42122 582061 42128 582073
rect 42832 582061 42838 582073
rect 42122 582033 42838 582061
rect 42122 582021 42128 582033
rect 42832 582021 42838 582033
rect 42890 582021 42896 582073
rect 42064 580837 42070 580889
rect 42122 580877 42128 580889
rect 43024 580877 43030 580889
rect 42122 580849 43030 580877
rect 42122 580837 42128 580849
rect 43024 580837 43030 580849
rect 43082 580837 43088 580889
rect 42160 579579 42166 579631
rect 42218 579619 42224 579631
rect 42928 579619 42934 579631
rect 42218 579591 42934 579619
rect 42218 579579 42224 579591
rect 42928 579579 42934 579591
rect 42986 579579 42992 579631
rect 42064 579431 42070 579483
rect 42122 579471 42128 579483
rect 47920 579471 47926 579483
rect 42122 579443 47926 579471
rect 42122 579431 42128 579443
rect 47920 579431 47926 579443
rect 47978 579431 47984 579483
rect 42064 578987 42070 579039
rect 42122 579027 42128 579039
rect 42448 579027 42454 579039
rect 42122 578999 42454 579027
rect 42122 578987 42128 578999
rect 42448 578987 42454 578999
rect 42506 578987 42512 579039
rect 672112 578913 672118 578965
rect 672170 578953 672176 578965
rect 679696 578953 679702 578965
rect 672170 578925 679702 578953
rect 672170 578913 672176 578925
rect 679696 578913 679702 578925
rect 679754 578913 679760 578965
rect 42160 578247 42166 578299
rect 42218 578287 42224 578299
rect 43024 578287 43030 578299
rect 42218 578259 43030 578287
rect 42218 578247 42224 578259
rect 43024 578247 43030 578259
rect 43082 578247 43088 578299
rect 42064 577507 42070 577559
rect 42122 577547 42128 577559
rect 42928 577547 42934 577559
rect 42122 577519 42934 577547
rect 42122 577507 42128 577519
rect 42928 577507 42934 577519
rect 42986 577507 42992 577559
rect 42160 575213 42166 575265
rect 42218 575253 42224 575265
rect 42448 575253 42454 575265
rect 42218 575225 42454 575253
rect 42218 575213 42224 575225
rect 42448 575213 42454 575225
rect 42506 575213 42512 575265
rect 42160 574695 42166 574747
rect 42218 574735 42224 574747
rect 43120 574735 43126 574747
rect 42218 574707 43126 574735
rect 42218 574695 42224 574707
rect 43120 574695 43126 574707
rect 43178 574695 43184 574747
rect 42064 574029 42070 574081
rect 42122 574069 42128 574081
rect 42832 574069 42838 574081
rect 42122 574041 42838 574069
rect 42122 574029 42128 574041
rect 42832 574029 42838 574041
rect 42890 574029 42896 574081
rect 42352 573289 42358 573341
rect 42410 573289 42416 573341
rect 42160 573215 42166 573267
rect 42218 573255 42224 573267
rect 42370 573255 42398 573289
rect 42218 573227 42398 573255
rect 42218 573215 42224 573227
rect 50320 573067 50326 573119
rect 50378 573107 50384 573119
rect 58960 573107 58966 573119
rect 50378 573079 58966 573107
rect 50378 573067 50384 573079
rect 58960 573067 58966 573079
rect 59018 573067 59024 573119
rect 47920 572993 47926 573045
rect 47978 573033 47984 573045
rect 59632 573033 59638 573045
rect 47978 573005 59638 573033
rect 47978 572993 47984 573005
rect 59632 572993 59638 573005
rect 59690 572993 59696 573045
rect 42064 570995 42070 571047
rect 42122 571035 42128 571047
rect 42928 571035 42934 571047
rect 42122 571007 42934 571035
rect 42122 570995 42128 571007
rect 42928 570995 42934 571007
rect 42986 570995 42992 571047
rect 42160 570921 42166 570973
rect 42218 570961 42224 570973
rect 43024 570961 43030 570973
rect 42218 570933 43030 570961
rect 42218 570921 42224 570933
rect 43024 570921 43030 570933
rect 43082 570921 43088 570973
rect 42160 570255 42166 570307
rect 42218 570295 42224 570307
rect 42832 570295 42838 570307
rect 42218 570267 42838 570295
rect 42218 570255 42224 570267
rect 42832 570255 42838 570267
rect 42890 570255 42896 570307
rect 56176 570181 56182 570233
rect 56234 570221 56240 570233
rect 60400 570221 60406 570233
rect 56234 570193 60406 570221
rect 56234 570181 56240 570193
rect 60400 570181 60406 570193
rect 60458 570181 60464 570233
rect 53200 570107 53206 570159
rect 53258 570147 53264 570159
rect 59152 570147 59158 570159
rect 53258 570119 59158 570147
rect 53258 570107 53264 570119
rect 59152 570107 59158 570119
rect 59210 570107 59216 570159
rect 42160 569737 42166 569789
rect 42218 569777 42224 569789
rect 45040 569777 45046 569789
rect 42218 569749 45046 569777
rect 42218 569737 42224 569749
rect 45040 569737 45046 569749
rect 45098 569737 45104 569789
rect 655504 567887 655510 567939
rect 655562 567927 655568 567939
rect 676048 567927 676054 567939
rect 655562 567899 676054 567927
rect 655562 567887 655568 567899
rect 676048 567887 676054 567899
rect 676106 567887 676112 567939
rect 655312 567739 655318 567791
rect 655370 567779 655376 567791
rect 676240 567779 676246 567791
rect 655370 567751 676246 567779
rect 655370 567739 655376 567751
rect 676240 567739 676246 567751
rect 676298 567739 676304 567791
rect 670864 567443 670870 567495
rect 670922 567483 670928 567495
rect 676048 567483 676054 567495
rect 670922 567455 676054 567483
rect 670922 567443 670928 567455
rect 676048 567443 676054 567455
rect 676106 567443 676112 567495
rect 655120 567369 655126 567421
rect 655178 567409 655184 567421
rect 676144 567409 676150 567421
rect 655178 567381 676150 567409
rect 655178 567369 655184 567381
rect 676144 567369 676150 567381
rect 676202 567369 676208 567421
rect 670096 567073 670102 567125
rect 670154 567113 670160 567125
rect 670576 567113 670582 567125
rect 670154 567085 670582 567113
rect 670154 567073 670160 567085
rect 670576 567073 670582 567085
rect 670634 567113 670640 567125
rect 676240 567113 676246 567125
rect 670634 567085 676246 567113
rect 670634 567073 670640 567085
rect 676240 567073 676246 567085
rect 676298 567073 676304 567125
rect 672400 566259 672406 566311
rect 672458 566299 672464 566311
rect 676240 566299 676246 566311
rect 672458 566271 676246 566299
rect 672458 566259 672464 566271
rect 676240 566259 676246 566271
rect 676298 566259 676304 566311
rect 669904 565889 669910 565941
rect 669962 565929 669968 565941
rect 670672 565929 670678 565941
rect 669962 565901 670678 565929
rect 669962 565889 669968 565901
rect 670672 565889 670678 565901
rect 670730 565929 670736 565941
rect 676048 565929 676054 565941
rect 670730 565901 676054 565929
rect 670730 565889 670736 565901
rect 676048 565889 676054 565901
rect 676106 565889 676112 565941
rect 672496 565371 672502 565423
rect 672554 565411 672560 565423
rect 676048 565411 676054 565423
rect 672554 565383 676054 565411
rect 672554 565371 672560 565383
rect 676048 565371 676054 565383
rect 676106 565371 676112 565423
rect 670960 561449 670966 561501
rect 671018 561489 671024 561501
rect 676048 561489 676054 561501
rect 671018 561461 676054 561489
rect 671018 561449 671024 561461
rect 676048 561449 676054 561461
rect 676106 561449 676112 561501
rect 673360 560857 673366 560909
rect 673418 560897 673424 560909
rect 676048 560897 676054 560909
rect 673418 560869 676054 560897
rect 673418 560857 673424 560869
rect 676048 560857 676054 560869
rect 676106 560857 676112 560909
rect 672592 560709 672598 560761
rect 672650 560749 672656 560761
rect 676240 560749 676246 560761
rect 672650 560721 676246 560749
rect 672650 560709 672656 560721
rect 676240 560709 676246 560721
rect 676298 560709 676304 560761
rect 673264 559377 673270 559429
rect 673322 559417 673328 559429
rect 676048 559417 676054 559429
rect 673322 559389 676054 559417
rect 673322 559377 673328 559389
rect 676048 559377 676054 559389
rect 676106 559377 676112 559429
rect 672784 559007 672790 559059
rect 672842 559047 672848 559059
rect 676048 559047 676054 559059
rect 672842 559019 676054 559047
rect 672842 559007 672848 559019
rect 676048 559007 676054 559019
rect 676106 559007 676112 559059
rect 672880 558637 672886 558689
rect 672938 558677 672944 558689
rect 676240 558677 676246 558689
rect 672938 558649 676246 558677
rect 672938 558637 672944 558649
rect 676240 558637 676246 558649
rect 676298 558637 676304 558689
rect 649840 555825 649846 555877
rect 649898 555865 649904 555877
rect 679792 555865 679798 555877
rect 649898 555837 679798 555865
rect 649898 555825 649904 555837
rect 679792 555825 679798 555837
rect 679850 555825 679856 555877
rect 653776 552865 653782 552917
rect 653834 552905 653840 552917
rect 675280 552905 675286 552917
rect 653834 552877 675286 552905
rect 653834 552865 653840 552877
rect 675280 552865 675286 552877
rect 675338 552865 675344 552917
rect 672880 549091 672886 549143
rect 672938 549131 672944 549143
rect 675280 549131 675286 549143
rect 672938 549103 675286 549131
rect 672938 549091 672944 549103
rect 675280 549091 675286 549103
rect 675338 549091 675344 549143
rect 673360 547907 673366 547959
rect 673418 547947 673424 547959
rect 675472 547947 675478 547959
rect 673418 547919 675478 547947
rect 673418 547907 673424 547919
rect 675472 547907 675478 547919
rect 675530 547907 675536 547959
rect 654160 547389 654166 547441
rect 654218 547429 654224 547441
rect 674896 547429 674902 547441
rect 654218 547401 674902 547429
rect 654218 547389 654224 547401
rect 674896 547389 674902 547401
rect 674954 547389 674960 547441
rect 656272 547315 656278 547367
rect 656330 547355 656336 547367
rect 674992 547355 674998 547367
rect 656330 547327 674998 547355
rect 656330 547315 656336 547327
rect 674992 547315 674998 547327
rect 675050 547315 675056 547367
rect 673264 547241 673270 547293
rect 673322 547281 673328 547293
rect 675280 547281 675286 547293
rect 673322 547253 675286 547281
rect 673322 547241 673328 547253
rect 675280 547241 675286 547253
rect 675338 547241 675344 547293
rect 672784 544873 672790 544925
rect 672842 544913 672848 544925
rect 675472 544913 675478 544925
rect 672842 544885 675478 544913
rect 672842 544873 672848 544885
rect 675472 544873 675478 544885
rect 675530 544873 675536 544925
rect 674992 543911 674998 543963
rect 675050 543951 675056 543963
rect 675376 543951 675382 543963
rect 675050 543923 675382 543951
rect 675050 543911 675056 543923
rect 675376 543911 675382 543923
rect 675434 543911 675440 543963
rect 673840 543689 673846 543741
rect 673898 543729 673904 543741
rect 675472 543729 675478 543741
rect 673898 543701 675478 543729
rect 673898 543689 673904 543701
rect 675472 543689 675478 543701
rect 675530 543689 675536 543741
rect 675184 542283 675190 542335
rect 675242 542323 675248 542335
rect 675376 542323 675382 542335
rect 675242 542295 675382 542323
rect 675242 542283 675248 542295
rect 675376 542283 675382 542295
rect 675434 542283 675440 542335
rect 674896 542061 674902 542113
rect 674954 542101 674960 542113
rect 675376 542101 675382 542113
rect 674954 542073 675382 542101
rect 674954 542061 674960 542073
rect 675376 542061 675382 542073
rect 675434 542061 675440 542113
rect 42928 541543 42934 541595
rect 42986 541583 42992 541595
rect 57712 541583 57718 541595
rect 42986 541555 57718 541583
rect 42986 541543 42992 541555
rect 57712 541543 57718 541555
rect 57770 541543 57776 541595
rect 42832 541469 42838 541521
rect 42890 541509 42896 541521
rect 57616 541509 57622 541521
rect 42890 541481 57622 541509
rect 42890 541469 42896 541481
rect 57616 541469 57622 541481
rect 57674 541469 57680 541521
rect 673936 538583 673942 538635
rect 673994 538623 674000 538635
rect 675472 538623 675478 538635
rect 673994 538595 675478 538623
rect 673994 538583 674000 538595
rect 675472 538583 675478 538595
rect 675530 538583 675536 538635
rect 42160 538435 42166 538487
rect 42218 538475 42224 538487
rect 42928 538475 42934 538487
rect 42218 538447 42934 538475
rect 42218 538435 42224 538447
rect 42928 538435 42934 538447
rect 42986 538435 42992 538487
rect 42160 537029 42166 537081
rect 42218 537069 42224 537081
rect 42832 537069 42838 537081
rect 42218 537041 42838 537069
rect 42218 537029 42224 537041
rect 42832 537029 42838 537041
rect 42890 537029 42896 537081
rect 42160 535697 42166 535749
rect 42218 535737 42224 535749
rect 43408 535737 43414 535749
rect 42218 535709 43414 535737
rect 42218 535697 42224 535709
rect 43408 535697 43414 535709
rect 43466 535697 43472 535749
rect 42064 526373 42070 526425
rect 42122 526413 42128 526425
rect 45040 526413 45046 526425
rect 42122 526385 45046 526413
rect 42122 526373 42128 526385
rect 45040 526373 45046 526385
rect 45098 526373 45104 526425
rect 655600 524523 655606 524575
rect 655658 524563 655664 524575
rect 676240 524563 676246 524575
rect 655658 524535 676246 524563
rect 655658 524523 655664 524535
rect 676240 524523 676246 524535
rect 676298 524523 676304 524575
rect 655408 524375 655414 524427
rect 655466 524415 655472 524427
rect 676336 524415 676342 524427
rect 655466 524387 676342 524415
rect 655466 524375 655472 524387
rect 676336 524375 676342 524387
rect 676394 524375 676400 524427
rect 50320 524301 50326 524353
rect 50378 524341 50384 524353
rect 58576 524341 58582 524353
rect 50378 524313 58582 524341
rect 50378 524301 50384 524313
rect 58576 524301 58582 524313
rect 58634 524301 58640 524353
rect 47920 524227 47926 524279
rect 47978 524267 47984 524279
rect 59344 524267 59350 524279
rect 47978 524239 59350 524267
rect 47978 524227 47984 524239
rect 59344 524227 59350 524239
rect 59402 524227 59408 524279
rect 655216 524153 655222 524205
rect 655274 524193 655280 524205
rect 676144 524193 676150 524205
rect 655274 524165 676150 524193
rect 655274 524153 655280 524165
rect 676144 524153 676150 524165
rect 676202 524153 676208 524205
rect 670864 524005 670870 524057
rect 670922 524045 670928 524057
rect 676048 524045 676054 524057
rect 670922 524017 676054 524045
rect 670922 524005 670928 524017
rect 676048 524005 676054 524017
rect 676106 524005 676112 524057
rect 672400 523857 672406 523909
rect 672458 523897 672464 523909
rect 676048 523897 676054 523909
rect 672458 523869 676054 523897
rect 672458 523857 672464 523869
rect 676048 523857 676054 523869
rect 676106 523857 676112 523909
rect 672496 521193 672502 521245
rect 672554 521233 672560 521245
rect 676240 521233 676246 521245
rect 672554 521205 676246 521233
rect 672554 521193 672560 521205
rect 676240 521193 676246 521205
rect 676298 521193 676304 521245
rect 673648 517641 673654 517693
rect 673706 517681 673712 517693
rect 676240 517681 676246 517693
rect 673706 517653 676246 517681
rect 673706 517641 673712 517653
rect 676240 517641 676246 517653
rect 676298 517641 676304 517693
rect 672976 516901 672982 516953
rect 673034 516941 673040 516953
rect 676048 516941 676054 516953
rect 673034 516913 676054 516941
rect 673034 516901 673040 516913
rect 676048 516901 676054 516913
rect 676106 516901 676112 516953
rect 672688 516457 672694 516509
rect 672746 516497 672752 516509
rect 676048 516497 676054 516509
rect 672746 516469 676054 516497
rect 672746 516457 672752 516469
rect 676048 516457 676054 516469
rect 676106 516457 676112 516509
rect 672208 516161 672214 516213
rect 672266 516201 672272 516213
rect 676240 516201 676246 516213
rect 672266 516173 676246 516201
rect 672266 516161 672272 516173
rect 676240 516161 676246 516173
rect 676298 516161 676304 516213
rect 672304 515421 672310 515473
rect 672362 515461 672368 515473
rect 676048 515461 676054 515473
rect 672362 515433 676054 515461
rect 672362 515421 672368 515433
rect 676048 515421 676054 515433
rect 676106 515421 676112 515473
rect 673168 514977 673174 515029
rect 673226 515017 673232 515029
rect 676048 515017 676054 515029
rect 673226 514989 676054 515017
rect 673226 514977 673232 514989
rect 676048 514977 676054 514989
rect 676106 514977 676112 515029
rect 673072 514459 673078 514511
rect 673130 514499 673136 514511
rect 676048 514499 676054 514511
rect 673130 514471 676054 514499
rect 673130 514459 673136 514471
rect 676048 514459 676054 514471
rect 676106 514459 676112 514511
rect 649936 512683 649942 512735
rect 649994 512723 650000 512735
rect 679984 512723 679990 512735
rect 649994 512695 679990 512723
rect 649994 512683 650000 512695
rect 679984 512683 679990 512695
rect 680042 512683 680048 512735
rect 676432 485303 676438 485355
rect 676490 485343 676496 485355
rect 676624 485343 676630 485355
rect 676490 485315 676630 485343
rect 676490 485303 676496 485315
rect 676624 485303 676630 485315
rect 676682 485303 676688 485355
rect 655504 481307 655510 481359
rect 655562 481347 655568 481359
rect 676240 481347 676246 481359
rect 655562 481319 676246 481347
rect 655562 481307 655568 481319
rect 676240 481307 676246 481319
rect 676298 481307 676304 481359
rect 655312 481159 655318 481211
rect 655370 481199 655376 481211
rect 676336 481199 676342 481211
rect 655370 481171 676342 481199
rect 655370 481159 655376 481171
rect 676336 481159 676342 481171
rect 676394 481159 676400 481211
rect 655120 480937 655126 480989
rect 655178 480977 655184 480989
rect 676144 480977 676150 480989
rect 655178 480949 676150 480977
rect 655178 480937 655184 480949
rect 676144 480937 676150 480949
rect 676202 480937 676208 480989
rect 670000 479383 670006 479435
rect 670058 479423 670064 479435
rect 676432 479423 676438 479435
rect 670058 479395 676438 479423
rect 670058 479383 670064 479395
rect 676432 479383 676438 479395
rect 676490 479383 676496 479435
rect 670288 479087 670294 479139
rect 670346 479127 670352 479139
rect 676624 479127 676630 479139
rect 670346 479099 676630 479127
rect 670346 479087 670352 479099
rect 676624 479087 676630 479099
rect 676682 479087 676688 479139
rect 675280 478643 675286 478695
rect 675338 478683 675344 478695
rect 676048 478683 676054 478695
rect 675338 478655 676054 478683
rect 675338 478643 675344 478655
rect 676048 478643 676054 478655
rect 676106 478643 676112 478695
rect 673648 478347 673654 478399
rect 673706 478387 673712 478399
rect 676240 478387 676246 478399
rect 673706 478359 676246 478387
rect 673706 478347 673712 478359
rect 676240 478347 676246 478359
rect 676298 478347 676304 478399
rect 673936 476793 673942 476845
rect 673994 476833 674000 476845
rect 676048 476833 676054 476845
rect 673994 476805 676054 476833
rect 673994 476793 674000 476805
rect 676048 476793 676054 476805
rect 676106 476793 676112 476845
rect 41776 476053 41782 476105
rect 41834 476093 41840 476105
rect 50320 476093 50326 476105
rect 41834 476065 50326 476093
rect 41834 476053 41840 476065
rect 50320 476053 50326 476065
rect 50378 476053 50384 476105
rect 41776 475535 41782 475587
rect 41834 475575 41840 475587
rect 47920 475575 47926 475587
rect 41834 475547 47926 475575
rect 41834 475535 41840 475547
rect 47920 475535 47926 475547
rect 47978 475535 47984 475587
rect 672880 474647 672886 474699
rect 672938 474687 672944 474699
rect 676048 474687 676054 474699
rect 672938 474659 676054 474687
rect 672938 474647 672944 474659
rect 676048 474647 676054 474659
rect 676106 474647 676112 474699
rect 41872 474573 41878 474625
rect 41930 474613 41936 474625
rect 43216 474613 43222 474625
rect 41930 474585 43222 474613
rect 41930 474573 41936 474585
rect 43216 474573 43222 474585
rect 43274 474573 43280 474625
rect 673264 474277 673270 474329
rect 673322 474317 673328 474329
rect 676240 474317 676246 474329
rect 673322 474289 676246 474317
rect 673322 474277 673328 474289
rect 676240 474277 676246 474289
rect 676298 474277 676304 474329
rect 673360 472797 673366 472849
rect 673418 472837 673424 472849
rect 676240 472837 676246 472849
rect 673418 472809 676246 472837
rect 673418 472797 673424 472809
rect 676240 472797 676246 472809
rect 676298 472797 676304 472849
rect 41776 472353 41782 472405
rect 41834 472393 41840 472405
rect 58960 472393 58966 472405
rect 41834 472365 58966 472393
rect 41834 472353 41840 472365
rect 58960 472353 58966 472365
rect 59018 472353 59024 472405
rect 672784 472205 672790 472257
rect 672842 472245 672848 472257
rect 676048 472245 676054 472257
rect 672842 472217 676054 472245
rect 672842 472205 672848 472217
rect 676048 472205 676054 472217
rect 676106 472205 676112 472257
rect 41776 471983 41782 472035
rect 41834 472023 41840 472035
rect 46000 472023 46006 472035
rect 41834 471995 46006 472023
rect 41834 471983 41840 471995
rect 46000 471983 46006 471995
rect 46058 471983 46064 472035
rect 673840 471613 673846 471665
rect 673898 471653 673904 471665
rect 676048 471653 676054 471665
rect 673898 471625 676054 471653
rect 673898 471613 673904 471625
rect 676048 471613 676054 471625
rect 676106 471613 676112 471665
rect 650032 469467 650038 469519
rect 650090 469507 650096 469519
rect 679792 469507 679798 469519
rect 650090 469479 679798 469507
rect 650090 469467 650096 469479
rect 679792 469467 679798 469479
rect 679850 469467 679856 469519
rect 41584 465249 41590 465301
rect 41642 465289 41648 465301
rect 43408 465289 43414 465301
rect 41642 465261 43414 465289
rect 41642 465249 41648 465261
rect 43408 465249 43414 465261
rect 43466 465249 43472 465301
rect 41776 463547 41782 463599
rect 41834 463587 41840 463599
rect 47920 463587 47926 463599
rect 41834 463559 47926 463587
rect 41834 463547 41840 463559
rect 47920 463547 47926 463559
rect 47978 463547 47984 463599
rect 34480 463103 34486 463155
rect 34538 463143 34544 463155
rect 41776 463143 41782 463155
rect 34538 463115 41782 463143
rect 34538 463103 34544 463115
rect 41776 463103 41782 463115
rect 41834 463103 41840 463155
rect 673648 440607 673654 440659
rect 673706 440647 673712 440659
rect 675376 440647 675382 440659
rect 673706 440619 675382 440647
rect 673706 440607 673712 440619
rect 675376 440607 675382 440619
rect 675434 440607 675440 440659
rect 41680 432023 41686 432075
rect 41738 432063 41744 432075
rect 62512 432063 62518 432075
rect 41738 432035 62518 432063
rect 41738 432023 41744 432035
rect 62512 432023 62518 432035
rect 62570 432023 62576 432075
rect 41776 429211 41782 429263
rect 41834 429251 41840 429263
rect 53200 429251 53206 429263
rect 41834 429223 53206 429251
rect 41834 429211 41840 429223
rect 53200 429211 53206 429223
rect 53258 429211 53264 429263
rect 673840 429137 673846 429189
rect 673898 429177 673904 429189
rect 675280 429177 675286 429189
rect 673898 429149 675286 429177
rect 673898 429137 673904 429149
rect 675280 429137 675286 429149
rect 675338 429137 675344 429189
rect 41584 428471 41590 428523
rect 41642 428511 41648 428523
rect 50320 428511 50326 428523
rect 41642 428483 50326 428511
rect 41642 428471 41648 428483
rect 50320 428471 50326 428483
rect 50378 428471 50384 428523
rect 41776 428175 41782 428227
rect 41834 428215 41840 428227
rect 48112 428215 48118 428227
rect 41834 428187 48118 428215
rect 41834 428175 41840 428187
rect 48112 428175 48118 428187
rect 48170 428175 48176 428227
rect 41584 426991 41590 427043
rect 41642 427031 41648 427043
rect 43312 427031 43318 427043
rect 41642 427003 43318 427031
rect 41642 426991 41648 427003
rect 43312 426991 43318 427003
rect 43370 426991 43376 427043
rect 41776 426621 41782 426673
rect 41834 426661 41840 426673
rect 43216 426661 43222 426673
rect 41834 426633 43222 426661
rect 41834 426621 41840 426633
rect 43216 426621 43222 426633
rect 43274 426621 43280 426673
rect 39664 426251 39670 426303
rect 39722 426291 39728 426303
rect 41680 426291 41686 426303
rect 39722 426263 41686 426291
rect 39722 426251 39728 426263
rect 41680 426251 41686 426263
rect 41738 426251 41744 426303
rect 41584 420405 41590 420457
rect 41642 420445 41648 420457
rect 43408 420445 43414 420457
rect 41642 420417 43414 420445
rect 41642 420405 41648 420417
rect 43408 420405 43414 420417
rect 43466 420405 43472 420457
rect 41584 417815 41590 417867
rect 41642 417855 41648 417867
rect 42832 417855 42838 417867
rect 41642 417827 42838 417855
rect 41642 417815 41648 417827
rect 42832 417815 42838 417827
rect 42890 417815 42896 417867
rect 41584 416483 41590 416535
rect 41642 416523 41648 416535
rect 48016 416523 48022 416535
rect 41642 416495 48022 416523
rect 41642 416483 41648 416495
rect 48016 416483 48022 416495
rect 48074 416483 48080 416535
rect 41680 414633 41686 414685
rect 41738 414673 41744 414685
rect 45328 414673 45334 414685
rect 41738 414645 45334 414673
rect 41738 414633 41744 414645
rect 45328 414633 45334 414645
rect 45386 414633 45392 414685
rect 41776 413819 41782 413871
rect 41834 413819 41840 413871
rect 41794 413575 41822 413819
rect 41776 413523 41782 413575
rect 41834 413523 41840 413575
rect 42064 410119 42070 410171
rect 42122 410159 42128 410171
rect 42736 410159 42742 410171
rect 42122 410131 42742 410159
rect 42122 410119 42128 410131
rect 42736 410119 42742 410131
rect 42794 410119 42800 410171
rect 42160 409823 42166 409875
rect 42218 409863 42224 409875
rect 42832 409863 42838 409875
rect 42218 409835 42838 409863
rect 42218 409823 42224 409835
rect 42832 409823 42838 409835
rect 42890 409823 42896 409875
rect 42064 408269 42070 408321
rect 42122 408309 42128 408321
rect 42832 408309 42838 408321
rect 42122 408281 42838 408309
rect 42122 408269 42128 408281
rect 42832 408269 42838 408281
rect 42890 408269 42896 408321
rect 42736 406049 42742 406101
rect 42794 406089 42800 406101
rect 58480 406089 58486 406101
rect 42794 406061 58486 406089
rect 42794 406049 42800 406061
rect 58480 406049 58486 406061
rect 58538 406049 58544 406101
rect 42832 402793 42838 402845
rect 42890 402833 42896 402845
rect 59632 402833 59638 402845
rect 42890 402805 59638 402833
rect 42890 402793 42896 402805
rect 59632 402793 59638 402805
rect 59690 402793 59696 402845
rect 53200 400277 53206 400329
rect 53258 400317 53264 400329
rect 59728 400317 59734 400329
rect 53258 400289 59734 400317
rect 53258 400277 53264 400289
rect 59728 400277 59734 400289
rect 59786 400277 59792 400329
rect 50320 400203 50326 400255
rect 50378 400243 50384 400255
rect 59536 400243 59542 400255
rect 50378 400215 59542 400243
rect 50378 400203 50384 400215
rect 59536 400203 59542 400215
rect 59594 400203 59600 400255
rect 48112 400129 48118 400181
rect 48170 400169 48176 400181
rect 59632 400169 59638 400181
rect 48170 400141 59638 400169
rect 48170 400129 48176 400141
rect 59632 400129 59638 400141
rect 59690 400129 59696 400181
rect 655504 394727 655510 394779
rect 655562 394767 655568 394779
rect 676144 394767 676150 394779
rect 655562 394739 676150 394767
rect 655562 394727 655568 394739
rect 676144 394727 676150 394739
rect 676202 394727 676208 394779
rect 655312 394653 655318 394705
rect 655370 394693 655376 394705
rect 676240 394693 676246 394705
rect 655370 394665 676246 394693
rect 655370 394653 655376 394665
rect 676240 394653 676246 394665
rect 676298 394653 676304 394705
rect 655120 394579 655126 394631
rect 655178 394619 655184 394631
rect 676336 394619 676342 394631
rect 655178 394591 676342 394619
rect 655178 394579 655184 394591
rect 676336 394579 676342 394591
rect 676394 394579 676400 394631
rect 42160 394505 42166 394557
rect 42218 394545 42224 394557
rect 57616 394545 57622 394557
rect 42218 394517 57622 394545
rect 42218 394505 42224 394517
rect 57616 394505 57622 394517
rect 57674 394505 57680 394557
rect 672592 393839 672598 393891
rect 672650 393879 672656 393891
rect 673840 393879 673846 393891
rect 672650 393851 673846 393879
rect 672650 393839 672656 393851
rect 673840 393839 673846 393851
rect 673898 393879 673904 393891
rect 676240 393879 676246 393891
rect 673898 393851 676246 393879
rect 673898 393839 673904 393851
rect 676240 393839 676246 393851
rect 676298 393839 676304 393891
rect 675376 393173 675382 393225
rect 675434 393213 675440 393225
rect 675856 393213 675862 393225
rect 675434 393185 675862 393213
rect 675434 393173 675440 393185
rect 675856 393173 675862 393185
rect 675914 393173 675920 393225
rect 675184 391693 675190 391745
rect 675242 391733 675248 391745
rect 676240 391733 676246 391745
rect 675242 391705 676246 391733
rect 675242 391693 675248 391705
rect 676240 391693 676246 391705
rect 676298 391693 676304 391745
rect 674032 389695 674038 389747
rect 674090 389735 674096 389747
rect 676048 389735 676054 389747
rect 674090 389707 676054 389735
rect 674090 389695 674096 389707
rect 676048 389695 676054 389707
rect 676106 389695 676112 389747
rect 674608 389103 674614 389155
rect 674666 389143 674672 389155
rect 676240 389143 676246 389155
rect 674666 389115 676246 389143
rect 674666 389103 674672 389115
rect 676240 389103 676246 389115
rect 676298 389103 676304 389155
rect 674896 388881 674902 388933
rect 674954 388921 674960 388933
rect 676048 388921 676054 388933
rect 674954 388893 676054 388921
rect 674954 388881 674960 388893
rect 676048 388881 676054 388893
rect 676106 388881 676112 388933
rect 675280 388807 675286 388859
rect 675338 388847 675344 388859
rect 676240 388847 676246 388859
rect 675338 388819 676246 388847
rect 675338 388807 675344 388819
rect 676240 388807 676246 388819
rect 676298 388807 676304 388859
rect 674128 387031 674134 387083
rect 674186 387071 674192 387083
rect 676240 387071 676246 387083
rect 674186 387043 676246 387071
rect 674186 387031 674192 387043
rect 676240 387031 676246 387043
rect 676298 387031 676304 387083
rect 674512 386735 674518 386787
rect 674570 386775 674576 386787
rect 676048 386775 676054 386787
rect 674570 386747 676054 386775
rect 674570 386735 674576 386747
rect 676048 386735 676054 386747
rect 676106 386735 676112 386787
rect 674416 386291 674422 386343
rect 674474 386331 674480 386343
rect 675952 386331 675958 386343
rect 674474 386303 675958 386331
rect 674474 386291 674480 386303
rect 675952 386291 675958 386303
rect 676010 386291 676016 386343
rect 674224 386069 674230 386121
rect 674282 386109 674288 386121
rect 676240 386109 676246 386121
rect 674282 386081 676246 386109
rect 674282 386069 674288 386081
rect 676240 386069 676246 386081
rect 676298 386069 676304 386121
rect 41776 385995 41782 386047
rect 41834 386035 41840 386047
rect 53200 386035 53206 386047
rect 41834 386007 53206 386035
rect 41834 385995 41840 386007
rect 53200 385995 53206 386007
rect 53258 385995 53264 386047
rect 674704 385995 674710 386047
rect 674762 386035 674768 386047
rect 675952 386035 675958 386047
rect 674762 386007 675958 386035
rect 674762 385995 674768 386007
rect 675952 385995 675958 386007
rect 676010 385995 676016 386047
rect 674800 385921 674806 385973
rect 674858 385961 674864 385973
rect 676048 385961 676054 385973
rect 674858 385933 676054 385961
rect 674858 385921 674864 385933
rect 676048 385921 676054 385933
rect 676106 385921 676112 385973
rect 41584 385255 41590 385307
rect 41642 385295 41648 385307
rect 50320 385295 50326 385307
rect 41642 385267 50326 385295
rect 41642 385255 41648 385267
rect 50320 385255 50326 385267
rect 50378 385255 50384 385307
rect 41776 384959 41782 385011
rect 41834 384999 41840 385011
rect 48208 384999 48214 385011
rect 41834 384971 48214 384999
rect 41834 384959 41840 384971
rect 48208 384959 48214 384971
rect 48266 384959 48272 385011
rect 41584 384737 41590 384789
rect 41642 384777 41648 384789
rect 43312 384777 43318 384789
rect 41642 384749 43318 384777
rect 41642 384737 41648 384749
rect 43312 384737 43318 384749
rect 43370 384737 43376 384789
rect 41584 383775 41590 383827
rect 41642 383815 41648 383827
rect 43312 383815 43318 383827
rect 41642 383787 43318 383815
rect 41642 383775 41648 383787
rect 43312 383775 43318 383787
rect 43370 383775 43376 383827
rect 41776 383479 41782 383531
rect 41834 383519 41840 383531
rect 43504 383519 43510 383531
rect 41834 383491 43510 383519
rect 41834 383479 41840 383491
rect 43504 383479 43510 383491
rect 43562 383479 43568 383531
rect 41584 383257 41590 383309
rect 41642 383297 41648 383309
rect 43216 383297 43222 383309
rect 41642 383269 43222 383297
rect 41642 383257 41648 383269
rect 43216 383257 43222 383269
rect 43274 383297 43280 383309
rect 45232 383297 45238 383309
rect 43274 383269 45238 383297
rect 43274 383257 43280 383269
rect 45232 383257 45238 383269
rect 45290 383257 45296 383309
rect 674320 383109 674326 383161
rect 674378 383149 674384 383161
rect 676240 383149 676246 383161
rect 674378 383121 676246 383149
rect 674378 383109 674384 383121
rect 676240 383109 676246 383121
rect 676298 383109 676304 383161
rect 650128 383035 650134 383087
rect 650186 383075 650192 383087
rect 679696 383075 679702 383087
rect 650186 383047 679702 383075
rect 650186 383035 650192 383047
rect 679696 383035 679702 383047
rect 679754 383035 679760 383087
rect 666640 382961 666646 383013
rect 666698 383001 666704 383013
rect 675856 383001 675862 383013
rect 666698 382973 675862 383001
rect 666698 382961 666704 382973
rect 675856 382961 675862 382973
rect 675914 382961 675920 383013
rect 41776 381999 41782 382051
rect 41834 382039 41840 382051
rect 43408 382039 43414 382051
rect 41834 382011 43414 382039
rect 41834 381999 41840 382011
rect 43408 381999 43414 382011
rect 43466 382039 43472 382051
rect 45424 382039 45430 382051
rect 43466 382011 45430 382039
rect 43466 381999 43472 382011
rect 45424 381999 45430 382011
rect 45482 381999 45488 382051
rect 674992 379409 674998 379461
rect 675050 379449 675056 379461
rect 675472 379449 675478 379461
rect 675050 379421 675478 379449
rect 675050 379409 675056 379421
rect 675472 379409 675478 379421
rect 675530 379409 675536 379461
rect 39952 377189 39958 377241
rect 40010 377229 40016 377241
rect 43408 377229 43414 377241
rect 40010 377201 43414 377229
rect 40010 377189 40016 377201
rect 43408 377189 43414 377201
rect 43466 377189 43472 377241
rect 674608 376523 674614 376575
rect 674666 376563 674672 376575
rect 675472 376563 675478 376575
rect 674666 376535 675478 376563
rect 674666 376523 674672 376535
rect 675472 376523 675478 376535
rect 675530 376523 675536 376575
rect 674512 375635 674518 375687
rect 674570 375675 674576 375687
rect 675376 375675 675382 375687
rect 674570 375647 675382 375675
rect 674570 375635 674576 375647
rect 675376 375635 675382 375647
rect 675434 375635 675440 375687
rect 674416 375191 674422 375243
rect 674474 375231 674480 375243
rect 675472 375231 675478 375243
rect 674474 375203 675478 375231
rect 674474 375191 674480 375203
rect 675472 375191 675478 375203
rect 675530 375191 675536 375243
rect 674800 374673 674806 374725
rect 674858 374713 674864 374725
rect 675376 374713 675382 374725
rect 674858 374685 675382 374713
rect 674858 374673 674864 374685
rect 675376 374673 675382 374685
rect 675434 374673 675440 374725
rect 41584 374451 41590 374503
rect 41642 374491 41648 374503
rect 42832 374491 42838 374503
rect 41642 374463 42838 374491
rect 41642 374451 41648 374463
rect 42832 374451 42838 374463
rect 42890 374451 42896 374503
rect 41584 373267 41590 373319
rect 41642 373307 41648 373319
rect 48112 373307 48118 373319
rect 41642 373279 48118 373307
rect 41642 373267 41648 373279
rect 48112 373267 48118 373279
rect 48170 373267 48176 373319
rect 674032 372157 674038 372209
rect 674090 372197 674096 372209
rect 675376 372197 675382 372209
rect 674090 372169 675382 372197
rect 674090 372157 674096 372169
rect 675376 372157 675382 372169
rect 675434 372157 675440 372209
rect 654160 371491 654166 371543
rect 654218 371531 654224 371543
rect 674992 371531 674998 371543
rect 654218 371503 674998 371531
rect 654218 371491 654224 371503
rect 674992 371491 674998 371503
rect 675050 371491 675056 371543
rect 674704 371417 674710 371469
rect 674762 371457 674768 371469
rect 675376 371457 675382 371469
rect 674762 371429 675382 371457
rect 674762 371417 674768 371429
rect 675376 371417 675382 371429
rect 675434 371417 675440 371469
rect 674224 370973 674230 371025
rect 674282 371013 674288 371025
rect 675376 371013 675382 371025
rect 674282 370985 675382 371013
rect 674282 370973 674288 370985
rect 675376 370973 675382 370985
rect 675434 370973 675440 371025
rect 41776 370603 41782 370655
rect 41834 370603 41840 370655
rect 41794 370359 41822 370603
rect 41776 370307 41782 370359
rect 41834 370307 41840 370359
rect 674320 370307 674326 370359
rect 674378 370347 674384 370359
rect 675472 370347 675478 370359
rect 674378 370319 675478 370347
rect 674378 370307 674384 370319
rect 675472 370307 675478 370319
rect 675530 370307 675536 370359
rect 674128 369123 674134 369175
rect 674186 369163 674192 369175
rect 675376 369163 675382 369175
rect 674186 369135 675382 369163
rect 674186 369123 674192 369135
rect 675376 369123 675382 369135
rect 675434 369123 675440 369175
rect 42064 366903 42070 366955
rect 42122 366943 42128 366955
rect 42736 366943 42742 366955
rect 42122 366915 42742 366943
rect 42122 366903 42128 366915
rect 42736 366903 42742 366915
rect 42794 366903 42800 366955
rect 42160 366681 42166 366733
rect 42218 366721 42224 366733
rect 42832 366721 42838 366733
rect 42218 366693 42838 366721
rect 42218 366681 42224 366693
rect 42832 366681 42838 366693
rect 42890 366681 42896 366733
rect 674896 365423 674902 365475
rect 674954 365463 674960 365475
rect 675472 365463 675478 365475
rect 674954 365435 675478 365463
rect 674954 365423 674960 365435
rect 675472 365423 675478 365435
rect 675530 365423 675536 365475
rect 42160 365053 42166 365105
rect 42218 365093 42224 365105
rect 42832 365093 42838 365105
rect 42218 365065 42838 365093
rect 42218 365053 42224 365065
rect 42832 365053 42838 365065
rect 42890 365053 42896 365105
rect 42736 362537 42742 362589
rect 42794 362577 42800 362589
rect 58288 362577 58294 362589
rect 42794 362549 58294 362577
rect 42794 362537 42800 362549
rect 58288 362537 58294 362549
rect 58346 362537 58352 362589
rect 660304 360835 660310 360887
rect 660362 360875 660368 360887
rect 666640 360875 666646 360887
rect 660362 360847 666646 360875
rect 660362 360835 660368 360847
rect 666640 360835 666646 360847
rect 666698 360835 666704 360887
rect 42832 359947 42838 359999
rect 42890 359987 42896 359999
rect 59152 359987 59158 359999
rect 42890 359959 59158 359987
rect 42890 359947 42896 359959
rect 59152 359947 59158 359959
rect 59210 359947 59216 359999
rect 53200 357061 53206 357113
rect 53258 357101 53264 357113
rect 58192 357101 58198 357113
rect 53258 357073 58198 357101
rect 53258 357061 53264 357073
rect 58192 357061 58198 357073
rect 58250 357061 58256 357113
rect 48208 356987 48214 357039
rect 48266 357027 48272 357039
rect 59632 357027 59638 357039
rect 48266 356999 59638 357027
rect 48266 356987 48272 356999
rect 59632 356987 59638 356999
rect 59690 356987 59696 357039
rect 50320 356913 50326 356965
rect 50378 356953 50384 356965
rect 58576 356953 58582 356965
rect 50378 356925 58582 356953
rect 50378 356913 50384 356925
rect 58576 356913 58582 356925
rect 58634 356913 58640 356965
rect 655216 351585 655222 351637
rect 655274 351625 655280 351637
rect 676048 351625 676054 351637
rect 655274 351597 676054 351625
rect 655274 351585 655280 351597
rect 676048 351585 676054 351597
rect 676106 351585 676112 351637
rect 655120 351511 655126 351563
rect 655178 351551 655184 351563
rect 676240 351551 676246 351563
rect 655178 351523 676246 351551
rect 655178 351511 655184 351523
rect 676240 351511 676246 351523
rect 676298 351511 676304 351563
rect 655408 351363 655414 351415
rect 655466 351403 655472 351415
rect 660304 351403 660310 351415
rect 655466 351375 660310 351403
rect 655466 351363 655472 351375
rect 660304 351363 660310 351375
rect 660362 351363 660368 351415
rect 42160 351289 42166 351341
rect 42218 351329 42224 351341
rect 57616 351329 57622 351341
rect 42218 351301 57622 351329
rect 42218 351289 42224 351301
rect 57616 351289 57622 351301
rect 57674 351289 57680 351341
rect 655312 348477 655318 348529
rect 655370 348517 655376 348529
rect 676048 348517 676054 348529
rect 655370 348489 676054 348517
rect 655370 348477 655376 348489
rect 676048 348477 676054 348489
rect 676106 348477 676112 348529
rect 674512 345591 674518 345643
rect 674570 345631 674576 345643
rect 676048 345631 676054 345643
rect 674570 345603 676054 345631
rect 674570 345591 674576 345603
rect 676048 345591 676054 345603
rect 676106 345591 676112 345643
rect 41776 342779 41782 342831
rect 41834 342819 41840 342831
rect 53200 342819 53206 342831
rect 41834 342791 53206 342819
rect 41834 342779 41840 342791
rect 53200 342779 53206 342791
rect 53258 342779 53264 342831
rect 674416 342779 674422 342831
rect 674474 342819 674480 342831
rect 676240 342819 676246 342831
rect 674474 342791 676246 342819
rect 674474 342779 674480 342791
rect 676240 342779 676246 342791
rect 676298 342779 676304 342831
rect 674704 342705 674710 342757
rect 674762 342745 674768 342757
rect 676048 342745 676054 342757
rect 674762 342717 676054 342745
rect 674762 342705 674768 342717
rect 676048 342705 676054 342717
rect 676106 342705 676112 342757
rect 41776 342261 41782 342313
rect 41834 342301 41840 342313
rect 50320 342301 50326 342313
rect 41834 342273 50326 342301
rect 41834 342261 41840 342273
rect 50320 342261 50326 342273
rect 50378 342261 50384 342313
rect 41776 341743 41782 341795
rect 41834 341783 41840 341795
rect 48208 341783 48214 341795
rect 41834 341755 48214 341783
rect 41834 341743 41840 341755
rect 48208 341743 48214 341755
rect 48266 341743 48272 341795
rect 41776 341373 41782 341425
rect 41834 341413 41840 341425
rect 43312 341413 43318 341425
rect 41834 341385 43318 341413
rect 41834 341373 41840 341385
rect 43312 341373 43318 341385
rect 43370 341373 43376 341425
rect 674800 341151 674806 341203
rect 674858 341191 674864 341203
rect 676048 341191 676054 341203
rect 674858 341163 676054 341191
rect 674858 341151 674864 341163
rect 676048 341151 676054 341163
rect 676106 341151 676112 341203
rect 41584 340559 41590 340611
rect 41642 340599 41648 340611
rect 43216 340599 43222 340611
rect 41642 340571 43222 340599
rect 41642 340559 41648 340571
rect 43216 340559 43222 340571
rect 43274 340559 43280 340611
rect 41776 340263 41782 340315
rect 41834 340303 41840 340315
rect 46192 340303 46198 340315
rect 41834 340275 46198 340303
rect 41834 340263 41840 340275
rect 46192 340263 46198 340275
rect 46250 340263 46256 340315
rect 41584 340041 41590 340093
rect 41642 340081 41648 340093
rect 43504 340081 43510 340093
rect 41642 340053 43510 340081
rect 41642 340041 41648 340053
rect 43504 340041 43510 340053
rect 43562 340081 43568 340093
rect 44368 340081 44374 340093
rect 43562 340053 44374 340081
rect 43562 340041 43568 340053
rect 44368 340041 44374 340053
rect 44426 340041 44432 340093
rect 674608 339967 674614 340019
rect 674666 340007 674672 340019
rect 675952 340007 675958 340019
rect 674666 339979 675958 340007
rect 674666 339967 674672 339979
rect 675952 339967 675958 339979
rect 676010 339967 676016 340019
rect 674992 339893 674998 339945
rect 675050 339933 675056 339945
rect 676240 339933 676246 339945
rect 675050 339905 676246 339933
rect 675050 339893 675056 339905
rect 676240 339893 676246 339905
rect 676298 339893 676304 339945
rect 674896 339819 674902 339871
rect 674954 339859 674960 339871
rect 676048 339859 676054 339871
rect 674954 339831 676054 339859
rect 674954 339819 674960 339831
rect 676048 339819 676054 339831
rect 676106 339819 676112 339871
rect 41584 339079 41590 339131
rect 41642 339119 41648 339131
rect 46096 339119 46102 339131
rect 41642 339091 46102 339119
rect 41642 339079 41648 339091
rect 46096 339079 46102 339091
rect 46154 339079 46160 339131
rect 41776 338857 41782 338909
rect 41834 338897 41840 338909
rect 43408 338897 43414 338909
rect 41834 338869 43414 338897
rect 41834 338857 41840 338869
rect 43408 338857 43414 338869
rect 43466 338897 43472 338909
rect 44464 338897 44470 338909
rect 43466 338869 44470 338897
rect 43466 338857 43472 338869
rect 44464 338857 44470 338869
rect 44522 338857 44528 338909
rect 650224 337007 650230 337059
rect 650282 337047 650288 337059
rect 679984 337047 679990 337059
rect 650282 337019 679990 337047
rect 650282 337007 650288 337019
rect 679984 337007 679990 337019
rect 680042 337007 680048 337059
rect 674512 335305 674518 335357
rect 674570 335345 674576 335357
rect 675184 335345 675190 335357
rect 674570 335317 675190 335345
rect 674570 335305 674576 335317
rect 675184 335305 675190 335317
rect 675242 335305 675248 335357
rect 674704 334787 674710 334839
rect 674762 334827 674768 334839
rect 675376 334827 675382 334839
rect 674762 334799 675382 334827
rect 674762 334787 674768 334799
rect 675376 334787 675382 334799
rect 675434 334787 675440 334839
rect 650416 334121 650422 334173
rect 650474 334161 650480 334173
rect 655408 334161 655414 334173
rect 650474 334133 655414 334161
rect 650474 334121 650480 334133
rect 655408 334121 655414 334133
rect 655466 334121 655472 334173
rect 674416 331679 674422 331731
rect 674474 331719 674480 331731
rect 675376 331719 675382 331731
rect 674474 331691 675382 331719
rect 674474 331679 674480 331691
rect 675376 331679 675382 331691
rect 675434 331679 675440 331731
rect 674992 330421 674998 330473
rect 675050 330461 675056 330473
rect 675472 330461 675478 330473
rect 675050 330433 675478 330461
rect 675050 330421 675056 330433
rect 675472 330421 675478 330433
rect 675530 330421 675536 330473
rect 41776 330347 41782 330399
rect 41834 330387 41840 330399
rect 45520 330387 45526 330399
rect 41834 330359 45526 330387
rect 41834 330347 41840 330359
rect 45520 330347 45526 330359
rect 45578 330347 45584 330399
rect 34480 329755 34486 329807
rect 34538 329795 34544 329807
rect 41776 329795 41782 329807
rect 34538 329767 41782 329795
rect 34538 329755 34544 329767
rect 41776 329755 41782 329767
rect 41834 329755 41840 329807
rect 654160 328275 654166 328327
rect 654218 328315 654224 328327
rect 675088 328315 675094 328327
rect 654218 328287 675094 328315
rect 654218 328275 654224 328287
rect 675088 328275 675094 328287
rect 675146 328275 675152 328327
rect 41776 327165 41782 327217
rect 41834 327165 41840 327217
rect 41794 326995 41822 327165
rect 674608 327091 674614 327143
rect 674666 327131 674672 327143
rect 675472 327131 675478 327143
rect 674666 327103 675478 327131
rect 674666 327091 674672 327103
rect 675472 327091 675478 327103
rect 675530 327091 675536 327143
rect 41776 326943 41782 326995
rect 41834 326943 41840 326995
rect 674800 326795 674806 326847
rect 674858 326835 674864 326847
rect 675376 326835 675382 326847
rect 674858 326807 675382 326835
rect 674858 326795 674864 326807
rect 675376 326795 675382 326807
rect 675434 326795 675440 326847
rect 674896 326129 674902 326181
rect 674954 326169 674960 326181
rect 675376 326169 675382 326181
rect 674954 326141 675382 326169
rect 674954 326129 674960 326141
rect 675376 326129 675382 326141
rect 675434 326129 675440 326181
rect 42160 323539 42166 323591
rect 42218 323579 42224 323591
rect 42448 323579 42454 323591
rect 42218 323551 42454 323579
rect 42218 323539 42224 323551
rect 42448 323539 42454 323551
rect 42506 323539 42512 323591
rect 42160 321689 42166 321741
rect 42218 321729 42224 321741
rect 42832 321729 42838 321741
rect 42218 321701 42838 321729
rect 42218 321689 42224 321701
rect 42832 321689 42838 321701
rect 42890 321689 42896 321741
rect 42448 319617 42454 319669
rect 42506 319657 42512 319669
rect 58480 319657 58486 319669
rect 42506 319629 58486 319657
rect 42506 319617 42512 319629
rect 58480 319617 58486 319629
rect 58538 319617 58544 319669
rect 42832 316731 42838 316783
rect 42890 316771 42896 316783
rect 59152 316771 59158 316783
rect 42890 316743 59158 316771
rect 42890 316731 42896 316743
rect 59152 316731 59158 316743
rect 59210 316731 59216 316783
rect 53200 313845 53206 313897
rect 53258 313885 53264 313897
rect 59728 313885 59734 313897
rect 53258 313857 59734 313885
rect 53258 313845 53264 313857
rect 59728 313845 59734 313857
rect 59786 313845 59792 313897
rect 50320 313771 50326 313823
rect 50378 313811 50384 313823
rect 59536 313811 59542 313823
rect 50378 313783 59542 313811
rect 50378 313771 50384 313783
rect 59536 313771 59542 313783
rect 59594 313771 59600 313823
rect 48208 313697 48214 313749
rect 48266 313737 48272 313749
rect 59632 313737 59638 313749
rect 48266 313709 59638 313737
rect 48266 313697 48272 313709
rect 59632 313697 59638 313709
rect 59690 313697 59696 313749
rect 42160 308073 42166 308125
rect 42218 308113 42224 308125
rect 59056 308113 59062 308125
rect 42218 308085 59062 308113
rect 42218 308073 42224 308085
rect 59056 308073 59062 308085
rect 59114 308073 59120 308125
rect 676240 305375 676246 305387
rect 659506 305347 676246 305375
rect 654064 305261 654070 305313
rect 654122 305301 654128 305313
rect 659506 305301 659534 305347
rect 676240 305335 676246 305347
rect 676298 305335 676304 305387
rect 654122 305273 659534 305301
rect 654122 305261 654128 305273
rect 653776 305187 653782 305239
rect 653834 305227 653840 305239
rect 676240 305227 676246 305239
rect 653834 305199 676246 305227
rect 653834 305187 653840 305199
rect 676240 305187 676246 305199
rect 676298 305187 676304 305239
rect 673360 304003 673366 304055
rect 673418 304043 673424 304055
rect 676048 304043 676054 304055
rect 673418 304015 676054 304043
rect 673418 304003 673424 304015
rect 676048 304003 676054 304015
rect 676106 304003 676112 304055
rect 673168 302967 673174 303019
rect 673226 303007 673232 303019
rect 676048 303007 676054 303019
rect 673226 302979 676054 303007
rect 673226 302967 673232 302979
rect 676048 302967 676054 302979
rect 676106 302967 676112 303019
rect 45328 302301 45334 302353
rect 45386 302341 45392 302353
rect 46480 302341 46486 302353
rect 45386 302313 46486 302341
rect 45386 302301 45392 302313
rect 46480 302301 46486 302313
rect 46538 302301 46544 302353
rect 654160 302301 654166 302353
rect 654218 302341 654224 302353
rect 676240 302341 676246 302353
rect 654218 302313 676246 302341
rect 654218 302301 654224 302313
rect 676240 302301 676246 302313
rect 676298 302301 676304 302353
rect 673264 301931 673270 301983
rect 673322 301971 673328 301983
rect 676048 301971 676054 301983
rect 673322 301943 676054 301971
rect 673322 301931 673328 301943
rect 676048 301931 676054 301943
rect 676106 301931 676112 301983
rect 46192 300895 46198 300947
rect 46250 300935 46256 300947
rect 46864 300935 46870 300947
rect 46250 300907 46870 300935
rect 46250 300895 46256 300907
rect 46864 300895 46870 300907
rect 46922 300935 46928 300947
rect 62704 300935 62710 300947
rect 46922 300907 62710 300935
rect 46922 300895 46928 300907
rect 62704 300895 62710 300907
rect 62762 300895 62768 300947
rect 39664 299637 39670 299689
rect 39722 299677 39728 299689
rect 46864 299677 46870 299689
rect 39722 299649 46870 299677
rect 39722 299637 39728 299649
rect 46864 299637 46870 299649
rect 46922 299637 46928 299689
rect 41776 299563 41782 299615
rect 41834 299603 41840 299615
rect 60208 299603 60214 299615
rect 41834 299575 60214 299603
rect 41834 299563 41840 299575
rect 60208 299563 60214 299575
rect 60266 299563 60272 299615
rect 46480 299489 46486 299541
rect 46538 299529 46544 299541
rect 54544 299529 54550 299541
rect 46538 299501 54550 299529
rect 46538 299489 46544 299501
rect 54544 299489 54550 299501
rect 54602 299489 54608 299541
rect 41776 298527 41782 298579
rect 41834 298567 41840 298579
rect 52816 298567 52822 298579
rect 41834 298539 52822 298567
rect 41834 298527 41840 298539
rect 52816 298527 52822 298539
rect 52874 298527 52880 298579
rect 41776 298157 41782 298209
rect 41834 298197 41840 298209
rect 43216 298197 43222 298209
rect 41834 298169 43222 298197
rect 41834 298157 41840 298169
rect 43216 298157 43222 298169
rect 43274 298157 43280 298209
rect 46096 298083 46102 298135
rect 46154 298123 46160 298135
rect 46864 298123 46870 298135
rect 46154 298095 46870 298123
rect 46154 298083 46160 298095
rect 46864 298083 46870 298095
rect 46922 298123 46928 298135
rect 62800 298123 62806 298135
rect 46922 298095 62806 298123
rect 46922 298083 46928 298095
rect 62800 298083 62806 298095
rect 62858 298083 62864 298135
rect 41776 297565 41782 297617
rect 41834 297605 41840 297617
rect 43216 297605 43222 297617
rect 41834 297577 43222 297605
rect 41834 297565 41840 297577
rect 43216 297565 43222 297577
rect 43274 297565 43280 297617
rect 41776 297047 41782 297099
rect 41834 297087 41840 297099
rect 46192 297087 46198 297099
rect 41834 297059 46198 297087
rect 41834 297047 41840 297059
rect 46192 297047 46198 297059
rect 46250 297047 46256 297099
rect 39856 296751 39862 296803
rect 39914 296791 39920 296803
rect 46864 296791 46870 296803
rect 39914 296763 46870 296791
rect 39914 296751 39920 296763
rect 46864 296751 46870 296763
rect 46922 296751 46928 296803
rect 41584 296677 41590 296729
rect 41642 296717 41648 296729
rect 57520 296717 57526 296729
rect 41642 296689 57526 296717
rect 41642 296677 41648 296689
rect 57520 296677 57526 296689
rect 57578 296677 57584 296729
rect 675184 296677 675190 296729
rect 675242 296717 675248 296729
rect 676048 296717 676054 296729
rect 675242 296689 676054 296717
rect 675242 296677 675248 296689
rect 676048 296677 676054 296689
rect 676106 296677 676112 296729
rect 41584 295863 41590 295915
rect 41642 295903 41648 295915
rect 46288 295903 46294 295915
rect 41642 295875 46294 295903
rect 41642 295863 41648 295875
rect 46288 295863 46294 295875
rect 46346 295863 46352 295915
rect 46096 293865 46102 293917
rect 46154 293905 46160 293917
rect 59632 293905 59638 293917
rect 46154 293877 59638 293905
rect 46154 293865 46160 293877
rect 59632 293865 59638 293877
rect 59690 293865 59696 293917
rect 48976 293791 48982 293843
rect 49034 293831 49040 293843
rect 58192 293831 58198 293843
rect 49034 293803 58198 293831
rect 49034 293791 49040 293803
rect 58192 293791 58198 293803
rect 58250 293791 58256 293843
rect 674992 293791 674998 293843
rect 675050 293831 675056 293843
rect 676048 293831 676054 293843
rect 675050 293803 676054 293831
rect 675050 293791 675056 293803
rect 676048 293791 676054 293803
rect 676106 293791 676112 293843
rect 679888 291759 679894 291771
rect 659506 291731 679894 291759
rect 650320 291645 650326 291697
rect 650378 291685 650384 291697
rect 659506 291685 659534 291731
rect 679888 291719 679894 291731
rect 679946 291719 679952 291771
rect 650378 291657 659534 291685
rect 650378 291645 650384 291657
rect 52816 291275 52822 291327
rect 52874 291315 52880 291327
rect 59632 291315 59638 291327
rect 52874 291287 59638 291315
rect 52874 291275 52880 291287
rect 59632 291275 59638 291287
rect 59690 291275 59696 291327
rect 54544 290979 54550 291031
rect 54602 291019 54608 291031
rect 54602 290991 60446 291019
rect 54602 290979 54608 290991
rect 44176 290905 44182 290957
rect 44234 290945 44240 290957
rect 59056 290945 59062 290957
rect 44234 290917 59062 290945
rect 44234 290905 44240 290917
rect 59056 290905 59062 290917
rect 59114 290905 59120 290957
rect 60418 290871 60446 290991
rect 63280 290871 63286 290883
rect 60418 290843 63286 290871
rect 63280 290831 63286 290843
rect 63338 290831 63344 290883
rect 675184 290387 675190 290439
rect 675242 290427 675248 290439
rect 675376 290427 675382 290439
rect 675242 290399 675382 290427
rect 675242 290387 675248 290399
rect 675376 290387 675382 290399
rect 675434 290387 675440 290439
rect 654160 289129 654166 289181
rect 654218 289169 654224 289181
rect 660880 289169 660886 289181
rect 654218 289141 660886 289169
rect 654218 289129 654224 289141
rect 660880 289129 660886 289141
rect 660938 289129 660944 289181
rect 45808 288019 45814 288071
rect 45866 288059 45872 288071
rect 59632 288059 59638 288071
rect 45866 288031 59638 288059
rect 45866 288019 45872 288031
rect 59632 288019 59638 288031
rect 59690 288019 59696 288071
rect 656560 287945 656566 287997
rect 656618 287985 656624 287997
rect 675184 287985 675190 287997
rect 656618 287957 675190 287985
rect 656618 287945 656624 287957
rect 675184 287945 675190 287957
rect 675242 287945 675248 287997
rect 41776 287131 41782 287183
rect 41834 287171 41840 287183
rect 44272 287171 44278 287183
rect 41834 287143 44278 287171
rect 41834 287131 41840 287143
rect 44272 287131 44278 287143
rect 44330 287131 44336 287183
rect 62224 286687 62230 286739
rect 62282 286727 62288 286739
rect 62896 286727 62902 286739
rect 62282 286699 62902 286727
rect 62282 286687 62288 286699
rect 62896 286687 62902 286699
rect 62954 286687 62960 286739
rect 34480 286539 34486 286591
rect 34538 286579 34544 286591
rect 41776 286579 41782 286591
rect 34538 286551 41782 286579
rect 34538 286539 34544 286551
rect 41776 286539 41782 286551
rect 41834 286539 41840 286591
rect 674992 286243 674998 286295
rect 675050 286283 675056 286295
rect 675376 286283 675382 286295
rect 675050 286255 675382 286283
rect 675050 286243 675056 286255
rect 675376 286243 675382 286255
rect 675434 286243 675440 286295
rect 48208 285207 48214 285259
rect 48266 285247 48272 285259
rect 59536 285247 59542 285259
rect 48266 285219 59542 285247
rect 48266 285207 48272 285219
rect 59536 285207 59542 285219
rect 59594 285207 59600 285259
rect 53200 285133 53206 285185
rect 53258 285173 53264 285185
rect 58096 285173 58102 285185
rect 53258 285145 58102 285173
rect 53258 285133 53264 285145
rect 58096 285133 58102 285145
rect 58154 285133 58160 285185
rect 653776 284245 653782 284297
rect 653834 284285 653840 284297
rect 658000 284285 658006 284297
rect 653834 284257 658006 284285
rect 653834 284245 653840 284257
rect 658000 284245 658006 284257
rect 658058 284245 658064 284297
rect 41776 284023 41782 284075
rect 41834 284023 41840 284075
rect 41794 283779 41822 284023
rect 41776 283727 41782 283779
rect 41834 283727 41840 283779
rect 45328 282543 45334 282595
rect 45386 282583 45392 282595
rect 59632 282583 59638 282595
rect 45386 282555 59638 282583
rect 45386 282543 45392 282555
rect 59632 282543 59638 282555
rect 59690 282543 59696 282595
rect 45616 282321 45622 282373
rect 45674 282361 45680 282373
rect 58960 282361 58966 282373
rect 45674 282333 58966 282361
rect 45674 282321 45680 282333
rect 58960 282321 58966 282333
rect 59018 282321 59024 282373
rect 56176 282247 56182 282299
rect 56234 282287 56240 282299
rect 57616 282287 57622 282299
rect 56234 282259 57622 282287
rect 56234 282247 56240 282259
rect 57616 282247 57622 282259
rect 57674 282247 57680 282299
rect 42160 281285 42166 281337
rect 42218 281325 42224 281337
rect 46096 281325 46102 281337
rect 42218 281297 46102 281325
rect 42218 281285 42224 281297
rect 46096 281285 46102 281297
rect 46154 281285 46160 281337
rect 45712 279435 45718 279487
rect 45770 279475 45776 279487
rect 59632 279475 59638 279487
rect 45770 279447 59638 279475
rect 45770 279435 45776 279447
rect 59632 279435 59638 279447
rect 59690 279435 59696 279487
rect 45904 279361 45910 279413
rect 45962 279401 45968 279413
rect 58192 279401 58198 279413
rect 45962 279373 58198 279401
rect 45962 279361 45968 279373
rect 58192 279361 58198 279373
rect 58250 279361 58256 279413
rect 654736 279361 654742 279413
rect 654794 279401 654800 279413
rect 663760 279401 663766 279413
rect 654794 279373 663766 279401
rect 654794 279361 654800 279373
rect 663760 279361 663766 279373
rect 663818 279361 663824 279413
rect 42160 279287 42166 279339
rect 42218 279327 42224 279339
rect 48976 279327 48982 279339
rect 42218 279299 48982 279327
rect 42218 279287 42224 279299
rect 48976 279287 48982 279299
rect 49034 279287 49040 279339
rect 313552 278325 313558 278377
rect 313610 278365 313616 278377
rect 404752 278365 404758 278377
rect 313610 278337 404758 278365
rect 313610 278325 313616 278337
rect 404752 278325 404758 278337
rect 404810 278325 404816 278377
rect 314896 278251 314902 278303
rect 314954 278291 314960 278303
rect 408304 278291 408310 278303
rect 314954 278263 408310 278291
rect 314954 278251 314960 278263
rect 408304 278251 408310 278263
rect 408362 278251 408368 278303
rect 316624 278177 316630 278229
rect 316682 278217 316688 278229
rect 411856 278217 411862 278229
rect 316682 278189 411862 278217
rect 316682 278177 316688 278189
rect 411856 278177 411862 278189
rect 411914 278177 411920 278229
rect 319504 278103 319510 278155
rect 319562 278143 319568 278155
rect 418960 278143 418966 278155
rect 319562 278115 418966 278143
rect 319562 278103 319568 278115
rect 418960 278103 418966 278115
rect 419018 278103 419024 278155
rect 320944 278029 320950 278081
rect 321002 278069 321008 278081
rect 422512 278069 422518 278081
rect 321002 278041 422518 278069
rect 321002 278029 321008 278041
rect 422512 278029 422518 278041
rect 422570 278029 422576 278081
rect 322096 277955 322102 278007
rect 322154 277995 322160 278007
rect 426256 277995 426262 278007
rect 322154 277967 426262 277995
rect 322154 277955 322160 277967
rect 426256 277955 426262 277967
rect 426314 277955 426320 278007
rect 63376 277881 63382 277933
rect 63434 277921 63440 277933
rect 381232 277921 381238 277933
rect 63434 277893 381238 277921
rect 63434 277881 63440 277893
rect 381232 277881 381238 277893
rect 381290 277881 381296 277933
rect 323824 277807 323830 277859
rect 323882 277847 323888 277859
rect 429904 277847 429910 277859
rect 323882 277819 429910 277847
rect 323882 277807 323888 277819
rect 429904 277807 429910 277819
rect 429962 277807 429968 277859
rect 326416 277733 326422 277785
rect 326474 277773 326480 277785
rect 437008 277773 437014 277785
rect 326474 277745 437014 277773
rect 326474 277733 326480 277745
rect 437008 277733 437014 277745
rect 437066 277733 437072 277785
rect 317872 277659 317878 277711
rect 317930 277699 317936 277711
rect 415696 277699 415702 277711
rect 317930 277671 415702 277699
rect 317930 277659 317936 277671
rect 415696 277659 415702 277671
rect 415754 277659 415760 277711
rect 329296 277585 329302 277637
rect 329354 277625 329360 277637
rect 444112 277625 444118 277637
rect 329354 277597 444118 277625
rect 329354 277585 329360 277597
rect 444112 277585 444118 277597
rect 444170 277585 444176 277637
rect 333616 277511 333622 277563
rect 333674 277551 333680 277563
rect 454768 277551 454774 277563
rect 333674 277523 454774 277551
rect 333674 277511 333680 277523
rect 454768 277511 454774 277523
rect 454826 277511 454832 277563
rect 336688 277437 336694 277489
rect 336746 277477 336752 277489
rect 461776 277477 461782 277489
rect 336746 277449 461782 277477
rect 336746 277437 336752 277449
rect 461776 277437 461782 277449
rect 461834 277437 461840 277489
rect 339280 277363 339286 277415
rect 339338 277403 339344 277415
rect 468880 277403 468886 277415
rect 339338 277375 468886 277403
rect 339338 277363 339344 277375
rect 468880 277363 468886 277375
rect 468938 277363 468944 277415
rect 342160 277289 342166 277341
rect 342218 277329 342224 277341
rect 475984 277329 475990 277341
rect 342218 277301 475990 277329
rect 342218 277289 342224 277301
rect 475984 277289 475990 277301
rect 476042 277289 476048 277341
rect 372496 277215 372502 277267
rect 372554 277255 372560 277267
rect 550480 277255 550486 277267
rect 372554 277227 550486 277255
rect 372554 277215 372560 277227
rect 550480 277215 550486 277227
rect 550538 277215 550544 277267
rect 373840 277141 373846 277193
rect 373898 277181 373904 277193
rect 554032 277181 554038 277193
rect 373898 277153 554038 277181
rect 373898 277141 373904 277153
rect 554032 277141 554038 277153
rect 554090 277141 554096 277193
rect 376816 277067 376822 277119
rect 376874 277107 376880 277119
rect 561136 277107 561142 277119
rect 376874 277079 561142 277107
rect 376874 277067 376880 277079
rect 561136 277067 561142 277079
rect 561194 277067 561200 277119
rect 377968 276993 377974 277045
rect 378026 277033 378032 277045
rect 564688 277033 564694 277045
rect 378026 277005 564694 277033
rect 378026 276993 378032 277005
rect 564688 276993 564694 277005
rect 564746 276993 564752 277045
rect 381040 276919 381046 276971
rect 381098 276959 381104 276971
rect 571696 276959 571702 276971
rect 381098 276931 571702 276959
rect 381098 276919 381104 276931
rect 571696 276919 571702 276931
rect 571754 276919 571760 276971
rect 379408 276845 379414 276897
rect 379466 276885 379472 276897
rect 568240 276885 568246 276897
rect 379466 276857 568246 276885
rect 379466 276845 379472 276857
rect 568240 276845 568246 276857
rect 568298 276845 568304 276897
rect 383632 276771 383638 276823
rect 383690 276811 383696 276823
rect 578800 276811 578806 276823
rect 383690 276783 578806 276811
rect 383690 276771 383696 276783
rect 578800 276771 578806 276783
rect 578858 276771 578864 276823
rect 382288 276697 382294 276749
rect 382346 276737 382352 276749
rect 575248 276737 575254 276749
rect 382346 276709 575254 276737
rect 382346 276697 382352 276709
rect 575248 276697 575254 276709
rect 575306 276697 575312 276749
rect 386512 276623 386518 276675
rect 386570 276663 386576 276675
rect 585904 276663 585910 276675
rect 386570 276635 585910 276663
rect 386570 276623 386576 276635
rect 585904 276623 585910 276635
rect 585962 276623 585968 276675
rect 390832 276549 390838 276601
rect 390890 276589 390896 276601
rect 596560 276589 596566 276601
rect 390890 276561 596566 276589
rect 390890 276549 390896 276561
rect 596560 276549 596566 276561
rect 596618 276549 596624 276601
rect 393904 276475 393910 276527
rect 393962 276515 393968 276527
rect 603664 276515 603670 276527
rect 393962 276487 603670 276515
rect 393962 276475 393968 276487
rect 603664 276475 603670 276487
rect 603722 276475 603728 276527
rect 284464 276401 284470 276453
rect 284522 276441 284528 276453
rect 332944 276441 332950 276453
rect 284522 276413 332950 276441
rect 284522 276401 284528 276413
rect 332944 276401 332950 276413
rect 333002 276401 333008 276453
rect 350224 276401 350230 276453
rect 350282 276441 350288 276453
rect 496048 276441 496054 276453
rect 350282 276413 496054 276441
rect 350282 276401 350288 276413
rect 496048 276401 496054 276413
rect 496106 276401 496112 276453
rect 286096 276327 286102 276379
rect 286154 276367 286160 276379
rect 336496 276367 336502 276379
rect 286154 276339 336502 276367
rect 286154 276327 286160 276339
rect 336496 276327 336502 276339
rect 336554 276327 336560 276379
rect 356176 276327 356182 276379
rect 356234 276367 356240 276379
rect 510256 276367 510262 276379
rect 356234 276339 510262 276367
rect 356234 276327 356240 276339
rect 510256 276327 510262 276339
rect 510314 276327 510320 276379
rect 288688 276253 288694 276305
rect 288746 276293 288752 276305
rect 343600 276293 343606 276305
rect 288746 276265 343606 276293
rect 288746 276253 288752 276265
rect 343600 276253 343606 276265
rect 343658 276253 343664 276305
rect 359152 276253 359158 276305
rect 359210 276293 359216 276305
rect 517360 276293 517366 276305
rect 359210 276265 517366 276293
rect 359210 276253 359216 276265
rect 517360 276253 517366 276265
rect 517418 276253 517424 276305
rect 287344 276179 287350 276231
rect 287402 276219 287408 276231
rect 340048 276219 340054 276231
rect 287402 276191 340054 276219
rect 287402 276179 287408 276191
rect 340048 276179 340054 276191
rect 340106 276179 340112 276231
rect 361744 276179 361750 276231
rect 361802 276219 361808 276231
rect 524464 276219 524470 276231
rect 361802 276191 524470 276219
rect 361802 276179 361808 276191
rect 524464 276179 524470 276191
rect 524522 276179 524528 276231
rect 291856 276105 291862 276157
rect 291914 276145 291920 276157
rect 350704 276145 350710 276157
rect 291914 276117 350710 276145
rect 291914 276105 291920 276117
rect 350704 276105 350710 276117
rect 350762 276105 350768 276157
rect 364624 276105 364630 276157
rect 364682 276145 364688 276157
rect 531568 276145 531574 276157
rect 364682 276117 531574 276145
rect 364682 276105 364688 276117
rect 531568 276105 531574 276117
rect 531626 276105 531632 276157
rect 290320 276031 290326 276083
rect 290378 276071 290384 276083
rect 347152 276071 347158 276083
rect 290378 276043 347158 276071
rect 290378 276031 290384 276043
rect 347152 276031 347158 276043
rect 347210 276031 347216 276083
rect 367696 276031 367702 276083
rect 367754 276071 367760 276083
rect 538672 276071 538678 276083
rect 367754 276043 538678 276071
rect 367754 276031 367760 276043
rect 538672 276031 538678 276043
rect 538730 276031 538736 276083
rect 293008 275957 293014 276009
rect 293066 275997 293072 276009
rect 354256 275997 354262 276009
rect 293066 275969 354262 275997
rect 293066 275957 293072 275969
rect 354256 275957 354262 275969
rect 354314 275957 354320 276009
rect 371056 275957 371062 276009
rect 371114 275997 371120 276009
rect 546928 275997 546934 276009
rect 371114 275969 546934 275997
rect 371114 275957 371120 275969
rect 546928 275957 546934 275969
rect 546986 275957 546992 276009
rect 294640 275883 294646 275935
rect 294698 275923 294704 275935
rect 357808 275923 357814 275935
rect 294698 275895 357814 275923
rect 294698 275883 294704 275895
rect 357808 275883 357814 275895
rect 357866 275883 357872 275935
rect 370288 275883 370294 275935
rect 370346 275923 370352 275935
rect 545776 275923 545782 275935
rect 370346 275895 545782 275923
rect 370346 275883 370352 275895
rect 545776 275883 545782 275895
rect 545834 275883 545840 275935
rect 295888 275809 295894 275861
rect 295946 275849 295952 275861
rect 361360 275849 361366 275861
rect 295946 275821 361366 275849
rect 295946 275809 295952 275821
rect 361360 275809 361366 275821
rect 361418 275809 361424 275861
rect 371920 275809 371926 275861
rect 371978 275849 371984 275861
rect 549328 275849 549334 275861
rect 371978 275821 549334 275849
rect 371978 275809 371984 275821
rect 549328 275809 549334 275821
rect 549386 275809 549392 275861
rect 297328 275735 297334 275787
rect 297386 275775 297392 275787
rect 364912 275775 364918 275787
rect 297386 275747 364918 275775
rect 297386 275735 297392 275747
rect 364912 275735 364918 275747
rect 364970 275735 364976 275787
rect 374608 275735 374614 275787
rect 374666 275775 374672 275787
rect 556336 275775 556342 275787
rect 374666 275747 556342 275775
rect 374666 275735 374672 275747
rect 556336 275735 556342 275747
rect 556394 275735 556400 275787
rect 298960 275661 298966 275713
rect 299018 275701 299024 275713
rect 368464 275701 368470 275713
rect 299018 275673 368470 275701
rect 299018 275661 299024 275673
rect 368464 275661 368470 275673
rect 368522 275661 368528 275713
rect 377488 275661 377494 275713
rect 377546 275701 377552 275713
rect 563440 275701 563446 275713
rect 377546 275673 563446 275701
rect 377546 275661 377552 275673
rect 563440 275661 563446 275673
rect 563498 275661 563504 275713
rect 297808 275587 297814 275639
rect 297866 275627 297872 275639
rect 366064 275627 366070 275639
rect 297866 275599 366070 275627
rect 297866 275587 297872 275599
rect 366064 275587 366070 275599
rect 366122 275587 366128 275639
rect 380560 275587 380566 275639
rect 380618 275627 380624 275639
rect 570544 275627 570550 275639
rect 380618 275599 570550 275627
rect 380618 275587 380624 275599
rect 570544 275587 570550 275599
rect 570602 275587 570608 275639
rect 299344 275513 299350 275565
rect 299402 275553 299408 275565
rect 369616 275553 369622 275565
rect 299402 275525 369622 275553
rect 299402 275513 299408 275525
rect 369616 275513 369622 275525
rect 369674 275513 369680 275565
rect 388912 275513 388918 275565
rect 388970 275553 388976 275565
rect 591856 275553 591862 275565
rect 388970 275525 591862 275553
rect 388970 275513 388976 275525
rect 591856 275513 591862 275525
rect 591914 275513 591920 275565
rect 301840 275439 301846 275491
rect 301898 275479 301904 275491
rect 375568 275479 375574 275491
rect 301898 275451 375574 275479
rect 301898 275439 301904 275451
rect 375568 275439 375574 275451
rect 375626 275439 375632 275491
rect 387760 275439 387766 275491
rect 387818 275479 387824 275491
rect 588304 275479 588310 275491
rect 387818 275451 588310 275479
rect 387818 275439 387824 275451
rect 588304 275439 588310 275451
rect 588362 275439 588368 275491
rect 303280 275365 303286 275417
rect 303338 275405 303344 275417
rect 379120 275405 379126 275417
rect 303338 275377 379126 275405
rect 303338 275365 303344 275377
rect 379120 275365 379126 275377
rect 379178 275365 379184 275417
rect 394672 275365 394678 275417
rect 394730 275405 394736 275417
rect 606064 275405 606070 275417
rect 394730 275377 606070 275405
rect 394730 275365 394736 275377
rect 606064 275365 606070 275377
rect 606122 275365 606128 275417
rect 306160 275291 306166 275343
rect 306218 275331 306224 275343
rect 386128 275331 386134 275343
rect 306218 275303 386134 275331
rect 306218 275291 306224 275303
rect 386128 275291 386134 275303
rect 386186 275291 386192 275343
rect 398224 275291 398230 275343
rect 398282 275331 398288 275343
rect 398282 275303 407870 275331
rect 398282 275291 398288 275303
rect 308752 275217 308758 275269
rect 308810 275257 308816 275269
rect 393232 275257 393238 275269
rect 308810 275229 393238 275257
rect 308810 275217 308816 275229
rect 393232 275217 393238 275229
rect 393290 275217 393296 275269
rect 400624 275217 400630 275269
rect 400682 275257 400688 275269
rect 407842 275257 407870 275303
rect 407920 275291 407926 275343
rect 407978 275331 407984 275343
rect 613072 275331 613078 275343
rect 407978 275303 613078 275331
rect 407978 275291 407984 275303
rect 613072 275291 613078 275303
rect 613130 275291 613136 275343
rect 614320 275257 614326 275269
rect 400682 275229 407774 275257
rect 407842 275229 614326 275257
rect 400682 275217 400688 275229
rect 310384 275143 310390 275195
rect 310442 275183 310448 275195
rect 396784 275183 396790 275195
rect 310442 275155 396790 275183
rect 310442 275143 310448 275155
rect 396784 275143 396790 275155
rect 396842 275143 396848 275195
rect 403216 275143 403222 275195
rect 403274 275183 403280 275195
rect 407746 275183 407774 275229
rect 614320 275217 614326 275229
rect 614378 275217 614384 275269
rect 620176 275183 620182 275195
rect 403274 275155 407678 275183
rect 407746 275155 620182 275183
rect 403274 275143 403280 275155
rect 313072 275069 313078 275121
rect 313130 275109 313136 275121
rect 403888 275109 403894 275121
rect 313130 275081 403894 275109
rect 313130 275069 313136 275081
rect 403888 275069 403894 275081
rect 403946 275069 403952 275121
rect 406384 275069 406390 275121
rect 406442 275109 406448 275121
rect 407650 275109 407678 275155
rect 620176 275143 620182 275155
rect 620234 275143 620240 275195
rect 627280 275109 627286 275121
rect 406442 275081 407582 275109
rect 407650 275081 627286 275109
rect 406442 275069 406448 275081
rect 314704 274995 314710 275047
rect 314762 275035 314768 275047
rect 407440 275035 407446 275047
rect 314762 275007 407446 275035
rect 314762 274995 314768 275007
rect 407440 274995 407446 275007
rect 407498 274995 407504 275047
rect 407554 275035 407582 275081
rect 627280 275069 627286 275081
rect 627338 275069 627344 275121
rect 634384 275035 634390 275047
rect 407554 275007 634390 275035
rect 634384 274995 634390 275007
rect 634442 274995 634448 275047
rect 283024 274921 283030 274973
rect 283082 274961 283088 274973
rect 329392 274961 329398 274973
rect 283082 274933 329398 274961
rect 283082 274921 283088 274933
rect 329392 274921 329398 274933
rect 329450 274921 329456 274973
rect 344560 274921 344566 274973
rect 344618 274961 344624 274973
rect 481936 274961 481942 274973
rect 344618 274933 481942 274961
rect 344618 274921 344624 274933
rect 481936 274921 481942 274933
rect 481994 274921 482000 274973
rect 281776 274847 281782 274899
rect 281834 274887 281840 274899
rect 325840 274887 325846 274899
rect 281834 274859 325846 274887
rect 281834 274847 281840 274859
rect 325840 274847 325846 274859
rect 325898 274847 325904 274899
rect 341680 274847 341686 274899
rect 341738 274887 341744 274899
rect 474832 274887 474838 274899
rect 341738 274859 474838 274887
rect 341738 274847 341744 274859
rect 474832 274847 474838 274859
rect 474890 274847 474896 274899
rect 339088 274773 339094 274825
rect 339146 274813 339152 274825
rect 467728 274813 467734 274825
rect 339146 274785 467734 274813
rect 339146 274773 339152 274785
rect 467728 274773 467734 274785
rect 467786 274773 467792 274825
rect 336016 274699 336022 274751
rect 336074 274739 336080 274751
rect 460624 274739 460630 274751
rect 336074 274711 460630 274739
rect 336074 274699 336080 274711
rect 460624 274699 460630 274711
rect 460682 274699 460688 274751
rect 333136 274625 333142 274677
rect 333194 274665 333200 274677
rect 453520 274665 453526 274677
rect 333194 274637 453526 274665
rect 333194 274625 333200 274637
rect 453520 274625 453526 274637
rect 453578 274625 453584 274677
rect 331888 274551 331894 274603
rect 331946 274591 331952 274603
rect 449968 274591 449974 274603
rect 331946 274563 449974 274591
rect 331946 274551 331952 274563
rect 449968 274551 449974 274563
rect 450026 274551 450032 274603
rect 328816 274477 328822 274529
rect 328874 274517 328880 274529
rect 442864 274517 442870 274529
rect 328874 274489 442870 274517
rect 328874 274477 328880 274489
rect 442864 274477 442870 274489
rect 442922 274477 442928 274529
rect 325936 274403 325942 274455
rect 325994 274443 326000 274455
rect 435856 274443 435862 274455
rect 325994 274415 435862 274443
rect 325994 274403 326000 274415
rect 435856 274403 435862 274415
rect 435914 274403 435920 274455
rect 321616 274329 321622 274381
rect 321674 274369 321680 274381
rect 425200 274369 425206 274381
rect 321674 274341 425206 274369
rect 321674 274329 321680 274341
rect 425200 274329 425206 274341
rect 425258 274329 425264 274381
rect 323344 274255 323350 274307
rect 323402 274295 323408 274307
rect 428752 274295 428758 274307
rect 323402 274267 428758 274295
rect 323402 274255 323408 274267
rect 428752 274255 428758 274267
rect 428810 274255 428816 274307
rect 318928 274181 318934 274233
rect 318986 274221 318992 274233
rect 418096 274221 418102 274233
rect 318986 274193 418102 274221
rect 318986 274181 318992 274193
rect 418096 274181 418102 274193
rect 418154 274181 418160 274233
rect 317296 274107 317302 274159
rect 317354 274147 317360 274159
rect 414544 274147 414550 274159
rect 317354 274119 414550 274147
rect 317354 274107 317360 274119
rect 414544 274107 414550 274119
rect 414602 274107 414608 274159
rect 347056 274033 347062 274085
rect 347114 274073 347120 274085
rect 401488 274073 401494 274085
rect 347114 274045 401494 274073
rect 347114 274033 347120 274045
rect 401488 274033 401494 274045
rect 401546 274033 401552 274085
rect 334288 273959 334294 274011
rect 334346 273999 334352 274011
rect 387376 273999 387382 274011
rect 334346 273971 387382 273999
rect 334346 273959 334352 273971
rect 387376 273959 387382 273971
rect 387434 273959 387440 274011
rect 397552 273959 397558 274011
rect 397610 273999 397616 274011
rect 407920 273999 407926 274011
rect 397610 273971 407926 273999
rect 397610 273959 397616 273971
rect 407920 273959 407926 273971
rect 407978 273959 407984 274011
rect 328336 273885 328342 273937
rect 328394 273925 328400 273937
rect 380272 273925 380278 273937
rect 328394 273897 380278 273925
rect 328394 273885 328400 273897
rect 380272 273885 380278 273897
rect 380330 273885 380336 273937
rect 343600 273811 343606 273863
rect 343658 273851 343664 273863
rect 394480 273851 394486 273863
rect 343658 273823 394486 273851
rect 343658 273811 343664 273823
rect 394480 273811 394486 273823
rect 394538 273811 394544 273863
rect 326800 273737 326806 273789
rect 326858 273777 326864 273789
rect 373168 273777 373174 273789
rect 326858 273749 373174 273777
rect 326858 273737 326864 273749
rect 373168 273737 373174 273749
rect 373226 273737 373232 273789
rect 673168 273663 673174 273715
rect 673226 273703 673232 273715
rect 679696 273703 679702 273715
rect 673226 273675 679702 273703
rect 673226 273663 673232 273675
rect 679696 273663 679702 273675
rect 679754 273663 679760 273715
rect 673264 273589 673270 273641
rect 673322 273629 673328 273641
rect 679792 273629 679798 273641
rect 673322 273601 679798 273629
rect 673322 273589 673328 273601
rect 679792 273589 679798 273601
rect 679850 273589 679856 273641
rect 160432 273515 160438 273567
rect 160490 273555 160496 273567
rect 207472 273555 207478 273567
rect 160490 273527 207478 273555
rect 160490 273515 160496 273527
rect 207472 273515 207478 273527
rect 207530 273515 207536 273567
rect 277744 273515 277750 273567
rect 277802 273555 277808 273567
rect 316432 273555 316438 273567
rect 277802 273527 316438 273555
rect 277802 273515 277808 273527
rect 316432 273515 316438 273527
rect 316490 273515 316496 273567
rect 349456 273515 349462 273567
rect 349514 273555 349520 273567
rect 493744 273555 493750 273567
rect 349514 273527 493750 273555
rect 349514 273515 349520 273527
rect 493744 273515 493750 273527
rect 493802 273515 493808 273567
rect 529840 273515 529846 273567
rect 529898 273555 529904 273567
rect 624976 273555 624982 273567
rect 529898 273527 624982 273555
rect 529898 273515 529904 273527
rect 624976 273515 624982 273527
rect 625034 273515 625040 273567
rect 108400 273441 108406 273493
rect 108458 273481 108464 273493
rect 109360 273481 109366 273493
rect 108458 273453 109366 273481
rect 108458 273441 108464 273453
rect 109360 273441 109366 273453
rect 109418 273441 109424 273493
rect 130864 273441 130870 273493
rect 130922 273481 130928 273493
rect 190096 273481 190102 273493
rect 130922 273453 190102 273481
rect 130922 273441 130928 273453
rect 190096 273441 190102 273453
rect 190154 273441 190160 273493
rect 193552 273441 193558 273493
rect 193610 273481 193616 273493
rect 221488 273481 221494 273493
rect 193610 273453 221494 273481
rect 193610 273441 193616 273453
rect 221488 273441 221494 273453
rect 221546 273441 221552 273493
rect 230128 273441 230134 273493
rect 230186 273481 230192 273493
rect 242896 273481 242902 273493
rect 230186 273453 242902 273481
rect 230186 273441 230192 273453
rect 242896 273441 242902 273453
rect 242954 273441 242960 273493
rect 275344 273441 275350 273493
rect 275402 273481 275408 273493
rect 310480 273481 310486 273493
rect 275402 273453 310486 273481
rect 275402 273441 275408 273453
rect 310480 273441 310486 273453
rect 310538 273441 310544 273493
rect 310576 273441 310582 273493
rect 310634 273481 310640 273493
rect 344752 273481 344758 273493
rect 310634 273453 344758 273481
rect 310634 273441 310640 273453
rect 344752 273441 344758 273453
rect 344810 273441 344816 273493
rect 350032 273441 350038 273493
rect 350090 273481 350096 273493
rect 494896 273481 494902 273493
rect 350090 273453 494902 273481
rect 350090 273441 350096 273453
rect 494896 273441 494902 273453
rect 494954 273441 494960 273493
rect 122608 273367 122614 273419
rect 122666 273407 122672 273419
rect 123760 273407 123766 273419
rect 122666 273379 123766 273407
rect 122666 273367 122672 273379
rect 123760 273367 123766 273379
rect 123818 273367 123824 273419
rect 142672 273367 142678 273419
rect 142730 273407 142736 273419
rect 209584 273407 209590 273419
rect 142730 273379 209590 273407
rect 142730 273367 142736 273379
rect 209584 273367 209590 273379
rect 209642 273367 209648 273419
rect 277072 273367 277078 273419
rect 277130 273407 277136 273419
rect 314032 273407 314038 273419
rect 277130 273379 314038 273407
rect 277130 273367 277136 273379
rect 314032 273367 314038 273379
rect 314090 273367 314096 273419
rect 337936 273367 337942 273419
rect 337994 273407 338000 273419
rect 341296 273407 341302 273419
rect 337994 273379 341302 273407
rect 337994 273367 338000 273379
rect 341296 273367 341302 273379
rect 341354 273367 341360 273419
rect 352432 273367 352438 273419
rect 352490 273407 352496 273419
rect 500848 273407 500854 273419
rect 352490 273379 500854 273407
rect 352490 273367 352496 273379
rect 500848 273367 500854 273379
rect 500906 273367 500912 273419
rect 135568 273293 135574 273345
rect 135626 273333 135632 273345
rect 209872 273333 209878 273345
rect 135626 273305 209878 273333
rect 135626 273293 135632 273305
rect 209872 273293 209878 273305
rect 209930 273293 209936 273345
rect 219568 273293 219574 273345
rect 219626 273333 219632 273345
rect 238672 273333 238678 273345
rect 219626 273305 238678 273333
rect 219626 273293 219632 273305
rect 238672 273293 238678 273305
rect 238730 273293 238736 273345
rect 279664 273293 279670 273345
rect 279722 273333 279728 273345
rect 321136 273333 321142 273345
rect 279722 273305 321142 273333
rect 279722 273293 279728 273305
rect 321136 273293 321142 273305
rect 321194 273293 321200 273345
rect 352624 273293 352630 273345
rect 352682 273333 352688 273345
rect 502000 273333 502006 273345
rect 352682 273305 502006 273333
rect 352682 273293 352688 273305
rect 502000 273293 502006 273305
rect 502058 273293 502064 273345
rect 68272 273219 68278 273271
rect 68330 273259 68336 273271
rect 142480 273259 142486 273271
rect 68330 273231 142486 273259
rect 68330 273219 68336 273231
rect 142480 273219 142486 273231
rect 142538 273219 142544 273271
rect 153328 273219 153334 273271
rect 153386 273259 153392 273271
rect 207376 273259 207382 273271
rect 153386 273231 207382 273259
rect 153386 273219 153392 273231
rect 207376 273219 207382 273231
rect 207434 273219 207440 273271
rect 278224 273219 278230 273271
rect 278282 273259 278288 273271
rect 317584 273259 317590 273271
rect 278282 273231 317590 273259
rect 278282 273219 278288 273231
rect 317584 273219 317590 273231
rect 317642 273219 317648 273271
rect 355504 273219 355510 273271
rect 355562 273259 355568 273271
rect 509104 273259 509110 273271
rect 355562 273231 509110 273259
rect 355562 273219 355568 273231
rect 509104 273219 509110 273231
rect 509162 273219 509168 273271
rect 132016 273145 132022 273197
rect 132074 273185 132080 273197
rect 209680 273185 209686 273197
rect 132074 273157 209686 273185
rect 132074 273145 132080 273157
rect 209680 273145 209686 273157
rect 209738 273145 209744 273197
rect 285616 273145 285622 273197
rect 285674 273185 285680 273197
rect 335344 273185 335350 273197
rect 285674 273157 335350 273185
rect 285674 273145 285680 273157
rect 335344 273145 335350 273157
rect 335402 273145 335408 273197
rect 355024 273145 355030 273197
rect 355082 273185 355088 273197
rect 507952 273185 507958 273197
rect 355082 273157 507958 273185
rect 355082 273145 355088 273157
rect 507952 273145 507958 273157
rect 508010 273145 508016 273197
rect 127312 273071 127318 273123
rect 127370 273111 127376 273123
rect 209968 273111 209974 273123
rect 127370 273083 209974 273111
rect 127370 273071 127376 273083
rect 209968 273071 209974 273083
rect 210026 273071 210032 273123
rect 220720 273071 220726 273123
rect 220778 273111 220784 273123
rect 239152 273111 239158 273123
rect 220778 273083 239158 273111
rect 220778 273071 220784 273083
rect 239152 273071 239158 273083
rect 239210 273071 239216 273123
rect 286768 273071 286774 273123
rect 286826 273111 286832 273123
rect 338896 273111 338902 273123
rect 286826 273083 338902 273111
rect 286826 273071 286832 273083
rect 338896 273071 338902 273083
rect 338954 273071 338960 273123
rect 358576 273071 358582 273123
rect 358634 273111 358640 273123
rect 358634 273083 375134 273111
rect 358634 273071 358640 273083
rect 125008 272997 125014 273049
rect 125066 273037 125072 273049
rect 207280 273037 207286 273049
rect 125066 273009 207286 273037
rect 125066 272997 125072 273009
rect 207280 272997 207286 273009
rect 207338 272997 207344 273049
rect 217168 272997 217174 273049
rect 217226 273037 217232 273049
rect 237616 273037 237622 273049
rect 217226 273009 237622 273037
rect 217226 272997 217232 273009
rect 237616 272997 237622 273009
rect 237674 272997 237680 273049
rect 284944 272997 284950 273049
rect 285002 273037 285008 273049
rect 334192 273037 334198 273049
rect 285002 273009 334198 273037
rect 285002 272997 285008 273009
rect 334192 272997 334198 273009
rect 334250 272997 334256 273049
rect 360976 272997 360982 273049
rect 361034 273037 361040 273049
rect 375106 273037 375134 273083
rect 375184 273071 375190 273123
rect 375242 273111 375248 273123
rect 514960 273111 514966 273123
rect 375242 273083 514966 273111
rect 375242 273071 375248 273083
rect 514960 273071 514966 273083
rect 515018 273071 515024 273123
rect 516208 273037 516214 273049
rect 361034 273009 375038 273037
rect 375106 273009 516214 273037
rect 361034 272997 361040 273009
rect 128464 272923 128470 272975
rect 128522 272963 128528 272975
rect 210160 272963 210166 272975
rect 128522 272935 210166 272963
rect 128522 272923 128528 272935
rect 210160 272923 210166 272935
rect 210218 272923 210224 272975
rect 216016 272923 216022 272975
rect 216074 272963 216080 272975
rect 236944 272963 236950 272975
rect 216074 272935 236950 272963
rect 216074 272923 216080 272935
rect 236944 272923 236950 272935
rect 237002 272923 237008 272975
rect 271024 272923 271030 272975
rect 271082 272963 271088 272975
rect 299920 272963 299926 272975
rect 271082 272935 299926 272963
rect 271082 272923 271088 272935
rect 299920 272923 299926 272935
rect 299978 272923 299984 272975
rect 305392 272923 305398 272975
rect 305450 272963 305456 272975
rect 358960 272963 358966 272975
rect 305450 272935 358966 272963
rect 305450 272923 305456 272935
rect 358960 272923 358966 272935
rect 359018 272923 359024 272975
rect 361264 272923 361270 272975
rect 361322 272963 361328 272975
rect 375010 272963 375038 273009
rect 516208 272997 516214 273009
rect 516266 272997 516272 273049
rect 522064 272963 522070 272975
rect 361322 272935 374942 272963
rect 375010 272935 522070 272963
rect 361322 272923 361328 272935
rect 123664 272849 123670 272901
rect 123722 272889 123728 272901
rect 209008 272889 209014 272901
rect 123722 272861 209014 272889
rect 123722 272849 123728 272861
rect 209008 272849 209014 272861
rect 209066 272849 209072 272901
rect 218320 272849 218326 272901
rect 218378 272889 218384 272901
rect 238096 272889 238102 272901
rect 218378 272861 238102 272889
rect 218378 272849 218384 272861
rect 238096 272849 238102 272861
rect 238154 272849 238160 272901
rect 289936 272849 289942 272901
rect 289994 272889 290000 272901
rect 346000 272889 346006 272901
rect 289994 272861 346006 272889
rect 289994 272849 290000 272861
rect 346000 272849 346006 272861
rect 346058 272849 346064 272901
rect 363568 272849 363574 272901
rect 363626 272889 363632 272901
rect 374914 272889 374942 272935
rect 522064 272923 522070 272935
rect 522122 272923 522128 272975
rect 523312 272889 523318 272901
rect 363626 272861 374846 272889
rect 374914 272861 523318 272889
rect 363626 272849 363632 272861
rect 116656 272775 116662 272827
rect 116714 272815 116720 272827
rect 207088 272815 207094 272827
rect 116714 272787 207094 272815
rect 116714 272775 116720 272787
rect 207088 272775 207094 272787
rect 207146 272775 207152 272827
rect 214768 272775 214774 272827
rect 214826 272815 214832 272827
rect 236464 272815 236470 272827
rect 214826 272787 236470 272815
rect 214826 272775 214832 272787
rect 236464 272775 236470 272787
rect 236522 272775 236528 272827
rect 292240 272775 292246 272827
rect 292298 272815 292304 272827
rect 351856 272815 351862 272827
rect 292298 272787 351862 272815
rect 292298 272775 292304 272787
rect 351856 272775 351862 272787
rect 351914 272775 351920 272827
rect 364144 272775 364150 272827
rect 364202 272815 364208 272827
rect 374818 272815 374846 272861
rect 523312 272849 523318 272861
rect 523370 272849 523376 272901
rect 529168 272815 529174 272827
rect 364202 272787 374750 272815
rect 374818 272787 529174 272815
rect 364202 272775 364208 272787
rect 120208 272701 120214 272753
rect 120266 272741 120272 272753
rect 207856 272741 207862 272753
rect 120266 272713 207862 272741
rect 120266 272701 120272 272713
rect 207856 272701 207862 272713
rect 207914 272701 207920 272753
rect 212464 272701 212470 272753
rect 212522 272741 212528 272753
rect 235696 272741 235702 272753
rect 212522 272713 235702 272741
rect 212522 272701 212528 272713
rect 235696 272701 235702 272713
rect 235754 272701 235760 272753
rect 292720 272701 292726 272753
rect 292778 272741 292784 272753
rect 353104 272741 353110 272753
rect 292778 272713 353110 272741
rect 292778 272701 292784 272713
rect 353104 272701 353110 272713
rect 353162 272701 353168 272753
rect 366544 272701 366550 272753
rect 366602 272741 366608 272753
rect 374722 272741 374750 272787
rect 529168 272775 529174 272787
rect 529226 272775 529232 272827
rect 530416 272741 530422 272753
rect 366602 272713 374654 272741
rect 374722 272713 530422 272741
rect 366602 272701 366608 272713
rect 113104 272627 113110 272679
rect 113162 272667 113168 272679
rect 206032 272667 206038 272679
rect 113162 272639 206038 272667
rect 113162 272627 113168 272639
rect 206032 272627 206038 272639
rect 206090 272627 206096 272679
rect 213616 272627 213622 272679
rect 213674 272667 213680 272679
rect 236272 272667 236278 272679
rect 213674 272639 236278 272667
rect 213674 272627 213680 272639
rect 236272 272627 236278 272639
rect 236330 272627 236336 272679
rect 295408 272627 295414 272679
rect 295466 272667 295472 272679
rect 360208 272667 360214 272679
rect 295466 272639 360214 272667
rect 295466 272627 295472 272639
rect 360208 272627 360214 272639
rect 360266 272627 360272 272679
rect 367120 272627 367126 272679
rect 367178 272667 367184 272679
rect 374626 272667 374654 272713
rect 530416 272701 530422 272713
rect 530474 272701 530480 272753
rect 536272 272667 536278 272679
rect 367178 272639 374558 272667
rect 374626 272639 536278 272667
rect 367178 272627 367184 272639
rect 110800 272553 110806 272605
rect 110858 272593 110864 272605
rect 205744 272593 205750 272605
rect 110858 272565 205750 272593
rect 110858 272553 110864 272565
rect 205744 272553 205750 272565
rect 205802 272553 205808 272605
rect 211216 272553 211222 272605
rect 211274 272593 211280 272605
rect 235024 272593 235030 272605
rect 211274 272565 235030 272593
rect 211274 272553 211280 272565
rect 235024 272553 235030 272565
rect 235082 272553 235088 272605
rect 270256 272553 270262 272605
rect 270314 272593 270320 272605
rect 297520 272593 297526 272605
rect 270314 272565 297526 272593
rect 270314 272553 270320 272565
rect 297520 272553 297526 272565
rect 297578 272553 297584 272605
rect 298288 272553 298294 272605
rect 298346 272593 298352 272605
rect 367216 272593 367222 272605
rect 298346 272565 367222 272593
rect 298346 272553 298352 272565
rect 367216 272553 367222 272565
rect 367274 272553 367280 272605
rect 372688 272553 372694 272605
rect 372746 272593 372752 272605
rect 374530 272593 374558 272639
rect 536272 272627 536278 272639
rect 536330 272627 536336 272679
rect 537424 272593 537430 272605
rect 372746 272565 374462 272593
rect 374530 272565 537430 272593
rect 372746 272553 372752 272565
rect 106096 272479 106102 272531
rect 106154 272519 106160 272531
rect 204016 272519 204022 272531
rect 106154 272491 204022 272519
rect 106154 272479 106160 272491
rect 204016 272479 204022 272491
rect 204074 272479 204080 272531
rect 208912 272479 208918 272531
rect 208970 272519 208976 272531
rect 234352 272519 234358 272531
rect 208970 272491 234358 272519
rect 208970 272479 208976 272491
rect 234352 272479 234358 272491
rect 234410 272479 234416 272531
rect 270544 272479 270550 272531
rect 270602 272519 270608 272531
rect 298672 272519 298678 272531
rect 270602 272491 298678 272519
rect 270602 272479 270608 272491
rect 298672 272479 298678 272491
rect 298730 272479 298736 272531
rect 301360 272479 301366 272531
rect 301418 272519 301424 272531
rect 374320 272519 374326 272531
rect 301418 272491 374326 272519
rect 301418 272479 301424 272491
rect 374320 272479 374326 272491
rect 374378 272479 374384 272531
rect 374434 272519 374462 272565
rect 537424 272553 537430 272565
rect 537482 272553 537488 272605
rect 551632 272519 551638 272531
rect 374434 272491 551638 272519
rect 551632 272479 551638 272491
rect 551690 272479 551696 272531
rect 103696 272405 103702 272457
rect 103754 272445 103760 272457
rect 203536 272445 203542 272457
rect 103754 272417 203542 272445
rect 103754 272405 103760 272417
rect 203536 272405 203542 272417
rect 203594 272405 203600 272457
rect 210064 272405 210070 272457
rect 210122 272445 210128 272457
rect 234544 272445 234550 272457
rect 210122 272417 234550 272445
rect 210122 272405 210128 272417
rect 234544 272405 234550 272417
rect 234602 272405 234608 272457
rect 236080 272405 236086 272457
rect 236138 272445 236144 272457
rect 245296 272445 245302 272457
rect 236138 272417 245302 272445
rect 236138 272405 236144 272417
rect 245296 272405 245302 272417
rect 245354 272405 245360 272457
rect 274192 272405 274198 272457
rect 274250 272445 274256 272457
rect 306928 272445 306934 272457
rect 274250 272417 306934 272445
rect 274250 272405 274256 272417
rect 306928 272405 306934 272417
rect 306986 272405 306992 272457
rect 307120 272405 307126 272457
rect 307178 272445 307184 272457
rect 388528 272445 388534 272457
rect 307178 272417 388534 272445
rect 307178 272405 307184 272417
rect 388528 272405 388534 272417
rect 388586 272405 388592 272457
rect 388624 272405 388630 272457
rect 388682 272445 388688 272457
rect 572944 272445 572950 272457
rect 388682 272417 572950 272445
rect 388682 272405 388688 272417
rect 572944 272405 572950 272417
rect 573002 272405 573008 272457
rect 98992 272331 98998 272383
rect 99050 272371 99056 272383
rect 199120 272371 199126 272383
rect 99050 272343 199126 272371
rect 99050 272331 99056 272343
rect 199120 272331 199126 272343
rect 199178 272331 199184 272383
rect 207664 272331 207670 272383
rect 207722 272371 207728 272383
rect 233872 272371 233878 272383
rect 207722 272343 233878 272371
rect 207722 272331 207728 272343
rect 233872 272331 233878 272343
rect 233930 272331 233936 272383
rect 234928 272331 234934 272383
rect 234986 272371 234992 272383
rect 244816 272371 244822 272383
rect 234986 272343 244822 272371
rect 234986 272331 234992 272343
rect 244816 272331 244822 272343
rect 244874 272331 244880 272383
rect 272752 272331 272758 272383
rect 272810 272371 272816 272383
rect 303472 272371 303478 272383
rect 272810 272343 303478 272371
rect 272810 272331 272816 272343
rect 303472 272331 303478 272343
rect 303530 272331 303536 272383
rect 303952 272331 303958 272383
rect 304010 272371 304016 272383
rect 381424 272371 381430 272383
rect 304010 272343 381430 272371
rect 304010 272331 304016 272343
rect 381424 272331 381430 272343
rect 381482 272331 381488 272383
rect 383440 272331 383446 272383
rect 383498 272371 383504 272383
rect 577648 272371 577654 272383
rect 383498 272343 577654 272371
rect 383498 272331 383504 272343
rect 577648 272331 577654 272343
rect 577706 272331 577712 272383
rect 96592 272257 96598 272309
rect 96650 272297 96656 272309
rect 201616 272297 201622 272309
rect 96650 272269 201622 272297
rect 96650 272257 96656 272269
rect 201616 272257 201622 272269
rect 201674 272257 201680 272309
rect 232528 272257 232534 272309
rect 232586 272297 232592 272309
rect 243664 272297 243670 272309
rect 232586 272269 243670 272297
rect 232586 272257 232592 272269
rect 243664 272257 243670 272269
rect 243722 272257 243728 272309
rect 275152 272257 275158 272309
rect 275210 272297 275216 272309
rect 309328 272297 309334 272309
rect 275210 272269 309334 272297
rect 275210 272257 275216 272269
rect 309328 272257 309334 272269
rect 309386 272257 309392 272309
rect 309904 272257 309910 272309
rect 309962 272297 309968 272309
rect 395632 272297 395638 272309
rect 309962 272269 395638 272297
rect 309962 272257 309968 272269
rect 395632 272257 395638 272269
rect 395690 272257 395696 272309
rect 395920 272257 395926 272309
rect 395978 272297 395984 272309
rect 608368 272297 608374 272309
rect 395978 272269 608374 272297
rect 395978 272257 395984 272269
rect 608368 272257 608374 272269
rect 608426 272257 608432 272309
rect 84784 272183 84790 272235
rect 84842 272223 84848 272235
rect 86320 272223 86326 272235
rect 84842 272195 86326 272223
rect 84842 272183 84848 272195
rect 86320 272183 86326 272195
rect 86378 272183 86384 272235
rect 104848 272183 104854 272235
rect 104906 272223 104912 272235
rect 106480 272223 106486 272235
rect 104906 272195 106486 272223
rect 104906 272183 104912 272195
rect 106480 272183 106486 272195
rect 106538 272183 106544 272235
rect 195664 272223 195670 272235
rect 175666 272195 195670 272223
rect 76528 272109 76534 272161
rect 76586 272149 76592 272161
rect 175666 272149 175694 272195
rect 195664 272183 195670 272195
rect 195722 272183 195728 272235
rect 198256 272183 198262 272235
rect 198314 272223 198320 272235
rect 224368 272223 224374 272235
rect 198314 272195 224374 272223
rect 198314 272183 198320 272195
rect 224368 272183 224374 272195
rect 224426 272183 224432 272235
rect 227824 272183 227830 272235
rect 227882 272223 227888 272235
rect 242128 272223 242134 272235
rect 227882 272195 242134 272223
rect 227882 272183 227888 272195
rect 242128 272183 242134 272195
rect 242186 272183 242192 272235
rect 273424 272183 273430 272235
rect 273482 272223 273488 272235
rect 305776 272223 305782 272235
rect 273482 272195 305782 272223
rect 273482 272183 273488 272195
rect 305776 272183 305782 272195
rect 305834 272183 305840 272235
rect 312784 272183 312790 272235
rect 312842 272223 312848 272235
rect 402736 272223 402742 272235
rect 312842 272195 402742 272223
rect 312842 272183 312848 272195
rect 402736 272183 402742 272195
rect 402794 272183 402800 272235
rect 406096 272183 406102 272235
rect 406154 272223 406160 272235
rect 413392 272223 413398 272235
rect 406154 272195 413398 272223
rect 406154 272183 406160 272195
rect 413392 272183 413398 272195
rect 413450 272183 413456 272235
rect 413488 272183 413494 272235
rect 413546 272223 413552 272235
rect 636784 272223 636790 272235
rect 413546 272195 636790 272223
rect 413546 272183 413552 272195
rect 636784 272183 636790 272195
rect 636842 272183 636848 272235
rect 76586 272121 175694 272149
rect 76586 272109 76592 272121
rect 194704 272109 194710 272161
rect 194762 272149 194768 272161
rect 224464 272149 224470 272161
rect 194762 272121 224470 272149
rect 194762 272109 194768 272121
rect 224464 272109 224470 272121
rect 224522 272109 224528 272161
rect 228976 272109 228982 272161
rect 229034 272149 229040 272161
rect 242416 272149 242422 272161
rect 229034 272121 242422 272149
rect 229034 272109 229040 272121
rect 242416 272109 242422 272121
rect 242474 272109 242480 272161
rect 276304 272109 276310 272161
rect 276362 272149 276368 272161
rect 312880 272149 312886 272161
rect 276362 272121 312886 272149
rect 276362 272109 276368 272121
rect 312880 272109 312886 272121
rect 312938 272109 312944 272161
rect 315472 272109 315478 272161
rect 315530 272149 315536 272161
rect 409840 272149 409846 272161
rect 315530 272121 409846 272149
rect 315530 272109 315536 272121
rect 409840 272109 409846 272121
rect 409898 272109 409904 272161
rect 411856 272109 411862 272161
rect 411914 272149 411920 272161
rect 643888 272149 643894 272161
rect 411914 272121 643894 272149
rect 411914 272109 411920 272121
rect 643888 272109 643894 272121
rect 643946 272109 643952 272161
rect 167536 272035 167542 272087
rect 167594 272075 167600 272087
rect 210640 272075 210646 272087
rect 167594 272047 210646 272075
rect 167594 272035 167600 272047
rect 210640 272035 210646 272047
rect 210698 272035 210704 272087
rect 298000 272035 298006 272087
rect 298058 272075 298064 272087
rect 327088 272075 327094 272087
rect 298058 272047 327094 272075
rect 298058 272035 298064 272047
rect 327088 272035 327094 272047
rect 327146 272035 327152 272087
rect 347248 272035 347254 272087
rect 347306 272075 347312 272087
rect 487792 272075 487798 272087
rect 347306 272047 487798 272075
rect 347306 272035 347312 272047
rect 487792 272035 487798 272047
rect 487850 272035 487856 272087
rect 174640 271961 174646 272013
rect 174698 272001 174704 272013
rect 210544 272001 210550 272013
rect 174698 271973 210550 272001
rect 174698 271961 174704 271973
rect 210544 271961 210550 271973
rect 210602 271961 210608 272013
rect 231376 271961 231382 272013
rect 231434 272001 231440 272013
rect 243088 272001 243094 272013
rect 231434 271973 243094 272001
rect 231434 271961 231440 271973
rect 243088 271961 243094 271973
rect 243146 271961 243152 272013
rect 299440 271961 299446 272013
rect 299498 272001 299504 272013
rect 328240 272001 328246 272013
rect 299498 271973 328246 272001
rect 299498 271961 299504 271973
rect 328240 271961 328246 271973
rect 328298 271961 328304 272013
rect 346480 271961 346486 272013
rect 346538 272001 346544 272013
rect 486640 272001 486646 272013
rect 346538 271973 486646 272001
rect 346538 271961 346544 271973
rect 486640 271961 486646 271973
rect 486698 271961 486704 272013
rect 159280 271887 159286 271939
rect 159338 271927 159344 271939
rect 192976 271927 192982 271939
rect 159338 271899 192982 271927
rect 159338 271887 159344 271899
rect 192976 271887 192982 271899
rect 193034 271887 193040 271939
rect 195856 271887 195862 271939
rect 195914 271927 195920 271939
rect 221680 271927 221686 271939
rect 195914 271899 221686 271927
rect 195914 271887 195920 271899
rect 221680 271887 221686 271899
rect 221738 271887 221744 271939
rect 233680 271887 233686 271939
rect 233738 271927 233744 271939
rect 244048 271927 244054 271939
rect 233738 271899 244054 271927
rect 233738 271887 233744 271899
rect 244048 271887 244054 271899
rect 244106 271887 244112 271939
rect 272272 271887 272278 271939
rect 272330 271927 272336 271939
rect 301936 271927 301942 271939
rect 272330 271899 301942 271927
rect 272330 271887 272336 271899
rect 301936 271887 301942 271899
rect 301994 271887 302000 271939
rect 302320 271887 302326 271939
rect 302378 271927 302384 271939
rect 324688 271927 324694 271939
rect 302378 271899 324694 271927
rect 302378 271887 302384 271899
rect 324688 271887 324694 271899
rect 324746 271887 324752 271939
rect 344080 271887 344086 271939
rect 344138 271927 344144 271939
rect 480688 271927 480694 271939
rect 344138 271899 480694 271927
rect 344138 271887 344144 271899
rect 480688 271887 480694 271899
rect 480746 271887 480752 271939
rect 191152 271813 191158 271865
rect 191210 271853 191216 271865
rect 227152 271853 227158 271865
rect 191210 271825 227158 271853
rect 191210 271813 191216 271825
rect 227152 271813 227158 271825
rect 227210 271813 227216 271865
rect 341488 271813 341494 271865
rect 341546 271853 341552 271865
rect 473680 271853 473686 271865
rect 341546 271825 473686 271853
rect 341546 271813 341552 271825
rect 473680 271813 473686 271825
rect 473738 271813 473744 271865
rect 101296 271739 101302 271791
rect 101354 271779 101360 271791
rect 103600 271779 103606 271791
rect 101354 271751 103606 271779
rect 101354 271739 101360 271751
rect 103600 271739 103606 271751
rect 103658 271739 103664 271791
rect 147376 271739 147382 271791
rect 147434 271779 147440 271791
rect 149680 271779 149686 271791
rect 147434 271751 149686 271779
rect 147434 271739 147440 271751
rect 149680 271739 149686 271751
rect 149738 271739 149744 271791
rect 192304 271739 192310 271791
rect 192362 271779 192368 271791
rect 224560 271779 224566 271791
rect 192362 271751 224566 271779
rect 192362 271739 192368 271751
rect 224560 271739 224566 271751
rect 224618 271739 224624 271791
rect 338608 271739 338614 271791
rect 338666 271779 338672 271791
rect 466576 271779 466582 271791
rect 338666 271751 466582 271779
rect 338666 271739 338672 271751
rect 466576 271739 466582 271751
rect 466634 271739 466640 271791
rect 166288 271665 166294 271717
rect 166346 271705 166352 271717
rect 198640 271705 198646 271717
rect 166346 271677 198646 271705
rect 166346 271665 166352 271677
rect 198640 271665 198646 271677
rect 198698 271665 198704 271717
rect 199408 271665 199414 271717
rect 199466 271705 199472 271717
rect 221584 271705 221590 271717
rect 199466 271677 221590 271705
rect 199466 271665 199472 271677
rect 221584 271665 221590 271677
rect 221642 271665 221648 271717
rect 335440 271665 335446 271717
rect 335498 271705 335504 271717
rect 459472 271705 459478 271717
rect 335498 271677 459478 271705
rect 335498 271665 335504 271677
rect 459472 271665 459478 271677
rect 459530 271665 459536 271717
rect 75280 271591 75286 271643
rect 75338 271631 75344 271643
rect 77680 271631 77686 271643
rect 75338 271603 77686 271631
rect 75338 271591 75344 271603
rect 77680 271591 77686 271603
rect 77738 271591 77744 271643
rect 129712 271591 129718 271643
rect 129770 271631 129776 271643
rect 132400 271631 132406 271643
rect 129770 271603 132406 271631
rect 129770 271591 129776 271603
rect 132400 271591 132406 271603
rect 132458 271591 132464 271643
rect 181744 271591 181750 271643
rect 181802 271631 181808 271643
rect 210448 271631 210454 271643
rect 181802 271603 210454 271631
rect 181802 271591 181808 271603
rect 210448 271591 210454 271603
rect 210506 271591 210512 271643
rect 332560 271591 332566 271643
rect 332618 271631 332624 271643
rect 452368 271631 452374 271643
rect 332618 271603 452374 271631
rect 332618 271591 332624 271603
rect 452368 271591 452374 271603
rect 452426 271591 452432 271643
rect 89488 271517 89494 271569
rect 89546 271557 89552 271569
rect 92080 271557 92086 271569
rect 89546 271529 92086 271557
rect 89546 271517 89552 271529
rect 92080 271517 92086 271529
rect 92138 271517 92144 271569
rect 150928 271517 150934 271569
rect 150986 271557 150992 271569
rect 152368 271557 152374 271569
rect 150986 271529 152374 271557
rect 150986 271517 150992 271529
rect 152368 271517 152374 271529
rect 152426 271517 152432 271569
rect 180496 271517 180502 271569
rect 180554 271557 180560 271569
rect 205168 271557 205174 271569
rect 180554 271529 205174 271557
rect 180554 271517 180560 271529
rect 205168 271517 205174 271529
rect 205226 271517 205232 271569
rect 329968 271517 329974 271569
rect 330026 271557 330032 271569
rect 445264 271557 445270 271569
rect 330026 271529 445270 271557
rect 330026 271517 330032 271529
rect 445264 271517 445270 271529
rect 445322 271517 445328 271569
rect 173392 271443 173398 271495
rect 173450 271483 173456 271495
rect 201520 271483 201526 271495
rect 173450 271455 201526 271483
rect 173450 271443 173456 271455
rect 201520 271443 201526 271455
rect 201578 271443 201584 271495
rect 201808 271443 201814 271495
rect 201866 271483 201872 271495
rect 223696 271483 223702 271495
rect 201866 271455 223702 271483
rect 201866 271443 201872 271455
rect 223696 271443 223702 271455
rect 223754 271443 223760 271495
rect 326896 271443 326902 271495
rect 326954 271483 326960 271495
rect 438160 271483 438166 271495
rect 326954 271455 438166 271483
rect 326954 271443 326960 271455
rect 438160 271443 438166 271455
rect 438218 271443 438224 271495
rect 185200 271369 185206 271421
rect 185258 271409 185264 271421
rect 210352 271409 210358 271421
rect 185258 271381 210358 271409
rect 185258 271369 185264 271381
rect 210352 271369 210358 271381
rect 210410 271369 210416 271421
rect 334096 271369 334102 271421
rect 334154 271409 334160 271421
rect 337744 271409 337750 271421
rect 334154 271381 337750 271409
rect 334154 271369 334160 271381
rect 337744 271369 337750 271381
rect 337802 271369 337808 271421
rect 346960 271369 346966 271421
rect 347018 271409 347024 271421
rect 431056 271409 431062 271421
rect 347018 271381 431062 271409
rect 347018 271369 347024 271381
rect 431056 271369 431062 271381
rect 431114 271369 431120 271421
rect 184048 271295 184054 271347
rect 184106 271335 184112 271347
rect 205936 271335 205942 271347
rect 184106 271307 205942 271335
rect 184106 271295 184112 271307
rect 205936 271295 205942 271307
rect 205994 271295 206000 271347
rect 321424 271295 321430 271347
rect 321482 271335 321488 271347
rect 423952 271335 423958 271347
rect 321482 271307 423958 271335
rect 321482 271295 321488 271307
rect 423952 271295 423958 271307
rect 424010 271295 424016 271347
rect 161584 271221 161590 271273
rect 161642 271261 161648 271273
rect 163888 271261 163894 271273
rect 161642 271233 163894 271261
rect 161642 271221 161648 271233
rect 163888 271221 163894 271233
rect 163946 271221 163952 271273
rect 188752 271221 188758 271273
rect 188810 271261 188816 271273
rect 210256 271261 210262 271273
rect 188810 271233 210262 271261
rect 188810 271221 188816 271233
rect 210256 271221 210262 271233
rect 210314 271221 210320 271273
rect 237232 271221 237238 271273
rect 237290 271261 237296 271273
rect 245584 271261 245590 271273
rect 237290 271233 245590 271261
rect 237290 271221 237296 271233
rect 245584 271221 245590 271233
rect 245642 271221 245648 271273
rect 318352 271221 318358 271273
rect 318410 271261 318416 271273
rect 416944 271261 416950 271273
rect 318410 271233 416950 271261
rect 318410 271221 318416 271233
rect 416944 271221 416950 271233
rect 417002 271221 417008 271273
rect 175792 271147 175798 271199
rect 175850 271187 175856 271199
rect 178288 271187 178294 271199
rect 175850 271159 178294 271187
rect 175850 271147 175856 271159
rect 178288 271147 178294 271159
rect 178346 271147 178352 271199
rect 187600 271147 187606 271199
rect 187658 271187 187664 271199
rect 205840 271187 205846 271199
rect 187658 271159 205846 271187
rect 187658 271147 187664 271159
rect 205840 271147 205846 271159
rect 205898 271147 205904 271199
rect 238480 271147 238486 271199
rect 238538 271187 238544 271199
rect 246064 271187 246070 271199
rect 238538 271159 246070 271187
rect 238538 271147 238544 271159
rect 246064 271147 246070 271159
rect 246122 271147 246128 271199
rect 324016 271147 324022 271199
rect 324074 271187 324080 271199
rect 346960 271187 346966 271199
rect 324074 271159 346966 271187
rect 324074 271147 324080 271159
rect 346960 271147 346966 271159
rect 347018 271147 347024 271199
rect 357904 271147 357910 271199
rect 357962 271187 357968 271199
rect 375184 271187 375190 271199
rect 357962 271159 375190 271187
rect 357962 271147 357968 271159
rect 375184 271147 375190 271159
rect 375242 271147 375248 271199
rect 409840 271147 409846 271199
rect 409898 271187 409904 271199
rect 413488 271187 413494 271199
rect 409898 271159 413494 271187
rect 409898 271147 409904 271159
rect 413488 271147 413494 271159
rect 413546 271147 413552 271199
rect 85936 271073 85942 271125
rect 85994 271113 86000 271125
rect 198544 271113 198550 271125
rect 85994 271085 198550 271113
rect 85994 271073 86000 271085
rect 198544 271073 198550 271085
rect 198602 271073 198608 271125
rect 205360 271073 205366 271125
rect 205418 271113 205424 271125
rect 232624 271113 232630 271125
rect 205418 271085 232630 271113
rect 205418 271073 205424 271085
rect 232624 271073 232630 271085
rect 232682 271073 232688 271125
rect 240784 271073 240790 271125
rect 240842 271113 240848 271125
rect 247216 271113 247222 271125
rect 240842 271085 247222 271113
rect 240842 271073 240848 271085
rect 247216 271073 247222 271085
rect 247274 271073 247280 271125
rect 221872 270999 221878 271051
rect 221930 271039 221936 271051
rect 239344 271039 239350 271051
rect 221930 271011 239350 271039
rect 221930 270999 221936 271011
rect 239344 270999 239350 271011
rect 239402 270999 239408 271051
rect 239536 270999 239542 271051
rect 239594 271039 239600 271051
rect 241264 271039 241270 271051
rect 239594 271011 241270 271039
rect 239594 270999 239600 271011
rect 241264 270999 241270 271011
rect 241322 270999 241328 271051
rect 241936 270999 241942 271051
rect 241994 271039 242000 271051
rect 247696 271039 247702 271051
rect 241994 271011 247702 271039
rect 241994 270999 242000 271011
rect 247696 270999 247702 271011
rect 247754 270999 247760 271051
rect 342736 270999 342742 271051
rect 342794 271039 342800 271051
rect 348304 271039 348310 271051
rect 342794 271011 348310 271039
rect 342794 270999 342800 271011
rect 348304 270999 348310 271011
rect 348362 270999 348368 271051
rect 223024 270925 223030 270977
rect 223082 270965 223088 270977
rect 240016 270965 240022 270977
rect 223082 270937 240022 270965
rect 223082 270925 223088 270937
rect 240016 270925 240022 270937
rect 240074 270925 240080 270977
rect 243184 270925 243190 270977
rect 243242 270965 243248 270977
rect 247984 270965 247990 270977
rect 243242 270937 247990 270965
rect 243242 270925 243248 270937
rect 247984 270925 247990 270937
rect 248042 270925 248048 270977
rect 224272 270851 224278 270903
rect 224330 270891 224336 270903
rect 240496 270891 240502 270903
rect 224330 270863 240502 270891
rect 224330 270851 224336 270863
rect 240496 270851 240502 270863
rect 240554 270851 240560 270903
rect 244336 270851 244342 270903
rect 244394 270891 244400 270903
rect 248656 270891 248662 270903
rect 244394 270863 248662 270891
rect 244394 270851 244400 270863
rect 248656 270851 248662 270863
rect 248714 270851 248720 270903
rect 225424 270777 225430 270829
rect 225482 270817 225488 270829
rect 241072 270817 241078 270829
rect 225482 270789 241078 270817
rect 225482 270777 225488 270789
rect 241072 270777 241078 270789
rect 241130 270777 241136 270829
rect 245488 270777 245494 270829
rect 245546 270817 245552 270829
rect 249136 270817 249142 270829
rect 245546 270789 249142 270817
rect 245546 270777 245552 270789
rect 249136 270777 249142 270789
rect 249194 270777 249200 270829
rect 94192 270703 94198 270755
rect 94250 270743 94256 270755
rect 94960 270743 94966 270755
rect 94250 270715 94966 270743
rect 94250 270703 94256 270715
rect 94960 270703 94966 270715
rect 95018 270703 95024 270755
rect 115504 270703 115510 270755
rect 115562 270743 115568 270755
rect 118000 270743 118006 270755
rect 115562 270715 118006 270743
rect 115562 270703 115568 270715
rect 118000 270703 118006 270715
rect 118058 270703 118064 270755
rect 119056 270703 119062 270755
rect 119114 270743 119120 270755
rect 120880 270743 120886 270755
rect 119114 270715 120886 270743
rect 119114 270703 119120 270715
rect 120880 270703 120886 270715
rect 120938 270703 120944 270755
rect 133264 270703 133270 270755
rect 133322 270743 133328 270755
rect 135280 270743 135286 270755
rect 133322 270715 135286 270743
rect 133322 270703 133328 270715
rect 135280 270703 135286 270715
rect 135338 270703 135344 270755
rect 136816 270703 136822 270755
rect 136874 270743 136880 270755
rect 138160 270743 138166 270755
rect 136874 270715 138166 270743
rect 136874 270703 136880 270715
rect 138160 270703 138166 270715
rect 138218 270703 138224 270755
rect 154480 270703 154486 270755
rect 154538 270743 154544 270755
rect 155440 270743 155446 270755
rect 154538 270715 155446 270743
rect 154538 270703 154544 270715
rect 155440 270703 155446 270715
rect 155498 270703 155504 270755
rect 165136 270703 165142 270755
rect 165194 270743 165200 270755
rect 166960 270743 166966 270755
rect 165194 270715 166966 270743
rect 165194 270703 165200 270715
rect 166960 270703 166966 270715
rect 167018 270703 167024 270755
rect 168688 270703 168694 270755
rect 168746 270743 168752 270755
rect 169840 270743 169846 270755
rect 168746 270715 169846 270743
rect 168746 270703 168752 270715
rect 169840 270703 169846 270715
rect 169898 270703 169904 270755
rect 179344 270703 179350 270755
rect 179402 270743 179408 270755
rect 181360 270743 181366 270755
rect 179402 270715 181366 270743
rect 179402 270703 179408 270715
rect 181360 270703 181366 270715
rect 181418 270703 181424 270755
rect 182896 270703 182902 270755
rect 182954 270743 182960 270755
rect 184240 270743 184246 270755
rect 182954 270715 184246 270743
rect 182954 270703 182960 270715
rect 184240 270703 184246 270715
rect 184298 270703 184304 270755
rect 185488 270703 185494 270755
rect 185546 270743 185552 270755
rect 186448 270743 186454 270755
rect 185546 270715 186454 270743
rect 185546 270703 185552 270715
rect 186448 270703 186454 270715
rect 186506 270703 186512 270755
rect 226576 270703 226582 270755
rect 226634 270743 226640 270755
rect 239536 270743 239542 270755
rect 226634 270715 239542 270743
rect 226634 270703 226640 270715
rect 239536 270703 239542 270715
rect 239594 270703 239600 270755
rect 239632 270703 239638 270755
rect 239690 270743 239696 270755
rect 246448 270743 246454 270755
rect 239690 270715 246454 270743
rect 239690 270703 239696 270715
rect 246448 270703 246454 270715
rect 246506 270703 246512 270755
rect 246736 270703 246742 270755
rect 246794 270743 246800 270755
rect 249616 270743 249622 270755
rect 246794 270715 249622 270743
rect 246794 270703 246800 270715
rect 249616 270703 249622 270715
rect 249674 270703 249680 270755
rect 351376 270703 351382 270755
rect 351434 270743 351440 270755
rect 355408 270743 355414 270755
rect 351434 270715 355414 270743
rect 351434 270703 351440 270715
rect 355408 270703 355414 270715
rect 355466 270703 355472 270755
rect 146224 270629 146230 270681
rect 146282 270669 146288 270681
rect 214960 270669 214966 270681
rect 146282 270641 214966 270669
rect 146282 270629 146288 270641
rect 214960 270629 214966 270641
rect 215018 270629 215024 270681
rect 280144 270629 280150 270681
rect 280202 270669 280208 270681
rect 322384 270669 322390 270681
rect 280202 270641 322390 270669
rect 280202 270629 280208 270641
rect 322384 270629 322390 270641
rect 322442 270629 322448 270681
rect 350704 270629 350710 270681
rect 350762 270669 350768 270681
rect 497296 270669 497302 270681
rect 350762 270641 497302 270669
rect 350762 270629 350768 270641
rect 497296 270629 497302 270641
rect 497354 270629 497360 270681
rect 137968 270555 137974 270607
rect 138026 270595 138032 270607
rect 212656 270595 212662 270607
rect 138026 270567 212662 270595
rect 138026 270555 138032 270567
rect 212656 270555 212662 270567
rect 212714 270555 212720 270607
rect 280624 270555 280630 270607
rect 280682 270595 280688 270607
rect 323536 270595 323542 270607
rect 280682 270567 323542 270595
rect 280682 270555 280688 270567
rect 323536 270555 323542 270567
rect 323594 270555 323600 270607
rect 351280 270555 351286 270607
rect 351338 270595 351344 270607
rect 498448 270595 498454 270607
rect 351338 270567 498454 270595
rect 351338 270555 351344 270567
rect 498448 270555 498454 270567
rect 498506 270555 498512 270607
rect 141520 270481 141526 270533
rect 141578 270521 141584 270533
rect 213808 270521 213814 270533
rect 141578 270493 213814 270521
rect 141578 270481 141584 270493
rect 213808 270481 213814 270493
rect 213866 270481 213872 270533
rect 264688 270481 264694 270533
rect 264746 270521 264752 270533
rect 283312 270521 283318 270533
rect 264746 270493 283318 270521
rect 264746 270481 264752 270493
rect 283312 270481 283318 270493
rect 283370 270481 283376 270533
rect 319984 270521 319990 270533
rect 283426 270493 319990 270521
rect 134416 270407 134422 270459
rect 134474 270447 134480 270459
rect 211888 270447 211894 270459
rect 134474 270419 211894 270447
rect 134474 270407 134480 270419
rect 211888 270407 211894 270419
rect 211946 270407 211952 270459
rect 253936 270407 253942 270459
rect 253994 270447 254000 270459
rect 257296 270447 257302 270459
rect 253994 270419 257302 270447
rect 253994 270407 254000 270419
rect 257296 270407 257302 270419
rect 257354 270407 257360 270459
rect 264880 270407 264886 270459
rect 264938 270447 264944 270459
rect 276400 270447 276406 270459
rect 264938 270419 276406 270447
rect 264938 270407 264944 270419
rect 276400 270407 276406 270419
rect 276458 270407 276464 270459
rect 279280 270407 279286 270459
rect 279338 270447 279344 270459
rect 283426 270447 283454 270493
rect 319984 270481 319990 270493
rect 320042 270481 320048 270533
rect 353680 270481 353686 270533
rect 353738 270521 353744 270533
rect 504400 270521 504406 270533
rect 353738 270493 504406 270521
rect 353738 270481 353744 270493
rect 504400 270481 504406 270493
rect 504458 270481 504464 270533
rect 279338 270419 283454 270447
rect 279338 270407 279344 270419
rect 283696 270407 283702 270459
rect 283754 270447 283760 270459
rect 330640 270447 330646 270459
rect 283754 270419 330646 270447
rect 283754 270407 283760 270419
rect 330640 270407 330646 270419
rect 330698 270407 330704 270459
rect 354064 270407 354070 270459
rect 354122 270447 354128 270459
rect 505552 270447 505558 270459
rect 354122 270419 505558 270447
rect 354122 270407 354128 270419
rect 505552 270407 505558 270419
rect 505610 270407 505616 270459
rect 121456 270333 121462 270385
rect 121514 270373 121520 270385
rect 208336 270373 208342 270385
rect 121514 270345 208342 270373
rect 121514 270333 121520 270345
rect 208336 270333 208342 270345
rect 208394 270333 208400 270385
rect 262480 270333 262486 270385
rect 262538 270373 262544 270385
rect 278608 270373 278614 270385
rect 262538 270345 278614 270373
rect 262538 270333 262544 270345
rect 278608 270333 278614 270345
rect 278666 270333 278672 270385
rect 284176 270333 284182 270385
rect 284234 270373 284240 270385
rect 331792 270373 331798 270385
rect 284234 270345 331798 270373
rect 284234 270333 284240 270345
rect 331792 270333 331798 270345
rect 331850 270333 331856 270385
rect 356752 270333 356758 270385
rect 356810 270373 356816 270385
rect 511504 270373 511510 270385
rect 356810 270345 511510 270373
rect 356810 270333 356816 270345
rect 511504 270333 511510 270345
rect 511562 270333 511568 270385
rect 117904 270259 117910 270311
rect 117962 270299 117968 270311
rect 207568 270299 207574 270311
rect 117962 270271 207574 270299
rect 117962 270259 117968 270271
rect 207568 270259 207574 270271
rect 207626 270259 207632 270311
rect 255280 270259 255286 270311
rect 255338 270299 255344 270311
rect 260848 270299 260854 270311
rect 255338 270271 260854 270299
rect 255338 270259 255344 270271
rect 260848 270259 260854 270271
rect 260906 270259 260912 270311
rect 266032 270259 266038 270311
rect 266090 270299 266096 270311
rect 286864 270299 286870 270311
rect 266090 270271 286870 270299
rect 266090 270259 266096 270271
rect 286864 270259 286870 270271
rect 286922 270259 286928 270311
rect 334096 270299 334102 270311
rect 286978 270271 334102 270299
rect 114352 270185 114358 270237
rect 114410 270225 114416 270237
rect 206416 270225 206422 270237
rect 114410 270197 206422 270225
rect 114410 270185 114416 270197
rect 206416 270185 206422 270197
rect 206474 270185 206480 270237
rect 210544 270185 210550 270237
rect 210602 270225 210608 270237
rect 222832 270225 222838 270237
rect 210602 270197 222838 270225
rect 210602 270185 210608 270197
rect 222832 270185 222838 270197
rect 222890 270185 222896 270237
rect 265360 270185 265366 270237
rect 265418 270225 265424 270237
rect 265418 270197 276350 270225
rect 265418 270185 265424 270197
rect 109552 270111 109558 270163
rect 109610 270151 109616 270163
rect 205264 270151 205270 270163
rect 109610 270123 205270 270151
rect 109610 270111 109616 270123
rect 205264 270111 205270 270123
rect 205322 270111 205328 270163
rect 210256 270111 210262 270163
rect 210314 270151 210320 270163
rect 226672 270151 226678 270163
rect 210314 270123 226678 270151
rect 210314 270111 210320 270123
rect 226672 270111 226678 270123
rect 226730 270111 226736 270163
rect 266512 270111 266518 270163
rect 266570 270151 266576 270163
rect 276322 270151 276350 270197
rect 276400 270185 276406 270237
rect 276458 270225 276464 270237
rect 284560 270225 284566 270237
rect 276458 270197 284566 270225
rect 276458 270185 276464 270197
rect 284560 270185 284566 270197
rect 284618 270185 284624 270237
rect 286288 270185 286294 270237
rect 286346 270225 286352 270237
rect 286978 270225 287006 270271
rect 334096 270259 334102 270271
rect 334154 270259 334160 270311
rect 356944 270259 356950 270311
rect 357002 270299 357008 270311
rect 512656 270299 512662 270311
rect 357002 270271 512662 270299
rect 357002 270259 357008 270271
rect 512656 270259 512662 270271
rect 512714 270259 512720 270311
rect 286346 270197 287006 270225
rect 286346 270185 286352 270197
rect 288496 270185 288502 270237
rect 288554 270225 288560 270237
rect 342448 270225 342454 270237
rect 288554 270197 342454 270225
rect 288554 270185 288560 270197
rect 342448 270185 342454 270197
rect 342506 270185 342512 270237
rect 359824 270185 359830 270237
rect 359882 270225 359888 270237
rect 519760 270225 519766 270237
rect 359882 270197 519766 270225
rect 359882 270185 359888 270197
rect 519760 270185 519766 270197
rect 519818 270185 519824 270237
rect 285712 270151 285718 270163
rect 266570 270123 276254 270151
rect 276322 270123 285718 270151
rect 266570 270111 266576 270123
rect 102544 270037 102550 270089
rect 102602 270077 102608 270089
rect 203344 270077 203350 270089
rect 102602 270049 203350 270077
rect 102602 270037 102608 270049
rect 203344 270037 203350 270049
rect 203402 270037 203408 270089
rect 210352 270037 210358 270089
rect 210410 270077 210416 270089
rect 225520 270077 225526 270089
rect 210410 270049 225526 270077
rect 210410 270037 210416 270049
rect 225520 270037 225526 270049
rect 225578 270037 225584 270089
rect 267280 270037 267286 270089
rect 267338 270077 267344 270089
rect 276226 270077 276254 270123
rect 285712 270111 285718 270123
rect 285770 270111 285776 270163
rect 287920 270111 287926 270163
rect 287978 270151 287984 270163
rect 337936 270151 337942 270163
rect 287978 270123 337942 270151
rect 287978 270111 287984 270123
rect 337936 270111 337942 270123
rect 337994 270111 338000 270163
rect 359344 270111 359350 270163
rect 359402 270151 359408 270163
rect 518512 270151 518518 270163
rect 359402 270123 518518 270151
rect 359402 270111 359408 270123
rect 518512 270111 518518 270123
rect 518570 270111 518576 270163
rect 288016 270077 288022 270089
rect 267338 270049 272126 270077
rect 276226 270049 288022 270077
rect 267338 270037 267344 270049
rect 107248 269963 107254 270015
rect 107306 270003 107312 270015
rect 204688 270003 204694 270015
rect 107306 269975 204694 270003
rect 107306 269963 107312 269975
rect 204688 269963 204694 269975
rect 204746 269963 204752 270015
rect 210448 269963 210454 270015
rect 210506 270003 210512 270015
rect 224752 270003 224758 270015
rect 210506 269975 224758 270003
rect 210506 269963 210512 269975
rect 224752 269963 224758 269975
rect 224810 269963 224816 270015
rect 267088 269963 267094 270015
rect 267146 270003 267152 270015
rect 272098 270003 272126 270049
rect 288016 270037 288022 270049
rect 288074 270037 288080 270089
rect 290608 270037 290614 270089
rect 290666 270077 290672 270089
rect 342736 270077 342742 270089
rect 290666 270049 342742 270077
rect 290666 270037 290672 270049
rect 342736 270037 342742 270049
rect 342794 270037 342800 270089
rect 362224 270037 362230 270089
rect 362282 270077 362288 270089
rect 525616 270077 525622 270089
rect 362282 270049 525622 270077
rect 362282 270037 362288 270049
rect 525616 270037 525622 270049
rect 525674 270037 525680 270089
rect 290416 270003 290422 270015
rect 267146 269975 272030 270003
rect 272098 269975 290422 270003
rect 267146 269963 267152 269975
rect 100144 269889 100150 269941
rect 100202 269929 100208 269941
rect 202864 269929 202870 269941
rect 100202 269901 202870 269929
rect 100202 269889 100208 269901
rect 202864 269889 202870 269901
rect 202922 269889 202928 269941
rect 205168 269889 205174 269941
rect 205226 269929 205232 269941
rect 224080 269929 224086 269941
rect 205226 269901 224086 269929
rect 205226 269889 205232 269901
rect 224080 269889 224086 269901
rect 224138 269889 224144 269941
rect 256240 269889 256246 269941
rect 256298 269929 256304 269941
rect 263248 269929 263254 269941
rect 256298 269901 263254 269929
rect 256298 269889 256304 269901
rect 263248 269889 263254 269901
rect 263306 269889 263312 269941
rect 267760 269889 267766 269941
rect 267818 269929 267824 269941
rect 272002 269929 272030 269975
rect 290416 269963 290422 269975
rect 290474 269963 290480 270015
rect 291088 269963 291094 270015
rect 291146 270003 291152 270015
rect 349552 270003 349558 270015
rect 291146 269975 349558 270003
rect 291146 269963 291152 269975
rect 349552 269963 349558 269975
rect 349610 269963 349616 270015
rect 362800 269963 362806 270015
rect 362858 270003 362864 270015
rect 526864 270003 526870 270015
rect 362858 269975 526870 270003
rect 362858 269963 362864 269975
rect 526864 269963 526870 269975
rect 526922 269963 526928 270015
rect 289264 269929 289270 269941
rect 267818 269901 271838 269929
rect 272002 269901 289270 269929
rect 267818 269889 267824 269901
rect 95440 269815 95446 269867
rect 95498 269855 95504 269867
rect 185680 269855 185686 269867
rect 95498 269827 185686 269855
rect 95498 269815 95504 269827
rect 185680 269815 185686 269827
rect 185738 269815 185744 269867
rect 205936 269815 205942 269867
rect 205994 269855 206000 269867
rect 225232 269855 225238 269867
rect 205994 269827 225238 269855
rect 205994 269815 206000 269827
rect 225232 269815 225238 269827
rect 225290 269815 225296 269867
rect 255760 269815 255766 269867
rect 255818 269855 255824 269867
rect 262096 269855 262102 269867
rect 255818 269827 262102 269855
rect 255818 269815 255824 269827
rect 262096 269815 262102 269827
rect 262154 269815 262160 269867
rect 269200 269815 269206 269867
rect 269258 269855 269264 269867
rect 271810 269855 271838 269901
rect 289264 269889 289270 269901
rect 289322 269889 289328 269941
rect 293968 269889 293974 269941
rect 294026 269929 294032 269941
rect 356656 269929 356662 269941
rect 294026 269901 356662 269929
rect 294026 269889 294032 269901
rect 356656 269889 356662 269901
rect 356714 269889 356720 269941
rect 365296 269889 365302 269941
rect 365354 269929 365360 269941
rect 532720 269929 532726 269941
rect 365354 269901 532726 269929
rect 365354 269889 365360 269901
rect 532720 269889 532726 269901
rect 532778 269889 532784 269941
rect 291568 269855 291574 269867
rect 269258 269827 271742 269855
rect 271810 269827 291574 269855
rect 269258 269815 269264 269827
rect 93040 269741 93046 269793
rect 93098 269781 93104 269793
rect 200944 269781 200950 269793
rect 93098 269753 200950 269781
rect 93098 269741 93104 269753
rect 200944 269741 200950 269753
rect 201002 269741 201008 269793
rect 205840 269741 205846 269793
rect 205898 269781 205904 269793
rect 226000 269781 226006 269793
rect 205898 269753 226006 269781
rect 205898 269741 205904 269753
rect 226000 269741 226006 269753
rect 226058 269741 226064 269793
rect 271714 269781 271742 269827
rect 291568 269815 291574 269827
rect 291626 269815 291632 269867
rect 293488 269815 293494 269867
rect 293546 269855 293552 269867
rect 351376 269855 351382 269867
rect 293546 269827 351382 269855
rect 293546 269815 293552 269827
rect 351376 269815 351382 269827
rect 351434 269815 351440 269867
rect 365680 269815 365686 269867
rect 365738 269855 365744 269867
rect 533872 269855 533878 269867
rect 365738 269827 533878 269855
rect 365738 269815 365744 269827
rect 533872 269815 533878 269827
rect 533930 269815 533936 269867
rect 295120 269781 295126 269793
rect 271714 269753 295126 269781
rect 295120 269741 295126 269753
rect 295178 269741 295184 269793
rect 297040 269741 297046 269793
rect 297098 269781 297104 269793
rect 363664 269781 363670 269793
rect 297098 269753 363670 269781
rect 297098 269741 297104 269753
rect 363664 269741 363670 269753
rect 363722 269741 363728 269793
rect 371248 269741 371254 269793
rect 371306 269781 371312 269793
rect 548080 269781 548086 269793
rect 371306 269753 548086 269781
rect 371306 269741 371312 269753
rect 548080 269741 548086 269753
rect 548138 269741 548144 269793
rect 90640 269667 90646 269719
rect 90698 269707 90704 269719
rect 199696 269707 199702 269719
rect 90698 269679 199702 269707
rect 90698 269667 90704 269679
rect 199696 269667 199702 269679
rect 199754 269667 199760 269719
rect 201520 269667 201526 269719
rect 201578 269707 201584 269719
rect 222352 269707 222358 269719
rect 201578 269679 222358 269707
rect 201578 269667 201584 269679
rect 222352 269667 222358 269679
rect 222410 269667 222416 269719
rect 259888 269667 259894 269719
rect 259946 269707 259952 269719
rect 271504 269707 271510 269719
rect 259946 269679 271510 269707
rect 259946 269667 259952 269679
rect 271504 269667 271510 269679
rect 271562 269667 271568 269719
rect 271600 269667 271606 269719
rect 271658 269707 271664 269719
rect 293776 269707 293782 269719
rect 271658 269679 293782 269707
rect 271658 269667 271664 269679
rect 293776 269667 293782 269679
rect 293834 269667 293840 269719
rect 299632 269667 299638 269719
rect 299690 269707 299696 269719
rect 370768 269707 370774 269719
rect 299690 269679 370774 269707
rect 299690 269667 299696 269679
rect 370768 269667 370774 269679
rect 370826 269667 370832 269719
rect 379888 269667 379894 269719
rect 379946 269707 379952 269719
rect 569392 269707 569398 269719
rect 379946 269679 569398 269707
rect 379946 269667 379952 269679
rect 569392 269667 569398 269679
rect 569450 269667 569456 269719
rect 83632 269593 83638 269645
rect 83690 269633 83696 269645
rect 198064 269633 198070 269645
rect 83690 269605 198070 269633
rect 83690 269593 83696 269605
rect 198064 269593 198070 269605
rect 198122 269593 198128 269645
rect 198640 269593 198646 269645
rect 198698 269633 198704 269645
rect 220528 269633 220534 269645
rect 198698 269605 220534 269633
rect 198698 269593 198704 269605
rect 220528 269593 220534 269605
rect 220586 269593 220592 269645
rect 249040 269593 249046 269645
rect 249098 269633 249104 269645
rect 250288 269633 250294 269645
rect 249098 269605 250294 269633
rect 249098 269593 249104 269605
rect 250288 269593 250294 269605
rect 250346 269593 250352 269645
rect 257680 269593 257686 269645
rect 257738 269633 257744 269645
rect 266800 269633 266806 269645
rect 257738 269605 266806 269633
rect 257738 269593 257744 269605
rect 266800 269593 266806 269605
rect 266858 269593 266864 269645
rect 269680 269593 269686 269645
rect 269738 269633 269744 269645
rect 296368 269633 296374 269645
rect 269738 269605 296374 269633
rect 269738 269593 269744 269605
rect 296368 269593 296374 269605
rect 296426 269593 296432 269645
rect 302608 269593 302614 269645
rect 302666 269633 302672 269645
rect 377872 269633 377878 269645
rect 302666 269605 377878 269633
rect 302666 269593 302672 269605
rect 377872 269593 377878 269605
rect 377930 269593 377936 269645
rect 384112 269593 384118 269645
rect 384170 269633 384176 269645
rect 580048 269633 580054 269645
rect 384170 269605 580054 269633
rect 384170 269593 384176 269605
rect 580048 269593 580054 269605
rect 580106 269593 580112 269645
rect 87184 269519 87190 269571
rect 87242 269559 87248 269571
rect 199024 269559 199030 269571
rect 87242 269531 199030 269559
rect 87242 269519 87248 269531
rect 199024 269519 199030 269531
rect 199082 269519 199088 269571
rect 206512 269519 206518 269571
rect 206570 269559 206576 269571
rect 233392 269559 233398 269571
rect 206570 269531 233398 269559
rect 206570 269519 206576 269531
rect 233392 269519 233398 269531
rect 233450 269519 233456 269571
rect 271504 269519 271510 269571
rect 271562 269559 271568 269571
rect 301072 269559 301078 269571
rect 271562 269531 301078 269559
rect 271562 269519 271568 269531
rect 301072 269519 301078 269531
rect 301130 269519 301136 269571
rect 305680 269519 305686 269571
rect 305738 269559 305744 269571
rect 384976 269559 384982 269571
rect 305738 269531 384982 269559
rect 305738 269519 305744 269531
rect 384976 269519 384982 269531
rect 385034 269519 385040 269571
rect 385360 269519 385366 269571
rect 385418 269559 385424 269571
rect 582352 269559 582358 269571
rect 385418 269531 582358 269559
rect 385418 269519 385424 269531
rect 582352 269519 582358 269531
rect 582410 269519 582416 269571
rect 81232 269445 81238 269497
rect 81290 269485 81296 269497
rect 196816 269485 196822 269497
rect 81290 269457 196822 269485
rect 81290 269445 81296 269457
rect 196816 269445 196822 269457
rect 196874 269445 196880 269497
rect 202960 269445 202966 269497
rect 203018 269485 203024 269497
rect 231952 269485 231958 269497
rect 203018 269457 231958 269485
rect 203018 269445 203024 269457
rect 231952 269445 231958 269457
rect 232010 269445 232016 269497
rect 260080 269445 260086 269497
rect 260138 269485 260144 269497
rect 272656 269485 272662 269497
rect 260138 269457 272662 269485
rect 260138 269445 260144 269457
rect 272656 269445 272662 269457
rect 272714 269445 272720 269497
rect 272944 269445 272950 269497
rect 273002 269485 273008 269497
rect 304624 269485 304630 269497
rect 273002 269457 304630 269485
rect 273002 269445 273008 269457
rect 304624 269445 304630 269457
rect 304682 269445 304688 269497
rect 308272 269445 308278 269497
rect 308330 269485 308336 269497
rect 392080 269485 392086 269497
rect 308330 269457 392086 269485
rect 308330 269445 308336 269457
rect 392080 269445 392086 269457
rect 392138 269445 392144 269497
rect 82384 269371 82390 269423
rect 82442 269411 82448 269423
rect 197392 269411 197398 269423
rect 82442 269383 197398 269411
rect 82442 269371 82448 269383
rect 197392 269371 197398 269383
rect 197450 269371 197456 269423
rect 204112 269371 204118 269423
rect 204170 269411 204176 269423
rect 232144 269411 232150 269423
rect 204170 269383 232150 269411
rect 204170 269371 204176 269383
rect 232144 269371 232150 269383
rect 232202 269371 232208 269423
rect 274672 269371 274678 269423
rect 274730 269411 274736 269423
rect 308176 269411 308182 269423
rect 274730 269383 308182 269411
rect 274730 269371 274736 269383
rect 308176 269371 308182 269383
rect 308234 269371 308240 269423
rect 311152 269371 311158 269423
rect 311210 269411 311216 269423
rect 399184 269411 399190 269423
rect 311210 269383 399190 269411
rect 311210 269371 311216 269383
rect 399184 269371 399190 269383
rect 399242 269371 399248 269423
rect 399952 269371 399958 269423
rect 400010 269411 400016 269423
rect 619024 269411 619030 269423
rect 400010 269383 619030 269411
rect 400010 269371 400016 269383
rect 619024 269371 619030 269383
rect 619082 269371 619088 269423
rect 74128 269297 74134 269349
rect 74186 269337 74192 269349
rect 194992 269337 194998 269349
rect 74186 269309 194998 269337
rect 74186 269297 74192 269309
rect 194992 269297 194998 269309
rect 195050 269297 195056 269349
rect 200656 269297 200662 269349
rect 200714 269337 200720 269349
rect 230992 269337 230998 269349
rect 200714 269309 230998 269337
rect 200714 269297 200720 269309
rect 230992 269297 230998 269309
rect 231050 269297 231056 269349
rect 258640 269297 258646 269349
rect 258698 269337 258704 269349
rect 269104 269337 269110 269349
rect 258698 269309 269110 269337
rect 258698 269297 258704 269309
rect 269104 269297 269110 269309
rect 269162 269297 269168 269349
rect 278896 269297 278902 269349
rect 278954 269337 278960 269349
rect 318832 269337 318838 269349
rect 278954 269309 318838 269337
rect 278954 269297 278960 269309
rect 318832 269297 318838 269309
rect 318890 269297 318896 269349
rect 319024 269297 319030 269349
rect 319082 269337 319088 269349
rect 406096 269337 406102 269349
rect 319082 269309 406102 269337
rect 319082 269297 319088 269309
rect 406096 269297 406102 269309
rect 406154 269297 406160 269349
rect 409648 269297 409654 269349
rect 409706 269337 409712 269349
rect 642640 269337 642646 269349
rect 409706 269309 642646 269337
rect 409706 269297 409712 269309
rect 642640 269297 642646 269309
rect 642698 269297 642704 269349
rect 67024 269223 67030 269275
rect 67082 269263 67088 269275
rect 192592 269263 192598 269275
rect 67082 269235 192598 269263
rect 67082 269223 67088 269235
rect 192592 269223 192598 269235
rect 192650 269223 192656 269275
rect 197104 269223 197110 269275
rect 197162 269263 197168 269275
rect 229552 269263 229558 269275
rect 197162 269235 229558 269263
rect 197162 269223 197168 269235
rect 229552 269223 229558 269235
rect 229610 269223 229616 269275
rect 257488 269223 257494 269275
rect 257546 269263 257552 269275
rect 265648 269263 265654 269275
rect 257546 269235 265654 269263
rect 257546 269223 257552 269235
rect 265648 269223 265654 269235
rect 265706 269223 265712 269275
rect 268624 269223 268630 269275
rect 268682 269263 268688 269275
rect 271600 269263 271606 269275
rect 268682 269235 271606 269263
rect 268682 269223 268688 269235
rect 271600 269223 271606 269235
rect 271658 269223 271664 269275
rect 275824 269223 275830 269275
rect 275882 269263 275888 269275
rect 311728 269263 311734 269275
rect 275882 269235 311734 269263
rect 275882 269223 275888 269235
rect 311728 269223 311734 269235
rect 311786 269223 311792 269275
rect 314224 269223 314230 269275
rect 314282 269263 314288 269275
rect 406288 269263 406294 269275
rect 314282 269235 406294 269263
rect 314282 269223 314288 269235
rect 406288 269223 406294 269235
rect 406346 269223 406352 269275
rect 408496 269223 408502 269275
rect 408554 269263 408560 269275
rect 640336 269263 640342 269275
rect 408554 269235 640342 269263
rect 408554 269223 408560 269235
rect 640336 269223 640342 269235
rect 640394 269223 640400 269275
rect 145072 269149 145078 269201
rect 145130 269189 145136 269201
rect 214480 269189 214486 269201
rect 145130 269161 214486 269189
rect 145130 269149 145136 269161
rect 214480 269149 214486 269161
rect 214538 269149 214544 269201
rect 262000 269149 262006 269201
rect 262058 269189 262064 269201
rect 277456 269189 277462 269201
rect 262058 269161 277462 269189
rect 262058 269149 262064 269161
rect 277456 269149 277462 269161
rect 277514 269149 277520 269201
rect 277552 269149 277558 269201
rect 277610 269189 277616 269201
rect 315280 269189 315286 269201
rect 277610 269161 315286 269189
rect 277610 269149 277616 269161
rect 315280 269149 315286 269161
rect 315338 269149 315344 269201
rect 348112 269149 348118 269201
rect 348170 269189 348176 269201
rect 490192 269189 490198 269201
rect 348170 269161 490198 269189
rect 348170 269149 348176 269161
rect 490192 269149 490198 269161
rect 490250 269149 490256 269201
rect 152176 269075 152182 269127
rect 152234 269115 152240 269127
rect 216688 269115 216694 269127
rect 152234 269087 216694 269115
rect 152234 269075 152240 269087
rect 216688 269075 216694 269087
rect 216746 269075 216752 269127
rect 253360 269075 253366 269127
rect 253418 269115 253424 269127
rect 256144 269115 256150 269127
rect 253418 269087 256150 269115
rect 253418 269075 253424 269087
rect 256144 269075 256150 269087
rect 256202 269075 256208 269127
rect 259408 269075 259414 269127
rect 259466 269115 259472 269127
rect 270352 269115 270358 269127
rect 259466 269087 270358 269115
rect 259466 269075 259472 269087
rect 270352 269075 270358 269087
rect 270410 269075 270416 269127
rect 295216 269075 295222 269127
rect 295274 269115 295280 269127
rect 305392 269115 305398 269127
rect 295274 269087 305398 269115
rect 295274 269075 295280 269087
rect 305392 269075 305398 269087
rect 305450 269075 305456 269127
rect 309232 269075 309238 269127
rect 309290 269115 309296 269127
rect 343600 269115 343606 269127
rect 309290 269087 343606 269115
rect 309290 269075 309296 269087
rect 343600 269075 343606 269087
rect 343658 269075 343664 269127
rect 348400 269075 348406 269127
rect 348458 269115 348464 269127
rect 491344 269115 491350 269127
rect 348458 269087 491350 269115
rect 348458 269075 348464 269087
rect 491344 269075 491350 269087
rect 491402 269075 491408 269127
rect 149776 269001 149782 269053
rect 149834 269041 149840 269053
rect 216208 269041 216214 269053
rect 149834 269013 216214 269041
rect 149834 269001 149840 269013
rect 216208 269001 216214 269013
rect 216266 269001 216272 269053
rect 261808 269001 261814 269053
rect 261866 269041 261872 269053
rect 276208 269041 276214 269053
rect 261866 269013 276214 269041
rect 261866 269001 261872 269013
rect 276208 269001 276214 269013
rect 276266 269001 276272 269053
rect 281296 269001 281302 269053
rect 281354 269041 281360 269053
rect 302320 269041 302326 269053
rect 281354 269013 302326 269041
rect 281354 269001 281360 269013
rect 302320 269001 302326 269013
rect 302378 269001 302384 269053
rect 306352 269001 306358 269053
rect 306410 269041 306416 269053
rect 334288 269041 334294 269053
rect 306410 269013 334294 269041
rect 306410 269001 306416 269013
rect 334288 269001 334294 269013
rect 334346 269001 334352 269053
rect 345424 269001 345430 269053
rect 345482 269041 345488 269053
rect 484240 269041 484246 269053
rect 345482 269013 484246 269041
rect 345482 269001 345488 269013
rect 484240 269001 484246 269013
rect 484298 269001 484304 269053
rect 148624 268927 148630 268979
rect 148682 268967 148688 268979
rect 215728 268967 215734 268979
rect 148682 268939 215734 268967
rect 148682 268927 148688 268939
rect 215728 268927 215734 268939
rect 215786 268927 215792 268979
rect 253168 268927 253174 268979
rect 253226 268967 253232 268979
rect 254992 268967 254998 268979
rect 253226 268939 254998 268967
rect 253226 268927 253232 268939
rect 254992 268927 254998 268939
rect 255050 268927 255056 268979
rect 261232 268927 261238 268979
rect 261290 268967 261296 268979
rect 275056 268967 275062 268979
rect 261290 268939 275062 268967
rect 261290 268927 261296 268939
rect 275056 268927 275062 268939
rect 275114 268927 275120 268979
rect 282064 268927 282070 268979
rect 282122 268967 282128 268979
rect 298000 268967 298006 268979
rect 282122 268939 298006 268967
rect 282122 268927 282128 268939
rect 298000 268927 298006 268939
rect 298058 268927 298064 268979
rect 300688 268927 300694 268979
rect 300746 268967 300752 268979
rect 326800 268967 326806 268979
rect 300746 268939 326806 268967
rect 300746 268927 300752 268939
rect 326800 268927 326806 268939
rect 326858 268927 326864 268979
rect 342640 268927 342646 268979
rect 342698 268967 342704 268979
rect 477136 268967 477142 268979
rect 342698 268939 477142 268967
rect 342698 268927 342704 268939
rect 477136 268927 477142 268939
rect 477194 268927 477200 268979
rect 155728 268853 155734 268905
rect 155786 268893 155792 268905
rect 217360 268893 217366 268905
rect 155786 268865 217366 268893
rect 155786 268853 155792 268865
rect 217360 268853 217366 268865
rect 217418 268853 217424 268905
rect 264112 268853 264118 268905
rect 264170 268893 264176 268905
rect 282160 268893 282166 268905
rect 264170 268865 282166 268893
rect 264170 268853 264176 268865
rect 282160 268853 282166 268865
rect 282218 268853 282224 268905
rect 303760 268853 303766 268905
rect 303818 268893 303824 268905
rect 328336 268893 328342 268905
rect 303818 268865 328342 268893
rect 303818 268853 303824 268865
rect 328336 268853 328342 268865
rect 328394 268853 328400 268905
rect 339760 268853 339766 268905
rect 339818 268893 339824 268905
rect 470128 268893 470134 268905
rect 339818 268865 470134 268893
rect 339818 268853 339824 268865
rect 470128 268853 470134 268865
rect 470186 268853 470192 268905
rect 42064 268779 42070 268831
rect 42122 268819 42128 268831
rect 44176 268819 44182 268831
rect 42122 268791 44182 268819
rect 42122 268779 42128 268791
rect 44176 268779 44182 268791
rect 44234 268779 44240 268831
rect 156880 268779 156886 268831
rect 156938 268819 156944 268831
rect 218128 268819 218134 268831
rect 156938 268791 218134 268819
rect 156938 268779 156944 268791
rect 218128 268779 218134 268791
rect 218186 268779 218192 268831
rect 258160 268779 258166 268831
rect 258218 268819 258224 268831
rect 267952 268819 267958 268831
rect 258218 268791 267958 268819
rect 258218 268779 258224 268791
rect 267952 268779 267958 268791
rect 268010 268779 268016 268831
rect 289168 268779 289174 268831
rect 289226 268819 289232 268831
rect 310576 268819 310582 268831
rect 289226 268791 310582 268819
rect 289226 268779 289232 268791
rect 310576 268779 310582 268791
rect 310634 268779 310640 268831
rect 336880 268779 336886 268831
rect 336938 268819 336944 268831
rect 463024 268819 463030 268831
rect 336938 268791 463030 268819
rect 336938 268779 336944 268791
rect 463024 268779 463030 268791
rect 463082 268779 463088 268831
rect 162832 268705 162838 268757
rect 162890 268745 162896 268757
rect 219280 268745 219286 268757
rect 162890 268717 219286 268745
rect 162890 268705 162896 268717
rect 219280 268705 219286 268717
rect 219338 268705 219344 268757
rect 268432 268705 268438 268757
rect 268490 268745 268496 268757
rect 292816 268745 292822 268757
rect 268490 268717 292822 268745
rect 268490 268705 268496 268717
rect 292816 268705 292822 268717
rect 292874 268705 292880 268757
rect 334288 268705 334294 268757
rect 334346 268745 334352 268757
rect 455920 268745 455926 268757
rect 334346 268717 455926 268745
rect 334346 268705 334352 268717
rect 455920 268705 455926 268717
rect 455978 268705 455984 268757
rect 163984 268631 163990 268683
rect 164042 268671 164048 268683
rect 219952 268671 219958 268683
rect 164042 268643 219958 268671
rect 164042 268631 164048 268643
rect 219952 268631 219958 268643
rect 220010 268631 220016 268683
rect 254608 268631 254614 268683
rect 254666 268671 254672 268683
rect 258544 268671 258550 268683
rect 254666 268643 258550 268671
rect 254666 268631 254672 268643
rect 258544 268631 258550 268643
rect 258602 268631 258608 268683
rect 260560 268631 260566 268683
rect 260618 268671 260624 268683
rect 273904 268671 273910 268683
rect 260618 268643 273910 268671
rect 260618 268631 260624 268643
rect 273904 268631 273910 268643
rect 273962 268631 273968 268683
rect 331216 268631 331222 268683
rect 331274 268671 331280 268683
rect 448816 268671 448822 268683
rect 331274 268643 448822 268671
rect 331274 268631 331280 268643
rect 448816 268631 448822 268643
rect 448874 268631 448880 268683
rect 169744 268557 169750 268609
rect 169802 268597 169808 268609
rect 221200 268597 221206 268609
rect 169802 268569 221206 268597
rect 169802 268557 169808 268569
rect 221200 268557 221206 268569
rect 221258 268557 221264 268609
rect 328336 268557 328342 268609
rect 328394 268597 328400 268609
rect 441712 268597 441718 268609
rect 328394 268569 441718 268597
rect 328394 268557 328400 268569
rect 441712 268557 441718 268569
rect 441770 268557 441776 268609
rect 171088 268483 171094 268535
rect 171146 268523 171152 268535
rect 221776 268523 221782 268535
rect 171146 268495 221782 268523
rect 171146 268483 171152 268495
rect 221776 268483 221782 268495
rect 221834 268483 221840 268535
rect 263632 268483 263638 268535
rect 263690 268523 263696 268535
rect 281008 268523 281014 268535
rect 263690 268495 281014 268523
rect 263690 268483 263696 268495
rect 281008 268483 281014 268495
rect 281066 268483 281072 268535
rect 325744 268483 325750 268535
rect 325802 268523 325808 268535
rect 434608 268523 434614 268535
rect 325802 268495 434614 268523
rect 325802 268483 325808 268495
rect 434608 268483 434614 268495
rect 434666 268483 434672 268535
rect 176944 268409 176950 268461
rect 177002 268449 177008 268461
rect 223408 268449 223414 268461
rect 177002 268421 223414 268449
rect 177002 268409 177008 268421
rect 223408 268409 223414 268421
rect 223466 268409 223472 268461
rect 322576 268409 322582 268461
rect 322634 268449 322640 268461
rect 427504 268449 427510 268461
rect 322634 268421 427510 268449
rect 322634 268409 322640 268421
rect 427504 268409 427510 268421
rect 427562 268409 427568 268461
rect 178192 268335 178198 268387
rect 178250 268375 178256 268387
rect 223600 268375 223606 268387
rect 178250 268347 223606 268375
rect 178250 268335 178256 268347
rect 223600 268335 223606 268347
rect 223658 268335 223664 268387
rect 247888 268335 247894 268387
rect 247946 268375 247952 268387
rect 249808 268375 249814 268387
rect 247946 268347 249814 268375
rect 247946 268335 247952 268347
rect 249808 268335 249814 268347
rect 249866 268335 249872 268387
rect 255088 268335 255094 268387
rect 255146 268375 255152 268387
rect 259696 268375 259702 268387
rect 255146 268347 259702 268375
rect 255146 268335 255152 268347
rect 259696 268335 259702 268347
rect 259754 268335 259760 268387
rect 262960 268335 262966 268387
rect 263018 268375 263024 268387
rect 279760 268375 279766 268387
rect 263018 268347 279766 268375
rect 263018 268335 263024 268347
rect 279760 268335 279766 268347
rect 279818 268335 279824 268387
rect 319696 268335 319702 268387
rect 319754 268375 319760 268387
rect 420496 268375 420502 268387
rect 319754 268347 420502 268375
rect 319754 268335 319760 268347
rect 420496 268335 420502 268347
rect 420554 268335 420560 268387
rect 185680 268261 185686 268313
rect 185738 268301 185744 268313
rect 201136 268301 201142 268313
rect 185738 268273 201142 268301
rect 185738 268261 185744 268273
rect 201136 268261 201142 268273
rect 201194 268261 201200 268313
rect 207472 268261 207478 268313
rect 207530 268301 207536 268313
rect 207530 268273 210974 268301
rect 207530 268261 207536 268273
rect 192976 268187 192982 268239
rect 193034 268227 193040 268239
rect 210832 268227 210838 268239
rect 193034 268199 210838 268227
rect 193034 268187 193040 268199
rect 210832 268187 210838 268199
rect 210890 268187 210896 268239
rect 190096 268113 190102 268165
rect 190154 268153 190160 268165
rect 210736 268153 210742 268165
rect 190154 268125 210742 268153
rect 190154 268113 190160 268125
rect 210736 268113 210742 268125
rect 210794 268113 210800 268165
rect 210946 268153 210974 268273
rect 211024 268261 211030 268313
rect 211082 268301 211088 268313
rect 218608 268301 218614 268313
rect 211082 268273 218614 268301
rect 211082 268261 211088 268273
rect 218608 268261 218614 268273
rect 218666 268261 218672 268313
rect 221488 268261 221494 268313
rect 221546 268301 221552 268313
rect 227824 268301 227830 268313
rect 221546 268273 227830 268301
rect 221546 268261 221552 268273
rect 227824 268261 227830 268273
rect 227882 268261 227888 268313
rect 312304 268261 312310 268313
rect 312362 268301 312368 268313
rect 347056 268301 347062 268313
rect 312362 268273 347062 268301
rect 312362 268261 312368 268273
rect 347056 268261 347062 268273
rect 347114 268261 347120 268313
rect 224368 268187 224374 268239
rect 224426 268227 224432 268239
rect 230032 268227 230038 268239
rect 224426 268199 230038 268227
rect 224426 268187 224432 268199
rect 230032 268187 230038 268199
rect 230090 268187 230096 268239
rect 257008 268187 257014 268239
rect 257066 268227 257072 268239
rect 264400 268227 264406 268239
rect 257066 268199 264406 268227
rect 257066 268187 257072 268199
rect 264400 268187 264406 268199
rect 264458 268187 264464 268239
rect 332368 268187 332374 268239
rect 332426 268227 332432 268239
rect 344848 268227 344854 268239
rect 332426 268199 344854 268227
rect 332426 268187 332432 268199
rect 344848 268187 344854 268199
rect 344906 268187 344912 268239
rect 345232 268187 345238 268239
rect 345290 268227 345296 268239
rect 354544 268227 354550 268239
rect 345290 268199 354550 268227
rect 345290 268187 345296 268199
rect 354544 268187 354550 268199
rect 354602 268187 354608 268239
rect 394384 268187 394390 268239
rect 394442 268227 394448 268239
rect 604816 268227 604822 268239
rect 394442 268199 604822 268227
rect 394442 268187 394448 268199
rect 604816 268187 604822 268199
rect 604874 268187 604880 268239
rect 218896 268153 218902 268165
rect 210946 268125 218902 268153
rect 218896 268113 218902 268125
rect 218954 268113 218960 268165
rect 223696 268113 223702 268165
rect 223754 268153 223760 268165
rect 231472 268153 231478 268165
rect 223754 268125 231478 268153
rect 223754 268113 223760 268125
rect 231472 268113 231478 268125
rect 231530 268113 231536 268165
rect 334960 268113 334966 268165
rect 335018 268153 335024 268165
rect 348496 268153 348502 268165
rect 335018 268125 348502 268153
rect 335018 268113 335024 268125
rect 348496 268113 348502 268125
rect 348554 268113 348560 268165
rect 207376 268039 207382 268091
rect 207434 268079 207440 268091
rect 216880 268079 216886 268091
rect 207434 268051 216886 268079
rect 207434 268039 207440 268051
rect 216880 268039 216886 268051
rect 216938 268039 216944 268091
rect 221584 268039 221590 268091
rect 221642 268079 221648 268091
rect 230512 268079 230518 268091
rect 221642 268051 230518 268079
rect 221642 268039 221648 268051
rect 230512 268039 230518 268051
rect 230570 268039 230576 268091
rect 252688 268039 252694 268091
rect 252746 268079 252752 268091
rect 253744 268079 253750 268091
rect 252746 268051 253750 268079
rect 252746 268039 252752 268051
rect 253744 268039 253750 268051
rect 253802 268039 253808 268091
rect 341008 268039 341014 268091
rect 341066 268079 341072 268091
rect 341066 268051 357134 268079
rect 341066 268039 341072 268051
rect 209872 267965 209878 268017
rect 209930 268005 209936 268017
rect 212368 268005 212374 268017
rect 209930 267977 212374 268005
rect 209930 267965 209936 267977
rect 212368 267965 212374 267977
rect 212426 267965 212432 268017
rect 221680 267965 221686 268017
rect 221738 268005 221744 268017
rect 229072 268005 229078 268017
rect 221738 267977 229078 268005
rect 221738 267965 221744 267977
rect 229072 267965 229078 267977
rect 229130 267965 229136 268017
rect 337840 267965 337846 268017
rect 337898 268005 337904 268017
rect 354256 268005 354262 268017
rect 337898 267977 354262 268005
rect 337898 267965 337904 267977
rect 354256 267965 354262 267977
rect 354314 267965 354320 268017
rect 357106 268005 357134 268051
rect 357520 268005 357526 268017
rect 357106 267977 357526 268005
rect 357520 267965 357526 267977
rect 357578 267965 357584 268017
rect 207280 267891 207286 267943
rect 207338 267931 207344 267943
rect 209488 267931 209494 267943
rect 207338 267903 209494 267931
rect 207338 267891 207344 267903
rect 209488 267891 209494 267903
rect 209546 267891 209552 267943
rect 210640 267891 210646 267943
rect 210698 267931 210704 267943
rect 221008 267931 221014 267943
rect 210698 267903 221014 267931
rect 210698 267891 210704 267903
rect 221008 267891 221014 267903
rect 221066 267891 221072 267943
rect 224464 267891 224470 267943
rect 224522 267931 224528 267943
rect 228400 267931 228406 267943
rect 224522 267903 228406 267931
rect 224522 267891 224528 267903
rect 228400 267891 228406 267903
rect 228458 267891 228464 267943
rect 343600 267891 343606 267943
rect 343658 267931 343664 267943
rect 343658 267903 354302 267931
rect 343658 267891 343664 267903
rect 199120 267817 199126 267869
rect 199178 267857 199184 267869
rect 202288 267857 202294 267869
rect 199178 267829 202294 267857
rect 199178 267817 199184 267829
rect 202288 267817 202294 267829
rect 202346 267817 202352 267869
rect 209680 267817 209686 267869
rect 209738 267857 209744 267869
rect 211408 267857 211414 267869
rect 209738 267829 211414 267857
rect 209738 267817 209744 267829
rect 211408 267817 211414 267829
rect 211466 267817 211472 267869
rect 224560 267817 224566 267869
rect 224618 267857 224624 267869
rect 227632 267857 227638 267869
rect 224618 267829 227638 267857
rect 224618 267817 224624 267829
rect 227632 267817 227638 267829
rect 227690 267817 227696 267869
rect 282544 267817 282550 267869
rect 282602 267857 282608 267869
rect 299440 267857 299446 267869
rect 282602 267829 299446 267857
rect 282602 267817 282608 267829
rect 299440 267817 299446 267829
rect 299498 267817 299504 267869
rect 317104 267817 317110 267869
rect 317162 267857 317168 267869
rect 319024 267857 319030 267869
rect 317162 267829 319030 267857
rect 317162 267817 317168 267829
rect 319024 267817 319030 267829
rect 319082 267817 319088 267869
rect 354274 267857 354302 267903
rect 354544 267891 354550 267943
rect 354602 267931 354608 267943
rect 385456 267931 385462 267943
rect 354602 267903 385462 267931
rect 354602 267891 354608 267903
rect 385456 267891 385462 267903
rect 385514 267891 385520 267943
rect 360688 267857 360694 267869
rect 354274 267829 360694 267857
rect 360688 267817 360694 267829
rect 360746 267817 360752 267869
rect 407248 267817 407254 267869
rect 407306 267857 407312 267869
rect 409840 267857 409846 267869
rect 407306 267829 409846 267857
rect 407306 267817 407312 267829
rect 409840 267817 409846 267829
rect 409898 267817 409904 267869
rect 409936 267817 409942 267869
rect 409994 267857 410000 267869
rect 411856 267857 411862 267869
rect 409994 267829 411862 267857
rect 409994 267817 410000 267829
rect 411856 267817 411862 267829
rect 411914 267817 411920 267869
rect 354832 267743 354838 267795
rect 354890 267783 354896 267795
rect 506704 267783 506710 267795
rect 354890 267755 506710 267783
rect 354890 267743 354896 267755
rect 506704 267743 506710 267755
rect 506762 267743 506768 267795
rect 357424 267669 357430 267721
rect 357482 267709 357488 267721
rect 513808 267709 513814 267721
rect 357482 267681 513814 267709
rect 357482 267669 357488 267681
rect 513808 267669 513814 267681
rect 513866 267669 513872 267721
rect 360304 267595 360310 267647
rect 360362 267635 360368 267647
rect 520912 267635 520918 267647
rect 360362 267607 520918 267635
rect 360362 267595 360368 267607
rect 520912 267595 520918 267607
rect 520970 267595 520976 267647
rect 363376 267521 363382 267573
rect 363434 267561 363440 267573
rect 528016 267561 528022 267573
rect 363434 267533 528022 267561
rect 363434 267521 363440 267533
rect 528016 267521 528022 267533
rect 528074 267521 528080 267573
rect 365968 267447 365974 267499
rect 366026 267487 366032 267499
rect 535120 267487 535126 267499
rect 366026 267459 535126 267487
rect 366026 267447 366032 267459
rect 535120 267447 535126 267459
rect 535178 267447 535184 267499
rect 368944 267373 368950 267425
rect 369002 267413 369008 267425
rect 542224 267413 542230 267425
rect 369002 267385 542230 267413
rect 369002 267373 369008 267385
rect 542224 267373 542230 267385
rect 542282 267373 542288 267425
rect 375088 267299 375094 267351
rect 375146 267339 375152 267351
rect 557584 267339 557590 267351
rect 375146 267311 557590 267339
rect 375146 267299 375152 267311
rect 557584 267299 557590 267311
rect 557642 267299 557648 267351
rect 384880 267225 384886 267277
rect 384938 267265 384944 267277
rect 581200 267265 581206 267277
rect 384938 267237 581206 267265
rect 384938 267225 384944 267237
rect 581200 267225 581206 267237
rect 581258 267225 581264 267277
rect 386032 267151 386038 267203
rect 386090 267191 386096 267203
rect 584752 267191 584758 267203
rect 386090 267163 584758 267191
rect 386090 267151 386096 267163
rect 584752 267151 584758 267163
rect 584810 267151 584816 267203
rect 296464 267077 296470 267129
rect 296522 267117 296528 267129
rect 362512 267117 362518 267129
rect 296522 267089 362518 267117
rect 296522 267077 296528 267089
rect 362512 267077 362518 267089
rect 362570 267077 362576 267129
rect 387952 267077 387958 267129
rect 388010 267117 388016 267129
rect 589456 267117 589462 267129
rect 388010 267089 589462 267117
rect 388010 267077 388016 267089
rect 589456 267077 589462 267089
rect 589514 267077 589520 267129
rect 300208 267003 300214 267055
rect 300266 267043 300272 267055
rect 372016 267043 372022 267055
rect 300266 267015 372022 267043
rect 300266 267003 300272 267015
rect 372016 267003 372022 267015
rect 372074 267003 372080 267055
rect 391984 267003 391990 267055
rect 392042 267043 392048 267055
rect 598960 267043 598966 267055
rect 392042 267015 598966 267043
rect 392042 267003 392048 267015
rect 598960 267003 598966 267015
rect 599018 267003 599024 267055
rect 302032 266929 302038 266981
rect 302090 266969 302096 266981
rect 376720 266969 376726 266981
rect 302090 266941 376726 266969
rect 302090 266929 302096 266941
rect 376720 266929 376726 266941
rect 376778 266929 376784 266981
rect 393232 266929 393238 266981
rect 393290 266969 393296 266981
rect 602512 266969 602518 266981
rect 393290 266941 602518 266969
rect 393290 266929 393296 266941
rect 602512 266929 602518 266941
rect 602570 266929 602576 266981
rect 304432 266855 304438 266907
rect 304490 266895 304496 266907
rect 382576 266895 382582 266907
rect 304490 266867 382582 266895
rect 304490 266855 304496 266867
rect 382576 266855 382582 266867
rect 382634 266855 382640 266907
rect 396304 266855 396310 266907
rect 396362 266895 396368 266907
rect 609520 266895 609526 266907
rect 396362 266867 609526 266895
rect 396362 266855 396368 266867
rect 609520 266855 609526 266867
rect 609578 266855 609584 266907
rect 305008 266781 305014 266833
rect 305066 266821 305072 266833
rect 383824 266821 383830 266833
rect 305066 266793 383830 266821
rect 305066 266781 305072 266793
rect 383824 266781 383830 266793
rect 383882 266781 383888 266833
rect 398896 266781 398902 266833
rect 398954 266821 398960 266833
rect 616624 266821 616630 266833
rect 398954 266793 616630 266821
rect 398954 266781 398960 266793
rect 616624 266781 616630 266793
rect 616682 266781 616688 266833
rect 308080 266707 308086 266759
rect 308138 266747 308144 266759
rect 390928 266747 390934 266759
rect 308138 266719 390934 266747
rect 308138 266707 308144 266719
rect 390928 266707 390934 266719
rect 390986 266707 390992 266759
rect 401776 266707 401782 266759
rect 401834 266747 401840 266759
rect 623728 266747 623734 266759
rect 401834 266719 623734 266747
rect 401834 266707 401840 266719
rect 623728 266707 623734 266719
rect 623786 266707 623792 266759
rect 307312 266633 307318 266685
rect 307370 266673 307376 266685
rect 389680 266673 389686 266685
rect 307370 266645 389686 266673
rect 307370 266633 307376 266645
rect 389680 266633 389686 266645
rect 389738 266633 389744 266685
rect 403696 266633 403702 266685
rect 403754 266673 403760 266685
rect 628432 266673 628438 266685
rect 403754 266645 628438 266673
rect 403754 266633 403760 266645
rect 628432 266633 628438 266645
rect 628490 266633 628496 266685
rect 310672 266559 310678 266611
rect 310730 266599 310736 266611
rect 398032 266599 398038 266611
rect 310730 266571 398038 266599
rect 310730 266559 310736 266571
rect 398032 266559 398038 266571
rect 398090 266559 398096 266611
rect 404944 266559 404950 266611
rect 405002 266599 405008 266611
rect 630832 266599 630838 266611
rect 405002 266571 630838 266599
rect 405002 266559 405008 266571
rect 630832 266559 630838 266571
rect 630890 266559 630896 266611
rect 315952 266485 315958 266537
rect 316010 266525 316016 266537
rect 408976 266525 408982 266537
rect 316010 266497 408982 266525
rect 316010 266485 316016 266497
rect 408976 266485 408982 266497
rect 409034 266485 409040 266537
rect 409168 266485 409174 266537
rect 409226 266525 409232 266537
rect 641488 266525 641494 266537
rect 409226 266497 641494 266525
rect 409226 266485 409232 266497
rect 641488 266485 641494 266497
rect 641546 266485 641552 266537
rect 187216 266411 187222 266463
rect 187274 266451 187280 266463
rect 189712 266451 189718 266463
rect 187274 266423 189718 266451
rect 187274 266411 187280 266423
rect 189712 266411 189718 266423
rect 189770 266411 189776 266463
rect 311632 266411 311638 266463
rect 311690 266451 311696 266463
rect 400336 266451 400342 266463
rect 311690 266423 400342 266451
rect 311690 266411 311696 266423
rect 400336 266411 400342 266423
rect 400394 266411 400400 266463
rect 407824 266411 407830 266463
rect 407882 266451 407888 266463
rect 637936 266451 637942 266463
rect 407882 266423 637942 266451
rect 407882 266411 407888 266423
rect 637936 266411 637942 266423
rect 637994 266411 638000 266463
rect 46096 266337 46102 266389
rect 46154 266377 46160 266389
rect 652240 266377 652246 266389
rect 46154 266349 652246 266377
rect 46154 266337 46160 266349
rect 652240 266337 652246 266349
rect 652298 266337 652304 266389
rect 351952 266263 351958 266315
rect 352010 266303 352016 266315
rect 499600 266303 499606 266315
rect 352010 266275 499606 266303
rect 352010 266263 352016 266275
rect 499600 266263 499606 266275
rect 499658 266263 499664 266315
rect 348880 266189 348886 266241
rect 348938 266229 348944 266241
rect 492592 266229 492598 266241
rect 348938 266201 492598 266229
rect 348938 266189 348944 266201
rect 492592 266189 492598 266201
rect 492650 266189 492656 266241
rect 346000 266115 346006 266167
rect 346058 266155 346064 266167
rect 485488 266155 485494 266167
rect 346058 266127 485494 266155
rect 346058 266115 346064 266127
rect 485488 266115 485494 266127
rect 485546 266115 485552 266167
rect 343312 266041 343318 266093
rect 343370 266081 343376 266093
rect 478384 266081 478390 266093
rect 343370 266053 478390 266081
rect 343370 266041 343376 266053
rect 478384 266041 478390 266053
rect 478442 266041 478448 266093
rect 340240 265967 340246 266019
rect 340298 266007 340304 266019
rect 471280 266007 471286 266019
rect 340298 265979 471286 266007
rect 340298 265967 340304 265979
rect 471280 265967 471286 265979
rect 471338 265967 471344 266019
rect 337360 265893 337366 265945
rect 337418 265933 337424 265945
rect 464176 265933 464182 265945
rect 337418 265905 464182 265933
rect 337418 265893 337424 265905
rect 464176 265893 464182 265905
rect 464234 265893 464240 265945
rect 334768 265819 334774 265871
rect 334826 265859 334832 265871
rect 457072 265859 457078 265871
rect 334826 265831 457078 265859
rect 334826 265819 334832 265831
rect 457072 265819 457078 265831
rect 457130 265819 457136 265871
rect 330448 265745 330454 265797
rect 330506 265785 330512 265797
rect 446416 265785 446422 265797
rect 330506 265757 446422 265785
rect 330506 265745 330512 265757
rect 446416 265745 446422 265757
rect 446474 265745 446480 265797
rect 327568 265671 327574 265723
rect 327626 265711 327632 265723
rect 439312 265711 439318 265723
rect 327626 265683 439318 265711
rect 327626 265671 327632 265683
rect 439312 265671 439318 265683
rect 439370 265671 439376 265723
rect 324496 265597 324502 265649
rect 324554 265637 324560 265649
rect 432304 265637 432310 265649
rect 324554 265609 432310 265637
rect 324554 265597 324560 265609
rect 432304 265597 432310 265609
rect 432362 265597 432368 265649
rect 320176 265523 320182 265575
rect 320234 265563 320240 265575
rect 320234 265535 407582 265563
rect 320234 265523 320240 265535
rect 407554 265415 407582 265535
rect 408976 265523 408982 265575
rect 409034 265563 409040 265575
rect 410992 265563 410998 265575
rect 409034 265535 410998 265563
rect 409034 265523 409040 265535
rect 410992 265523 410998 265535
rect 411050 265523 411056 265575
rect 483088 265489 483094 265501
rect 437746 265461 483094 265489
rect 421648 265415 421654 265427
rect 407554 265387 421654 265415
rect 421648 265375 421654 265387
rect 421706 265375 421712 265427
rect 385456 265301 385462 265353
rect 385514 265341 385520 265353
rect 437746 265341 437774 265461
rect 483088 265449 483094 265461
rect 483146 265449 483152 265501
rect 385514 265313 437774 265341
rect 385514 265301 385520 265313
rect 23056 265005 23062 265057
rect 23114 265045 23120 265057
rect 46096 265045 46102 265057
rect 23114 265017 46102 265045
rect 23114 265005 23120 265017
rect 46096 265005 46102 265017
rect 46154 265005 46160 265057
rect 46192 264931 46198 264983
rect 46250 264971 46256 264983
rect 669808 264971 669814 264983
rect 46250 264943 669814 264971
rect 46250 264931 46256 264943
rect 669808 264931 669814 264943
rect 669866 264931 669872 264983
rect 360688 264857 360694 264909
rect 360746 264897 360752 264909
rect 479536 264897 479542 264909
rect 360746 264869 479542 264897
rect 360746 264857 360752 264869
rect 479536 264857 479542 264869
rect 479594 264857 479600 264909
rect 357520 264783 357526 264835
rect 357578 264823 357584 264835
rect 472432 264823 472438 264835
rect 357578 264795 472438 264823
rect 357578 264783 357584 264795
rect 472432 264783 472438 264795
rect 472490 264783 472496 264835
rect 354256 264709 354262 264761
rect 354314 264749 354320 264761
rect 465328 264749 465334 264761
rect 354314 264721 465334 264749
rect 354314 264709 354320 264721
rect 465328 264709 465334 264721
rect 465386 264709 465392 264761
rect 348496 264635 348502 264687
rect 348554 264675 348560 264687
rect 458224 264675 458230 264687
rect 348554 264647 458230 264675
rect 348554 264635 348560 264647
rect 458224 264635 458230 264647
rect 458282 264635 458288 264687
rect 331120 264561 331126 264613
rect 331178 264601 331184 264613
rect 447664 264601 447670 264613
rect 331178 264573 447670 264601
rect 331178 264561 331184 264573
rect 447664 264561 447670 264573
rect 447722 264561 447728 264613
rect 344848 264487 344854 264539
rect 344906 264527 344912 264539
rect 451216 264527 451222 264539
rect 344906 264499 451222 264527
rect 344906 264487 344912 264499
rect 451216 264487 451222 264499
rect 451274 264487 451280 264539
rect 328048 264413 328054 264465
rect 328106 264453 328112 264465
rect 440560 264453 440566 264465
rect 328106 264425 440566 264453
rect 328106 264413 328112 264425
rect 440560 264413 440566 264425
rect 440618 264413 440624 264465
rect 408016 264117 408022 264169
rect 408074 264157 408080 264169
rect 412816 264157 412822 264169
rect 408074 264129 412822 264157
rect 408074 264117 408080 264129
rect 412816 264117 412822 264129
rect 412874 264117 412880 264169
rect 324976 264043 324982 264095
rect 325034 264083 325040 264095
rect 433456 264083 433462 264095
rect 325034 264055 433462 264083
rect 325034 264043 325040 264055
rect 433456 264043 433462 264055
rect 433514 264043 433520 264095
rect 389440 263969 389446 264021
rect 389498 264009 389504 264021
rect 593008 264009 593014 264021
rect 389498 263981 593014 264009
rect 389498 263969 389504 263981
rect 593008 263969 593014 263981
rect 593066 263969 593072 264021
rect 392272 263895 392278 263947
rect 392330 263935 392336 263947
rect 600112 263935 600118 263947
rect 392330 263907 600118 263935
rect 392330 263895 392336 263907
rect 600112 263895 600118 263907
rect 600170 263895 600176 263947
rect 395440 263821 395446 263873
rect 395498 263861 395504 263873
rect 607216 263861 607222 263873
rect 395498 263833 607222 263861
rect 395498 263821 395504 263833
rect 607216 263821 607222 263833
rect 607274 263821 607280 263873
rect 399664 263747 399670 263799
rect 399722 263787 399728 263799
rect 617872 263787 617878 263799
rect 399722 263759 617878 263787
rect 399722 263747 399728 263759
rect 617872 263747 617878 263759
rect 617930 263747 617936 263799
rect 401104 263673 401110 263725
rect 401162 263713 401168 263725
rect 621424 263713 621430 263725
rect 401162 263685 621430 263713
rect 401162 263673 401168 263685
rect 621424 263673 621430 263685
rect 621482 263673 621488 263725
rect 23344 263599 23350 263651
rect 23402 263639 23408 263651
rect 46192 263639 46198 263651
rect 23402 263611 46198 263639
rect 23402 263599 23408 263611
rect 46192 263599 46198 263611
rect 46250 263599 46256 263651
rect 406864 263599 406870 263651
rect 406922 263639 406928 263651
rect 427600 263639 427606 263651
rect 406922 263611 427606 263639
rect 406922 263599 406928 263611
rect 427600 263599 427606 263611
rect 427658 263599 427664 263651
rect 631984 263639 631990 263651
rect 427810 263611 631990 263639
rect 23248 263525 23254 263577
rect 23306 263565 23312 263577
rect 46288 263565 46294 263577
rect 23306 263537 46294 263565
rect 23306 263525 23312 263537
rect 46288 263525 46294 263537
rect 46346 263525 46352 263577
rect 405424 263525 405430 263577
rect 405482 263565 405488 263577
rect 427810 263565 427838 263611
rect 631984 263599 631990 263611
rect 632042 263599 632048 263651
rect 405482 263537 427838 263565
rect 405482 263525 405488 263537
rect 427888 263525 427894 263577
rect 427946 263565 427952 263577
rect 635536 263565 635542 263577
rect 427946 263537 635542 263565
rect 427946 263525 427952 263537
rect 635536 263525 635542 263537
rect 635594 263525 635600 263577
rect 412816 263451 412822 263503
rect 412874 263491 412880 263503
rect 639088 263491 639094 263503
rect 412874 263463 639094 263491
rect 412874 263451 412880 263463
rect 639088 263451 639094 263463
rect 639146 263451 639152 263503
rect 656368 262415 656374 262467
rect 656426 262455 656432 262467
rect 676048 262455 676054 262467
rect 656426 262427 676054 262455
rect 656426 262415 656432 262427
rect 676048 262415 676054 262427
rect 676106 262415 676112 262467
rect 656176 262267 656182 262319
rect 656234 262307 656240 262319
rect 676240 262307 676246 262319
rect 656234 262279 676246 262307
rect 656234 262267 656240 262279
rect 676240 262267 676246 262279
rect 676298 262267 676304 262319
rect 23152 262119 23158 262171
rect 23210 262159 23216 262171
rect 46192 262159 46198 262171
rect 23210 262131 46198 262159
rect 23210 262119 23216 262131
rect 46192 262119 46198 262131
rect 46250 262119 46256 262171
rect 420400 262119 420406 262171
rect 420458 262159 420464 262171
rect 606160 262159 606166 262171
rect 420458 262131 606166 262159
rect 420458 262119 420464 262131
rect 606160 262119 606166 262131
rect 606218 262119 606224 262171
rect 673360 261601 673366 261653
rect 673418 261641 673424 261653
rect 676048 261641 676054 261653
rect 673418 261613 676054 261641
rect 673418 261601 673424 261613
rect 676048 261601 676054 261613
rect 676106 261601 676112 261653
rect 656080 259455 656086 259507
rect 656138 259495 656144 259507
rect 676240 259495 676246 259507
rect 656138 259467 676246 259495
rect 656138 259455 656144 259467
rect 676240 259455 676246 259467
rect 676298 259455 676304 259507
rect 420400 259233 420406 259285
rect 420458 259273 420464 259285
rect 606256 259273 606262 259285
rect 420458 259245 606262 259273
rect 420458 259233 420464 259245
rect 606256 259233 606262 259245
rect 606314 259233 606320 259285
rect 674704 256939 674710 256991
rect 674762 256979 674768 256991
rect 676048 256979 676054 256991
rect 674762 256951 676054 256979
rect 674762 256939 674768 256951
rect 676048 256939 676054 256951
rect 676106 256939 676112 256991
rect 40240 256347 40246 256399
rect 40298 256387 40304 256399
rect 48208 256387 48214 256399
rect 40298 256359 48214 256387
rect 40298 256347 40304 256359
rect 48208 256347 48214 256359
rect 48266 256347 48272 256399
rect 420400 256347 420406 256399
rect 420458 256387 420464 256399
rect 606352 256387 606358 256399
rect 420458 256359 606358 256387
rect 420458 256347 420464 256359
rect 606352 256347 606358 256359
rect 606410 256347 606416 256399
rect 41776 255385 41782 255437
rect 41834 255425 41840 255437
rect 53200 255425 53206 255437
rect 41834 255397 53206 255425
rect 41834 255385 41840 255397
rect 53200 255385 53206 255397
rect 53258 255385 53264 255437
rect 48016 255015 48022 255067
rect 48074 255055 48080 255067
rect 186352 255055 186358 255067
rect 48074 255027 186358 255055
rect 48074 255015 48080 255027
rect 186352 255015 186358 255027
rect 186410 255015 186416 255067
rect 41776 254941 41782 254993
rect 41834 254981 41840 254993
rect 43216 254981 43222 254993
rect 41834 254953 43222 254981
rect 41834 254941 41840 254953
rect 43216 254941 43222 254953
rect 43274 254941 43280 254993
rect 47536 254941 47542 254993
rect 47594 254981 47600 254993
rect 185968 254981 185974 254993
rect 47594 254953 185974 254981
rect 47594 254941 47600 254953
rect 185968 254941 185974 254953
rect 186026 254941 186032 254993
rect 48112 254867 48118 254919
rect 48170 254907 48176 254919
rect 186544 254907 186550 254919
rect 48170 254879 186550 254907
rect 48170 254867 48176 254879
rect 186544 254867 186550 254879
rect 186602 254867 186608 254919
rect 41776 254423 41782 254475
rect 41834 254463 41840 254475
rect 43216 254463 43222 254475
rect 41834 254435 43222 254463
rect 41834 254423 41840 254435
rect 43216 254423 43222 254435
rect 43274 254423 43280 254475
rect 675088 253609 675094 253661
rect 675146 253649 675152 253661
rect 676240 253649 676246 253661
rect 675146 253621 676246 253649
rect 675146 253609 675152 253621
rect 676240 253609 676246 253621
rect 676298 253609 676304 253661
rect 674896 253535 674902 253587
rect 674954 253575 674960 253587
rect 675952 253575 675958 253587
rect 674954 253547 675958 253575
rect 674954 253535 674960 253547
rect 675952 253535 675958 253547
rect 676010 253535 676016 253587
rect 41584 253461 41590 253513
rect 41642 253501 41648 253513
rect 56176 253501 56182 253513
rect 41642 253473 56182 253501
rect 41642 253461 41648 253473
rect 56176 253461 56182 253473
rect 56234 253461 56240 253513
rect 420400 253461 420406 253513
rect 420458 253501 420464 253513
rect 603280 253501 603286 253513
rect 420458 253473 603286 253501
rect 420458 253461 420464 253473
rect 603280 253461 603286 253473
rect 603338 253461 603344 253513
rect 675280 253461 675286 253513
rect 675338 253501 675344 253513
rect 676048 253501 676054 253513
rect 675338 253473 676054 253501
rect 675338 253461 675344 253473
rect 676048 253461 676054 253473
rect 676106 253461 676112 253513
rect 141040 252425 141046 252477
rect 141098 252465 141104 252477
rect 174256 252465 174262 252477
rect 141098 252437 174262 252465
rect 141098 252425 141104 252437
rect 174256 252425 174262 252437
rect 174314 252425 174320 252477
rect 97840 252351 97846 252403
rect 97898 252391 97904 252403
rect 156880 252391 156886 252403
rect 97898 252363 156886 252391
rect 97898 252351 97904 252363
rect 156880 252351 156886 252363
rect 156938 252351 156944 252403
rect 94960 252277 94966 252329
rect 95018 252317 95024 252329
rect 154000 252317 154006 252329
rect 95018 252289 154006 252317
rect 95018 252277 95024 252289
rect 154000 252277 154006 252289
rect 154058 252277 154064 252329
rect 103600 252203 103606 252255
rect 103658 252243 103664 252255
rect 165520 252243 165526 252255
rect 103658 252215 165526 252243
rect 103658 252203 103664 252215
rect 165520 252203 165526 252215
rect 165578 252203 165584 252255
rect 106480 252129 106486 252181
rect 106538 252169 106544 252181
rect 171280 252169 171286 252181
rect 106538 252141 171286 252169
rect 106538 252129 106544 252141
rect 171280 252129 171286 252141
rect 171338 252129 171344 252181
rect 109360 252055 109366 252107
rect 109418 252095 109424 252107
rect 179920 252095 179926 252107
rect 109418 252067 179926 252095
rect 109418 252055 109424 252067
rect 179920 252055 179926 252067
rect 179978 252055 179984 252107
rect 56080 251981 56086 252033
rect 56138 252021 56144 252033
rect 186448 252021 186454 252033
rect 56138 251993 186454 252021
rect 56138 251981 56144 251993
rect 186448 251981 186454 251993
rect 186506 251981 186512 252033
rect 674512 250723 674518 250775
rect 674570 250763 674576 250775
rect 675952 250763 675958 250775
rect 674570 250735 675958 250763
rect 674570 250723 674576 250735
rect 675952 250723 675958 250735
rect 676010 250723 676016 250775
rect 674608 250649 674614 250701
rect 674666 250689 674672 250701
rect 676240 250689 676246 250701
rect 674666 250661 676246 250689
rect 674666 250649 674672 250661
rect 676240 250649 676246 250661
rect 676298 250649 676304 250701
rect 420400 250575 420406 250627
rect 420458 250615 420464 250627
rect 603376 250615 603382 250627
rect 420458 250587 603382 250615
rect 420458 250575 420464 250587
rect 603376 250575 603382 250587
rect 603434 250575 603440 250627
rect 674992 250575 674998 250627
rect 675050 250615 675056 250627
rect 676048 250615 676054 250627
rect 675050 250587 676054 250615
rect 675050 250575 675056 250587
rect 676048 250575 676054 250587
rect 676106 250575 676112 250627
rect 135280 249909 135286 249961
rect 135338 249949 135344 249961
rect 145552 249949 145558 249961
rect 135338 249921 145558 249949
rect 135338 249909 135344 249921
rect 145552 249909 145558 249921
rect 145610 249909 145616 249961
rect 138160 249835 138166 249887
rect 138218 249875 138224 249887
rect 171472 249875 171478 249887
rect 138218 249847 171478 249875
rect 138218 249835 138224 249847
rect 171472 249835 171478 249847
rect 171530 249835 171536 249887
rect 118000 249761 118006 249813
rect 118058 249801 118064 249813
rect 156976 249801 156982 249813
rect 118058 249773 156982 249801
rect 118058 249761 118064 249773
rect 156976 249761 156982 249773
rect 157034 249761 157040 249813
rect 123760 249687 123766 249739
rect 123818 249727 123824 249739
rect 162736 249727 162742 249739
rect 123818 249699 162742 249727
rect 123818 249687 123824 249699
rect 162736 249687 162742 249699
rect 162794 249687 162800 249739
rect 126640 249613 126646 249665
rect 126698 249653 126704 249665
rect 168496 249653 168502 249665
rect 126698 249625 168502 249653
rect 126698 249613 126704 249625
rect 168496 249613 168502 249625
rect 168554 249613 168560 249665
rect 120880 249539 120886 249591
rect 120938 249579 120944 249591
rect 165616 249579 165622 249591
rect 120938 249551 165622 249579
rect 120938 249539 120944 249551
rect 165616 249539 165622 249551
rect 165674 249539 165680 249591
rect 132400 249465 132406 249517
rect 132458 249505 132464 249517
rect 180112 249505 180118 249517
rect 132458 249477 180118 249505
rect 132458 249465 132464 249477
rect 180112 249465 180118 249477
rect 180170 249465 180176 249517
rect 92080 249391 92086 249443
rect 92138 249431 92144 249443
rect 159760 249431 159766 249443
rect 92138 249403 159766 249431
rect 92138 249391 92144 249403
rect 159760 249391 159766 249403
rect 159818 249391 159824 249443
rect 77680 249317 77686 249369
rect 77738 249357 77744 249369
rect 145360 249357 145366 249369
rect 77738 249329 145366 249357
rect 77738 249317 77744 249329
rect 145360 249317 145366 249329
rect 145418 249317 145424 249369
rect 86320 249243 86326 249295
rect 86378 249283 86384 249295
rect 177040 249283 177046 249295
rect 86378 249255 177046 249283
rect 86378 249243 86384 249255
rect 177040 249243 177046 249255
rect 177098 249243 177104 249295
rect 80560 249169 80566 249221
rect 80618 249209 80624 249221
rect 182800 249209 182806 249221
rect 80618 249181 182806 249209
rect 80618 249169 80624 249181
rect 182800 249169 182806 249181
rect 182858 249169 182864 249221
rect 47920 249095 47926 249147
rect 47978 249135 47984 249147
rect 186736 249135 186742 249147
rect 47978 249107 186742 249135
rect 47978 249095 47984 249107
rect 186736 249095 186742 249107
rect 186794 249095 186800 249147
rect 646672 249095 646678 249147
rect 646730 249135 646736 249147
rect 679984 249135 679990 249147
rect 646730 249107 679990 249135
rect 646730 249095 646736 249107
rect 679984 249095 679990 249107
rect 680042 249095 680048 249147
rect 420304 247763 420310 247815
rect 420362 247803 420368 247815
rect 603472 247803 603478 247815
rect 420362 247775 603478 247803
rect 420362 247763 420368 247775
rect 603472 247763 603478 247775
rect 603530 247763 603536 247815
rect 420400 247689 420406 247741
rect 420458 247729 420464 247741
rect 629200 247729 629206 247741
rect 420458 247701 629206 247729
rect 420458 247689 420464 247701
rect 629200 247689 629206 247701
rect 629258 247689 629264 247741
rect 675760 247097 675766 247149
rect 675818 247097 675824 247149
rect 112240 246653 112246 246705
rect 112298 246693 112304 246705
rect 185776 246693 185782 246705
rect 112298 246665 185782 246693
rect 112298 246653 112304 246665
rect 185776 246653 185782 246665
rect 185834 246653 185840 246705
rect 675088 246653 675094 246705
rect 675146 246693 675152 246705
rect 675472 246693 675478 246705
rect 675146 246665 675478 246693
rect 675146 246653 675152 246665
rect 675472 246653 675478 246665
rect 675530 246653 675536 246705
rect 675778 246631 675806 247097
rect 47632 246579 47638 246631
rect 47690 246619 47696 246631
rect 186064 246619 186070 246631
rect 47690 246591 186070 246619
rect 47690 246579 47696 246591
rect 186064 246579 186070 246591
rect 186122 246579 186128 246631
rect 675760 246579 675766 246631
rect 675818 246579 675824 246631
rect 47728 246505 47734 246557
rect 47786 246545 47792 246557
rect 186256 246545 186262 246557
rect 47786 246517 186262 246545
rect 47786 246505 47792 246517
rect 186256 246505 186262 246517
rect 186314 246505 186320 246557
rect 47440 246431 47446 246483
rect 47498 246471 47504 246483
rect 186160 246471 186166 246483
rect 47498 246443 186166 246471
rect 47498 246431 47504 246443
rect 186160 246431 186166 246443
rect 186218 246431 186224 246483
rect 47824 246357 47830 246409
rect 47882 246397 47888 246409
rect 186640 246397 186646 246409
rect 47882 246369 186646 246397
rect 47882 246357 47888 246369
rect 186640 246357 186646 246369
rect 186698 246357 186704 246409
rect 45520 246283 45526 246335
rect 45578 246323 45584 246335
rect 186832 246323 186838 246335
rect 45578 246295 186838 246323
rect 45578 246283 45584 246295
rect 186832 246283 186838 246295
rect 186890 246283 186896 246335
rect 44272 246209 44278 246261
rect 44330 246249 44336 246261
rect 187024 246249 187030 246261
rect 44330 246221 187030 246249
rect 44330 246209 44336 246221
rect 187024 246209 187030 246221
rect 187082 246209 187088 246261
rect 674704 245395 674710 245447
rect 674762 245435 674768 245447
rect 675376 245435 675382 245447
rect 674762 245407 675382 245435
rect 674762 245395 674768 245407
rect 675376 245395 675382 245407
rect 675434 245395 675440 245447
rect 41584 244951 41590 245003
rect 41642 244991 41648 245003
rect 145456 244991 145462 245003
rect 41642 244963 145462 244991
rect 41642 244951 41648 244963
rect 145456 244951 145462 244963
rect 145514 244951 145520 245003
rect 44752 244877 44758 244929
rect 44810 244917 44816 244929
rect 186928 244917 186934 244929
rect 44810 244889 186934 244917
rect 44810 244877 44816 244889
rect 186928 244877 186934 244889
rect 186986 244877 186992 244929
rect 41776 244803 41782 244855
rect 41834 244843 41840 244855
rect 145648 244843 145654 244855
rect 41834 244815 145654 244843
rect 41834 244803 41840 244815
rect 145648 244803 145654 244815
rect 145706 244803 145712 244855
rect 420400 244803 420406 244855
rect 420458 244843 420464 244855
rect 629296 244843 629302 244855
rect 420458 244815 629302 244843
rect 420458 244803 420464 244815
rect 629296 244803 629302 244815
rect 629354 244803 629360 244855
rect 674896 242879 674902 242931
rect 674954 242919 674960 242931
rect 675376 242919 675382 242931
rect 674954 242891 675382 242919
rect 674954 242879 674960 242891
rect 675376 242879 675382 242891
rect 675434 242879 675440 242931
rect 44656 242805 44662 242857
rect 44714 242845 44720 242857
rect 185680 242845 185686 242857
rect 44714 242817 185686 242845
rect 44714 242805 44720 242817
rect 185680 242805 185686 242817
rect 185738 242805 185744 242857
rect 44560 242731 44566 242783
rect 44618 242771 44624 242783
rect 185584 242771 185590 242783
rect 44618 242743 185590 242771
rect 44618 242731 44624 242743
rect 185584 242731 185590 242743
rect 185642 242731 185648 242783
rect 44848 242657 44854 242709
rect 44906 242697 44912 242709
rect 185872 242697 185878 242709
rect 44906 242669 185878 242697
rect 44906 242657 44912 242669
rect 185872 242657 185878 242669
rect 185930 242657 185936 242709
rect 41584 242583 41590 242635
rect 41642 242623 41648 242635
rect 142576 242623 142582 242635
rect 41642 242595 142582 242623
rect 41642 242583 41648 242595
rect 142576 242583 142582 242595
rect 142634 242583 142640 242635
rect 675184 242287 675190 242339
rect 675242 242327 675248 242339
rect 675376 242327 675382 242339
rect 675242 242299 675382 242327
rect 675242 242287 675248 242299
rect 675376 242287 675382 242299
rect 675434 242287 675440 242339
rect 420400 241917 420406 241969
rect 420458 241957 420464 241969
rect 600400 241957 600406 241969
rect 420458 241929 600406 241957
rect 420458 241917 420464 241929
rect 600400 241917 600406 241929
rect 600458 241917 600464 241969
rect 655888 241843 655894 241895
rect 655946 241883 655952 241895
rect 675088 241883 675094 241895
rect 655946 241855 675094 241883
rect 655946 241843 655952 241855
rect 675088 241843 675094 241855
rect 675146 241843 675152 241895
rect 674992 241769 674998 241821
rect 675050 241809 675056 241821
rect 675376 241809 675382 241821
rect 675050 241781 675382 241809
rect 675050 241769 675056 241781
rect 675376 241769 675382 241781
rect 675434 241769 675440 241821
rect 41776 240807 41782 240859
rect 41834 240807 41840 240859
rect 41794 240563 41822 240807
rect 41776 240511 41782 240563
rect 41834 240511 41840 240563
rect 380848 239919 380854 239971
rect 380906 239959 380912 239971
rect 412048 239959 412054 239971
rect 380906 239931 412054 239959
rect 380906 239919 380912 239931
rect 412048 239919 412054 239931
rect 412106 239919 412112 239971
rect 409552 239845 409558 239897
rect 409610 239885 409616 239897
rect 412144 239885 412150 239897
rect 409610 239857 412150 239885
rect 409610 239845 409616 239857
rect 412144 239845 412150 239857
rect 412202 239845 412208 239897
rect 357136 239771 357142 239823
rect 357194 239811 357200 239823
rect 434608 239811 434614 239823
rect 357194 239783 434614 239811
rect 357194 239771 357200 239783
rect 434608 239771 434614 239783
rect 434666 239771 434672 239823
rect 377296 239697 377302 239749
rect 377354 239737 377360 239749
rect 446704 239737 446710 239749
rect 377354 239709 446710 239737
rect 377354 239697 377360 239709
rect 446704 239697 446710 239709
rect 446762 239697 446768 239749
rect 385360 239623 385366 239675
rect 385418 239663 385424 239675
rect 470896 239663 470902 239675
rect 385418 239635 470902 239663
rect 385418 239623 385424 239635
rect 470896 239623 470902 239635
rect 470954 239623 470960 239675
rect 374416 239549 374422 239601
rect 374474 239589 374480 239601
rect 488272 239589 488278 239601
rect 374474 239561 488278 239589
rect 374474 239549 374480 239561
rect 488272 239549 488278 239561
rect 488330 239549 488336 239601
rect 334288 239475 334294 239527
rect 334346 239515 334352 239527
rect 458800 239515 458806 239527
rect 334346 239487 458806 239515
rect 334346 239475 334352 239487
rect 458800 239475 458806 239487
rect 458858 239475 458864 239527
rect 394672 239401 394678 239453
rect 394730 239441 394736 239453
rect 532816 239441 532822 239453
rect 394730 239413 532822 239441
rect 394730 239401 394736 239413
rect 532816 239401 532822 239413
rect 532874 239401 532880 239453
rect 397744 239327 397750 239379
rect 397802 239367 397808 239379
rect 541456 239367 541462 239379
rect 397802 239339 541462 239367
rect 397802 239327 397808 239339
rect 541456 239327 541462 239339
rect 541514 239327 541520 239379
rect 406000 239253 406006 239305
rect 406058 239293 406064 239305
rect 550864 239293 550870 239305
rect 406058 239265 550870 239293
rect 406058 239253 406064 239265
rect 550864 239253 550870 239265
rect 550922 239253 550928 239305
rect 420400 239179 420406 239231
rect 420458 239219 420464 239231
rect 599152 239219 599158 239231
rect 420458 239191 599158 239219
rect 420458 239179 420464 239191
rect 599152 239179 599158 239191
rect 599210 239179 599216 239231
rect 350416 239105 350422 239157
rect 350474 239145 350480 239157
rect 508624 239145 508630 239157
rect 350474 239117 508630 239145
rect 350474 239105 350480 239117
rect 508624 239105 508630 239117
rect 508682 239105 508688 239157
rect 368560 239031 368566 239083
rect 368618 239071 368624 239083
rect 544816 239071 544822 239083
rect 368618 239043 544822 239071
rect 368618 239031 368624 239043
rect 544816 239031 544822 239043
rect 544874 239031 544880 239083
rect 324400 238957 324406 239009
rect 324458 238997 324464 239009
rect 455056 238997 455062 239009
rect 324458 238969 455062 238997
rect 324458 238957 324464 238969
rect 455056 238957 455062 238969
rect 455114 238957 455120 239009
rect 323920 238883 323926 238935
rect 323978 238923 323984 238935
rect 455152 238923 455158 238935
rect 323978 238895 455158 238923
rect 323978 238883 323984 238895
rect 455152 238883 455158 238895
rect 455210 238883 455216 238935
rect 326704 238809 326710 238861
rect 326762 238849 326768 238861
rect 462544 238849 462550 238861
rect 326762 238821 462550 238849
rect 326762 238809 326768 238821
rect 462544 238809 462550 238821
rect 462602 238809 462608 238861
rect 328912 238735 328918 238787
rect 328970 238775 328976 238787
rect 464752 238775 464758 238787
rect 328970 238747 464758 238775
rect 328970 238735 328976 238747
rect 464752 238735 464758 238747
rect 464810 238735 464816 238787
rect 329872 238661 329878 238713
rect 329930 238701 329936 238713
rect 468592 238701 468598 238713
rect 329930 238673 468598 238701
rect 329930 238661 329936 238673
rect 468592 238661 468598 238673
rect 468650 238661 468656 238713
rect 332656 238587 332662 238639
rect 332714 238627 332720 238639
rect 474640 238627 474646 238639
rect 332714 238599 474646 238627
rect 332714 238587 332720 238599
rect 474640 238587 474646 238599
rect 474698 238587 474704 238639
rect 674608 238587 674614 238639
rect 674666 238627 674672 238639
rect 675376 238627 675382 238639
rect 674666 238599 675382 238627
rect 674666 238587 674672 238599
rect 675376 238587 675382 238599
rect 675434 238587 675440 238639
rect 335728 238513 335734 238565
rect 335786 238553 335792 238565
rect 480688 238553 480694 238565
rect 335786 238525 480694 238553
rect 335786 238513 335792 238525
rect 480688 238513 480694 238525
rect 480746 238513 480752 238565
rect 336688 238439 336694 238491
rect 336746 238479 336752 238491
rect 478096 238479 478102 238491
rect 336746 238451 478102 238479
rect 336746 238439 336752 238451
rect 478096 238439 478102 238451
rect 478154 238439 478160 238491
rect 338992 238365 338998 238417
rect 339050 238405 339056 238417
rect 486736 238405 486742 238417
rect 339050 238377 486742 238405
rect 339050 238365 339056 238377
rect 486736 238365 486742 238377
rect 486794 238365 486800 238417
rect 341776 238291 341782 238343
rect 341834 238331 341840 238343
rect 492784 238331 492790 238343
rect 341834 238303 492790 238331
rect 341834 238291 341840 238303
rect 492784 238291 492790 238303
rect 492842 238291 492848 238343
rect 345328 238217 345334 238269
rect 345386 238257 345392 238269
rect 500272 238257 500278 238269
rect 345386 238229 500278 238257
rect 345386 238217 345392 238229
rect 500272 238217 500278 238229
rect 500330 238217 500336 238269
rect 346672 238143 346678 238195
rect 346730 238183 346736 238195
rect 503344 238183 503350 238195
rect 346730 238155 503350 238183
rect 346730 238143 346736 238155
rect 503344 238143 503350 238155
rect 503402 238143 503408 238195
rect 349936 238069 349942 238121
rect 349994 238109 350000 238121
rect 509392 238109 509398 238121
rect 349994 238081 509398 238109
rect 349994 238069 350000 238081
rect 509392 238069 509398 238081
rect 509450 238069 509456 238121
rect 353488 237995 353494 238047
rect 353546 238035 353552 238047
rect 514672 238035 514678 238047
rect 353546 238007 514678 238035
rect 353546 237995 353552 238007
rect 514672 237995 514678 238007
rect 514730 237995 514736 238047
rect 352720 237921 352726 237973
rect 352778 237961 352784 237973
rect 512752 237961 512758 237973
rect 352778 237933 512758 237961
rect 352778 237921 352784 237933
rect 512752 237921 512758 237933
rect 512810 237921 512816 237973
rect 355696 237847 355702 237899
rect 355754 237887 355760 237899
rect 522160 237887 522166 237899
rect 355754 237859 522166 237887
rect 355754 237847 355760 237859
rect 522160 237847 522166 237859
rect 522218 237847 522224 237899
rect 363088 237773 363094 237825
rect 363146 237813 363152 237825
rect 535120 237813 535126 237825
rect 363146 237785 535126 237813
rect 363146 237773 363152 237785
rect 535120 237773 535126 237785
rect 535178 237773 535184 237825
rect 275344 237699 275350 237751
rect 275402 237739 275408 237751
rect 357520 237739 357526 237751
rect 275402 237711 357526 237739
rect 275402 237699 275408 237711
rect 357520 237699 357526 237711
rect 357578 237699 357584 237751
rect 361744 237699 361750 237751
rect 361802 237739 361808 237751
rect 533488 237739 533494 237751
rect 361802 237711 533494 237739
rect 361802 237699 361808 237711
rect 533488 237699 533494 237711
rect 533546 237699 533552 237751
rect 277072 237625 277078 237677
rect 277130 237665 277136 237677
rect 363664 237665 363670 237677
rect 277130 237637 363670 237665
rect 277130 237625 277136 237637
rect 363664 237625 363670 237637
rect 363722 237625 363728 237677
rect 364432 237625 364438 237677
rect 364490 237665 364496 237677
rect 535792 237665 535798 237677
rect 364490 237637 535798 237665
rect 364490 237625 364496 237637
rect 535792 237625 535798 237637
rect 535850 237625 535856 237677
rect 365872 237551 365878 237603
rect 365930 237591 365936 237603
rect 541072 237591 541078 237603
rect 365930 237563 541078 237591
rect 365930 237551 365936 237563
rect 541072 237551 541078 237563
rect 541130 237551 541136 237603
rect 674512 237551 674518 237603
rect 674570 237591 674576 237603
rect 675376 237591 675382 237603
rect 674570 237563 675382 237591
rect 674570 237551 674576 237563
rect 675376 237551 675382 237563
rect 675434 237551 675440 237603
rect 320848 237477 320854 237529
rect 320906 237517 320912 237529
rect 450448 237517 450454 237529
rect 320906 237489 450454 237517
rect 320906 237477 320912 237489
rect 450448 237477 450454 237489
rect 450506 237477 450512 237529
rect 317584 237403 317590 237455
rect 317642 237443 317648 237455
rect 444496 237443 444502 237455
rect 317642 237415 444502 237443
rect 317642 237403 317648 237415
rect 444496 237403 444502 237415
rect 444554 237403 444560 237455
rect 317104 237329 317110 237381
rect 317162 237369 317168 237381
rect 441424 237369 441430 237381
rect 317162 237341 441430 237369
rect 317162 237329 317168 237341
rect 441424 237329 441430 237341
rect 441482 237329 441488 237381
rect 314800 237255 314806 237307
rect 314858 237295 314864 237307
rect 438352 237295 438358 237307
rect 314858 237267 438358 237295
rect 314858 237255 314864 237267
rect 438352 237255 438358 237267
rect 438410 237255 438416 237307
rect 311536 237181 311542 237233
rect 311594 237221 311600 237233
rect 432400 237221 432406 237233
rect 311594 237193 432406 237221
rect 311594 237181 311600 237193
rect 432400 237181 432406 237193
rect 432458 237181 432464 237233
rect 308560 237107 308566 237159
rect 308618 237147 308624 237159
rect 426352 237147 426358 237159
rect 308618 237119 426358 237147
rect 308618 237107 308624 237119
rect 426352 237107 426358 237119
rect 426410 237107 426416 237159
rect 310768 237033 310774 237085
rect 310826 237073 310832 237085
rect 428656 237073 428662 237085
rect 310826 237045 428662 237073
rect 310826 237033 310832 237045
rect 428656 237033 428662 237045
rect 428714 237033 428720 237085
rect 305776 236959 305782 237011
rect 305834 236999 305840 237011
rect 420304 236999 420310 237011
rect 305834 236971 420310 236999
rect 305834 236959 305840 236971
rect 420304 236959 420310 236971
rect 420362 236959 420368 237011
rect 298960 236885 298966 236937
rect 299018 236925 299024 236937
rect 404464 236925 404470 236937
rect 299018 236897 404470 236925
rect 299018 236885 299024 236897
rect 404464 236885 404470 236897
rect 404522 236885 404528 236937
rect 405904 236885 405910 236937
rect 405962 236925 405968 236937
rect 414448 236925 414454 236937
rect 405962 236897 414454 236925
rect 405962 236885 405968 236897
rect 414448 236885 414454 236897
rect 414506 236885 414512 236937
rect 279856 236811 279862 236863
rect 279914 236851 279920 236863
rect 370480 236851 370486 236863
rect 279914 236823 370486 236851
rect 279914 236811 279920 236823
rect 370480 236811 370486 236823
rect 370538 236811 370544 236863
rect 386992 236811 386998 236863
rect 387050 236851 387056 236863
rect 387568 236851 387574 236863
rect 387050 236823 387574 236851
rect 387050 236811 387056 236823
rect 387568 236811 387574 236823
rect 387626 236811 387632 236863
rect 397072 236811 397078 236863
rect 397130 236851 397136 236863
rect 397648 236851 397654 236863
rect 397130 236823 397654 236851
rect 397130 236811 397136 236823
rect 397648 236811 397654 236823
rect 397706 236811 397712 236863
rect 398032 236811 398038 236863
rect 398090 236851 398096 236863
rect 413584 236851 413590 236863
rect 398090 236823 413590 236851
rect 398090 236811 398096 236823
rect 413584 236811 413590 236823
rect 413642 236811 413648 236863
rect 278416 236737 278422 236789
rect 278474 236777 278480 236789
rect 366736 236777 366742 236789
rect 278474 236749 366742 236777
rect 278474 236737 278480 236749
rect 366736 236737 366742 236749
rect 366794 236737 366800 236789
rect 396976 236737 396982 236789
rect 397034 236777 397040 236789
rect 413392 236777 413398 236789
rect 397034 236749 413398 236777
rect 397034 236737 397040 236749
rect 413392 236737 413398 236749
rect 413450 236737 413456 236789
rect 379792 236663 379798 236715
rect 379850 236703 379856 236715
rect 398320 236703 398326 236715
rect 379850 236675 398326 236703
rect 379850 236663 379856 236675
rect 398320 236663 398326 236675
rect 398378 236663 398384 236715
rect 410704 236367 410710 236419
rect 410762 236407 410768 236419
rect 442192 236407 442198 236419
rect 410762 236379 442198 236407
rect 410762 236367 410768 236379
rect 442192 236367 442198 236379
rect 442250 236367 442256 236419
rect 390736 236293 390742 236345
rect 390794 236333 390800 236345
rect 492016 236333 492022 236345
rect 390794 236305 492022 236333
rect 390794 236293 390800 236305
rect 492016 236293 492022 236305
rect 492074 236293 492080 236345
rect 394576 236219 394582 236271
rect 394634 236259 394640 236271
rect 505648 236259 505654 236271
rect 394634 236231 505654 236259
rect 394634 236219 394640 236231
rect 505648 236219 505654 236231
rect 505706 236219 505712 236271
rect 382384 236145 382390 236197
rect 382442 236185 382448 236197
rect 397360 236185 397366 236197
rect 382442 236157 397366 236185
rect 382442 236145 382448 236157
rect 397360 236145 397366 236157
rect 397418 236145 397424 236197
rect 400336 236145 400342 236197
rect 400394 236185 400400 236197
rect 523792 236185 523798 236197
rect 400394 236157 523798 236185
rect 400394 236145 400400 236157
rect 523792 236145 523798 236157
rect 523850 236145 523856 236197
rect 251056 236071 251062 236123
rect 251114 236111 251120 236123
rect 273712 236111 273718 236123
rect 251114 236083 273718 236111
rect 251114 236071 251120 236083
rect 273712 236071 273718 236083
rect 273770 236071 273776 236123
rect 277552 236071 277558 236123
rect 277610 236111 277616 236123
rect 313936 236111 313942 236123
rect 277610 236083 313942 236111
rect 277610 236071 277616 236083
rect 313936 236071 313942 236083
rect 313994 236071 314000 236123
rect 326128 236071 326134 236123
rect 326186 236111 326192 236123
rect 334288 236111 334294 236123
rect 326186 236083 334294 236111
rect 326186 236071 326192 236083
rect 334288 236071 334294 236083
rect 334346 236071 334352 236123
rect 341200 236071 341206 236123
rect 341258 236111 341264 236123
rect 374416 236111 374422 236123
rect 341258 236083 374422 236111
rect 341258 236071 341264 236083
rect 374416 236071 374422 236083
rect 374474 236071 374480 236123
rect 376336 236071 376342 236123
rect 376394 236111 376400 236123
rect 376394 236083 406142 236111
rect 376394 236071 376400 236083
rect 208432 235997 208438 236049
rect 208490 236037 208496 236049
rect 223216 236037 223222 236049
rect 208490 236009 223222 236037
rect 208490 235997 208496 236009
rect 223216 235997 223222 236009
rect 223274 235997 223280 236049
rect 247984 235997 247990 236049
rect 248042 236037 248048 236049
rect 273616 236037 273622 236049
rect 248042 236009 273622 236037
rect 248042 235997 248048 236009
rect 273616 235997 273622 236009
rect 273674 235997 273680 236049
rect 276112 235997 276118 236049
rect 276170 236037 276176 236049
rect 308272 236037 308278 236049
rect 276170 236009 308278 236037
rect 276170 235997 276176 236009
rect 308272 235997 308278 236009
rect 308330 235997 308336 236049
rect 313840 235997 313846 236049
rect 313898 236037 313904 236049
rect 357136 236037 357142 236049
rect 313898 236009 357142 236037
rect 313898 235997 313904 236009
rect 357136 235997 357142 236009
rect 357194 235997 357200 236049
rect 371824 235997 371830 236049
rect 371882 236037 371888 236049
rect 406000 236037 406006 236049
rect 371882 236009 406006 236037
rect 371882 235997 371888 236009
rect 406000 235997 406006 236009
rect 406058 235997 406064 236049
rect 146992 235923 146998 235975
rect 147050 235963 147056 235975
rect 151216 235963 151222 235975
rect 147050 235935 151222 235963
rect 147050 235923 147056 235935
rect 151216 235923 151222 235935
rect 151274 235923 151280 235975
rect 207472 235923 207478 235975
rect 207530 235963 207536 235975
rect 223984 235963 223990 235975
rect 207530 235935 223990 235963
rect 207530 235923 207536 235935
rect 223984 235923 223990 235935
rect 224042 235923 224048 235975
rect 243280 235923 243286 235975
rect 243338 235963 243344 235975
rect 271024 235963 271030 235975
rect 243338 235935 271030 235963
rect 243338 235923 243344 235935
rect 271024 235923 271030 235935
rect 271082 235923 271088 235975
rect 280624 235923 280630 235975
rect 280682 235963 280688 235975
rect 320848 235963 320854 235975
rect 280682 235935 320854 235963
rect 280682 235923 280688 235935
rect 320848 235923 320854 235935
rect 320906 235923 320912 235975
rect 386704 235923 386710 235975
rect 386762 235963 386768 235975
rect 405616 235963 405622 235975
rect 386762 235935 405622 235963
rect 386762 235923 386768 235935
rect 405616 235923 405622 235935
rect 405674 235923 405680 235975
rect 406114 235963 406142 236083
rect 410032 236071 410038 236123
rect 410090 236111 410096 236123
rect 584560 236111 584566 236123
rect 410090 236083 584566 236111
rect 410090 236071 410096 236083
rect 584560 236071 584566 236083
rect 584618 236071 584624 236123
rect 406288 235997 406294 236049
rect 406346 236037 406352 236049
rect 415408 236037 415414 236049
rect 406346 236009 415414 236037
rect 406346 235997 406352 236009
rect 415408 235997 415414 236009
rect 415466 235997 415472 236049
rect 413872 235963 413878 235975
rect 406114 235935 413878 235963
rect 413872 235923 413878 235935
rect 413930 235923 413936 235975
rect 209680 235849 209686 235901
rect 209738 235889 209744 235901
rect 226192 235889 226198 235901
rect 209738 235861 226198 235889
rect 209738 235849 209744 235861
rect 226192 235849 226198 235861
rect 226250 235849 226256 235901
rect 234256 235849 234262 235901
rect 234314 235889 234320 235901
rect 264880 235889 264886 235901
rect 234314 235861 264886 235889
rect 234314 235849 234320 235861
rect 264880 235849 264886 235861
rect 264938 235849 264944 235901
rect 279280 235849 279286 235901
rect 279338 235889 279344 235901
rect 319600 235889 319606 235901
rect 279338 235861 319606 235889
rect 279338 235849 279344 235861
rect 319600 235849 319606 235861
rect 319658 235849 319664 235901
rect 326224 235849 326230 235901
rect 326282 235889 326288 235901
rect 460240 235889 460246 235901
rect 326282 235861 460246 235889
rect 326282 235849 326288 235861
rect 460240 235849 460246 235861
rect 460298 235849 460304 235901
rect 208912 235775 208918 235827
rect 208970 235815 208976 235827
rect 226960 235815 226966 235827
rect 208970 235787 226966 235815
rect 208970 235775 208976 235787
rect 226960 235775 226966 235787
rect 227018 235775 227024 235827
rect 237520 235775 237526 235827
rect 237578 235815 237584 235827
rect 268624 235815 268630 235827
rect 237578 235787 268630 235815
rect 237578 235775 237584 235787
rect 268624 235775 268630 235787
rect 268682 235775 268688 235827
rect 290320 235775 290326 235827
rect 290378 235815 290384 235827
rect 334096 235815 334102 235827
rect 290378 235787 334102 235815
rect 290378 235775 290384 235787
rect 334096 235775 334102 235787
rect 334154 235775 334160 235827
rect 343504 235775 343510 235827
rect 343562 235815 343568 235827
rect 495760 235815 495766 235827
rect 343562 235787 495766 235815
rect 343562 235775 343568 235787
rect 495760 235775 495766 235787
rect 495818 235775 495824 235827
rect 211216 235701 211222 235753
rect 211274 235741 211280 235753
rect 229264 235741 229270 235753
rect 211274 235713 229270 235741
rect 211274 235701 211280 235713
rect 229264 235701 229270 235713
rect 229322 235701 229328 235753
rect 231184 235701 231190 235753
rect 231242 235741 231248 235753
rect 259024 235741 259030 235753
rect 231242 235713 259030 235741
rect 231242 235701 231248 235713
rect 259024 235701 259030 235713
rect 259082 235701 259088 235753
rect 262864 235701 262870 235753
rect 262922 235741 262928 235753
rect 305104 235741 305110 235753
rect 262922 235713 305110 235741
rect 262922 235701 262928 235713
rect 305104 235701 305110 235713
rect 305162 235701 305168 235753
rect 317200 235701 317206 235753
rect 317258 235741 317264 235753
rect 410704 235741 410710 235753
rect 317258 235713 410710 235741
rect 317258 235701 317264 235713
rect 410704 235701 410710 235713
rect 410762 235701 410768 235753
rect 413680 235741 413686 235753
rect 410818 235713 413686 235741
rect 210640 235627 210646 235679
rect 210698 235667 210704 235679
rect 230032 235667 230038 235679
rect 210698 235639 230038 235667
rect 210698 235627 210704 235639
rect 230032 235627 230038 235639
rect 230090 235627 230096 235679
rect 239344 235627 239350 235679
rect 239402 235667 239408 235679
rect 287344 235667 287350 235679
rect 239402 235639 287350 235667
rect 239402 235627 239408 235639
rect 287344 235627 287350 235639
rect 287402 235627 287408 235679
rect 311152 235627 311158 235679
rect 311210 235667 311216 235679
rect 311210 235639 405566 235667
rect 311210 235627 311216 235639
rect 210064 235553 210070 235605
rect 210122 235593 210128 235605
rect 227824 235593 227830 235605
rect 210122 235565 227830 235593
rect 210122 235553 210128 235565
rect 227824 235553 227830 235565
rect 227882 235553 227888 235605
rect 236464 235553 236470 235605
rect 236522 235593 236528 235605
rect 282928 235593 282934 235605
rect 236522 235565 282934 235593
rect 236522 235553 236528 235565
rect 282928 235553 282934 235565
rect 282986 235553 282992 235605
rect 287056 235553 287062 235605
rect 287114 235593 287120 235605
rect 318160 235593 318166 235605
rect 287114 235565 318166 235593
rect 287114 235553 287120 235565
rect 318160 235553 318166 235565
rect 318218 235553 318224 235605
rect 358000 235553 358006 235605
rect 358058 235593 358064 235605
rect 400336 235593 400342 235605
rect 358058 235565 400342 235593
rect 358058 235553 358064 235565
rect 400336 235553 400342 235565
rect 400394 235553 400400 235605
rect 405538 235593 405566 235639
rect 405616 235627 405622 235679
rect 405674 235667 405680 235679
rect 410818 235667 410846 235713
rect 413680 235701 413686 235713
rect 413738 235701 413744 235753
rect 405674 235639 410846 235667
rect 405674 235627 405680 235639
rect 412144 235627 412150 235679
rect 412202 235667 412208 235679
rect 590416 235667 590422 235679
rect 412202 235639 590422 235667
rect 412202 235627 412208 235639
rect 590416 235627 590422 235639
rect 590474 235627 590480 235679
rect 408976 235593 408982 235605
rect 405538 235565 408982 235593
rect 408976 235553 408982 235565
rect 409034 235553 409040 235605
rect 409168 235553 409174 235605
rect 409226 235593 409232 235605
rect 588784 235593 588790 235605
rect 409226 235565 588790 235593
rect 409226 235553 409232 235565
rect 588784 235553 588790 235565
rect 588842 235553 588848 235605
rect 212944 235479 212950 235531
rect 213002 235519 213008 235531
rect 232336 235519 232342 235531
rect 213002 235491 232342 235519
rect 213002 235479 213008 235491
rect 232336 235479 232342 235491
rect 232394 235479 232400 235531
rect 238000 235479 238006 235531
rect 238058 235519 238064 235531
rect 285904 235519 285910 235531
rect 238058 235491 285910 235519
rect 238058 235479 238064 235491
rect 285904 235479 285910 235491
rect 285962 235479 285968 235531
rect 299824 235479 299830 235531
rect 299882 235519 299888 235531
rect 354256 235519 354262 235531
rect 299882 235491 354262 235519
rect 299882 235479 299888 235491
rect 354256 235479 354262 235491
rect 354314 235479 354320 235531
rect 394960 235479 394966 235531
rect 395018 235519 395024 235531
rect 587344 235519 587350 235531
rect 395018 235491 587350 235519
rect 395018 235479 395024 235491
rect 587344 235479 587350 235491
rect 587402 235479 587408 235531
rect 211984 235405 211990 235457
rect 212042 235445 212048 235457
rect 233008 235445 233014 235457
rect 212042 235417 233014 235445
rect 212042 235405 212048 235417
rect 233008 235405 233014 235417
rect 233066 235405 233072 235457
rect 242128 235405 242134 235457
rect 242186 235445 242192 235457
rect 293392 235445 293398 235457
rect 242186 235417 293398 235445
rect 242186 235405 242192 235417
rect 293392 235405 293398 235417
rect 293450 235405 293456 235457
rect 294832 235405 294838 235457
rect 294890 235445 294896 235457
rect 337648 235445 337654 235457
rect 294890 235417 337654 235445
rect 294890 235405 294896 235417
rect 337648 235405 337654 235417
rect 337706 235405 337712 235457
rect 339472 235405 339478 235457
rect 339530 235445 339536 235457
rect 395056 235445 395062 235457
rect 339530 235417 395062 235445
rect 339530 235405 339536 235417
rect 395056 235405 395062 235417
rect 395114 235405 395120 235457
rect 396784 235405 396790 235457
rect 396842 235445 396848 235457
rect 587632 235445 587638 235457
rect 396842 235417 587638 235445
rect 396842 235405 396848 235417
rect 587632 235405 587638 235417
rect 587690 235405 587696 235457
rect 206992 235331 206998 235383
rect 207050 235371 207056 235383
rect 221776 235371 221782 235383
rect 207050 235343 221782 235371
rect 207050 235331 207056 235343
rect 221776 235331 221782 235343
rect 221834 235331 221840 235383
rect 223888 235331 223894 235383
rect 223946 235371 223952 235383
rect 244720 235371 244726 235383
rect 223946 235343 244726 235371
rect 223946 235331 223952 235343
rect 244720 235331 244726 235343
rect 244778 235331 244784 235383
rect 249712 235331 249718 235383
rect 249770 235371 249776 235383
rect 302320 235371 302326 235383
rect 249770 235343 302326 235371
rect 249770 235331 249776 235343
rect 302320 235331 302326 235343
rect 302378 235331 302384 235383
rect 304816 235331 304822 235383
rect 304874 235371 304880 235383
rect 362608 235371 362614 235383
rect 304874 235343 362614 235371
rect 304874 235331 304880 235343
rect 362608 235331 362614 235343
rect 362666 235331 362672 235383
rect 393424 235331 393430 235383
rect 393482 235371 393488 235383
rect 587056 235371 587062 235383
rect 393482 235343 587062 235371
rect 393482 235331 393488 235343
rect 587056 235331 587062 235343
rect 587114 235331 587120 235383
rect 214192 235257 214198 235309
rect 214250 235297 214256 235309
rect 235312 235297 235318 235309
rect 214250 235269 235318 235297
rect 214250 235257 214256 235269
rect 235312 235257 235318 235269
rect 235370 235257 235376 235309
rect 288880 235257 288886 235309
rect 288938 235297 288944 235309
rect 346864 235297 346870 235309
rect 288938 235269 346870 235297
rect 288938 235257 288944 235269
rect 346864 235257 346870 235269
rect 346922 235257 346928 235309
rect 392176 235257 392182 235309
rect 392234 235297 392240 235309
rect 585520 235297 585526 235309
rect 392234 235269 585526 235297
rect 392234 235257 392240 235269
rect 585520 235257 585526 235269
rect 585578 235257 585584 235309
rect 209296 235183 209302 235235
rect 209354 235223 209360 235235
rect 228496 235223 228502 235235
rect 209354 235195 228502 235223
rect 209354 235183 209360 235195
rect 228496 235183 228502 235195
rect 228554 235183 228560 235235
rect 229744 235183 229750 235235
rect 229802 235223 229808 235235
rect 253552 235223 253558 235235
rect 229802 235195 253558 235223
rect 229802 235183 229808 235195
rect 253552 235183 253558 235195
rect 253610 235183 253616 235235
rect 257488 235183 257494 235235
rect 257546 235223 257552 235235
rect 308176 235223 308182 235235
rect 257546 235195 308182 235223
rect 257546 235183 257552 235195
rect 308176 235183 308182 235195
rect 308234 235183 308240 235235
rect 334960 235183 334966 235235
rect 335018 235223 335024 235235
rect 391696 235223 391702 235235
rect 335018 235195 391702 235223
rect 335018 235183 335024 235195
rect 391696 235183 391702 235195
rect 391754 235183 391760 235235
rect 396304 235183 396310 235235
rect 396362 235223 396368 235235
rect 588592 235223 588598 235235
rect 396362 235195 588598 235223
rect 396362 235183 396368 235195
rect 588592 235183 588598 235195
rect 588650 235183 588656 235235
rect 211600 235109 211606 235161
rect 211658 235149 211664 235161
rect 230704 235149 230710 235161
rect 211658 235121 230710 235149
rect 211658 235109 211664 235121
rect 230704 235109 230710 235121
rect 230762 235109 230768 235161
rect 232912 235109 232918 235161
rect 232970 235149 232976 235161
rect 262000 235149 262006 235161
rect 232970 235121 262006 235149
rect 232970 235109 232976 235121
rect 262000 235109 262006 235121
rect 262058 235109 262064 235161
rect 266128 235109 266134 235161
rect 266186 235149 266192 235161
rect 324208 235149 324214 235161
rect 266186 235121 324214 235149
rect 266186 235109 266192 235121
rect 324208 235109 324214 235121
rect 324266 235109 324272 235161
rect 332176 235109 332182 235161
rect 332234 235149 332240 235161
rect 385360 235149 385366 235161
rect 332234 235121 385366 235149
rect 332234 235109 332240 235121
rect 385360 235109 385366 235121
rect 385418 235109 385424 235161
rect 387664 235109 387670 235161
rect 387722 235149 387728 235161
rect 583408 235149 583414 235161
rect 387722 235121 583414 235149
rect 387722 235109 387728 235121
rect 583408 235109 583414 235121
rect 583466 235109 583472 235161
rect 207856 235035 207862 235087
rect 207914 235075 207920 235087
rect 215920 235075 215926 235087
rect 207914 235047 215926 235075
rect 207914 235035 207920 235047
rect 215920 235035 215926 235047
rect 215978 235035 215984 235087
rect 220624 235035 220630 235087
rect 220682 235075 220688 235087
rect 241840 235075 241846 235087
rect 220682 235047 241846 235075
rect 220682 235035 220688 235047
rect 241840 235035 241846 235047
rect 241898 235035 241904 235087
rect 246640 235035 246646 235087
rect 246698 235075 246704 235087
rect 299248 235075 299254 235087
rect 246698 235047 299254 235075
rect 246698 235035 246704 235047
rect 299248 235035 299254 235047
rect 299306 235035 299312 235087
rect 309328 235035 309334 235087
rect 309386 235075 309392 235087
rect 368848 235075 368854 235087
rect 309386 235047 368854 235075
rect 309386 235035 309392 235047
rect 368848 235035 368854 235047
rect 368906 235035 368912 235087
rect 394864 235035 394870 235087
rect 394922 235075 394928 235087
rect 596080 235075 596086 235087
rect 394922 235047 596086 235075
rect 394922 235035 394928 235047
rect 596080 235035 596086 235047
rect 596138 235035 596144 235087
rect 211024 234961 211030 235013
rect 211082 235001 211088 235013
rect 231568 235001 231574 235013
rect 211082 234973 231574 235001
rect 211082 234961 211088 234973
rect 231568 234961 231574 234973
rect 231626 234961 231632 235013
rect 243856 234961 243862 235013
rect 243914 235001 243920 235013
rect 296464 235001 296470 235013
rect 243914 234973 296470 235001
rect 243914 234961 243920 234973
rect 296464 234961 296470 234973
rect 296522 234961 296528 235013
rect 298000 234961 298006 235013
rect 298058 235001 298064 235013
rect 362416 235001 362422 235013
rect 298058 234973 362422 235001
rect 298058 234961 298064 234973
rect 362416 234961 362422 234973
rect 362474 234961 362480 235013
rect 362512 234961 362518 235013
rect 362570 235001 362576 235013
rect 394672 235001 394678 235013
rect 362570 234973 394678 235001
rect 362570 234961 362576 234973
rect 394672 234961 394678 234973
rect 394730 234961 394736 235013
rect 398992 234961 398998 235013
rect 399050 235001 399056 235013
rect 605968 235001 605974 235013
rect 399050 234973 605974 235001
rect 399050 234961 399056 234973
rect 605968 234961 605974 234973
rect 606026 234961 606032 235013
rect 213424 234887 213430 234939
rect 213482 234927 213488 234939
rect 213482 234899 225470 234927
rect 213482 234887 213488 234899
rect 208720 234813 208726 234865
rect 208778 234853 208784 234865
rect 224752 234853 224758 234865
rect 208778 234825 224758 234853
rect 208778 234813 208784 234825
rect 224752 234813 224758 234825
rect 224810 234813 224816 234865
rect 204400 234739 204406 234791
rect 204458 234779 204464 234791
rect 215824 234779 215830 234791
rect 204458 234751 215830 234779
rect 204458 234739 204464 234751
rect 215824 234739 215830 234751
rect 215882 234739 215888 234791
rect 225442 234779 225470 234899
rect 235696 234887 235702 234939
rect 235754 234927 235760 234939
rect 266896 234927 266902 234939
rect 235754 234899 266902 234927
rect 235754 234887 235760 234899
rect 266896 234887 266902 234899
rect 266954 234887 266960 234939
rect 268912 234887 268918 234939
rect 268970 234927 268976 234939
rect 331408 234927 331414 234939
rect 268970 234899 331414 234927
rect 268970 234887 268976 234899
rect 331408 234887 331414 234899
rect 331466 234887 331472 234939
rect 333424 234887 333430 234939
rect 333482 234927 333488 234939
rect 394768 234927 394774 234939
rect 333482 234899 394774 234927
rect 333482 234887 333488 234899
rect 394768 234887 394774 234899
rect 394826 234887 394832 234939
rect 398608 234887 398614 234939
rect 398666 234927 398672 234939
rect 605296 234927 605302 234939
rect 398666 234899 605302 234927
rect 398666 234887 398672 234899
rect 605296 234887 605302 234899
rect 605354 234887 605360 234939
rect 225520 234813 225526 234865
rect 225578 234853 225584 234865
rect 260176 234853 260182 234865
rect 225578 234825 260182 234853
rect 225578 234813 225584 234825
rect 260176 234813 260182 234825
rect 260234 234813 260240 234865
rect 260272 234813 260278 234865
rect 260330 234853 260336 234865
rect 323056 234853 323062 234865
rect 260330 234825 323062 234853
rect 260330 234813 260336 234825
rect 323056 234813 323062 234825
rect 323114 234813 323120 234865
rect 327664 234813 327670 234865
rect 327722 234853 327728 234865
rect 392464 234853 392470 234865
rect 327722 234825 392470 234853
rect 327722 234813 327728 234825
rect 392464 234813 392470 234825
rect 392522 234813 392528 234865
rect 403600 234813 403606 234865
rect 403658 234853 403664 234865
rect 615856 234853 615862 234865
rect 403658 234825 615862 234853
rect 403658 234813 403664 234825
rect 615856 234813 615862 234825
rect 615914 234813 615920 234865
rect 236080 234779 236086 234791
rect 225442 234751 236086 234779
rect 236080 234739 236086 234751
rect 236138 234739 236144 234791
rect 254224 234739 254230 234791
rect 254282 234779 254288 234791
rect 306640 234779 306646 234791
rect 254282 234751 306646 234779
rect 254282 234739 254288 234751
rect 306640 234739 306646 234751
rect 306698 234739 306704 234791
rect 321616 234739 321622 234791
rect 321674 234779 321680 234791
rect 387280 234779 387286 234791
rect 321674 234751 387286 234779
rect 321674 234739 321680 234751
rect 387280 234739 387286 234751
rect 387338 234739 387344 234791
rect 406672 234739 406678 234791
rect 406730 234779 406736 234791
rect 621808 234779 621814 234791
rect 406730 234751 621814 234779
rect 406730 234739 406736 234751
rect 621808 234739 621814 234751
rect 621866 234739 621872 234791
rect 202864 234665 202870 234717
rect 202922 234705 202928 234717
rect 214864 234705 214870 234717
rect 202922 234677 214870 234705
rect 202922 234665 202928 234677
rect 214864 234665 214870 234677
rect 214922 234665 214928 234717
rect 225136 234665 225142 234717
rect 225194 234705 225200 234717
rect 247696 234705 247702 234717
rect 225194 234677 247702 234705
rect 225194 234665 225200 234677
rect 247696 234665 247702 234677
rect 247754 234665 247760 234717
rect 251152 234665 251158 234717
rect 251210 234705 251216 234717
rect 304144 234705 304150 234717
rect 251210 234677 304150 234705
rect 251210 234665 251216 234677
rect 304144 234665 304150 234677
rect 304202 234665 304208 234717
rect 315280 234665 315286 234717
rect 315338 234705 315344 234717
rect 394672 234705 394678 234717
rect 315338 234677 394678 234705
rect 315338 234665 315344 234677
rect 394672 234665 394678 234677
rect 394730 234665 394736 234717
rect 408112 234665 408118 234717
rect 408170 234705 408176 234717
rect 624880 234705 624886 234717
rect 408170 234677 624886 234705
rect 408170 234665 408176 234677
rect 624880 234665 624886 234677
rect 624938 234665 624944 234717
rect 204784 234591 204790 234643
rect 204842 234631 204848 234643
rect 204842 234603 213662 234631
rect 204842 234591 204848 234603
rect 202000 234517 202006 234569
rect 202058 234557 202064 234569
rect 213424 234557 213430 234569
rect 202058 234529 213430 234557
rect 202058 234517 202064 234529
rect 213424 234517 213430 234529
rect 213482 234517 213488 234569
rect 203248 234443 203254 234495
rect 203306 234483 203312 234495
rect 207760 234483 207766 234495
rect 203306 234455 207766 234483
rect 203306 234443 203312 234455
rect 207760 234443 207766 234455
rect 207818 234443 207824 234495
rect 206128 234369 206134 234421
rect 206186 234409 206192 234421
rect 213634 234409 213662 234603
rect 222352 234591 222358 234643
rect 222410 234631 222416 234643
rect 222410 234603 227534 234631
rect 222410 234591 222416 234603
rect 227506 234557 227534 234603
rect 240208 234591 240214 234643
rect 240266 234631 240272 234643
rect 264688 234631 264694 234643
rect 240266 234603 264694 234631
rect 240266 234591 240272 234603
rect 264688 234591 264694 234603
rect 264746 234591 264752 234643
rect 267472 234591 267478 234643
rect 267530 234631 267536 234643
rect 285040 234631 285046 234643
rect 267530 234603 285046 234631
rect 267530 234591 267536 234603
rect 285040 234591 285046 234603
rect 285098 234591 285104 234643
rect 286672 234591 286678 234643
rect 286730 234631 286736 234643
rect 326800 234631 326806 234643
rect 286730 234603 326806 234631
rect 286730 234591 286736 234603
rect 326800 234591 326806 234603
rect 326858 234591 326864 234643
rect 329296 234591 329302 234643
rect 329354 234631 329360 234643
rect 449296 234631 449302 234643
rect 329354 234603 449302 234631
rect 329354 234591 329360 234603
rect 449296 234591 449302 234603
rect 449354 234591 449360 234643
rect 243952 234557 243958 234569
rect 227506 234529 243958 234557
rect 243952 234517 243958 234529
rect 244010 234517 244016 234569
rect 250576 234557 250582 234569
rect 247666 234529 250582 234557
rect 215920 234443 215926 234495
rect 215978 234483 215984 234495
rect 225520 234483 225526 234495
rect 215978 234455 225526 234483
rect 215978 234443 215984 234455
rect 225520 234443 225526 234455
rect 225578 234443 225584 234495
rect 235600 234443 235606 234495
rect 235658 234483 235664 234495
rect 247666 234483 247694 234529
rect 250576 234517 250582 234529
rect 250634 234517 250640 234569
rect 255280 234517 255286 234569
rect 255338 234557 255344 234569
rect 278224 234557 278230 234569
rect 255338 234529 278230 234557
rect 255338 234517 255344 234529
rect 278224 234517 278230 234529
rect 278282 234517 278288 234569
rect 283888 234517 283894 234569
rect 283946 234557 283952 234569
rect 320656 234557 320662 234569
rect 283946 234529 320662 234557
rect 283946 234517 283952 234529
rect 320656 234517 320662 234529
rect 320714 234517 320720 234569
rect 323536 234517 323542 234569
rect 323594 234557 323600 234569
rect 434896 234557 434902 234569
rect 323594 234529 434902 234557
rect 323594 234517 323600 234529
rect 434896 234517 434902 234529
rect 434954 234517 434960 234569
rect 235658 234455 247694 234483
rect 235658 234443 235664 234455
rect 250480 234443 250486 234495
rect 250538 234483 250544 234495
rect 267952 234483 267958 234495
rect 250538 234455 267958 234483
rect 250538 234443 250544 234455
rect 267952 234443 267958 234455
rect 268010 234443 268016 234495
rect 273040 234443 273046 234495
rect 273098 234483 273104 234495
rect 304720 234483 304726 234495
rect 273098 234455 304726 234483
rect 273098 234443 273104 234455
rect 304720 234443 304726 234455
rect 304778 234443 304784 234495
rect 313840 234483 313846 234495
rect 306658 234455 313846 234483
rect 219376 234409 219382 234421
rect 206186 234381 211358 234409
rect 213634 234381 219382 234409
rect 206186 234369 206192 234381
rect 206512 234295 206518 234347
rect 206570 234335 206576 234347
rect 211330 234335 211358 234381
rect 219376 234369 219382 234381
rect 219434 234369 219440 234421
rect 237040 234369 237046 234421
rect 237098 234409 237104 234421
rect 258064 234409 258070 234421
rect 237098 234381 258070 234409
rect 237098 234369 237104 234381
rect 258064 234369 258070 234381
rect 258122 234369 258128 234421
rect 262480 234369 262486 234421
rect 262538 234409 262544 234421
rect 290896 234409 290902 234421
rect 262538 234381 290902 234409
rect 262538 234369 262544 234381
rect 290896 234369 290902 234381
rect 290954 234369 290960 234421
rect 292912 234369 292918 234421
rect 292970 234409 292976 234421
rect 306658 234409 306686 234455
rect 313840 234443 313846 234455
rect 313898 234443 313904 234495
rect 314416 234443 314422 234495
rect 314474 234483 314480 234495
rect 426160 234483 426166 234495
rect 314474 234455 426166 234483
rect 314474 234443 314480 234455
rect 426160 234443 426166 234455
rect 426218 234443 426224 234495
rect 292970 234381 306686 234409
rect 292970 234369 292976 234381
rect 312688 234369 312694 234421
rect 312746 234409 312752 234421
rect 407440 234409 407446 234421
rect 312746 234381 407446 234409
rect 312746 234369 312752 234381
rect 407440 234369 407446 234381
rect 407498 234369 407504 234421
rect 408976 234369 408982 234421
rect 409034 234409 409040 234421
rect 410608 234409 410614 234421
rect 409034 234381 410614 234409
rect 409034 234369 409040 234381
rect 410608 234369 410614 234381
rect 410666 234369 410672 234421
rect 221008 234335 221014 234347
rect 206570 234307 211262 234335
rect 211330 234307 221014 234335
rect 206570 234295 206576 234307
rect 200272 234221 200278 234273
rect 200330 234261 200336 234273
rect 210352 234261 210358 234273
rect 200330 234233 210358 234261
rect 200330 234221 200336 234233
rect 210352 234221 210358 234233
rect 210410 234221 210416 234273
rect 211234 234261 211262 234307
rect 221008 234295 221014 234307
rect 221066 234295 221072 234347
rect 239824 234295 239830 234347
rect 239882 234335 239888 234347
rect 260464 234335 260470 234347
rect 239882 234307 260470 234335
rect 239882 234295 239888 234307
rect 260464 234295 260470 234307
rect 260522 234295 260528 234347
rect 271600 234295 271606 234347
rect 271658 234335 271664 234347
rect 302224 234335 302230 234347
rect 271658 234307 302230 234335
rect 271658 234295 271664 234307
rect 302224 234295 302230 234307
rect 302282 234295 302288 234347
rect 308464 234295 308470 234347
rect 308522 234335 308528 234347
rect 414736 234335 414742 234347
rect 308522 234307 414742 234335
rect 308522 234295 308528 234307
rect 414736 234295 414742 234307
rect 414794 234295 414800 234347
rect 222448 234261 222454 234273
rect 211234 234233 222454 234261
rect 222448 234221 222454 234233
rect 222506 234221 222512 234273
rect 242896 234221 242902 234273
rect 242954 234261 242960 234273
rect 260752 234261 260758 234273
rect 242954 234233 260758 234261
rect 242954 234221 242960 234233
rect 260752 234221 260758 234233
rect 260810 234221 260816 234273
rect 261232 234221 261238 234273
rect 261290 234261 261296 234273
rect 288016 234261 288022 234273
rect 261290 234233 288022 234261
rect 261290 234221 261296 234233
rect 288016 234221 288022 234233
rect 288074 234221 288080 234273
rect 295216 234221 295222 234273
rect 295274 234261 295280 234273
rect 348688 234261 348694 234273
rect 295274 234233 348694 234261
rect 295274 234221 295280 234233
rect 348688 234221 348694 234233
rect 348746 234221 348752 234273
rect 352144 234221 352150 234273
rect 352202 234261 352208 234273
rect 401104 234261 401110 234273
rect 352202 234233 401110 234261
rect 352202 234221 352208 234233
rect 401104 234221 401110 234233
rect 401162 234221 401168 234273
rect 407248 234221 407254 234273
rect 407306 234261 407312 234273
rect 503920 234261 503926 234273
rect 407306 234233 503926 234261
rect 407306 234221 407312 234233
rect 503920 234221 503926 234233
rect 503978 234221 503984 234273
rect 200176 234147 200182 234199
rect 200234 234187 200240 234199
rect 208816 234187 208822 234199
rect 200234 234159 208822 234187
rect 200234 234147 200240 234159
rect 208816 234147 208822 234159
rect 208874 234147 208880 234199
rect 256528 234147 256534 234199
rect 256586 234187 256592 234199
rect 278032 234187 278038 234199
rect 256586 234159 278038 234187
rect 256586 234147 256592 234159
rect 278032 234147 278038 234159
rect 278090 234147 278096 234199
rect 283984 234147 283990 234199
rect 284042 234187 284048 234199
rect 311248 234187 311254 234199
rect 284042 234159 311254 234187
rect 284042 234147 284048 234159
rect 311248 234147 311254 234159
rect 311306 234147 311312 234199
rect 318352 234147 318358 234199
rect 318410 234187 318416 234199
rect 371632 234187 371638 234199
rect 318410 234159 371638 234187
rect 318410 234147 318416 234159
rect 371632 234147 371638 234159
rect 371690 234147 371696 234199
rect 378544 234147 378550 234199
rect 378602 234187 378608 234199
rect 399184 234187 399190 234199
rect 378602 234159 399190 234187
rect 378602 234147 378608 234159
rect 399184 234147 399190 234159
rect 399242 234147 399248 234199
rect 403504 234147 403510 234199
rect 403562 234187 403568 234199
rect 495376 234187 495382 234199
rect 403562 234159 495382 234187
rect 403562 234147 403568 234159
rect 495376 234147 495382 234159
rect 495434 234147 495440 234199
rect 198736 234073 198742 234125
rect 198794 234113 198800 234125
rect 207376 234113 207382 234125
rect 198794 234085 207382 234113
rect 198794 234073 198800 234085
rect 207376 234073 207382 234085
rect 207434 234073 207440 234125
rect 207760 234073 207766 234125
rect 207818 234113 207824 234125
rect 216496 234113 216502 234125
rect 207818 234085 216502 234113
rect 207818 234073 207824 234085
rect 216496 234073 216502 234085
rect 216554 234073 216560 234125
rect 244336 234073 244342 234125
rect 244394 234113 244400 234125
rect 263824 234113 263830 234125
rect 244394 234085 263830 234113
rect 244394 234073 244400 234085
rect 263824 234073 263830 234085
rect 263882 234073 263888 234125
rect 268528 234073 268534 234125
rect 268586 234113 268592 234125
rect 293776 234113 293782 234125
rect 268586 234085 293782 234113
rect 268586 234073 268592 234085
rect 293776 234073 293782 234085
rect 293834 234073 293840 234125
rect 295696 234073 295702 234125
rect 295754 234113 295760 234125
rect 341200 234113 341206 234125
rect 295754 234085 341206 234113
rect 295754 234073 295760 234085
rect 341200 234073 341206 234085
rect 341258 234073 341264 234125
rect 345904 234073 345910 234125
rect 345962 234113 345968 234125
rect 400144 234113 400150 234125
rect 345962 234085 400150 234113
rect 345962 234073 345968 234085
rect 400144 234073 400150 234085
rect 400202 234073 400208 234125
rect 401776 234073 401782 234125
rect 401834 234113 401840 234125
rect 484624 234113 484630 234125
rect 401834 234085 484630 234113
rect 401834 234073 401840 234085
rect 484624 234073 484630 234085
rect 484682 234073 484688 234125
rect 198352 233999 198358 234051
rect 198410 234039 198416 234051
rect 205936 234039 205942 234051
rect 198410 234011 205942 234039
rect 198410 233999 198416 234011
rect 205936 233999 205942 234011
rect 205994 233999 206000 234051
rect 218704 234039 218710 234051
rect 206818 234011 218710 234039
rect 197488 233925 197494 233977
rect 197546 233965 197552 233977
rect 204304 233965 204310 233977
rect 197546 233937 204310 233965
rect 197546 233925 197552 233937
rect 204304 233925 204310 233937
rect 204362 233925 204368 233977
rect 205552 233925 205558 233977
rect 205610 233965 205616 233977
rect 206818 233965 206846 234011
rect 218704 233999 218710 234011
rect 218762 233999 218768 234051
rect 247408 233999 247414 234051
rect 247466 234039 247472 234051
rect 266320 234039 266326 234051
rect 247466 234011 266326 234039
rect 247466 233999 247472 234011
rect 266320 233999 266326 234011
rect 266378 233999 266384 234051
rect 267088 233999 267094 234051
rect 267146 234039 267152 234051
rect 290992 234039 290998 234051
rect 267146 234011 290998 234039
rect 267146 233999 267152 234011
rect 290992 233999 290998 234011
rect 291050 233999 291056 234051
rect 301648 233999 301654 234051
rect 301706 234039 301712 234051
rect 344080 234039 344086 234051
rect 301706 234011 344086 234039
rect 301706 233999 301712 234011
rect 344080 233999 344086 234011
rect 344138 233999 344144 234051
rect 344368 233999 344374 234051
rect 344426 234039 344432 234051
rect 394864 234039 394870 234051
rect 344426 234011 394870 234039
rect 344426 233999 344432 234011
rect 394864 233999 394870 234011
rect 394922 233999 394928 234051
rect 396688 233999 396694 234051
rect 396746 234039 396752 234051
rect 475216 234039 475222 234051
rect 396746 234011 475222 234039
rect 396746 233999 396752 234011
rect 475216 233999 475222 234011
rect 475274 233999 475280 234051
rect 205610 233937 206846 233965
rect 205610 233925 205616 233937
rect 206896 233925 206902 233977
rect 206954 233965 206960 233977
rect 220240 233965 220246 233977
rect 206954 233937 220246 233965
rect 206954 233925 206960 233937
rect 220240 233925 220246 233937
rect 220298 233925 220304 233977
rect 259792 233925 259798 233977
rect 259850 233965 259856 233977
rect 281488 233965 281494 233977
rect 259850 233937 281494 233965
rect 259850 233925 259856 233937
rect 281488 233925 281494 233937
rect 281546 233925 281552 233977
rect 305200 233925 305206 233977
rect 305258 233965 305264 233977
rect 351376 233965 351382 233977
rect 305258 233937 351382 233965
rect 305258 233925 305264 233937
rect 351376 233925 351382 233937
rect 351434 233925 351440 233977
rect 361264 233925 361270 233977
rect 361322 233965 361328 233977
rect 432016 233965 432022 233977
rect 361322 233937 432022 233965
rect 361322 233925 361328 233937
rect 432016 233925 432022 233937
rect 432074 233925 432080 233977
rect 199120 233851 199126 233903
rect 199178 233891 199184 233903
rect 205072 233891 205078 233903
rect 199178 233863 205078 233891
rect 199178 233851 199184 233863
rect 205072 233851 205078 233863
rect 205130 233851 205136 233903
rect 205168 233851 205174 233903
rect 205226 233891 205232 233903
rect 205226 233863 215678 233891
rect 205226 233851 205232 233863
rect 196912 233777 196918 233829
rect 196970 233817 196976 233829
rect 202864 233817 202870 233829
rect 196970 233789 202870 233817
rect 196970 233777 196976 233789
rect 202864 233777 202870 233789
rect 202922 233777 202928 233829
rect 204208 233777 204214 233829
rect 204266 233817 204272 233829
rect 215536 233817 215542 233829
rect 204266 233789 215542 233817
rect 204266 233777 204272 233789
rect 215536 233777 215542 233789
rect 215594 233777 215600 233829
rect 196528 233703 196534 233755
rect 196586 233743 196592 233755
rect 200560 233743 200566 233755
rect 196586 233715 200566 233743
rect 196586 233703 196592 233715
rect 200560 233703 200566 233715
rect 200618 233703 200624 233755
rect 201520 233703 201526 233755
rect 201578 233743 201584 233755
rect 211888 233743 211894 233755
rect 201578 233715 211894 233743
rect 201578 233703 201584 233715
rect 211888 233703 211894 233715
rect 211946 233703 211952 233755
rect 195664 233629 195670 233681
rect 195722 233669 195728 233681
rect 201328 233669 201334 233681
rect 195722 233641 201334 233669
rect 195722 233629 195728 233641
rect 201328 233629 201334 233641
rect 201386 233629 201392 233681
rect 202480 233629 202486 233681
rect 202538 233669 202544 233681
rect 212560 233669 212566 233681
rect 202538 233641 212566 233669
rect 202538 233629 202544 233641
rect 212560 233629 212566 233641
rect 212618 233629 212624 233681
rect 215650 233669 215678 233863
rect 258352 233851 258358 233903
rect 258410 233891 258416 233903
rect 278704 233891 278710 233903
rect 258410 233863 278710 233891
rect 258410 233851 258416 233863
rect 278704 233851 278710 233863
rect 278762 233851 278768 233903
rect 296080 233851 296086 233903
rect 296138 233891 296144 233903
rect 339760 233891 339766 233903
rect 296138 233863 339766 233891
rect 296138 233851 296144 233863
rect 339760 233851 339766 233863
rect 339818 233851 339824 233903
rect 370288 233851 370294 233903
rect 370346 233891 370352 233903
rect 427888 233891 427894 233903
rect 370346 233863 427894 233891
rect 370346 233851 370352 233863
rect 427888 233851 427894 233863
rect 427946 233851 427952 233903
rect 215824 233777 215830 233829
rect 215882 233817 215888 233829
rect 217936 233817 217942 233829
rect 215882 233789 217942 233817
rect 215882 233777 215888 233789
rect 217936 233777 217942 233789
rect 217994 233777 218000 233829
rect 253456 233777 253462 233829
rect 253514 233817 253520 233829
rect 270832 233817 270838 233829
rect 253514 233789 270838 233817
rect 253514 233777 253520 233789
rect 270832 233777 270838 233789
rect 270890 233777 270896 233829
rect 294448 233777 294454 233829
rect 294506 233817 294512 233829
rect 331216 233817 331222 233829
rect 294506 233789 331222 233817
rect 294506 233777 294512 233789
rect 331216 233777 331222 233789
rect 331274 233777 331280 233829
rect 354928 233777 354934 233829
rect 354986 233817 354992 233829
rect 354986 233789 397454 233817
rect 354986 233777 354992 233789
rect 285136 233703 285142 233755
rect 285194 233743 285200 233755
rect 323152 233743 323158 233755
rect 285194 233715 323158 233743
rect 285194 233703 285200 233715
rect 323152 233703 323158 233715
rect 323210 233703 323216 233755
rect 338032 233703 338038 233755
rect 338090 233743 338096 233755
rect 386224 233743 386230 233755
rect 338090 233715 386230 233743
rect 338090 233703 338096 233715
rect 386224 233703 386230 233715
rect 386282 233703 386288 233755
rect 397426 233743 397454 233789
rect 398224 233777 398230 233829
rect 398282 233817 398288 233829
rect 405808 233817 405814 233829
rect 398282 233789 405814 233817
rect 398282 233777 398288 233789
rect 405808 233777 405814 233789
rect 405866 233777 405872 233829
rect 407440 233777 407446 233829
rect 407498 233817 407504 233829
rect 423280 233817 423286 233829
rect 407498 233789 423286 233817
rect 407498 233777 407504 233789
rect 423280 233777 423286 233789
rect 423338 233777 423344 233829
rect 407536 233743 407542 233755
rect 397426 233715 407542 233743
rect 407536 233703 407542 233715
rect 407594 233703 407600 233755
rect 217168 233669 217174 233681
rect 215650 233641 217174 233669
rect 217168 233629 217174 233641
rect 217226 233629 217232 233681
rect 306256 233629 306262 233681
rect 306314 233669 306320 233681
rect 344464 233669 344470 233681
rect 306314 233641 344470 233669
rect 306314 233629 306320 233641
rect 344464 233629 344470 233641
rect 344522 233629 344528 233681
rect 363472 233629 363478 233681
rect 363530 233669 363536 233681
rect 364144 233669 364150 233681
rect 363530 233641 364150 233669
rect 363530 233629 363536 233641
rect 364144 233629 364150 233641
rect 364202 233629 364208 233681
rect 383632 233629 383638 233681
rect 383690 233669 383696 233681
rect 408112 233669 408118 233681
rect 383690 233641 408118 233669
rect 383690 233629 383696 233641
rect 408112 233629 408118 233641
rect 408170 233629 408176 233681
rect 192880 233555 192886 233607
rect 192938 233595 192944 233607
rect 195280 233595 195286 233607
rect 192938 233567 195286 233595
rect 192938 233555 192944 233567
rect 195280 233555 195286 233567
rect 195338 233555 195344 233607
rect 195568 233555 195574 233607
rect 195626 233595 195632 233607
rect 199792 233595 199798 233607
rect 195626 233567 199798 233595
rect 195626 233555 195632 233567
rect 199792 233555 199798 233567
rect 199850 233555 199856 233607
rect 201040 233555 201046 233607
rect 201098 233595 201104 233607
rect 209680 233595 209686 233607
rect 201098 233567 209686 233595
rect 201098 233555 201104 233567
rect 209680 233555 209686 233567
rect 209738 233555 209744 233607
rect 228400 233555 228406 233607
rect 228458 233595 228464 233607
rect 238096 233595 238102 233607
rect 228458 233567 238102 233595
rect 228458 233555 228464 233567
rect 238096 233555 238102 233567
rect 238154 233555 238160 233607
rect 259888 233555 259894 233607
rect 259946 233595 259952 233607
rect 267760 233595 267766 233607
rect 259946 233567 267766 233595
rect 259946 233555 259952 233567
rect 267760 233555 267766 233567
rect 267818 233555 267824 233607
rect 302896 233555 302902 233607
rect 302954 233595 302960 233607
rect 337360 233595 337366 233607
rect 302954 233567 337366 233595
rect 302954 233555 302960 233567
rect 337360 233555 337366 233567
rect 337418 233555 337424 233607
rect 348880 233555 348886 233607
rect 348938 233595 348944 233607
rect 394576 233595 394582 233607
rect 348938 233567 394582 233595
rect 348938 233555 348944 233567
rect 394576 233555 394582 233567
rect 394634 233555 394640 233607
rect 194224 233481 194230 233533
rect 194282 233521 194288 233533
rect 198352 233521 198358 233533
rect 194282 233493 198358 233521
rect 194282 233481 194288 233493
rect 198352 233481 198358 233493
rect 198410 233481 198416 233533
rect 200656 233481 200662 233533
rect 200714 233521 200720 233533
rect 208144 233521 208150 233533
rect 200714 233493 208150 233521
rect 200714 233481 200720 233493
rect 208144 233481 208150 233493
rect 208202 233481 208208 233533
rect 240592 233481 240598 233533
rect 240650 233521 240656 233533
rect 290416 233521 290422 233533
rect 240650 233493 290422 233521
rect 240650 233481 240656 233493
rect 290416 233481 290422 233493
rect 290474 233481 290480 233533
rect 297232 233481 297238 233533
rect 297290 233521 297296 233533
rect 328336 233521 328342 233533
rect 297290 233493 328342 233521
rect 297290 233481 297296 233493
rect 328336 233481 328342 233493
rect 328394 233481 328400 233533
rect 338608 233481 338614 233533
rect 338666 233521 338672 233533
rect 466480 233521 466486 233533
rect 338666 233493 466486 233521
rect 338666 233481 338672 233493
rect 466480 233481 466486 233493
rect 466538 233481 466544 233533
rect 194608 233407 194614 233459
rect 194666 233447 194672 233459
rect 196048 233447 196054 233459
rect 194666 233419 196054 233447
rect 194666 233407 194672 233419
rect 196048 233407 196054 233419
rect 196106 233407 196112 233459
rect 196144 233407 196150 233459
rect 196202 233447 196208 233459
rect 199120 233447 199126 233459
rect 196202 233419 199126 233447
rect 196202 233407 196208 233419
rect 199120 233407 199126 233419
rect 199178 233407 199184 233459
rect 199696 233407 199702 233459
rect 199754 233447 199760 233459
rect 206608 233447 206614 233459
rect 199754 233419 206614 233447
rect 199754 233407 199760 233419
rect 206608 233407 206614 233419
rect 206666 233407 206672 233459
rect 264400 233407 264406 233459
rect 264458 233447 264464 233459
rect 272848 233447 272854 233459
rect 264458 233419 272854 233447
rect 264458 233407 264464 233419
rect 272848 233407 272854 233419
rect 272906 233407 272912 233459
rect 287440 233407 287446 233459
rect 287498 233447 287504 233459
rect 311152 233447 311158 233459
rect 287498 233419 311158 233447
rect 287498 233407 287504 233419
rect 311152 233407 311158 233419
rect 311210 233407 311216 233459
rect 320272 233407 320278 233459
rect 320330 233447 320336 233459
rect 448240 233447 448246 233459
rect 320330 233419 448246 233447
rect 320330 233407 320336 233419
rect 448240 233407 448246 233419
rect 448298 233407 448304 233459
rect 192400 233333 192406 233385
rect 192458 233373 192464 233385
rect 193744 233373 193750 233385
rect 192458 233345 193750 233373
rect 192458 233333 192464 233345
rect 193744 233333 193750 233345
rect 193802 233333 193808 233385
rect 193840 233333 193846 233385
rect 193898 233373 193904 233385
rect 196816 233373 196822 233385
rect 193898 233345 196822 233373
rect 193898 233333 193904 233345
rect 196816 233333 196822 233345
rect 196874 233333 196880 233385
rect 197968 233333 197974 233385
rect 198026 233373 198032 233385
rect 203632 233373 203638 233385
rect 198026 233345 203638 233373
rect 198026 233333 198032 233345
rect 203632 233333 203638 233345
rect 203690 233333 203696 233385
rect 203920 233333 203926 233385
rect 203978 233373 203984 233385
rect 214192 233373 214198 233385
rect 203978 233345 214198 233373
rect 203978 233333 203984 233345
rect 214192 233333 214198 233345
rect 214250 233333 214256 233385
rect 226672 233333 226678 233385
rect 226730 233373 226736 233385
rect 236752 233373 236758 233385
rect 226730 233345 236758 233373
rect 226730 233333 226736 233345
rect 236752 233333 236758 233345
rect 236810 233333 236816 233385
rect 261616 233333 261622 233385
rect 261674 233373 261680 233385
rect 269008 233373 269014 233385
rect 261674 233345 269014 233373
rect 261674 233333 261680 233345
rect 269008 233333 269014 233345
rect 269066 233333 269072 233385
rect 270448 233333 270454 233385
rect 270506 233373 270512 233385
rect 275056 233373 275062 233385
rect 270506 233345 275062 233373
rect 270506 233333 270512 233345
rect 275056 233333 275062 233345
rect 275114 233333 275120 233385
rect 288400 233333 288406 233385
rect 288458 233373 288464 233385
rect 311056 233373 311062 233385
rect 288458 233345 311062 233373
rect 288458 233333 288464 233345
rect 311056 233333 311062 233345
rect 311114 233333 311120 233385
rect 324784 233333 324790 233385
rect 324842 233373 324848 233385
rect 327760 233373 327766 233385
rect 324842 233345 327766 233373
rect 324842 233333 324848 233345
rect 327760 233333 327766 233345
rect 327818 233333 327824 233385
rect 328528 233333 328534 233385
rect 328586 233373 328592 233385
rect 331120 233373 331126 233385
rect 328586 233345 331126 233373
rect 328586 233333 328592 233345
rect 331120 233333 331126 233345
rect 331178 233333 331184 233385
rect 335344 233333 335350 233385
rect 335402 233373 335408 233385
rect 463600 233373 463606 233385
rect 335402 233345 463606 233373
rect 335402 233333 335408 233345
rect 463600 233333 463606 233345
rect 463658 233333 463664 233385
rect 193456 233259 193462 233311
rect 193514 233299 193520 233311
rect 194608 233299 194614 233311
rect 193514 233271 194614 233299
rect 193514 233259 193520 233271
rect 194608 233259 194614 233271
rect 194666 233259 194672 233311
rect 195184 233259 195190 233311
rect 195242 233299 195248 233311
rect 197488 233299 197494 233311
rect 195242 233271 197494 233299
rect 195242 233259 195248 233271
rect 197488 233259 197494 233271
rect 197546 233259 197552 233311
rect 197872 233259 197878 233311
rect 197930 233299 197936 233311
rect 202096 233299 202102 233311
rect 197930 233271 202102 233299
rect 197930 233259 197936 233271
rect 202096 233259 202102 233271
rect 202154 233259 202160 233311
rect 202384 233259 202390 233311
rect 202442 233299 202448 233311
rect 211120 233299 211126 233311
rect 202442 233271 211126 233299
rect 202442 233259 202448 233271
rect 211120 233259 211126 233271
rect 211178 233259 211184 233311
rect 257968 233259 257974 233311
rect 258026 233299 258032 233311
rect 269488 233299 269494 233311
rect 258026 233271 269494 233299
rect 258026 233259 258032 233271
rect 269488 233259 269494 233271
rect 269546 233259 269552 233311
rect 270256 233259 270262 233311
rect 270314 233299 270320 233311
rect 273520 233299 273526 233311
rect 270314 233271 273526 233299
rect 270314 233259 270320 233271
rect 273520 233259 273526 233271
rect 273578 233259 273584 233311
rect 297136 233259 297142 233311
rect 297194 233299 297200 233311
rect 319408 233299 319414 233311
rect 297194 233271 319414 233299
rect 297194 233259 297200 233271
rect 319408 233259 319414 233271
rect 319466 233259 319472 233311
rect 319888 233259 319894 233311
rect 319946 233299 319952 233311
rect 377296 233299 377302 233311
rect 319946 233271 377302 233299
rect 319946 233259 319952 233271
rect 377296 233259 377302 233271
rect 377354 233259 377360 233311
rect 386320 233259 386326 233311
rect 386378 233299 386384 233311
rect 388720 233299 388726 233311
rect 386378 233271 388726 233299
rect 386378 233259 386384 233271
rect 388720 233259 388726 233271
rect 388778 233259 388784 233311
rect 395920 233259 395926 233311
rect 395978 233299 395984 233311
rect 400240 233299 400246 233311
rect 395978 233271 400246 233299
rect 395978 233259 395984 233271
rect 400240 233259 400246 233271
rect 400298 233259 400304 233311
rect 401200 233259 401206 233311
rect 401258 233299 401264 233311
rect 408880 233299 408886 233311
rect 401258 233271 408886 233299
rect 401258 233259 401264 233271
rect 408880 233259 408886 233271
rect 408938 233259 408944 233311
rect 259120 233185 259126 233237
rect 259178 233225 259184 233237
rect 328144 233225 328150 233237
rect 259178 233197 328150 233225
rect 259178 233185 259184 233197
rect 328144 233185 328150 233197
rect 328202 233185 328208 233237
rect 340816 233185 340822 233237
rect 340874 233225 340880 233237
rect 491248 233225 491254 233237
rect 340874 233197 491254 233225
rect 340874 233185 340880 233197
rect 491248 233185 491254 233197
rect 491306 233185 491312 233237
rect 495376 233185 495382 233237
rect 495434 233225 495440 233237
rect 614992 233225 614998 233237
rect 495434 233197 614998 233225
rect 495434 233185 495440 233197
rect 614992 233185 614998 233197
rect 615050 233185 615056 233237
rect 262096 233111 262102 233163
rect 262154 233151 262160 233163
rect 334192 233151 334198 233163
rect 262154 233123 334198 233151
rect 262154 233111 262160 233123
rect 334192 233111 334198 233123
rect 334250 233111 334256 233163
rect 347056 233111 347062 233163
rect 347114 233151 347120 233163
rect 501040 233151 501046 233163
rect 347114 233123 501046 233151
rect 347114 233111 347120 233123
rect 501040 233111 501046 233123
rect 501098 233111 501104 233163
rect 265744 233037 265750 233089
rect 265802 233077 265808 233089
rect 338032 233077 338038 233089
rect 265802 233049 338038 233077
rect 265802 233037 265808 233049
rect 338032 233037 338038 233049
rect 338090 233037 338096 233089
rect 350320 233037 350326 233089
rect 350378 233077 350384 233089
rect 507088 233077 507094 233089
rect 350378 233049 507094 233077
rect 350378 233037 350384 233049
rect 507088 233037 507094 233049
rect 507146 233037 507152 233089
rect 260656 232963 260662 233015
rect 260714 233003 260720 233015
rect 331312 233003 331318 233015
rect 260714 232975 331318 233003
rect 260714 232963 260720 232975
rect 331312 232963 331318 232975
rect 331370 232963 331376 233015
rect 353104 232963 353110 233015
rect 353162 233003 353168 233015
rect 513136 233003 513142 233015
rect 353162 232975 513142 233003
rect 353162 232963 353168 232975
rect 513136 232963 513142 232975
rect 513194 232963 513200 233015
rect 289936 232889 289942 232941
rect 289994 232929 290000 232941
rect 382864 232929 382870 232941
rect 289994 232901 382870 232929
rect 289994 232889 290000 232901
rect 382864 232889 382870 232901
rect 382922 232889 382928 232941
rect 410032 232889 410038 232941
rect 410090 232929 410096 232941
rect 572080 232929 572086 232941
rect 410090 232901 572086 232929
rect 410090 232889 410096 232901
rect 572080 232889 572086 232901
rect 572138 232889 572144 232941
rect 263920 232815 263926 232867
rect 263978 232855 263984 232867
rect 337264 232855 337270 232867
rect 263978 232827 337270 232855
rect 263978 232815 263984 232827
rect 337264 232815 337270 232827
rect 337322 232815 337328 232867
rect 356272 232815 356278 232867
rect 356330 232855 356336 232867
rect 519184 232855 519190 232867
rect 356330 232827 519190 232855
rect 356330 232815 356336 232827
rect 519184 232815 519190 232827
rect 519242 232815 519248 232867
rect 216592 232741 216598 232793
rect 216650 232781 216656 232793
rect 242128 232781 242134 232793
rect 216650 232753 242134 232781
rect 216650 232741 216656 232753
rect 242128 232741 242134 232753
rect 242186 232741 242192 232793
rect 265168 232741 265174 232793
rect 265226 232781 265232 232793
rect 340240 232781 340246 232793
rect 265226 232753 340246 232781
rect 265226 232741 265232 232753
rect 340240 232741 340246 232753
rect 340298 232741 340304 232793
rect 359056 232741 359062 232793
rect 359114 232781 359120 232793
rect 525232 232781 525238 232793
rect 359114 232753 525238 232781
rect 359114 232741 359120 232753
rect 525232 232741 525238 232753
rect 525290 232741 525296 232793
rect 237616 232667 237622 232719
rect 237674 232707 237680 232719
rect 284368 232707 284374 232719
rect 237674 232679 284374 232707
rect 237674 232667 237680 232679
rect 284368 232667 284374 232679
rect 284426 232667 284432 232719
rect 295312 232667 295318 232719
rect 295370 232707 295376 232719
rect 397360 232707 397366 232719
rect 295370 232679 397366 232707
rect 295370 232667 295376 232679
rect 397360 232667 397366 232679
rect 397418 232667 397424 232719
rect 399184 232667 399190 232719
rect 399242 232707 399248 232719
rect 566704 232707 566710 232719
rect 399242 232679 566710 232707
rect 399242 232667 399248 232679
rect 566704 232667 566710 232679
rect 566762 232667 566768 232719
rect 218032 232593 218038 232645
rect 218090 232633 218096 232645
rect 245104 232633 245110 232645
rect 218090 232605 245110 232633
rect 218090 232593 218096 232605
rect 245104 232593 245110 232605
rect 245162 232593 245168 232645
rect 268432 232593 268438 232645
rect 268490 232633 268496 232645
rect 346288 232633 346294 232645
rect 268490 232605 346294 232633
rect 268490 232593 268496 232605
rect 346288 232593 346294 232605
rect 346346 232593 346352 232645
rect 352336 232633 352342 232645
rect 346690 232605 352342 232633
rect 219760 232519 219766 232571
rect 219818 232559 219824 232571
rect 248080 232559 248086 232571
rect 219818 232531 248086 232559
rect 219818 232519 219824 232531
rect 248080 232519 248086 232531
rect 248138 232519 248144 232571
rect 266608 232519 266614 232571
rect 266666 232559 266672 232571
rect 343216 232559 343222 232571
rect 266666 232531 343222 232559
rect 266666 232519 266672 232531
rect 343216 232519 343222 232531
rect 343274 232519 343280 232571
rect 221104 232445 221110 232497
rect 221162 232485 221168 232497
rect 251152 232485 251158 232497
rect 221162 232457 251158 232485
rect 221162 232445 221168 232457
rect 251152 232445 251158 232457
rect 251210 232445 251216 232497
rect 271216 232445 271222 232497
rect 271274 232485 271280 232497
rect 346690 232485 346718 232605
rect 352336 232593 352342 232605
rect 352394 232593 352400 232645
rect 362128 232593 362134 232645
rect 362186 232633 362192 232645
rect 531280 232633 531286 232645
rect 362186 232605 531286 232633
rect 362186 232593 362192 232605
rect 531280 232593 531286 232605
rect 531338 232593 531344 232645
rect 356080 232559 356086 232571
rect 271274 232457 346718 232485
rect 346786 232531 356086 232559
rect 271274 232445 271280 232457
rect 222544 232371 222550 232423
rect 222602 232411 222608 232423
rect 254224 232411 254230 232423
rect 222602 232383 254230 232411
rect 222602 232371 222608 232383
rect 254224 232371 254230 232383
rect 254282 232371 254288 232423
rect 274864 232371 274870 232423
rect 274922 232411 274928 232423
rect 346786 232411 346814 232531
rect 356080 232519 356086 232531
rect 356138 232519 356144 232571
rect 365392 232519 365398 232571
rect 365450 232559 365456 232571
rect 537232 232559 537238 232571
rect 365450 232531 537238 232559
rect 365450 232519 365456 232531
rect 537232 232519 537238 232531
rect 537290 232519 537296 232571
rect 366256 232445 366262 232497
rect 366314 232485 366320 232497
rect 542608 232485 542614 232497
rect 366314 232457 542614 232485
rect 366314 232445 366320 232457
rect 542608 232445 542614 232457
rect 542666 232445 542672 232497
rect 349360 232411 349366 232423
rect 274922 232383 346814 232411
rect 346882 232383 349366 232411
rect 274922 232371 274928 232383
rect 222928 232297 222934 232349
rect 222986 232337 222992 232349
rect 255664 232337 255670 232349
rect 222986 232309 255670 232337
rect 222986 232297 222992 232309
rect 255664 232297 255670 232309
rect 255722 232297 255728 232349
rect 269680 232297 269686 232349
rect 269738 232337 269744 232349
rect 346882 232337 346910 232383
rect 349360 232371 349366 232383
rect 349418 232371 349424 232423
rect 365008 232371 365014 232423
rect 365066 232411 365072 232423
rect 539536 232411 539542 232423
rect 365066 232383 539542 232411
rect 365066 232371 365072 232383
rect 539536 232371 539542 232383
rect 539594 232371 539600 232423
rect 269738 232309 346910 232337
rect 269738 232297 269744 232309
rect 346960 232297 346966 232349
rect 347018 232337 347024 232349
rect 361360 232337 361366 232349
rect 347018 232309 361366 232337
rect 347018 232297 347024 232309
rect 361360 232297 361366 232309
rect 361418 232297 361424 232349
rect 368176 232297 368182 232349
rect 368234 232337 368240 232349
rect 543376 232337 543382 232349
rect 368234 232309 543382 232337
rect 368234 232297 368240 232309
rect 543376 232297 543382 232309
rect 543434 232297 543440 232349
rect 224272 232223 224278 232275
rect 224330 232263 224336 232275
rect 257200 232263 257206 232275
rect 224330 232235 257206 232263
rect 224330 232223 224336 232235
rect 257200 232223 257206 232235
rect 257258 232223 257264 232275
rect 274192 232223 274198 232275
rect 274250 232263 274256 232275
rect 358288 232263 358294 232275
rect 274250 232235 358294 232263
rect 274250 232223 274256 232235
rect 358288 232223 358294 232235
rect 358346 232223 358352 232275
rect 369520 232223 369526 232275
rect 369578 232263 369584 232275
rect 548560 232263 548566 232275
rect 369578 232235 548566 232263
rect 369578 232223 369584 232235
rect 548560 232223 548566 232235
rect 548618 232223 548624 232275
rect 226288 232149 226294 232201
rect 226346 232189 226352 232201
rect 261712 232189 261718 232201
rect 226346 232161 261718 232189
rect 226346 232149 226352 232161
rect 261712 232149 261718 232161
rect 261770 232149 261776 232201
rect 272944 232149 272950 232201
rect 273002 232189 273008 232201
rect 355312 232189 355318 232201
rect 273002 232161 355318 232189
rect 273002 232149 273008 232161
rect 355312 232149 355318 232161
rect 355370 232149 355376 232201
rect 368080 232149 368086 232201
rect 368138 232189 368144 232201
rect 545584 232189 545590 232201
rect 368138 232161 545590 232189
rect 368138 232149 368144 232161
rect 545584 232149 545590 232161
rect 545642 232149 545648 232201
rect 227056 232075 227062 232127
rect 227114 232115 227120 232127
rect 263248 232115 263254 232127
rect 227114 232087 263254 232115
rect 227114 232075 227120 232087
rect 263248 232075 263254 232087
rect 263306 232075 263312 232127
rect 277456 232075 277462 232127
rect 277514 232115 277520 232127
rect 364432 232115 364438 232127
rect 277514 232087 364438 232115
rect 277514 232075 277520 232087
rect 364432 232075 364438 232087
rect 364490 232075 364496 232127
rect 372688 232075 372694 232127
rect 372746 232115 372752 232127
rect 552400 232115 552406 232127
rect 372746 232087 552406 232115
rect 372746 232075 372752 232087
rect 552400 232075 552406 232087
rect 552458 232075 552464 232127
rect 233872 232001 233878 232053
rect 233930 232041 233936 232053
rect 274480 232041 274486 232053
rect 233930 232013 274486 232041
rect 233930 232001 233936 232013
rect 274480 232001 274486 232013
rect 274538 232001 274544 232053
rect 275728 232001 275734 232053
rect 275786 232041 275792 232053
rect 346960 232041 346966 232053
rect 275786 232013 346966 232041
rect 275786 232001 275792 232013
rect 346960 232001 346966 232013
rect 347018 232001 347024 232053
rect 354256 232001 354262 232053
rect 354314 232041 354320 232053
rect 367120 232041 367126 232053
rect 354314 232013 367126 232041
rect 354314 232001 354320 232013
rect 367120 232001 367126 232013
rect 367178 232001 367184 232053
rect 372304 232001 372310 232053
rect 372362 232041 372368 232053
rect 554704 232041 554710 232053
rect 372362 232013 554710 232041
rect 372362 232001 372368 232013
rect 554704 232001 554710 232013
rect 554762 232001 554768 232053
rect 234832 231927 234838 231979
rect 234890 231967 234896 231979
rect 278320 231967 278326 231979
rect 234890 231939 278326 231967
rect 234890 231927 234896 231939
rect 278320 231927 278326 231939
rect 278378 231927 278384 231979
rect 278992 231927 278998 231979
rect 279050 231967 279056 231979
rect 367408 231967 367414 231979
rect 279050 231939 367414 231967
rect 279050 231927 279056 231939
rect 367408 231927 367414 231939
rect 367466 231927 367472 231979
rect 375760 231927 375766 231979
rect 375818 231967 375824 231979
rect 558448 231967 558454 231979
rect 375818 231939 558454 231967
rect 375818 231927 375824 231939
rect 558448 231927 558454 231939
rect 558506 231927 558512 231979
rect 233200 231853 233206 231905
rect 233258 231893 233264 231905
rect 275344 231893 275350 231905
rect 233258 231865 275350 231893
rect 233258 231853 233264 231865
rect 275344 231853 275350 231865
rect 275402 231853 275408 231905
rect 280240 231853 280246 231905
rect 280298 231893 280304 231905
rect 370384 231893 370390 231905
rect 280298 231865 370390 231893
rect 280298 231853 280304 231865
rect 370384 231853 370390 231865
rect 370442 231853 370448 231905
rect 374512 231853 374518 231905
rect 374570 231893 374576 231905
rect 557008 231893 557014 231905
rect 374570 231865 557014 231893
rect 374570 231853 374576 231865
rect 557008 231853 557014 231865
rect 557066 231853 557072 231905
rect 235984 231779 235990 231831
rect 236042 231819 236048 231831
rect 281296 231819 281302 231831
rect 236042 231791 281302 231819
rect 236042 231779 236048 231791
rect 281296 231779 281302 231791
rect 281354 231779 281360 231831
rect 281968 231779 281974 231831
rect 282026 231819 282032 231831
rect 373456 231819 373462 231831
rect 282026 231791 373462 231819
rect 282026 231779 282032 231791
rect 373456 231779 373462 231791
rect 373514 231779 373520 231831
rect 378928 231779 378934 231831
rect 378986 231819 378992 231831
rect 564496 231819 564502 231831
rect 378986 231791 564502 231819
rect 378986 231779 378992 231791
rect 564496 231779 564502 231791
rect 564554 231779 564560 231831
rect 258736 231705 258742 231757
rect 258794 231745 258800 231757
rect 326704 231745 326710 231757
rect 258794 231717 326710 231745
rect 258794 231705 258800 231717
rect 326704 231705 326710 231717
rect 326762 231705 326768 231757
rect 337552 231705 337558 231757
rect 337610 231745 337616 231757
rect 485200 231745 485206 231757
rect 337610 231717 485206 231745
rect 337610 231705 337616 231717
rect 485200 231705 485206 231717
rect 485258 231705 485264 231757
rect 255760 231631 255766 231683
rect 255818 231671 255824 231683
rect 320560 231671 320566 231683
rect 255818 231643 320566 231671
rect 255818 231631 255824 231643
rect 320560 231631 320566 231643
rect 320618 231631 320624 231683
rect 334864 231631 334870 231683
rect 334922 231671 334928 231683
rect 479152 231671 479158 231683
rect 334922 231643 479158 231671
rect 334922 231631 334928 231643
rect 479152 231631 479158 231643
rect 479210 231631 479216 231683
rect 257584 231557 257590 231609
rect 257642 231597 257648 231609
rect 325168 231597 325174 231609
rect 257642 231569 325174 231597
rect 257642 231557 257648 231569
rect 325168 231557 325174 231569
rect 325226 231557 325232 231609
rect 327088 231557 327094 231609
rect 327146 231597 327152 231609
rect 464080 231597 464086 231609
rect 327146 231569 464086 231597
rect 327146 231557 327152 231569
rect 464080 231557 464086 231569
rect 464138 231557 464144 231609
rect 248368 231483 248374 231535
rect 248426 231523 248432 231535
rect 305488 231523 305494 231535
rect 248426 231495 305494 231523
rect 248426 231483 248432 231495
rect 305488 231483 305494 231495
rect 305546 231483 305552 231535
rect 312208 231483 312214 231535
rect 312266 231523 312272 231535
rect 433840 231523 433846 231535
rect 312266 231495 433846 231523
rect 312266 231483 312272 231495
rect 433840 231483 433846 231495
rect 433898 231483 433904 231535
rect 281200 231409 281206 231461
rect 281258 231449 281264 231461
rect 289648 231449 289654 231461
rect 281258 231421 289654 231449
rect 281258 231409 281264 231421
rect 289648 231409 289654 231421
rect 289706 231409 289712 231461
rect 290800 231409 290806 231461
rect 290858 231449 290864 231461
rect 374608 231449 374614 231461
rect 290858 231421 374614 231449
rect 290858 231409 290864 231421
rect 374608 231409 374614 231421
rect 374666 231409 374672 231461
rect 403120 231409 403126 231461
rect 403178 231449 403184 231461
rect 520720 231449 520726 231461
rect 403178 231421 520726 231449
rect 403178 231409 403184 231421
rect 520720 231409 520726 231421
rect 520778 231409 520784 231461
rect 292528 231335 292534 231387
rect 292586 231375 292592 231387
rect 379984 231375 379990 231387
rect 292586 231347 379990 231375
rect 292586 231335 292592 231347
rect 379984 231335 379990 231347
rect 380042 231335 380048 231387
rect 400144 231335 400150 231387
rect 400202 231375 400208 231387
rect 499600 231375 499606 231387
rect 400202 231347 499606 231375
rect 400202 231335 400208 231347
rect 499600 231335 499606 231347
rect 499658 231335 499664 231387
rect 245200 231261 245206 231313
rect 245258 231301 245264 231313
rect 299440 231301 299446 231313
rect 245258 231273 299446 231301
rect 245258 231261 245264 231273
rect 299440 231261 299446 231273
rect 299498 231261 299504 231313
rect 300208 231261 300214 231313
rect 300266 231301 300272 231313
rect 385840 231301 385846 231313
rect 300266 231273 385846 231301
rect 300266 231261 300272 231273
rect 385840 231261 385846 231273
rect 385898 231261 385904 231313
rect 395056 231261 395062 231313
rect 395114 231301 395120 231313
rect 485968 231301 485974 231313
rect 395114 231273 485974 231301
rect 395114 231261 395120 231273
rect 485968 231261 485974 231273
rect 486026 231261 486032 231313
rect 293488 231187 293494 231239
rect 293546 231227 293552 231239
rect 365104 231227 365110 231239
rect 293546 231199 365110 231227
rect 293546 231187 293552 231199
rect 365104 231187 365110 231199
rect 365162 231187 365168 231239
rect 394768 231187 394774 231239
rect 394826 231227 394832 231239
rect 473872 231227 473878 231239
rect 394826 231199 473878 231227
rect 394826 231187 394832 231199
rect 473872 231187 473878 231199
rect 473930 231187 473936 231239
rect 256144 231113 256150 231165
rect 256202 231153 256208 231165
rect 322096 231153 322102 231165
rect 256202 231125 322102 231153
rect 256202 231113 256208 231125
rect 322096 231113 322102 231125
rect 322154 231113 322160 231165
rect 337360 231113 337366 231165
rect 337418 231153 337424 231165
rect 337418 231125 414686 231153
rect 337418 231113 337424 231125
rect 252976 231039 252982 231091
rect 253034 231079 253040 231091
rect 314512 231079 314518 231091
rect 253034 231051 314518 231079
rect 253034 231039 253040 231051
rect 314512 231039 314518 231051
rect 314570 231039 314576 231091
rect 344464 231039 344470 231091
rect 344522 231079 344528 231091
rect 344522 231051 407534 231079
rect 344522 231039 344528 231051
rect 290608 230965 290614 231017
rect 290666 231005 290672 231017
rect 297424 231005 297430 231017
rect 290666 230977 297430 231005
rect 290666 230965 290672 230977
rect 297424 230965 297430 230977
rect 297482 230965 297488 231017
rect 308176 230965 308182 231017
rect 308234 231005 308240 231017
rect 323632 231005 323638 231017
rect 308234 230977 323638 231005
rect 308234 230965 308240 230977
rect 323632 230965 323638 230977
rect 323690 230965 323696 231017
rect 328336 230965 328342 231017
rect 328394 231005 328400 231017
rect 401392 231005 401398 231017
rect 328394 230977 401398 231005
rect 328394 230965 328400 230977
rect 401392 230965 401398 230977
rect 401450 230965 401456 231017
rect 323056 230891 323062 230943
rect 323114 230931 323120 230943
rect 329584 230931 329590 230943
rect 323114 230903 329590 230931
rect 323114 230891 323120 230903
rect 329584 230891 329590 230903
rect 329642 230891 329648 230943
rect 331216 230891 331222 230943
rect 331274 230931 331280 230943
rect 395344 230931 395350 230943
rect 331274 230903 395350 230931
rect 331274 230891 331280 230903
rect 395344 230891 395350 230903
rect 395402 230891 395408 230943
rect 407506 230931 407534 231051
rect 414658 231005 414686 231125
rect 414736 231113 414742 231165
rect 414794 231153 414800 231165
rect 424048 231153 424054 231165
rect 414794 231125 424054 231153
rect 414794 231113 414800 231125
rect 424048 231113 424054 231125
rect 424106 231113 424112 231165
rect 415696 231005 415702 231017
rect 414658 230977 415702 231005
rect 415696 230965 415702 230977
rect 415754 230965 415760 231017
rect 419536 230931 419542 230943
rect 407506 230903 419542 230931
rect 419536 230891 419542 230903
rect 419594 230891 419600 230943
rect 282544 230817 282550 230869
rect 282602 230857 282608 230869
rect 300592 230857 300598 230869
rect 282602 230829 300598 230857
rect 282602 230817 282608 230829
rect 300592 230817 300598 230829
rect 300650 230817 300656 230869
rect 326800 230817 326806 230869
rect 326858 230857 326864 230869
rect 380176 230857 380182 230869
rect 326858 230829 380182 230857
rect 326858 230817 326864 230829
rect 380176 230817 380182 230829
rect 380234 230817 380240 230869
rect 387280 230817 387286 230869
rect 387338 230857 387344 230869
rect 449680 230857 449686 230869
rect 387338 230829 449686 230857
rect 387338 230817 387344 230829
rect 449680 230817 449686 230829
rect 449738 230817 449744 230869
rect 319600 230743 319606 230795
rect 319658 230783 319664 230795
rect 365008 230783 365014 230795
rect 319658 230755 365014 230783
rect 319658 230743 319664 230755
rect 365008 230743 365014 230755
rect 365066 230743 365072 230795
rect 367120 230743 367126 230795
rect 367178 230783 367184 230795
rect 409648 230783 409654 230795
rect 367178 230755 409654 230783
rect 367178 230743 367184 230755
rect 409648 230743 409654 230755
rect 409706 230743 409712 230795
rect 313936 230669 313942 230721
rect 313994 230709 314000 230721
rect 362128 230709 362134 230721
rect 313994 230681 362134 230709
rect 313994 230669 314000 230681
rect 362128 230669 362134 230681
rect 362186 230669 362192 230721
rect 362608 230669 362614 230721
rect 362666 230709 362672 230721
rect 416464 230709 416470 230721
rect 362666 230681 416470 230709
rect 362666 230669 362672 230681
rect 416464 230669 416470 230681
rect 416522 230669 416528 230721
rect 302320 230595 302326 230647
rect 302378 230635 302384 230647
rect 308560 230635 308566 230647
rect 302378 230607 308566 230635
rect 302378 230595 302384 230607
rect 308560 230595 308566 230607
rect 308618 230595 308624 230647
rect 320656 230595 320662 230647
rect 320714 230635 320720 230647
rect 374224 230635 374230 230647
rect 320714 230607 374230 230635
rect 320714 230595 320720 230607
rect 374224 230595 374230 230607
rect 374282 230595 374288 230647
rect 306640 230521 306646 230573
rect 306698 230561 306704 230573
rect 317584 230561 317590 230573
rect 306698 230533 317590 230561
rect 306698 230521 306704 230533
rect 317584 230521 317590 230533
rect 317642 230521 317648 230573
rect 323152 230521 323158 230573
rect 323210 230561 323216 230573
rect 377104 230561 377110 230573
rect 323210 230533 377110 230561
rect 323210 230521 323216 230533
rect 377104 230521 377110 230533
rect 377162 230521 377168 230573
rect 147472 230447 147478 230499
rect 147530 230487 147536 230499
rect 154096 230487 154102 230499
rect 147530 230459 154102 230487
rect 147530 230447 147536 230459
rect 154096 230447 154102 230459
rect 154154 230447 154160 230499
rect 299248 230447 299254 230499
rect 299306 230487 299312 230499
rect 302512 230487 302518 230499
rect 299306 230459 302518 230487
rect 299306 230447 299312 230459
rect 302512 230447 302518 230459
rect 302570 230447 302576 230499
rect 304144 230447 304150 230499
rect 304202 230487 304208 230499
rect 311632 230487 311638 230499
rect 304202 230459 311638 230487
rect 304202 230447 304208 230459
rect 311632 230447 311638 230459
rect 311690 230447 311696 230499
rect 320848 230447 320854 230499
rect 320906 230487 320912 230499
rect 368176 230487 368182 230499
rect 320906 230459 368182 230487
rect 320906 230447 320912 230459
rect 368176 230447 368182 230459
rect 368234 230447 368240 230499
rect 426160 230447 426166 230499
rect 426218 230487 426224 230499
rect 436144 230487 436150 230499
rect 426218 230459 436150 230487
rect 426218 230447 426224 230459
rect 436144 230447 436150 230459
rect 436202 230447 436208 230499
rect 246160 230373 246166 230425
rect 246218 230413 246224 230425
rect 298672 230413 298678 230425
rect 246218 230385 298678 230413
rect 246218 230373 246224 230385
rect 298672 230373 298678 230385
rect 298730 230373 298736 230425
rect 313456 230373 313462 230425
rect 313514 230413 313520 230425
rect 436912 230413 436918 230425
rect 313514 230385 436918 230413
rect 313514 230373 313520 230385
rect 436912 230373 436918 230385
rect 436970 230373 436976 230425
rect 241072 230299 241078 230351
rect 241130 230339 241136 230351
rect 291952 230339 291958 230351
rect 241130 230311 291958 230339
rect 241130 230299 241136 230311
rect 291952 230299 291958 230311
rect 292010 230299 292016 230351
rect 314896 230299 314902 230351
rect 314954 230339 314960 230351
rect 439984 230339 439990 230351
rect 314954 230311 439990 230339
rect 314954 230299 314960 230311
rect 439984 230299 439990 230311
rect 440042 230299 440048 230351
rect 245776 230225 245782 230277
rect 245834 230265 245840 230277
rect 300976 230265 300982 230277
rect 245834 230237 300982 230265
rect 245834 230225 245840 230237
rect 300976 230225 300982 230237
rect 301034 230225 301040 230277
rect 317968 230225 317974 230277
rect 318026 230265 318032 230277
rect 445936 230265 445942 230277
rect 318026 230237 445942 230265
rect 318026 230225 318032 230237
rect 445936 230225 445942 230237
rect 445994 230225 446000 230277
rect 451984 230265 451990 230277
rect 449218 230237 451990 230265
rect 248944 230151 248950 230203
rect 249002 230191 249008 230203
rect 304816 230191 304822 230203
rect 249002 230163 304822 230191
rect 249002 230151 249008 230163
rect 304816 230151 304822 230163
rect 304874 230151 304880 230203
rect 321232 230151 321238 230203
rect 321290 230191 321296 230203
rect 449218 230191 449246 230237
rect 451984 230225 451990 230237
rect 452042 230225 452048 230277
rect 321290 230163 449246 230191
rect 321290 230151 321296 230163
rect 449296 230151 449302 230203
rect 449354 230191 449360 230203
rect 466384 230191 466390 230203
rect 449354 230163 466390 230191
rect 449354 230151 449360 230163
rect 466384 230151 466390 230163
rect 466442 230151 466448 230203
rect 251920 230077 251926 230129
rect 251978 230117 251984 230129
rect 310768 230117 310774 230129
rect 251978 230089 310774 230117
rect 251978 230077 251984 230089
rect 310768 230077 310774 230089
rect 310826 230077 310832 230129
rect 325744 230077 325750 230129
rect 325802 230117 325808 230129
rect 461008 230117 461014 230129
rect 325802 230089 461014 230117
rect 325802 230077 325808 230089
rect 461008 230077 461014 230089
rect 461066 230077 461072 230129
rect 463600 230077 463606 230129
rect 463658 230117 463664 230129
rect 478384 230117 478390 230129
rect 463658 230089 478390 230117
rect 463658 230077 463664 230089
rect 478384 230077 478390 230089
rect 478442 230077 478448 230129
rect 248752 230003 248758 230055
rect 248810 230043 248816 230055
rect 307024 230043 307030 230055
rect 248810 230015 307030 230043
rect 248810 230003 248816 230015
rect 307024 230003 307030 230015
rect 307082 230003 307088 230055
rect 324016 230003 324022 230055
rect 324074 230043 324080 230055
rect 458032 230043 458038 230055
rect 324074 230015 458038 230043
rect 324074 230003 324080 230015
rect 458032 230003 458038 230015
rect 458090 230003 458096 230055
rect 466480 230003 466486 230055
rect 466538 230043 466544 230055
rect 484432 230043 484438 230055
rect 466538 230015 484438 230043
rect 466538 230003 466544 230015
rect 484432 230003 484438 230015
rect 484490 230003 484496 230055
rect 503920 230003 503926 230055
rect 503978 230043 503984 230055
rect 622672 230043 622678 230055
rect 503978 230015 622678 230043
rect 503978 230003 503984 230015
rect 622672 230003 622678 230015
rect 622730 230003 622736 230055
rect 227440 229929 227446 229981
rect 227498 229969 227504 229981
rect 264784 229969 264790 229981
rect 227498 229941 264790 229969
rect 227498 229929 227504 229941
rect 264784 229929 264790 229941
rect 264842 229929 264848 229981
rect 290896 229929 290902 229981
rect 290954 229969 290960 229981
rect 331888 229969 331894 229981
rect 290954 229941 331894 229969
rect 290954 229929 290960 229941
rect 331888 229929 331894 229941
rect 331946 229929 331952 229981
rect 434896 229929 434902 229981
rect 434954 229969 434960 229981
rect 454288 229969 454294 229981
rect 434954 229941 454294 229969
rect 434954 229929 434960 229941
rect 454288 229929 454294 229941
rect 454346 229929 454352 229981
rect 475216 229929 475222 229981
rect 475274 229969 475280 229981
rect 601456 229969 601462 229981
rect 475274 229941 601462 229969
rect 475274 229929 475280 229941
rect 601456 229929 601462 229941
rect 601514 229929 601520 229981
rect 250192 229855 250198 229907
rect 250250 229895 250256 229907
rect 310000 229895 310006 229907
rect 250250 229867 310006 229895
rect 250250 229855 250256 229867
rect 310000 229855 310006 229867
rect 310058 229855 310064 229907
rect 331600 229855 331606 229907
rect 331658 229895 331664 229907
rect 473104 229895 473110 229907
rect 331658 229867 473110 229895
rect 331658 229855 331664 229867
rect 473104 229855 473110 229867
rect 473162 229855 473168 229907
rect 480880 229855 480886 229907
rect 480938 229895 480944 229907
rect 609040 229895 609046 229907
rect 480938 229867 609046 229895
rect 480938 229855 480944 229867
rect 609040 229855 609046 229867
rect 609098 229855 609104 229907
rect 147088 229781 147094 229833
rect 147146 229821 147152 229833
rect 151408 229821 151414 229833
rect 147146 229793 151414 229821
rect 147146 229781 147152 229793
rect 151408 229781 151414 229793
rect 151466 229781 151472 229833
rect 251536 229781 251542 229833
rect 251594 229821 251600 229833
rect 313072 229821 313078 229833
rect 251594 229793 313078 229821
rect 251594 229781 251600 229793
rect 313072 229781 313078 229793
rect 313130 229781 313136 229833
rect 336304 229781 336310 229833
rect 336362 229821 336368 229833
rect 482128 229821 482134 229833
rect 336362 229793 482134 229821
rect 336362 229781 336368 229793
rect 482128 229781 482134 229793
rect 482186 229781 482192 229833
rect 484624 229781 484630 229833
rect 484682 229821 484688 229833
rect 612112 229821 612118 229833
rect 484682 229793 612118 229821
rect 484682 229781 484688 229793
rect 612112 229781 612118 229793
rect 612170 229781 612176 229833
rect 254800 229707 254806 229759
rect 254858 229747 254864 229759
rect 319120 229747 319126 229759
rect 254858 229719 319126 229747
rect 254858 229707 254864 229719
rect 319120 229707 319126 229719
rect 319178 229707 319184 229759
rect 348496 229707 348502 229759
rect 348554 229747 348560 229759
rect 504016 229747 504022 229759
rect 348554 229719 504022 229747
rect 348554 229707 348560 229719
rect 504016 229707 504022 229719
rect 504074 229707 504080 229759
rect 215248 229633 215254 229685
rect 215306 229673 215312 229685
rect 239056 229673 239062 229685
rect 215306 229645 239062 229673
rect 215306 229633 215312 229645
rect 239056 229633 239062 229645
rect 239114 229633 239120 229685
rect 244240 229633 244246 229685
rect 244298 229673 244304 229685
rect 298000 229673 298006 229685
rect 244298 229645 298006 229673
rect 244298 229633 244304 229645
rect 298000 229633 298006 229645
rect 298058 229633 298064 229685
rect 298384 229633 298390 229685
rect 298442 229673 298448 229685
rect 406768 229673 406774 229685
rect 298442 229645 406774 229673
rect 298442 229633 298448 229645
rect 406768 229633 406774 229645
rect 406826 229633 406832 229685
rect 409840 229633 409846 229685
rect 409898 229673 409904 229685
rect 565936 229673 565942 229685
rect 409898 229645 565942 229673
rect 409898 229633 409904 229645
rect 565936 229633 565942 229645
rect 565994 229633 566000 229685
rect 220144 229559 220150 229611
rect 220202 229599 220208 229611
rect 249712 229599 249718 229611
rect 220202 229571 249718 229599
rect 220202 229559 220208 229571
rect 249712 229559 249718 229571
rect 249770 229559 249776 229611
rect 253072 229559 253078 229611
rect 253130 229599 253136 229611
rect 316144 229599 316150 229611
rect 253130 229571 316150 229599
rect 253130 229559 253136 229571
rect 316144 229559 316150 229571
rect 316202 229559 316208 229611
rect 351760 229559 351766 229611
rect 351818 229599 351824 229611
rect 510160 229599 510166 229611
rect 351818 229571 510166 229599
rect 351818 229559 351824 229571
rect 510160 229559 510166 229571
rect 510218 229559 510224 229611
rect 221584 229485 221590 229537
rect 221642 229525 221648 229537
rect 252592 229525 252598 229537
rect 221642 229497 252598 229525
rect 221642 229485 221648 229497
rect 252592 229485 252598 229497
rect 252650 229485 252656 229537
rect 255184 229485 255190 229537
rect 255242 229525 255248 229537
rect 316816 229525 316822 229537
rect 255242 229497 316822 229525
rect 255242 229485 255248 229497
rect 316816 229485 316822 229497
rect 316874 229485 316880 229537
rect 354832 229485 354838 229537
rect 354890 229525 354896 229537
rect 516112 229525 516118 229537
rect 354890 229497 516118 229525
rect 354890 229485 354896 229497
rect 516112 229485 516118 229497
rect 516170 229485 516176 229537
rect 264304 229411 264310 229463
rect 264362 229451 264368 229463
rect 334960 229451 334966 229463
rect 264362 229423 334966 229451
rect 264362 229411 264368 229423
rect 334960 229411 334966 229423
rect 335018 229411 335024 229463
rect 357616 229411 357622 229463
rect 357674 229451 357680 229463
rect 357674 229423 377294 229451
rect 357674 229411 357680 229423
rect 230320 229337 230326 229389
rect 230378 229377 230384 229389
rect 269296 229377 269302 229389
rect 230378 229349 269302 229377
rect 230378 229337 230384 229349
rect 269296 229337 269302 229349
rect 269354 229337 269360 229389
rect 273520 229337 273526 229389
rect 273578 229377 273584 229389
rect 347056 229377 347062 229389
rect 273578 229349 347062 229377
rect 273578 229337 273584 229349
rect 347056 229337 347062 229349
rect 347114 229337 347120 229389
rect 369520 229377 369526 229389
rect 357106 229349 369526 229377
rect 231856 229263 231862 229315
rect 231914 229303 231920 229315
rect 272272 229303 272278 229315
rect 231914 229275 272278 229303
rect 231914 229263 231920 229275
rect 272272 229263 272278 229275
rect 272330 229263 272336 229315
rect 283504 229263 283510 229315
rect 283562 229303 283568 229315
rect 357106 229303 357134 229349
rect 369520 229337 369526 229349
rect 369578 229337 369584 229389
rect 369904 229337 369910 229389
rect 369962 229377 369968 229389
rect 377266 229377 377294 229423
rect 380080 229411 380086 229463
rect 380138 229451 380144 229463
rect 538864 229451 538870 229463
rect 380138 229423 538870 229451
rect 380138 229411 380144 229423
rect 538864 229411 538870 229423
rect 538922 229411 538928 229463
rect 522160 229377 522166 229389
rect 369962 229349 374654 229377
rect 377266 229349 522166 229377
rect 369962 229337 369968 229349
rect 283562 229275 357134 229303
rect 283562 229263 283568 229275
rect 357424 229263 357430 229315
rect 357482 229303 357488 229315
rect 374512 229303 374518 229315
rect 357482 229275 374518 229303
rect 357482 229263 357488 229275
rect 374512 229263 374518 229275
rect 374570 229263 374576 229315
rect 374626 229303 374654 229349
rect 522160 229337 522166 229349
rect 522218 229337 522224 229389
rect 546352 229303 546358 229315
rect 374626 229275 546358 229303
rect 546352 229263 546358 229275
rect 546410 229263 546416 229315
rect 233488 229189 233494 229241
rect 233546 229229 233552 229241
rect 276784 229229 276790 229241
rect 233546 229201 276790 229229
rect 233546 229189 233552 229201
rect 276784 229189 276790 229201
rect 276842 229189 276848 229241
rect 282160 229189 282166 229241
rect 282218 229229 282224 229241
rect 371248 229229 371254 229241
rect 282218 229201 371254 229229
rect 282218 229189 282224 229201
rect 371248 229189 371254 229201
rect 371306 229189 371312 229241
rect 374320 229189 374326 229241
rect 374378 229229 374384 229241
rect 555280 229229 555286 229241
rect 374378 229201 555286 229229
rect 374378 229189 374384 229201
rect 555280 229189 555286 229201
rect 555338 229189 555344 229241
rect 231952 229115 231958 229167
rect 232010 229155 232016 229167
rect 273808 229155 273814 229167
rect 232010 229127 273814 229155
rect 232010 229115 232016 229127
rect 273808 229115 273814 229127
rect 273866 229115 273872 229167
rect 287920 229115 287926 229167
rect 287978 229155 287984 229167
rect 374416 229155 374422 229167
rect 287978 229127 374422 229155
rect 287978 229115 287984 229127
rect 374416 229115 374422 229127
rect 374474 229115 374480 229167
rect 377200 229115 377206 229167
rect 377258 229155 377264 229167
rect 561424 229155 561430 229167
rect 377258 229127 561430 229155
rect 377258 229115 377264 229127
rect 561424 229115 561430 229127
rect 561482 229115 561488 229167
rect 238384 229041 238390 229093
rect 238442 229081 238448 229093
rect 283600 229081 283606 229093
rect 238442 229053 283606 229081
rect 238442 229041 238448 229053
rect 283600 229041 283606 229053
rect 283658 229041 283664 229093
rect 284752 229041 284758 229093
rect 284810 229081 284816 229093
rect 371536 229081 371542 229093
rect 284810 229053 371542 229081
rect 284810 229041 284816 229053
rect 371536 229041 371542 229053
rect 371594 229041 371600 229093
rect 376816 229041 376822 229093
rect 376874 229081 376880 229093
rect 563632 229081 563638 229093
rect 376874 229053 563638 229081
rect 376874 229041 376880 229053
rect 563632 229041 563638 229053
rect 563690 229041 563696 229093
rect 235216 228967 235222 229019
rect 235274 229007 235280 229019
rect 279856 229007 279862 229019
rect 235274 228979 279862 229007
rect 235274 228967 235280 228979
rect 279856 228967 279862 228979
rect 279914 228967 279920 229019
rect 286288 228967 286294 229019
rect 286346 229007 286352 229019
rect 357424 229007 357430 229019
rect 286346 228979 357430 229007
rect 286346 228967 286352 228979
rect 357424 228967 357430 228979
rect 357482 228967 357488 229019
rect 357520 228967 357526 229019
rect 357578 229007 357584 229019
rect 359920 229007 359926 229019
rect 357578 228979 359926 229007
rect 357578 228967 357584 228979
rect 359920 228967 359926 228979
rect 359978 228967 359984 229019
rect 368944 228967 368950 229019
rect 369002 229007 369008 229019
rect 370480 229007 370486 229019
rect 369002 228979 370486 229007
rect 369002 228967 369008 228979
rect 370480 228967 370486 228979
rect 370538 228967 370544 229019
rect 380464 228967 380470 229019
rect 380522 229007 380528 229019
rect 567472 229007 567478 229019
rect 380522 228979 567478 229007
rect 380522 228967 380528 228979
rect 567472 228967 567478 228979
rect 567530 228967 567536 229019
rect 242512 228893 242518 228945
rect 242570 228933 242576 228945
rect 294928 228933 294934 228945
rect 242570 228905 294934 228933
rect 242570 228893 242576 228905
rect 294928 228893 294934 228905
rect 294986 228893 294992 228945
rect 308944 228893 308950 228945
rect 309002 228933 309008 228945
rect 427792 228933 427798 228945
rect 309002 228905 427798 228933
rect 309002 228893 309008 228905
rect 427792 228893 427798 228905
rect 427850 228893 427856 228945
rect 427888 228893 427894 228945
rect 427946 228933 427952 228945
rect 547888 228933 547894 228945
rect 427946 228905 547894 228933
rect 427946 228893 427952 228905
rect 547888 228893 547894 228905
rect 547946 228893 547952 228945
rect 241648 228819 241654 228871
rect 241706 228859 241712 228871
rect 289744 228859 289750 228871
rect 241706 228831 289750 228859
rect 241706 228819 241712 228831
rect 289744 228819 289750 228831
rect 289802 228819 289808 228871
rect 310672 228819 310678 228871
rect 310730 228859 310736 228871
rect 430864 228859 430870 228871
rect 310730 228831 430870 228859
rect 310730 228819 310736 228831
rect 430864 228819 430870 228831
rect 430922 228819 430928 228871
rect 432016 228819 432022 228871
rect 432074 228859 432080 228871
rect 529744 228859 529750 228871
rect 432074 228831 529750 228859
rect 432074 228819 432080 228831
rect 529744 228819 529750 228831
rect 529802 228819 529808 228871
rect 239728 228745 239734 228797
rect 239786 228785 239792 228797
rect 288880 228785 288886 228797
rect 239786 228757 288886 228785
rect 239786 228745 239792 228757
rect 288880 228745 288886 228757
rect 288938 228745 288944 228797
rect 306160 228745 306166 228797
rect 306218 228785 306224 228797
rect 421840 228785 421846 228797
rect 306218 228757 421846 228785
rect 306218 228745 306224 228757
rect 421840 228745 421846 228757
rect 421898 228745 421904 228797
rect 228880 228671 228886 228723
rect 228938 228711 228944 228723
rect 267856 228711 267862 228723
rect 228938 228683 267862 228711
rect 228938 228671 228944 228683
rect 267856 228671 267862 228683
rect 267914 228671 267920 228723
rect 304432 228671 304438 228723
rect 304490 228711 304496 228723
rect 418768 228711 418774 228723
rect 304490 228683 418774 228711
rect 304490 228671 304496 228683
rect 418768 228671 418774 228683
rect 418826 228671 418832 228723
rect 455056 228671 455062 228723
rect 455114 228711 455120 228723
rect 455728 228711 455734 228723
rect 455114 228683 455734 228711
rect 455114 228671 455120 228683
rect 455728 228671 455734 228683
rect 455786 228671 455792 228723
rect 230608 228597 230614 228649
rect 230666 228637 230672 228649
rect 270736 228637 270742 228649
rect 230666 228609 270742 228637
rect 230666 228597 230672 228609
rect 270736 228597 270742 228609
rect 270794 228597 270800 228649
rect 291472 228597 291478 228649
rect 291530 228637 291536 228649
rect 382960 228637 382966 228649
rect 291530 228609 382966 228637
rect 291530 228597 291536 228609
rect 382960 228597 382966 228609
rect 383018 228597 383024 228649
rect 407536 228597 407542 228649
rect 407594 228637 407600 228649
rect 517648 228637 517654 228649
rect 407594 228609 517654 228637
rect 407594 228597 407600 228609
rect 517648 228597 517654 228609
rect 517706 228597 517712 228649
rect 190192 228523 190198 228575
rect 190250 228563 190256 228575
rect 192304 228563 192310 228575
rect 190250 228535 192310 228563
rect 190250 228523 190256 228535
rect 192304 228523 192310 228535
rect 192362 228523 192368 228575
rect 228784 228523 228790 228575
rect 228842 228563 228848 228575
rect 266224 228563 266230 228575
rect 228842 228535 266230 228563
rect 228842 228523 228848 228535
rect 266224 228523 266230 228535
rect 266282 228523 266288 228575
rect 266320 228523 266326 228575
rect 266378 228563 266384 228575
rect 301744 228563 301750 228575
rect 266378 228535 301750 228563
rect 266378 228523 266384 228535
rect 301744 228523 301750 228535
rect 301802 228523 301808 228575
rect 303472 228523 303478 228575
rect 303530 228563 303536 228575
rect 413488 228563 413494 228575
rect 303530 228535 413494 228563
rect 303530 228523 303536 228535
rect 413488 228523 413494 228535
rect 413546 228523 413552 228575
rect 455152 228523 455158 228575
rect 455210 228563 455216 228575
rect 456496 228563 456502 228575
rect 455210 228535 456502 228563
rect 455210 228523 455216 228535
rect 456496 228523 456502 228535
rect 456554 228523 456560 228575
rect 535792 228523 535798 228575
rect 535850 228563 535856 228575
rect 538000 228563 538006 228575
rect 535850 228535 538006 228563
rect 535850 228523 535856 228535
rect 538000 228523 538006 228535
rect 538058 228523 538064 228575
rect 544336 228523 544342 228575
rect 544394 228563 544400 228575
rect 547120 228563 547126 228575
rect 544394 228535 547126 228563
rect 544394 228523 544400 228535
rect 547120 228523 547126 228535
rect 547178 228523 547184 228575
rect 556144 228523 556150 228575
rect 556202 228563 556208 228575
rect 557680 228563 557686 228575
rect 556202 228535 557686 228563
rect 556202 228523 556208 228535
rect 557680 228523 557686 228535
rect 557738 228523 557744 228575
rect 567376 228523 567382 228575
rect 567434 228563 567440 228575
rect 569008 228563 569014 228575
rect 567434 228535 569014 228563
rect 567434 228523 567440 228535
rect 569008 228523 569014 228535
rect 569066 228523 569072 228575
rect 224368 228449 224374 228501
rect 224426 228489 224432 228501
rect 258736 228489 258742 228501
rect 224426 228461 258742 228489
rect 224426 228449 224432 228461
rect 258736 228449 258742 228461
rect 258794 228449 258800 228501
rect 260464 228449 260470 228501
rect 260522 228489 260528 228501
rect 286672 228489 286678 228501
rect 260522 228461 286678 228489
rect 260522 228449 260528 228461
rect 286672 228449 286678 228461
rect 286730 228449 286736 228501
rect 289360 228449 289366 228501
rect 289418 228489 289424 228501
rect 380080 228489 380086 228501
rect 289418 228461 380086 228489
rect 289418 228449 289424 228461
rect 380080 228449 380086 228461
rect 380138 228449 380144 228501
rect 405328 228449 405334 228501
rect 405386 228489 405392 228501
rect 502576 228489 502582 228501
rect 405386 228461 502582 228489
rect 405386 228449 405392 228461
rect 502576 228449 502582 228461
rect 502634 228449 502640 228501
rect 250576 228375 250582 228427
rect 250634 228415 250640 228427
rect 277552 228415 277558 228427
rect 250634 228387 277558 228415
rect 250634 228375 250640 228387
rect 277552 228375 277558 228387
rect 277610 228375 277616 228427
rect 288016 228375 288022 228427
rect 288074 228415 288080 228427
rect 328912 228415 328918 228427
rect 288074 228387 328918 228415
rect 288074 228375 288080 228387
rect 328912 228375 328918 228387
rect 328970 228375 328976 228427
rect 331120 228375 331126 228427
rect 331178 228415 331184 228427
rect 467056 228415 467062 228427
rect 331178 228387 467062 228415
rect 331178 228375 331184 228387
rect 467056 228375 467062 228387
rect 467114 228375 467120 228427
rect 535792 228375 535798 228427
rect 535850 228415 535856 228427
rect 537904 228415 537910 228427
rect 535850 228387 537910 228415
rect 535850 228375 535856 228387
rect 537904 228375 537910 228387
rect 537962 228375 537968 228427
rect 260752 228301 260758 228353
rect 260810 228341 260816 228353
rect 292624 228341 292630 228353
rect 260810 228313 292630 228341
rect 260810 228301 260816 228313
rect 292624 228301 292630 228313
rect 292682 228301 292688 228353
rect 293872 228301 293878 228353
rect 293930 228341 293936 228353
rect 380272 228341 380278 228353
rect 293930 228313 380278 228341
rect 293930 228301 293936 228313
rect 380272 228301 380278 228313
rect 380330 228301 380336 228353
rect 391696 228301 391702 228353
rect 391754 228341 391760 228353
rect 476944 228341 476950 228353
rect 391754 228313 476950 228341
rect 391754 228301 391760 228313
rect 476944 228301 476950 228313
rect 477002 228301 477008 228353
rect 270832 228227 270838 228279
rect 270890 228267 270896 228279
rect 313840 228267 313846 228279
rect 270890 228239 313846 228267
rect 270890 228227 270896 228239
rect 313840 228227 313846 228239
rect 313898 228227 313904 228279
rect 313936 228227 313942 228279
rect 313994 228267 314000 228279
rect 392368 228267 392374 228279
rect 313994 228239 392374 228267
rect 313994 228227 314000 228239
rect 392368 228227 392374 228239
rect 392426 228227 392432 228279
rect 392464 228227 392470 228279
rect 392522 228267 392528 228279
rect 461872 228267 461878 228279
rect 392522 228239 461878 228267
rect 392522 228227 392528 228239
rect 461872 228227 461878 228239
rect 461930 228227 461936 228279
rect 267952 228153 267958 228205
rect 268010 228193 268016 228205
rect 307696 228193 307702 228205
rect 268010 228165 307702 228193
rect 268010 228153 268016 228165
rect 307696 228153 307702 228165
rect 307754 228153 307760 228205
rect 311056 228153 311062 228205
rect 311114 228193 311120 228205
rect 383248 228193 383254 228205
rect 311114 228165 383254 228193
rect 311114 228153 311120 228165
rect 383248 228153 383254 228165
rect 383306 228153 383312 228205
rect 394672 228153 394678 228205
rect 394730 228193 394736 228205
rect 437680 228193 437686 228205
rect 394730 228165 437686 228193
rect 394730 228153 394736 228165
rect 437680 228153 437686 228165
rect 437738 228153 437744 228205
rect 269488 228079 269494 228131
rect 269546 228119 269552 228131
rect 322960 228119 322966 228131
rect 269546 228091 322966 228119
rect 269546 228079 269552 228091
rect 322960 228079 322966 228091
rect 323018 228079 323024 228131
rect 344080 228079 344086 228131
rect 344138 228119 344144 228131
rect 412720 228119 412726 228131
rect 344138 228091 412726 228119
rect 344138 228079 344144 228091
rect 412720 228079 412726 228091
rect 412778 228079 412784 228131
rect 258064 228005 258070 228057
rect 258122 228045 258128 228057
rect 280624 228045 280630 228057
rect 258122 228017 280630 228045
rect 258122 228005 258128 228017
rect 280624 228005 280630 228017
rect 280682 228005 280688 228057
rect 290992 228005 290998 228057
rect 291050 228045 291056 228057
rect 341008 228045 341014 228057
rect 291050 228017 341014 228045
rect 291050 228005 291056 228017
rect 341008 228005 341014 228017
rect 341066 228005 341072 228057
rect 341200 228005 341206 228057
rect 341258 228045 341264 228057
rect 398320 228045 398326 228057
rect 341258 228017 398326 228045
rect 341258 228005 341264 228017
rect 398320 228005 398326 228017
rect 398378 228005 398384 228057
rect 263824 227931 263830 227983
rect 263882 227971 263888 227983
rect 295696 227971 295702 227983
rect 263882 227943 295702 227971
rect 263882 227931 263888 227943
rect 295696 227931 295702 227943
rect 295754 227931 295760 227983
rect 308272 227931 308278 227983
rect 308330 227971 308336 227983
rect 359152 227971 359158 227983
rect 308330 227943 359158 227971
rect 308330 227931 308336 227943
rect 359152 227931 359158 227943
rect 359210 227931 359216 227983
rect 368848 227931 368854 227983
rect 368906 227971 368912 227983
rect 425584 227971 425590 227983
rect 368906 227943 425590 227971
rect 368906 227931 368912 227943
rect 425584 227931 425590 227943
rect 425642 227931 425648 227983
rect 293776 227857 293782 227909
rect 293834 227897 293840 227909
rect 343984 227897 343990 227909
rect 293834 227869 343990 227897
rect 293834 227857 293840 227869
rect 343984 227857 343990 227869
rect 344042 227857 344048 227909
rect 302224 227783 302230 227835
rect 302282 227823 302288 227835
rect 350032 227823 350038 227835
rect 302282 227795 350038 227823
rect 302282 227783 302288 227795
rect 350032 227783 350038 227795
rect 350090 227783 350096 227835
rect 247024 227709 247030 227761
rect 247082 227749 247088 227761
rect 303952 227749 303958 227761
rect 247082 227721 303958 227749
rect 247082 227709 247088 227721
rect 303952 227709 303958 227721
rect 304010 227709 304016 227761
rect 304720 227709 304726 227761
rect 304778 227749 304784 227761
rect 353104 227749 353110 227761
rect 304778 227721 353110 227749
rect 304778 227709 304784 227721
rect 353104 227709 353110 227721
rect 353162 227709 353168 227761
rect 387760 227709 387766 227761
rect 387818 227749 387824 227761
rect 396208 227749 396214 227761
rect 387818 227721 396214 227749
rect 387818 227709 387824 227721
rect 396208 227709 396214 227721
rect 396266 227709 396272 227761
rect 281488 227635 281494 227687
rect 281546 227675 281552 227687
rect 325840 227675 325846 227687
rect 281546 227647 325846 227675
rect 281546 227635 281552 227647
rect 325840 227635 325846 227647
rect 325898 227635 325904 227687
rect 149392 227561 149398 227613
rect 149450 227601 149456 227613
rect 177136 227601 177142 227613
rect 149450 227573 177142 227601
rect 149450 227561 149456 227573
rect 177136 227561 177142 227573
rect 177194 227561 177200 227613
rect 278032 227561 278038 227613
rect 278090 227601 278096 227613
rect 319888 227601 319894 227613
rect 278090 227573 319894 227601
rect 278090 227561 278096 227573
rect 319888 227561 319894 227573
rect 319946 227561 319952 227613
rect 319984 227561 319990 227613
rect 320042 227601 320048 227613
rect 403696 227601 403702 227613
rect 320042 227573 403702 227601
rect 320042 227561 320048 227573
rect 403696 227561 403702 227573
rect 403754 227561 403760 227613
rect 423280 227561 423286 227613
rect 423338 227601 423344 227613
rect 433168 227601 433174 227613
rect 423338 227573 433174 227601
rect 423338 227561 423344 227573
rect 433168 227561 433174 227573
rect 433226 227561 433232 227613
rect 187120 227487 187126 227539
rect 187178 227527 187184 227539
rect 190768 227527 190774 227539
rect 187178 227499 190774 227527
rect 187178 227487 187184 227499
rect 190768 227487 190774 227499
rect 190826 227487 190832 227539
rect 216112 227487 216118 227539
rect 216170 227527 216176 227539
rect 239824 227527 239830 227539
rect 216170 227499 239830 227527
rect 216170 227487 216176 227499
rect 239824 227487 239830 227499
rect 239882 227487 239888 227539
rect 249328 227487 249334 227539
rect 249386 227527 249392 227539
rect 306256 227527 306262 227539
rect 249386 227499 306262 227527
rect 249386 227487 249392 227499
rect 306256 227487 306262 227499
rect 306314 227487 306320 227539
rect 311248 227487 311254 227539
rect 311306 227527 311312 227539
rect 375760 227527 375766 227539
rect 311306 227499 375766 227527
rect 311306 227487 311312 227499
rect 375760 227487 375766 227499
rect 375818 227487 375824 227539
rect 389488 227487 389494 227539
rect 389546 227527 389552 227539
rect 587152 227527 587158 227539
rect 389546 227499 587158 227527
rect 389546 227487 389552 227499
rect 587152 227487 587158 227499
rect 587210 227487 587216 227539
rect 590704 227487 590710 227539
rect 590762 227527 590768 227539
rect 594640 227527 594646 227539
rect 590762 227499 594646 227527
rect 590762 227487 590768 227499
rect 594640 227487 594646 227499
rect 594698 227487 594704 227539
rect 629296 227487 629302 227539
rect 629354 227527 629360 227539
rect 634000 227527 634006 227539
rect 629354 227499 634006 227527
rect 629354 227487 629360 227499
rect 634000 227487 634006 227499
rect 634058 227487 634064 227539
rect 213040 227413 213046 227465
rect 213098 227453 213104 227465
rect 233776 227453 233782 227465
rect 213098 227425 233782 227453
rect 213098 227413 213104 227425
rect 233776 227413 233782 227425
rect 233834 227413 233840 227465
rect 238768 227413 238774 227465
rect 238826 227453 238832 227465
rect 252208 227453 252214 227465
rect 238826 227425 252214 227453
rect 238826 227413 238832 227425
rect 252208 227413 252214 227425
rect 252266 227413 252272 227465
rect 253840 227413 253846 227465
rect 253898 227453 253904 227465
rect 315376 227453 315382 227465
rect 253898 227425 315382 227453
rect 253898 227413 253904 227425
rect 315376 227413 315382 227425
rect 315434 227413 315440 227465
rect 318160 227413 318166 227465
rect 318218 227453 318224 227465
rect 381808 227453 381814 227465
rect 318218 227425 381814 227453
rect 318218 227413 318224 227425
rect 381808 227413 381814 227425
rect 381866 227413 381872 227465
rect 390448 227413 390454 227465
rect 390506 227453 390512 227465
rect 390506 227425 588542 227453
rect 390506 227413 390512 227425
rect 217456 227339 217462 227391
rect 217514 227379 217520 227391
rect 241264 227379 241270 227391
rect 217514 227351 241270 227379
rect 217514 227339 217520 227351
rect 241264 227339 241270 227351
rect 241322 227339 241328 227391
rect 244720 227339 244726 227391
rect 244778 227379 244784 227391
rect 254896 227379 254902 227391
rect 244778 227351 254902 227379
rect 244778 227339 244784 227351
rect 254896 227339 254902 227351
rect 254954 227339 254960 227391
rect 311152 227339 311158 227391
rect 311210 227379 311216 227391
rect 384016 227379 384022 227391
rect 311210 227351 384022 227379
rect 311210 227339 311216 227351
rect 384016 227339 384022 227351
rect 384074 227339 384080 227391
rect 388528 227339 388534 227391
rect 388586 227379 388592 227391
rect 585616 227379 585622 227391
rect 388586 227351 585622 227379
rect 388586 227339 388592 227351
rect 585616 227339 585622 227351
rect 585674 227339 585680 227391
rect 588514 227379 588542 227425
rect 588592 227413 588598 227465
rect 588650 227453 588656 227465
rect 600784 227453 600790 227465
rect 588650 227425 600790 227453
rect 588650 227413 588656 227425
rect 600784 227413 600790 227425
rect 600842 227413 600848 227465
rect 606352 227413 606358 227465
rect 606410 227453 606416 227465
rect 638512 227453 638518 227465
rect 606410 227425 638518 227453
rect 606410 227413 606416 227425
rect 638512 227413 638518 227425
rect 638570 227413 638576 227465
rect 589360 227379 589366 227391
rect 588514 227351 589366 227379
rect 589360 227339 589366 227351
rect 589418 227339 589424 227391
rect 219472 227265 219478 227317
rect 219530 227305 219536 227317
rect 245872 227305 245878 227317
rect 219530 227277 245878 227305
rect 219530 227265 219536 227277
rect 245872 227265 245878 227277
rect 245930 227265 245936 227317
rect 275056 227265 275062 227317
rect 275114 227305 275120 227317
rect 348592 227305 348598 227317
rect 275114 227277 348598 227305
rect 275114 227265 275120 227277
rect 348592 227265 348598 227277
rect 348650 227265 348656 227317
rect 388912 227265 388918 227317
rect 388970 227305 388976 227317
rect 586384 227305 586390 227317
rect 388970 227277 586390 227305
rect 388970 227265 388976 227277
rect 586384 227265 586390 227277
rect 586442 227265 586448 227317
rect 588784 227265 588790 227317
rect 588842 227305 588848 227317
rect 626416 227305 626422 227317
rect 588842 227277 626422 227305
rect 588842 227265 588848 227277
rect 626416 227265 626422 227277
rect 626474 227265 626480 227317
rect 217840 227191 217846 227243
rect 217898 227231 217904 227243
rect 242896 227231 242902 227243
rect 217898 227203 242902 227231
rect 217898 227191 217904 227203
rect 242896 227191 242902 227203
rect 242954 227191 242960 227243
rect 271984 227191 271990 227243
rect 272042 227231 272048 227243
rect 351568 227231 351574 227243
rect 272042 227203 351574 227231
rect 272042 227191 272048 227203
rect 351568 227191 351574 227203
rect 351626 227191 351632 227243
rect 398896 227191 398902 227243
rect 398954 227231 398960 227243
rect 584848 227231 584854 227243
rect 398954 227203 584854 227231
rect 398954 227191 398960 227203
rect 584848 227191 584854 227203
rect 584906 227191 584912 227243
rect 587440 227191 587446 227243
rect 587498 227231 587504 227243
rect 630160 227231 630166 227243
rect 587498 227203 630166 227231
rect 587498 227191 587504 227203
rect 630160 227191 630166 227203
rect 630218 227191 630224 227243
rect 220336 227117 220342 227169
rect 220394 227157 220400 227169
rect 247408 227157 247414 227169
rect 220394 227129 247414 227157
rect 220394 227117 220400 227129
rect 247408 227117 247414 227129
rect 247466 227117 247472 227169
rect 264688 227117 264694 227169
rect 264746 227157 264752 227169
rect 288112 227157 288118 227169
rect 264746 227129 288118 227157
rect 264746 227117 264752 227129
rect 288112 227117 288118 227129
rect 288170 227117 288176 227169
rect 289648 227117 289654 227169
rect 289706 227157 289712 227169
rect 369616 227157 369622 227169
rect 289706 227129 369622 227157
rect 289706 227117 289712 227129
rect 369616 227117 369622 227129
rect 369674 227117 369680 227169
rect 390064 227117 390070 227169
rect 390122 227157 390128 227169
rect 588592 227157 588598 227169
rect 390122 227129 588598 227157
rect 390122 227117 390128 227129
rect 588592 227117 588598 227129
rect 588650 227117 588656 227169
rect 590896 227117 590902 227169
rect 590954 227157 590960 227169
rect 630928 227157 630934 227169
rect 590954 227129 630934 227157
rect 590954 227117 590960 227129
rect 630928 227117 630934 227129
rect 630986 227117 630992 227169
rect 215728 227043 215734 227095
rect 215786 227083 215792 227095
rect 238384 227083 238390 227095
rect 215786 227055 238390 227083
rect 215786 227043 215792 227055
rect 238384 227043 238390 227055
rect 238442 227043 238448 227095
rect 276688 227043 276694 227095
rect 276746 227083 276752 227095
rect 360592 227083 360598 227095
rect 276746 227055 360598 227083
rect 276746 227043 276752 227055
rect 360592 227043 360598 227055
rect 360650 227043 360656 227095
rect 390832 227043 390838 227095
rect 390890 227083 390896 227095
rect 590128 227083 590134 227095
rect 390890 227055 590134 227083
rect 390890 227043 390896 227055
rect 590128 227043 590134 227055
rect 590186 227043 590192 227095
rect 590416 227043 590422 227095
rect 590474 227083 590480 227095
rect 632368 227083 632374 227095
rect 590474 227055 632374 227083
rect 590474 227043 590480 227055
rect 632368 227043 632374 227055
rect 632426 227043 632432 227095
rect 238096 226969 238102 227021
rect 238154 227009 238160 227021
rect 264016 227009 264022 227021
rect 238154 226981 264022 227009
rect 238154 226969 238160 226981
rect 264016 226969 264022 226981
rect 264074 226969 264080 227021
rect 275248 226969 275254 227021
rect 275306 227009 275312 227021
rect 357616 227009 357622 227021
rect 275306 226981 357622 227009
rect 275306 226969 275312 226981
rect 357616 226969 357622 226981
rect 357674 226969 357680 227021
rect 359824 226969 359830 227021
rect 359882 227009 359888 227021
rect 359882 226981 392414 227009
rect 359882 226969 359888 226981
rect 221680 226895 221686 226947
rect 221738 226935 221744 226947
rect 250384 226935 250390 226947
rect 221738 226907 250390 226935
rect 221738 226895 221744 226907
rect 250384 226895 250390 226907
rect 250442 226895 250448 226947
rect 253552 226895 253558 226947
rect 253610 226935 253616 226947
rect 266992 226935 266998 226947
rect 253610 226907 266998 226935
rect 253610 226895 253616 226907
rect 266992 226895 266998 226907
rect 267050 226895 267056 226947
rect 273424 226895 273430 226947
rect 273482 226935 273488 226947
rect 354544 226935 354550 226947
rect 273482 226907 354550 226935
rect 273482 226895 273488 226907
rect 354544 226895 354550 226907
rect 354602 226895 354608 226947
rect 354640 226895 354646 226947
rect 354698 226935 354704 226947
rect 392176 226935 392182 226947
rect 354698 226907 392182 226935
rect 354698 226895 354704 226907
rect 392176 226895 392182 226907
rect 392234 226895 392240 226947
rect 392386 226935 392414 226981
rect 392656 226969 392662 227021
rect 392714 227009 392720 227021
rect 593968 227009 593974 227021
rect 392714 226981 593974 227009
rect 392714 226969 392720 226981
rect 593968 226969 593974 226981
rect 594026 226969 594032 227021
rect 599152 226969 599158 227021
rect 599210 226969 599216 227021
rect 603376 226969 603382 227021
rect 603434 227009 603440 227021
rect 636880 227009 636886 227021
rect 603434 226981 636886 227009
rect 603434 226969 603440 226981
rect 636880 226969 636886 226981
rect 636938 226969 636944 227021
rect 393136 226935 393142 226947
rect 392386 226907 393142 226935
rect 393136 226895 393142 226907
rect 393194 226895 393200 226947
rect 587344 226895 587350 226947
rect 587402 226935 587408 226947
rect 598480 226935 598486 226947
rect 587402 226907 598486 226935
rect 587402 226895 587408 226907
rect 598480 226895 598486 226907
rect 598538 226895 598544 226947
rect 599170 226935 599198 226969
rect 633136 226935 633142 226947
rect 599170 226907 633142 226935
rect 633136 226895 633142 226907
rect 633194 226895 633200 226947
rect 224944 226821 224950 226873
rect 225002 226861 225008 226873
rect 256432 226861 256438 226873
rect 225002 226833 256438 226861
rect 225002 226821 225008 226833
rect 256432 226821 256438 226833
rect 256490 226821 256496 226873
rect 324208 226821 324214 226873
rect 324266 226861 324272 226873
rect 339472 226861 339478 226873
rect 324266 226833 339478 226861
rect 324266 226821 324272 226833
rect 339472 226821 339478 226833
rect 339530 226821 339536 226873
rect 365104 226821 365110 226873
rect 365162 226861 365168 226873
rect 365162 226833 395486 226861
rect 365162 226821 365168 226833
rect 223312 226747 223318 226799
rect 223370 226787 223376 226799
rect 253456 226787 253462 226799
rect 223370 226759 253462 226787
rect 223370 226747 223376 226759
rect 253456 226747 253462 226759
rect 253514 226747 253520 226799
rect 279760 226747 279766 226799
rect 279818 226787 279824 226799
rect 298192 226787 298198 226799
rect 279818 226759 298198 226787
rect 279818 226747 279824 226759
rect 298192 226747 298198 226759
rect 298250 226747 298256 226799
rect 298384 226747 298390 226799
rect 298442 226787 298448 226799
rect 366736 226787 366742 226799
rect 298442 226759 366742 226787
rect 298442 226747 298448 226759
rect 366736 226747 366742 226759
rect 366794 226747 366800 226799
rect 372688 226787 372694 226799
rect 367042 226759 372694 226787
rect 226576 226673 226582 226725
rect 226634 226713 226640 226725
rect 259408 226713 259414 226725
rect 226634 226685 259414 226713
rect 226634 226673 226640 226685
rect 259408 226673 259414 226685
rect 259466 226673 259472 226725
rect 284656 226673 284662 226725
rect 284714 226713 284720 226725
rect 298096 226713 298102 226725
rect 284714 226685 298102 226713
rect 284714 226673 284720 226685
rect 298096 226673 298102 226685
rect 298154 226673 298160 226725
rect 300592 226673 300598 226725
rect 300650 226713 300656 226725
rect 367042 226713 367070 226759
rect 372688 226747 372694 226759
rect 372746 226747 372752 226799
rect 374608 226747 374614 226799
rect 374666 226787 374672 226799
rect 391504 226787 391510 226799
rect 374666 226759 391510 226787
rect 374666 226747 374672 226759
rect 391504 226747 391510 226759
rect 391562 226747 391568 226799
rect 395458 226787 395486 226833
rect 395536 226821 395542 226873
rect 395594 226861 395600 226873
rect 599152 226861 599158 226873
rect 395594 226833 599158 226861
rect 395594 226821 395600 226833
rect 599152 226821 599158 226833
rect 599210 226821 599216 226873
rect 600400 226821 600406 226873
rect 600458 226861 600464 226873
rect 634672 226861 634678 226873
rect 600458 226833 634678 226861
rect 600458 226821 600464 226833
rect 634672 226821 634678 226833
rect 634730 226821 634736 226873
rect 396112 226787 396118 226799
rect 395458 226759 396118 226787
rect 396112 226747 396118 226759
rect 396170 226747 396176 226799
rect 400816 226747 400822 226799
rect 400874 226787 400880 226799
rect 419152 226787 419158 226799
rect 400874 226759 419158 226787
rect 400874 226747 400880 226759
rect 419152 226747 419158 226759
rect 419210 226747 419216 226799
rect 419248 226747 419254 226799
rect 419306 226787 419312 226799
rect 419306 226759 603230 226787
rect 419306 226747 419312 226759
rect 378736 226713 378742 226725
rect 300650 226685 367070 226713
rect 367138 226685 378742 226713
rect 300650 226673 300656 226685
rect 227920 226599 227926 226651
rect 227978 226639 227984 226651
rect 262480 226639 262486 226651
rect 227978 226611 262486 226639
rect 227978 226599 227984 226611
rect 262480 226599 262486 226611
rect 262538 226599 262544 226651
rect 264880 226599 264886 226651
rect 264938 226639 264944 226651
rect 276112 226639 276118 226651
rect 264938 226611 276118 226639
rect 264938 226599 264944 226611
rect 276112 226599 276118 226611
rect 276170 226599 276176 226651
rect 285712 226599 285718 226651
rect 285770 226639 285776 226651
rect 367138 226639 367166 226685
rect 378736 226673 378742 226685
rect 378794 226673 378800 226725
rect 380272 226673 380278 226725
rect 380330 226713 380336 226725
rect 397648 226713 397654 226725
rect 380330 226685 397654 226713
rect 380330 226673 380336 226685
rect 397648 226673 397654 226685
rect 397706 226673 397712 226725
rect 402160 226673 402166 226725
rect 402218 226713 402224 226725
rect 418864 226713 418870 226725
rect 402218 226685 418870 226713
rect 402218 226673 402224 226685
rect 418864 226673 418870 226685
rect 418922 226673 418928 226725
rect 423346 226685 429134 226713
rect 285770 226611 367166 226639
rect 285770 226599 285776 226611
rect 374416 226599 374422 226651
rect 374474 226639 374480 226651
rect 385552 226639 385558 226651
rect 374474 226611 385558 226639
rect 374474 226599 374480 226611
rect 385552 226599 385558 226611
rect 385610 226599 385616 226651
rect 397168 226599 397174 226651
rect 397226 226639 397232 226651
rect 423346 226639 423374 226685
rect 397226 226611 423374 226639
rect 429106 226639 429134 226685
rect 587632 226673 587638 226725
rect 587690 226713 587696 226725
rect 602224 226713 602230 226725
rect 587690 226685 602230 226713
rect 587690 226673 587696 226685
rect 602224 226673 602230 226685
rect 602282 226673 602288 226725
rect 603202 226713 603230 226759
rect 603280 226747 603286 226799
rect 603338 226787 603344 226799
rect 637744 226787 637750 226799
rect 603338 226759 637750 226787
rect 603338 226747 603344 226759
rect 637744 226747 637750 226759
rect 637802 226747 637808 226799
rect 603664 226713 603670 226725
rect 603202 226685 603670 226713
rect 603664 226673 603670 226685
rect 603722 226673 603728 226725
rect 606256 226673 606262 226725
rect 606314 226713 606320 226725
rect 639184 226713 639190 226725
rect 606314 226685 639190 226713
rect 606314 226673 606320 226685
rect 639184 226673 639190 226685
rect 639242 226673 639248 226725
rect 602992 226639 602998 226651
rect 429106 226611 602998 226639
rect 397226 226599 397232 226611
rect 602992 226599 602998 226611
rect 603050 226599 603056 226651
rect 606160 226599 606166 226651
rect 606218 226639 606224 226651
rect 639952 226639 639958 226651
rect 606218 226611 639958 226639
rect 606218 226599 606224 226611
rect 639952 226599 639958 226611
rect 640010 226599 640016 226651
rect 229552 226525 229558 226577
rect 229610 226565 229616 226577
rect 265552 226565 265558 226577
rect 229610 226537 265558 226565
rect 229610 226525 229616 226537
rect 265552 226525 265558 226537
rect 265610 226525 265616 226577
rect 271024 226525 271030 226577
rect 271082 226565 271088 226577
rect 294256 226565 294262 226577
rect 271082 226537 294262 226565
rect 271082 226525 271088 226537
rect 294256 226525 294262 226537
rect 294314 226525 294320 226577
rect 297424 226525 297430 226577
rect 297482 226565 297488 226577
rect 390064 226565 390070 226577
rect 297482 226537 390070 226565
rect 297482 226525 297488 226537
rect 390064 226525 390070 226537
rect 390122 226525 390128 226577
rect 392176 226525 392182 226577
rect 392234 226565 392240 226577
rect 392234 226537 402494 226565
rect 392234 226525 392240 226537
rect 231088 226451 231094 226503
rect 231146 226491 231152 226503
rect 268528 226491 268534 226503
rect 231146 226463 268534 226491
rect 231146 226451 231152 226463
rect 268528 226451 268534 226463
rect 268586 226451 268592 226503
rect 288496 226451 288502 226503
rect 288554 226491 288560 226503
rect 384784 226491 384790 226503
rect 288554 226463 384790 226491
rect 288554 226451 288560 226463
rect 384784 226451 384790 226463
rect 384842 226451 384848 226503
rect 385744 226451 385750 226503
rect 385802 226491 385808 226503
rect 398800 226491 398806 226503
rect 385802 226463 398806 226491
rect 385802 226451 385808 226463
rect 398800 226451 398806 226463
rect 398858 226451 398864 226503
rect 232528 226377 232534 226429
rect 232586 226417 232592 226429
rect 271600 226417 271606 226429
rect 232586 226389 271606 226417
rect 232586 226377 232592 226389
rect 271600 226377 271606 226389
rect 271658 226377 271664 226429
rect 272848 226377 272854 226429
rect 272906 226417 272912 226429
rect 282544 226417 282550 226429
rect 272906 226389 282550 226417
rect 272906 226377 272912 226389
rect 282544 226377 282550 226389
rect 282602 226377 282608 226429
rect 298096 226377 298102 226429
rect 298154 226417 298160 226429
rect 378064 226417 378070 226429
rect 298154 226389 378070 226417
rect 298154 226377 298160 226389
rect 378064 226377 378070 226389
rect 378122 226377 378128 226429
rect 379888 226377 379894 226429
rect 379946 226417 379952 226429
rect 387760 226417 387766 226429
rect 379946 226389 387766 226417
rect 379946 226377 379952 226389
rect 387760 226377 387766 226389
rect 387818 226377 387824 226429
rect 388144 226377 388150 226429
rect 388202 226417 388208 226429
rect 398896 226417 398902 226429
rect 388202 226389 398902 226417
rect 388202 226377 388208 226389
rect 398896 226377 398902 226389
rect 398954 226377 398960 226429
rect 402466 226417 402494 226537
rect 402544 226525 402550 226577
rect 402602 226565 402608 226577
rect 402602 226537 419006 226565
rect 402602 226525 402608 226537
rect 404944 226451 404950 226503
rect 405002 226491 405008 226503
rect 405002 226463 418910 226491
rect 405002 226451 405008 226463
rect 408208 226417 408214 226429
rect 402466 226389 408214 226417
rect 408208 226377 408214 226389
rect 408266 226377 408272 226429
rect 213808 226303 213814 226355
rect 213866 226343 213872 226355
rect 237520 226343 237526 226355
rect 213866 226315 237526 226343
rect 213866 226303 213872 226315
rect 237520 226303 237526 226315
rect 237578 226303 237584 226355
rect 244816 226303 244822 226355
rect 244874 226343 244880 226355
rect 244874 226315 252158 226343
rect 244874 226303 244880 226315
rect 147088 226229 147094 226281
rect 147146 226269 147152 226281
rect 151312 226269 151318 226281
rect 147146 226241 151318 226269
rect 147146 226229 147152 226241
rect 151312 226229 151318 226241
rect 151370 226229 151376 226281
rect 217072 226229 217078 226281
rect 217130 226269 217136 226281
rect 243568 226269 243574 226281
rect 217130 226241 243574 226269
rect 217130 226229 217136 226241
rect 243568 226229 243574 226241
rect 243626 226229 243632 226281
rect 246544 226229 246550 226281
rect 246602 226269 246608 226281
rect 252130 226269 252158 226315
rect 252208 226303 252214 226355
rect 252266 226343 252272 226355
rect 285136 226343 285142 226355
rect 252266 226315 285142 226343
rect 252266 226303 252272 226315
rect 285136 226303 285142 226315
rect 285194 226303 285200 226355
rect 291568 226303 291574 226355
rect 291626 226343 291632 226355
rect 390832 226343 390838 226355
rect 291626 226315 390838 226343
rect 291626 226303 291632 226315
rect 390832 226303 390838 226315
rect 390890 226303 390896 226355
rect 402832 226343 402838 226355
rect 397762 226315 402838 226343
rect 297232 226269 297238 226281
rect 246602 226241 252062 226269
rect 252130 226241 297238 226269
rect 246602 226229 246608 226241
rect 42256 226155 42262 226207
rect 42314 226195 42320 226207
rect 45808 226195 45814 226207
rect 42314 226167 45814 226195
rect 42314 226155 42320 226167
rect 45808 226155 45814 226167
rect 45866 226155 45872 226207
rect 215632 226155 215638 226207
rect 215690 226195 215696 226207
rect 240592 226195 240598 226207
rect 215690 226167 240598 226195
rect 215690 226155 215696 226167
rect 240592 226155 240598 226167
rect 240650 226155 240656 226207
rect 243952 226155 243958 226207
rect 244010 226195 244016 226207
rect 251920 226195 251926 226207
rect 244010 226167 251926 226195
rect 244010 226155 244016 226167
rect 251920 226155 251926 226167
rect 251978 226155 251984 226207
rect 151120 226081 151126 226133
rect 151178 226121 151184 226133
rect 187120 226121 187126 226133
rect 151178 226093 187126 226121
rect 151178 226081 151184 226093
rect 187120 226081 187126 226093
rect 187178 226081 187184 226133
rect 218320 226081 218326 226133
rect 218378 226121 218384 226133
rect 246640 226121 246646 226133
rect 218378 226093 246646 226121
rect 218378 226081 218384 226093
rect 246640 226081 246646 226093
rect 246698 226081 246704 226133
rect 252034 226121 252062 226241
rect 297232 226229 297238 226241
rect 297290 226229 297296 226281
rect 297616 226229 297622 226281
rect 297674 226269 297680 226281
rect 397762 226269 397790 226315
rect 402832 226303 402838 226315
rect 402890 226303 402896 226355
rect 408016 226303 408022 226355
rect 408074 226343 408080 226355
rect 418882 226343 418910 226463
rect 418978 226417 419006 226537
rect 419152 226525 419158 226577
rect 419210 226565 419216 226577
rect 609808 226565 609814 226577
rect 419210 226537 609814 226565
rect 419210 226525 419216 226537
rect 609808 226525 609814 226537
rect 609866 226525 609872 226577
rect 419056 226451 419062 226503
rect 419114 226491 419120 226503
rect 612784 226491 612790 226503
rect 419114 226463 612790 226491
rect 419114 226451 419120 226463
rect 612784 226451 612790 226463
rect 612842 226451 612848 226503
rect 613552 226417 613558 226429
rect 418978 226389 613558 226417
rect 613552 226377 613558 226389
rect 613610 226377 613616 226429
rect 629200 226377 629206 226429
rect 629258 226417 629264 226429
rect 635440 226417 635446 226429
rect 629258 226389 635446 226417
rect 629258 226377 629264 226389
rect 635440 226377 635446 226389
rect 635498 226377 635504 226429
rect 618064 226343 618070 226355
rect 408074 226315 408974 226343
rect 418882 226315 618070 226343
rect 408074 226303 408080 226315
rect 297674 226241 397790 226269
rect 297674 226229 297680 226241
rect 397840 226229 397846 226281
rect 397898 226269 397904 226281
rect 400240 226269 400246 226281
rect 397898 226241 400246 226269
rect 397898 226229 397904 226241
rect 400240 226229 400246 226241
rect 400298 226229 400304 226281
rect 408946 226269 408974 226315
rect 618064 226303 618070 226315
rect 618122 226303 618128 226355
rect 624112 226269 624118 226281
rect 408946 226241 624118 226269
rect 624112 226229 624118 226241
rect 624170 226229 624176 226281
rect 252112 226155 252118 226207
rect 252170 226195 252176 226207
rect 291184 226195 291190 226207
rect 252170 226167 291190 226195
rect 252170 226155 252176 226167
rect 291184 226155 291190 226167
rect 291242 226155 291248 226207
rect 301264 226155 301270 226207
rect 301322 226195 301328 226207
rect 301322 226167 410366 226195
rect 301322 226155 301328 226167
rect 300208 226121 300214 226133
rect 252034 226093 300214 226121
rect 300208 226081 300214 226093
rect 300266 226081 300272 226133
rect 300688 226081 300694 226133
rect 300746 226121 300752 226133
rect 408976 226121 408982 226133
rect 300746 226093 408982 226121
rect 300746 226081 300752 226093
rect 408976 226081 408982 226093
rect 409034 226081 409040 226133
rect 410338 226121 410366 226167
rect 410416 226155 410422 226207
rect 410474 226195 410480 226207
rect 629392 226195 629398 226207
rect 410474 226167 629398 226195
rect 410474 226155 410480 226167
rect 629392 226155 629398 226167
rect 629450 226155 629456 226207
rect 411280 226121 411286 226133
rect 410338 226093 411286 226121
rect 411280 226081 411286 226093
rect 411338 226081 411344 226133
rect 411664 226081 411670 226133
rect 411722 226121 411728 226133
rect 631696 226121 631702 226133
rect 411722 226093 631702 226121
rect 411722 226081 411728 226093
rect 631696 226081 631702 226093
rect 631754 226081 631760 226133
rect 214576 226007 214582 226059
rect 214634 226047 214640 226059
rect 236848 226047 236854 226059
rect 214634 226019 236854 226047
rect 214634 226007 214640 226019
rect 236848 226007 236854 226019
rect 236906 226007 236912 226059
rect 241840 226007 241846 226059
rect 241898 226047 241904 226059
rect 248848 226047 248854 226059
rect 241898 226019 248854 226047
rect 241898 226007 241904 226019
rect 248848 226007 248854 226019
rect 248906 226007 248912 226059
rect 257104 226007 257110 226059
rect 257162 226047 257168 226059
rect 257162 226019 266846 226047
rect 257162 226007 257168 226019
rect 212368 225933 212374 225985
rect 212426 225973 212432 225985
rect 234544 225973 234550 225985
rect 212426 225945 234550 225973
rect 212426 225933 212432 225945
rect 234544 225933 234550 225945
rect 234602 225933 234608 225985
rect 236752 225933 236758 225985
rect 236810 225973 236816 225985
rect 261040 225973 261046 225985
rect 236810 225945 261046 225973
rect 236810 225933 236816 225945
rect 261040 225933 261046 225945
rect 261098 225933 261104 225985
rect 266818 225973 266846 226019
rect 266896 226007 266902 226059
rect 266954 226047 266960 226059
rect 279088 226047 279094 226059
rect 266954 226019 279094 226047
rect 266954 226007 266960 226019
rect 279088 226007 279094 226019
rect 279146 226007 279152 226059
rect 282544 226007 282550 226059
rect 282602 226047 282608 226059
rect 336400 226047 336406 226059
rect 282602 226019 336406 226047
rect 282602 226007 282608 226019
rect 336400 226007 336406 226019
rect 336458 226007 336464 226059
rect 379888 226047 379894 226059
rect 368626 226019 379894 226047
rect 321328 225973 321334 225985
rect 266818 225945 321334 225973
rect 321328 225933 321334 225945
rect 321386 225933 321392 225985
rect 334096 225933 334102 225985
rect 334154 225973 334160 225985
rect 368626 225973 368654 226019
rect 379888 226007 379894 226019
rect 379946 226007 379952 226059
rect 379984 226007 379990 226059
rect 380042 226047 380048 226059
rect 394576 226047 394582 226059
rect 380042 226019 394582 226047
rect 380042 226007 380048 226019
rect 394576 226007 394582 226019
rect 394634 226007 394640 226059
rect 398800 226007 398806 226059
rect 398858 226047 398864 226059
rect 579568 226047 579574 226059
rect 398858 226019 579574 226047
rect 398858 226007 398864 226019
rect 579568 226007 579574 226019
rect 579626 226007 579632 226059
rect 584560 226007 584566 226059
rect 584618 226047 584624 226059
rect 628624 226047 628630 226059
rect 584618 226019 628630 226047
rect 584618 226007 584624 226019
rect 628624 226007 628630 226019
rect 628682 226007 628688 226059
rect 334154 225945 368654 225973
rect 374338 225945 382910 225973
rect 334154 225933 334160 225945
rect 218800 225859 218806 225911
rect 218858 225899 218864 225911
rect 244336 225899 244342 225911
rect 218858 225871 244342 225899
rect 218858 225859 218864 225871
rect 244336 225859 244342 225871
rect 244394 225859 244400 225911
rect 262000 225859 262006 225911
rect 262058 225899 262064 225911
rect 273040 225899 273046 225911
rect 262058 225871 273046 225899
rect 262058 225859 262064 225871
rect 273040 225859 273046 225871
rect 273098 225859 273104 225911
rect 330448 225899 330454 225911
rect 278530 225871 330454 225899
rect 241744 225785 241750 225837
rect 241802 225825 241808 225837
rect 252112 225825 252118 225837
rect 241802 225797 252118 225825
rect 241802 225785 241808 225797
rect 252112 225785 252118 225797
rect 252170 225785 252176 225837
rect 267760 225785 267766 225837
rect 267818 225825 267824 225837
rect 278416 225825 278422 225837
rect 267818 225797 278422 225825
rect 267818 225785 267824 225797
rect 278416 225785 278422 225797
rect 278474 225785 278480 225837
rect 247696 225711 247702 225763
rect 247754 225751 247760 225763
rect 257968 225751 257974 225763
rect 247754 225723 257974 225751
rect 247754 225711 247760 225723
rect 257968 225711 257974 225723
rect 258026 225711 258032 225763
rect 269008 225711 269014 225763
rect 269066 225751 269072 225763
rect 278530 225751 278558 225871
rect 330448 225859 330454 225871
rect 330506 225859 330512 225911
rect 331408 225859 331414 225911
rect 331466 225899 331472 225911
rect 345520 225899 345526 225911
rect 331466 225871 345526 225899
rect 331466 225859 331472 225871
rect 345520 225859 345526 225871
rect 345578 225859 345584 225911
rect 346864 225859 346870 225911
rect 346922 225899 346928 225911
rect 374338 225899 374366 225945
rect 346922 225871 374366 225899
rect 346922 225859 346928 225871
rect 278608 225785 278614 225837
rect 278666 225825 278672 225837
rect 327376 225825 327382 225837
rect 278666 225797 327382 225825
rect 278666 225785 278672 225797
rect 327376 225785 327382 225797
rect 327434 225785 327440 225837
rect 374512 225785 374518 225837
rect 374570 225825 374576 225837
rect 382576 225825 382582 225837
rect 374570 225797 382582 225825
rect 374570 225785 374576 225797
rect 382576 225785 382582 225797
rect 382634 225785 382640 225837
rect 382882 225825 382910 225945
rect 382960 225933 382966 225985
rect 383018 225973 383024 225985
rect 388624 225973 388630 225985
rect 383018 225945 388630 225973
rect 383018 225933 383024 225945
rect 388624 225933 388630 225945
rect 388682 225933 388688 225985
rect 388720 225933 388726 225985
rect 388778 225973 388784 225985
rect 388778 225945 398846 225973
rect 388778 225933 388784 225945
rect 386992 225899 386998 225911
rect 385762 225871 386998 225899
rect 385762 225825 385790 225871
rect 386992 225859 386998 225871
rect 387050 225859 387056 225911
rect 387376 225859 387382 225911
rect 387434 225899 387440 225911
rect 398704 225899 398710 225911
rect 387434 225871 398710 225899
rect 387434 225859 387440 225871
rect 398704 225859 398710 225871
rect 398762 225859 398768 225911
rect 382882 225797 385790 225825
rect 385840 225785 385846 225837
rect 385898 225825 385904 225837
rect 398608 225825 398614 225837
rect 385898 225797 398614 225825
rect 385898 225785 385904 225797
rect 398608 225785 398614 225797
rect 398666 225785 398672 225837
rect 398818 225825 398846 225945
rect 398896 225933 398902 225985
rect 398954 225973 398960 225985
rect 582640 225973 582646 225985
rect 398954 225945 582646 225973
rect 398954 225933 398960 225945
rect 582640 225933 582646 225945
rect 582698 225933 582704 225985
rect 603472 225933 603478 225985
rect 603530 225973 603536 225985
rect 636208 225973 636214 225985
rect 603530 225945 636214 225973
rect 603530 225933 603536 225945
rect 636208 225933 636214 225945
rect 636266 225933 636272 225985
rect 400240 225859 400246 225911
rect 400298 225899 400304 225911
rect 419248 225899 419254 225911
rect 400298 225871 419254 225899
rect 400298 225859 400304 225871
rect 419248 225859 419254 225871
rect 419306 225859 419312 225911
rect 581104 225825 581110 225837
rect 398818 225797 581110 225825
rect 581104 225785 581110 225797
rect 581162 225785 581168 225837
rect 591472 225785 591478 225837
rect 591530 225825 591536 225837
rect 591530 225797 599054 225825
rect 591530 225785 591536 225797
rect 269066 225723 278558 225751
rect 269066 225711 269072 225723
rect 285040 225711 285046 225763
rect 285098 225751 285104 225763
rect 342544 225751 342550 225763
rect 285098 225723 342550 225751
rect 285098 225711 285104 225723
rect 342544 225711 342550 225723
rect 342602 225711 342608 225763
rect 365680 225711 365686 225763
rect 365738 225751 365744 225763
rect 393808 225751 393814 225763
rect 365738 225723 393814 225751
rect 365738 225711 365744 225723
rect 393808 225711 393814 225723
rect 393866 225711 393872 225763
rect 396208 225711 396214 225763
rect 396266 225751 396272 225763
rect 584080 225751 584086 225763
rect 396266 225723 584086 225751
rect 396266 225711 396272 225723
rect 584080 225711 584086 225723
rect 584138 225711 584144 225763
rect 587056 225711 587062 225763
rect 587114 225751 587120 225763
rect 595408 225751 595414 225763
rect 587114 225723 595414 225751
rect 587114 225711 587120 225723
rect 595408 225711 595414 225723
rect 595466 225711 595472 225763
rect 599026 225751 599054 225797
rect 627856 225751 627862 225763
rect 599026 225723 627862 225751
rect 627856 225711 627862 225723
rect 627914 225711 627920 225763
rect 278224 225637 278230 225689
rect 278282 225677 278288 225689
rect 318352 225677 318358 225689
rect 278282 225649 318358 225677
rect 278282 225637 278288 225649
rect 318352 225637 318358 225649
rect 318410 225637 318416 225689
rect 321712 225637 321718 225689
rect 321770 225677 321776 225689
rect 451216 225677 451222 225689
rect 321770 225649 451222 225677
rect 321770 225637 321776 225649
rect 451216 225637 451222 225649
rect 451274 225637 451280 225689
rect 273712 225563 273718 225615
rect 273770 225603 273776 225615
rect 309328 225603 309334 225615
rect 273770 225575 309334 225603
rect 273770 225563 273776 225575
rect 309328 225563 309334 225575
rect 309386 225563 309392 225615
rect 315760 225563 315766 225615
rect 315818 225603 315824 225615
rect 439120 225603 439126 225615
rect 315818 225575 439126 225603
rect 315818 225563 315824 225575
rect 439120 225563 439126 225575
rect 439178 225563 439184 225615
rect 273616 225489 273622 225541
rect 273674 225529 273680 225541
rect 303184 225529 303190 225541
rect 273674 225501 303190 225529
rect 273674 225489 273680 225501
rect 303184 225489 303190 225501
rect 303242 225489 303248 225541
rect 309904 225489 309910 225541
rect 309962 225529 309968 225541
rect 427024 225529 427030 225541
rect 309962 225501 427030 225529
rect 309962 225489 309968 225501
rect 427024 225489 427030 225501
rect 427082 225489 427088 225541
rect 585520 225489 585526 225541
rect 585578 225529 585584 225541
rect 592336 225529 592342 225541
rect 585578 225501 592342 225529
rect 585578 225489 585584 225501
rect 592336 225489 592342 225501
rect 592394 225489 592400 225541
rect 259024 225415 259030 225467
rect 259082 225455 259088 225467
rect 269968 225455 269974 225467
rect 259082 225427 269974 225455
rect 259082 225415 259088 225427
rect 269968 225415 269974 225427
rect 270026 225415 270032 225467
rect 306736 225415 306742 225467
rect 306794 225455 306800 225467
rect 420976 225455 420982 225467
rect 306794 225427 420982 225455
rect 306794 225415 306800 225427
rect 420976 225415 420982 225427
rect 421034 225415 421040 225467
rect 303856 225341 303862 225393
rect 303914 225381 303920 225393
rect 415024 225381 415030 225393
rect 303914 225353 415030 225381
rect 303914 225341 303920 225353
rect 415024 225341 415030 225353
rect 415082 225341 415088 225393
rect 302128 225267 302134 225319
rect 302186 225307 302192 225319
rect 411952 225307 411958 225319
rect 302186 225279 411958 225307
rect 302186 225267 302192 225279
rect 411952 225267 411958 225279
rect 412010 225267 412016 225319
rect 278704 225193 278710 225245
rect 278762 225233 278768 225245
rect 324400 225233 324406 225245
rect 278762 225205 324406 225233
rect 278762 225193 278768 225205
rect 324400 225193 324406 225205
rect 324458 225193 324464 225245
rect 351376 225193 351382 225245
rect 351434 225233 351440 225245
rect 418000 225233 418006 225245
rect 351434 225205 418006 225233
rect 351434 225193 351440 225205
rect 418000 225193 418006 225205
rect 418058 225193 418064 225245
rect 305104 225119 305110 225171
rect 305162 225159 305168 225171
rect 333520 225159 333526 225171
rect 305162 225131 333526 225159
rect 305162 225119 305168 225131
rect 333520 225119 333526 225131
rect 333578 225119 333584 225171
rect 339760 225119 339766 225171
rect 339818 225159 339824 225171
rect 399952 225159 399958 225171
rect 339818 225131 399958 225159
rect 339818 225119 339824 225131
rect 399952 225119 399958 225131
rect 400010 225119 400016 225171
rect 408880 225119 408886 225171
rect 408938 225159 408944 225171
rect 610480 225159 610486 225171
rect 408938 225131 610486 225159
rect 408938 225119 408944 225131
rect 610480 225119 610486 225131
rect 610538 225119 610544 225171
rect 252688 225045 252694 225097
rect 252746 225085 252752 225097
rect 312304 225085 312310 225097
rect 252746 225057 312310 225085
rect 252746 225045 252752 225057
rect 312304 225045 312310 225057
rect 312362 225045 312368 225097
rect 337648 225045 337654 225097
rect 337706 225085 337712 225097
rect 396880 225085 396886 225097
rect 337706 225057 396886 225085
rect 337706 225045 337712 225057
rect 396880 225045 396886 225057
rect 396938 225045 396944 225097
rect 398608 225045 398614 225097
rect 398666 225085 398672 225097
rect 398666 225057 399326 225085
rect 398666 225045 398672 225057
rect 348688 224971 348694 225023
rect 348746 225011 348752 225023
rect 399088 225011 399094 225023
rect 348746 224983 399094 225011
rect 348746 224971 348752 224983
rect 399088 224971 399094 224983
rect 399146 224971 399152 225023
rect 399298 225011 399326 225057
rect 399376 225045 399382 225097
rect 399434 225085 399440 225097
rect 606736 225085 606742 225097
rect 399434 225057 606742 225085
rect 399434 225045 399440 225057
rect 606736 225045 606742 225057
rect 606794 225045 606800 225097
rect 407440 225011 407446 225023
rect 399298 224983 407446 225011
rect 407440 224971 407446 224983
rect 407498 224971 407504 225023
rect 369424 224897 369430 224949
rect 369482 224937 369488 224949
rect 405136 224937 405142 224949
rect 369482 224909 405142 224937
rect 369482 224897 369488 224909
rect 405136 224897 405142 224909
rect 405194 224897 405200 224949
rect 149488 224823 149494 224875
rect 149546 224863 149552 224875
rect 174160 224863 174166 224875
rect 149546 224835 174166 224863
rect 149546 224823 149552 224835
rect 174160 224823 174166 224835
rect 174218 224823 174224 224875
rect 362800 224823 362806 224875
rect 362858 224863 362864 224875
rect 402160 224863 402166 224875
rect 362858 224835 402166 224863
rect 362858 224823 362864 224835
rect 402160 224823 402166 224835
rect 402218 224823 402224 224875
rect 149392 224749 149398 224801
rect 149450 224789 149456 224801
rect 159856 224789 159862 224801
rect 149450 224761 159862 224789
rect 149450 224749 149456 224761
rect 159856 224749 159862 224761
rect 159914 224749 159920 224801
rect 277936 224749 277942 224801
rect 277994 224789 278000 224801
rect 363664 224789 363670 224801
rect 277994 224761 363670 224789
rect 277994 224749 278000 224761
rect 363664 224749 363670 224761
rect 363722 224749 363728 224801
rect 371536 224749 371542 224801
rect 371594 224789 371600 224801
rect 379504 224789 379510 224801
rect 371594 224761 379510 224789
rect 371594 224749 371600 224761
rect 379504 224749 379510 224761
rect 379562 224749 379568 224801
rect 380080 224749 380086 224801
rect 380138 224789 380144 224801
rect 388624 224789 388630 224801
rect 380138 224761 388630 224789
rect 380138 224749 380144 224761
rect 388624 224749 388630 224761
rect 388682 224749 388688 224801
rect 388720 224749 388726 224801
rect 388778 224789 388784 224801
rect 389296 224789 389302 224801
rect 388778 224761 389302 224789
rect 388778 224749 388784 224761
rect 389296 224749 389302 224761
rect 389354 224749 389360 224801
rect 392272 224749 392278 224801
rect 392330 224789 392336 224801
rect 392330 224761 408974 224789
rect 392330 224749 392336 224761
rect 268624 224675 268630 224727
rect 268682 224715 268688 224727
rect 282064 224715 282070 224727
rect 268682 224687 282070 224715
rect 268682 224675 268688 224687
rect 282064 224675 282070 224687
rect 282122 224675 282128 224727
rect 362416 224675 362422 224727
rect 362474 224715 362480 224727
rect 369424 224715 369430 224727
rect 362474 224687 369430 224715
rect 362474 224675 362480 224687
rect 369424 224675 369430 224687
rect 369482 224675 369488 224727
rect 369520 224675 369526 224727
rect 369578 224715 369584 224727
rect 376432 224715 376438 224727
rect 369578 224687 376438 224715
rect 369578 224675 369584 224687
rect 376432 224675 376438 224687
rect 376490 224675 376496 224727
rect 382864 224675 382870 224727
rect 382922 224715 382928 224727
rect 386320 224715 386326 224727
rect 382922 224687 386326 224715
rect 382922 224675 382928 224687
rect 386320 224675 386326 224687
rect 386378 224675 386384 224727
rect 397456 224675 397462 224727
rect 397514 224715 397520 224727
rect 400624 224715 400630 224727
rect 397514 224687 400630 224715
rect 397514 224675 397520 224687
rect 400624 224675 400630 224687
rect 400682 224675 400688 224727
rect 408946 224715 408974 224761
rect 593104 224715 593110 224727
rect 408946 224687 593110 224715
rect 593104 224675 593110 224687
rect 593162 224675 593168 224727
rect 596080 224675 596086 224727
rect 596138 224715 596144 224727
rect 597712 224715 597718 224727
rect 596138 224687 597718 224715
rect 596138 224675 596144 224687
rect 597712 224675 597718 224687
rect 597770 224675 597776 224727
rect 316336 224601 316342 224653
rect 316394 224641 316400 224653
rect 441424 224641 441430 224653
rect 316394 224613 441430 224641
rect 316394 224601 316400 224613
rect 441424 224601 441430 224613
rect 441482 224601 441488 224653
rect 319312 224527 319318 224579
rect 319370 224567 319376 224579
rect 447472 224567 447478 224579
rect 319370 224539 447478 224567
rect 319370 224527 319376 224539
rect 447472 224527 447478 224539
rect 447530 224527 447536 224579
rect 323248 224453 323254 224505
rect 323306 224493 323312 224505
rect 452752 224493 452758 224505
rect 323306 224465 452758 224493
rect 323306 224453 323312 224465
rect 452752 224453 452758 224465
rect 452810 224453 452816 224505
rect 322288 224379 322294 224431
rect 322346 224419 322352 224431
rect 453424 224419 453430 224431
rect 322346 224391 453430 224419
rect 322346 224379 322352 224391
rect 453424 224379 453430 224391
rect 453482 224379 453488 224431
rect 325264 224305 325270 224357
rect 325322 224345 325328 224357
rect 459568 224345 459574 224357
rect 325322 224317 459574 224345
rect 325322 224305 325328 224317
rect 459568 224305 459574 224317
rect 459626 224305 459632 224357
rect 328240 224231 328246 224283
rect 328298 224271 328304 224283
rect 465616 224271 465622 224283
rect 328298 224243 465622 224271
rect 328298 224231 328304 224243
rect 465616 224231 465622 224243
rect 465674 224231 465680 224283
rect 331504 224157 331510 224209
rect 331562 224197 331568 224209
rect 471568 224197 471574 224209
rect 331562 224169 471574 224197
rect 331562 224157 331568 224169
rect 471568 224157 471574 224169
rect 471626 224157 471632 224209
rect 553264 224157 553270 224209
rect 553322 224197 553328 224209
rect 555376 224197 555382 224209
rect 553322 224169 555382 224197
rect 553322 224157 553328 224169
rect 555376 224157 555382 224169
rect 555434 224157 555440 224209
rect 330736 224083 330742 224135
rect 330794 224123 330800 224135
rect 467824 224123 467830 224135
rect 330794 224095 467830 224123
rect 330794 224083 330800 224095
rect 467824 224083 467830 224095
rect 467882 224083 467888 224135
rect 334480 224009 334486 224061
rect 334538 224049 334544 224061
rect 477616 224049 477622 224061
rect 334538 224021 477622 224049
rect 334538 224009 334544 224021
rect 477616 224009 477622 224021
rect 477674 224009 477680 224061
rect 337168 223935 337174 223987
rect 337226 223975 337232 223987
rect 483760 223975 483766 223987
rect 337226 223947 483766 223975
rect 337226 223935 337232 223947
rect 483760 223935 483766 223947
rect 483818 223935 483824 223987
rect 340432 223861 340438 223913
rect 340490 223901 340496 223913
rect 489712 223901 489718 223913
rect 340490 223873 489718 223901
rect 340490 223861 340496 223873
rect 489712 223861 489718 223873
rect 489770 223861 489776 223913
rect 343600 223787 343606 223839
rect 343658 223827 343664 223839
rect 497296 223827 497302 223839
rect 343658 223799 497302 223827
rect 343658 223787 343664 223799
rect 497296 223787 497302 223799
rect 497354 223787 497360 223839
rect 261904 223713 261910 223765
rect 261962 223753 261968 223765
rect 332656 223753 332662 223765
rect 261962 223725 332662 223753
rect 261962 223713 261968 223725
rect 332656 223713 332662 223725
rect 332714 223713 332720 223765
rect 346576 223713 346582 223765
rect 346634 223753 346640 223765
rect 501808 223753 501814 223765
rect 346634 223725 501814 223753
rect 346634 223713 346640 223725
rect 501808 223713 501814 223725
rect 501866 223713 501872 223765
rect 263536 223639 263542 223691
rect 263594 223679 263600 223691
rect 335728 223679 335734 223691
rect 263594 223651 335734 223679
rect 263594 223639 263600 223651
rect 335728 223639 335734 223651
rect 335786 223639 335792 223691
rect 349552 223639 349558 223691
rect 349610 223679 349616 223691
rect 507856 223679 507862 223691
rect 349610 223651 507862 223679
rect 349610 223639 349616 223651
rect 507856 223639 507862 223651
rect 507914 223639 507920 223691
rect 268048 223565 268054 223617
rect 268106 223605 268112 223617
rect 344848 223605 344854 223617
rect 268106 223577 344854 223605
rect 268106 223565 268112 223577
rect 344848 223565 344854 223577
rect 344906 223565 344912 223617
rect 348016 223565 348022 223617
rect 348074 223605 348080 223617
rect 504784 223605 504790 223617
rect 348074 223577 504790 223605
rect 348074 223565 348080 223577
rect 504784 223565 504790 223577
rect 504842 223565 504848 223617
rect 266512 223491 266518 223543
rect 266570 223531 266576 223543
rect 341776 223531 341782 223543
rect 266570 223503 341782 223531
rect 266570 223491 266576 223503
rect 341776 223491 341782 223503
rect 341834 223491 341840 223543
rect 348112 223491 348118 223543
rect 348170 223531 348176 223543
rect 506320 223531 506326 223543
rect 348170 223503 506326 223531
rect 348170 223491 348176 223503
rect 506320 223491 506326 223503
rect 506378 223491 506384 223543
rect 264592 223417 264598 223469
rect 264650 223457 264656 223469
rect 338704 223457 338710 223469
rect 264650 223429 338710 223457
rect 264650 223417 264656 223429
rect 338704 223417 338710 223429
rect 338762 223417 338768 223469
rect 351088 223417 351094 223469
rect 351146 223457 351152 223469
rect 510832 223457 510838 223469
rect 351146 223429 510838 223457
rect 351146 223417 351152 223429
rect 510832 223417 510838 223429
rect 510890 223417 510896 223469
rect 270928 223343 270934 223395
rect 270986 223383 270992 223395
rect 350800 223383 350806 223395
rect 270986 223355 350806 223383
rect 270986 223343 270992 223355
rect 350800 223343 350806 223355
rect 350858 223343 350864 223395
rect 352528 223343 352534 223395
rect 352586 223383 352592 223395
rect 513904 223383 513910 223395
rect 352586 223355 513910 223383
rect 352586 223343 352592 223355
rect 513904 223343 513910 223355
rect 513962 223343 513968 223395
rect 269392 223269 269398 223321
rect 269450 223309 269456 223321
rect 347728 223309 347734 223321
rect 269450 223281 347734 223309
rect 269450 223269 269456 223281
rect 347728 223269 347734 223281
rect 347786 223269 347792 223321
rect 351184 223269 351190 223321
rect 351242 223309 351248 223321
rect 512368 223309 512374 223321
rect 351242 223281 512374 223309
rect 351242 223269 351248 223281
rect 512368 223269 512374 223281
rect 512426 223269 512432 223321
rect 272560 223195 272566 223247
rect 272618 223235 272624 223247
rect 353872 223235 353878 223247
rect 272618 223207 353878 223235
rect 272618 223195 272624 223207
rect 353872 223195 353878 223207
rect 353930 223195 353936 223247
rect 354064 223195 354070 223247
rect 354122 223235 354128 223247
rect 516976 223235 516982 223247
rect 354122 223207 516982 223235
rect 354122 223195 354128 223207
rect 516976 223195 516982 223207
rect 517034 223195 517040 223247
rect 313360 223121 313366 223173
rect 313418 223161 313424 223173
rect 435376 223161 435382 223173
rect 313418 223133 435382 223161
rect 313418 223121 313424 223133
rect 435376 223121 435382 223133
rect 435434 223121 435440 223173
rect 310288 223047 310294 223099
rect 310346 223087 310352 223099
rect 429328 223087 429334 223099
rect 310346 223059 429334 223087
rect 310346 223047 310352 223059
rect 429328 223047 429334 223059
rect 429386 223047 429392 223099
rect 307216 222973 307222 223025
rect 307274 223013 307280 223025
rect 423280 223013 423286 223025
rect 307274 222985 423286 223013
rect 307274 222973 307280 222985
rect 423280 222973 423286 222985
rect 423338 222973 423344 223025
rect 312592 222899 312598 222951
rect 312650 222939 312656 222951
rect 431536 222939 431542 222951
rect 312650 222911 431542 222939
rect 312650 222899 312656 222911
rect 431536 222899 431542 222911
rect 431594 222899 431600 222951
rect 307984 222825 307990 222877
rect 308042 222865 308048 222877
rect 422512 222865 422518 222877
rect 308042 222837 422518 222865
rect 308042 222825 308048 222837
rect 422512 222825 422518 222837
rect 422570 222825 422576 222877
rect 304240 222751 304246 222803
rect 304298 222791 304304 222803
rect 417232 222791 417238 222803
rect 304298 222763 417238 222791
rect 304298 222751 304304 222763
rect 417232 222751 417238 222763
rect 417290 222751 417296 222803
rect 286192 222677 286198 222729
rect 286250 222717 286256 222729
rect 381040 222717 381046 222729
rect 286250 222689 381046 222717
rect 286250 222677 286256 222689
rect 381040 222677 381046 222689
rect 381098 222677 381104 222729
rect 401104 222677 401110 222729
rect 401162 222717 401168 222729
rect 511600 222717 511606 222729
rect 401162 222689 511606 222717
rect 401162 222677 401168 222689
rect 511600 222677 511606 222689
rect 511658 222677 511664 222729
rect 302800 222603 302806 222655
rect 302858 222643 302864 222655
rect 414256 222643 414262 222655
rect 302858 222615 414262 222643
rect 302858 222603 302864 222615
rect 414256 222603 414262 222615
rect 414314 222603 414320 222655
rect 301936 222529 301942 222581
rect 301994 222569 302000 222581
rect 410512 222569 410518 222581
rect 301994 222541 410518 222569
rect 301994 222529 302000 222541
rect 410512 222529 410518 222541
rect 410570 222529 410576 222581
rect 410608 222529 410614 222581
rect 410666 222569 410672 222581
rect 430096 222569 430102 222581
rect 410666 222541 430102 222569
rect 410666 222529 410672 222541
rect 430096 222529 430102 222541
rect 430154 222529 430160 222581
rect 281584 222455 281590 222507
rect 281642 222495 281648 222507
rect 371920 222495 371926 222507
rect 281642 222467 371926 222495
rect 281642 222455 281648 222467
rect 371920 222455 371926 222467
rect 371978 222455 371984 222507
rect 394864 222455 394870 222507
rect 394922 222495 394928 222507
rect 496528 222495 496534 222507
rect 394922 222467 496534 222495
rect 394922 222455 394928 222467
rect 496528 222455 496534 222467
rect 496586 222455 496592 222507
rect 283120 222381 283126 222433
rect 283178 222421 283184 222433
rect 374992 222421 374998 222433
rect 283178 222393 374998 222421
rect 283178 222381 283184 222393
rect 374992 222381 374998 222393
rect 375050 222381 375056 222433
rect 386224 222381 386230 222433
rect 386282 222421 386288 222433
rect 482896 222421 482902 222433
rect 386282 222393 482902 222421
rect 386282 222381 386288 222393
rect 482896 222381 482902 222393
rect 482954 222381 482960 222433
rect 274096 222307 274102 222359
rect 274154 222347 274160 222359
rect 356848 222347 356854 222359
rect 274154 222319 356854 222347
rect 274154 222307 274160 222319
rect 356848 222307 356854 222319
rect 356906 222307 356912 222359
rect 371632 222307 371638 222359
rect 371690 222347 371696 222359
rect 443728 222347 443734 222359
rect 371690 222319 443734 222347
rect 371690 222307 371696 222319
rect 443728 222307 443734 222319
rect 443786 222307 443792 222359
rect 149392 221863 149398 221915
rect 149450 221903 149456 221915
rect 171376 221903 171382 221915
rect 149450 221875 171382 221903
rect 149450 221863 149456 221875
rect 171376 221863 171382 221875
rect 171434 221863 171440 221915
rect 149488 221789 149494 221841
rect 149546 221829 149552 221841
rect 182896 221829 182902 221841
rect 149546 221801 182902 221829
rect 149546 221789 149552 221801
rect 182896 221789 182902 221801
rect 182954 221789 182960 221841
rect 145648 221715 145654 221767
rect 145706 221755 145712 221767
rect 184336 221755 184342 221767
rect 145706 221727 184342 221755
rect 145706 221715 145712 221727
rect 184336 221715 184342 221727
rect 184394 221715 184400 221767
rect 478096 221715 478102 221767
rect 478154 221755 478160 221767
rect 479968 221755 479974 221767
rect 478154 221727 479974 221755
rect 478154 221715 478160 221727
rect 479968 221715 479974 221727
rect 480026 221715 480032 221767
rect 512752 221715 512758 221767
rect 512810 221755 512816 221767
rect 515392 221755 515398 221767
rect 512810 221727 515398 221755
rect 512810 221715 512816 221727
rect 515392 221715 515398 221727
rect 515450 221715 515456 221767
rect 655984 219347 655990 219399
rect 656042 219387 656048 219399
rect 676240 219387 676246 219399
rect 656042 219359 676246 219387
rect 656042 219347 656048 219359
rect 676240 219347 676246 219359
rect 676298 219347 676304 219399
rect 655792 219199 655798 219251
rect 655850 219239 655856 219251
rect 676240 219239 676246 219251
rect 655850 219211 676246 219239
rect 655850 219199 655856 219211
rect 676240 219199 676246 219211
rect 676298 219199 676304 219251
rect 149392 219051 149398 219103
rect 149450 219091 149456 219103
rect 162640 219091 162646 219103
rect 149450 219063 162646 219091
rect 149450 219051 149456 219063
rect 162640 219051 162646 219063
rect 162698 219051 162704 219103
rect 655600 219051 655606 219103
rect 655658 219091 655664 219103
rect 676048 219091 676054 219103
rect 655658 219063 676054 219091
rect 655658 219051 655664 219063
rect 676048 219051 676054 219063
rect 676106 219051 676112 219103
rect 149488 218977 149494 219029
rect 149546 219017 149552 219029
rect 168400 219017 168406 219029
rect 149546 218989 168406 219017
rect 149546 218977 149552 218989
rect 168400 218977 168406 218989
rect 168458 218977 168464 219029
rect 149392 218903 149398 218955
rect 149450 218943 149456 218955
rect 180016 218943 180022 218955
rect 149450 218915 180022 218943
rect 149450 218903 149456 218915
rect 180016 218903 180022 218915
rect 180074 218903 180080 218955
rect 143056 218829 143062 218881
rect 143114 218869 143120 218881
rect 184336 218869 184342 218881
rect 143114 218841 184342 218869
rect 143114 218829 143120 218841
rect 184336 218829 184342 218841
rect 184394 218829 184400 218881
rect 147280 217719 147286 217771
rect 147338 217759 147344 217771
rect 151792 217759 151798 217771
rect 147338 217731 151798 217759
rect 147338 217719 147344 217731
rect 151792 217719 151798 217731
rect 151850 217719 151856 217771
rect 149392 216017 149398 216069
rect 149450 216057 149456 216069
rect 177232 216057 177238 216069
rect 149450 216029 177238 216057
rect 149450 216017 149456 216029
rect 177232 216017 177238 216029
rect 177290 216017 177296 216069
rect 41776 213279 41782 213331
rect 41834 213319 41840 213331
rect 45904 213319 45910 213331
rect 41834 213291 45910 213319
rect 41834 213279 41840 213291
rect 45904 213279 45910 213291
rect 45962 213279 45968 213331
rect 149488 213205 149494 213257
rect 149546 213245 149552 213257
rect 159952 213245 159958 213257
rect 149546 213217 159958 213245
rect 149546 213205 149552 213217
rect 159952 213205 159958 213217
rect 160010 213205 160016 213257
rect 674704 213205 674710 213257
rect 674762 213245 674768 213257
rect 676240 213245 676246 213257
rect 674762 213217 676246 213245
rect 674762 213205 674768 213217
rect 676240 213205 676246 213217
rect 676298 213205 676304 213257
rect 149392 213131 149398 213183
rect 149450 213171 149456 213183
rect 174352 213171 174358 213183
rect 149450 213143 174358 213171
rect 149450 213131 149456 213143
rect 174352 213131 174358 213143
rect 174410 213131 174416 213183
rect 675184 213131 675190 213183
rect 675242 213171 675248 213183
rect 676048 213171 676054 213183
rect 675242 213143 676054 213171
rect 675242 213131 675248 213143
rect 676048 213131 676054 213143
rect 676106 213131 676112 213183
rect 41584 212909 41590 212961
rect 41642 212949 41648 212961
rect 45712 212949 45718 212961
rect 41642 212921 45718 212949
rect 41642 212909 41648 212921
rect 45712 212909 45718 212921
rect 45770 212909 45776 212961
rect 146896 212761 146902 212813
rect 146954 212801 146960 212813
rect 151984 212801 151990 212813
rect 146954 212773 151990 212801
rect 146954 212761 146960 212773
rect 151984 212761 151990 212773
rect 152042 212761 152048 212813
rect 41776 212169 41782 212221
rect 41834 212209 41840 212221
rect 45616 212209 45622 212221
rect 41834 212181 45622 212209
rect 41834 212169 41840 212181
rect 45616 212169 45622 212181
rect 45674 212169 45680 212221
rect 41776 211725 41782 211777
rect 41834 211765 41840 211777
rect 43216 211765 43222 211777
rect 41834 211737 43222 211765
rect 41834 211725 41840 211737
rect 43216 211725 43222 211737
rect 43274 211725 43280 211777
rect 41584 211429 41590 211481
rect 41642 211469 41648 211481
rect 44848 211469 44854 211481
rect 41642 211441 44854 211469
rect 41642 211429 41648 211441
rect 44848 211429 44854 211441
rect 44906 211429 44912 211481
rect 147088 210985 147094 211037
rect 147146 211025 147152 211037
rect 151696 211025 151702 211037
rect 147146 210997 151702 211025
rect 147146 210985 147152 210997
rect 151696 210985 151702 210997
rect 151754 210985 151760 211037
rect 41776 210689 41782 210741
rect 41834 210729 41840 210741
rect 50512 210729 50518 210741
rect 41834 210701 50518 210729
rect 41834 210689 41840 210701
rect 50512 210689 50518 210701
rect 50570 210689 50576 210741
rect 147472 210319 147478 210371
rect 147530 210359 147536 210371
rect 151600 210359 151606 210371
rect 147530 210331 151606 210359
rect 147530 210319 147536 210331
rect 151600 210319 151606 210331
rect 151658 210319 151664 210371
rect 674800 210319 674806 210371
rect 674858 210359 674864 210371
rect 676048 210359 676054 210371
rect 674858 210331 676054 210359
rect 674858 210319 674864 210331
rect 676048 210319 676054 210331
rect 676106 210319 676112 210371
rect 674896 210245 674902 210297
rect 674954 210285 674960 210297
rect 676240 210285 676246 210297
rect 674954 210257 676246 210285
rect 674954 210245 674960 210257
rect 676240 210245 676246 210257
rect 676298 210245 676304 210297
rect 41776 210171 41782 210223
rect 41834 210211 41840 210223
rect 46192 210211 46198 210223
rect 41834 210183 46198 210211
rect 41834 210171 41840 210183
rect 46192 210171 46198 210183
rect 46250 210171 46256 210223
rect 41584 209949 41590 210001
rect 41642 209989 41648 210001
rect 50320 209989 50326 210001
rect 41642 209961 50326 209989
rect 41642 209949 41648 209961
rect 50320 209949 50326 209961
rect 50378 209949 50384 210001
rect 41584 209357 41590 209409
rect 41642 209397 41648 209409
rect 46096 209397 46102 209409
rect 41642 209369 46102 209397
rect 41642 209357 41648 209369
rect 46096 209357 46102 209369
rect 46154 209357 46160 209409
rect 147184 207877 147190 207929
rect 147242 207917 147248 207929
rect 151504 207917 151510 207929
rect 147242 207889 151510 207917
rect 147242 207877 147248 207889
rect 151504 207877 151510 207889
rect 151562 207877 151568 207929
rect 646768 207507 646774 207559
rect 646826 207547 646832 207559
rect 679888 207547 679894 207559
rect 646826 207519 679894 207547
rect 646826 207507 646832 207519
rect 679888 207507 679894 207519
rect 679946 207507 679952 207559
rect 674032 207433 674038 207485
rect 674090 207473 674096 207485
rect 675952 207473 675958 207485
rect 674090 207445 675958 207473
rect 674090 207433 674096 207445
rect 675952 207433 675958 207445
rect 676010 207433 676016 207485
rect 146896 207359 146902 207411
rect 146954 207399 146960 207411
rect 151888 207399 151894 207411
rect 146954 207371 151894 207399
rect 146954 207359 146960 207371
rect 151888 207359 151894 207371
rect 151946 207359 151952 207411
rect 674992 207359 674998 207411
rect 675050 207399 675056 207411
rect 676048 207399 676054 207411
rect 675050 207371 676054 207399
rect 675050 207359 675056 207371
rect 676048 207359 676054 207371
rect 676106 207359 676112 207411
rect 146896 206249 146902 206301
rect 146954 206289 146960 206301
rect 152080 206289 152086 206301
rect 146954 206261 152086 206289
rect 146954 206249 146960 206261
rect 152080 206249 152086 206261
rect 152138 206249 152144 206301
rect 185776 205879 185782 205931
rect 185834 205919 185840 205931
rect 186256 205919 186262 205931
rect 185834 205891 186262 205919
rect 185834 205879 185840 205891
rect 186256 205879 186262 205891
rect 186314 205879 186320 205931
rect 674608 205435 674614 205487
rect 674666 205475 674672 205487
rect 674800 205475 674806 205487
rect 674666 205447 674806 205475
rect 674666 205435 674672 205447
rect 674800 205435 674806 205447
rect 674858 205435 674864 205487
rect 149488 204473 149494 204525
rect 149546 204513 149552 204525
rect 165712 204513 165718 204525
rect 149546 204485 165718 204513
rect 149546 204473 149552 204485
rect 165712 204473 165718 204485
rect 165770 204473 165776 204525
rect 149392 204177 149398 204229
rect 149450 204217 149456 204229
rect 157072 204217 157078 204229
rect 149450 204189 157078 204217
rect 149450 204177 149456 204189
rect 157072 204177 157078 204189
rect 157130 204177 157136 204229
rect 147856 202845 147862 202897
rect 147914 202885 147920 202897
rect 154192 202885 154198 202897
rect 147914 202857 154198 202885
rect 147914 202845 147920 202857
rect 154192 202845 154198 202857
rect 154250 202845 154256 202897
rect 675088 202401 675094 202453
rect 675146 202441 675152 202453
rect 675376 202441 675382 202453
rect 675146 202413 675382 202441
rect 675146 202401 675152 202413
rect 675376 202401 675382 202413
rect 675434 202401 675440 202453
rect 41872 201661 41878 201713
rect 41930 201701 41936 201713
rect 44752 201701 44758 201713
rect 41930 201673 44758 201701
rect 41930 201661 41936 201673
rect 44752 201661 44758 201673
rect 44810 201661 44816 201713
rect 149392 201587 149398 201639
rect 149450 201627 149456 201639
rect 182992 201627 182998 201639
rect 149450 201599 182998 201627
rect 149450 201587 149456 201599
rect 182992 201587 182998 201599
rect 183050 201587 183056 201639
rect 41584 201513 41590 201565
rect 41642 201553 41648 201565
rect 44656 201553 44662 201565
rect 41642 201525 44662 201553
rect 41642 201513 41648 201525
rect 44656 201513 44662 201525
rect 44714 201513 44720 201565
rect 143056 201513 143062 201565
rect 143114 201553 143120 201565
rect 184336 201553 184342 201565
rect 143114 201525 184342 201553
rect 143114 201513 143120 201525
rect 184336 201513 184342 201525
rect 184394 201513 184400 201565
rect 674704 201365 674710 201417
rect 674762 201405 674768 201417
rect 675184 201405 675190 201417
rect 674762 201377 675190 201405
rect 674762 201365 674768 201377
rect 675184 201365 675190 201377
rect 675242 201365 675248 201417
rect 41584 200921 41590 200973
rect 41642 200961 41648 200973
rect 44560 200961 44566 200973
rect 41642 200933 44566 200961
rect 41642 200921 41648 200933
rect 44560 200921 44566 200933
rect 44618 200921 44624 200973
rect 149392 200477 149398 200529
rect 149450 200517 149456 200529
rect 160048 200517 160054 200529
rect 149450 200489 160054 200517
rect 149450 200477 149456 200489
rect 160048 200477 160054 200489
rect 160106 200477 160112 200529
rect 674992 199515 674998 199567
rect 675050 199555 675056 199567
rect 675472 199555 675478 199567
rect 675050 199527 675478 199555
rect 675050 199515 675056 199527
rect 675472 199515 675478 199527
rect 675530 199515 675536 199567
rect 147568 199293 147574 199345
rect 147626 199333 147632 199345
rect 152176 199333 152182 199345
rect 147626 199305 152182 199333
rect 147626 199293 147632 199305
rect 152176 199293 152182 199305
rect 152234 199293 152240 199345
rect 181360 198627 181366 198679
rect 181418 198667 181424 198679
rect 184336 198667 184342 198679
rect 181418 198639 184342 198667
rect 181418 198627 181424 198639
rect 184336 198627 184342 198639
rect 184394 198627 184400 198679
rect 660880 198627 660886 198679
rect 660938 198667 660944 198679
rect 675088 198667 675094 198679
rect 660938 198639 675094 198667
rect 660938 198627 660944 198639
rect 675088 198627 675094 198639
rect 675146 198627 675152 198679
rect 178288 198553 178294 198605
rect 178346 198593 178352 198605
rect 184432 198593 184438 198605
rect 178346 198565 184438 198593
rect 178346 198553 178352 198565
rect 184432 198553 184438 198565
rect 184490 198553 184496 198605
rect 674800 198553 674806 198605
rect 674858 198593 674864 198605
rect 675472 198593 675478 198605
rect 674858 198565 675478 198593
rect 674858 198553 674864 198565
rect 675472 198553 675478 198565
rect 675530 198553 675536 198605
rect 674608 198183 674614 198235
rect 674666 198223 674672 198235
rect 675376 198223 675382 198235
rect 674666 198195 675382 198223
rect 674666 198183 674672 198195
rect 675376 198183 675382 198195
rect 675434 198183 675440 198235
rect 674896 197665 674902 197717
rect 674954 197705 674960 197717
rect 675376 197705 675382 197717
rect 674954 197677 675382 197705
rect 674954 197665 674960 197677
rect 675376 197665 675382 197677
rect 675434 197665 675440 197717
rect 41776 197591 41782 197643
rect 41834 197591 41840 197643
rect 41794 197421 41822 197591
rect 41776 197369 41782 197421
rect 41834 197369 41840 197421
rect 147280 195963 147286 196015
rect 147338 196003 147344 196015
rect 171568 196003 171574 196015
rect 147338 195975 171574 196003
rect 147338 195963 147344 195975
rect 171568 195963 171574 195975
rect 171626 195963 171632 196015
rect 149392 195889 149398 195941
rect 149450 195929 149456 195941
rect 174448 195929 174454 195941
rect 149450 195901 174454 195929
rect 149450 195889 149456 195901
rect 174448 195889 174454 195901
rect 174506 195889 174512 195941
rect 149296 195815 149302 195867
rect 149354 195855 149360 195867
rect 180208 195855 180214 195867
rect 149354 195827 180214 195855
rect 149354 195815 149360 195827
rect 180208 195815 180214 195827
rect 180266 195815 180272 195867
rect 166960 195741 166966 195793
rect 167018 195781 167024 195793
rect 184528 195781 184534 195793
rect 167018 195753 184534 195781
rect 167018 195741 167024 195753
rect 184528 195741 184534 195753
rect 184586 195741 184592 195793
rect 169840 195667 169846 195719
rect 169898 195707 169904 195719
rect 184432 195707 184438 195719
rect 169898 195679 184438 195707
rect 169898 195667 169904 195679
rect 184432 195667 184438 195679
rect 184490 195667 184496 195719
rect 172720 195593 172726 195645
rect 172778 195633 172784 195645
rect 184336 195633 184342 195645
rect 172778 195605 184342 195633
rect 172778 195593 172784 195605
rect 184336 195593 184342 195605
rect 184394 195593 184400 195645
rect 674032 194335 674038 194387
rect 674090 194375 674096 194387
rect 675376 194375 675382 194387
rect 674090 194347 675382 194375
rect 674090 194335 674096 194347
rect 675376 194335 675382 194347
rect 675434 194335 675440 194387
rect 149392 193077 149398 193129
rect 149450 193117 149456 193129
rect 165808 193117 165814 193129
rect 149450 193089 165814 193117
rect 149450 193077 149456 193089
rect 165808 193077 165814 193089
rect 165866 193077 165872 193129
rect 149488 193003 149494 193055
rect 149546 193043 149552 193055
rect 168592 193043 168598 193055
rect 149546 193015 168598 193043
rect 149546 193003 149552 193015
rect 168592 193003 168598 193015
rect 168650 193003 168656 193055
rect 152368 192929 152374 192981
rect 152426 192969 152432 192981
rect 184624 192969 184630 192981
rect 152426 192941 184630 192969
rect 152426 192929 152432 192941
rect 184624 192929 184630 192941
rect 184682 192929 184688 192981
rect 155440 192855 155446 192907
rect 155498 192895 155504 192907
rect 184528 192895 184534 192907
rect 155498 192867 184534 192895
rect 155498 192855 155504 192867
rect 184528 192855 184534 192867
rect 184586 192855 184592 192907
rect 158128 192781 158134 192833
rect 158186 192821 158192 192833
rect 184336 192821 184342 192833
rect 158186 192793 184342 192821
rect 158186 192781 158192 192793
rect 184336 192781 184342 192793
rect 184394 192781 184400 192833
rect 163888 192707 163894 192759
rect 163946 192747 163952 192759
rect 184432 192747 184438 192759
rect 163946 192719 184438 192747
rect 163946 192707 163952 192719
rect 184432 192707 184438 192719
rect 184490 192707 184496 192759
rect 149392 190191 149398 190243
rect 149450 190231 149456 190243
rect 157168 190231 157174 190243
rect 149450 190203 157174 190231
rect 149450 190191 149456 190203
rect 157168 190191 157174 190203
rect 157226 190191 157232 190243
rect 149488 190117 149494 190169
rect 149546 190157 149552 190169
rect 162832 190157 162838 190169
rect 149546 190129 162838 190157
rect 149546 190117 149552 190129
rect 162832 190117 162838 190129
rect 162890 190117 162896 190169
rect 143920 190043 143926 190095
rect 143978 190083 143984 190095
rect 184528 190083 184534 190095
rect 143978 190055 184534 190083
rect 143978 190043 143984 190055
rect 184528 190043 184534 190055
rect 184586 190043 184592 190095
rect 149680 189969 149686 190021
rect 149738 190009 149744 190021
rect 184336 190009 184342 190021
rect 149738 189981 184342 190009
rect 149738 189969 149744 189981
rect 184336 189969 184342 189981
rect 184394 189969 184400 190021
rect 171472 189895 171478 189947
rect 171530 189935 171536 189947
rect 184432 189935 184438 189947
rect 171530 189907 184438 189935
rect 171530 189895 171536 189907
rect 184432 189895 184438 189907
rect 184490 189895 184496 189947
rect 174256 189821 174262 189873
rect 174314 189861 174320 189873
rect 184336 189861 184342 189873
rect 174314 189833 184342 189861
rect 174314 189821 174320 189833
rect 184336 189821 184342 189833
rect 184394 189821 184400 189873
rect 147664 189525 147670 189577
rect 147722 189565 147728 189577
rect 154288 189565 154294 189577
rect 147722 189537 154294 189565
rect 147722 189525 147728 189537
rect 154288 189525 154294 189537
rect 154346 189525 154352 189577
rect 145552 187157 145558 187209
rect 145610 187197 145616 187209
rect 184336 187197 184342 187209
rect 145610 187169 184342 187197
rect 145610 187157 145616 187169
rect 184336 187157 184342 187169
rect 184394 187157 184400 187209
rect 162736 187083 162742 187135
rect 162794 187123 162800 187135
rect 184528 187123 184534 187135
rect 162794 187095 184534 187123
rect 162794 187083 162800 187095
rect 184528 187083 184534 187095
rect 184586 187083 184592 187135
rect 168496 187009 168502 187061
rect 168554 187049 168560 187061
rect 184432 187049 184438 187061
rect 168554 187021 184438 187049
rect 168554 187009 168560 187021
rect 184432 187009 184438 187021
rect 184490 187009 184496 187061
rect 180112 186935 180118 186987
rect 180170 186975 180176 186987
rect 185392 186975 185398 186987
rect 180170 186947 185398 186975
rect 180170 186935 180176 186947
rect 185392 186935 185398 186947
rect 185450 186935 185456 186987
rect 156976 184271 156982 184323
rect 157034 184311 157040 184323
rect 184432 184311 184438 184323
rect 157034 184283 184438 184311
rect 157034 184271 157040 184283
rect 184432 184271 184438 184283
rect 184490 184271 184496 184323
rect 165616 184197 165622 184249
rect 165674 184237 165680 184249
rect 184336 184237 184342 184249
rect 165674 184209 184342 184237
rect 165674 184197 165680 184209
rect 184336 184197 184342 184209
rect 184394 184197 184400 184249
rect 179920 184123 179926 184175
rect 179978 184163 179984 184175
rect 184528 184163 184534 184175
rect 179978 184135 184534 184163
rect 179978 184123 179984 184135
rect 184528 184123 184534 184135
rect 184586 184123 184592 184175
rect 645136 183087 645142 183139
rect 645194 183127 645200 183139
rect 649360 183127 649366 183139
rect 645194 183099 649366 183127
rect 645194 183087 645200 183099
rect 649360 183087 649366 183099
rect 649418 183087 649424 183139
rect 149392 182939 149398 182991
rect 149450 182979 149456 182991
rect 185968 182979 185974 182991
rect 149450 182951 185974 182979
rect 149450 182939 149456 182951
rect 185968 182939 185974 182951
rect 186026 182939 186032 182991
rect 149296 182865 149302 182917
rect 149354 182905 149360 182917
rect 186160 182905 186166 182917
rect 149354 182877 186166 182905
rect 149354 182865 149360 182877
rect 186160 182865 186166 182877
rect 186218 182865 186224 182917
rect 42160 182347 42166 182399
rect 42218 182387 42224 182399
rect 45328 182387 45334 182399
rect 42218 182359 45334 182387
rect 42218 182347 42224 182359
rect 45328 182347 45334 182359
rect 45386 182347 45392 182399
rect 149488 181533 149494 181585
rect 149546 181573 149552 181585
rect 177328 181573 177334 181585
rect 149546 181545 177334 181573
rect 149546 181533 149552 181545
rect 177328 181533 177334 181545
rect 177386 181533 177392 181585
rect 149392 181459 149398 181511
rect 149450 181499 149456 181511
rect 183088 181499 183094 181511
rect 149450 181471 183094 181499
rect 149450 181459 149456 181471
rect 183088 181459 183094 181471
rect 183146 181459 183152 181511
rect 154000 181385 154006 181437
rect 154058 181425 154064 181437
rect 184624 181425 184630 181437
rect 154058 181397 184630 181425
rect 154058 181385 154064 181397
rect 184624 181385 184630 181397
rect 184682 181385 184688 181437
rect 156880 181311 156886 181363
rect 156938 181351 156944 181363
rect 184528 181351 184534 181363
rect 156938 181323 184534 181351
rect 156938 181311 156944 181323
rect 184528 181311 184534 181323
rect 184586 181311 184592 181363
rect 165520 181237 165526 181289
rect 165578 181277 165584 181289
rect 184432 181277 184438 181289
rect 165578 181249 184438 181277
rect 165578 181237 165584 181249
rect 184432 181237 184438 181249
rect 184490 181237 184496 181289
rect 171280 181163 171286 181215
rect 171338 181203 171344 181215
rect 184336 181203 184342 181215
rect 171338 181175 184342 181203
rect 171338 181163 171344 181175
rect 184336 181163 184342 181175
rect 184394 181163 184400 181215
rect 149584 179979 149590 180031
rect 149642 180019 149648 180031
rect 185392 180019 185398 180031
rect 149642 179991 185398 180019
rect 149642 179979 149648 179991
rect 185392 179979 185398 179991
rect 185450 179979 185456 180031
rect 645136 179387 645142 179439
rect 645194 179427 645200 179439
rect 649456 179427 649462 179439
rect 645194 179399 649462 179427
rect 645194 179387 645200 179399
rect 649456 179387 649462 179399
rect 649514 179387 649520 179439
rect 149488 178721 149494 178773
rect 149546 178761 149552 178773
rect 162736 178761 162742 178773
rect 149546 178733 162742 178761
rect 149546 178721 149552 178733
rect 162736 178721 162742 178733
rect 162794 178721 162800 178773
rect 149392 178647 149398 178699
rect 149450 178687 149456 178699
rect 168496 178687 168502 178699
rect 149450 178659 168502 178687
rect 149450 178647 149456 178659
rect 168496 178647 168502 178659
rect 168554 178647 168560 178699
rect 149296 178573 149302 178625
rect 149354 178613 149360 178625
rect 171472 178613 171478 178625
rect 149354 178585 171478 178613
rect 149354 178573 149360 178585
rect 171472 178573 171478 178585
rect 171530 178573 171536 178625
rect 159760 178499 159766 178551
rect 159818 178539 159824 178551
rect 184336 178539 184342 178551
rect 159818 178511 184342 178539
rect 159818 178499 159824 178511
rect 184336 178499 184342 178511
rect 184394 178499 184400 178551
rect 182800 178425 182806 178477
rect 182858 178465 182864 178477
rect 184528 178465 184534 178477
rect 182858 178437 184534 178465
rect 182858 178425 182864 178437
rect 184528 178425 184534 178437
rect 184586 178425 184592 178477
rect 177040 178351 177046 178403
rect 177098 178391 177104 178403
rect 184432 178391 184438 178403
rect 177098 178363 184438 178391
rect 177098 178351 177104 178363
rect 184432 178351 184438 178363
rect 184490 178351 184496 178403
rect 149392 175761 149398 175813
rect 149450 175801 149456 175813
rect 156880 175801 156886 175813
rect 149450 175773 156886 175801
rect 149450 175761 149456 175773
rect 156880 175761 156886 175773
rect 156938 175761 156944 175813
rect 149488 175687 149494 175739
rect 149546 175727 149552 175739
rect 165520 175727 165526 175739
rect 149546 175699 165526 175727
rect 149546 175687 149552 175699
rect 165520 175687 165526 175699
rect 165578 175687 165584 175739
rect 145456 175613 145462 175665
rect 145514 175653 145520 175665
rect 184432 175653 184438 175665
rect 145514 175625 184438 175653
rect 145514 175613 145520 175625
rect 184432 175613 184438 175625
rect 184490 175613 184496 175665
rect 145360 175539 145366 175591
rect 145418 175579 145424 175591
rect 184336 175579 184342 175591
rect 145418 175551 184342 175579
rect 145418 175539 145424 175551
rect 184336 175539 184342 175551
rect 184394 175539 184400 175591
rect 645136 174873 645142 174925
rect 645194 174913 645200 174925
rect 649552 174913 649558 174925
rect 645194 174885 649558 174913
rect 645194 174873 645200 174885
rect 649552 174873 649558 174885
rect 649610 174873 649616 174925
rect 147760 174355 147766 174407
rect 147818 174395 147824 174407
rect 154000 174395 154006 174407
rect 147818 174367 154006 174395
rect 147818 174355 147824 174367
rect 154000 174355 154006 174367
rect 154058 174355 154064 174407
rect 149200 174207 149206 174259
rect 149258 174247 149264 174259
rect 186064 174247 186070 174259
rect 149258 174219 186070 174247
rect 149258 174207 149264 174219
rect 186064 174207 186070 174219
rect 186122 174207 186128 174259
rect 655696 173171 655702 173223
rect 655754 173211 655760 173223
rect 676240 173211 676246 173223
rect 655754 173183 676246 173211
rect 655754 173171 655760 173183
rect 676240 173171 676246 173183
rect 676298 173171 676304 173223
rect 655504 173023 655510 173075
rect 655562 173063 655568 173075
rect 676144 173063 676150 173075
rect 655562 173035 676150 173063
rect 655562 173023 655568 173035
rect 676144 173023 676150 173035
rect 676202 173023 676208 173075
rect 655408 172801 655414 172853
rect 655466 172841 655472 172853
rect 676048 172841 676054 172853
rect 655466 172813 676054 172841
rect 655466 172801 655472 172813
rect 676048 172801 676054 172813
rect 676106 172801 676112 172853
rect 148720 172727 148726 172779
rect 148778 172767 148784 172779
rect 184528 172767 184534 172779
rect 148778 172739 184534 172767
rect 148778 172727 148784 172739
rect 184528 172727 184534 172739
rect 184586 172727 184592 172779
rect 148336 172653 148342 172705
rect 148394 172693 148400 172705
rect 184336 172693 184342 172705
rect 148394 172665 184342 172693
rect 148394 172653 148400 172665
rect 184336 172653 184342 172665
rect 184394 172653 184400 172705
rect 148912 172579 148918 172631
rect 148970 172619 148976 172631
rect 184624 172619 184630 172631
rect 148970 172591 184630 172619
rect 148970 172579 148976 172591
rect 184624 172579 184630 172591
rect 184682 172579 184688 172631
rect 148528 172505 148534 172557
rect 148586 172545 148592 172557
rect 184432 172545 184438 172557
rect 148586 172517 184438 172545
rect 148586 172505 148592 172517
rect 184432 172505 184438 172517
rect 184490 172505 184496 172557
rect 645136 171025 645142 171077
rect 645194 171065 645200 171077
rect 649648 171065 649654 171077
rect 645194 171037 649654 171065
rect 645194 171025 645200 171037
rect 649648 171025 649654 171037
rect 649706 171025 649712 171077
rect 672592 169915 672598 169967
rect 672650 169955 672656 169967
rect 673840 169955 673846 169967
rect 672650 169927 673846 169955
rect 672650 169915 672656 169927
rect 673840 169915 673846 169927
rect 673898 169955 673904 169967
rect 676048 169955 676054 169967
rect 673898 169927 676054 169955
rect 673898 169915 673904 169927
rect 676048 169915 676054 169927
rect 676106 169915 676112 169967
rect 148432 169841 148438 169893
rect 148490 169881 148496 169893
rect 184528 169881 184534 169893
rect 148490 169853 184534 169881
rect 148490 169841 148496 169853
rect 184528 169841 184534 169853
rect 184586 169841 184592 169893
rect 148624 169767 148630 169819
rect 148682 169807 148688 169819
rect 184624 169807 184630 169819
rect 148682 169779 184630 169807
rect 148682 169767 148688 169779
rect 184624 169767 184630 169779
rect 184682 169767 184688 169819
rect 148240 169693 148246 169745
rect 148298 169733 148304 169745
rect 184336 169733 184342 169745
rect 148298 169705 184342 169733
rect 148298 169693 148304 169705
rect 184336 169693 184342 169705
rect 184394 169693 184400 169745
rect 151216 169619 151222 169671
rect 151274 169659 151280 169671
rect 184432 169659 184438 169671
rect 151274 169631 184438 169659
rect 151274 169619 151280 169631
rect 184432 169619 184438 169631
rect 184490 169619 184496 169671
rect 673456 169027 673462 169079
rect 673514 169067 673520 169079
rect 676048 169067 676054 169079
rect 673514 169039 676054 169067
rect 673514 169027 673520 169039
rect 676048 169027 676054 169039
rect 676106 169027 676112 169079
rect 645136 168213 645142 168265
rect 645194 168253 645200 168265
rect 649840 168253 649846 168265
rect 645194 168225 649846 168253
rect 645194 168213 645200 168225
rect 649840 168213 649846 168225
rect 649898 168213 649904 168265
rect 149008 166955 149014 167007
rect 149066 166995 149072 167007
rect 184528 166995 184534 167007
rect 149066 166967 184534 166995
rect 149066 166955 149072 166967
rect 184528 166955 184534 166967
rect 184586 166955 184592 167007
rect 148816 166881 148822 166933
rect 148874 166921 148880 166933
rect 184336 166921 184342 166933
rect 148874 166893 184342 166921
rect 148874 166881 148880 166893
rect 184336 166881 184342 166893
rect 184394 166881 184400 166933
rect 149392 166807 149398 166859
rect 149450 166847 149456 166859
rect 184432 166847 184438 166859
rect 149450 166819 184438 166847
rect 149450 166807 149456 166819
rect 184432 166807 184438 166819
rect 184490 166807 184496 166859
rect 151408 164069 151414 164121
rect 151466 164109 151472 164121
rect 184528 164109 184534 164121
rect 151466 164081 184534 164109
rect 151466 164069 151472 164081
rect 184528 164069 184534 164081
rect 184586 164069 184592 164121
rect 154096 163995 154102 164047
rect 154154 164035 154160 164047
rect 184336 164035 184342 164047
rect 154154 164007 184342 164035
rect 154154 163995 154160 164007
rect 184336 163995 184342 164007
rect 184394 163995 184400 164047
rect 174160 163921 174166 163973
rect 174218 163961 174224 163973
rect 184432 163961 184438 163973
rect 174218 163933 184438 163961
rect 174218 163921 174224 163933
rect 184432 163921 184438 163933
rect 184490 163921 184496 163973
rect 177136 163847 177142 163899
rect 177194 163887 177200 163899
rect 184336 163887 184342 163899
rect 177194 163859 184342 163887
rect 177194 163847 177200 163859
rect 184336 163847 184342 163859
rect 184394 163847 184400 163899
rect 645136 163329 645142 163381
rect 645194 163369 645200 163381
rect 649936 163369 649942 163381
rect 645194 163341 649942 163369
rect 645194 163329 645200 163341
rect 649936 163329 649942 163341
rect 649994 163329 650000 163381
rect 676240 161593 676246 161605
rect 659506 161565 676246 161593
rect 646864 161479 646870 161531
rect 646922 161519 646928 161531
rect 659506 161519 659534 161565
rect 676240 161553 676246 161565
rect 676298 161553 676304 161605
rect 646922 161491 659534 161519
rect 646922 161479 646928 161491
rect 647056 161405 647062 161457
rect 647114 161445 647120 161457
rect 676240 161445 676246 161457
rect 647114 161417 676246 161445
rect 647114 161405 647120 161417
rect 676240 161405 676246 161417
rect 676298 161405 676304 161457
rect 646960 161331 646966 161383
rect 647018 161371 647024 161383
rect 676144 161371 676150 161383
rect 647018 161343 676150 161371
rect 647018 161331 647024 161343
rect 676144 161331 676150 161343
rect 676202 161331 676208 161383
rect 674128 161257 674134 161309
rect 674186 161297 674192 161309
rect 676048 161297 676054 161309
rect 674186 161269 676054 161297
rect 674186 161257 674192 161269
rect 676048 161257 676054 161269
rect 676106 161257 676112 161309
rect 182896 161183 182902 161235
rect 182954 161223 182960 161235
rect 184624 161223 184630 161235
rect 182954 161195 184630 161223
rect 182954 161183 182960 161195
rect 184624 161183 184630 161195
rect 184682 161183 184688 161235
rect 159856 161109 159862 161161
rect 159914 161149 159920 161161
rect 184432 161149 184438 161161
rect 159914 161121 184438 161149
rect 159914 161109 159920 161121
rect 184432 161109 184438 161121
rect 184490 161109 184496 161161
rect 171376 161035 171382 161087
rect 171434 161075 171440 161087
rect 184528 161075 184534 161087
rect 171434 161047 184534 161075
rect 171434 161035 171440 161047
rect 184528 161035 184534 161047
rect 184586 161035 184592 161087
rect 151312 160961 151318 161013
rect 151370 161001 151376 161013
rect 184336 161001 184342 161013
rect 151370 160973 184342 161001
rect 151370 160961 151376 160973
rect 184336 160961 184342 160973
rect 184394 160961 184400 161013
rect 645136 159703 645142 159755
rect 645194 159743 645200 159755
rect 650032 159743 650038 159755
rect 645194 159715 650038 159743
rect 645194 159703 645200 159715
rect 650032 159703 650038 159715
rect 650090 159703 650096 159755
rect 147088 158445 147094 158497
rect 147146 158485 147152 158497
rect 151408 158485 151414 158497
rect 147146 158457 151414 158485
rect 147146 158445 147152 158457
rect 151408 158445 151414 158457
rect 151466 158445 151472 158497
rect 151792 158371 151798 158423
rect 151850 158411 151856 158423
rect 184528 158411 184534 158423
rect 151850 158383 184534 158411
rect 151850 158371 151856 158383
rect 184528 158371 184534 158383
rect 184586 158371 184592 158423
rect 162640 158297 162646 158349
rect 162698 158337 162704 158349
rect 184432 158337 184438 158349
rect 162698 158309 184438 158337
rect 162698 158297 162704 158309
rect 184432 158297 184438 158309
rect 184490 158297 184496 158349
rect 168400 158223 168406 158275
rect 168458 158263 168464 158275
rect 184336 158263 184342 158275
rect 168458 158235 184342 158263
rect 168458 158223 168464 158235
rect 184336 158223 184342 158235
rect 184394 158223 184400 158275
rect 180016 158149 180022 158201
rect 180074 158189 180080 158201
rect 184624 158189 184630 158201
rect 180074 158161 184630 158189
rect 180074 158149 180080 158161
rect 184624 158149 184630 158161
rect 184682 158149 184688 158201
rect 149392 157631 149398 157683
rect 149450 157671 149456 157683
rect 159760 157671 159766 157683
rect 149450 157643 159766 157671
rect 149450 157631 149456 157643
rect 159760 157631 159766 157643
rect 159818 157631 159824 157683
rect 147088 156151 147094 156203
rect 147146 156191 147152 156203
rect 151216 156191 151222 156203
rect 147146 156163 151222 156191
rect 147146 156151 147152 156163
rect 151216 156151 151222 156163
rect 151274 156151 151280 156203
rect 645136 156003 645142 156055
rect 645194 156043 645200 156055
rect 650128 156043 650134 156055
rect 645194 156015 650134 156043
rect 645194 156003 645200 156015
rect 650128 156003 650134 156015
rect 650186 156003 650192 156055
rect 149392 155707 149398 155759
rect 149450 155747 149456 155759
rect 182800 155747 182806 155759
rect 149450 155719 182806 155747
rect 149450 155707 149456 155719
rect 182800 155707 182806 155719
rect 182858 155707 182864 155759
rect 151984 155485 151990 155537
rect 152042 155525 152048 155537
rect 184624 155525 184630 155537
rect 152042 155497 184630 155525
rect 152042 155485 152048 155497
rect 184624 155485 184630 155497
rect 184682 155485 184688 155537
rect 658000 155485 658006 155537
rect 658058 155525 658064 155537
rect 675088 155525 675094 155537
rect 658058 155497 675094 155525
rect 658058 155485 658064 155497
rect 675088 155485 675094 155497
rect 675146 155485 675152 155537
rect 159952 155411 159958 155463
rect 160010 155451 160016 155463
rect 184336 155451 184342 155463
rect 160010 155423 184342 155451
rect 160010 155411 160016 155423
rect 184336 155411 184342 155423
rect 184394 155411 184400 155463
rect 174352 155337 174358 155389
rect 174410 155377 174416 155389
rect 184432 155377 184438 155389
rect 174410 155349 184438 155377
rect 174410 155337 174416 155349
rect 184432 155337 184438 155349
rect 184490 155337 184496 155389
rect 177232 155263 177238 155315
rect 177290 155303 177296 155315
rect 184528 155303 184534 155315
rect 177290 155275 184534 155303
rect 177290 155263 177296 155275
rect 184528 155263 184534 155275
rect 184586 155263 184592 155315
rect 674128 153339 674134 153391
rect 674186 153379 674192 153391
rect 675376 153379 675382 153391
rect 674186 153351 675382 153379
rect 674186 153339 674192 153351
rect 675376 153339 675382 153351
rect 675434 153339 675440 153391
rect 149488 152747 149494 152799
rect 149546 152787 149552 152799
rect 172816 152787 172822 152799
rect 149546 152759 172822 152787
rect 149546 152747 149552 152759
rect 172816 152747 172822 152759
rect 172874 152747 172880 152799
rect 149392 152673 149398 152725
rect 149450 152713 149456 152725
rect 179920 152713 179926 152725
rect 149450 152685 179926 152713
rect 149450 152673 149456 152685
rect 179920 152673 179926 152685
rect 179978 152673 179984 152725
rect 151888 152599 151894 152651
rect 151946 152639 151952 152651
rect 184528 152639 184534 152651
rect 151946 152611 184534 152639
rect 151946 152599 151952 152611
rect 184528 152599 184534 152611
rect 184586 152599 184592 152651
rect 151600 152525 151606 152577
rect 151658 152565 151664 152577
rect 184432 152565 184438 152577
rect 151658 152537 184438 152565
rect 151658 152525 151664 152537
rect 184432 152525 184438 152537
rect 184490 152525 184496 152577
rect 645136 152525 645142 152577
rect 645194 152565 645200 152577
rect 650224 152565 650230 152577
rect 645194 152537 650230 152565
rect 645194 152525 645200 152537
rect 650224 152525 650230 152537
rect 650282 152525 650288 152577
rect 151696 152451 151702 152503
rect 151754 152491 151760 152503
rect 184336 152491 184342 152503
rect 151754 152463 184342 152491
rect 151754 152451 151760 152463
rect 184336 152451 184342 152463
rect 184394 152451 184400 152503
rect 149392 149935 149398 149987
rect 149450 149975 149456 149987
rect 174256 149975 174262 149987
rect 149450 149947 174262 149975
rect 149450 149935 149456 149947
rect 174256 149935 174262 149947
rect 174314 149935 174320 149987
rect 149488 149861 149494 149913
rect 149546 149901 149552 149913
rect 177040 149901 177046 149913
rect 149546 149873 177046 149901
rect 149546 149861 149552 149873
rect 177040 149861 177046 149873
rect 177098 149861 177104 149913
rect 149680 149787 149686 149839
rect 149738 149827 149744 149839
rect 180016 149827 180022 149839
rect 149738 149799 180022 149827
rect 149738 149787 149744 149799
rect 180016 149787 180022 149799
rect 180074 149787 180080 149839
rect 151504 149713 151510 149765
rect 151562 149753 151568 149765
rect 184336 149753 184342 149765
rect 151562 149725 184342 149753
rect 151562 149713 151568 149725
rect 184336 149713 184342 149725
rect 184394 149713 184400 149765
rect 152080 149639 152086 149691
rect 152138 149679 152144 149691
rect 184432 149679 184438 149691
rect 152138 149651 184438 149679
rect 152138 149639 152144 149651
rect 184432 149639 184438 149651
rect 184490 149639 184496 149691
rect 157072 149565 157078 149617
rect 157130 149605 157136 149617
rect 184528 149605 184534 149617
rect 157130 149577 184534 149605
rect 157130 149565 157136 149577
rect 184528 149565 184534 149577
rect 184586 149565 184592 149617
rect 165712 149491 165718 149543
rect 165770 149531 165776 149543
rect 184336 149531 184342 149543
rect 165770 149503 184342 149531
rect 165770 149491 165776 149503
rect 184336 149491 184342 149503
rect 184394 149491 184400 149543
rect 675184 149121 675190 149173
rect 675242 149161 675248 149173
rect 675376 149161 675382 149173
rect 675242 149133 675382 149161
rect 675242 149121 675248 149133
rect 675376 149121 675382 149133
rect 675434 149121 675440 149173
rect 645136 148159 645142 148211
rect 645194 148199 645200 148211
rect 650320 148199 650326 148211
rect 645194 148171 650326 148199
rect 645194 148159 645200 148171
rect 650320 148159 650326 148171
rect 650378 148159 650384 148211
rect 149008 147863 149014 147915
rect 149066 147903 149072 147915
rect 149200 147903 149206 147915
rect 149066 147875 149206 147903
rect 149066 147863 149072 147875
rect 149200 147863 149206 147875
rect 149258 147863 149264 147915
rect 149200 147419 149206 147471
rect 149258 147459 149264 147471
rect 149392 147459 149398 147471
rect 149258 147431 149398 147459
rect 149258 147419 149264 147431
rect 149392 147419 149398 147431
rect 149450 147419 149456 147471
rect 149392 146975 149398 147027
rect 149450 147015 149456 147027
rect 168400 147015 168406 147027
rect 149450 146987 168406 147015
rect 149450 146975 149456 146987
rect 168400 146975 168406 146987
rect 168458 146975 168464 147027
rect 149488 146901 149494 146953
rect 149546 146941 149552 146953
rect 171376 146941 171382 146953
rect 149546 146913 171382 146941
rect 149546 146901 149552 146913
rect 171376 146901 171382 146913
rect 171434 146901 171440 146953
rect 182992 146827 182998 146879
rect 183050 146867 183056 146879
rect 186736 146867 186742 146879
rect 183050 146839 186742 146867
rect 183050 146827 183056 146839
rect 186736 146827 186742 146839
rect 186794 146827 186800 146879
rect 154192 146753 154198 146805
rect 154250 146793 154256 146805
rect 184336 146793 184342 146805
rect 154250 146765 184342 146793
rect 154250 146753 154256 146765
rect 184336 146753 184342 146765
rect 184394 146753 184400 146805
rect 160048 146679 160054 146731
rect 160106 146719 160112 146731
rect 184432 146719 184438 146731
rect 160106 146691 184438 146719
rect 160106 146679 160112 146691
rect 184432 146679 184438 146691
rect 184490 146679 184496 146731
rect 152176 146605 152182 146657
rect 152234 146645 152240 146657
rect 184528 146645 184534 146657
rect 152234 146617 184534 146645
rect 152234 146605 152240 146617
rect 184528 146605 184534 146617
rect 184586 146605 184592 146657
rect 673456 146087 673462 146139
rect 673514 146127 673520 146139
rect 675376 146127 675382 146139
rect 673514 146099 675382 146127
rect 673514 146087 673520 146099
rect 675376 146087 675382 146099
rect 675434 146087 675440 146139
rect 149392 144089 149398 144141
rect 149450 144129 149456 144141
rect 162928 144129 162934 144141
rect 149450 144101 162934 144129
rect 149450 144089 149456 144101
rect 162928 144089 162934 144101
rect 162986 144089 162992 144141
rect 149488 144015 149494 144067
rect 149546 144055 149552 144067
rect 165712 144055 165718 144067
rect 149546 144027 165718 144055
rect 149546 144015 149552 144027
rect 165712 144015 165718 144027
rect 165770 144015 165776 144067
rect 168592 143941 168598 143993
rect 168650 143981 168656 143993
rect 184528 143981 184534 143993
rect 168650 143953 184534 143981
rect 168650 143941 168656 143953
rect 184528 143941 184534 143953
rect 184586 143941 184592 143993
rect 171568 143867 171574 143919
rect 171626 143907 171632 143919
rect 184432 143907 184438 143919
rect 171626 143879 184438 143907
rect 171626 143867 171632 143879
rect 184432 143867 184438 143879
rect 184490 143867 184496 143919
rect 174448 143793 174454 143845
rect 174506 143833 174512 143845
rect 184336 143833 184342 143845
rect 174506 143805 184342 143833
rect 174506 143793 174512 143805
rect 184336 143793 184342 143805
rect 184394 143793 184400 143845
rect 180208 143719 180214 143771
rect 180266 143759 180272 143771
rect 185392 143759 185398 143771
rect 180266 143731 185398 143759
rect 180266 143719 180272 143731
rect 185392 143719 185398 143731
rect 185450 143719 185456 143771
rect 149488 142313 149494 142365
rect 149546 142353 149552 142365
rect 159856 142353 159862 142365
rect 149546 142325 159862 142353
rect 149546 142313 149552 142325
rect 159856 142313 159862 142325
rect 159914 142313 159920 142365
rect 149392 141795 149398 141847
rect 149450 141835 149456 141847
rect 156976 141835 156982 141847
rect 149450 141807 156982 141835
rect 149450 141795 149456 141807
rect 156976 141795 156982 141807
rect 157034 141795 157040 141847
rect 147088 141203 147094 141255
rect 147146 141243 147152 141255
rect 154096 141243 154102 141255
rect 147146 141215 154102 141243
rect 147146 141203 147152 141215
rect 154096 141203 154102 141215
rect 154154 141203 154160 141255
rect 146896 141055 146902 141107
rect 146954 141095 146960 141107
rect 151120 141095 151126 141107
rect 146954 141067 151126 141095
rect 146954 141055 146960 141067
rect 151120 141055 151126 141067
rect 151178 141055 151184 141107
rect 154288 141055 154294 141107
rect 154346 141095 154352 141107
rect 184624 141095 184630 141107
rect 154346 141067 184630 141095
rect 154346 141055 154352 141067
rect 184624 141055 184630 141067
rect 184682 141055 184688 141107
rect 157168 140981 157174 141033
rect 157226 141021 157232 141033
rect 184528 141021 184534 141033
rect 157226 140993 184534 141021
rect 157226 140981 157232 140993
rect 184528 140981 184534 140993
rect 184586 140981 184592 141033
rect 162832 140907 162838 140959
rect 162890 140947 162896 140959
rect 184432 140947 184438 140959
rect 162890 140919 184438 140947
rect 162890 140907 162896 140919
rect 184432 140907 184438 140919
rect 184490 140907 184496 140959
rect 165808 140833 165814 140885
rect 165866 140873 165872 140885
rect 184336 140873 184342 140885
rect 165866 140845 184342 140873
rect 165866 140833 165872 140845
rect 184336 140833 184342 140845
rect 184394 140833 184400 140885
rect 149392 138243 149398 138295
rect 149450 138283 149456 138295
rect 162640 138283 162646 138295
rect 149450 138255 162646 138283
rect 149450 138243 149456 138255
rect 162640 138243 162646 138255
rect 162698 138243 162704 138295
rect 172816 136763 172822 136815
rect 172874 136803 172880 136815
rect 185680 136803 185686 136815
rect 172874 136775 185686 136803
rect 172874 136763 172880 136775
rect 185680 136763 185686 136775
rect 185738 136763 185744 136815
rect 149392 135431 149398 135483
rect 149450 135471 149456 135483
rect 174160 135471 174166 135483
rect 149450 135443 174166 135471
rect 149450 135431 149456 135443
rect 174160 135431 174166 135443
rect 174218 135431 174224 135483
rect 149680 135357 149686 135409
rect 149738 135397 149744 135409
rect 182896 135397 182902 135409
rect 149738 135369 182902 135397
rect 149738 135357 149744 135369
rect 182896 135357 182902 135369
rect 182954 135357 182960 135409
rect 162736 135283 162742 135335
rect 162794 135323 162800 135335
rect 184336 135323 184342 135335
rect 162794 135295 184342 135323
rect 162794 135283 162800 135295
rect 184336 135283 184342 135295
rect 184394 135283 184400 135335
rect 183088 134913 183094 134965
rect 183146 134953 183152 134965
rect 184528 134953 184534 134965
rect 183146 134925 184534 134953
rect 183146 134913 183152 134925
rect 184528 134913 184534 134925
rect 184586 134913 184592 134965
rect 177328 134839 177334 134891
rect 177386 134879 177392 134891
rect 184432 134879 184438 134891
rect 177386 134851 184438 134879
rect 177386 134839 177392 134851
rect 184432 134839 184438 134851
rect 184490 134839 184496 134891
rect 148816 133951 148822 134003
rect 148874 133991 148880 134003
rect 149584 133991 149590 134003
rect 148874 133963 149590 133991
rect 148874 133951 148880 133963
rect 149584 133951 149590 133963
rect 149642 133951 149648 134003
rect 148912 132915 148918 132967
rect 148970 132955 148976 132967
rect 149680 132955 149686 132967
rect 148970 132927 149686 132955
rect 148970 132915 148976 132927
rect 149680 132915 149686 132927
rect 149738 132915 149744 132967
rect 149392 132471 149398 132523
rect 149450 132511 149456 132523
rect 171280 132511 171286 132523
rect 149450 132483 171286 132511
rect 149450 132471 149456 132483
rect 171280 132471 171286 132483
rect 171338 132471 171344 132523
rect 156880 132397 156886 132449
rect 156938 132437 156944 132449
rect 184624 132437 184630 132449
rect 156938 132409 184630 132437
rect 156938 132397 156944 132409
rect 184624 132397 184630 132409
rect 184682 132397 184688 132449
rect 165520 132323 165526 132375
rect 165578 132363 165584 132375
rect 184528 132363 184534 132375
rect 165578 132335 184534 132363
rect 165578 132323 165584 132335
rect 184528 132323 184534 132335
rect 184586 132323 184592 132375
rect 168496 132249 168502 132301
rect 168554 132289 168560 132301
rect 184432 132289 184438 132301
rect 168554 132261 184438 132289
rect 168554 132249 168560 132261
rect 184432 132249 184438 132261
rect 184490 132249 184496 132301
rect 171472 132175 171478 132227
rect 171530 132215 171536 132227
rect 184336 132215 184342 132227
rect 171530 132187 184342 132215
rect 171530 132175 171536 132187
rect 184336 132175 184342 132187
rect 184394 132175 184400 132227
rect 149392 129659 149398 129711
rect 149450 129699 149456 129711
rect 165616 129699 165622 129711
rect 149450 129671 165622 129699
rect 149450 129659 149456 129671
rect 165616 129659 165622 129671
rect 165674 129659 165680 129711
rect 149296 129585 149302 129637
rect 149354 129625 149360 129637
rect 177232 129625 177238 129637
rect 149354 129597 177238 129625
rect 149354 129585 149360 129597
rect 177232 129585 177238 129597
rect 177290 129585 177296 129637
rect 655312 129585 655318 129637
rect 655370 129625 655376 129637
rect 676240 129625 676246 129637
rect 655370 129597 676246 129625
rect 655370 129585 655376 129597
rect 676240 129585 676246 129597
rect 676298 129585 676304 129637
rect 149200 129511 149206 129563
rect 149258 129551 149264 129563
rect 184432 129551 184438 129563
rect 149258 129523 184438 129551
rect 149258 129511 149264 129523
rect 184432 129511 184438 129523
rect 184490 129511 184496 129563
rect 149488 129437 149494 129489
rect 149546 129477 149552 129489
rect 184528 129477 184534 129489
rect 149546 129449 184534 129477
rect 149546 129437 149552 129449
rect 184528 129437 184534 129449
rect 184586 129437 184592 129489
rect 149104 129363 149110 129415
rect 149162 129403 149168 129415
rect 184624 129403 184630 129415
rect 149162 129375 184630 129403
rect 149162 129363 149168 129375
rect 184624 129363 184630 129375
rect 184682 129363 184688 129415
rect 154000 129289 154006 129341
rect 154058 129329 154064 129341
rect 184336 129329 184342 129341
rect 154058 129301 184342 129329
rect 154058 129289 154064 129301
rect 184336 129289 184342 129301
rect 184394 129289 184400 129341
rect 655216 127069 655222 127121
rect 655274 127109 655280 127121
rect 676240 127109 676246 127121
rect 655274 127081 676246 127109
rect 655274 127069 655280 127081
rect 676240 127069 676246 127081
rect 676298 127069 676304 127121
rect 655120 126921 655126 126973
rect 655178 126961 655184 126973
rect 676336 126961 676342 126973
rect 655178 126933 676342 126961
rect 655178 126921 655184 126933
rect 676336 126921 676342 126933
rect 676394 126921 676400 126973
rect 647920 126773 647926 126825
rect 647978 126813 647984 126825
rect 676144 126813 676150 126825
rect 647978 126785 676150 126813
rect 647978 126773 647984 126785
rect 676144 126773 676150 126785
rect 676202 126773 676208 126825
rect 149392 126699 149398 126751
rect 149450 126739 149456 126751
rect 156880 126739 156886 126751
rect 149450 126711 156886 126739
rect 149450 126699 149456 126711
rect 156880 126699 156886 126711
rect 156938 126699 156944 126751
rect 646576 126699 646582 126751
rect 646634 126739 646640 126751
rect 676048 126739 676054 126751
rect 646634 126711 676054 126739
rect 646634 126699 646640 126711
rect 676048 126699 676054 126711
rect 676106 126699 676112 126751
rect 148528 126625 148534 126677
rect 148586 126665 148592 126677
rect 184528 126665 184534 126677
rect 148586 126637 184534 126665
rect 148586 126625 148592 126637
rect 184528 126625 184534 126637
rect 184586 126625 184592 126677
rect 148720 126551 148726 126603
rect 148778 126591 148784 126603
rect 184432 126591 184438 126603
rect 148778 126563 184438 126591
rect 148778 126551 148784 126563
rect 184432 126551 184438 126563
rect 184490 126551 184496 126603
rect 148912 126477 148918 126529
rect 148970 126517 148976 126529
rect 184336 126517 184342 126529
rect 148970 126489 184342 126517
rect 148970 126477 148976 126489
rect 184336 126477 184342 126489
rect 184394 126477 184400 126529
rect 673840 126329 673846 126381
rect 673898 126369 673904 126381
rect 676048 126369 676054 126381
rect 673898 126341 676054 126369
rect 673898 126329 673904 126341
rect 676048 126329 676054 126341
rect 676106 126329 676112 126381
rect 675184 123961 675190 124013
rect 675242 124001 675248 124013
rect 676048 124001 676054 124013
rect 675242 123973 676054 124001
rect 675242 123961 675248 123973
rect 676048 123961 676054 123973
rect 676106 123961 676112 124013
rect 148432 123887 148438 123939
rect 148490 123927 148496 123939
rect 154192 123927 154198 123939
rect 148490 123899 154198 123927
rect 148490 123887 148496 123899
rect 154192 123887 154198 123899
rect 154250 123887 154256 123939
rect 646480 123887 646486 123939
rect 646538 123927 646544 123939
rect 676240 123927 676246 123939
rect 646538 123899 676246 123927
rect 646538 123887 646544 123899
rect 676240 123887 676246 123899
rect 676298 123887 676304 123939
rect 148240 123813 148246 123865
rect 148298 123853 148304 123865
rect 184624 123853 184630 123865
rect 148298 123825 184630 123853
rect 148298 123813 148304 123825
rect 184624 123813 184630 123825
rect 184682 123813 184688 123865
rect 148528 123739 148534 123791
rect 148586 123779 148592 123791
rect 184432 123779 184438 123791
rect 148586 123751 184438 123779
rect 148586 123739 148592 123751
rect 184432 123739 184438 123751
rect 184490 123739 184496 123791
rect 148624 123665 148630 123717
rect 148682 123705 148688 123717
rect 184336 123705 184342 123717
rect 148682 123677 184342 123705
rect 148682 123665 148688 123677
rect 184336 123665 184342 123677
rect 184394 123665 184400 123717
rect 149680 123591 149686 123643
rect 149738 123631 149744 123643
rect 184528 123631 184534 123643
rect 149738 123603 184534 123631
rect 149738 123591 149744 123603
rect 184528 123591 184534 123603
rect 184586 123591 184592 123643
rect 674608 121149 674614 121201
rect 674666 121189 674672 121201
rect 675952 121189 675958 121201
rect 674666 121161 675958 121189
rect 674666 121149 674672 121161
rect 675952 121149 675958 121161
rect 676010 121149 676016 121201
rect 674704 121075 674710 121127
rect 674762 121115 674768 121127
rect 676240 121115 676246 121127
rect 674762 121087 676246 121115
rect 674762 121075 674768 121087
rect 676240 121075 676246 121087
rect 676298 121075 676304 121127
rect 674992 121001 674998 121053
rect 675050 121041 675056 121053
rect 676048 121041 676054 121053
rect 675050 121013 676054 121041
rect 675050 121001 675056 121013
rect 676048 121001 676054 121013
rect 676106 121001 676112 121053
rect 148336 120927 148342 120979
rect 148394 120967 148400 120979
rect 184432 120967 184438 120979
rect 148394 120939 184438 120967
rect 148394 120927 148400 120939
rect 184432 120927 184438 120939
rect 184490 120927 184496 120979
rect 149488 120853 149494 120905
rect 149546 120893 149552 120905
rect 184528 120893 184534 120905
rect 149546 120865 184534 120893
rect 149546 120853 149552 120865
rect 184528 120853 184534 120865
rect 184586 120853 184592 120905
rect 171376 120779 171382 120831
rect 171434 120819 171440 120831
rect 184624 120819 184630 120831
rect 171434 120791 184630 120819
rect 171434 120779 171440 120791
rect 184624 120779 184630 120791
rect 184682 120779 184688 120831
rect 174256 120705 174262 120757
rect 174314 120745 174320 120757
rect 184336 120745 184342 120757
rect 174314 120717 184342 120745
rect 174314 120705 174320 120717
rect 184336 120705 184342 120717
rect 184394 120705 184400 120757
rect 180016 120631 180022 120683
rect 180074 120671 180080 120683
rect 186256 120671 186262 120683
rect 180074 120643 186262 120671
rect 180074 120631 180080 120643
rect 186256 120631 186262 120643
rect 186314 120631 186320 120683
rect 674320 119891 674326 119943
rect 674378 119931 674384 119943
rect 676048 119931 676054 119943
rect 674378 119903 676054 119931
rect 674378 119891 674384 119903
rect 676048 119891 676054 119903
rect 676106 119891 676112 119943
rect 674800 118559 674806 118611
rect 674858 118599 674864 118611
rect 676240 118599 676246 118611
rect 674858 118571 676246 118599
rect 674858 118559 674864 118571
rect 676240 118559 676246 118571
rect 676298 118559 676304 118611
rect 646192 118411 646198 118463
rect 646250 118451 646256 118463
rect 676240 118451 676246 118463
rect 646250 118423 676246 118451
rect 646250 118411 646256 118423
rect 676240 118411 676246 118423
rect 676298 118411 676304 118463
rect 149392 118263 149398 118315
rect 149450 118303 149456 118315
rect 168496 118303 168502 118315
rect 149450 118275 168502 118303
rect 149450 118263 149456 118275
rect 168496 118263 168502 118275
rect 168554 118263 168560 118315
rect 149488 118189 149494 118241
rect 149546 118229 149552 118241
rect 174352 118229 174358 118241
rect 149546 118201 174358 118229
rect 149546 118189 149552 118201
rect 174352 118189 174358 118201
rect 174410 118189 174416 118241
rect 674416 118189 674422 118241
rect 674474 118229 674480 118241
rect 675952 118229 675958 118241
rect 674474 118201 675958 118229
rect 674474 118189 674480 118201
rect 675952 118189 675958 118201
rect 676010 118189 676016 118241
rect 149392 118115 149398 118167
rect 149450 118155 149456 118167
rect 180112 118155 180118 118167
rect 149450 118127 180118 118155
rect 149450 118115 149456 118127
rect 180112 118115 180118 118127
rect 180170 118115 180176 118167
rect 674896 118115 674902 118167
rect 674954 118155 674960 118167
rect 676048 118155 676054 118167
rect 674954 118127 676054 118155
rect 674954 118115 674960 118127
rect 676048 118115 676054 118127
rect 676106 118115 676112 118167
rect 159856 118041 159862 118093
rect 159914 118081 159920 118093
rect 184624 118081 184630 118093
rect 159914 118053 184630 118081
rect 159914 118041 159920 118053
rect 184624 118041 184630 118053
rect 184682 118041 184688 118093
rect 162928 117967 162934 118019
rect 162986 118007 162992 118019
rect 184528 118007 184534 118019
rect 162986 117979 184534 118007
rect 162986 117967 162992 117979
rect 184528 117967 184534 117979
rect 184586 117967 184592 118019
rect 165712 117893 165718 117945
rect 165770 117933 165776 117945
rect 184432 117933 184438 117945
rect 165770 117905 184438 117933
rect 165770 117893 165776 117905
rect 184432 117893 184438 117905
rect 184490 117893 184496 117945
rect 168400 117819 168406 117871
rect 168458 117859 168464 117871
rect 184336 117859 184342 117871
rect 168458 117831 184342 117859
rect 168458 117819 168464 117831
rect 184336 117819 184342 117831
rect 184394 117819 184400 117871
rect 647728 115451 647734 115503
rect 647786 115491 647792 115503
rect 676240 115491 676246 115503
rect 647786 115463 676246 115491
rect 647786 115451 647792 115463
rect 676240 115451 676246 115463
rect 676298 115451 676304 115503
rect 149392 115303 149398 115355
rect 149450 115343 149456 115355
rect 162736 115343 162742 115355
rect 149450 115315 162742 115343
rect 149450 115303 149456 115315
rect 162736 115303 162742 115315
rect 162794 115303 162800 115355
rect 647824 115303 647830 115355
rect 647882 115343 647888 115355
rect 676144 115343 676150 115355
rect 647882 115315 676150 115343
rect 647882 115303 647888 115315
rect 676144 115303 676150 115315
rect 676202 115303 676208 115355
rect 149488 115229 149494 115281
rect 149546 115269 149552 115281
rect 165520 115269 165526 115281
rect 149546 115241 165526 115269
rect 149546 115229 149552 115241
rect 165520 115229 165526 115241
rect 165578 115229 165584 115281
rect 647920 115229 647926 115281
rect 647978 115269 647984 115281
rect 665296 115269 665302 115281
rect 647978 115241 665302 115269
rect 647978 115229 647984 115241
rect 665296 115229 665302 115241
rect 665354 115229 665360 115281
rect 151408 115155 151414 115207
rect 151466 115195 151472 115207
rect 184624 115195 184630 115207
rect 151466 115167 184630 115195
rect 151466 115155 151472 115167
rect 184624 115155 184630 115167
rect 184682 115155 184688 115207
rect 154096 115081 154102 115133
rect 154154 115121 154160 115133
rect 184432 115121 184438 115133
rect 154154 115093 184438 115121
rect 154154 115081 154160 115093
rect 184432 115081 184438 115093
rect 184490 115081 184496 115133
rect 156976 115007 156982 115059
rect 157034 115047 157040 115059
rect 184336 115047 184342 115059
rect 157034 115019 184342 115047
rect 157034 115007 157040 115019
rect 184336 115007 184342 115019
rect 184394 115007 184400 115059
rect 159760 114933 159766 114985
rect 159818 114973 159824 114985
rect 184528 114973 184534 114985
rect 159818 114945 184534 114973
rect 159818 114933 159824 114945
rect 184528 114933 184534 114945
rect 184586 114933 184592 114985
rect 663760 114637 663766 114689
rect 663818 114677 663824 114689
rect 675376 114677 675382 114689
rect 663818 114649 675382 114677
rect 663818 114637 663824 114649
rect 675376 114637 675382 114649
rect 675434 114637 675440 114689
rect 177232 113897 177238 113949
rect 177290 113937 177296 113949
rect 184720 113937 184726 113949
rect 177290 113909 184726 113937
rect 177290 113897 177296 113909
rect 184720 113897 184726 113909
rect 184778 113897 184784 113949
rect 149488 112713 149494 112765
rect 149546 112753 149552 112765
rect 159856 112753 159862 112765
rect 149546 112725 159862 112753
rect 149546 112713 149552 112725
rect 159856 112713 159862 112725
rect 159914 112713 159920 112765
rect 149392 112343 149398 112395
rect 149450 112383 149456 112395
rect 177136 112383 177142 112395
rect 149450 112355 177142 112383
rect 149450 112343 149456 112355
rect 177136 112343 177142 112355
rect 177194 112343 177200 112395
rect 151216 112269 151222 112321
rect 151274 112309 151280 112321
rect 184336 112309 184342 112321
rect 151274 112281 184342 112309
rect 151274 112269 151280 112281
rect 184336 112269 184342 112281
rect 184394 112269 184400 112321
rect 182800 112195 182806 112247
rect 182858 112235 182864 112247
rect 184528 112235 184534 112247
rect 182858 112207 184534 112235
rect 182858 112195 182864 112207
rect 184528 112195 184534 112207
rect 184586 112195 184592 112247
rect 674608 110271 674614 110323
rect 674666 110311 674672 110323
rect 675376 110311 675382 110323
rect 674666 110283 675382 110311
rect 674666 110271 674672 110283
rect 675376 110271 675382 110283
rect 675434 110271 675440 110323
rect 674704 109679 674710 109731
rect 674762 109719 674768 109731
rect 675472 109719 675478 109731
rect 674762 109691 675478 109719
rect 674762 109679 674768 109691
rect 675472 109679 675478 109691
rect 675530 109679 675536 109731
rect 149392 109531 149398 109583
rect 149450 109571 149456 109583
rect 156976 109571 156982 109583
rect 149450 109543 156982 109571
rect 149450 109531 149456 109543
rect 156976 109531 156982 109543
rect 157034 109531 157040 109583
rect 162640 109383 162646 109435
rect 162698 109423 162704 109435
rect 184336 109423 184342 109435
rect 162698 109395 184342 109423
rect 162698 109383 162704 109395
rect 184336 109383 184342 109395
rect 184394 109383 184400 109435
rect 179920 109309 179926 109361
rect 179978 109349 179984 109361
rect 185296 109349 185302 109361
rect 179978 109321 185302 109349
rect 179978 109309 179984 109321
rect 185296 109309 185302 109321
rect 185354 109309 185360 109361
rect 177040 109235 177046 109287
rect 177098 109275 177104 109287
rect 184432 109275 184438 109287
rect 177098 109247 184438 109275
rect 177098 109235 177104 109247
rect 184432 109235 184438 109247
rect 184490 109235 184496 109287
rect 674896 109013 674902 109065
rect 674954 109053 674960 109065
rect 675376 109053 675382 109065
rect 674954 109025 675382 109053
rect 674954 109013 674960 109025
rect 675376 109013 675382 109025
rect 675434 109013 675440 109065
rect 147856 108347 147862 108399
rect 147914 108387 147920 108399
rect 154000 108387 154006 108399
rect 147914 108359 154006 108387
rect 147914 108347 147920 108359
rect 154000 108347 154006 108359
rect 154058 108347 154064 108399
rect 154192 107977 154198 108029
rect 154250 108017 154256 108029
rect 184624 108017 184630 108029
rect 154250 107989 184630 108017
rect 154250 107977 154256 107989
rect 184624 107977 184630 107989
rect 184682 107977 184688 108029
rect 147184 107163 147190 107215
rect 147242 107203 147248 107215
rect 151120 107203 151126 107215
rect 147242 107175 151126 107203
rect 147242 107163 147248 107175
rect 151120 107163 151126 107175
rect 151178 107163 151184 107215
rect 182896 106497 182902 106549
rect 182954 106537 182960 106549
rect 186640 106537 186646 106549
rect 182954 106509 186646 106537
rect 182954 106497 182960 106509
rect 186640 106497 186646 106509
rect 186698 106497 186704 106549
rect 171280 106423 171286 106475
rect 171338 106463 171344 106475
rect 184528 106463 184534 106475
rect 171338 106435 184534 106463
rect 171338 106423 171344 106435
rect 184528 106423 184534 106435
rect 184586 106423 184592 106475
rect 174160 106349 174166 106401
rect 174218 106389 174224 106401
rect 184336 106389 184342 106401
rect 174218 106361 184342 106389
rect 174218 106349 174224 106361
rect 184336 106349 184342 106361
rect 184394 106349 184400 106401
rect 149584 106275 149590 106327
rect 149642 106315 149648 106327
rect 184432 106315 184438 106327
rect 149642 106287 184438 106315
rect 149642 106275 149648 106287
rect 184432 106275 184438 106287
rect 184490 106275 184496 106327
rect 674896 105905 674902 105957
rect 674954 105945 674960 105957
rect 675472 105945 675478 105957
rect 674954 105917 675478 105945
rect 674954 105905 674960 105917
rect 675472 105905 675478 105917
rect 675530 105905 675536 105957
rect 674320 105239 674326 105291
rect 674378 105279 674384 105291
rect 675376 105279 675382 105291
rect 674378 105251 675382 105279
rect 674378 105239 674384 105251
rect 675376 105239 675382 105251
rect 675434 105239 675440 105291
rect 674416 104721 674422 104773
rect 674474 104761 674480 104773
rect 675376 104761 675382 104773
rect 674474 104733 675382 104761
rect 674474 104721 674480 104733
rect 675376 104721 675382 104733
rect 675434 104721 675440 104773
rect 654064 104499 654070 104551
rect 654122 104539 654128 104551
rect 665584 104539 665590 104551
rect 654122 104511 665590 104539
rect 654122 104499 654128 104511
rect 665584 104499 665590 104511
rect 665642 104499 665648 104551
rect 645904 103833 645910 103885
rect 645962 103873 645968 103885
rect 657520 103873 657526 103885
rect 645962 103845 657526 103873
rect 645962 103833 645968 103845
rect 657520 103833 657526 103845
rect 657578 103833 657584 103885
rect 647920 103759 647926 103811
rect 647978 103799 647984 103811
rect 661168 103799 661174 103811
rect 647978 103771 661174 103799
rect 647978 103759 647984 103771
rect 661168 103759 661174 103771
rect 661226 103759 661232 103811
rect 149104 103611 149110 103663
rect 149162 103651 149168 103663
rect 184528 103651 184534 103663
rect 149162 103623 184534 103651
rect 149162 103611 149168 103623
rect 184528 103611 184534 103623
rect 184586 103611 184592 103663
rect 149008 103537 149014 103589
rect 149066 103577 149072 103589
rect 184336 103577 184342 103589
rect 149066 103549 184342 103577
rect 149066 103537 149072 103549
rect 184336 103537 184342 103549
rect 184394 103537 184400 103589
rect 165616 103463 165622 103515
rect 165674 103503 165680 103515
rect 184432 103503 184438 103515
rect 165674 103475 184438 103503
rect 165674 103463 165680 103475
rect 184432 103463 184438 103475
rect 184490 103463 184496 103515
rect 645136 102057 645142 102109
rect 645194 102097 645200 102109
rect 652432 102097 652438 102109
rect 645194 102069 652438 102097
rect 645194 102057 645200 102069
rect 652432 102057 652438 102069
rect 652490 102057 652496 102109
rect 149392 100799 149398 100851
rect 149450 100839 149456 100851
rect 168400 100839 168406 100851
rect 149450 100811 168406 100839
rect 149450 100799 149456 100811
rect 168400 100799 168406 100811
rect 168458 100799 168464 100851
rect 149680 100725 149686 100777
rect 149738 100765 149744 100777
rect 184528 100765 184534 100777
rect 149738 100737 184534 100765
rect 149738 100725 149744 100737
rect 184528 100725 184534 100737
rect 184586 100725 184592 100777
rect 149296 100651 149302 100703
rect 149354 100691 149360 100703
rect 184432 100691 184438 100703
rect 149354 100663 184438 100691
rect 149354 100651 149360 100663
rect 184432 100651 184438 100663
rect 184490 100651 184496 100703
rect 156880 100577 156886 100629
rect 156938 100617 156944 100629
rect 184336 100617 184342 100629
rect 156938 100589 184342 100617
rect 156938 100577 156944 100589
rect 184336 100577 184342 100589
rect 184394 100577 184400 100629
rect 149392 97987 149398 98039
rect 149450 98027 149456 98039
rect 184240 98027 184246 98039
rect 149450 97999 184246 98027
rect 149450 97987 149456 97999
rect 184240 97987 184246 97999
rect 184298 97987 184304 98039
rect 149488 97913 149494 97965
rect 149546 97953 149552 97965
rect 186160 97953 186166 97965
rect 149546 97925 186166 97953
rect 149546 97913 149552 97925
rect 186160 97913 186166 97925
rect 186218 97913 186224 97965
rect 647920 97913 647926 97965
rect 647978 97953 647984 97965
rect 662512 97953 662518 97965
rect 647978 97925 662518 97953
rect 647978 97913 647984 97925
rect 662512 97913 662518 97925
rect 662570 97913 662576 97965
rect 148528 97839 148534 97891
rect 148586 97879 148592 97891
rect 184336 97879 184342 97891
rect 148586 97851 184342 97879
rect 148586 97839 148592 97851
rect 184336 97839 184342 97851
rect 184394 97839 184400 97891
rect 148624 97765 148630 97817
rect 148682 97805 148688 97817
rect 184432 97805 184438 97817
rect 148682 97777 184438 97805
rect 148682 97765 148688 97777
rect 184432 97765 184438 97777
rect 184490 97765 184496 97817
rect 168496 97691 168502 97743
rect 168554 97731 168560 97743
rect 184528 97731 184534 97743
rect 168554 97703 184534 97731
rect 168554 97691 168560 97703
rect 184528 97691 184534 97703
rect 184586 97691 184592 97743
rect 640720 96507 640726 96559
rect 640778 96547 640784 96559
rect 654064 96547 654070 96559
rect 640778 96519 654070 96547
rect 640778 96507 640784 96519
rect 654064 96507 654070 96519
rect 654122 96507 654128 96559
rect 645424 95915 645430 95967
rect 645482 95955 645488 95967
rect 653680 95955 653686 95967
rect 645482 95927 653686 95955
rect 645482 95915 645488 95927
rect 653680 95915 653686 95927
rect 653738 95915 653744 95967
rect 149488 95101 149494 95153
rect 149546 95141 149552 95153
rect 166672 95141 166678 95153
rect 149546 95113 166678 95141
rect 149546 95101 149552 95113
rect 166672 95101 166678 95113
rect 166730 95101 166736 95153
rect 149392 95027 149398 95079
rect 149450 95067 149456 95079
rect 179920 95067 179926 95079
rect 149450 95039 179926 95067
rect 149450 95027 149456 95039
rect 179920 95027 179926 95039
rect 179978 95027 179984 95079
rect 162736 94953 162742 95005
rect 162794 94993 162800 95005
rect 184528 94993 184534 95005
rect 162794 94965 184534 94993
rect 162794 94953 162800 94965
rect 184528 94953 184534 94965
rect 184586 94953 184592 95005
rect 165520 94879 165526 94931
rect 165578 94919 165584 94931
rect 184432 94919 184438 94931
rect 165578 94891 184438 94919
rect 165578 94879 165584 94891
rect 184432 94879 184438 94891
rect 184490 94879 184496 94931
rect 174352 94805 174358 94857
rect 174410 94845 174416 94857
rect 184336 94845 184342 94857
rect 174410 94817 184342 94845
rect 174410 94805 174416 94817
rect 184336 94805 184342 94817
rect 184394 94805 184400 94857
rect 180112 94583 180118 94635
rect 180170 94623 180176 94635
rect 184624 94623 184630 94635
rect 180170 94595 184630 94623
rect 180170 94583 180176 94595
rect 184624 94583 184630 94595
rect 184682 94583 184688 94635
rect 646768 92659 646774 92711
rect 646826 92699 646832 92711
rect 663088 92699 663094 92711
rect 646826 92671 663094 92699
rect 646826 92659 646832 92671
rect 663088 92659 663094 92671
rect 663146 92659 663152 92711
rect 149392 92363 149398 92415
rect 149450 92403 149456 92415
rect 159568 92403 159574 92415
rect 149450 92375 159574 92403
rect 149450 92363 149456 92375
rect 159568 92363 159574 92375
rect 159626 92363 159632 92415
rect 646480 92363 646486 92415
rect 646538 92403 646544 92415
rect 660688 92403 660694 92415
rect 646538 92375 660694 92403
rect 646538 92363 646544 92375
rect 660688 92363 660694 92375
rect 660746 92363 660752 92415
rect 645520 92289 645526 92341
rect 645578 92329 645584 92341
rect 661744 92329 661750 92341
rect 645578 92301 661750 92329
rect 645578 92289 645584 92301
rect 661744 92289 661750 92301
rect 661802 92289 661808 92341
rect 646864 92215 646870 92267
rect 646922 92255 646928 92267
rect 659824 92255 659830 92267
rect 646922 92227 659830 92255
rect 646922 92215 646928 92227
rect 659824 92215 659830 92227
rect 659882 92215 659888 92267
rect 149488 92141 149494 92193
rect 149546 92181 149552 92193
rect 162352 92181 162358 92193
rect 149546 92153 162358 92181
rect 149546 92141 149552 92153
rect 162352 92141 162358 92153
rect 162410 92141 162416 92193
rect 647056 92141 647062 92193
rect 647114 92181 647120 92193
rect 658864 92181 658870 92193
rect 647114 92153 658870 92181
rect 647114 92141 647120 92153
rect 658864 92141 658870 92153
rect 658922 92141 658928 92193
rect 148336 92067 148342 92119
rect 148394 92107 148400 92119
rect 184528 92107 184534 92119
rect 148394 92079 184534 92107
rect 148394 92067 148400 92079
rect 184528 92067 184534 92079
rect 184586 92067 184592 92119
rect 148720 91993 148726 92045
rect 148778 92033 148784 92045
rect 184432 92033 184438 92045
rect 148778 92005 184438 92033
rect 148778 91993 148784 92005
rect 184432 91993 184438 92005
rect 184490 91993 184496 92045
rect 159856 91919 159862 91971
rect 159914 91959 159920 91971
rect 184336 91959 184342 91971
rect 159914 91931 184342 91959
rect 159914 91919 159920 91931
rect 184336 91919 184342 91931
rect 184394 91919 184400 91971
rect 177136 91845 177142 91897
rect 177194 91885 177200 91897
rect 184624 91885 184630 91897
rect 177194 91857 184630 91885
rect 177194 91845 177200 91857
rect 184624 91845 184630 91857
rect 184682 91845 184688 91897
rect 148816 89181 148822 89233
rect 148874 89221 148880 89233
rect 184624 89221 184630 89233
rect 148874 89193 184630 89221
rect 148874 89181 148880 89193
rect 184624 89181 184630 89193
rect 184682 89181 184688 89233
rect 151120 89107 151126 89159
rect 151178 89147 151184 89159
rect 184528 89147 184534 89159
rect 151178 89119 184534 89147
rect 151178 89107 151184 89119
rect 184528 89107 184534 89119
rect 184586 89107 184592 89159
rect 154000 89033 154006 89085
rect 154058 89073 154064 89085
rect 184432 89073 184438 89085
rect 154058 89045 184438 89073
rect 154058 89033 154064 89045
rect 184432 89033 184438 89045
rect 184490 89033 184496 89085
rect 156976 88959 156982 89011
rect 157034 88999 157040 89011
rect 184336 88999 184342 89011
rect 157034 88971 184342 88999
rect 157034 88959 157040 88971
rect 184336 88959 184342 88971
rect 184394 88959 184400 89011
rect 645904 87479 645910 87531
rect 645962 87519 645968 87531
rect 650896 87519 650902 87531
rect 645962 87491 650902 87519
rect 645962 87479 645968 87491
rect 650896 87479 650902 87491
rect 650954 87479 650960 87531
rect 647920 87257 647926 87309
rect 647978 87297 647984 87309
rect 658000 87297 658006 87309
rect 647978 87269 658006 87297
rect 647978 87257 647984 87269
rect 658000 87257 658006 87269
rect 658058 87257 658064 87309
rect 647152 87035 647158 87087
rect 647210 87075 647216 87087
rect 663280 87075 663286 87087
rect 647210 87047 663286 87075
rect 647210 87035 647216 87047
rect 663280 87035 663286 87047
rect 663338 87035 663344 87087
rect 149488 86739 149494 86791
rect 149546 86779 149552 86791
rect 156400 86779 156406 86791
rect 149546 86751 156406 86779
rect 149546 86739 149552 86751
rect 156400 86739 156406 86751
rect 156458 86739 156464 86791
rect 148720 86443 148726 86495
rect 148778 86483 148784 86495
rect 154096 86483 154102 86495
rect 148778 86455 154102 86483
rect 148778 86443 148784 86455
rect 154096 86443 154102 86455
rect 154154 86443 154160 86495
rect 148432 86369 148438 86421
rect 148490 86409 148496 86421
rect 184528 86409 184534 86421
rect 148490 86381 184534 86409
rect 148490 86369 148496 86381
rect 184528 86369 184534 86381
rect 184586 86369 184592 86421
rect 148240 86295 148246 86347
rect 148298 86335 148304 86347
rect 184336 86335 184342 86347
rect 148298 86307 184342 86335
rect 148298 86295 148304 86307
rect 184336 86295 184342 86307
rect 184394 86295 184400 86347
rect 148912 86221 148918 86273
rect 148970 86261 148976 86273
rect 184432 86261 184438 86273
rect 148970 86233 184438 86261
rect 148970 86221 148976 86233
rect 184432 86221 184438 86233
rect 184490 86221 184496 86273
rect 645904 84001 645910 84053
rect 645962 84041 645968 84053
rect 657040 84041 657046 84053
rect 645962 84013 657046 84041
rect 645962 84001 645968 84013
rect 657040 84001 657046 84013
rect 657098 84001 657104 84053
rect 146992 83557 146998 83609
rect 147050 83597 147056 83609
rect 151120 83597 151126 83609
rect 147050 83569 151126 83597
rect 147050 83557 147056 83569
rect 151120 83557 151126 83569
rect 151178 83557 151184 83609
rect 646768 83557 646774 83609
rect 646826 83597 646832 83609
rect 651760 83597 651766 83609
rect 646826 83569 651766 83597
rect 646826 83557 646832 83569
rect 651760 83557 651766 83569
rect 651818 83557 651824 83609
rect 166672 83483 166678 83535
rect 166730 83523 166736 83535
rect 184432 83523 184438 83535
rect 166730 83495 184438 83523
rect 166730 83483 166736 83495
rect 184432 83483 184438 83495
rect 184490 83483 184496 83535
rect 168400 83409 168406 83461
rect 168458 83449 168464 83461
rect 184336 83449 184342 83461
rect 168458 83421 184342 83449
rect 168458 83409 168464 83421
rect 184336 83409 184342 83421
rect 184394 83409 184400 83461
rect 647920 81855 647926 81907
rect 647978 81895 647984 81907
rect 663280 81895 663286 81907
rect 647978 81867 663286 81895
rect 647978 81855 647984 81867
rect 663280 81855 663286 81867
rect 663338 81855 663344 81907
rect 657040 81633 657046 81685
rect 657098 81673 657104 81685
rect 658576 81673 658582 81685
rect 657098 81645 658582 81673
rect 657098 81633 657104 81645
rect 658576 81633 658582 81645
rect 658634 81633 658640 81685
rect 647824 81559 647830 81611
rect 647882 81599 647888 81611
rect 662416 81599 662422 81611
rect 647882 81571 662422 81599
rect 647882 81559 647888 81571
rect 662416 81559 662422 81571
rect 662474 81559 662480 81611
rect 647728 81485 647734 81537
rect 647786 81525 647792 81537
rect 663472 81525 663478 81537
rect 647786 81497 663478 81525
rect 647786 81485 647792 81497
rect 663472 81485 663478 81497
rect 663530 81485 663536 81537
rect 647920 80745 647926 80797
rect 647978 80785 647984 80797
rect 662512 80785 662518 80797
rect 647978 80757 662518 80785
rect 647978 80745 647984 80757
rect 662512 80745 662518 80757
rect 662570 80745 662576 80797
rect 659440 80671 659446 80723
rect 659498 80711 659504 80723
rect 659536 80711 659542 80723
rect 659498 80683 659542 80711
rect 659498 80671 659504 80683
rect 659536 80671 659542 80683
rect 659594 80671 659600 80723
rect 149584 80597 149590 80649
rect 149642 80637 149648 80649
rect 184432 80637 184438 80649
rect 149642 80609 184438 80637
rect 149642 80597 149648 80609
rect 184432 80597 184438 80609
rect 184490 80597 184496 80649
rect 159568 80523 159574 80575
rect 159626 80563 159632 80575
rect 184528 80563 184534 80575
rect 159626 80535 184534 80563
rect 159626 80523 159632 80535
rect 184528 80523 184534 80535
rect 184586 80523 184592 80575
rect 162352 80449 162358 80501
rect 162410 80489 162416 80501
rect 184336 80489 184342 80501
rect 162410 80461 184342 80489
rect 162410 80449 162416 80461
rect 184336 80449 184342 80461
rect 184394 80449 184400 80501
rect 179920 80375 179926 80427
rect 179978 80415 179984 80427
rect 184624 80415 184630 80427
rect 179978 80387 184630 80415
rect 179978 80375 179984 80387
rect 184624 80375 184630 80387
rect 184682 80375 184688 80427
rect 149296 77711 149302 77763
rect 149354 77751 149360 77763
rect 184432 77751 184438 77763
rect 149354 77723 184438 77751
rect 149354 77711 149360 77723
rect 184432 77711 184438 77723
rect 184490 77711 184496 77763
rect 646960 77711 646966 77763
rect 647018 77751 647024 77763
rect 658288 77751 658294 77763
rect 647018 77723 658294 77751
rect 647018 77711 647024 77723
rect 658288 77711 658294 77723
rect 658346 77711 658352 77763
rect 149392 77637 149398 77689
rect 149450 77677 149456 77689
rect 184624 77677 184630 77689
rect 149450 77649 184630 77677
rect 149450 77637 149456 77649
rect 184624 77637 184630 77649
rect 184682 77637 184688 77689
rect 646576 77637 646582 77689
rect 646634 77677 646640 77689
rect 659440 77677 659446 77689
rect 646634 77649 659446 77677
rect 646634 77637 646640 77649
rect 659440 77637 659446 77649
rect 659498 77637 659504 77689
rect 149200 77563 149206 77615
rect 149258 77603 149264 77615
rect 184336 77603 184342 77615
rect 149258 77575 184342 77603
rect 149258 77563 149264 77575
rect 184336 77563 184342 77575
rect 184394 77563 184400 77615
rect 646672 77563 646678 77615
rect 646730 77603 646736 77615
rect 661744 77603 661750 77615
rect 646730 77575 661750 77603
rect 646730 77563 646736 77575
rect 661744 77563 661750 77575
rect 661802 77563 661808 77615
rect 156400 77489 156406 77541
rect 156458 77529 156464 77541
rect 184528 77529 184534 77541
rect 156458 77501 184534 77529
rect 156458 77489 156464 77501
rect 184528 77489 184534 77501
rect 184586 77489 184592 77541
rect 647920 77489 647926 77541
rect 647978 77529 647984 77541
rect 656944 77529 656950 77541
rect 647978 77501 656950 77529
rect 647978 77489 647984 77501
rect 656944 77489 656950 77501
rect 657002 77489 657008 77541
rect 646000 76083 646006 76135
rect 646058 76123 646064 76135
rect 657520 76123 657526 76135
rect 646058 76095 657526 76123
rect 646058 76083 646064 76095
rect 657520 76083 657526 76095
rect 657578 76083 657584 76135
rect 647152 74899 647158 74951
rect 647210 74939 647216 74951
rect 660112 74939 660118 74951
rect 647210 74911 660118 74939
rect 647210 74899 647216 74911
rect 660112 74899 660118 74911
rect 660170 74899 660176 74951
rect 148624 74825 148630 74877
rect 148682 74865 148688 74877
rect 184528 74865 184534 74877
rect 148682 74837 184534 74865
rect 148682 74825 148688 74837
rect 184528 74825 184534 74837
rect 184586 74825 184592 74877
rect 148912 74751 148918 74803
rect 148970 74791 148976 74803
rect 184624 74791 184630 74803
rect 148970 74763 184630 74791
rect 148970 74751 148976 74763
rect 184624 74751 184630 74763
rect 184682 74751 184688 74803
rect 151120 74677 151126 74729
rect 151178 74717 151184 74729
rect 184432 74717 184438 74729
rect 151178 74689 184438 74717
rect 151178 74677 151184 74689
rect 184432 74677 184438 74689
rect 184490 74677 184496 74729
rect 154096 74603 154102 74655
rect 154154 74643 154160 74655
rect 184336 74643 184342 74655
rect 154154 74615 184342 74643
rect 154154 74603 154160 74615
rect 184336 74603 184342 74615
rect 184394 74603 184400 74655
rect 647920 72087 647926 72139
rect 647978 72127 647984 72139
rect 660688 72127 660694 72139
rect 647978 72099 660694 72127
rect 647978 72087 647984 72099
rect 660688 72087 660694 72099
rect 660746 72087 660752 72139
rect 148240 71939 148246 71991
rect 148298 71979 148304 71991
rect 184336 71979 184342 71991
rect 148298 71951 184342 71979
rect 148298 71939 148304 71951
rect 184336 71939 184342 71951
rect 184394 71939 184400 71991
rect 149584 71865 149590 71917
rect 149642 71905 149648 71917
rect 184432 71905 184438 71917
rect 149642 71877 184438 71905
rect 149642 71865 149648 71877
rect 184432 71865 184438 71877
rect 184490 71865 184496 71917
rect 149680 71791 149686 71843
rect 149738 71831 149744 71843
rect 184528 71831 184534 71843
rect 149738 71803 184534 71831
rect 149738 71791 149744 71803
rect 184528 71791 184534 71803
rect 184586 71791 184592 71843
rect 647920 69571 647926 69623
rect 647978 69611 647984 69623
rect 661456 69611 661462 69623
rect 647978 69583 661462 69611
rect 647978 69571 647984 69583
rect 661456 69571 661462 69583
rect 661514 69571 661520 69623
rect 148816 69053 148822 69105
rect 148874 69093 148880 69105
rect 184336 69093 184342 69105
rect 148874 69065 184342 69093
rect 148874 69053 148880 69065
rect 184336 69053 184342 69065
rect 184394 69053 184400 69105
rect 149584 68979 149590 69031
rect 149642 69019 149648 69031
rect 184432 69019 184438 69031
rect 149642 68991 184438 69019
rect 149642 68979 149648 68991
rect 184432 68979 184438 68991
rect 184490 68979 184496 69031
rect 149296 68905 149302 68957
rect 149354 68945 149360 68957
rect 184528 68945 184534 68957
rect 149354 68917 184534 68945
rect 149354 68905 149360 68917
rect 184528 68905 184534 68917
rect 184586 68905 184592 68957
rect 149200 68831 149206 68883
rect 149258 68871 149264 68883
rect 184336 68871 184342 68883
rect 149258 68843 184342 68871
rect 149258 68831 149264 68843
rect 184336 68831 184342 68843
rect 184394 68831 184400 68883
rect 149104 66167 149110 66219
rect 149162 66207 149168 66219
rect 184528 66207 184534 66219
rect 149162 66179 184534 66207
rect 149162 66167 149168 66179
rect 184528 66167 184534 66179
rect 184586 66167 184592 66219
rect 646000 66167 646006 66219
rect 646058 66207 646064 66219
rect 652336 66207 652342 66219
rect 646058 66179 652342 66207
rect 646058 66167 646064 66179
rect 652336 66167 652342 66179
rect 652394 66167 652400 66219
rect 149488 66093 149494 66145
rect 149546 66133 149552 66145
rect 184624 66133 184630 66145
rect 149546 66105 184630 66133
rect 149546 66093 149552 66105
rect 184624 66093 184630 66105
rect 184682 66093 184688 66145
rect 149392 66019 149398 66071
rect 149450 66059 149456 66071
rect 184432 66059 184438 66071
rect 149450 66031 184438 66059
rect 149450 66019 149456 66031
rect 184432 66019 184438 66031
rect 184490 66019 184496 66071
rect 149008 65945 149014 65997
rect 149066 65985 149072 65997
rect 184336 65985 184342 65997
rect 149066 65957 184342 65985
rect 149066 65945 149072 65957
rect 184336 65945 184342 65957
rect 184394 65945 184400 65997
rect 647920 63429 647926 63481
rect 647978 63469 647984 63481
rect 663184 63469 663190 63481
rect 647978 63441 663190 63469
rect 647978 63429 647984 63441
rect 663184 63429 663190 63441
rect 663242 63429 663248 63481
rect 149584 63281 149590 63333
rect 149642 63321 149648 63333
rect 184432 63321 184438 63333
rect 149642 63293 184438 63321
rect 149642 63281 149648 63293
rect 184432 63281 184438 63293
rect 184490 63281 184496 63333
rect 149488 63207 149494 63259
rect 149546 63247 149552 63259
rect 184528 63247 184534 63259
rect 149546 63219 184534 63247
rect 149546 63207 149552 63219
rect 184528 63207 184534 63219
rect 184586 63207 184592 63259
rect 149392 63133 149398 63185
rect 149450 63173 149456 63185
rect 184624 63173 184630 63185
rect 149450 63145 184630 63173
rect 149450 63133 149456 63145
rect 184624 63133 184630 63145
rect 184682 63133 184688 63185
rect 149200 63059 149206 63111
rect 149258 63099 149264 63111
rect 184336 63099 184342 63111
rect 149258 63071 184342 63099
rect 149258 63059 149264 63071
rect 184336 63059 184342 63071
rect 184394 63059 184400 63111
rect 647920 60987 647926 61039
rect 647978 61027 647984 61039
rect 663376 61027 663382 61039
rect 647978 60999 663382 61027
rect 647978 60987 647984 60999
rect 663376 60987 663382 60999
rect 663434 60987 663440 61039
rect 149392 60395 149398 60447
rect 149450 60435 149456 60447
rect 184528 60435 184534 60447
rect 149450 60407 184534 60435
rect 149450 60395 149456 60407
rect 184528 60395 184534 60407
rect 184586 60395 184592 60447
rect 149296 60321 149302 60373
rect 149354 60361 149360 60373
rect 184336 60361 184342 60373
rect 149354 60333 184342 60361
rect 149354 60321 149360 60333
rect 184336 60321 184342 60333
rect 184394 60321 184400 60373
rect 149488 60247 149494 60299
rect 149546 60287 149552 60299
rect 184432 60287 184438 60299
rect 149546 60259 184438 60287
rect 149546 60247 149552 60259
rect 184432 60247 184438 60259
rect 184490 60247 184496 60299
rect 646000 59063 646006 59115
rect 646058 59103 646064 59115
rect 652240 59103 652246 59115
rect 646058 59075 652246 59103
rect 646058 59063 646064 59075
rect 652240 59063 652246 59075
rect 652298 59063 652304 59115
rect 149392 58989 149398 59041
rect 149450 59029 149456 59041
rect 184336 59029 184342 59041
rect 149450 59001 184342 59029
rect 149450 58989 149456 59001
rect 184336 58989 184342 59001
rect 184394 58989 184400 59041
rect 149392 57509 149398 57561
rect 149450 57549 149456 57561
rect 184336 57549 184342 57561
rect 149450 57521 184342 57549
rect 149450 57509 149456 57521
rect 184336 57509 184342 57521
rect 184394 57509 184400 57561
rect 149392 56177 149398 56229
rect 149450 56217 149456 56229
rect 184432 56217 184438 56229
rect 149450 56189 184438 56217
rect 149450 56177 149456 56189
rect 184432 56177 184438 56189
rect 184490 56177 184496 56229
rect 149488 56103 149494 56155
rect 149546 56143 149552 56155
rect 184336 56143 184342 56155
rect 149546 56115 184342 56143
rect 149546 56103 149552 56115
rect 184336 56103 184342 56115
rect 184394 56103 184400 56155
rect 149680 54623 149686 54675
rect 149738 54663 149744 54675
rect 184336 54663 184342 54675
rect 149738 54635 184342 54663
rect 149738 54623 149744 54635
rect 184336 54623 184342 54635
rect 184394 54623 184400 54675
rect 149392 53217 149398 53269
rect 149450 53257 149456 53269
rect 184336 53257 184342 53269
rect 149450 53229 184342 53257
rect 149450 53217 149456 53229
rect 184336 53217 184342 53229
rect 184394 53217 184400 53269
rect 418768 48407 418774 48459
rect 418826 48447 418832 48459
rect 424048 48447 424054 48459
rect 418826 48419 424054 48447
rect 418826 48407 418832 48419
rect 424048 48407 424054 48419
rect 424106 48407 424112 48459
rect 480976 48111 480982 48163
rect 481034 48151 481040 48163
rect 527920 48151 527926 48163
rect 481034 48123 527926 48151
rect 481034 48111 481040 48123
rect 527920 48111 527926 48123
rect 527978 48111 527984 48163
rect 460336 48037 460342 48089
rect 460394 48077 460400 48089
rect 510352 48077 510358 48089
rect 460394 48049 510358 48077
rect 460394 48037 460400 48049
rect 510352 48037 510358 48049
rect 510410 48037 510416 48089
rect 305296 47963 305302 48015
rect 305354 48003 305360 48015
rect 354832 48003 354838 48015
rect 305354 47975 354838 48003
rect 305354 47963 305360 47975
rect 354832 47963 354838 47975
rect 354890 47963 354896 48015
rect 426160 47963 426166 48015
rect 426218 48003 426224 48015
rect 492976 48003 492982 48015
rect 426218 47975 492982 48003
rect 426218 47963 426224 47975
rect 492976 47963 492982 47975
rect 493034 47963 493040 48015
rect 311056 47889 311062 47941
rect 311114 47929 311120 47941
rect 371920 47929 371926 47941
rect 311114 47901 371926 47929
rect 311114 47889 311120 47901
rect 371920 47889 371926 47901
rect 371978 47889 371984 47941
rect 405520 47889 405526 47941
rect 405578 47929 405584 47941
rect 441328 47929 441334 47941
rect 405578 47901 441334 47929
rect 405578 47889 405584 47901
rect 441328 47889 441334 47901
rect 441386 47889 441392 47941
rect 472240 47889 472246 47941
rect 472298 47929 472304 47941
rect 562480 47929 562486 47941
rect 472298 47901 562486 47929
rect 472298 47889 472304 47901
rect 562480 47889 562486 47901
rect 562538 47889 562544 47941
rect 302896 47815 302902 47867
rect 302954 47855 302960 47867
rect 506800 47855 506806 47867
rect 302954 47827 506806 47855
rect 302954 47815 302960 47827
rect 506800 47815 506806 47827
rect 506858 47815 506864 47867
rect 320176 47741 320182 47793
rect 320234 47781 320240 47793
rect 529264 47781 529270 47793
rect 320234 47753 529270 47781
rect 320234 47741 320240 47753
rect 529264 47741 529270 47753
rect 529322 47741 529328 47793
rect 233680 47667 233686 47719
rect 233738 47707 233744 47719
rect 475504 47707 475510 47719
rect 233738 47679 475510 47707
rect 233738 47667 233744 47679
rect 475504 47667 475510 47679
rect 475562 47667 475568 47719
rect 268528 47593 268534 47645
rect 268586 47633 268592 47645
rect 520624 47633 520630 47645
rect 268586 47605 520630 47633
rect 268586 47593 268592 47605
rect 520624 47593 520630 47605
rect 520682 47593 520688 47645
rect 250960 47519 250966 47571
rect 251018 47559 251024 47571
rect 521200 47559 521206 47571
rect 251018 47531 521206 47559
rect 251018 47519 251024 47531
rect 521200 47519 521206 47531
rect 521258 47519 521264 47571
rect 145360 47075 145366 47127
rect 145418 47115 145424 47127
rect 199120 47115 199126 47127
rect 145418 47087 199126 47115
rect 145418 47075 145424 47087
rect 199120 47075 199126 47087
rect 199178 47075 199184 47127
rect 328336 46705 328342 46757
rect 328394 46745 328400 46757
rect 337456 46745 337462 46757
rect 328394 46717 337462 46745
rect 328394 46705 328400 46717
rect 337456 46705 337462 46717
rect 337514 46705 337520 46757
rect 464848 46409 464854 46461
rect 464906 46449 464912 46461
rect 475696 46449 475702 46461
rect 464906 46421 475702 46449
rect 464906 46409 464912 46421
rect 475696 46409 475702 46421
rect 475754 46409 475760 46461
rect 207376 46187 207382 46239
rect 207434 46227 207440 46239
rect 216400 46227 216406 46239
rect 207434 46199 216406 46227
rect 207434 46187 207440 46199
rect 216400 46187 216406 46199
rect 216458 46187 216464 46239
rect 539728 46187 539734 46239
rect 539786 46227 539792 46239
rect 545200 46227 545206 46239
rect 539786 46199 545206 46227
rect 539786 46187 539792 46199
rect 545200 46187 545206 46199
rect 545258 46187 545264 46239
rect 401776 46113 401782 46165
rect 401834 46153 401840 46165
rect 406768 46153 406774 46165
rect 401834 46125 406774 46153
rect 401834 46113 401840 46125
rect 406768 46113 406774 46125
rect 406826 46113 406832 46165
rect 506800 44855 506806 44907
rect 506858 44895 506864 44907
rect 512176 44895 512182 44907
rect 506858 44867 512182 44895
rect 506858 44855 506864 44867
rect 512176 44855 512182 44867
rect 512234 44855 512240 44907
rect 630736 43671 630742 43723
rect 630794 43711 630800 43723
rect 640720 43711 640726 43723
rect 630794 43683 640726 43711
rect 630794 43671 630800 43683
rect 640720 43671 640726 43683
rect 640778 43671 640784 43723
rect 285808 43227 285814 43279
rect 285866 43267 285872 43279
rect 518704 43267 518710 43279
rect 285866 43239 518710 43267
rect 285866 43227 285872 43239
rect 518704 43227 518710 43239
rect 518762 43227 518768 43279
rect 302896 43153 302902 43205
rect 302954 43193 302960 43205
rect 305296 43193 305302 43205
rect 302954 43165 305302 43193
rect 302954 43153 302960 43165
rect 305296 43153 305302 43165
rect 305354 43153 305360 43205
rect 403216 43153 403222 43205
rect 403274 43193 403280 43205
rect 418768 43193 418774 43205
rect 403274 43165 418774 43193
rect 403274 43153 403280 43165
rect 418768 43153 418774 43165
rect 418826 43153 418832 43205
rect 444880 43153 444886 43205
rect 444938 43193 444944 43205
rect 458608 43193 458614 43205
rect 444938 43165 458614 43193
rect 444938 43153 444944 43165
rect 458608 43153 458614 43165
rect 458666 43153 458672 43205
rect 357712 42117 357718 42169
rect 357770 42157 357776 42169
rect 357770 42129 377294 42157
rect 357770 42117 357776 42129
rect 307216 42043 307222 42095
rect 307274 42083 307280 42095
rect 311056 42083 311062 42095
rect 307274 42055 311062 42083
rect 307274 42043 307280 42055
rect 311056 42043 311062 42055
rect 311114 42043 311120 42095
rect 362032 42043 362038 42095
rect 362090 42083 362096 42095
rect 365968 42083 365974 42095
rect 362090 42055 365974 42083
rect 362090 42043 362096 42055
rect 365968 42043 365974 42055
rect 366026 42043 366032 42095
rect 377266 42083 377294 42129
rect 401776 42083 401782 42095
rect 377266 42055 401782 42083
rect 401776 42043 401782 42055
rect 401834 42043 401840 42095
rect 471664 42043 471670 42095
rect 471722 42083 471728 42095
rect 480976 42083 480982 42095
rect 471722 42055 480982 42083
rect 471722 42043 471728 42055
rect 480976 42043 480982 42055
rect 481034 42043 481040 42095
rect 186256 41969 186262 42021
rect 186314 42009 186320 42021
rect 187024 42009 187030 42021
rect 186314 41981 187030 42009
rect 186314 41969 186320 41981
rect 187024 41969 187030 41981
rect 187082 41969 187088 42021
rect 194320 41969 194326 42021
rect 194378 42009 194384 42021
rect 630736 42009 630742 42021
rect 194378 41981 630742 42009
rect 194378 41969 194384 41981
rect 630736 41969 630742 41981
rect 630794 41969 630800 42021
rect 514000 41747 514006 41799
rect 514058 41787 514064 41799
rect 514864 41787 514870 41799
rect 514058 41759 514870 41787
rect 514058 41747 514064 41759
rect 514864 41747 514870 41759
rect 514922 41747 514928 41799
rect 186256 41451 186262 41503
rect 186314 41491 186320 41503
rect 207376 41491 207382 41503
rect 186314 41463 207382 41491
rect 186314 41451 186320 41463
rect 207376 41451 207382 41463
rect 207434 41451 207440 41503
rect 403216 37495 403222 37507
rect 397426 37467 403222 37495
rect 365872 37381 365878 37433
rect 365930 37421 365936 37433
rect 397426 37421 397454 37467
rect 403216 37455 403222 37467
rect 403274 37455 403280 37507
rect 365930 37393 397454 37421
rect 365930 37381 365936 37393
rect 475504 37381 475510 37433
rect 475562 37421 475568 37433
rect 514000 37421 514006 37433
rect 475562 37393 514006 37421
rect 475562 37381 475568 37393
rect 514000 37381 514006 37393
rect 514058 37381 514064 37433
rect 365968 37307 365974 37359
rect 366026 37347 366032 37359
rect 389200 37347 389206 37359
rect 366026 37319 389206 37347
rect 366026 37307 366032 37319
rect 389200 37307 389206 37319
rect 389258 37307 389264 37359
rect 420784 34495 420790 34547
rect 420842 34535 420848 34547
rect 444880 34535 444886 34547
rect 420842 34507 444886 34535
rect 420842 34495 420848 34507
rect 444880 34495 444886 34507
rect 444938 34495 444944 34547
<< via1 >>
rect 287926 993609 287978 993661
rect 291286 993609 291338 993661
rect 175606 992795 175658 992847
rect 178486 992795 178538 992847
rect 129526 984951 129578 985003
rect 132406 984951 132458 985003
rect 399574 983471 399626 983523
rect 432022 983471 432074 983523
rect 178582 982953 178634 983005
rect 184246 982953 184298 983005
rect 392470 982879 392522 982931
rect 394582 982805 394634 982857
rect 649462 982879 649514 982931
rect 652246 981991 652298 982043
rect 649462 981917 649514 981969
rect 656662 981917 656714 981969
rect 652246 979179 652298 979231
rect 679702 979179 679754 979231
rect 656662 974887 656714 974939
rect 671062 974887 671114 974939
rect 671062 963935 671114 963987
rect 677590 963935 677642 963987
rect 40150 961863 40202 961915
rect 60022 961863 60074 961915
rect 677494 959051 677546 959103
rect 679702 959051 679754 959103
rect 653782 944325 653834 944377
rect 676822 944325 676874 944377
rect 654262 878613 654314 878665
rect 676246 878613 676298 878665
rect 654166 878539 654218 878591
rect 676150 878539 676202 878591
rect 654070 878465 654122 878517
rect 676342 878465 676394 878517
rect 673366 878391 673418 878443
rect 676054 878391 676106 878443
rect 670870 877207 670922 877259
rect 676246 877207 676298 877259
rect 670966 876171 671018 876223
rect 676246 876171 676298 876223
rect 674038 872693 674090 872745
rect 676246 872693 676298 872745
rect 674326 872619 674378 872671
rect 676054 872619 676106 872671
rect 674134 870103 674186 870155
rect 676054 870103 676106 870155
rect 674902 869881 674954 869933
rect 676246 869881 676298 869933
rect 675094 869807 675146 869859
rect 676054 869807 676106 869859
rect 674998 869733 675050 869785
rect 679702 869733 679754 869785
rect 675190 869659 675242 869711
rect 679798 869659 679850 869711
rect 674518 866995 674570 867047
rect 676246 866995 676298 867047
rect 649462 866921 649514 866973
rect 679798 866921 679850 866973
rect 674614 864257 674666 864309
rect 679894 864257 679946 864309
rect 674998 864183 675050 864235
rect 680182 864183 680234 864235
rect 675286 864109 675338 864161
rect 680278 864109 680330 864161
rect 654262 864035 654314 864087
rect 675478 864035 675530 864087
rect 674230 863147 674282 863199
rect 680086 863147 680138 863199
rect 674422 863073 674474 863125
rect 679990 863073 680042 863125
rect 675190 862407 675242 862459
rect 675382 862407 675434 862459
rect 674902 861963 674954 862015
rect 675382 861963 675434 862015
rect 674614 861815 674666 861867
rect 674902 861815 674954 861867
rect 656374 861223 656426 861275
rect 674614 861223 674666 861275
rect 654838 861149 654890 861201
rect 675190 861149 675242 861201
rect 674998 859521 675050 859573
rect 675478 859521 675530 859573
rect 674902 858707 674954 858759
rect 675382 858707 675434 858759
rect 674038 858263 674090 858315
rect 674998 858263 675050 858315
rect 674230 858115 674282 858167
rect 675478 858115 675530 858167
rect 674422 857671 674474 857723
rect 675382 857671 675434 857723
rect 674998 855155 675050 855207
rect 675382 855155 675434 855207
rect 675094 854489 675146 854541
rect 675382 854489 675434 854541
rect 674902 853971 674954 854023
rect 675382 853971 675434 854023
rect 674518 853157 674570 853209
rect 675478 853157 675530 853209
rect 675190 852713 675242 852765
rect 675382 852713 675434 852765
rect 674134 852121 674186 852173
rect 675382 852121 675434 852173
rect 674614 850863 674666 850915
rect 675382 850863 675434 850915
rect 674326 850123 674378 850175
rect 675478 850123 675530 850175
rect 675190 848421 675242 848473
rect 675478 848421 675530 848473
rect 41782 817933 41834 817985
rect 47542 817933 47594 817985
rect 41782 817267 41834 817319
rect 44758 817267 44810 817319
rect 41590 816527 41642 816579
rect 44854 816527 44906 816579
rect 41782 815787 41834 815839
rect 43222 815787 43274 815839
rect 41782 814825 41834 814877
rect 44662 814825 44714 814877
rect 41590 813567 41642 813619
rect 44566 813567 44618 813619
rect 41878 808757 41930 808809
rect 42742 808757 42794 808809
rect 41878 807055 41930 807107
rect 43030 807055 43082 807107
rect 41398 806981 41450 807033
rect 43126 806981 43178 807033
rect 41590 806759 41642 806811
rect 42838 806759 42890 806811
rect 41590 806463 41642 806515
rect 42934 806463 42986 806515
rect 37366 806315 37418 806367
rect 42646 806315 42698 806367
rect 41590 805131 41642 805183
rect 47446 805131 47498 805183
rect 34390 804909 34442 804961
rect 41878 804909 41930 804961
rect 40150 801357 40202 801409
rect 43414 801357 43466 801409
rect 40246 801283 40298 801335
rect 43318 801283 43370 801335
rect 41974 801061 42026 801113
rect 43510 801061 43562 801113
rect 41782 800987 41834 801039
rect 42070 800987 42122 801039
rect 41782 800765 41834 800817
rect 43030 800765 43082 800817
rect 43606 800765 43658 800817
rect 42646 800617 42698 800669
rect 43030 800617 43082 800669
rect 57622 800617 57674 800669
rect 43126 800543 43178 800595
rect 43414 800469 43466 800521
rect 43318 799211 43370 799263
rect 43606 799211 43658 799263
rect 42166 798915 42218 798967
rect 42646 798915 42698 798967
rect 42166 797879 42218 797931
rect 43318 797879 43370 797931
rect 42166 797065 42218 797117
rect 42742 797065 42794 797117
rect 42742 796917 42794 796969
rect 43510 796917 43562 796969
rect 42070 796251 42122 796303
rect 43030 796251 43082 796303
rect 43030 796103 43082 796155
rect 43414 796103 43466 796155
rect 42166 795659 42218 795711
rect 42934 795659 42986 795711
rect 42646 795511 42698 795563
rect 42934 795511 42986 795563
rect 42166 795215 42218 795267
rect 42838 795215 42890 795267
rect 42838 795067 42890 795119
rect 43606 795067 43658 795119
rect 42646 794919 42698 794971
rect 43702 794919 43754 794971
rect 42070 794475 42122 794527
rect 43030 794475 43082 794527
rect 42166 793735 42218 793787
rect 42742 793735 42794 793787
rect 42646 792107 42698 792159
rect 42838 792107 42890 792159
rect 42550 791885 42602 791937
rect 42646 791811 42698 791863
rect 42070 791441 42122 791493
rect 42550 791441 42602 791493
rect 42166 790775 42218 790827
rect 42646 790775 42698 790827
rect 43318 789739 43370 789791
rect 58006 789739 58058 789791
rect 42070 789591 42122 789643
rect 43126 789591 43178 789643
rect 42646 789147 42698 789199
rect 58198 789147 58250 789199
rect 44854 789073 44906 789125
rect 58390 789073 58442 789125
rect 42262 787815 42314 787867
rect 43030 787815 43082 787867
rect 42166 787223 42218 787275
rect 42934 787223 42986 787275
rect 42166 785891 42218 785943
rect 42646 785891 42698 785943
rect 44758 785595 44810 785647
rect 58678 785595 58730 785647
rect 47542 785225 47594 785277
rect 59638 785225 59690 785277
rect 654166 774717 654218 774769
rect 675382 774791 675434 774843
rect 41782 774643 41834 774695
rect 47638 774643 47690 774695
rect 41590 773903 41642 773955
rect 44758 773903 44810 773955
rect 41782 773459 41834 773511
rect 44950 773459 45002 773511
rect 41590 773385 41642 773437
rect 43222 773385 43274 773437
rect 41782 772571 41834 772623
rect 43222 772571 43274 772623
rect 41590 772127 41642 772179
rect 62038 772127 62090 772179
rect 43126 771905 43178 771957
rect 61846 771905 61898 771957
rect 654838 771905 654890 771957
rect 674998 771905 675050 771957
rect 656182 771831 656234 771883
rect 675094 771831 675146 771883
rect 674230 771313 674282 771365
rect 675382 771313 675434 771365
rect 41782 769611 41834 769663
rect 43126 769611 43178 769663
rect 674422 766799 674474 766851
rect 675382 766799 675434 766851
rect 674134 766281 674186 766333
rect 675478 766281 675530 766333
rect 674326 765689 674378 765741
rect 675478 765689 675530 765741
rect 675094 765245 675146 765297
rect 675382 765245 675434 765297
rect 41782 765097 41834 765149
rect 42742 765097 42794 765149
rect 674518 765097 674570 765149
rect 675478 765097 675530 765149
rect 674902 763691 674954 763743
rect 675382 763691 675434 763743
rect 41590 763543 41642 763595
rect 42934 763543 42986 763595
rect 674998 763469 675050 763521
rect 675382 763469 675434 763521
rect 41590 763395 41642 763447
rect 42838 763395 42890 763447
rect 41782 762063 41834 762115
rect 47542 762063 47594 762115
rect 674998 761841 675050 761893
rect 675382 761841 675434 761893
rect 40246 760287 40298 760339
rect 41014 760287 41066 760339
rect 674902 760287 674954 760339
rect 675382 760287 675434 760339
rect 37366 760213 37418 760265
rect 41782 760213 41834 760265
rect 40150 758067 40202 758119
rect 43606 758067 43658 758119
rect 42262 757919 42314 757971
rect 43510 757919 43562 757971
rect 41974 757845 42026 757897
rect 43414 757845 43466 757897
rect 41878 757771 41930 757823
rect 42166 757771 42218 757823
rect 43318 757771 43370 757823
rect 41878 757549 41930 757601
rect 42742 756365 42794 756417
rect 42358 756143 42410 756195
rect 42166 755699 42218 755751
rect 43126 755699 43178 755751
rect 43126 755551 43178 755603
rect 43318 755551 43370 755603
rect 42070 754663 42122 754715
rect 43318 754663 43370 754715
rect 42166 753849 42218 753901
rect 42934 753849 42986 753901
rect 42934 753701 42986 753753
rect 43414 753701 43466 753753
rect 42166 752591 42218 752643
rect 42838 752591 42890 752643
rect 42070 752369 42122 752421
rect 43414 752369 43466 752421
rect 42070 751851 42122 751903
rect 42358 751999 42410 752051
rect 42358 751851 42410 751903
rect 43126 751851 43178 751903
rect 43030 751777 43082 751829
rect 43510 751777 43562 751829
rect 42838 751629 42890 751681
rect 43126 751629 43178 751681
rect 42358 751555 42410 751607
rect 42838 751481 42890 751533
rect 42166 751259 42218 751311
rect 42934 751259 42986 751311
rect 42166 750519 42218 750571
rect 43030 750519 43082 750571
rect 43318 748743 43370 748795
rect 57910 748743 57962 748795
rect 42166 748151 42218 748203
rect 42838 748151 42890 748203
rect 42166 747559 42218 747611
rect 43606 747559 43658 747611
rect 42166 746227 42218 746279
rect 42934 746227 42986 746279
rect 42358 746079 42410 746131
rect 44854 746079 44906 746131
rect 42358 745931 42410 745983
rect 54646 745931 54698 745983
rect 54742 745931 54794 745983
rect 57622 745931 57674 745983
rect 44950 745339 45002 745391
rect 59254 745339 59306 745391
rect 43414 745265 43466 745317
rect 59638 745265 59690 745317
rect 42166 744599 42218 744651
rect 43030 744599 43082 744651
rect 42166 744007 42218 744059
rect 43126 744007 43178 744059
rect 42070 743341 42122 743393
rect 42838 743341 42890 743393
rect 47638 742971 47690 743023
rect 59638 742971 59690 743023
rect 44758 742897 44810 742949
rect 59734 742897 59786 742949
rect 42166 742749 42218 742801
rect 42358 742749 42410 742801
rect 41782 731427 41834 731479
rect 50326 731427 50378 731479
rect 41590 730687 41642 730739
rect 47734 730687 47786 730739
rect 41782 730317 41834 730369
rect 44758 730317 44810 730369
rect 41590 730169 41642 730221
rect 43222 730169 43274 730221
rect 41590 729207 41642 729259
rect 43702 729207 43754 729259
rect 41206 728837 41258 728889
rect 62230 728837 62282 728889
rect 40438 728763 40490 728815
rect 62422 728763 62474 728815
rect 654166 728689 654218 728741
rect 675286 728689 675338 728741
rect 41590 728615 41642 728667
rect 43510 728615 43562 728667
rect 41782 727875 41834 727927
rect 43414 727875 43466 727927
rect 654262 727135 654314 727187
rect 674614 727135 674666 727187
rect 41782 726099 41834 726151
rect 42934 726099 42986 726151
rect 673270 724915 673322 724967
rect 675478 724915 675530 724967
rect 654166 724323 654218 724375
rect 673942 724323 673994 724375
rect 673942 723361 673994 723413
rect 675286 723361 675338 723413
rect 674518 722399 674570 722451
rect 675382 722399 675434 722451
rect 41590 721363 41642 721415
rect 43126 721363 43178 721415
rect 674038 721141 674090 721193
rect 675478 721141 675530 721193
rect 674614 720845 674666 720897
rect 675382 720845 675434 720897
rect 672886 720697 672938 720749
rect 675478 720697 675530 720749
rect 41590 720401 41642 720453
rect 42838 720401 42890 720453
rect 41590 720179 41642 720231
rect 43030 720179 43082 720231
rect 674518 719291 674570 719343
rect 675382 719291 675434 719343
rect 41590 718699 41642 718751
rect 47638 718699 47690 718751
rect 675286 715591 675338 715643
rect 675382 715591 675434 715643
rect 675382 715369 675434 715421
rect 675574 715295 675626 715347
rect 41974 714629 42026 714681
rect 43318 714629 43370 714681
rect 41782 714555 41834 714607
rect 41878 714555 41930 714607
rect 43606 714555 43658 714607
rect 41782 714333 41834 714385
rect 42262 714259 42314 714311
rect 43222 714259 43274 714311
rect 673366 714185 673418 714237
rect 679702 714185 679754 714237
rect 42838 712853 42890 712905
rect 43126 712853 43178 712905
rect 43222 712557 43274 712609
rect 43510 712557 43562 712609
rect 42070 712483 42122 712535
rect 42934 712483 42986 712535
rect 42934 712335 42986 712387
rect 43318 712335 43370 712387
rect 43318 712187 43370 712239
rect 43702 712187 43754 712239
rect 42166 711225 42218 711277
rect 43702 711225 43754 711277
rect 42070 710633 42122 710685
rect 42838 710633 42890 710685
rect 42838 710485 42890 710537
rect 43606 710485 43658 710537
rect 674038 709893 674090 709945
rect 675670 709893 675722 709945
rect 42166 709597 42218 709649
rect 43510 709597 43562 709649
rect 42070 709375 42122 709427
rect 43030 709375 43082 709427
rect 43030 708783 43082 708835
rect 42166 708635 42218 708687
rect 42838 708635 42890 708687
rect 42166 708191 42218 708243
rect 42742 708191 42794 708243
rect 42742 708043 42794 708095
rect 42070 707229 42122 707281
rect 42934 707229 42986 707281
rect 42358 705527 42410 705579
rect 42742 705527 42794 705579
rect 42166 705083 42218 705135
rect 42358 705083 42410 705135
rect 43702 704861 43754 704913
rect 58390 704861 58442 704913
rect 42166 704491 42218 704543
rect 42838 704491 42890 704543
rect 42070 703751 42122 703803
rect 43126 703751 43178 703803
rect 42166 703233 42218 703285
rect 43030 703233 43082 703285
rect 655606 703011 655658 703063
rect 676246 703011 676298 703063
rect 655222 702863 655274 702915
rect 676246 702863 676298 702915
rect 43510 702641 43562 702693
rect 58774 702641 58826 702693
rect 44758 702567 44810 702619
rect 58678 702567 58730 702619
rect 42070 700791 42122 700843
rect 42934 700791 42986 700843
rect 669526 700791 669578 700843
rect 670870 700791 670922 700843
rect 676246 700791 676298 700843
rect 42166 700199 42218 700251
rect 42742 700199 42794 700251
rect 670678 700051 670730 700103
rect 676246 700051 676298 700103
rect 655414 699829 655466 699881
rect 676054 699829 676106 699881
rect 50326 699755 50378 699807
rect 59254 699755 59306 699807
rect 47734 699681 47786 699733
rect 58870 699681 58922 699733
rect 670966 699681 671018 699733
rect 676054 699681 676106 699733
rect 42070 699533 42122 699585
rect 42838 699533 42890 699585
rect 674230 699163 674282 699215
rect 676246 699163 676298 699215
rect 670870 699089 670922 699141
rect 676054 699089 676106 699141
rect 674998 698941 675050 698993
rect 676054 698941 676106 698993
rect 669718 696943 669770 696995
rect 670966 696943 671018 696995
rect 674902 696869 674954 696921
rect 676054 696869 676106 696921
rect 674422 696795 674474 696847
rect 675958 696795 676010 696847
rect 674902 696647 674954 696699
rect 676246 696647 676298 696699
rect 674326 693983 674378 694035
rect 676054 693983 676106 694035
rect 674134 693613 674186 693665
rect 676054 693613 676106 693665
rect 670774 691171 670826 691223
rect 679702 691171 679754 691223
rect 674326 689765 674378 689817
rect 675670 689765 675722 689817
rect 674998 689395 675050 689447
rect 675574 689395 675626 689447
rect 649462 688359 649514 688411
rect 679990 688359 680042 688411
rect 41782 688211 41834 688263
rect 53206 688211 53258 688263
rect 41590 687471 41642 687523
rect 50326 687471 50378 687523
rect 41782 687175 41834 687227
rect 47830 687175 47882 687227
rect 41590 686953 41642 687005
rect 43318 686953 43370 687005
rect 674038 686213 674090 686265
rect 675382 686213 675434 686265
rect 41590 685991 41642 686043
rect 43510 685991 43562 686043
rect 656374 685547 656426 685599
rect 674038 685547 674090 685599
rect 41782 685325 41834 685377
rect 43222 685325 43274 685377
rect 44758 685325 44810 685377
rect 672406 685325 672458 685377
rect 675478 685325 675530 685377
rect 41590 684511 41642 684563
rect 43318 684511 43370 684563
rect 41782 684141 41834 684193
rect 43414 684141 43466 684193
rect 44950 684141 45002 684193
rect 41782 682735 41834 682787
rect 43126 682735 43178 682787
rect 672694 682069 672746 682121
rect 675478 682069 675530 682121
rect 672982 681255 673034 681307
rect 675382 681255 675434 681307
rect 655990 681181 656042 681233
rect 674902 681181 674954 681233
rect 654454 681107 654506 681159
rect 674422 681107 674474 681159
rect 672214 680737 672266 680789
rect 675382 680737 675434 680789
rect 674902 679627 674954 679679
rect 675286 679627 675338 679679
rect 675190 679035 675242 679087
rect 674998 678813 675050 678865
rect 673078 677555 673130 677607
rect 675382 677555 675434 677607
rect 41590 677259 41642 677311
rect 42934 677259 42986 677311
rect 41782 677185 41834 677237
rect 42838 677185 42890 677237
rect 672502 677037 672554 677089
rect 675478 677037 675530 677089
rect 673174 676667 673226 676719
rect 675478 676667 675530 676719
rect 674422 676149 674474 676201
rect 675286 676149 675338 676201
rect 41782 675705 41834 675757
rect 47734 675705 47786 675757
rect 672310 675113 672362 675165
rect 675478 675113 675530 675165
rect 42742 671043 42794 671095
rect 59638 671043 59690 671095
rect 42262 670747 42314 670799
rect 42166 670525 42218 670577
rect 674902 669637 674954 669689
rect 675574 669637 675626 669689
rect 674998 669563 675050 669615
rect 675478 669563 675530 669615
rect 42166 669119 42218 669171
rect 43126 669119 43178 669171
rect 42838 668527 42890 668579
rect 43126 668527 43178 668579
rect 42166 668453 42218 668505
rect 42742 668453 42794 668505
rect 42166 667269 42218 667321
rect 43030 667269 43082 667321
rect 42070 665863 42122 665915
rect 43126 665863 43178 665915
rect 42166 665641 42218 665693
rect 43222 665641 43274 665693
rect 42166 665419 42218 665471
rect 42742 665419 42794 665471
rect 42070 664605 42122 664657
rect 42934 664605 42986 664657
rect 42166 664161 42218 664213
rect 42838 664161 42890 664213
rect 42070 661645 42122 661697
rect 43030 661645 43082 661697
rect 42166 661127 42218 661179
rect 42742 661127 42794 661179
rect 42166 660239 42218 660291
rect 43126 660239 43178 660291
rect 42070 659647 42122 659699
rect 42358 659647 42410 659699
rect 47830 659425 47882 659477
rect 59158 659425 59210 659477
rect 43222 659351 43274 659403
rect 58774 659351 58826 659403
rect 42166 657945 42218 657997
rect 42934 657945 42986 657997
rect 670774 657575 670826 657627
rect 676054 657575 676106 657627
rect 42166 657427 42218 657479
rect 42838 657427 42890 657479
rect 655510 657131 655562 657183
rect 676150 657131 676202 657183
rect 655318 656983 655370 657035
rect 676246 656983 676298 657035
rect 673750 656909 673802 656961
rect 676054 656909 676106 656961
rect 655126 656835 655178 656887
rect 676342 656835 676394 656887
rect 42166 656761 42218 656813
rect 43030 656761 43082 656813
rect 53206 656613 53258 656665
rect 58198 656613 58250 656665
rect 50326 656539 50378 656591
rect 58390 656539 58442 656591
rect 670678 656465 670730 656517
rect 676054 656465 676106 656517
rect 42166 656095 42218 656147
rect 45046 656095 45098 656147
rect 670870 656021 670922 656073
rect 676054 656021 676106 656073
rect 670966 655725 671018 655777
rect 676246 655725 676298 655777
rect 652246 655281 652298 655333
rect 670966 655281 671018 655333
rect 649750 655207 649802 655259
rect 670678 655207 670730 655259
rect 670774 654763 670826 654815
rect 676246 654763 676298 654815
rect 674614 653727 674666 653779
rect 676054 653727 676106 653779
rect 674518 650841 674570 650893
rect 676054 650841 676106 650893
rect 673270 649213 673322 649265
rect 676246 649213 676298 649265
rect 672886 648029 672938 648081
rect 676054 648029 676106 648081
rect 649558 645143 649610 645195
rect 679798 645143 679850 645195
rect 41590 644847 41642 644899
rect 53206 644847 53258 644899
rect 41590 644255 41642 644307
rect 50326 644255 50378 644307
rect 41782 643959 41834 644011
rect 47926 643959 47978 644011
rect 41590 643737 41642 643789
rect 43510 643737 43562 643789
rect 41590 642775 41642 642827
rect 43222 642775 43274 642827
rect 43126 642479 43178 642531
rect 61942 642479 61994 642531
rect 43414 642257 43466 642309
rect 45142 642257 45194 642309
rect 654166 642183 654218 642235
rect 675190 642183 675242 642235
rect 41590 641295 41642 641347
rect 43318 641295 43370 641347
rect 41590 639667 41642 639719
rect 43030 639667 43082 639719
rect 670966 637817 671018 637869
rect 675382 637817 675434 637869
rect 673366 637077 673418 637129
rect 675478 637077 675530 637129
rect 655798 636633 655850 636685
rect 675190 636633 675242 636685
rect 673270 636485 673322 636537
rect 675382 636485 675434 636537
rect 655894 635005 655946 635057
rect 674998 635005 675050 635057
rect 41782 634191 41834 634243
rect 43126 634191 43178 634243
rect 41782 633895 41834 633947
rect 42934 633895 42986 633947
rect 672790 633599 672842 633651
rect 675382 633599 675434 633651
rect 41782 632489 41834 632541
rect 47830 632489 47882 632541
rect 672886 632341 672938 632393
rect 675478 632341 675530 632393
rect 672598 630713 672650 630765
rect 675286 630713 675338 630765
rect 674998 630639 675050 630691
rect 675478 630639 675530 630691
rect 41878 627975 41930 628027
rect 42838 627827 42890 627879
rect 54646 627827 54698 627879
rect 41878 627753 41930 627805
rect 43126 626643 43178 626695
rect 42934 626495 42986 626547
rect 43126 626495 43178 626547
rect 42166 625903 42218 625955
rect 43030 625903 43082 625955
rect 43030 625755 43082 625807
rect 42070 625237 42122 625289
rect 42838 625237 42890 625289
rect 54646 624793 54698 624845
rect 58966 624793 59018 624845
rect 42166 624053 42218 624105
rect 43030 624053 43082 624105
rect 42070 622647 42122 622699
rect 43126 622647 43178 622699
rect 42166 622499 42218 622551
rect 43414 622499 43466 622551
rect 42070 622203 42122 622255
rect 42838 622203 42890 622255
rect 42166 621463 42218 621515
rect 42934 621463 42986 621515
rect 42166 618429 42218 618481
rect 42838 618429 42890 618481
rect 42166 617763 42218 617815
rect 43030 617763 43082 617815
rect 42838 616357 42890 616409
rect 58198 616357 58250 616409
rect 47926 616283 47978 616335
rect 58966 616283 59018 616335
rect 43414 616209 43466 616261
rect 59638 616209 59690 616261
rect 42166 614803 42218 614855
rect 42934 614803 42986 614855
rect 42166 614211 42218 614263
rect 43126 614211 43178 614263
rect 655606 613915 655658 613967
rect 676246 613915 676298 613967
rect 655414 613767 655466 613819
rect 676150 613767 676202 613819
rect 655222 613619 655274 613671
rect 676054 613619 676106 613671
rect 42070 613471 42122 613523
rect 43030 613471 43082 613523
rect 53206 613397 53258 613449
rect 59638 613397 59690 613449
rect 50326 613323 50378 613375
rect 59542 613323 59594 613375
rect 673750 613175 673802 613227
rect 676054 613175 676106 613227
rect 42166 612953 42218 613005
rect 42838 612953 42890 613005
rect 672118 612583 672170 612635
rect 676054 612583 676106 612635
rect 669814 611843 669866 611895
rect 670870 611843 670922 611895
rect 676246 611843 676298 611895
rect 670582 611621 670634 611673
rect 676054 611621 676106 611673
rect 669622 611103 669674 611155
rect 670774 611103 670826 611155
rect 676054 611103 676106 611155
rect 670678 610585 670730 610637
rect 676054 610585 676106 610637
rect 672406 607181 672458 607233
rect 676054 607181 676106 607233
rect 672694 606663 672746 606715
rect 676054 606663 676106 606715
rect 672982 606293 673034 606345
rect 676246 606293 676298 606345
rect 672310 605701 672362 605753
rect 676054 605701 676106 605753
rect 672502 605109 672554 605161
rect 676054 605109 676106 605161
rect 672214 604665 672266 604717
rect 676054 604665 676106 604717
rect 673078 604369 673130 604421
rect 676246 604369 676298 604421
rect 673174 603629 673226 603681
rect 676054 603629 676106 603681
rect 654550 602001 654602 602053
rect 675382 602001 675434 602053
rect 649654 601927 649706 601979
rect 679990 601927 680042 601979
rect 41782 601335 41834 601387
rect 53206 601335 53258 601387
rect 41782 600743 41834 600795
rect 50326 600743 50378 600795
rect 43318 600447 43370 600499
rect 62326 600447 62378 600499
rect 41782 600373 41834 600425
rect 43222 600373 43274 600425
rect 41782 599781 41834 599833
rect 43222 599781 43274 599833
rect 39766 599411 39818 599463
rect 43318 599411 43370 599463
rect 41782 599263 41834 599315
rect 43318 599263 43370 599315
rect 40342 599189 40394 599241
rect 62134 599189 62186 599241
rect 41590 599041 41642 599093
rect 56182 599041 56234 599093
rect 41782 598301 41834 598353
rect 46102 598301 46154 598353
rect 41590 596599 41642 596651
rect 43126 596599 43178 596651
rect 674902 596303 674954 596355
rect 675382 596303 675434 596355
rect 654166 593343 654218 593395
rect 674902 593343 674954 593395
rect 673654 593269 673706 593321
rect 675382 593269 675434 593321
rect 672982 592677 673034 592729
rect 675478 592677 675530 592729
rect 672310 592085 672362 592137
rect 675382 592085 675434 592137
rect 41782 590975 41834 591027
rect 43030 590975 43082 591027
rect 41782 590827 41834 590879
rect 42934 590827 42986 590879
rect 654358 590457 654410 590509
rect 674998 590457 675050 590509
rect 673174 588977 673226 589029
rect 675382 588977 675434 589029
rect 672214 588533 672266 588585
rect 675382 588533 675434 588585
rect 674902 588089 674954 588141
rect 675382 588089 675434 588141
rect 673078 587941 673130 587993
rect 675478 587941 675530 587993
rect 41590 587497 41642 587549
rect 56086 587497 56138 587549
rect 672694 586461 672746 586513
rect 675382 586461 675434 586513
rect 674998 586239 675050 586291
rect 675478 586239 675530 586291
rect 41878 584759 41930 584811
rect 42838 584685 42890 584737
rect 58966 584685 59018 584737
rect 41878 584537 41930 584589
rect 42070 582687 42122 582739
rect 43126 582687 43178 582739
rect 42070 582021 42122 582073
rect 42838 582021 42890 582073
rect 42070 580837 42122 580889
rect 43030 580837 43082 580889
rect 42166 579579 42218 579631
rect 42934 579579 42986 579631
rect 42070 579431 42122 579483
rect 47926 579431 47978 579483
rect 42070 578987 42122 579039
rect 42454 578987 42506 579039
rect 672118 578913 672170 578965
rect 679702 578913 679754 578965
rect 42166 578247 42218 578299
rect 43030 578247 43082 578299
rect 42070 577507 42122 577559
rect 42934 577507 42986 577559
rect 42166 575213 42218 575265
rect 42454 575213 42506 575265
rect 42166 574695 42218 574747
rect 43126 574695 43178 574747
rect 42070 574029 42122 574081
rect 42838 574029 42890 574081
rect 42358 573289 42410 573341
rect 42166 573215 42218 573267
rect 50326 573067 50378 573119
rect 58966 573067 59018 573119
rect 47926 572993 47978 573045
rect 59638 572993 59690 573045
rect 42070 570995 42122 571047
rect 42934 570995 42986 571047
rect 42166 570921 42218 570973
rect 43030 570921 43082 570973
rect 42166 570255 42218 570307
rect 42838 570255 42890 570307
rect 56182 570181 56234 570233
rect 60406 570181 60458 570233
rect 53206 570107 53258 570159
rect 59158 570107 59210 570159
rect 42166 569737 42218 569789
rect 45046 569737 45098 569789
rect 655510 567887 655562 567939
rect 676054 567887 676106 567939
rect 655318 567739 655370 567791
rect 676246 567739 676298 567791
rect 670870 567443 670922 567495
rect 676054 567443 676106 567495
rect 655126 567369 655178 567421
rect 676150 567369 676202 567421
rect 670102 567073 670154 567125
rect 670582 567073 670634 567125
rect 676246 567073 676298 567125
rect 672406 566259 672458 566311
rect 676246 566259 676298 566311
rect 669910 565889 669962 565941
rect 670678 565889 670730 565941
rect 676054 565889 676106 565941
rect 672502 565371 672554 565423
rect 676054 565371 676106 565423
rect 670966 561449 671018 561501
rect 676054 561449 676106 561501
rect 673366 560857 673418 560909
rect 676054 560857 676106 560909
rect 672598 560709 672650 560761
rect 676246 560709 676298 560761
rect 673270 559377 673322 559429
rect 676054 559377 676106 559429
rect 672790 559007 672842 559059
rect 676054 559007 676106 559059
rect 672886 558637 672938 558689
rect 676246 558637 676298 558689
rect 649846 555825 649898 555877
rect 679798 555825 679850 555877
rect 653782 552865 653834 552917
rect 675286 552865 675338 552917
rect 672886 549091 672938 549143
rect 675286 549091 675338 549143
rect 673366 547907 673418 547959
rect 675478 547907 675530 547959
rect 654166 547389 654218 547441
rect 674902 547389 674954 547441
rect 656278 547315 656330 547367
rect 674998 547315 675050 547367
rect 673270 547241 673322 547293
rect 675286 547241 675338 547293
rect 672790 544873 672842 544925
rect 675478 544873 675530 544925
rect 674998 543911 675050 543963
rect 675382 543911 675434 543963
rect 673846 543689 673898 543741
rect 675478 543689 675530 543741
rect 675190 542283 675242 542335
rect 675382 542283 675434 542335
rect 674902 542061 674954 542113
rect 675382 542061 675434 542113
rect 42934 541543 42986 541595
rect 57718 541543 57770 541595
rect 42838 541469 42890 541521
rect 57622 541469 57674 541521
rect 673942 538583 673994 538635
rect 675478 538583 675530 538635
rect 42166 538435 42218 538487
rect 42934 538435 42986 538487
rect 42166 537029 42218 537081
rect 42838 537029 42890 537081
rect 42166 535697 42218 535749
rect 43414 535697 43466 535749
rect 42070 526373 42122 526425
rect 45046 526373 45098 526425
rect 655606 524523 655658 524575
rect 676246 524523 676298 524575
rect 655414 524375 655466 524427
rect 676342 524375 676394 524427
rect 50326 524301 50378 524353
rect 58582 524301 58634 524353
rect 47926 524227 47978 524279
rect 59350 524227 59402 524279
rect 655222 524153 655274 524205
rect 676150 524153 676202 524205
rect 670870 524005 670922 524057
rect 676054 524005 676106 524057
rect 672406 523857 672458 523909
rect 676054 523857 676106 523909
rect 672502 521193 672554 521245
rect 676246 521193 676298 521245
rect 673654 517641 673706 517693
rect 676246 517641 676298 517693
rect 672982 516901 673034 516953
rect 676054 516901 676106 516953
rect 672694 516457 672746 516509
rect 676054 516457 676106 516509
rect 672214 516161 672266 516213
rect 676246 516161 676298 516213
rect 672310 515421 672362 515473
rect 676054 515421 676106 515473
rect 673174 514977 673226 515029
rect 676054 514977 676106 515029
rect 673078 514459 673130 514511
rect 676054 514459 676106 514511
rect 649942 512683 649994 512735
rect 679990 512683 680042 512735
rect 676438 485303 676490 485355
rect 676630 485303 676682 485355
rect 655510 481307 655562 481359
rect 676246 481307 676298 481359
rect 655318 481159 655370 481211
rect 676342 481159 676394 481211
rect 655126 480937 655178 480989
rect 676150 480937 676202 480989
rect 670006 479383 670058 479435
rect 676438 479383 676490 479435
rect 670294 479087 670346 479139
rect 676630 479087 676682 479139
rect 675286 478643 675338 478695
rect 676054 478643 676106 478695
rect 673654 478347 673706 478399
rect 676246 478347 676298 478399
rect 673942 476793 673994 476845
rect 676054 476793 676106 476845
rect 41782 476053 41834 476105
rect 50326 476053 50378 476105
rect 41782 475535 41834 475587
rect 47926 475535 47978 475587
rect 672886 474647 672938 474699
rect 676054 474647 676106 474699
rect 41878 474573 41930 474625
rect 43222 474573 43274 474625
rect 673270 474277 673322 474329
rect 676246 474277 676298 474329
rect 673366 472797 673418 472849
rect 676246 472797 676298 472849
rect 41782 472353 41834 472405
rect 58966 472353 59018 472405
rect 672790 472205 672842 472257
rect 676054 472205 676106 472257
rect 41782 471983 41834 472035
rect 46006 471983 46058 472035
rect 673846 471613 673898 471665
rect 676054 471613 676106 471665
rect 650038 469467 650090 469519
rect 679798 469467 679850 469519
rect 41590 465249 41642 465301
rect 43414 465249 43466 465301
rect 41782 463547 41834 463599
rect 47926 463547 47978 463599
rect 34486 463103 34538 463155
rect 41782 463103 41834 463155
rect 673654 440607 673706 440659
rect 675382 440607 675434 440659
rect 41686 432023 41738 432075
rect 62518 432023 62570 432075
rect 41782 429211 41834 429263
rect 53206 429211 53258 429263
rect 673846 429137 673898 429189
rect 675286 429137 675338 429189
rect 41590 428471 41642 428523
rect 50326 428471 50378 428523
rect 41782 428175 41834 428227
rect 48118 428175 48170 428227
rect 41590 426991 41642 427043
rect 43318 426991 43370 427043
rect 41782 426621 41834 426673
rect 43222 426621 43274 426673
rect 39670 426251 39722 426303
rect 41686 426251 41738 426303
rect 41590 420405 41642 420457
rect 43414 420405 43466 420457
rect 41590 417815 41642 417867
rect 42838 417815 42890 417867
rect 41590 416483 41642 416535
rect 48022 416483 48074 416535
rect 41686 414633 41738 414685
rect 45334 414633 45386 414685
rect 41782 413819 41834 413871
rect 41782 413523 41834 413575
rect 42070 410119 42122 410171
rect 42742 410119 42794 410171
rect 42166 409823 42218 409875
rect 42838 409823 42890 409875
rect 42070 408269 42122 408321
rect 42838 408269 42890 408321
rect 42742 406049 42794 406101
rect 58486 406049 58538 406101
rect 42838 402793 42890 402845
rect 59638 402793 59690 402845
rect 53206 400277 53258 400329
rect 59734 400277 59786 400329
rect 50326 400203 50378 400255
rect 59542 400203 59594 400255
rect 48118 400129 48170 400181
rect 59638 400129 59690 400181
rect 655510 394727 655562 394779
rect 676150 394727 676202 394779
rect 655318 394653 655370 394705
rect 676246 394653 676298 394705
rect 655126 394579 655178 394631
rect 676342 394579 676394 394631
rect 42166 394505 42218 394557
rect 57622 394505 57674 394557
rect 672598 393839 672650 393891
rect 673846 393839 673898 393891
rect 676246 393839 676298 393891
rect 675382 393173 675434 393225
rect 675862 393173 675914 393225
rect 675190 391693 675242 391745
rect 676246 391693 676298 391745
rect 674038 389695 674090 389747
rect 676054 389695 676106 389747
rect 674614 389103 674666 389155
rect 676246 389103 676298 389155
rect 674902 388881 674954 388933
rect 676054 388881 676106 388933
rect 675286 388807 675338 388859
rect 676246 388807 676298 388859
rect 674134 387031 674186 387083
rect 676246 387031 676298 387083
rect 674518 386735 674570 386787
rect 676054 386735 676106 386787
rect 674422 386291 674474 386343
rect 675958 386291 676010 386343
rect 674230 386069 674282 386121
rect 676246 386069 676298 386121
rect 41782 385995 41834 386047
rect 53206 385995 53258 386047
rect 674710 385995 674762 386047
rect 675958 385995 676010 386047
rect 674806 385921 674858 385973
rect 676054 385921 676106 385973
rect 41590 385255 41642 385307
rect 50326 385255 50378 385307
rect 41782 384959 41834 385011
rect 48214 384959 48266 385011
rect 41590 384737 41642 384789
rect 43318 384737 43370 384789
rect 41590 383775 41642 383827
rect 43318 383775 43370 383827
rect 41782 383479 41834 383531
rect 43510 383479 43562 383531
rect 41590 383257 41642 383309
rect 43222 383257 43274 383309
rect 45238 383257 45290 383309
rect 674326 383109 674378 383161
rect 676246 383109 676298 383161
rect 650134 383035 650186 383087
rect 679702 383035 679754 383087
rect 666646 382961 666698 383013
rect 675862 382961 675914 383013
rect 41782 381999 41834 382051
rect 43414 381999 43466 382051
rect 45430 381999 45482 382051
rect 674998 379409 675050 379461
rect 675478 379409 675530 379461
rect 39958 377189 40010 377241
rect 43414 377189 43466 377241
rect 674614 376523 674666 376575
rect 675478 376523 675530 376575
rect 674518 375635 674570 375687
rect 675382 375635 675434 375687
rect 674422 375191 674474 375243
rect 675478 375191 675530 375243
rect 674806 374673 674858 374725
rect 675382 374673 675434 374725
rect 41590 374451 41642 374503
rect 42838 374451 42890 374503
rect 41590 373267 41642 373319
rect 48118 373267 48170 373319
rect 674038 372157 674090 372209
rect 675382 372157 675434 372209
rect 654166 371491 654218 371543
rect 674998 371491 675050 371543
rect 674710 371417 674762 371469
rect 675382 371417 675434 371469
rect 674230 370973 674282 371025
rect 675382 370973 675434 371025
rect 41782 370603 41834 370655
rect 41782 370307 41834 370359
rect 674326 370307 674378 370359
rect 675478 370307 675530 370359
rect 674134 369123 674186 369175
rect 675382 369123 675434 369175
rect 42070 366903 42122 366955
rect 42742 366903 42794 366955
rect 42166 366681 42218 366733
rect 42838 366681 42890 366733
rect 674902 365423 674954 365475
rect 675478 365423 675530 365475
rect 42166 365053 42218 365105
rect 42838 365053 42890 365105
rect 42742 362537 42794 362589
rect 58294 362537 58346 362589
rect 660310 360835 660362 360887
rect 666646 360835 666698 360887
rect 42838 359947 42890 359999
rect 59158 359947 59210 359999
rect 53206 357061 53258 357113
rect 58198 357061 58250 357113
rect 48214 356987 48266 357039
rect 59638 356987 59690 357039
rect 50326 356913 50378 356965
rect 58582 356913 58634 356965
rect 655222 351585 655274 351637
rect 676054 351585 676106 351637
rect 655126 351511 655178 351563
rect 676246 351511 676298 351563
rect 655414 351363 655466 351415
rect 660310 351363 660362 351415
rect 42166 351289 42218 351341
rect 57622 351289 57674 351341
rect 655318 348477 655370 348529
rect 676054 348477 676106 348529
rect 674518 345591 674570 345643
rect 676054 345591 676106 345643
rect 41782 342779 41834 342831
rect 53206 342779 53258 342831
rect 674422 342779 674474 342831
rect 676246 342779 676298 342831
rect 674710 342705 674762 342757
rect 676054 342705 676106 342757
rect 41782 342261 41834 342313
rect 50326 342261 50378 342313
rect 41782 341743 41834 341795
rect 48214 341743 48266 341795
rect 41782 341373 41834 341425
rect 43318 341373 43370 341425
rect 674806 341151 674858 341203
rect 676054 341151 676106 341203
rect 41590 340559 41642 340611
rect 43222 340559 43274 340611
rect 41782 340263 41834 340315
rect 46198 340263 46250 340315
rect 41590 340041 41642 340093
rect 43510 340041 43562 340093
rect 44374 340041 44426 340093
rect 674614 339967 674666 340019
rect 675958 339967 676010 340019
rect 674998 339893 675050 339945
rect 676246 339893 676298 339945
rect 674902 339819 674954 339871
rect 676054 339819 676106 339871
rect 41590 339079 41642 339131
rect 46102 339079 46154 339131
rect 41782 338857 41834 338909
rect 43414 338857 43466 338909
rect 44470 338857 44522 338909
rect 650230 337007 650282 337059
rect 679990 337007 680042 337059
rect 674518 335305 674570 335357
rect 675190 335305 675242 335357
rect 674710 334787 674762 334839
rect 675382 334787 675434 334839
rect 650422 334121 650474 334173
rect 655414 334121 655466 334173
rect 674422 331679 674474 331731
rect 675382 331679 675434 331731
rect 674998 330421 675050 330473
rect 675478 330421 675530 330473
rect 41782 330347 41834 330399
rect 45526 330347 45578 330399
rect 34486 329755 34538 329807
rect 41782 329755 41834 329807
rect 654166 328275 654218 328327
rect 675094 328275 675146 328327
rect 41782 327165 41834 327217
rect 674614 327091 674666 327143
rect 675478 327091 675530 327143
rect 41782 326943 41834 326995
rect 674806 326795 674858 326847
rect 675382 326795 675434 326847
rect 674902 326129 674954 326181
rect 675382 326129 675434 326181
rect 42166 323539 42218 323591
rect 42454 323539 42506 323591
rect 42166 321689 42218 321741
rect 42838 321689 42890 321741
rect 42454 319617 42506 319669
rect 58486 319617 58538 319669
rect 42838 316731 42890 316783
rect 59158 316731 59210 316783
rect 53206 313845 53258 313897
rect 59734 313845 59786 313897
rect 50326 313771 50378 313823
rect 59542 313771 59594 313823
rect 48214 313697 48266 313749
rect 59638 313697 59690 313749
rect 42166 308073 42218 308125
rect 59062 308073 59114 308125
rect 654070 305261 654122 305313
rect 676246 305335 676298 305387
rect 653782 305187 653834 305239
rect 676246 305187 676298 305239
rect 673366 304003 673418 304055
rect 676054 304003 676106 304055
rect 673174 302967 673226 303019
rect 676054 302967 676106 303019
rect 45334 302301 45386 302353
rect 46486 302301 46538 302353
rect 654166 302301 654218 302353
rect 676246 302301 676298 302353
rect 673270 301931 673322 301983
rect 676054 301931 676106 301983
rect 46198 300895 46250 300947
rect 46870 300895 46922 300947
rect 62710 300895 62762 300947
rect 39670 299637 39722 299689
rect 46870 299637 46922 299689
rect 41782 299563 41834 299615
rect 60214 299563 60266 299615
rect 46486 299489 46538 299541
rect 54550 299489 54602 299541
rect 41782 298527 41834 298579
rect 52822 298527 52874 298579
rect 41782 298157 41834 298209
rect 43222 298157 43274 298209
rect 46102 298083 46154 298135
rect 46870 298083 46922 298135
rect 62806 298083 62858 298135
rect 41782 297565 41834 297617
rect 43222 297565 43274 297617
rect 41782 297047 41834 297099
rect 46198 297047 46250 297099
rect 39862 296751 39914 296803
rect 46870 296751 46922 296803
rect 41590 296677 41642 296729
rect 57526 296677 57578 296729
rect 675190 296677 675242 296729
rect 676054 296677 676106 296729
rect 41590 295863 41642 295915
rect 46294 295863 46346 295915
rect 46102 293865 46154 293917
rect 59638 293865 59690 293917
rect 48982 293791 49034 293843
rect 58198 293791 58250 293843
rect 674998 293791 675050 293843
rect 676054 293791 676106 293843
rect 650326 291645 650378 291697
rect 679894 291719 679946 291771
rect 52822 291275 52874 291327
rect 59638 291275 59690 291327
rect 54550 290979 54602 291031
rect 44182 290905 44234 290957
rect 59062 290905 59114 290957
rect 63286 290831 63338 290883
rect 675190 290387 675242 290439
rect 675382 290387 675434 290439
rect 654166 289129 654218 289181
rect 660886 289129 660938 289181
rect 45814 288019 45866 288071
rect 59638 288019 59690 288071
rect 656566 287945 656618 287997
rect 675190 287945 675242 287997
rect 41782 287131 41834 287183
rect 44278 287131 44330 287183
rect 62230 286687 62282 286739
rect 62902 286687 62954 286739
rect 34486 286539 34538 286591
rect 41782 286539 41834 286591
rect 674998 286243 675050 286295
rect 675382 286243 675434 286295
rect 48214 285207 48266 285259
rect 59542 285207 59594 285259
rect 53206 285133 53258 285185
rect 58102 285133 58154 285185
rect 653782 284245 653834 284297
rect 658006 284245 658058 284297
rect 41782 284023 41834 284075
rect 41782 283727 41834 283779
rect 45334 282543 45386 282595
rect 59638 282543 59690 282595
rect 45622 282321 45674 282373
rect 58966 282321 59018 282373
rect 56182 282247 56234 282299
rect 57622 282247 57674 282299
rect 42166 281285 42218 281337
rect 46102 281285 46154 281337
rect 45718 279435 45770 279487
rect 59638 279435 59690 279487
rect 45910 279361 45962 279413
rect 58198 279361 58250 279413
rect 654742 279361 654794 279413
rect 663766 279361 663818 279413
rect 42166 279287 42218 279339
rect 48982 279287 49034 279339
rect 313558 278325 313610 278377
rect 404758 278325 404810 278377
rect 314902 278251 314954 278303
rect 408310 278251 408362 278303
rect 316630 278177 316682 278229
rect 411862 278177 411914 278229
rect 319510 278103 319562 278155
rect 418966 278103 419018 278155
rect 320950 278029 321002 278081
rect 422518 278029 422570 278081
rect 322102 277955 322154 278007
rect 426262 277955 426314 278007
rect 63382 277881 63434 277933
rect 381238 277881 381290 277933
rect 323830 277807 323882 277859
rect 429910 277807 429962 277859
rect 326422 277733 326474 277785
rect 437014 277733 437066 277785
rect 317878 277659 317930 277711
rect 415702 277659 415754 277711
rect 329302 277585 329354 277637
rect 444118 277585 444170 277637
rect 333622 277511 333674 277563
rect 454774 277511 454826 277563
rect 336694 277437 336746 277489
rect 461782 277437 461834 277489
rect 339286 277363 339338 277415
rect 468886 277363 468938 277415
rect 342166 277289 342218 277341
rect 475990 277289 476042 277341
rect 372502 277215 372554 277267
rect 550486 277215 550538 277267
rect 373846 277141 373898 277193
rect 554038 277141 554090 277193
rect 376822 277067 376874 277119
rect 561142 277067 561194 277119
rect 377974 276993 378026 277045
rect 564694 276993 564746 277045
rect 381046 276919 381098 276971
rect 571702 276919 571754 276971
rect 379414 276845 379466 276897
rect 568246 276845 568298 276897
rect 383638 276771 383690 276823
rect 578806 276771 578858 276823
rect 382294 276697 382346 276749
rect 575254 276697 575306 276749
rect 386518 276623 386570 276675
rect 585910 276623 585962 276675
rect 390838 276549 390890 276601
rect 596566 276549 596618 276601
rect 393910 276475 393962 276527
rect 603670 276475 603722 276527
rect 284470 276401 284522 276453
rect 332950 276401 333002 276453
rect 350230 276401 350282 276453
rect 496054 276401 496106 276453
rect 286102 276327 286154 276379
rect 336502 276327 336554 276379
rect 356182 276327 356234 276379
rect 510262 276327 510314 276379
rect 288694 276253 288746 276305
rect 343606 276253 343658 276305
rect 359158 276253 359210 276305
rect 517366 276253 517418 276305
rect 287350 276179 287402 276231
rect 340054 276179 340106 276231
rect 361750 276179 361802 276231
rect 524470 276179 524522 276231
rect 291862 276105 291914 276157
rect 350710 276105 350762 276157
rect 364630 276105 364682 276157
rect 531574 276105 531626 276157
rect 290326 276031 290378 276083
rect 347158 276031 347210 276083
rect 367702 276031 367754 276083
rect 538678 276031 538730 276083
rect 293014 275957 293066 276009
rect 354262 275957 354314 276009
rect 371062 275957 371114 276009
rect 546934 275957 546986 276009
rect 294646 275883 294698 275935
rect 357814 275883 357866 275935
rect 370294 275883 370346 275935
rect 545782 275883 545834 275935
rect 295894 275809 295946 275861
rect 361366 275809 361418 275861
rect 371926 275809 371978 275861
rect 549334 275809 549386 275861
rect 297334 275735 297386 275787
rect 364918 275735 364970 275787
rect 374614 275735 374666 275787
rect 556342 275735 556394 275787
rect 298966 275661 299018 275713
rect 368470 275661 368522 275713
rect 377494 275661 377546 275713
rect 563446 275661 563498 275713
rect 297814 275587 297866 275639
rect 366070 275587 366122 275639
rect 380566 275587 380618 275639
rect 570550 275587 570602 275639
rect 299350 275513 299402 275565
rect 369622 275513 369674 275565
rect 388918 275513 388970 275565
rect 591862 275513 591914 275565
rect 301846 275439 301898 275491
rect 375574 275439 375626 275491
rect 387766 275439 387818 275491
rect 588310 275439 588362 275491
rect 303286 275365 303338 275417
rect 379126 275365 379178 275417
rect 394678 275365 394730 275417
rect 606070 275365 606122 275417
rect 306166 275291 306218 275343
rect 386134 275291 386186 275343
rect 398230 275291 398282 275343
rect 308758 275217 308810 275269
rect 393238 275217 393290 275269
rect 400630 275217 400682 275269
rect 407926 275291 407978 275343
rect 613078 275291 613130 275343
rect 310390 275143 310442 275195
rect 396790 275143 396842 275195
rect 403222 275143 403274 275195
rect 614326 275217 614378 275269
rect 313078 275069 313130 275121
rect 403894 275069 403946 275121
rect 406390 275069 406442 275121
rect 620182 275143 620234 275195
rect 314710 274995 314762 275047
rect 407446 274995 407498 275047
rect 627286 275069 627338 275121
rect 634390 274995 634442 275047
rect 283030 274921 283082 274973
rect 329398 274921 329450 274973
rect 344566 274921 344618 274973
rect 481942 274921 481994 274973
rect 281782 274847 281834 274899
rect 325846 274847 325898 274899
rect 341686 274847 341738 274899
rect 474838 274847 474890 274899
rect 339094 274773 339146 274825
rect 467734 274773 467786 274825
rect 336022 274699 336074 274751
rect 460630 274699 460682 274751
rect 333142 274625 333194 274677
rect 453526 274625 453578 274677
rect 331894 274551 331946 274603
rect 449974 274551 450026 274603
rect 328822 274477 328874 274529
rect 442870 274477 442922 274529
rect 325942 274403 325994 274455
rect 435862 274403 435914 274455
rect 321622 274329 321674 274381
rect 425206 274329 425258 274381
rect 323350 274255 323402 274307
rect 428758 274255 428810 274307
rect 318934 274181 318986 274233
rect 418102 274181 418154 274233
rect 317302 274107 317354 274159
rect 414550 274107 414602 274159
rect 347062 274033 347114 274085
rect 401494 274033 401546 274085
rect 334294 273959 334346 274011
rect 387382 273959 387434 274011
rect 397558 273959 397610 274011
rect 407926 273959 407978 274011
rect 328342 273885 328394 273937
rect 380278 273885 380330 273937
rect 343606 273811 343658 273863
rect 394486 273811 394538 273863
rect 326806 273737 326858 273789
rect 373174 273737 373226 273789
rect 673174 273663 673226 273715
rect 679702 273663 679754 273715
rect 673270 273589 673322 273641
rect 679798 273589 679850 273641
rect 160438 273515 160490 273567
rect 207478 273515 207530 273567
rect 277750 273515 277802 273567
rect 316438 273515 316490 273567
rect 349462 273515 349514 273567
rect 493750 273515 493802 273567
rect 529846 273515 529898 273567
rect 624982 273515 625034 273567
rect 108406 273441 108458 273493
rect 109366 273441 109418 273493
rect 130870 273441 130922 273493
rect 190102 273441 190154 273493
rect 193558 273441 193610 273493
rect 221494 273441 221546 273493
rect 230134 273441 230186 273493
rect 242902 273441 242954 273493
rect 275350 273441 275402 273493
rect 310486 273441 310538 273493
rect 310582 273441 310634 273493
rect 344758 273441 344810 273493
rect 350038 273441 350090 273493
rect 494902 273441 494954 273493
rect 122614 273367 122666 273419
rect 123766 273367 123818 273419
rect 142678 273367 142730 273419
rect 209590 273367 209642 273419
rect 277078 273367 277130 273419
rect 314038 273367 314090 273419
rect 337942 273367 337994 273419
rect 341302 273367 341354 273419
rect 352438 273367 352490 273419
rect 500854 273367 500906 273419
rect 135574 273293 135626 273345
rect 209878 273293 209930 273345
rect 219574 273293 219626 273345
rect 238678 273293 238730 273345
rect 279670 273293 279722 273345
rect 321142 273293 321194 273345
rect 352630 273293 352682 273345
rect 502006 273293 502058 273345
rect 68278 273219 68330 273271
rect 142486 273219 142538 273271
rect 153334 273219 153386 273271
rect 207382 273219 207434 273271
rect 278230 273219 278282 273271
rect 317590 273219 317642 273271
rect 355510 273219 355562 273271
rect 509110 273219 509162 273271
rect 132022 273145 132074 273197
rect 209686 273145 209738 273197
rect 285622 273145 285674 273197
rect 335350 273145 335402 273197
rect 355030 273145 355082 273197
rect 507958 273145 508010 273197
rect 127318 273071 127370 273123
rect 209974 273071 210026 273123
rect 220726 273071 220778 273123
rect 239158 273071 239210 273123
rect 286774 273071 286826 273123
rect 338902 273071 338954 273123
rect 358582 273071 358634 273123
rect 125014 272997 125066 273049
rect 207286 272997 207338 273049
rect 217174 272997 217226 273049
rect 237622 272997 237674 273049
rect 284950 272997 285002 273049
rect 334198 272997 334250 273049
rect 360982 272997 361034 273049
rect 375190 273071 375242 273123
rect 514966 273071 515018 273123
rect 128470 272923 128522 272975
rect 210166 272923 210218 272975
rect 216022 272923 216074 272975
rect 236950 272923 237002 272975
rect 271030 272923 271082 272975
rect 299926 272923 299978 272975
rect 305398 272923 305450 272975
rect 358966 272923 359018 272975
rect 361270 272923 361322 272975
rect 516214 272997 516266 273049
rect 123670 272849 123722 272901
rect 209014 272849 209066 272901
rect 218326 272849 218378 272901
rect 238102 272849 238154 272901
rect 289942 272849 289994 272901
rect 346006 272849 346058 272901
rect 363574 272849 363626 272901
rect 522070 272923 522122 272975
rect 116662 272775 116714 272827
rect 207094 272775 207146 272827
rect 214774 272775 214826 272827
rect 236470 272775 236522 272827
rect 292246 272775 292298 272827
rect 351862 272775 351914 272827
rect 364150 272775 364202 272827
rect 523318 272849 523370 272901
rect 120214 272701 120266 272753
rect 207862 272701 207914 272753
rect 212470 272701 212522 272753
rect 235702 272701 235754 272753
rect 292726 272701 292778 272753
rect 353110 272701 353162 272753
rect 366550 272701 366602 272753
rect 529174 272775 529226 272827
rect 113110 272627 113162 272679
rect 206038 272627 206090 272679
rect 213622 272627 213674 272679
rect 236278 272627 236330 272679
rect 295414 272627 295466 272679
rect 360214 272627 360266 272679
rect 367126 272627 367178 272679
rect 530422 272701 530474 272753
rect 110806 272553 110858 272605
rect 205750 272553 205802 272605
rect 211222 272553 211274 272605
rect 235030 272553 235082 272605
rect 270262 272553 270314 272605
rect 297526 272553 297578 272605
rect 298294 272553 298346 272605
rect 367222 272553 367274 272605
rect 372694 272553 372746 272605
rect 536278 272627 536330 272679
rect 106102 272479 106154 272531
rect 204022 272479 204074 272531
rect 208918 272479 208970 272531
rect 234358 272479 234410 272531
rect 270550 272479 270602 272531
rect 298678 272479 298730 272531
rect 301366 272479 301418 272531
rect 374326 272479 374378 272531
rect 537430 272553 537482 272605
rect 551638 272479 551690 272531
rect 103702 272405 103754 272457
rect 203542 272405 203594 272457
rect 210070 272405 210122 272457
rect 234550 272405 234602 272457
rect 236086 272405 236138 272457
rect 245302 272405 245354 272457
rect 274198 272405 274250 272457
rect 306934 272405 306986 272457
rect 307126 272405 307178 272457
rect 388534 272405 388586 272457
rect 388630 272405 388682 272457
rect 572950 272405 573002 272457
rect 98998 272331 99050 272383
rect 199126 272331 199178 272383
rect 207670 272331 207722 272383
rect 233878 272331 233930 272383
rect 234934 272331 234986 272383
rect 244822 272331 244874 272383
rect 272758 272331 272810 272383
rect 303478 272331 303530 272383
rect 303958 272331 304010 272383
rect 381430 272331 381482 272383
rect 383446 272331 383498 272383
rect 577654 272331 577706 272383
rect 96598 272257 96650 272309
rect 201622 272257 201674 272309
rect 232534 272257 232586 272309
rect 243670 272257 243722 272309
rect 275158 272257 275210 272309
rect 309334 272257 309386 272309
rect 309910 272257 309962 272309
rect 395638 272257 395690 272309
rect 395926 272257 395978 272309
rect 608374 272257 608426 272309
rect 84790 272183 84842 272235
rect 86326 272183 86378 272235
rect 104854 272183 104906 272235
rect 106486 272183 106538 272235
rect 76534 272109 76586 272161
rect 195670 272183 195722 272235
rect 198262 272183 198314 272235
rect 224374 272183 224426 272235
rect 227830 272183 227882 272235
rect 242134 272183 242186 272235
rect 273430 272183 273482 272235
rect 305782 272183 305834 272235
rect 312790 272183 312842 272235
rect 402742 272183 402794 272235
rect 406102 272183 406154 272235
rect 413398 272183 413450 272235
rect 413494 272183 413546 272235
rect 636790 272183 636842 272235
rect 194710 272109 194762 272161
rect 224470 272109 224522 272161
rect 228982 272109 229034 272161
rect 242422 272109 242474 272161
rect 276310 272109 276362 272161
rect 312886 272109 312938 272161
rect 315478 272109 315530 272161
rect 409846 272109 409898 272161
rect 411862 272109 411914 272161
rect 643894 272109 643946 272161
rect 167542 272035 167594 272087
rect 210646 272035 210698 272087
rect 298006 272035 298058 272087
rect 327094 272035 327146 272087
rect 347254 272035 347306 272087
rect 487798 272035 487850 272087
rect 174646 271961 174698 272013
rect 210550 271961 210602 272013
rect 231382 271961 231434 272013
rect 243094 271961 243146 272013
rect 299446 271961 299498 272013
rect 328246 271961 328298 272013
rect 346486 271961 346538 272013
rect 486646 271961 486698 272013
rect 159286 271887 159338 271939
rect 192982 271887 193034 271939
rect 195862 271887 195914 271939
rect 221686 271887 221738 271939
rect 233686 271887 233738 271939
rect 244054 271887 244106 271939
rect 272278 271887 272330 271939
rect 301942 271887 301994 271939
rect 302326 271887 302378 271939
rect 324694 271887 324746 271939
rect 344086 271887 344138 271939
rect 480694 271887 480746 271939
rect 191158 271813 191210 271865
rect 227158 271813 227210 271865
rect 341494 271813 341546 271865
rect 473686 271813 473738 271865
rect 101302 271739 101354 271791
rect 103606 271739 103658 271791
rect 147382 271739 147434 271791
rect 149686 271739 149738 271791
rect 192310 271739 192362 271791
rect 224566 271739 224618 271791
rect 338614 271739 338666 271791
rect 466582 271739 466634 271791
rect 166294 271665 166346 271717
rect 198646 271665 198698 271717
rect 199414 271665 199466 271717
rect 221590 271665 221642 271717
rect 335446 271665 335498 271717
rect 459478 271665 459530 271717
rect 75286 271591 75338 271643
rect 77686 271591 77738 271643
rect 129718 271591 129770 271643
rect 132406 271591 132458 271643
rect 181750 271591 181802 271643
rect 210454 271591 210506 271643
rect 332566 271591 332618 271643
rect 452374 271591 452426 271643
rect 89494 271517 89546 271569
rect 92086 271517 92138 271569
rect 150934 271517 150986 271569
rect 152374 271517 152426 271569
rect 180502 271517 180554 271569
rect 205174 271517 205226 271569
rect 329974 271517 330026 271569
rect 445270 271517 445322 271569
rect 173398 271443 173450 271495
rect 201526 271443 201578 271495
rect 201814 271443 201866 271495
rect 223702 271443 223754 271495
rect 326902 271443 326954 271495
rect 438166 271443 438218 271495
rect 185206 271369 185258 271421
rect 210358 271369 210410 271421
rect 334102 271369 334154 271421
rect 337750 271369 337802 271421
rect 346966 271369 347018 271421
rect 431062 271369 431114 271421
rect 184054 271295 184106 271347
rect 205942 271295 205994 271347
rect 321430 271295 321482 271347
rect 423958 271295 424010 271347
rect 161590 271221 161642 271273
rect 163894 271221 163946 271273
rect 188758 271221 188810 271273
rect 210262 271221 210314 271273
rect 237238 271221 237290 271273
rect 245590 271221 245642 271273
rect 318358 271221 318410 271273
rect 416950 271221 417002 271273
rect 175798 271147 175850 271199
rect 178294 271147 178346 271199
rect 187606 271147 187658 271199
rect 205846 271147 205898 271199
rect 238486 271147 238538 271199
rect 246070 271147 246122 271199
rect 324022 271147 324074 271199
rect 346966 271147 347018 271199
rect 357910 271147 357962 271199
rect 375190 271147 375242 271199
rect 409846 271147 409898 271199
rect 413494 271147 413546 271199
rect 85942 271073 85994 271125
rect 198550 271073 198602 271125
rect 205366 271073 205418 271125
rect 232630 271073 232682 271125
rect 240790 271073 240842 271125
rect 247222 271073 247274 271125
rect 221878 270999 221930 271051
rect 239350 270999 239402 271051
rect 239542 270999 239594 271051
rect 241270 270999 241322 271051
rect 241942 270999 241994 271051
rect 247702 270999 247754 271051
rect 342742 270999 342794 271051
rect 348310 270999 348362 271051
rect 223030 270925 223082 270977
rect 240022 270925 240074 270977
rect 243190 270925 243242 270977
rect 247990 270925 248042 270977
rect 224278 270851 224330 270903
rect 240502 270851 240554 270903
rect 244342 270851 244394 270903
rect 248662 270851 248714 270903
rect 225430 270777 225482 270829
rect 241078 270777 241130 270829
rect 245494 270777 245546 270829
rect 249142 270777 249194 270829
rect 94198 270703 94250 270755
rect 94966 270703 95018 270755
rect 115510 270703 115562 270755
rect 118006 270703 118058 270755
rect 119062 270703 119114 270755
rect 120886 270703 120938 270755
rect 133270 270703 133322 270755
rect 135286 270703 135338 270755
rect 136822 270703 136874 270755
rect 138166 270703 138218 270755
rect 154486 270703 154538 270755
rect 155446 270703 155498 270755
rect 165142 270703 165194 270755
rect 166966 270703 167018 270755
rect 168694 270703 168746 270755
rect 169846 270703 169898 270755
rect 179350 270703 179402 270755
rect 181366 270703 181418 270755
rect 182902 270703 182954 270755
rect 184246 270703 184298 270755
rect 185494 270703 185546 270755
rect 186454 270703 186506 270755
rect 226582 270703 226634 270755
rect 239542 270703 239594 270755
rect 239638 270703 239690 270755
rect 246454 270703 246506 270755
rect 246742 270703 246794 270755
rect 249622 270703 249674 270755
rect 351382 270703 351434 270755
rect 355414 270703 355466 270755
rect 146230 270629 146282 270681
rect 214966 270629 215018 270681
rect 280150 270629 280202 270681
rect 322390 270629 322442 270681
rect 350710 270629 350762 270681
rect 497302 270629 497354 270681
rect 137974 270555 138026 270607
rect 212662 270555 212714 270607
rect 280630 270555 280682 270607
rect 323542 270555 323594 270607
rect 351286 270555 351338 270607
rect 498454 270555 498506 270607
rect 141526 270481 141578 270533
rect 213814 270481 213866 270533
rect 264694 270481 264746 270533
rect 283318 270481 283370 270533
rect 134422 270407 134474 270459
rect 211894 270407 211946 270459
rect 253942 270407 253994 270459
rect 257302 270407 257354 270459
rect 264886 270407 264938 270459
rect 276406 270407 276458 270459
rect 279286 270407 279338 270459
rect 319990 270481 320042 270533
rect 353686 270481 353738 270533
rect 504406 270481 504458 270533
rect 283702 270407 283754 270459
rect 330646 270407 330698 270459
rect 354070 270407 354122 270459
rect 505558 270407 505610 270459
rect 121462 270333 121514 270385
rect 208342 270333 208394 270385
rect 262486 270333 262538 270385
rect 278614 270333 278666 270385
rect 284182 270333 284234 270385
rect 331798 270333 331850 270385
rect 356758 270333 356810 270385
rect 511510 270333 511562 270385
rect 117910 270259 117962 270311
rect 207574 270259 207626 270311
rect 255286 270259 255338 270311
rect 260854 270259 260906 270311
rect 266038 270259 266090 270311
rect 286870 270259 286922 270311
rect 114358 270185 114410 270237
rect 206422 270185 206474 270237
rect 210550 270185 210602 270237
rect 222838 270185 222890 270237
rect 265366 270185 265418 270237
rect 109558 270111 109610 270163
rect 205270 270111 205322 270163
rect 210262 270111 210314 270163
rect 226678 270111 226730 270163
rect 266518 270111 266570 270163
rect 276406 270185 276458 270237
rect 284566 270185 284618 270237
rect 286294 270185 286346 270237
rect 334102 270259 334154 270311
rect 356950 270259 357002 270311
rect 512662 270259 512714 270311
rect 288502 270185 288554 270237
rect 342454 270185 342506 270237
rect 359830 270185 359882 270237
rect 519766 270185 519818 270237
rect 102550 270037 102602 270089
rect 203350 270037 203402 270089
rect 210358 270037 210410 270089
rect 225526 270037 225578 270089
rect 267286 270037 267338 270089
rect 285718 270111 285770 270163
rect 287926 270111 287978 270163
rect 337942 270111 337994 270163
rect 359350 270111 359402 270163
rect 518518 270111 518570 270163
rect 107254 269963 107306 270015
rect 204694 269963 204746 270015
rect 210454 269963 210506 270015
rect 224758 269963 224810 270015
rect 267094 269963 267146 270015
rect 288022 270037 288074 270089
rect 290614 270037 290666 270089
rect 342742 270037 342794 270089
rect 362230 270037 362282 270089
rect 525622 270037 525674 270089
rect 100150 269889 100202 269941
rect 202870 269889 202922 269941
rect 205174 269889 205226 269941
rect 224086 269889 224138 269941
rect 256246 269889 256298 269941
rect 263254 269889 263306 269941
rect 267766 269889 267818 269941
rect 290422 269963 290474 270015
rect 291094 269963 291146 270015
rect 349558 269963 349610 270015
rect 362806 269963 362858 270015
rect 526870 269963 526922 270015
rect 95446 269815 95498 269867
rect 185686 269815 185738 269867
rect 205942 269815 205994 269867
rect 225238 269815 225290 269867
rect 255766 269815 255818 269867
rect 262102 269815 262154 269867
rect 269206 269815 269258 269867
rect 289270 269889 289322 269941
rect 293974 269889 294026 269941
rect 356662 269889 356714 269941
rect 365302 269889 365354 269941
rect 532726 269889 532778 269941
rect 93046 269741 93098 269793
rect 200950 269741 201002 269793
rect 205846 269741 205898 269793
rect 226006 269741 226058 269793
rect 291574 269815 291626 269867
rect 293494 269815 293546 269867
rect 351382 269815 351434 269867
rect 365686 269815 365738 269867
rect 533878 269815 533930 269867
rect 295126 269741 295178 269793
rect 297046 269741 297098 269793
rect 363670 269741 363722 269793
rect 371254 269741 371306 269793
rect 548086 269741 548138 269793
rect 90646 269667 90698 269719
rect 199702 269667 199754 269719
rect 201526 269667 201578 269719
rect 222358 269667 222410 269719
rect 259894 269667 259946 269719
rect 271510 269667 271562 269719
rect 271606 269667 271658 269719
rect 293782 269667 293834 269719
rect 299638 269667 299690 269719
rect 370774 269667 370826 269719
rect 379894 269667 379946 269719
rect 569398 269667 569450 269719
rect 83638 269593 83690 269645
rect 198070 269593 198122 269645
rect 198646 269593 198698 269645
rect 220534 269593 220586 269645
rect 249046 269593 249098 269645
rect 250294 269593 250346 269645
rect 257686 269593 257738 269645
rect 266806 269593 266858 269645
rect 269686 269593 269738 269645
rect 296374 269593 296426 269645
rect 302614 269593 302666 269645
rect 377878 269593 377930 269645
rect 384118 269593 384170 269645
rect 580054 269593 580106 269645
rect 87190 269519 87242 269571
rect 199030 269519 199082 269571
rect 206518 269519 206570 269571
rect 233398 269519 233450 269571
rect 271510 269519 271562 269571
rect 301078 269519 301130 269571
rect 305686 269519 305738 269571
rect 384982 269519 385034 269571
rect 385366 269519 385418 269571
rect 582358 269519 582410 269571
rect 81238 269445 81290 269497
rect 196822 269445 196874 269497
rect 202966 269445 203018 269497
rect 231958 269445 232010 269497
rect 260086 269445 260138 269497
rect 272662 269445 272714 269497
rect 272950 269445 273002 269497
rect 304630 269445 304682 269497
rect 308278 269445 308330 269497
rect 392086 269445 392138 269497
rect 82390 269371 82442 269423
rect 197398 269371 197450 269423
rect 204118 269371 204170 269423
rect 232150 269371 232202 269423
rect 274678 269371 274730 269423
rect 308182 269371 308234 269423
rect 311158 269371 311210 269423
rect 399190 269371 399242 269423
rect 399958 269371 400010 269423
rect 619030 269371 619082 269423
rect 74134 269297 74186 269349
rect 194998 269297 195050 269349
rect 200662 269297 200714 269349
rect 230998 269297 231050 269349
rect 258646 269297 258698 269349
rect 269110 269297 269162 269349
rect 278902 269297 278954 269349
rect 318838 269297 318890 269349
rect 319030 269297 319082 269349
rect 406102 269297 406154 269349
rect 409654 269297 409706 269349
rect 642646 269297 642698 269349
rect 67030 269223 67082 269275
rect 192598 269223 192650 269275
rect 197110 269223 197162 269275
rect 229558 269223 229610 269275
rect 257494 269223 257546 269275
rect 265654 269223 265706 269275
rect 268630 269223 268682 269275
rect 271606 269223 271658 269275
rect 275830 269223 275882 269275
rect 311734 269223 311786 269275
rect 314230 269223 314282 269275
rect 406294 269223 406346 269275
rect 408502 269223 408554 269275
rect 640342 269223 640394 269275
rect 145078 269149 145130 269201
rect 214486 269149 214538 269201
rect 262006 269149 262058 269201
rect 277462 269149 277514 269201
rect 277558 269149 277610 269201
rect 315286 269149 315338 269201
rect 348118 269149 348170 269201
rect 490198 269149 490250 269201
rect 152182 269075 152234 269127
rect 216694 269075 216746 269127
rect 253366 269075 253418 269127
rect 256150 269075 256202 269127
rect 259414 269075 259466 269127
rect 270358 269075 270410 269127
rect 295222 269075 295274 269127
rect 305398 269075 305450 269127
rect 309238 269075 309290 269127
rect 343606 269075 343658 269127
rect 348406 269075 348458 269127
rect 491350 269075 491402 269127
rect 149782 269001 149834 269053
rect 216214 269001 216266 269053
rect 261814 269001 261866 269053
rect 276214 269001 276266 269053
rect 281302 269001 281354 269053
rect 302326 269001 302378 269053
rect 306358 269001 306410 269053
rect 334294 269001 334346 269053
rect 345430 269001 345482 269053
rect 484246 269001 484298 269053
rect 148630 268927 148682 268979
rect 215734 268927 215786 268979
rect 253174 268927 253226 268979
rect 254998 268927 255050 268979
rect 261238 268927 261290 268979
rect 275062 268927 275114 268979
rect 282070 268927 282122 268979
rect 298006 268927 298058 268979
rect 300694 268927 300746 268979
rect 326806 268927 326858 268979
rect 342646 268927 342698 268979
rect 477142 268927 477194 268979
rect 155734 268853 155786 268905
rect 217366 268853 217418 268905
rect 264118 268853 264170 268905
rect 282166 268853 282218 268905
rect 303766 268853 303818 268905
rect 328342 268853 328394 268905
rect 339766 268853 339818 268905
rect 470134 268853 470186 268905
rect 42070 268779 42122 268831
rect 44182 268779 44234 268831
rect 156886 268779 156938 268831
rect 218134 268779 218186 268831
rect 258166 268779 258218 268831
rect 267958 268779 268010 268831
rect 289174 268779 289226 268831
rect 310582 268779 310634 268831
rect 336886 268779 336938 268831
rect 463030 268779 463082 268831
rect 162838 268705 162890 268757
rect 219286 268705 219338 268757
rect 268438 268705 268490 268757
rect 292822 268705 292874 268757
rect 334294 268705 334346 268757
rect 455926 268705 455978 268757
rect 163990 268631 164042 268683
rect 219958 268631 220010 268683
rect 254614 268631 254666 268683
rect 258550 268631 258602 268683
rect 260566 268631 260618 268683
rect 273910 268631 273962 268683
rect 331222 268631 331274 268683
rect 448822 268631 448874 268683
rect 169750 268557 169802 268609
rect 221206 268557 221258 268609
rect 328342 268557 328394 268609
rect 441718 268557 441770 268609
rect 171094 268483 171146 268535
rect 221782 268483 221834 268535
rect 263638 268483 263690 268535
rect 281014 268483 281066 268535
rect 325750 268483 325802 268535
rect 434614 268483 434666 268535
rect 176950 268409 177002 268461
rect 223414 268409 223466 268461
rect 322582 268409 322634 268461
rect 427510 268409 427562 268461
rect 178198 268335 178250 268387
rect 223606 268335 223658 268387
rect 247894 268335 247946 268387
rect 249814 268335 249866 268387
rect 255094 268335 255146 268387
rect 259702 268335 259754 268387
rect 262966 268335 263018 268387
rect 279766 268335 279818 268387
rect 319702 268335 319754 268387
rect 420502 268335 420554 268387
rect 185686 268261 185738 268313
rect 201142 268261 201194 268313
rect 207478 268261 207530 268313
rect 192982 268187 193034 268239
rect 210838 268187 210890 268239
rect 190102 268113 190154 268165
rect 210742 268113 210794 268165
rect 211030 268261 211082 268313
rect 218614 268261 218666 268313
rect 221494 268261 221546 268313
rect 227830 268261 227882 268313
rect 312310 268261 312362 268313
rect 347062 268261 347114 268313
rect 224374 268187 224426 268239
rect 230038 268187 230090 268239
rect 257014 268187 257066 268239
rect 264406 268187 264458 268239
rect 332374 268187 332426 268239
rect 344854 268187 344906 268239
rect 345238 268187 345290 268239
rect 354550 268187 354602 268239
rect 394390 268187 394442 268239
rect 604822 268187 604874 268239
rect 218902 268113 218954 268165
rect 223702 268113 223754 268165
rect 231478 268113 231530 268165
rect 334966 268113 335018 268165
rect 348502 268113 348554 268165
rect 207382 268039 207434 268091
rect 216886 268039 216938 268091
rect 221590 268039 221642 268091
rect 230518 268039 230570 268091
rect 252694 268039 252746 268091
rect 253750 268039 253802 268091
rect 341014 268039 341066 268091
rect 209878 267965 209930 268017
rect 212374 267965 212426 268017
rect 221686 267965 221738 268017
rect 229078 267965 229130 268017
rect 337846 267965 337898 268017
rect 354262 267965 354314 268017
rect 357526 267965 357578 268017
rect 207286 267891 207338 267943
rect 209494 267891 209546 267943
rect 210646 267891 210698 267943
rect 221014 267891 221066 267943
rect 224470 267891 224522 267943
rect 228406 267891 228458 267943
rect 343606 267891 343658 267943
rect 199126 267817 199178 267869
rect 202294 267817 202346 267869
rect 209686 267817 209738 267869
rect 211414 267817 211466 267869
rect 224566 267817 224618 267869
rect 227638 267817 227690 267869
rect 282550 267817 282602 267869
rect 299446 267817 299498 267869
rect 317110 267817 317162 267869
rect 319030 267817 319082 267869
rect 354550 267891 354602 267943
rect 385462 267891 385514 267943
rect 360694 267817 360746 267869
rect 407254 267817 407306 267869
rect 409846 267817 409898 267869
rect 409942 267817 409994 267869
rect 411862 267817 411914 267869
rect 354838 267743 354890 267795
rect 506710 267743 506762 267795
rect 357430 267669 357482 267721
rect 513814 267669 513866 267721
rect 360310 267595 360362 267647
rect 520918 267595 520970 267647
rect 363382 267521 363434 267573
rect 528022 267521 528074 267573
rect 365974 267447 366026 267499
rect 535126 267447 535178 267499
rect 368950 267373 369002 267425
rect 542230 267373 542282 267425
rect 375094 267299 375146 267351
rect 557590 267299 557642 267351
rect 384886 267225 384938 267277
rect 581206 267225 581258 267277
rect 386038 267151 386090 267203
rect 584758 267151 584810 267203
rect 296470 267077 296522 267129
rect 362518 267077 362570 267129
rect 387958 267077 388010 267129
rect 589462 267077 589514 267129
rect 300214 267003 300266 267055
rect 372022 267003 372074 267055
rect 391990 267003 392042 267055
rect 598966 267003 599018 267055
rect 302038 266929 302090 266981
rect 376726 266929 376778 266981
rect 393238 266929 393290 266981
rect 602518 266929 602570 266981
rect 304438 266855 304490 266907
rect 382582 266855 382634 266907
rect 396310 266855 396362 266907
rect 609526 266855 609578 266907
rect 305014 266781 305066 266833
rect 383830 266781 383882 266833
rect 398902 266781 398954 266833
rect 616630 266781 616682 266833
rect 308086 266707 308138 266759
rect 390934 266707 390986 266759
rect 401782 266707 401834 266759
rect 623734 266707 623786 266759
rect 307318 266633 307370 266685
rect 389686 266633 389738 266685
rect 403702 266633 403754 266685
rect 628438 266633 628490 266685
rect 310678 266559 310730 266611
rect 398038 266559 398090 266611
rect 404950 266559 405002 266611
rect 630838 266559 630890 266611
rect 315958 266485 316010 266537
rect 408982 266485 409034 266537
rect 409174 266485 409226 266537
rect 641494 266485 641546 266537
rect 187222 266411 187274 266463
rect 189718 266411 189770 266463
rect 311638 266411 311690 266463
rect 400342 266411 400394 266463
rect 407830 266411 407882 266463
rect 637942 266411 637994 266463
rect 46102 266337 46154 266389
rect 652246 266337 652298 266389
rect 351958 266263 352010 266315
rect 499606 266263 499658 266315
rect 348886 266189 348938 266241
rect 492598 266189 492650 266241
rect 346006 266115 346058 266167
rect 485494 266115 485546 266167
rect 343318 266041 343370 266093
rect 478390 266041 478442 266093
rect 340246 265967 340298 266019
rect 471286 265967 471338 266019
rect 337366 265893 337418 265945
rect 464182 265893 464234 265945
rect 334774 265819 334826 265871
rect 457078 265819 457130 265871
rect 330454 265745 330506 265797
rect 446422 265745 446474 265797
rect 327574 265671 327626 265723
rect 439318 265671 439370 265723
rect 324502 265597 324554 265649
rect 432310 265597 432362 265649
rect 320182 265523 320234 265575
rect 408982 265523 409034 265575
rect 410998 265523 411050 265575
rect 421654 265375 421706 265427
rect 385462 265301 385514 265353
rect 483094 265449 483146 265501
rect 23062 265005 23114 265057
rect 46102 265005 46154 265057
rect 46198 264931 46250 264983
rect 669814 264931 669866 264983
rect 360694 264857 360746 264909
rect 479542 264857 479594 264909
rect 357526 264783 357578 264835
rect 472438 264783 472490 264835
rect 354262 264709 354314 264761
rect 465334 264709 465386 264761
rect 348502 264635 348554 264687
rect 458230 264635 458282 264687
rect 331126 264561 331178 264613
rect 447670 264561 447722 264613
rect 344854 264487 344906 264539
rect 451222 264487 451274 264539
rect 328054 264413 328106 264465
rect 440566 264413 440618 264465
rect 408022 264117 408074 264169
rect 412822 264117 412874 264169
rect 324982 264043 325034 264095
rect 433462 264043 433514 264095
rect 389446 263969 389498 264021
rect 593014 263969 593066 264021
rect 392278 263895 392330 263947
rect 600118 263895 600170 263947
rect 395446 263821 395498 263873
rect 607222 263821 607274 263873
rect 399670 263747 399722 263799
rect 617878 263747 617930 263799
rect 401110 263673 401162 263725
rect 621430 263673 621482 263725
rect 23350 263599 23402 263651
rect 46198 263599 46250 263651
rect 406870 263599 406922 263651
rect 427606 263599 427658 263651
rect 23254 263525 23306 263577
rect 46294 263525 46346 263577
rect 405430 263525 405482 263577
rect 631990 263599 632042 263651
rect 427894 263525 427946 263577
rect 635542 263525 635594 263577
rect 412822 263451 412874 263503
rect 639094 263451 639146 263503
rect 656374 262415 656426 262467
rect 676054 262415 676106 262467
rect 656182 262267 656234 262319
rect 676246 262267 676298 262319
rect 23158 262119 23210 262171
rect 46198 262119 46250 262171
rect 420406 262119 420458 262171
rect 606166 262119 606218 262171
rect 673366 261601 673418 261653
rect 676054 261601 676106 261653
rect 656086 259455 656138 259507
rect 676246 259455 676298 259507
rect 420406 259233 420458 259285
rect 606262 259233 606314 259285
rect 674710 256939 674762 256991
rect 676054 256939 676106 256991
rect 40246 256347 40298 256399
rect 48214 256347 48266 256399
rect 420406 256347 420458 256399
rect 606358 256347 606410 256399
rect 41782 255385 41834 255437
rect 53206 255385 53258 255437
rect 48022 255015 48074 255067
rect 186358 255015 186410 255067
rect 41782 254941 41834 254993
rect 43222 254941 43274 254993
rect 47542 254941 47594 254993
rect 185974 254941 186026 254993
rect 48118 254867 48170 254919
rect 186550 254867 186602 254919
rect 41782 254423 41834 254475
rect 43222 254423 43274 254475
rect 675094 253609 675146 253661
rect 676246 253609 676298 253661
rect 674902 253535 674954 253587
rect 675958 253535 676010 253587
rect 41590 253461 41642 253513
rect 56182 253461 56234 253513
rect 420406 253461 420458 253513
rect 603286 253461 603338 253513
rect 675286 253461 675338 253513
rect 676054 253461 676106 253513
rect 141046 252425 141098 252477
rect 174262 252425 174314 252477
rect 97846 252351 97898 252403
rect 156886 252351 156938 252403
rect 94966 252277 95018 252329
rect 154006 252277 154058 252329
rect 103606 252203 103658 252255
rect 165526 252203 165578 252255
rect 106486 252129 106538 252181
rect 171286 252129 171338 252181
rect 109366 252055 109418 252107
rect 179926 252055 179978 252107
rect 56086 251981 56138 252033
rect 186454 251981 186506 252033
rect 674518 250723 674570 250775
rect 675958 250723 676010 250775
rect 674614 250649 674666 250701
rect 676246 250649 676298 250701
rect 420406 250575 420458 250627
rect 603382 250575 603434 250627
rect 674998 250575 675050 250627
rect 676054 250575 676106 250627
rect 135286 249909 135338 249961
rect 145558 249909 145610 249961
rect 138166 249835 138218 249887
rect 171478 249835 171530 249887
rect 118006 249761 118058 249813
rect 156982 249761 157034 249813
rect 123766 249687 123818 249739
rect 162742 249687 162794 249739
rect 126646 249613 126698 249665
rect 168502 249613 168554 249665
rect 120886 249539 120938 249591
rect 165622 249539 165674 249591
rect 132406 249465 132458 249517
rect 180118 249465 180170 249517
rect 92086 249391 92138 249443
rect 159766 249391 159818 249443
rect 77686 249317 77738 249369
rect 145366 249317 145418 249369
rect 86326 249243 86378 249295
rect 177046 249243 177098 249295
rect 80566 249169 80618 249221
rect 182806 249169 182858 249221
rect 47926 249095 47978 249147
rect 186742 249095 186794 249147
rect 646678 249095 646730 249147
rect 679990 249095 680042 249147
rect 420310 247763 420362 247815
rect 603478 247763 603530 247815
rect 420406 247689 420458 247741
rect 629206 247689 629258 247741
rect 675766 247097 675818 247149
rect 112246 246653 112298 246705
rect 185782 246653 185834 246705
rect 675094 246653 675146 246705
rect 675478 246653 675530 246705
rect 47638 246579 47690 246631
rect 186070 246579 186122 246631
rect 675766 246579 675818 246631
rect 47734 246505 47786 246557
rect 186262 246505 186314 246557
rect 47446 246431 47498 246483
rect 186166 246431 186218 246483
rect 47830 246357 47882 246409
rect 186646 246357 186698 246409
rect 45526 246283 45578 246335
rect 186838 246283 186890 246335
rect 44278 246209 44330 246261
rect 187030 246209 187082 246261
rect 674710 245395 674762 245447
rect 675382 245395 675434 245447
rect 41590 244951 41642 245003
rect 145462 244951 145514 245003
rect 44758 244877 44810 244929
rect 186934 244877 186986 244929
rect 41782 244803 41834 244855
rect 145654 244803 145706 244855
rect 420406 244803 420458 244855
rect 629302 244803 629354 244855
rect 674902 242879 674954 242931
rect 675382 242879 675434 242931
rect 44662 242805 44714 242857
rect 185686 242805 185738 242857
rect 44566 242731 44618 242783
rect 185590 242731 185642 242783
rect 44854 242657 44906 242709
rect 185878 242657 185930 242709
rect 41590 242583 41642 242635
rect 142582 242583 142634 242635
rect 675190 242287 675242 242339
rect 675382 242287 675434 242339
rect 420406 241917 420458 241969
rect 600406 241917 600458 241969
rect 655894 241843 655946 241895
rect 675094 241843 675146 241895
rect 674998 241769 675050 241821
rect 675382 241769 675434 241821
rect 41782 240807 41834 240859
rect 41782 240511 41834 240563
rect 380854 239919 380906 239971
rect 412054 239919 412106 239971
rect 409558 239845 409610 239897
rect 412150 239845 412202 239897
rect 357142 239771 357194 239823
rect 434614 239771 434666 239823
rect 377302 239697 377354 239749
rect 446710 239697 446762 239749
rect 385366 239623 385418 239675
rect 470902 239623 470954 239675
rect 374422 239549 374474 239601
rect 488278 239549 488330 239601
rect 334294 239475 334346 239527
rect 458806 239475 458858 239527
rect 394678 239401 394730 239453
rect 532822 239401 532874 239453
rect 397750 239327 397802 239379
rect 541462 239327 541514 239379
rect 406006 239253 406058 239305
rect 550870 239253 550922 239305
rect 420406 239179 420458 239231
rect 599158 239179 599210 239231
rect 350422 239105 350474 239157
rect 508630 239105 508682 239157
rect 368566 239031 368618 239083
rect 544822 239031 544874 239083
rect 324406 238957 324458 239009
rect 455062 238957 455114 239009
rect 323926 238883 323978 238935
rect 455158 238883 455210 238935
rect 326710 238809 326762 238861
rect 462550 238809 462602 238861
rect 328918 238735 328970 238787
rect 464758 238735 464810 238787
rect 329878 238661 329930 238713
rect 468598 238661 468650 238713
rect 332662 238587 332714 238639
rect 474646 238587 474698 238639
rect 674614 238587 674666 238639
rect 675382 238587 675434 238639
rect 335734 238513 335786 238565
rect 480694 238513 480746 238565
rect 336694 238439 336746 238491
rect 478102 238439 478154 238491
rect 338998 238365 339050 238417
rect 486742 238365 486794 238417
rect 341782 238291 341834 238343
rect 492790 238291 492842 238343
rect 345334 238217 345386 238269
rect 500278 238217 500330 238269
rect 346678 238143 346730 238195
rect 503350 238143 503402 238195
rect 349942 238069 349994 238121
rect 509398 238069 509450 238121
rect 353494 237995 353546 238047
rect 514678 237995 514730 238047
rect 352726 237921 352778 237973
rect 512758 237921 512810 237973
rect 355702 237847 355754 237899
rect 522166 237847 522218 237899
rect 363094 237773 363146 237825
rect 535126 237773 535178 237825
rect 275350 237699 275402 237751
rect 357526 237699 357578 237751
rect 361750 237699 361802 237751
rect 533494 237699 533546 237751
rect 277078 237625 277130 237677
rect 363670 237625 363722 237677
rect 364438 237625 364490 237677
rect 535798 237625 535850 237677
rect 365878 237551 365930 237603
rect 541078 237551 541130 237603
rect 674518 237551 674570 237603
rect 675382 237551 675434 237603
rect 320854 237477 320906 237529
rect 450454 237477 450506 237529
rect 317590 237403 317642 237455
rect 444502 237403 444554 237455
rect 317110 237329 317162 237381
rect 441430 237329 441482 237381
rect 314806 237255 314858 237307
rect 438358 237255 438410 237307
rect 311542 237181 311594 237233
rect 432406 237181 432458 237233
rect 308566 237107 308618 237159
rect 426358 237107 426410 237159
rect 310774 237033 310826 237085
rect 428662 237033 428714 237085
rect 305782 236959 305834 237011
rect 420310 236959 420362 237011
rect 298966 236885 299018 236937
rect 404470 236885 404522 236937
rect 405910 236885 405962 236937
rect 414454 236885 414506 236937
rect 279862 236811 279914 236863
rect 370486 236811 370538 236863
rect 386998 236811 387050 236863
rect 387574 236811 387626 236863
rect 397078 236811 397130 236863
rect 397654 236811 397706 236863
rect 398038 236811 398090 236863
rect 413590 236811 413642 236863
rect 278422 236737 278474 236789
rect 366742 236737 366794 236789
rect 396982 236737 397034 236789
rect 413398 236737 413450 236789
rect 379798 236663 379850 236715
rect 398326 236663 398378 236715
rect 410710 236367 410762 236419
rect 442198 236367 442250 236419
rect 390742 236293 390794 236345
rect 492022 236293 492074 236345
rect 394582 236219 394634 236271
rect 505654 236219 505706 236271
rect 382390 236145 382442 236197
rect 397366 236145 397418 236197
rect 400342 236145 400394 236197
rect 523798 236145 523850 236197
rect 251062 236071 251114 236123
rect 273718 236071 273770 236123
rect 277558 236071 277610 236123
rect 313942 236071 313994 236123
rect 326134 236071 326186 236123
rect 334294 236071 334346 236123
rect 341206 236071 341258 236123
rect 374422 236071 374474 236123
rect 376342 236071 376394 236123
rect 208438 235997 208490 236049
rect 223222 235997 223274 236049
rect 247990 235997 248042 236049
rect 273622 235997 273674 236049
rect 276118 235997 276170 236049
rect 308278 235997 308330 236049
rect 313846 235997 313898 236049
rect 357142 235997 357194 236049
rect 371830 235997 371882 236049
rect 406006 235997 406058 236049
rect 146998 235923 147050 235975
rect 151222 235923 151274 235975
rect 207478 235923 207530 235975
rect 223990 235923 224042 235975
rect 243286 235923 243338 235975
rect 271030 235923 271082 235975
rect 280630 235923 280682 235975
rect 320854 235923 320906 235975
rect 386710 235923 386762 235975
rect 405622 235923 405674 235975
rect 410038 236071 410090 236123
rect 584566 236071 584618 236123
rect 406294 235997 406346 236049
rect 415414 235997 415466 236049
rect 413878 235923 413930 235975
rect 209686 235849 209738 235901
rect 226198 235849 226250 235901
rect 234262 235849 234314 235901
rect 264886 235849 264938 235901
rect 279286 235849 279338 235901
rect 319606 235849 319658 235901
rect 326230 235849 326282 235901
rect 460246 235849 460298 235901
rect 208918 235775 208970 235827
rect 226966 235775 227018 235827
rect 237526 235775 237578 235827
rect 268630 235775 268682 235827
rect 290326 235775 290378 235827
rect 334102 235775 334154 235827
rect 343510 235775 343562 235827
rect 495766 235775 495818 235827
rect 211222 235701 211274 235753
rect 229270 235701 229322 235753
rect 231190 235701 231242 235753
rect 259030 235701 259082 235753
rect 262870 235701 262922 235753
rect 305110 235701 305162 235753
rect 317206 235701 317258 235753
rect 410710 235701 410762 235753
rect 210646 235627 210698 235679
rect 230038 235627 230090 235679
rect 239350 235627 239402 235679
rect 287350 235627 287402 235679
rect 311158 235627 311210 235679
rect 210070 235553 210122 235605
rect 227830 235553 227882 235605
rect 236470 235553 236522 235605
rect 282934 235553 282986 235605
rect 287062 235553 287114 235605
rect 318166 235553 318218 235605
rect 358006 235553 358058 235605
rect 400342 235553 400394 235605
rect 405622 235627 405674 235679
rect 413686 235701 413738 235753
rect 412150 235627 412202 235679
rect 590422 235627 590474 235679
rect 408982 235553 409034 235605
rect 409174 235553 409226 235605
rect 588790 235553 588842 235605
rect 212950 235479 213002 235531
rect 232342 235479 232394 235531
rect 238006 235479 238058 235531
rect 285910 235479 285962 235531
rect 299830 235479 299882 235531
rect 354262 235479 354314 235531
rect 394966 235479 395018 235531
rect 587350 235479 587402 235531
rect 211990 235405 212042 235457
rect 233014 235405 233066 235457
rect 242134 235405 242186 235457
rect 293398 235405 293450 235457
rect 294838 235405 294890 235457
rect 337654 235405 337706 235457
rect 339478 235405 339530 235457
rect 395062 235405 395114 235457
rect 396790 235405 396842 235457
rect 587638 235405 587690 235457
rect 206998 235331 207050 235383
rect 221782 235331 221834 235383
rect 223894 235331 223946 235383
rect 244726 235331 244778 235383
rect 249718 235331 249770 235383
rect 302326 235331 302378 235383
rect 304822 235331 304874 235383
rect 362614 235331 362666 235383
rect 393430 235331 393482 235383
rect 587062 235331 587114 235383
rect 214198 235257 214250 235309
rect 235318 235257 235370 235309
rect 288886 235257 288938 235309
rect 346870 235257 346922 235309
rect 392182 235257 392234 235309
rect 585526 235257 585578 235309
rect 209302 235183 209354 235235
rect 228502 235183 228554 235235
rect 229750 235183 229802 235235
rect 253558 235183 253610 235235
rect 257494 235183 257546 235235
rect 308182 235183 308234 235235
rect 334966 235183 335018 235235
rect 391702 235183 391754 235235
rect 396310 235183 396362 235235
rect 588598 235183 588650 235235
rect 211606 235109 211658 235161
rect 230710 235109 230762 235161
rect 232918 235109 232970 235161
rect 262006 235109 262058 235161
rect 266134 235109 266186 235161
rect 324214 235109 324266 235161
rect 332182 235109 332234 235161
rect 385366 235109 385418 235161
rect 387670 235109 387722 235161
rect 583414 235109 583466 235161
rect 207862 235035 207914 235087
rect 215926 235035 215978 235087
rect 220630 235035 220682 235087
rect 241846 235035 241898 235087
rect 246646 235035 246698 235087
rect 299254 235035 299306 235087
rect 309334 235035 309386 235087
rect 368854 235035 368906 235087
rect 394870 235035 394922 235087
rect 596086 235035 596138 235087
rect 211030 234961 211082 235013
rect 231574 234961 231626 235013
rect 243862 234961 243914 235013
rect 296470 234961 296522 235013
rect 298006 234961 298058 235013
rect 362422 234961 362474 235013
rect 362518 234961 362570 235013
rect 394678 234961 394730 235013
rect 398998 234961 399050 235013
rect 605974 234961 606026 235013
rect 213430 234887 213482 234939
rect 208726 234813 208778 234865
rect 224758 234813 224810 234865
rect 204406 234739 204458 234791
rect 215830 234739 215882 234791
rect 235702 234887 235754 234939
rect 266902 234887 266954 234939
rect 268918 234887 268970 234939
rect 331414 234887 331466 234939
rect 333430 234887 333482 234939
rect 394774 234887 394826 234939
rect 398614 234887 398666 234939
rect 605302 234887 605354 234939
rect 225526 234813 225578 234865
rect 260182 234813 260234 234865
rect 260278 234813 260330 234865
rect 323062 234813 323114 234865
rect 327670 234813 327722 234865
rect 392470 234813 392522 234865
rect 403606 234813 403658 234865
rect 615862 234813 615914 234865
rect 236086 234739 236138 234791
rect 254230 234739 254282 234791
rect 306646 234739 306698 234791
rect 321622 234739 321674 234791
rect 387286 234739 387338 234791
rect 406678 234739 406730 234791
rect 621814 234739 621866 234791
rect 202870 234665 202922 234717
rect 214870 234665 214922 234717
rect 225142 234665 225194 234717
rect 247702 234665 247754 234717
rect 251158 234665 251210 234717
rect 304150 234665 304202 234717
rect 315286 234665 315338 234717
rect 394678 234665 394730 234717
rect 408118 234665 408170 234717
rect 624886 234665 624938 234717
rect 204790 234591 204842 234643
rect 202006 234517 202058 234569
rect 213430 234517 213482 234569
rect 203254 234443 203306 234495
rect 207766 234443 207818 234495
rect 206134 234369 206186 234421
rect 222358 234591 222410 234643
rect 240214 234591 240266 234643
rect 264694 234591 264746 234643
rect 267478 234591 267530 234643
rect 285046 234591 285098 234643
rect 286678 234591 286730 234643
rect 326806 234591 326858 234643
rect 329302 234591 329354 234643
rect 449302 234591 449354 234643
rect 243958 234517 244010 234569
rect 215926 234443 215978 234495
rect 225526 234443 225578 234495
rect 235606 234443 235658 234495
rect 250582 234517 250634 234569
rect 255286 234517 255338 234569
rect 278230 234517 278282 234569
rect 283894 234517 283946 234569
rect 320662 234517 320714 234569
rect 323542 234517 323594 234569
rect 434902 234517 434954 234569
rect 250486 234443 250538 234495
rect 267958 234443 268010 234495
rect 273046 234443 273098 234495
rect 304726 234443 304778 234495
rect 206518 234295 206570 234347
rect 219382 234369 219434 234421
rect 237046 234369 237098 234421
rect 258070 234369 258122 234421
rect 262486 234369 262538 234421
rect 290902 234369 290954 234421
rect 292918 234369 292970 234421
rect 313846 234443 313898 234495
rect 314422 234443 314474 234495
rect 426166 234443 426218 234495
rect 312694 234369 312746 234421
rect 407446 234369 407498 234421
rect 408982 234369 409034 234421
rect 410614 234369 410666 234421
rect 200278 234221 200330 234273
rect 210358 234221 210410 234273
rect 221014 234295 221066 234347
rect 239830 234295 239882 234347
rect 260470 234295 260522 234347
rect 271606 234295 271658 234347
rect 302230 234295 302282 234347
rect 308470 234295 308522 234347
rect 414742 234295 414794 234347
rect 222454 234221 222506 234273
rect 242902 234221 242954 234273
rect 260758 234221 260810 234273
rect 261238 234221 261290 234273
rect 288022 234221 288074 234273
rect 295222 234221 295274 234273
rect 348694 234221 348746 234273
rect 352150 234221 352202 234273
rect 401110 234221 401162 234273
rect 407254 234221 407306 234273
rect 503926 234221 503978 234273
rect 200182 234147 200234 234199
rect 208822 234147 208874 234199
rect 256534 234147 256586 234199
rect 278038 234147 278090 234199
rect 283990 234147 284042 234199
rect 311254 234147 311306 234199
rect 318358 234147 318410 234199
rect 371638 234147 371690 234199
rect 378550 234147 378602 234199
rect 399190 234147 399242 234199
rect 403510 234147 403562 234199
rect 495382 234147 495434 234199
rect 198742 234073 198794 234125
rect 207382 234073 207434 234125
rect 207766 234073 207818 234125
rect 216502 234073 216554 234125
rect 244342 234073 244394 234125
rect 263830 234073 263882 234125
rect 268534 234073 268586 234125
rect 293782 234073 293834 234125
rect 295702 234073 295754 234125
rect 341206 234073 341258 234125
rect 345910 234073 345962 234125
rect 400150 234073 400202 234125
rect 401782 234073 401834 234125
rect 484630 234073 484682 234125
rect 198358 233999 198410 234051
rect 205942 233999 205994 234051
rect 197494 233925 197546 233977
rect 204310 233925 204362 233977
rect 205558 233925 205610 233977
rect 218710 233999 218762 234051
rect 247414 233999 247466 234051
rect 266326 233999 266378 234051
rect 267094 233999 267146 234051
rect 290998 233999 291050 234051
rect 301654 233999 301706 234051
rect 344086 233999 344138 234051
rect 344374 233999 344426 234051
rect 394870 233999 394922 234051
rect 396694 233999 396746 234051
rect 475222 233999 475274 234051
rect 206902 233925 206954 233977
rect 220246 233925 220298 233977
rect 259798 233925 259850 233977
rect 281494 233925 281546 233977
rect 305206 233925 305258 233977
rect 351382 233925 351434 233977
rect 361270 233925 361322 233977
rect 432022 233925 432074 233977
rect 199126 233851 199178 233903
rect 205078 233851 205130 233903
rect 205174 233851 205226 233903
rect 196918 233777 196970 233829
rect 202870 233777 202922 233829
rect 204214 233777 204266 233829
rect 215542 233777 215594 233829
rect 196534 233703 196586 233755
rect 200566 233703 200618 233755
rect 201526 233703 201578 233755
rect 211894 233703 211946 233755
rect 195670 233629 195722 233681
rect 201334 233629 201386 233681
rect 202486 233629 202538 233681
rect 212566 233629 212618 233681
rect 258358 233851 258410 233903
rect 278710 233851 278762 233903
rect 296086 233851 296138 233903
rect 339766 233851 339818 233903
rect 370294 233851 370346 233903
rect 427894 233851 427946 233903
rect 215830 233777 215882 233829
rect 217942 233777 217994 233829
rect 253462 233777 253514 233829
rect 270838 233777 270890 233829
rect 294454 233777 294506 233829
rect 331222 233777 331274 233829
rect 354934 233777 354986 233829
rect 285142 233703 285194 233755
rect 323158 233703 323210 233755
rect 338038 233703 338090 233755
rect 386230 233703 386282 233755
rect 398230 233777 398282 233829
rect 405814 233777 405866 233829
rect 407446 233777 407498 233829
rect 423286 233777 423338 233829
rect 407542 233703 407594 233755
rect 217174 233629 217226 233681
rect 306262 233629 306314 233681
rect 344470 233629 344522 233681
rect 363478 233629 363530 233681
rect 364150 233629 364202 233681
rect 383638 233629 383690 233681
rect 408118 233629 408170 233681
rect 192886 233555 192938 233607
rect 195286 233555 195338 233607
rect 195574 233555 195626 233607
rect 199798 233555 199850 233607
rect 201046 233555 201098 233607
rect 209686 233555 209738 233607
rect 228406 233555 228458 233607
rect 238102 233555 238154 233607
rect 259894 233555 259946 233607
rect 267766 233555 267818 233607
rect 302902 233555 302954 233607
rect 337366 233555 337418 233607
rect 348886 233555 348938 233607
rect 394582 233555 394634 233607
rect 194230 233481 194282 233533
rect 198358 233481 198410 233533
rect 200662 233481 200714 233533
rect 208150 233481 208202 233533
rect 240598 233481 240650 233533
rect 290422 233481 290474 233533
rect 297238 233481 297290 233533
rect 328342 233481 328394 233533
rect 338614 233481 338666 233533
rect 466486 233481 466538 233533
rect 194614 233407 194666 233459
rect 196054 233407 196106 233459
rect 196150 233407 196202 233459
rect 199126 233407 199178 233459
rect 199702 233407 199754 233459
rect 206614 233407 206666 233459
rect 264406 233407 264458 233459
rect 272854 233407 272906 233459
rect 287446 233407 287498 233459
rect 311158 233407 311210 233459
rect 320278 233407 320330 233459
rect 448246 233407 448298 233459
rect 192406 233333 192458 233385
rect 193750 233333 193802 233385
rect 193846 233333 193898 233385
rect 196822 233333 196874 233385
rect 197974 233333 198026 233385
rect 203638 233333 203690 233385
rect 203926 233333 203978 233385
rect 214198 233333 214250 233385
rect 226678 233333 226730 233385
rect 236758 233333 236810 233385
rect 261622 233333 261674 233385
rect 269014 233333 269066 233385
rect 270454 233333 270506 233385
rect 275062 233333 275114 233385
rect 288406 233333 288458 233385
rect 311062 233333 311114 233385
rect 324790 233333 324842 233385
rect 327766 233333 327818 233385
rect 328534 233333 328586 233385
rect 331126 233333 331178 233385
rect 335350 233333 335402 233385
rect 463606 233333 463658 233385
rect 193462 233259 193514 233311
rect 194614 233259 194666 233311
rect 195190 233259 195242 233311
rect 197494 233259 197546 233311
rect 197878 233259 197930 233311
rect 202102 233259 202154 233311
rect 202390 233259 202442 233311
rect 211126 233259 211178 233311
rect 257974 233259 258026 233311
rect 269494 233259 269546 233311
rect 270262 233259 270314 233311
rect 273526 233259 273578 233311
rect 297142 233259 297194 233311
rect 319414 233259 319466 233311
rect 319894 233259 319946 233311
rect 377302 233259 377354 233311
rect 386326 233259 386378 233311
rect 388726 233259 388778 233311
rect 395926 233259 395978 233311
rect 400246 233259 400298 233311
rect 401206 233259 401258 233311
rect 408886 233259 408938 233311
rect 259126 233185 259178 233237
rect 328150 233185 328202 233237
rect 340822 233185 340874 233237
rect 491254 233185 491306 233237
rect 495382 233185 495434 233237
rect 614998 233185 615050 233237
rect 262102 233111 262154 233163
rect 334198 233111 334250 233163
rect 347062 233111 347114 233163
rect 501046 233111 501098 233163
rect 265750 233037 265802 233089
rect 338038 233037 338090 233089
rect 350326 233037 350378 233089
rect 507094 233037 507146 233089
rect 260662 232963 260714 233015
rect 331318 232963 331370 233015
rect 353110 232963 353162 233015
rect 513142 232963 513194 233015
rect 289942 232889 289994 232941
rect 382870 232889 382922 232941
rect 410038 232889 410090 232941
rect 572086 232889 572138 232941
rect 263926 232815 263978 232867
rect 337270 232815 337322 232867
rect 356278 232815 356330 232867
rect 519190 232815 519242 232867
rect 216598 232741 216650 232793
rect 242134 232741 242186 232793
rect 265174 232741 265226 232793
rect 340246 232741 340298 232793
rect 359062 232741 359114 232793
rect 525238 232741 525290 232793
rect 237622 232667 237674 232719
rect 284374 232667 284426 232719
rect 295318 232667 295370 232719
rect 397366 232667 397418 232719
rect 399190 232667 399242 232719
rect 566710 232667 566762 232719
rect 218038 232593 218090 232645
rect 245110 232593 245162 232645
rect 268438 232593 268490 232645
rect 346294 232593 346346 232645
rect 219766 232519 219818 232571
rect 248086 232519 248138 232571
rect 266614 232519 266666 232571
rect 343222 232519 343274 232571
rect 221110 232445 221162 232497
rect 251158 232445 251210 232497
rect 271222 232445 271274 232497
rect 352342 232593 352394 232645
rect 362134 232593 362186 232645
rect 531286 232593 531338 232645
rect 222550 232371 222602 232423
rect 254230 232371 254282 232423
rect 274870 232371 274922 232423
rect 356086 232519 356138 232571
rect 365398 232519 365450 232571
rect 537238 232519 537290 232571
rect 366262 232445 366314 232497
rect 542614 232445 542666 232497
rect 222934 232297 222986 232349
rect 255670 232297 255722 232349
rect 269686 232297 269738 232349
rect 349366 232371 349418 232423
rect 365014 232371 365066 232423
rect 539542 232371 539594 232423
rect 346966 232297 347018 232349
rect 361366 232297 361418 232349
rect 368182 232297 368234 232349
rect 543382 232297 543434 232349
rect 224278 232223 224330 232275
rect 257206 232223 257258 232275
rect 274198 232223 274250 232275
rect 358294 232223 358346 232275
rect 369526 232223 369578 232275
rect 548566 232223 548618 232275
rect 226294 232149 226346 232201
rect 261718 232149 261770 232201
rect 272950 232149 273002 232201
rect 355318 232149 355370 232201
rect 368086 232149 368138 232201
rect 545590 232149 545642 232201
rect 227062 232075 227114 232127
rect 263254 232075 263306 232127
rect 277462 232075 277514 232127
rect 364438 232075 364490 232127
rect 372694 232075 372746 232127
rect 552406 232075 552458 232127
rect 233878 232001 233930 232053
rect 274486 232001 274538 232053
rect 275734 232001 275786 232053
rect 346966 232001 347018 232053
rect 354262 232001 354314 232053
rect 367126 232001 367178 232053
rect 372310 232001 372362 232053
rect 554710 232001 554762 232053
rect 234838 231927 234890 231979
rect 278326 231927 278378 231979
rect 278998 231927 279050 231979
rect 367414 231927 367466 231979
rect 375766 231927 375818 231979
rect 558454 231927 558506 231979
rect 233206 231853 233258 231905
rect 275350 231853 275402 231905
rect 280246 231853 280298 231905
rect 370390 231853 370442 231905
rect 374518 231853 374570 231905
rect 557014 231853 557066 231905
rect 235990 231779 236042 231831
rect 281302 231779 281354 231831
rect 281974 231779 282026 231831
rect 373462 231779 373514 231831
rect 378934 231779 378986 231831
rect 564502 231779 564554 231831
rect 258742 231705 258794 231757
rect 326710 231705 326762 231757
rect 337558 231705 337610 231757
rect 485206 231705 485258 231757
rect 255766 231631 255818 231683
rect 320566 231631 320618 231683
rect 334870 231631 334922 231683
rect 479158 231631 479210 231683
rect 257590 231557 257642 231609
rect 325174 231557 325226 231609
rect 327094 231557 327146 231609
rect 464086 231557 464138 231609
rect 248374 231483 248426 231535
rect 305494 231483 305546 231535
rect 312214 231483 312266 231535
rect 433846 231483 433898 231535
rect 281206 231409 281258 231461
rect 289654 231409 289706 231461
rect 290806 231409 290858 231461
rect 374614 231409 374666 231461
rect 403126 231409 403178 231461
rect 520726 231409 520778 231461
rect 292534 231335 292586 231387
rect 379990 231335 380042 231387
rect 400150 231335 400202 231387
rect 499606 231335 499658 231387
rect 245206 231261 245258 231313
rect 299446 231261 299498 231313
rect 300214 231261 300266 231313
rect 385846 231261 385898 231313
rect 395062 231261 395114 231313
rect 485974 231261 486026 231313
rect 293494 231187 293546 231239
rect 365110 231187 365162 231239
rect 394774 231187 394826 231239
rect 473878 231187 473930 231239
rect 256150 231113 256202 231165
rect 322102 231113 322154 231165
rect 337366 231113 337418 231165
rect 252982 231039 253034 231091
rect 314518 231039 314570 231091
rect 344470 231039 344522 231091
rect 290614 230965 290666 231017
rect 297430 230965 297482 231017
rect 308182 230965 308234 231017
rect 323638 230965 323690 231017
rect 328342 230965 328394 231017
rect 401398 230965 401450 231017
rect 323062 230891 323114 230943
rect 329590 230891 329642 230943
rect 331222 230891 331274 230943
rect 395350 230891 395402 230943
rect 414742 231113 414794 231165
rect 424054 231113 424106 231165
rect 415702 230965 415754 231017
rect 419542 230891 419594 230943
rect 282550 230817 282602 230869
rect 300598 230817 300650 230869
rect 326806 230817 326858 230869
rect 380182 230817 380234 230869
rect 387286 230817 387338 230869
rect 449686 230817 449738 230869
rect 319606 230743 319658 230795
rect 365014 230743 365066 230795
rect 367126 230743 367178 230795
rect 409654 230743 409706 230795
rect 313942 230669 313994 230721
rect 362134 230669 362186 230721
rect 362614 230669 362666 230721
rect 416470 230669 416522 230721
rect 302326 230595 302378 230647
rect 308566 230595 308618 230647
rect 320662 230595 320714 230647
rect 374230 230595 374282 230647
rect 306646 230521 306698 230573
rect 317590 230521 317642 230573
rect 323158 230521 323210 230573
rect 377110 230521 377162 230573
rect 147478 230447 147530 230499
rect 154102 230447 154154 230499
rect 299254 230447 299306 230499
rect 302518 230447 302570 230499
rect 304150 230447 304202 230499
rect 311638 230447 311690 230499
rect 320854 230447 320906 230499
rect 368182 230447 368234 230499
rect 426166 230447 426218 230499
rect 436150 230447 436202 230499
rect 246166 230373 246218 230425
rect 298678 230373 298730 230425
rect 313462 230373 313514 230425
rect 436918 230373 436970 230425
rect 241078 230299 241130 230351
rect 291958 230299 292010 230351
rect 314902 230299 314954 230351
rect 439990 230299 440042 230351
rect 245782 230225 245834 230277
rect 300982 230225 301034 230277
rect 317974 230225 318026 230277
rect 445942 230225 445994 230277
rect 248950 230151 249002 230203
rect 304822 230151 304874 230203
rect 321238 230151 321290 230203
rect 451990 230225 452042 230277
rect 449302 230151 449354 230203
rect 466390 230151 466442 230203
rect 251926 230077 251978 230129
rect 310774 230077 310826 230129
rect 325750 230077 325802 230129
rect 461014 230077 461066 230129
rect 463606 230077 463658 230129
rect 478390 230077 478442 230129
rect 248758 230003 248810 230055
rect 307030 230003 307082 230055
rect 324022 230003 324074 230055
rect 458038 230003 458090 230055
rect 466486 230003 466538 230055
rect 484438 230003 484490 230055
rect 503926 230003 503978 230055
rect 622678 230003 622730 230055
rect 227446 229929 227498 229981
rect 264790 229929 264842 229981
rect 290902 229929 290954 229981
rect 331894 229929 331946 229981
rect 434902 229929 434954 229981
rect 454294 229929 454346 229981
rect 475222 229929 475274 229981
rect 601462 229929 601514 229981
rect 250198 229855 250250 229907
rect 310006 229855 310058 229907
rect 331606 229855 331658 229907
rect 473110 229855 473162 229907
rect 480886 229855 480938 229907
rect 609046 229855 609098 229907
rect 147094 229781 147146 229833
rect 151414 229781 151466 229833
rect 251542 229781 251594 229833
rect 313078 229781 313130 229833
rect 336310 229781 336362 229833
rect 482134 229781 482186 229833
rect 484630 229781 484682 229833
rect 612118 229781 612170 229833
rect 254806 229707 254858 229759
rect 319126 229707 319178 229759
rect 348502 229707 348554 229759
rect 504022 229707 504074 229759
rect 215254 229633 215306 229685
rect 239062 229633 239114 229685
rect 244246 229633 244298 229685
rect 298006 229633 298058 229685
rect 298390 229633 298442 229685
rect 406774 229633 406826 229685
rect 409846 229633 409898 229685
rect 565942 229633 565994 229685
rect 220150 229559 220202 229611
rect 249718 229559 249770 229611
rect 253078 229559 253130 229611
rect 316150 229559 316202 229611
rect 351766 229559 351818 229611
rect 510166 229559 510218 229611
rect 221590 229485 221642 229537
rect 252598 229485 252650 229537
rect 255190 229485 255242 229537
rect 316822 229485 316874 229537
rect 354838 229485 354890 229537
rect 516118 229485 516170 229537
rect 264310 229411 264362 229463
rect 334966 229411 335018 229463
rect 357622 229411 357674 229463
rect 230326 229337 230378 229389
rect 269302 229337 269354 229389
rect 273526 229337 273578 229389
rect 347062 229337 347114 229389
rect 231862 229263 231914 229315
rect 272278 229263 272330 229315
rect 283510 229263 283562 229315
rect 369526 229337 369578 229389
rect 369910 229337 369962 229389
rect 380086 229411 380138 229463
rect 538870 229411 538922 229463
rect 357430 229263 357482 229315
rect 374518 229263 374570 229315
rect 522166 229337 522218 229389
rect 546358 229263 546410 229315
rect 233494 229189 233546 229241
rect 276790 229189 276842 229241
rect 282166 229189 282218 229241
rect 371254 229189 371306 229241
rect 374326 229189 374378 229241
rect 555286 229189 555338 229241
rect 231958 229115 232010 229167
rect 273814 229115 273866 229167
rect 287926 229115 287978 229167
rect 374422 229115 374474 229167
rect 377206 229115 377258 229167
rect 561430 229115 561482 229167
rect 238390 229041 238442 229093
rect 283606 229041 283658 229093
rect 284758 229041 284810 229093
rect 371542 229041 371594 229093
rect 376822 229041 376874 229093
rect 563638 229041 563690 229093
rect 235222 228967 235274 229019
rect 279862 228967 279914 229019
rect 286294 228967 286346 229019
rect 357430 228967 357482 229019
rect 357526 228967 357578 229019
rect 359926 228967 359978 229019
rect 368950 228967 369002 229019
rect 370486 228967 370538 229019
rect 380470 228967 380522 229019
rect 567478 228967 567530 229019
rect 242518 228893 242570 228945
rect 294934 228893 294986 228945
rect 308950 228893 309002 228945
rect 427798 228893 427850 228945
rect 427894 228893 427946 228945
rect 547894 228893 547946 228945
rect 241654 228819 241706 228871
rect 289750 228819 289802 228871
rect 310678 228819 310730 228871
rect 430870 228819 430922 228871
rect 432022 228819 432074 228871
rect 529750 228819 529802 228871
rect 239734 228745 239786 228797
rect 288886 228745 288938 228797
rect 306166 228745 306218 228797
rect 421846 228745 421898 228797
rect 228886 228671 228938 228723
rect 267862 228671 267914 228723
rect 304438 228671 304490 228723
rect 418774 228671 418826 228723
rect 455062 228671 455114 228723
rect 455734 228671 455786 228723
rect 230614 228597 230666 228649
rect 270742 228597 270794 228649
rect 291478 228597 291530 228649
rect 382966 228597 383018 228649
rect 407542 228597 407594 228649
rect 517654 228597 517706 228649
rect 190198 228523 190250 228575
rect 192310 228523 192362 228575
rect 228790 228523 228842 228575
rect 266230 228523 266282 228575
rect 266326 228523 266378 228575
rect 301750 228523 301802 228575
rect 303478 228523 303530 228575
rect 413494 228523 413546 228575
rect 455158 228523 455210 228575
rect 456502 228523 456554 228575
rect 535798 228523 535850 228575
rect 538006 228523 538058 228575
rect 544342 228523 544394 228575
rect 547126 228523 547178 228575
rect 556150 228523 556202 228575
rect 557686 228523 557738 228575
rect 567382 228523 567434 228575
rect 569014 228523 569066 228575
rect 224374 228449 224426 228501
rect 258742 228449 258794 228501
rect 260470 228449 260522 228501
rect 286678 228449 286730 228501
rect 289366 228449 289418 228501
rect 380086 228449 380138 228501
rect 405334 228449 405386 228501
rect 502582 228449 502634 228501
rect 250582 228375 250634 228427
rect 277558 228375 277610 228427
rect 288022 228375 288074 228427
rect 328918 228375 328970 228427
rect 331126 228375 331178 228427
rect 467062 228375 467114 228427
rect 535798 228375 535850 228427
rect 537910 228375 537962 228427
rect 260758 228301 260810 228353
rect 292630 228301 292682 228353
rect 293878 228301 293930 228353
rect 380278 228301 380330 228353
rect 391702 228301 391754 228353
rect 476950 228301 477002 228353
rect 270838 228227 270890 228279
rect 313846 228227 313898 228279
rect 313942 228227 313994 228279
rect 392374 228227 392426 228279
rect 392470 228227 392522 228279
rect 461878 228227 461930 228279
rect 267958 228153 268010 228205
rect 307702 228153 307754 228205
rect 311062 228153 311114 228205
rect 383254 228153 383306 228205
rect 394678 228153 394730 228205
rect 437686 228153 437738 228205
rect 269494 228079 269546 228131
rect 322966 228079 323018 228131
rect 344086 228079 344138 228131
rect 412726 228079 412778 228131
rect 258070 228005 258122 228057
rect 280630 228005 280682 228057
rect 290998 228005 291050 228057
rect 341014 228005 341066 228057
rect 341206 228005 341258 228057
rect 398326 228005 398378 228057
rect 263830 227931 263882 227983
rect 295702 227931 295754 227983
rect 308278 227931 308330 227983
rect 359158 227931 359210 227983
rect 368854 227931 368906 227983
rect 425590 227931 425642 227983
rect 293782 227857 293834 227909
rect 343990 227857 344042 227909
rect 302230 227783 302282 227835
rect 350038 227783 350090 227835
rect 247030 227709 247082 227761
rect 303958 227709 304010 227761
rect 304726 227709 304778 227761
rect 353110 227709 353162 227761
rect 387766 227709 387818 227761
rect 396214 227709 396266 227761
rect 281494 227635 281546 227687
rect 325846 227635 325898 227687
rect 149398 227561 149450 227613
rect 177142 227561 177194 227613
rect 278038 227561 278090 227613
rect 319894 227561 319946 227613
rect 319990 227561 320042 227613
rect 403702 227561 403754 227613
rect 423286 227561 423338 227613
rect 433174 227561 433226 227613
rect 187126 227487 187178 227539
rect 190774 227487 190826 227539
rect 216118 227487 216170 227539
rect 239830 227487 239882 227539
rect 249334 227487 249386 227539
rect 306262 227487 306314 227539
rect 311254 227487 311306 227539
rect 375766 227487 375818 227539
rect 389494 227487 389546 227539
rect 587158 227487 587210 227539
rect 590710 227487 590762 227539
rect 594646 227487 594698 227539
rect 629302 227487 629354 227539
rect 634006 227487 634058 227539
rect 213046 227413 213098 227465
rect 233782 227413 233834 227465
rect 238774 227413 238826 227465
rect 252214 227413 252266 227465
rect 253846 227413 253898 227465
rect 315382 227413 315434 227465
rect 318166 227413 318218 227465
rect 381814 227413 381866 227465
rect 390454 227413 390506 227465
rect 217462 227339 217514 227391
rect 241270 227339 241322 227391
rect 244726 227339 244778 227391
rect 254902 227339 254954 227391
rect 311158 227339 311210 227391
rect 384022 227339 384074 227391
rect 388534 227339 388586 227391
rect 585622 227339 585674 227391
rect 588598 227413 588650 227465
rect 600790 227413 600842 227465
rect 606358 227413 606410 227465
rect 638518 227413 638570 227465
rect 589366 227339 589418 227391
rect 219478 227265 219530 227317
rect 245878 227265 245930 227317
rect 275062 227265 275114 227317
rect 348598 227265 348650 227317
rect 388918 227265 388970 227317
rect 586390 227265 586442 227317
rect 588790 227265 588842 227317
rect 626422 227265 626474 227317
rect 217846 227191 217898 227243
rect 242902 227191 242954 227243
rect 271990 227191 272042 227243
rect 351574 227191 351626 227243
rect 398902 227191 398954 227243
rect 584854 227191 584906 227243
rect 587446 227191 587498 227243
rect 630166 227191 630218 227243
rect 220342 227117 220394 227169
rect 247414 227117 247466 227169
rect 264694 227117 264746 227169
rect 288118 227117 288170 227169
rect 289654 227117 289706 227169
rect 369622 227117 369674 227169
rect 390070 227117 390122 227169
rect 588598 227117 588650 227169
rect 590902 227117 590954 227169
rect 630934 227117 630986 227169
rect 215734 227043 215786 227095
rect 238390 227043 238442 227095
rect 276694 227043 276746 227095
rect 360598 227043 360650 227095
rect 390838 227043 390890 227095
rect 590134 227043 590186 227095
rect 590422 227043 590474 227095
rect 632374 227043 632426 227095
rect 238102 226969 238154 227021
rect 264022 226969 264074 227021
rect 275254 226969 275306 227021
rect 357622 226969 357674 227021
rect 359830 226969 359882 227021
rect 221686 226895 221738 226947
rect 250390 226895 250442 226947
rect 253558 226895 253610 226947
rect 266998 226895 267050 226947
rect 273430 226895 273482 226947
rect 354550 226895 354602 226947
rect 354646 226895 354698 226947
rect 392182 226895 392234 226947
rect 392662 226969 392714 227021
rect 593974 226969 594026 227021
rect 599158 226969 599210 227021
rect 603382 226969 603434 227021
rect 636886 226969 636938 227021
rect 393142 226895 393194 226947
rect 587350 226895 587402 226947
rect 598486 226895 598538 226947
rect 633142 226895 633194 226947
rect 224950 226821 225002 226873
rect 256438 226821 256490 226873
rect 324214 226821 324266 226873
rect 339478 226821 339530 226873
rect 365110 226821 365162 226873
rect 223318 226747 223370 226799
rect 253462 226747 253514 226799
rect 279766 226747 279818 226799
rect 298198 226747 298250 226799
rect 298390 226747 298442 226799
rect 366742 226747 366794 226799
rect 226582 226673 226634 226725
rect 259414 226673 259466 226725
rect 284662 226673 284714 226725
rect 298102 226673 298154 226725
rect 300598 226673 300650 226725
rect 372694 226747 372746 226799
rect 374614 226747 374666 226799
rect 391510 226747 391562 226799
rect 395542 226821 395594 226873
rect 599158 226821 599210 226873
rect 600406 226821 600458 226873
rect 634678 226821 634730 226873
rect 396118 226747 396170 226799
rect 400822 226747 400874 226799
rect 419158 226747 419210 226799
rect 419254 226747 419306 226799
rect 227926 226599 227978 226651
rect 262486 226599 262538 226651
rect 264886 226599 264938 226651
rect 276118 226599 276170 226651
rect 285718 226599 285770 226651
rect 378742 226673 378794 226725
rect 380278 226673 380330 226725
rect 397654 226673 397706 226725
rect 402166 226673 402218 226725
rect 418870 226673 418922 226725
rect 374422 226599 374474 226651
rect 385558 226599 385610 226651
rect 397174 226599 397226 226651
rect 587638 226673 587690 226725
rect 602230 226673 602282 226725
rect 603286 226747 603338 226799
rect 637750 226747 637802 226799
rect 603670 226673 603722 226725
rect 606262 226673 606314 226725
rect 639190 226673 639242 226725
rect 602998 226599 603050 226651
rect 606166 226599 606218 226651
rect 639958 226599 640010 226651
rect 229558 226525 229610 226577
rect 265558 226525 265610 226577
rect 271030 226525 271082 226577
rect 294262 226525 294314 226577
rect 297430 226525 297482 226577
rect 390070 226525 390122 226577
rect 392182 226525 392234 226577
rect 231094 226451 231146 226503
rect 268534 226451 268586 226503
rect 288502 226451 288554 226503
rect 384790 226451 384842 226503
rect 385750 226451 385802 226503
rect 398806 226451 398858 226503
rect 232534 226377 232586 226429
rect 271606 226377 271658 226429
rect 272854 226377 272906 226429
rect 282550 226377 282602 226429
rect 298102 226377 298154 226429
rect 378070 226377 378122 226429
rect 379894 226377 379946 226429
rect 387766 226377 387818 226429
rect 388150 226377 388202 226429
rect 398902 226377 398954 226429
rect 402550 226525 402602 226577
rect 404950 226451 405002 226503
rect 408214 226377 408266 226429
rect 213814 226303 213866 226355
rect 237526 226303 237578 226355
rect 244822 226303 244874 226355
rect 147094 226229 147146 226281
rect 151318 226229 151370 226281
rect 217078 226229 217130 226281
rect 243574 226229 243626 226281
rect 246550 226229 246602 226281
rect 252214 226303 252266 226355
rect 285142 226303 285194 226355
rect 291574 226303 291626 226355
rect 390838 226303 390890 226355
rect 42262 226155 42314 226207
rect 45814 226155 45866 226207
rect 215638 226155 215690 226207
rect 240598 226155 240650 226207
rect 243958 226155 244010 226207
rect 251926 226155 251978 226207
rect 151126 226081 151178 226133
rect 187126 226081 187178 226133
rect 218326 226081 218378 226133
rect 246646 226081 246698 226133
rect 297238 226229 297290 226281
rect 297622 226229 297674 226281
rect 402838 226303 402890 226355
rect 408022 226303 408074 226355
rect 419158 226525 419210 226577
rect 609814 226525 609866 226577
rect 419062 226451 419114 226503
rect 612790 226451 612842 226503
rect 613558 226377 613610 226429
rect 629206 226377 629258 226429
rect 635446 226377 635498 226429
rect 397846 226229 397898 226281
rect 400246 226229 400298 226281
rect 618070 226303 618122 226355
rect 624118 226229 624170 226281
rect 252118 226155 252170 226207
rect 291190 226155 291242 226207
rect 301270 226155 301322 226207
rect 300214 226081 300266 226133
rect 300694 226081 300746 226133
rect 408982 226081 409034 226133
rect 410422 226155 410474 226207
rect 629398 226155 629450 226207
rect 411286 226081 411338 226133
rect 411670 226081 411722 226133
rect 631702 226081 631754 226133
rect 214582 226007 214634 226059
rect 236854 226007 236906 226059
rect 241846 226007 241898 226059
rect 248854 226007 248906 226059
rect 257110 226007 257162 226059
rect 212374 225933 212426 225985
rect 234550 225933 234602 225985
rect 236758 225933 236810 225985
rect 261046 225933 261098 225985
rect 266902 226007 266954 226059
rect 279094 226007 279146 226059
rect 282550 226007 282602 226059
rect 336406 226007 336458 226059
rect 321334 225933 321386 225985
rect 334102 225933 334154 225985
rect 379894 226007 379946 226059
rect 379990 226007 380042 226059
rect 394582 226007 394634 226059
rect 398806 226007 398858 226059
rect 579574 226007 579626 226059
rect 584566 226007 584618 226059
rect 628630 226007 628682 226059
rect 218806 225859 218858 225911
rect 244342 225859 244394 225911
rect 262006 225859 262058 225911
rect 273046 225859 273098 225911
rect 241750 225785 241802 225837
rect 252118 225785 252170 225837
rect 267766 225785 267818 225837
rect 278422 225785 278474 225837
rect 247702 225711 247754 225763
rect 257974 225711 258026 225763
rect 269014 225711 269066 225763
rect 330454 225859 330506 225911
rect 331414 225859 331466 225911
rect 345526 225859 345578 225911
rect 346870 225859 346922 225911
rect 278614 225785 278666 225837
rect 327382 225785 327434 225837
rect 374518 225785 374570 225837
rect 382582 225785 382634 225837
rect 382966 225933 383018 225985
rect 388630 225933 388682 225985
rect 388726 225933 388778 225985
rect 386998 225859 387050 225911
rect 387382 225859 387434 225911
rect 398710 225859 398762 225911
rect 385846 225785 385898 225837
rect 398614 225785 398666 225837
rect 398902 225933 398954 225985
rect 582646 225933 582698 225985
rect 603478 225933 603530 225985
rect 636214 225933 636266 225985
rect 400246 225859 400298 225911
rect 419254 225859 419306 225911
rect 581110 225785 581162 225837
rect 591478 225785 591530 225837
rect 285046 225711 285098 225763
rect 342550 225711 342602 225763
rect 365686 225711 365738 225763
rect 393814 225711 393866 225763
rect 396214 225711 396266 225763
rect 584086 225711 584138 225763
rect 587062 225711 587114 225763
rect 595414 225711 595466 225763
rect 627862 225711 627914 225763
rect 278230 225637 278282 225689
rect 318358 225637 318410 225689
rect 321718 225637 321770 225689
rect 451222 225637 451274 225689
rect 273718 225563 273770 225615
rect 309334 225563 309386 225615
rect 315766 225563 315818 225615
rect 439126 225563 439178 225615
rect 273622 225489 273674 225541
rect 303190 225489 303242 225541
rect 309910 225489 309962 225541
rect 427030 225489 427082 225541
rect 585526 225489 585578 225541
rect 592342 225489 592394 225541
rect 259030 225415 259082 225467
rect 269974 225415 270026 225467
rect 306742 225415 306794 225467
rect 420982 225415 421034 225467
rect 303862 225341 303914 225393
rect 415030 225341 415082 225393
rect 302134 225267 302186 225319
rect 411958 225267 412010 225319
rect 278710 225193 278762 225245
rect 324406 225193 324458 225245
rect 351382 225193 351434 225245
rect 418006 225193 418058 225245
rect 305110 225119 305162 225171
rect 333526 225119 333578 225171
rect 339766 225119 339818 225171
rect 399958 225119 400010 225171
rect 408886 225119 408938 225171
rect 610486 225119 610538 225171
rect 252694 225045 252746 225097
rect 312310 225045 312362 225097
rect 337654 225045 337706 225097
rect 396886 225045 396938 225097
rect 398614 225045 398666 225097
rect 348694 224971 348746 225023
rect 399094 224971 399146 225023
rect 399382 225045 399434 225097
rect 606742 225045 606794 225097
rect 407446 224971 407498 225023
rect 369430 224897 369482 224949
rect 405142 224897 405194 224949
rect 149494 224823 149546 224875
rect 174166 224823 174218 224875
rect 362806 224823 362858 224875
rect 402166 224823 402218 224875
rect 149398 224749 149450 224801
rect 159862 224749 159914 224801
rect 277942 224749 277994 224801
rect 363670 224749 363722 224801
rect 371542 224749 371594 224801
rect 379510 224749 379562 224801
rect 380086 224749 380138 224801
rect 388630 224749 388682 224801
rect 388726 224749 388778 224801
rect 389302 224749 389354 224801
rect 392278 224749 392330 224801
rect 268630 224675 268682 224727
rect 282070 224675 282122 224727
rect 362422 224675 362474 224727
rect 369430 224675 369482 224727
rect 369526 224675 369578 224727
rect 376438 224675 376490 224727
rect 382870 224675 382922 224727
rect 386326 224675 386378 224727
rect 397462 224675 397514 224727
rect 400630 224675 400682 224727
rect 593110 224675 593162 224727
rect 596086 224675 596138 224727
rect 597718 224675 597770 224727
rect 316342 224601 316394 224653
rect 441430 224601 441482 224653
rect 319318 224527 319370 224579
rect 447478 224527 447530 224579
rect 323254 224453 323306 224505
rect 452758 224453 452810 224505
rect 322294 224379 322346 224431
rect 453430 224379 453482 224431
rect 325270 224305 325322 224357
rect 459574 224305 459626 224357
rect 328246 224231 328298 224283
rect 465622 224231 465674 224283
rect 331510 224157 331562 224209
rect 471574 224157 471626 224209
rect 553270 224157 553322 224209
rect 555382 224157 555434 224209
rect 330742 224083 330794 224135
rect 467830 224083 467882 224135
rect 334486 224009 334538 224061
rect 477622 224009 477674 224061
rect 337174 223935 337226 223987
rect 483766 223935 483818 223987
rect 340438 223861 340490 223913
rect 489718 223861 489770 223913
rect 343606 223787 343658 223839
rect 497302 223787 497354 223839
rect 261910 223713 261962 223765
rect 332662 223713 332714 223765
rect 346582 223713 346634 223765
rect 501814 223713 501866 223765
rect 263542 223639 263594 223691
rect 335734 223639 335786 223691
rect 349558 223639 349610 223691
rect 507862 223639 507914 223691
rect 268054 223565 268106 223617
rect 344854 223565 344906 223617
rect 348022 223565 348074 223617
rect 504790 223565 504842 223617
rect 266518 223491 266570 223543
rect 341782 223491 341834 223543
rect 348118 223491 348170 223543
rect 506326 223491 506378 223543
rect 264598 223417 264650 223469
rect 338710 223417 338762 223469
rect 351094 223417 351146 223469
rect 510838 223417 510890 223469
rect 270934 223343 270986 223395
rect 350806 223343 350858 223395
rect 352534 223343 352586 223395
rect 513910 223343 513962 223395
rect 269398 223269 269450 223321
rect 347734 223269 347786 223321
rect 351190 223269 351242 223321
rect 512374 223269 512426 223321
rect 272566 223195 272618 223247
rect 353878 223195 353930 223247
rect 354070 223195 354122 223247
rect 516982 223195 517034 223247
rect 313366 223121 313418 223173
rect 435382 223121 435434 223173
rect 310294 223047 310346 223099
rect 429334 223047 429386 223099
rect 307222 222973 307274 223025
rect 423286 222973 423338 223025
rect 312598 222899 312650 222951
rect 431542 222899 431594 222951
rect 307990 222825 308042 222877
rect 422518 222825 422570 222877
rect 304246 222751 304298 222803
rect 417238 222751 417290 222803
rect 286198 222677 286250 222729
rect 381046 222677 381098 222729
rect 401110 222677 401162 222729
rect 511606 222677 511658 222729
rect 302806 222603 302858 222655
rect 414262 222603 414314 222655
rect 301942 222529 301994 222581
rect 410518 222529 410570 222581
rect 410614 222529 410666 222581
rect 430102 222529 430154 222581
rect 281590 222455 281642 222507
rect 371926 222455 371978 222507
rect 394870 222455 394922 222507
rect 496534 222455 496586 222507
rect 283126 222381 283178 222433
rect 374998 222381 375050 222433
rect 386230 222381 386282 222433
rect 482902 222381 482954 222433
rect 274102 222307 274154 222359
rect 356854 222307 356906 222359
rect 371638 222307 371690 222359
rect 443734 222307 443786 222359
rect 149398 221863 149450 221915
rect 171382 221863 171434 221915
rect 149494 221789 149546 221841
rect 182902 221789 182954 221841
rect 145654 221715 145706 221767
rect 184342 221715 184394 221767
rect 478102 221715 478154 221767
rect 479974 221715 480026 221767
rect 512758 221715 512810 221767
rect 515398 221715 515450 221767
rect 655990 219347 656042 219399
rect 676246 219347 676298 219399
rect 655798 219199 655850 219251
rect 676246 219199 676298 219251
rect 149398 219051 149450 219103
rect 162646 219051 162698 219103
rect 655606 219051 655658 219103
rect 676054 219051 676106 219103
rect 149494 218977 149546 219029
rect 168406 218977 168458 219029
rect 149398 218903 149450 218955
rect 180022 218903 180074 218955
rect 143062 218829 143114 218881
rect 184342 218829 184394 218881
rect 147286 217719 147338 217771
rect 151798 217719 151850 217771
rect 149398 216017 149450 216069
rect 177238 216017 177290 216069
rect 41782 213279 41834 213331
rect 45910 213279 45962 213331
rect 149494 213205 149546 213257
rect 159958 213205 160010 213257
rect 674710 213205 674762 213257
rect 676246 213205 676298 213257
rect 149398 213131 149450 213183
rect 174358 213131 174410 213183
rect 675190 213131 675242 213183
rect 676054 213131 676106 213183
rect 41590 212909 41642 212961
rect 45718 212909 45770 212961
rect 146902 212761 146954 212813
rect 151990 212761 152042 212813
rect 41782 212169 41834 212221
rect 45622 212169 45674 212221
rect 41782 211725 41834 211777
rect 43222 211725 43274 211777
rect 41590 211429 41642 211481
rect 44854 211429 44906 211481
rect 147094 210985 147146 211037
rect 151702 210985 151754 211037
rect 41782 210689 41834 210741
rect 50518 210689 50570 210741
rect 147478 210319 147530 210371
rect 151606 210319 151658 210371
rect 674806 210319 674858 210371
rect 676054 210319 676106 210371
rect 674902 210245 674954 210297
rect 676246 210245 676298 210297
rect 41782 210171 41834 210223
rect 46198 210171 46250 210223
rect 41590 209949 41642 210001
rect 50326 209949 50378 210001
rect 41590 209357 41642 209409
rect 46102 209357 46154 209409
rect 147190 207877 147242 207929
rect 151510 207877 151562 207929
rect 646774 207507 646826 207559
rect 679894 207507 679946 207559
rect 674038 207433 674090 207485
rect 675958 207433 676010 207485
rect 146902 207359 146954 207411
rect 151894 207359 151946 207411
rect 674998 207359 675050 207411
rect 676054 207359 676106 207411
rect 146902 206249 146954 206301
rect 152086 206249 152138 206301
rect 185782 205879 185834 205931
rect 186262 205879 186314 205931
rect 674614 205435 674666 205487
rect 674806 205435 674858 205487
rect 149494 204473 149546 204525
rect 165718 204473 165770 204525
rect 149398 204177 149450 204229
rect 157078 204177 157130 204229
rect 147862 202845 147914 202897
rect 154198 202845 154250 202897
rect 675094 202401 675146 202453
rect 675382 202401 675434 202453
rect 41878 201661 41930 201713
rect 44758 201661 44810 201713
rect 149398 201587 149450 201639
rect 182998 201587 183050 201639
rect 41590 201513 41642 201565
rect 44662 201513 44714 201565
rect 143062 201513 143114 201565
rect 184342 201513 184394 201565
rect 674710 201365 674762 201417
rect 675190 201365 675242 201417
rect 41590 200921 41642 200973
rect 44566 200921 44618 200973
rect 149398 200477 149450 200529
rect 160054 200477 160106 200529
rect 674998 199515 675050 199567
rect 675478 199515 675530 199567
rect 147574 199293 147626 199345
rect 152182 199293 152234 199345
rect 181366 198627 181418 198679
rect 184342 198627 184394 198679
rect 660886 198627 660938 198679
rect 675094 198627 675146 198679
rect 178294 198553 178346 198605
rect 184438 198553 184490 198605
rect 674806 198553 674858 198605
rect 675478 198553 675530 198605
rect 674614 198183 674666 198235
rect 675382 198183 675434 198235
rect 674902 197665 674954 197717
rect 675382 197665 675434 197717
rect 41782 197591 41834 197643
rect 41782 197369 41834 197421
rect 147286 195963 147338 196015
rect 171574 195963 171626 196015
rect 149398 195889 149450 195941
rect 174454 195889 174506 195941
rect 149302 195815 149354 195867
rect 180214 195815 180266 195867
rect 166966 195741 167018 195793
rect 184534 195741 184586 195793
rect 169846 195667 169898 195719
rect 184438 195667 184490 195719
rect 172726 195593 172778 195645
rect 184342 195593 184394 195645
rect 674038 194335 674090 194387
rect 675382 194335 675434 194387
rect 149398 193077 149450 193129
rect 165814 193077 165866 193129
rect 149494 193003 149546 193055
rect 168598 193003 168650 193055
rect 152374 192929 152426 192981
rect 184630 192929 184682 192981
rect 155446 192855 155498 192907
rect 184534 192855 184586 192907
rect 158134 192781 158186 192833
rect 184342 192781 184394 192833
rect 163894 192707 163946 192759
rect 184438 192707 184490 192759
rect 149398 190191 149450 190243
rect 157174 190191 157226 190243
rect 149494 190117 149546 190169
rect 162838 190117 162890 190169
rect 143926 190043 143978 190095
rect 184534 190043 184586 190095
rect 149686 189969 149738 190021
rect 184342 189969 184394 190021
rect 171478 189895 171530 189947
rect 184438 189895 184490 189947
rect 174262 189821 174314 189873
rect 184342 189821 184394 189873
rect 147670 189525 147722 189577
rect 154294 189525 154346 189577
rect 145558 187157 145610 187209
rect 184342 187157 184394 187209
rect 162742 187083 162794 187135
rect 184534 187083 184586 187135
rect 168502 187009 168554 187061
rect 184438 187009 184490 187061
rect 180118 186935 180170 186987
rect 185398 186935 185450 186987
rect 156982 184271 157034 184323
rect 184438 184271 184490 184323
rect 165622 184197 165674 184249
rect 184342 184197 184394 184249
rect 179926 184123 179978 184175
rect 184534 184123 184586 184175
rect 645142 183087 645194 183139
rect 649366 183087 649418 183139
rect 149398 182939 149450 182991
rect 185974 182939 186026 182991
rect 149302 182865 149354 182917
rect 186166 182865 186218 182917
rect 42166 182347 42218 182399
rect 45334 182347 45386 182399
rect 149494 181533 149546 181585
rect 177334 181533 177386 181585
rect 149398 181459 149450 181511
rect 183094 181459 183146 181511
rect 154006 181385 154058 181437
rect 184630 181385 184682 181437
rect 156886 181311 156938 181363
rect 184534 181311 184586 181363
rect 165526 181237 165578 181289
rect 184438 181237 184490 181289
rect 171286 181163 171338 181215
rect 184342 181163 184394 181215
rect 149590 179979 149642 180031
rect 185398 179979 185450 180031
rect 645142 179387 645194 179439
rect 649462 179387 649514 179439
rect 149494 178721 149546 178773
rect 162742 178721 162794 178773
rect 149398 178647 149450 178699
rect 168502 178647 168554 178699
rect 149302 178573 149354 178625
rect 171478 178573 171530 178625
rect 159766 178499 159818 178551
rect 184342 178499 184394 178551
rect 182806 178425 182858 178477
rect 184534 178425 184586 178477
rect 177046 178351 177098 178403
rect 184438 178351 184490 178403
rect 149398 175761 149450 175813
rect 156886 175761 156938 175813
rect 149494 175687 149546 175739
rect 165526 175687 165578 175739
rect 145462 175613 145514 175665
rect 184438 175613 184490 175665
rect 145366 175539 145418 175591
rect 184342 175539 184394 175591
rect 645142 174873 645194 174925
rect 649558 174873 649610 174925
rect 147766 174355 147818 174407
rect 154006 174355 154058 174407
rect 149206 174207 149258 174259
rect 186070 174207 186122 174259
rect 655702 173171 655754 173223
rect 676246 173171 676298 173223
rect 655510 173023 655562 173075
rect 676150 173023 676202 173075
rect 655414 172801 655466 172853
rect 676054 172801 676106 172853
rect 148726 172727 148778 172779
rect 184534 172727 184586 172779
rect 148342 172653 148394 172705
rect 184342 172653 184394 172705
rect 148918 172579 148970 172631
rect 184630 172579 184682 172631
rect 148534 172505 148586 172557
rect 184438 172505 184490 172557
rect 645142 171025 645194 171077
rect 649654 171025 649706 171077
rect 672598 169915 672650 169967
rect 673846 169915 673898 169967
rect 676054 169915 676106 169967
rect 148438 169841 148490 169893
rect 184534 169841 184586 169893
rect 148630 169767 148682 169819
rect 184630 169767 184682 169819
rect 148246 169693 148298 169745
rect 184342 169693 184394 169745
rect 151222 169619 151274 169671
rect 184438 169619 184490 169671
rect 673462 169027 673514 169079
rect 676054 169027 676106 169079
rect 645142 168213 645194 168265
rect 649846 168213 649898 168265
rect 149014 166955 149066 167007
rect 184534 166955 184586 167007
rect 148822 166881 148874 166933
rect 184342 166881 184394 166933
rect 149398 166807 149450 166859
rect 184438 166807 184490 166859
rect 151414 164069 151466 164121
rect 184534 164069 184586 164121
rect 154102 163995 154154 164047
rect 184342 163995 184394 164047
rect 174166 163921 174218 163973
rect 184438 163921 184490 163973
rect 177142 163847 177194 163899
rect 184342 163847 184394 163899
rect 645142 163329 645194 163381
rect 649942 163329 649994 163381
rect 646870 161479 646922 161531
rect 676246 161553 676298 161605
rect 647062 161405 647114 161457
rect 676246 161405 676298 161457
rect 646966 161331 647018 161383
rect 676150 161331 676202 161383
rect 674134 161257 674186 161309
rect 676054 161257 676106 161309
rect 182902 161183 182954 161235
rect 184630 161183 184682 161235
rect 159862 161109 159914 161161
rect 184438 161109 184490 161161
rect 171382 161035 171434 161087
rect 184534 161035 184586 161087
rect 151318 160961 151370 161013
rect 184342 160961 184394 161013
rect 645142 159703 645194 159755
rect 650038 159703 650090 159755
rect 147094 158445 147146 158497
rect 151414 158445 151466 158497
rect 151798 158371 151850 158423
rect 184534 158371 184586 158423
rect 162646 158297 162698 158349
rect 184438 158297 184490 158349
rect 168406 158223 168458 158275
rect 184342 158223 184394 158275
rect 180022 158149 180074 158201
rect 184630 158149 184682 158201
rect 149398 157631 149450 157683
rect 159766 157631 159818 157683
rect 147094 156151 147146 156203
rect 151222 156151 151274 156203
rect 645142 156003 645194 156055
rect 650134 156003 650186 156055
rect 149398 155707 149450 155759
rect 182806 155707 182858 155759
rect 151990 155485 152042 155537
rect 184630 155485 184682 155537
rect 658006 155485 658058 155537
rect 675094 155485 675146 155537
rect 159958 155411 160010 155463
rect 184342 155411 184394 155463
rect 174358 155337 174410 155389
rect 184438 155337 184490 155389
rect 177238 155263 177290 155315
rect 184534 155263 184586 155315
rect 674134 153339 674186 153391
rect 675382 153339 675434 153391
rect 149494 152747 149546 152799
rect 172822 152747 172874 152799
rect 149398 152673 149450 152725
rect 179926 152673 179978 152725
rect 151894 152599 151946 152651
rect 184534 152599 184586 152651
rect 151606 152525 151658 152577
rect 184438 152525 184490 152577
rect 645142 152525 645194 152577
rect 650230 152525 650282 152577
rect 151702 152451 151754 152503
rect 184342 152451 184394 152503
rect 149398 149935 149450 149987
rect 174262 149935 174314 149987
rect 149494 149861 149546 149913
rect 177046 149861 177098 149913
rect 149686 149787 149738 149839
rect 180022 149787 180074 149839
rect 151510 149713 151562 149765
rect 184342 149713 184394 149765
rect 152086 149639 152138 149691
rect 184438 149639 184490 149691
rect 157078 149565 157130 149617
rect 184534 149565 184586 149617
rect 165718 149491 165770 149543
rect 184342 149491 184394 149543
rect 675190 149121 675242 149173
rect 675382 149121 675434 149173
rect 645142 148159 645194 148211
rect 650326 148159 650378 148211
rect 149014 147863 149066 147915
rect 149206 147863 149258 147915
rect 149206 147419 149258 147471
rect 149398 147419 149450 147471
rect 149398 146975 149450 147027
rect 168406 146975 168458 147027
rect 149494 146901 149546 146953
rect 171382 146901 171434 146953
rect 182998 146827 183050 146879
rect 186742 146827 186794 146879
rect 154198 146753 154250 146805
rect 184342 146753 184394 146805
rect 160054 146679 160106 146731
rect 184438 146679 184490 146731
rect 152182 146605 152234 146657
rect 184534 146605 184586 146657
rect 673462 146087 673514 146139
rect 675382 146087 675434 146139
rect 149398 144089 149450 144141
rect 162934 144089 162986 144141
rect 149494 144015 149546 144067
rect 165718 144015 165770 144067
rect 168598 143941 168650 143993
rect 184534 143941 184586 143993
rect 171574 143867 171626 143919
rect 184438 143867 184490 143919
rect 174454 143793 174506 143845
rect 184342 143793 184394 143845
rect 180214 143719 180266 143771
rect 185398 143719 185450 143771
rect 149494 142313 149546 142365
rect 159862 142313 159914 142365
rect 149398 141795 149450 141847
rect 156982 141795 157034 141847
rect 147094 141203 147146 141255
rect 154102 141203 154154 141255
rect 146902 141055 146954 141107
rect 151126 141055 151178 141107
rect 154294 141055 154346 141107
rect 184630 141055 184682 141107
rect 157174 140981 157226 141033
rect 184534 140981 184586 141033
rect 162838 140907 162890 140959
rect 184438 140907 184490 140959
rect 165814 140833 165866 140885
rect 184342 140833 184394 140885
rect 149398 138243 149450 138295
rect 162646 138243 162698 138295
rect 172822 136763 172874 136815
rect 185686 136763 185738 136815
rect 149398 135431 149450 135483
rect 174166 135431 174218 135483
rect 149686 135357 149738 135409
rect 182902 135357 182954 135409
rect 162742 135283 162794 135335
rect 184342 135283 184394 135335
rect 183094 134913 183146 134965
rect 184534 134913 184586 134965
rect 177334 134839 177386 134891
rect 184438 134839 184490 134891
rect 148822 133951 148874 134003
rect 149590 133951 149642 134003
rect 148918 132915 148970 132967
rect 149686 132915 149738 132967
rect 149398 132471 149450 132523
rect 171286 132471 171338 132523
rect 156886 132397 156938 132449
rect 184630 132397 184682 132449
rect 165526 132323 165578 132375
rect 184534 132323 184586 132375
rect 168502 132249 168554 132301
rect 184438 132249 184490 132301
rect 171478 132175 171530 132227
rect 184342 132175 184394 132227
rect 149398 129659 149450 129711
rect 165622 129659 165674 129711
rect 149302 129585 149354 129637
rect 177238 129585 177290 129637
rect 655318 129585 655370 129637
rect 676246 129585 676298 129637
rect 149206 129511 149258 129563
rect 184438 129511 184490 129563
rect 149494 129437 149546 129489
rect 184534 129437 184586 129489
rect 149110 129363 149162 129415
rect 184630 129363 184682 129415
rect 154006 129289 154058 129341
rect 184342 129289 184394 129341
rect 655222 127069 655274 127121
rect 676246 127069 676298 127121
rect 655126 126921 655178 126973
rect 676342 126921 676394 126973
rect 647926 126773 647978 126825
rect 676150 126773 676202 126825
rect 149398 126699 149450 126751
rect 156886 126699 156938 126751
rect 646582 126699 646634 126751
rect 676054 126699 676106 126751
rect 148534 126625 148586 126677
rect 184534 126625 184586 126677
rect 148726 126551 148778 126603
rect 184438 126551 184490 126603
rect 148918 126477 148970 126529
rect 184342 126477 184394 126529
rect 673846 126329 673898 126381
rect 676054 126329 676106 126381
rect 675190 123961 675242 124013
rect 676054 123961 676106 124013
rect 148438 123887 148490 123939
rect 154198 123887 154250 123939
rect 646486 123887 646538 123939
rect 676246 123887 676298 123939
rect 148246 123813 148298 123865
rect 184630 123813 184682 123865
rect 148534 123739 148586 123791
rect 184438 123739 184490 123791
rect 148630 123665 148682 123717
rect 184342 123665 184394 123717
rect 149686 123591 149738 123643
rect 184534 123591 184586 123643
rect 674614 121149 674666 121201
rect 675958 121149 676010 121201
rect 674710 121075 674762 121127
rect 676246 121075 676298 121127
rect 674998 121001 675050 121053
rect 676054 121001 676106 121053
rect 148342 120927 148394 120979
rect 184438 120927 184490 120979
rect 149494 120853 149546 120905
rect 184534 120853 184586 120905
rect 171382 120779 171434 120831
rect 184630 120779 184682 120831
rect 174262 120705 174314 120757
rect 184342 120705 184394 120757
rect 180022 120631 180074 120683
rect 186262 120631 186314 120683
rect 674326 119891 674378 119943
rect 676054 119891 676106 119943
rect 674806 118559 674858 118611
rect 676246 118559 676298 118611
rect 646198 118411 646250 118463
rect 676246 118411 676298 118463
rect 149398 118263 149450 118315
rect 168502 118263 168554 118315
rect 149494 118189 149546 118241
rect 174358 118189 174410 118241
rect 674422 118189 674474 118241
rect 675958 118189 676010 118241
rect 149398 118115 149450 118167
rect 180118 118115 180170 118167
rect 674902 118115 674954 118167
rect 676054 118115 676106 118167
rect 159862 118041 159914 118093
rect 184630 118041 184682 118093
rect 162934 117967 162986 118019
rect 184534 117967 184586 118019
rect 165718 117893 165770 117945
rect 184438 117893 184490 117945
rect 168406 117819 168458 117871
rect 184342 117819 184394 117871
rect 647734 115451 647786 115503
rect 676246 115451 676298 115503
rect 149398 115303 149450 115355
rect 162742 115303 162794 115355
rect 647830 115303 647882 115355
rect 676150 115303 676202 115355
rect 149494 115229 149546 115281
rect 165526 115229 165578 115281
rect 647926 115229 647978 115281
rect 665302 115229 665354 115281
rect 151414 115155 151466 115207
rect 184630 115155 184682 115207
rect 154102 115081 154154 115133
rect 184438 115081 184490 115133
rect 156982 115007 157034 115059
rect 184342 115007 184394 115059
rect 159766 114933 159818 114985
rect 184534 114933 184586 114985
rect 663766 114637 663818 114689
rect 675382 114637 675434 114689
rect 177238 113897 177290 113949
rect 184726 113897 184778 113949
rect 149494 112713 149546 112765
rect 159862 112713 159914 112765
rect 149398 112343 149450 112395
rect 177142 112343 177194 112395
rect 151222 112269 151274 112321
rect 184342 112269 184394 112321
rect 182806 112195 182858 112247
rect 184534 112195 184586 112247
rect 674614 110271 674666 110323
rect 675382 110271 675434 110323
rect 674710 109679 674762 109731
rect 675478 109679 675530 109731
rect 149398 109531 149450 109583
rect 156982 109531 157034 109583
rect 162646 109383 162698 109435
rect 184342 109383 184394 109435
rect 179926 109309 179978 109361
rect 185302 109309 185354 109361
rect 177046 109235 177098 109287
rect 184438 109235 184490 109287
rect 674902 109013 674954 109065
rect 675382 109013 675434 109065
rect 147862 108347 147914 108399
rect 154006 108347 154058 108399
rect 154198 107977 154250 108029
rect 184630 107977 184682 108029
rect 147190 107163 147242 107215
rect 151126 107163 151178 107215
rect 182902 106497 182954 106549
rect 186646 106497 186698 106549
rect 171286 106423 171338 106475
rect 184534 106423 184586 106475
rect 174166 106349 174218 106401
rect 184342 106349 184394 106401
rect 149590 106275 149642 106327
rect 184438 106275 184490 106327
rect 674902 105905 674954 105957
rect 675478 105905 675530 105957
rect 674326 105239 674378 105291
rect 675382 105239 675434 105291
rect 674422 104721 674474 104773
rect 675382 104721 675434 104773
rect 654070 104499 654122 104551
rect 665590 104499 665642 104551
rect 645910 103833 645962 103885
rect 657526 103833 657578 103885
rect 647926 103759 647978 103811
rect 661174 103759 661226 103811
rect 149110 103611 149162 103663
rect 184534 103611 184586 103663
rect 149014 103537 149066 103589
rect 184342 103537 184394 103589
rect 165622 103463 165674 103515
rect 184438 103463 184490 103515
rect 645142 102057 645194 102109
rect 652438 102057 652490 102109
rect 149398 100799 149450 100851
rect 168406 100799 168458 100851
rect 149686 100725 149738 100777
rect 184534 100725 184586 100777
rect 149302 100651 149354 100703
rect 184438 100651 184490 100703
rect 156886 100577 156938 100629
rect 184342 100577 184394 100629
rect 149398 97987 149450 98039
rect 184246 97987 184298 98039
rect 149494 97913 149546 97965
rect 186166 97913 186218 97965
rect 647926 97913 647978 97965
rect 662518 97913 662570 97965
rect 148534 97839 148586 97891
rect 184342 97839 184394 97891
rect 148630 97765 148682 97817
rect 184438 97765 184490 97817
rect 168502 97691 168554 97743
rect 184534 97691 184586 97743
rect 640726 96507 640778 96559
rect 654070 96507 654122 96559
rect 645430 95915 645482 95967
rect 653686 95915 653738 95967
rect 149494 95101 149546 95153
rect 166678 95101 166730 95153
rect 149398 95027 149450 95079
rect 179926 95027 179978 95079
rect 162742 94953 162794 95005
rect 184534 94953 184586 95005
rect 165526 94879 165578 94931
rect 184438 94879 184490 94931
rect 174358 94805 174410 94857
rect 184342 94805 184394 94857
rect 180118 94583 180170 94635
rect 184630 94583 184682 94635
rect 646774 92659 646826 92711
rect 663094 92659 663146 92711
rect 149398 92363 149450 92415
rect 159574 92363 159626 92415
rect 646486 92363 646538 92415
rect 660694 92363 660746 92415
rect 645526 92289 645578 92341
rect 661750 92289 661802 92341
rect 646870 92215 646922 92267
rect 659830 92215 659882 92267
rect 149494 92141 149546 92193
rect 162358 92141 162410 92193
rect 647062 92141 647114 92193
rect 658870 92141 658922 92193
rect 148342 92067 148394 92119
rect 184534 92067 184586 92119
rect 148726 91993 148778 92045
rect 184438 91993 184490 92045
rect 159862 91919 159914 91971
rect 184342 91919 184394 91971
rect 177142 91845 177194 91897
rect 184630 91845 184682 91897
rect 148822 89181 148874 89233
rect 184630 89181 184682 89233
rect 151126 89107 151178 89159
rect 184534 89107 184586 89159
rect 154006 89033 154058 89085
rect 184438 89033 184490 89085
rect 156982 88959 157034 89011
rect 184342 88959 184394 89011
rect 645910 87479 645962 87531
rect 650902 87479 650954 87531
rect 647926 87257 647978 87309
rect 658006 87257 658058 87309
rect 647158 87035 647210 87087
rect 663286 87035 663338 87087
rect 149494 86739 149546 86791
rect 156406 86739 156458 86791
rect 148726 86443 148778 86495
rect 154102 86443 154154 86495
rect 148438 86369 148490 86421
rect 184534 86369 184586 86421
rect 148246 86295 148298 86347
rect 184342 86295 184394 86347
rect 148918 86221 148970 86273
rect 184438 86221 184490 86273
rect 645910 84001 645962 84053
rect 657046 84001 657098 84053
rect 146998 83557 147050 83609
rect 151126 83557 151178 83609
rect 646774 83557 646826 83609
rect 651766 83557 651818 83609
rect 166678 83483 166730 83535
rect 184438 83483 184490 83535
rect 168406 83409 168458 83461
rect 184342 83409 184394 83461
rect 647926 81855 647978 81907
rect 663286 81855 663338 81907
rect 657046 81633 657098 81685
rect 658582 81633 658634 81685
rect 647830 81559 647882 81611
rect 662422 81559 662474 81611
rect 647734 81485 647786 81537
rect 663478 81485 663530 81537
rect 647926 80745 647978 80797
rect 662518 80745 662570 80797
rect 659446 80671 659498 80723
rect 659542 80671 659594 80723
rect 149590 80597 149642 80649
rect 184438 80597 184490 80649
rect 159574 80523 159626 80575
rect 184534 80523 184586 80575
rect 162358 80449 162410 80501
rect 184342 80449 184394 80501
rect 179926 80375 179978 80427
rect 184630 80375 184682 80427
rect 149302 77711 149354 77763
rect 184438 77711 184490 77763
rect 646966 77711 647018 77763
rect 658294 77711 658346 77763
rect 149398 77637 149450 77689
rect 184630 77637 184682 77689
rect 646582 77637 646634 77689
rect 659446 77637 659498 77689
rect 149206 77563 149258 77615
rect 184342 77563 184394 77615
rect 646678 77563 646730 77615
rect 661750 77563 661802 77615
rect 156406 77489 156458 77541
rect 184534 77489 184586 77541
rect 647926 77489 647978 77541
rect 656950 77489 657002 77541
rect 646006 76083 646058 76135
rect 657526 76083 657578 76135
rect 647158 74899 647210 74951
rect 660118 74899 660170 74951
rect 148630 74825 148682 74877
rect 184534 74825 184586 74877
rect 148918 74751 148970 74803
rect 184630 74751 184682 74803
rect 151126 74677 151178 74729
rect 184438 74677 184490 74729
rect 154102 74603 154154 74655
rect 184342 74603 184394 74655
rect 647926 72087 647978 72139
rect 660694 72087 660746 72139
rect 148246 71939 148298 71991
rect 184342 71939 184394 71991
rect 149590 71865 149642 71917
rect 184438 71865 184490 71917
rect 149686 71791 149738 71843
rect 184534 71791 184586 71843
rect 647926 69571 647978 69623
rect 661462 69571 661514 69623
rect 148822 69053 148874 69105
rect 184342 69053 184394 69105
rect 149590 68979 149642 69031
rect 184438 68979 184490 69031
rect 149302 68905 149354 68957
rect 184534 68905 184586 68957
rect 149206 68831 149258 68883
rect 184342 68831 184394 68883
rect 149110 66167 149162 66219
rect 184534 66167 184586 66219
rect 646006 66167 646058 66219
rect 652342 66167 652394 66219
rect 149494 66093 149546 66145
rect 184630 66093 184682 66145
rect 149398 66019 149450 66071
rect 184438 66019 184490 66071
rect 149014 65945 149066 65997
rect 184342 65945 184394 65997
rect 647926 63429 647978 63481
rect 663190 63429 663242 63481
rect 149590 63281 149642 63333
rect 184438 63281 184490 63333
rect 149494 63207 149546 63259
rect 184534 63207 184586 63259
rect 149398 63133 149450 63185
rect 184630 63133 184682 63185
rect 149206 63059 149258 63111
rect 184342 63059 184394 63111
rect 647926 60987 647978 61039
rect 663382 60987 663434 61039
rect 149398 60395 149450 60447
rect 184534 60395 184586 60447
rect 149302 60321 149354 60373
rect 184342 60321 184394 60373
rect 149494 60247 149546 60299
rect 184438 60247 184490 60299
rect 646006 59063 646058 59115
rect 652246 59063 652298 59115
rect 149398 58989 149450 59041
rect 184342 58989 184394 59041
rect 149398 57509 149450 57561
rect 184342 57509 184394 57561
rect 149398 56177 149450 56229
rect 184438 56177 184490 56229
rect 149494 56103 149546 56155
rect 184342 56103 184394 56155
rect 149686 54623 149738 54675
rect 184342 54623 184394 54675
rect 149398 53217 149450 53269
rect 184342 53217 184394 53269
rect 418774 48407 418826 48459
rect 424054 48407 424106 48459
rect 480982 48111 481034 48163
rect 527926 48111 527978 48163
rect 460342 48037 460394 48089
rect 510358 48037 510410 48089
rect 305302 47963 305354 48015
rect 354838 47963 354890 48015
rect 426166 47963 426218 48015
rect 492982 47963 493034 48015
rect 311062 47889 311114 47941
rect 371926 47889 371978 47941
rect 405526 47889 405578 47941
rect 441334 47889 441386 47941
rect 472246 47889 472298 47941
rect 562486 47889 562538 47941
rect 302902 47815 302954 47867
rect 506806 47815 506858 47867
rect 320182 47741 320234 47793
rect 529270 47741 529322 47793
rect 233686 47667 233738 47719
rect 475510 47667 475562 47719
rect 268534 47593 268586 47645
rect 520630 47593 520682 47645
rect 250966 47519 251018 47571
rect 521206 47519 521258 47571
rect 145366 47075 145418 47127
rect 199126 47075 199178 47127
rect 328342 46705 328394 46757
rect 337462 46705 337514 46757
rect 464854 46409 464906 46461
rect 475702 46409 475754 46461
rect 207382 46187 207434 46239
rect 216406 46187 216458 46239
rect 539734 46187 539786 46239
rect 545206 46187 545258 46239
rect 401782 46113 401834 46165
rect 406774 46113 406826 46165
rect 506806 44855 506858 44907
rect 512182 44855 512234 44907
rect 630742 43671 630794 43723
rect 640726 43671 640778 43723
rect 285814 43227 285866 43279
rect 518710 43227 518762 43279
rect 302902 43153 302954 43205
rect 305302 43153 305354 43205
rect 403222 43153 403274 43205
rect 418774 43153 418826 43205
rect 444886 43153 444938 43205
rect 458614 43153 458666 43205
rect 357718 42117 357770 42169
rect 307222 42043 307274 42095
rect 311062 42043 311114 42095
rect 362038 42043 362090 42095
rect 365974 42043 366026 42095
rect 401782 42043 401834 42095
rect 471670 42043 471722 42095
rect 480982 42043 481034 42095
rect 186262 41969 186314 42021
rect 187030 41969 187082 42021
rect 194326 41969 194378 42021
rect 630742 41969 630794 42021
rect 514006 41747 514058 41799
rect 514870 41747 514922 41799
rect 186262 41451 186314 41503
rect 207382 41451 207434 41503
rect 365878 37381 365930 37433
rect 403222 37455 403274 37507
rect 475510 37381 475562 37433
rect 514006 37381 514058 37433
rect 365974 37307 366026 37359
rect 389206 37307 389258 37359
rect 420790 34495 420842 34547
rect 444886 34495 444938 34547
<< metal2 >>
rect 175604 997770 175660 997779
rect 486740 997770 486796 997779
rect 175604 997705 175660 997714
rect 80564 997178 80620 997187
rect 80564 997113 80620 997122
rect 129524 997178 129580 997187
rect 129524 997113 129580 997122
rect 80578 982979 80606 997113
rect 129538 985009 129566 997113
rect 175618 992853 175646 997705
rect 175606 992847 175658 992853
rect 175606 992789 175658 992795
rect 178486 992847 178538 992853
rect 178486 992789 178538 992795
rect 178498 987840 178526 992789
rect 178498 987812 178622 987840
rect 129526 985003 129578 985009
rect 129526 984945 129578 984951
rect 132406 985003 132458 985009
rect 132406 984945 132458 984951
rect 132418 982979 132446 984945
rect 178594 983011 178622 987812
rect 178582 983005 178634 983011
rect 80564 982970 80620 982979
rect 80564 982905 80620 982914
rect 132404 982970 132460 982979
rect 184246 983005 184298 983011
rect 178582 982947 178634 982953
rect 184244 982970 184246 982979
rect 233218 982979 233246 997742
rect 238964 997178 239020 997187
rect 238964 997113 239020 997122
rect 238978 983127 239006 997113
rect 238964 983118 239020 983127
rect 238964 983053 239020 983062
rect 239938 982979 239966 997742
rect 285058 982979 285086 997742
rect 291298 993667 291326 997742
rect 486740 997705 486796 997714
rect 538580 997770 538636 997779
rect 538580 997705 538636 997714
rect 639380 997770 639436 997779
rect 639380 997705 639436 997714
rect 293108 997178 293164 997187
rect 293108 997113 293164 997122
rect 432020 997178 432076 997187
rect 432020 997113 432076 997122
rect 287926 993661 287978 993667
rect 287926 993603 287978 993609
rect 291286 993661 291338 993667
rect 291286 993603 291338 993609
rect 287938 983127 287966 993603
rect 287924 983118 287980 983127
rect 287924 983053 287980 983062
rect 293122 982979 293150 997113
rect 432034 983529 432062 997113
rect 399574 983523 399626 983529
rect 399574 983465 399626 983471
rect 432022 983523 432074 983529
rect 432022 983465 432074 983471
rect 399586 982979 399614 983465
rect 486754 982979 486782 997705
rect 538594 982979 538622 997705
rect 639394 982979 639422 997705
rect 184298 982970 184300 982979
rect 132404 982905 132460 982914
rect 184244 982905 184300 982914
rect 233204 982970 233260 982979
rect 233204 982905 233260 982914
rect 239924 982970 239980 982979
rect 239924 982905 239980 982914
rect 285044 982970 285100 982979
rect 285044 982905 285100 982914
rect 293108 982970 293164 982979
rect 293108 982905 293164 982914
rect 392468 982970 392524 982979
rect 392468 982905 392470 982914
rect 392522 982905 392524 982914
rect 394580 982970 394636 982979
rect 394580 982905 394636 982914
rect 399572 982970 399628 982979
rect 399572 982905 399628 982914
rect 486740 982970 486796 982979
rect 486740 982905 486796 982914
rect 538580 982970 538636 982979
rect 538580 982905 538636 982914
rect 639380 982970 639436 982979
rect 639380 982905 639436 982914
rect 649462 982931 649514 982937
rect 392470 982873 392522 982879
rect 394594 982863 394622 982905
rect 649462 982873 649514 982879
rect 394582 982857 394634 982863
rect 394582 982799 394634 982805
rect 649474 981975 649502 982873
rect 652246 982043 652298 982049
rect 652246 981985 652298 981991
rect 649462 981969 649514 981975
rect 649462 981911 649514 981917
rect 652258 979237 652286 981985
rect 656662 981969 656714 981975
rect 656662 981911 656714 981917
rect 652246 979231 652298 979237
rect 652246 979173 652298 979179
rect 656674 974945 656702 981911
rect 679702 979231 679754 979237
rect 679702 979173 679754 979179
rect 656662 974939 656714 974945
rect 656662 974881 656714 974887
rect 671062 974939 671114 974945
rect 671062 974881 671114 974887
rect 671074 963993 671102 974881
rect 671062 963987 671114 963993
rect 671062 963929 671114 963935
rect 677590 963987 677642 963993
rect 677590 963929 677642 963935
rect 40148 961954 40204 961963
rect 40148 961889 40150 961898
rect 40202 961889 40204 961898
rect 60022 961915 60074 961921
rect 40150 961857 40202 961863
rect 60022 961857 60074 961863
rect 60034 961815 60062 961857
rect 60020 961806 60076 961815
rect 60020 961741 60076 961750
rect 653780 959142 653836 959151
rect 653780 959077 653836 959086
rect 677494 959103 677546 959109
rect 653794 944383 653822 959077
rect 677494 959045 677546 959051
rect 677506 948916 677534 959045
rect 677602 958818 677630 963929
rect 679714 959109 679742 979173
rect 679702 959103 679754 959109
rect 679702 959045 679754 959051
rect 677506 948888 677616 948916
rect 653782 944377 653834 944383
rect 676822 944377 676874 944383
rect 653782 944319 653834 944325
rect 676820 944342 676822 944351
rect 676874 944342 676876 944351
rect 676820 944277 676876 944286
rect 676340 880258 676396 880267
rect 676340 880193 676396 880202
rect 676148 879666 676204 879675
rect 676148 879601 676204 879610
rect 654262 878665 654314 878671
rect 654262 878607 654314 878613
rect 654166 878591 654218 878597
rect 654166 878533 654218 878539
rect 654070 878517 654122 878523
rect 654070 878459 654122 878465
rect 654082 867687 654110 878459
rect 654178 868871 654206 878533
rect 654164 868862 654220 868871
rect 654164 868797 654220 868806
rect 654068 867678 654124 867687
rect 654068 867613 654124 867622
rect 649462 866973 649514 866979
rect 649462 866915 649514 866921
rect 649474 861134 649502 866915
rect 654274 866503 654302 878607
rect 676162 878597 676190 879601
rect 676244 879222 676300 879231
rect 676244 879157 676300 879166
rect 676258 878671 676286 879157
rect 676246 878665 676298 878671
rect 676246 878607 676298 878613
rect 676150 878591 676202 878597
rect 676150 878533 676202 878539
rect 676354 878523 676382 880193
rect 676342 878517 676394 878523
rect 676052 878482 676108 878491
rect 673366 878443 673418 878449
rect 676342 878459 676394 878465
rect 676052 878417 676054 878426
rect 673366 878385 673418 878391
rect 676106 878417 676108 878426
rect 676054 878385 676106 878391
rect 670870 877259 670922 877265
rect 670870 877201 670922 877207
rect 654260 866494 654316 866503
rect 654260 866429 654316 866438
rect 654260 864126 654316 864135
rect 654260 864061 654262 864070
rect 654314 864061 654316 864070
rect 654262 864029 654314 864035
rect 654836 862942 654892 862951
rect 654836 862877 654892 862886
rect 654850 861207 654878 862877
rect 656372 861906 656428 861915
rect 656372 861841 656428 861850
rect 656386 861281 656414 861841
rect 656374 861275 656426 861281
rect 656374 861217 656426 861223
rect 654838 861201 654890 861207
rect 654838 861143 654890 861149
rect 649378 861106 649502 861134
rect 41782 817985 41834 817991
rect 41780 817950 41782 817959
rect 47542 817985 47594 817991
rect 41834 817950 41836 817959
rect 47542 817927 47594 817933
rect 41780 817885 41836 817894
rect 41780 817358 41836 817367
rect 41780 817293 41782 817302
rect 41834 817293 41836 817302
rect 44758 817319 44810 817325
rect 41782 817261 41834 817267
rect 44758 817261 44810 817267
rect 41588 816618 41644 816627
rect 41588 816553 41590 816562
rect 41642 816553 41644 816562
rect 41590 816521 41642 816527
rect 41780 815878 41836 815887
rect 41780 815813 41782 815822
rect 41834 815813 41836 815822
rect 43222 815839 43274 815845
rect 41782 815781 41834 815787
rect 43222 815781 43274 815787
rect 41780 814916 41836 814925
rect 41780 814851 41782 814860
rect 41834 814851 41836 814860
rect 41782 814819 41834 814825
rect 41588 813658 41644 813667
rect 41588 813593 41590 813602
rect 41642 813593 41644 813602
rect 41590 813561 41642 813567
rect 42068 812918 42124 812927
rect 42068 812853 42124 812862
rect 34484 812474 34540 812483
rect 34484 812409 34540 812418
rect 34388 810254 34444 810263
rect 34388 810189 34444 810198
rect 28820 805666 28876 805675
rect 28820 805601 28876 805610
rect 28834 805231 28862 805601
rect 28820 805222 28876 805231
rect 28820 805157 28876 805166
rect 34402 804967 34430 810189
rect 34498 805083 34526 812409
rect 37364 811734 37420 811743
rect 37364 811669 37420 811678
rect 37378 806373 37406 811669
rect 41972 811364 42028 811373
rect 41972 811299 42028 811308
rect 41780 810846 41836 810855
rect 41780 810781 41836 810790
rect 40148 809662 40204 809671
rect 40148 809597 40204 809606
rect 37366 806367 37418 806373
rect 37366 806309 37418 806315
rect 34484 805074 34540 805083
rect 34484 805009 34540 805018
rect 34390 804961 34442 804967
rect 34390 804903 34442 804909
rect 40162 801415 40190 809597
rect 40244 809514 40300 809523
rect 40244 809449 40300 809458
rect 40150 801409 40202 801415
rect 40150 801351 40202 801357
rect 40258 801341 40286 809449
rect 41588 808182 41644 808191
rect 41588 808117 41644 808126
rect 41396 807146 41452 807155
rect 41396 807081 41452 807090
rect 41410 807039 41438 807081
rect 41398 807033 41450 807039
rect 41398 806975 41450 806981
rect 41602 806817 41630 808117
rect 41590 806811 41642 806817
rect 41590 806753 41642 806759
rect 41588 806702 41644 806711
rect 41588 806637 41644 806646
rect 41602 806521 41630 806637
rect 41590 806515 41642 806521
rect 41590 806457 41642 806463
rect 41588 806110 41644 806119
rect 41588 806045 41644 806054
rect 41602 805231 41630 806045
rect 41588 805222 41644 805231
rect 41588 805157 41590 805166
rect 41642 805157 41644 805166
rect 41590 805125 41642 805131
rect 40246 801335 40298 801341
rect 40246 801277 40298 801283
rect 41794 801045 41822 810781
rect 41876 808922 41932 808931
rect 41876 808857 41932 808866
rect 41890 808815 41918 808857
rect 41878 808809 41930 808815
rect 41878 808751 41930 808757
rect 41876 807886 41932 807895
rect 41876 807821 41932 807830
rect 41890 807113 41918 807821
rect 41878 807107 41930 807113
rect 41878 807049 41930 807055
rect 41878 804961 41930 804967
rect 41878 804903 41930 804909
rect 41890 801087 41918 804903
rect 41986 801119 42014 811299
rect 41974 801113 42026 801119
rect 41876 801078 41932 801087
rect 41782 801039 41834 801045
rect 41974 801055 42026 801061
rect 42082 801045 42110 812853
rect 42742 808809 42794 808815
rect 42742 808751 42794 808757
rect 42646 806367 42698 806373
rect 42646 806309 42698 806315
rect 41876 801013 41932 801022
rect 42070 801039 42122 801045
rect 41782 800981 41834 800987
rect 42070 800981 42122 800987
rect 41782 800817 41834 800823
rect 42658 800791 42686 806309
rect 41782 800759 41834 800765
rect 42644 800782 42700 800791
rect 41794 800236 41822 800759
rect 42644 800717 42700 800726
rect 42646 800669 42698 800675
rect 42646 800611 42698 800617
rect 42658 798973 42686 800611
rect 42166 798967 42218 798973
rect 42166 798909 42218 798915
rect 42646 798967 42698 798973
rect 42646 798909 42698 798915
rect 42178 798386 42206 798909
rect 42644 798858 42700 798867
rect 42644 798793 42700 798802
rect 42166 797931 42218 797937
rect 42166 797873 42218 797879
rect 42178 797761 42206 797873
rect 42166 797117 42218 797123
rect 42166 797059 42218 797065
rect 42178 796565 42206 797059
rect 42070 796303 42122 796309
rect 42070 796245 42122 796251
rect 42082 795944 42110 796245
rect 42166 795711 42218 795717
rect 42166 795653 42218 795659
rect 42178 795352 42206 795653
rect 42658 795569 42686 798793
rect 42754 797123 42782 808751
rect 43030 807107 43082 807113
rect 43030 807049 43082 807055
rect 42838 806811 42890 806817
rect 42838 806753 42890 806759
rect 42742 797117 42794 797123
rect 42742 797059 42794 797065
rect 42742 796969 42794 796975
rect 42742 796911 42794 796917
rect 42646 795563 42698 795569
rect 42646 795505 42698 795511
rect 42166 795267 42218 795273
rect 42166 795209 42218 795215
rect 42178 794725 42206 795209
rect 42646 794971 42698 794977
rect 42646 794913 42698 794919
rect 42070 794527 42122 794533
rect 42070 794469 42122 794475
rect 42082 794094 42110 794469
rect 42166 793787 42218 793793
rect 42166 793729 42218 793735
rect 42178 793502 42206 793729
rect 42658 792165 42686 794913
rect 42754 793793 42782 796911
rect 42850 795273 42878 806753
rect 42934 806515 42986 806521
rect 42934 806457 42986 806463
rect 42946 795717 42974 806457
rect 43042 800823 43070 807049
rect 43126 807033 43178 807039
rect 43126 806975 43178 806981
rect 43030 800817 43082 800823
rect 43030 800759 43082 800765
rect 43030 800669 43082 800675
rect 43030 800611 43082 800617
rect 43042 796309 43070 800611
rect 43138 800601 43166 806975
rect 43126 800595 43178 800601
rect 43126 800537 43178 800543
rect 43124 800486 43180 800495
rect 43124 800421 43180 800430
rect 43030 796303 43082 796309
rect 43030 796245 43082 796251
rect 43030 796155 43082 796161
rect 43030 796097 43082 796103
rect 42934 795711 42986 795717
rect 42934 795653 42986 795659
rect 42934 795563 42986 795569
rect 42934 795505 42986 795511
rect 42838 795267 42890 795273
rect 42838 795209 42890 795215
rect 42838 795119 42890 795125
rect 42838 795061 42890 795067
rect 42742 793787 42794 793793
rect 42742 793729 42794 793735
rect 42850 792165 42878 795061
rect 42646 792159 42698 792165
rect 42646 792101 42698 792107
rect 42838 792159 42890 792165
rect 42838 792101 42890 792107
rect 42550 791937 42602 791943
rect 42550 791879 42602 791885
rect 42562 791499 42590 791879
rect 42646 791863 42698 791869
rect 42646 791805 42698 791811
rect 42070 791493 42122 791499
rect 42070 791435 42122 791441
rect 42550 791493 42602 791499
rect 42550 791435 42602 791441
rect 42082 791060 42110 791435
rect 42658 790833 42686 791805
rect 42166 790827 42218 790833
rect 42166 790769 42218 790775
rect 42646 790827 42698 790833
rect 42646 790769 42698 790775
rect 42178 790394 42206 790769
rect 42164 790274 42220 790283
rect 42164 790209 42220 790218
rect 42178 789757 42206 790209
rect 42070 789643 42122 789649
rect 42070 789585 42122 789591
rect 42082 789210 42110 789585
rect 42646 789199 42698 789205
rect 42646 789141 42698 789147
rect 42262 787867 42314 787873
rect 42262 787809 42314 787815
rect 42274 787374 42302 787809
rect 42192 787346 42302 787374
rect 42166 787275 42218 787281
rect 42166 787217 42218 787223
rect 42178 786694 42206 787217
rect 41780 786426 41836 786435
rect 41780 786361 41836 786370
rect 41794 786102 41822 786361
rect 42658 785949 42686 789141
rect 42946 787281 42974 795505
rect 43042 794533 43070 796097
rect 43030 794527 43082 794533
rect 43030 794469 43082 794475
rect 43028 793974 43084 793983
rect 43028 793909 43084 793918
rect 43042 787873 43070 793909
rect 43138 789649 43166 800421
rect 43126 789643 43178 789649
rect 43126 789585 43178 789591
rect 43030 787867 43082 787873
rect 43030 787809 43082 787815
rect 42934 787275 42986 787281
rect 42934 787217 42986 787223
rect 42166 785943 42218 785949
rect 42166 785885 42218 785891
rect 42646 785943 42698 785949
rect 42646 785885 42698 785891
rect 42178 785510 42206 785885
rect 41780 774734 41836 774743
rect 41780 774669 41782 774678
rect 41834 774669 41836 774678
rect 41782 774637 41834 774643
rect 41588 773994 41644 774003
rect 41588 773929 41590 773938
rect 41642 773929 41644 773938
rect 41590 773897 41642 773903
rect 41780 773550 41836 773559
rect 41780 773485 41782 773494
rect 41834 773485 41836 773494
rect 41782 773453 41834 773459
rect 43234 773443 43262 815781
rect 44662 814877 44714 814883
rect 44662 814819 44714 814825
rect 44566 813619 44618 813625
rect 44566 813561 44618 813567
rect 43414 801409 43466 801415
rect 43414 801351 43466 801357
rect 43318 801335 43370 801341
rect 43318 801277 43370 801283
rect 43330 799269 43358 801277
rect 43426 800643 43454 801351
rect 43510 801113 43562 801119
rect 43510 801055 43562 801061
rect 43412 800634 43468 800643
rect 43412 800569 43468 800578
rect 43414 800521 43466 800527
rect 43414 800463 43466 800469
rect 43318 799263 43370 799269
rect 43318 799205 43370 799211
rect 43318 797931 43370 797937
rect 43318 797873 43370 797879
rect 43330 789797 43358 797873
rect 43426 796161 43454 800463
rect 43522 796975 43550 801055
rect 43606 800817 43658 800823
rect 43606 800759 43658 800765
rect 43618 800654 43646 800759
rect 43618 800626 43742 800654
rect 43606 799263 43658 799269
rect 43606 799205 43658 799211
rect 43510 796969 43562 796975
rect 43510 796911 43562 796917
rect 43414 796155 43466 796161
rect 43414 796097 43466 796103
rect 43618 795125 43646 799205
rect 43606 795119 43658 795125
rect 43606 795061 43658 795067
rect 43714 794977 43742 800626
rect 43702 794971 43754 794977
rect 43702 794913 43754 794919
rect 43318 789791 43370 789797
rect 43318 789733 43370 789739
rect 41590 773437 41642 773443
rect 41588 773402 41590 773411
rect 43222 773437 43274 773443
rect 41642 773402 41644 773411
rect 43222 773379 43274 773385
rect 41588 773337 41644 773346
rect 41780 772662 41836 772671
rect 41780 772597 41782 772606
rect 41834 772597 41836 772606
rect 43222 772623 43274 772629
rect 41782 772565 41834 772571
rect 43222 772565 43274 772571
rect 41588 772366 41644 772375
rect 41588 772301 41644 772310
rect 41602 772185 41630 772301
rect 41590 772179 41642 772185
rect 41590 772121 41642 772127
rect 41602 770895 41630 772121
rect 43126 771957 43178 771963
rect 43124 771922 43126 771931
rect 43178 771922 43180 771931
rect 43124 771857 43180 771866
rect 41588 770886 41644 770895
rect 41588 770821 41644 770830
rect 41780 769702 41836 769711
rect 41780 769637 41782 769646
rect 41834 769637 41836 769646
rect 43126 769663 43178 769669
rect 41782 769605 41834 769611
rect 43126 769605 43178 769611
rect 37364 768518 37420 768527
rect 37364 768453 37420 768462
rect 28820 762450 28876 762459
rect 28820 762385 28876 762394
rect 28834 762015 28862 762385
rect 28820 762006 28876 762015
rect 28820 761941 28876 761950
rect 37378 760271 37406 768453
rect 42260 768222 42316 768231
rect 42260 768157 42316 768166
rect 41876 767630 41932 767639
rect 41876 767565 41932 767574
rect 40244 766446 40300 766455
rect 40244 766381 40300 766390
rect 40148 766298 40204 766307
rect 40148 766233 40204 766242
rect 37366 760265 37418 760271
rect 37366 760207 37418 760213
rect 40162 758125 40190 766233
rect 40258 760345 40286 766381
rect 41588 765558 41644 765567
rect 41588 765493 41644 765502
rect 41602 763601 41630 765493
rect 41780 765188 41836 765197
rect 41780 765123 41782 765132
rect 41834 765123 41836 765132
rect 41782 765091 41834 765097
rect 41590 763595 41642 763601
rect 41590 763537 41642 763543
rect 41588 763486 41644 763495
rect 41588 763421 41590 763430
rect 41642 763421 41644 763430
rect 41590 763389 41642 763395
rect 41780 762154 41836 762163
rect 41780 762089 41782 762098
rect 41834 762089 41836 762098
rect 41782 762057 41834 762063
rect 40246 760339 40298 760345
rect 40246 760281 40298 760287
rect 41014 760339 41066 760345
rect 41014 760281 41066 760287
rect 41026 760239 41054 760281
rect 41782 760265 41834 760271
rect 41012 760230 41068 760239
rect 41782 760207 41834 760213
rect 41012 760165 41068 760174
rect 40150 758119 40202 758125
rect 40150 758061 40202 758067
rect 41794 758019 41822 760207
rect 41780 758010 41836 758019
rect 41780 757945 41836 757954
rect 41890 757829 41918 767565
rect 42068 767186 42124 767195
rect 42068 767121 42124 767130
rect 41972 764226 42028 764235
rect 41972 764161 42028 764170
rect 41986 757903 42014 764161
rect 41974 757897 42026 757903
rect 42082 757871 42110 767121
rect 42164 764670 42220 764679
rect 42164 764605 42220 764614
rect 41974 757839 42026 757845
rect 42068 757862 42124 757871
rect 41878 757823 41930 757829
rect 42178 757829 42206 764605
rect 42274 757977 42302 768157
rect 42742 765149 42794 765155
rect 42742 765091 42794 765097
rect 42262 757971 42314 757977
rect 42262 757913 42314 757919
rect 42068 757797 42124 757806
rect 42166 757823 42218 757829
rect 41878 757765 41930 757771
rect 42166 757765 42218 757771
rect 41878 757601 41930 757607
rect 41878 757543 41930 757549
rect 41890 757020 41918 757543
rect 42754 756423 42782 765091
rect 42934 763595 42986 763601
rect 42934 763537 42986 763543
rect 42838 763447 42890 763453
rect 42838 763389 42890 763395
rect 42742 756417 42794 756423
rect 42742 756359 42794 756365
rect 42358 756195 42410 756201
rect 42358 756137 42410 756143
rect 42166 755751 42218 755757
rect 42166 755693 42218 755699
rect 42178 755205 42206 755693
rect 42070 754715 42122 754721
rect 42070 754657 42122 754663
rect 42082 754578 42110 754657
rect 42166 753901 42218 753907
rect 42166 753843 42218 753849
rect 42178 753365 42206 753843
rect 42082 752427 42110 752728
rect 42166 752643 42218 752649
rect 42166 752585 42218 752591
rect 42070 752421 42122 752427
rect 42070 752363 42122 752369
rect 42178 752169 42206 752585
rect 42370 752057 42398 756137
rect 42850 752649 42878 763389
rect 42946 753907 42974 763537
rect 43138 755757 43166 769605
rect 43126 755751 43178 755757
rect 43126 755693 43178 755699
rect 43126 755603 43178 755609
rect 43126 755545 43178 755551
rect 42934 753901 42986 753907
rect 42934 753843 42986 753849
rect 42934 753753 42986 753759
rect 42934 753695 42986 753701
rect 42838 752643 42890 752649
rect 42838 752585 42890 752591
rect 42836 752534 42892 752543
rect 42836 752469 42892 752478
rect 42358 752051 42410 752057
rect 42358 751993 42410 751999
rect 42070 751903 42122 751909
rect 42070 751845 42122 751851
rect 42358 751903 42410 751909
rect 42358 751845 42410 751851
rect 42082 751544 42110 751845
rect 42370 751613 42398 751845
rect 42850 751687 42878 752469
rect 42838 751681 42890 751687
rect 42838 751623 42890 751629
rect 42358 751607 42410 751613
rect 42358 751549 42410 751555
rect 42838 751533 42890 751539
rect 42838 751475 42890 751481
rect 42166 751311 42218 751317
rect 42166 751253 42218 751259
rect 42178 750878 42206 751253
rect 42166 750571 42218 750577
rect 42166 750513 42218 750519
rect 42178 750329 42206 750513
rect 42850 748209 42878 751475
rect 42946 751317 42974 753695
rect 43138 751909 43166 755545
rect 43126 751903 43178 751909
rect 43126 751845 43178 751851
rect 43030 751829 43082 751835
rect 43030 751771 43082 751777
rect 42934 751311 42986 751317
rect 42934 751253 42986 751259
rect 42932 751202 42988 751211
rect 42932 751137 42988 751146
rect 42166 748203 42218 748209
rect 42166 748145 42218 748151
rect 42838 748203 42890 748209
rect 42838 748145 42890 748151
rect 42178 747844 42206 748145
rect 42166 747611 42218 747617
rect 42166 747553 42218 747559
rect 42178 747178 42206 747553
rect 42836 747354 42892 747363
rect 42836 747289 42892 747298
rect 41780 747058 41836 747067
rect 41780 746993 41836 747002
rect 41794 746557 41822 746993
rect 42166 746279 42218 746285
rect 42166 746221 42218 746227
rect 42178 745994 42206 746221
rect 42274 746137 42398 746156
rect 42274 746131 42410 746137
rect 42274 746128 42358 746131
rect 42358 746073 42410 746079
rect 42358 745983 42410 745989
rect 42358 745925 42410 745931
rect 42166 744651 42218 744657
rect 42166 744593 42218 744599
rect 42178 744144 42206 744593
rect 42166 744059 42218 744065
rect 42166 744001 42218 744007
rect 42178 743521 42206 744001
rect 42070 743393 42122 743399
rect 42070 743335 42122 743341
rect 42082 742886 42110 743335
rect 42370 742807 42398 745925
rect 42850 743399 42878 747289
rect 42946 746285 42974 751137
rect 43042 750577 43070 751771
rect 43126 751681 43178 751687
rect 43126 751623 43178 751629
rect 43030 750571 43082 750577
rect 43030 750513 43082 750519
rect 43028 748834 43084 748843
rect 43028 748769 43084 748778
rect 42934 746279 42986 746285
rect 42934 746221 42986 746227
rect 43042 744657 43070 748769
rect 43030 744651 43082 744657
rect 43030 744593 43082 744599
rect 43138 744065 43166 751623
rect 43126 744059 43178 744065
rect 43126 744001 43178 744007
rect 42838 743393 42890 743399
rect 42838 743335 42890 743341
rect 42166 742801 42218 742807
rect 42166 742743 42218 742749
rect 42358 742801 42410 742807
rect 42358 742743 42410 742749
rect 42178 742325 42206 742743
rect 41780 731518 41836 731527
rect 41780 731453 41782 731462
rect 41834 731453 41836 731462
rect 41782 731421 41834 731427
rect 41588 730778 41644 730787
rect 41588 730713 41590 730722
rect 41642 730713 41644 730722
rect 41590 730681 41642 730687
rect 41780 730408 41836 730417
rect 41780 730343 41782 730352
rect 41834 730343 41836 730352
rect 41782 730311 41834 730317
rect 43234 730227 43262 772565
rect 43606 758119 43658 758125
rect 43606 758061 43658 758067
rect 43510 757971 43562 757977
rect 43510 757913 43562 757919
rect 43414 757897 43466 757903
rect 43414 757839 43466 757845
rect 43318 757823 43370 757829
rect 43318 757765 43370 757771
rect 43330 755609 43358 757765
rect 43318 755603 43370 755609
rect 43318 755545 43370 755551
rect 43318 754715 43370 754721
rect 43318 754657 43370 754663
rect 43330 748801 43358 754657
rect 43426 753759 43454 757839
rect 43414 753753 43466 753759
rect 43414 753695 43466 753701
rect 43414 752421 43466 752427
rect 43414 752363 43466 752369
rect 43318 748795 43370 748801
rect 43318 748737 43370 748743
rect 43426 745323 43454 752363
rect 43522 751835 43550 757913
rect 43510 751829 43562 751835
rect 43510 751771 43562 751777
rect 43618 747617 43646 758061
rect 43606 747611 43658 747617
rect 43606 747553 43658 747559
rect 43414 745317 43466 745323
rect 43414 745259 43466 745265
rect 41590 730221 41642 730227
rect 41588 730186 41590 730195
rect 43222 730221 43274 730227
rect 41642 730186 41644 730195
rect 43222 730163 43274 730169
rect 41588 730121 41644 730130
rect 41204 729298 41260 729307
rect 41204 729233 41260 729242
rect 41588 729298 41644 729307
rect 41588 729233 41590 729242
rect 41218 728895 41246 729233
rect 41642 729233 41644 729242
rect 43702 729259 43754 729265
rect 41590 729201 41642 729207
rect 43702 729201 43754 729207
rect 41206 728889 41258 728895
rect 41206 728831 41258 728837
rect 40438 728815 40490 728821
rect 40438 728757 40490 728763
rect 40450 728715 40478 728757
rect 40436 728706 40492 728715
rect 40436 728641 40492 728650
rect 41588 728706 41644 728715
rect 41588 728641 41590 728650
rect 41642 728641 41644 728650
rect 43510 728667 43562 728673
rect 41590 728609 41642 728615
rect 43510 728609 43562 728615
rect 41780 727966 41836 727975
rect 41780 727901 41782 727910
rect 41834 727901 41836 727910
rect 43414 727927 43466 727933
rect 41782 727869 41834 727875
rect 43414 727869 43466 727875
rect 34484 726782 34540 726791
rect 34484 726717 34540 726726
rect 28820 719234 28876 719243
rect 28820 719169 28876 719178
rect 28834 718799 28862 719169
rect 28820 718790 28876 718799
rect 28820 718725 28876 718734
rect 34498 717763 34526 726717
rect 41780 726486 41836 726495
rect 41780 726421 41836 726430
rect 41794 726157 41822 726421
rect 41782 726151 41834 726157
rect 41782 726093 41834 726099
rect 42934 726151 42986 726157
rect 42934 726093 42986 726099
rect 37364 725302 37420 725311
rect 37364 725237 37420 725246
rect 37378 718651 37406 725237
rect 41972 725006 42028 725015
rect 41972 724941 42028 724950
rect 41780 724414 41836 724423
rect 41780 724349 41836 724358
rect 40148 723230 40204 723239
rect 40148 723165 40204 723174
rect 37364 718642 37420 718651
rect 37364 718577 37420 718586
rect 34484 717754 34540 717763
rect 34484 717689 34540 717698
rect 40162 716875 40190 723165
rect 40244 723082 40300 723091
rect 40244 723017 40300 723026
rect 40258 717023 40286 723017
rect 41588 722342 41644 722351
rect 41588 722277 41644 722286
rect 41602 721421 41630 722277
rect 41590 721415 41642 721421
rect 41590 721357 41642 721363
rect 41588 720862 41644 720871
rect 41588 720797 41644 720806
rect 41602 720459 41630 720797
rect 41590 720453 41642 720459
rect 41590 720395 41642 720401
rect 41588 720270 41644 720279
rect 41588 720205 41590 720214
rect 41642 720205 41644 720214
rect 41590 720173 41642 720179
rect 41588 718790 41644 718799
rect 41588 718725 41590 718734
rect 41642 718725 41644 718734
rect 41590 718693 41642 718699
rect 40244 717014 40300 717023
rect 40244 716949 40300 716958
rect 40148 716866 40204 716875
rect 40148 716801 40204 716810
rect 41794 714613 41822 724349
rect 41876 721972 41932 721981
rect 41876 721907 41932 721916
rect 41890 714613 41918 721907
rect 41986 714687 42014 724941
rect 42260 721454 42316 721463
rect 42260 721389 42316 721398
rect 41974 714681 42026 714687
rect 41974 714623 42026 714629
rect 41782 714607 41834 714613
rect 41782 714549 41834 714555
rect 41878 714607 41930 714613
rect 41878 714549 41930 714555
rect 41782 714385 41834 714391
rect 41782 714327 41834 714333
rect 41794 713845 41822 714327
rect 42274 714317 42302 721389
rect 42838 720453 42890 720459
rect 42838 720395 42890 720401
rect 42262 714311 42314 714317
rect 42262 714253 42314 714259
rect 42850 713004 42878 720395
rect 42754 712976 42878 713004
rect 42070 712535 42122 712541
rect 42070 712477 42122 712483
rect 42082 712028 42110 712477
rect 42178 711283 42206 711374
rect 42166 711277 42218 711283
rect 42166 711219 42218 711225
rect 42070 710685 42122 710691
rect 42070 710627 42122 710633
rect 42082 710178 42110 710627
rect 42166 709649 42218 709655
rect 42166 709591 42218 709597
rect 42178 709512 42206 709591
rect 42070 709427 42122 709433
rect 42070 709369 42122 709375
rect 42082 708994 42110 709369
rect 42166 708687 42218 708693
rect 42166 708629 42218 708635
rect 42178 708328 42206 708629
rect 42754 708249 42782 712976
rect 42838 712905 42890 712911
rect 42838 712847 42890 712853
rect 42850 710691 42878 712847
rect 42946 712541 42974 726093
rect 43126 721415 43178 721421
rect 43126 721357 43178 721363
rect 43030 720231 43082 720237
rect 43030 720173 43082 720179
rect 42934 712535 42986 712541
rect 42934 712477 42986 712483
rect 42934 712387 42986 712393
rect 42934 712329 42986 712335
rect 42838 710685 42890 710691
rect 42838 710627 42890 710633
rect 42838 710537 42890 710543
rect 42838 710479 42890 710485
rect 42850 708693 42878 710479
rect 42838 708687 42890 708693
rect 42838 708629 42890 708635
rect 42836 708578 42892 708587
rect 42836 708513 42892 708522
rect 42166 708243 42218 708249
rect 42166 708185 42218 708191
rect 42742 708243 42794 708249
rect 42742 708185 42794 708191
rect 42178 707662 42206 708185
rect 42742 708095 42794 708101
rect 42742 708037 42794 708043
rect 42070 707281 42122 707287
rect 42070 707223 42122 707229
rect 42082 707144 42110 707223
rect 42754 705585 42782 708037
rect 42358 705579 42410 705585
rect 42358 705521 42410 705527
rect 42742 705579 42794 705585
rect 42742 705521 42794 705527
rect 42370 705141 42398 705521
rect 42740 705470 42796 705479
rect 42740 705405 42796 705414
rect 42166 705135 42218 705141
rect 42166 705077 42218 705083
rect 42358 705135 42410 705141
rect 42358 705077 42410 705083
rect 42178 704628 42206 705077
rect 42166 704543 42218 704549
rect 42166 704485 42218 704491
rect 42178 704001 42206 704485
rect 42070 703803 42122 703809
rect 42070 703745 42122 703751
rect 42082 703370 42110 703745
rect 42166 703285 42218 703291
rect 42166 703227 42218 703233
rect 42178 702778 42206 703227
rect 41780 701326 41836 701335
rect 41780 701261 41836 701270
rect 41794 700965 41822 701261
rect 42070 700843 42122 700849
rect 42070 700785 42122 700791
rect 42082 700336 42110 700785
rect 42754 700257 42782 705405
rect 42850 704549 42878 708513
rect 42946 707287 42974 712329
rect 43042 709433 43070 720173
rect 43138 712911 43166 721357
rect 43318 714681 43370 714687
rect 43318 714623 43370 714629
rect 43222 714311 43274 714317
rect 43222 714253 43274 714259
rect 43126 712905 43178 712911
rect 43126 712847 43178 712853
rect 43234 712708 43262 714253
rect 43138 712680 43262 712708
rect 43030 709427 43082 709433
rect 43030 709369 43082 709375
rect 43138 709008 43166 712680
rect 43222 712609 43274 712615
rect 43222 712551 43274 712557
rect 43042 708980 43166 709008
rect 43042 708841 43070 708980
rect 43124 708874 43180 708883
rect 43030 708835 43082 708841
rect 43124 708809 43180 708818
rect 43030 708777 43082 708783
rect 43028 708726 43084 708735
rect 43028 708661 43084 708670
rect 42934 707281 42986 707287
rect 42934 707223 42986 707229
rect 42932 705914 42988 705923
rect 42932 705849 42988 705858
rect 42838 704543 42890 704549
rect 42838 704485 42890 704491
rect 42836 702066 42892 702075
rect 42836 702001 42892 702010
rect 42166 700251 42218 700257
rect 42166 700193 42218 700199
rect 42742 700251 42794 700257
rect 42742 700193 42794 700199
rect 42178 699670 42206 700193
rect 42850 699591 42878 702001
rect 42946 700849 42974 705849
rect 43042 703291 43070 708661
rect 43138 703809 43166 708809
rect 43126 703803 43178 703809
rect 43126 703745 43178 703751
rect 43030 703285 43082 703291
rect 43030 703227 43082 703233
rect 42934 700843 42986 700849
rect 42934 700785 42986 700791
rect 42070 699585 42122 699591
rect 42070 699527 42122 699533
rect 42838 699585 42890 699591
rect 42838 699527 42890 699533
rect 42082 699152 42110 699527
rect 41780 688302 41836 688311
rect 41780 688237 41782 688246
rect 41834 688237 41836 688246
rect 41782 688205 41834 688211
rect 41588 687562 41644 687571
rect 41588 687497 41590 687506
rect 41642 687497 41644 687506
rect 41590 687465 41642 687471
rect 41780 687266 41836 687275
rect 41780 687201 41782 687210
rect 41834 687201 41836 687210
rect 41782 687169 41834 687175
rect 41590 687005 41642 687011
rect 41588 686970 41590 686979
rect 41642 686970 41644 686979
rect 41588 686905 41644 686914
rect 41588 686082 41644 686091
rect 41588 686017 41590 686026
rect 41642 686017 41644 686026
rect 41590 685985 41642 685991
rect 43234 685383 43262 712551
rect 43330 712393 43358 714623
rect 43318 712387 43370 712393
rect 43318 712329 43370 712335
rect 43318 712239 43370 712245
rect 43318 712181 43370 712187
rect 43330 687011 43358 712181
rect 43318 687005 43370 687011
rect 43318 686947 43370 686953
rect 41782 685377 41834 685383
rect 41780 685342 41782 685351
rect 43222 685377 43274 685383
rect 41834 685342 41836 685351
rect 43222 685319 43274 685325
rect 41780 685277 41836 685286
rect 41588 684602 41644 684611
rect 41588 684537 41590 684546
rect 41642 684537 41644 684546
rect 43318 684563 43370 684569
rect 41590 684505 41642 684511
rect 43318 684505 43370 684511
rect 41782 684193 41834 684199
rect 41780 684158 41782 684167
rect 41834 684158 41836 684167
rect 41780 684093 41836 684102
rect 41780 683270 41836 683279
rect 41780 683205 41836 683214
rect 41794 682793 41822 683205
rect 41782 682787 41834 682793
rect 41782 682729 41834 682735
rect 43126 682787 43178 682793
rect 43126 682729 43178 682735
rect 42260 681198 42316 681207
rect 42260 681133 42316 681142
rect 41588 679126 41644 679135
rect 41588 679061 41644 679070
rect 41602 677317 41630 679061
rect 41590 677311 41642 677317
rect 41590 677253 41642 677259
rect 41780 677276 41836 677285
rect 41780 677211 41782 677220
rect 41834 677211 41836 677220
rect 41782 677179 41834 677185
rect 41780 676758 41836 676767
rect 41780 676693 41836 676702
rect 28820 676018 28876 676027
rect 28820 675953 28876 675962
rect 28834 675583 28862 675953
rect 41794 675805 41822 676693
rect 41780 675796 41836 675805
rect 41780 675731 41782 675740
rect 41834 675731 41836 675740
rect 41782 675699 41834 675705
rect 28820 675574 28876 675583
rect 28820 675509 28876 675518
rect 42274 670805 42302 681133
rect 42934 677311 42986 677317
rect 42934 677253 42986 677259
rect 42838 677237 42890 677243
rect 42838 677179 42890 677185
rect 42742 671095 42794 671101
rect 42742 671037 42794 671043
rect 42262 670799 42314 670805
rect 42262 670741 42314 670747
rect 42166 670577 42218 670583
rect 42166 670519 42218 670525
rect 42178 670440 42206 670519
rect 42166 669171 42218 669177
rect 42166 669113 42218 669119
rect 42178 668590 42206 669113
rect 42754 668511 42782 671037
rect 42850 668585 42878 677179
rect 42946 671054 42974 677253
rect 42946 671026 43070 671054
rect 42932 668618 42988 668627
rect 42838 668579 42890 668585
rect 42932 668553 42988 668562
rect 42838 668521 42890 668527
rect 42166 668505 42218 668511
rect 42166 668447 42218 668453
rect 42742 668505 42794 668511
rect 42742 668447 42794 668453
rect 42836 668470 42892 668479
rect 42178 667961 42206 668447
rect 42836 668405 42892 668414
rect 42740 668322 42796 668331
rect 42740 668257 42796 668266
rect 42166 667321 42218 667327
rect 42166 667263 42218 667269
rect 42178 666740 42206 667263
rect 42070 665915 42122 665921
rect 42070 665857 42122 665863
rect 42082 665556 42110 665857
rect 42178 665699 42206 666148
rect 42166 665693 42218 665699
rect 42166 665635 42218 665641
rect 42754 665477 42782 668257
rect 42166 665471 42218 665477
rect 42166 665413 42218 665419
rect 42742 665471 42794 665477
rect 42742 665413 42794 665419
rect 42178 664925 42206 665413
rect 42740 665362 42796 665371
rect 42740 665297 42796 665306
rect 42070 664657 42122 664663
rect 42070 664599 42122 664605
rect 42082 664298 42110 664599
rect 42166 664213 42218 664219
rect 42166 664155 42218 664161
rect 42178 663706 42206 664155
rect 42356 662402 42412 662411
rect 42356 662337 42412 662346
rect 42070 661697 42122 661703
rect 42070 661639 42122 661645
rect 42082 661264 42110 661639
rect 42166 661179 42218 661185
rect 42166 661121 42218 661127
rect 42178 660598 42206 661121
rect 42166 660291 42218 660297
rect 42166 660233 42218 660239
rect 42178 659932 42206 660233
rect 42370 659705 42398 662337
rect 42754 661185 42782 665297
rect 42850 664219 42878 668405
rect 42946 664663 42974 668553
rect 43042 667327 43070 671026
rect 43138 669177 43166 682729
rect 43330 679694 43358 684505
rect 43426 684199 43454 727869
rect 43522 712615 43550 728609
rect 43606 714607 43658 714613
rect 43606 714549 43658 714555
rect 43510 712609 43562 712615
rect 43510 712551 43562 712557
rect 43618 710543 43646 714549
rect 43714 712245 43742 729201
rect 43702 712239 43754 712245
rect 43702 712181 43754 712187
rect 43702 711277 43754 711283
rect 43702 711219 43754 711225
rect 43606 710537 43658 710543
rect 43606 710479 43658 710485
rect 43510 709649 43562 709655
rect 43510 709591 43562 709597
rect 43522 702699 43550 709591
rect 43714 704919 43742 711219
rect 43702 704913 43754 704919
rect 43702 704855 43754 704861
rect 43510 702693 43562 702699
rect 43510 702635 43562 702641
rect 43510 686043 43562 686049
rect 43510 685985 43562 685991
rect 43414 684193 43466 684199
rect 43414 684135 43466 684141
rect 43330 679666 43454 679694
rect 43126 669171 43178 669177
rect 43126 669113 43178 669119
rect 43126 668579 43178 668585
rect 43126 668521 43178 668527
rect 43030 667321 43082 667327
rect 43030 667263 43082 667269
rect 43028 666250 43084 666259
rect 43028 666185 43084 666194
rect 42934 664657 42986 664663
rect 42934 664599 42986 664605
rect 42932 664326 42988 664335
rect 42932 664261 42988 664270
rect 42838 664213 42890 664219
rect 42838 664155 42890 664161
rect 42836 664030 42892 664039
rect 42836 663965 42892 663974
rect 42742 661179 42794 661185
rect 42742 661121 42794 661127
rect 42070 659699 42122 659705
rect 42070 659641 42122 659647
rect 42358 659699 42410 659705
rect 42358 659641 42410 659647
rect 42082 659414 42110 659641
rect 42166 657997 42218 658003
rect 42166 657939 42218 657945
rect 42178 657564 42206 657939
rect 42850 657485 42878 663965
rect 42946 658003 42974 664261
rect 43042 661703 43070 666185
rect 43138 665921 43166 668521
rect 43126 665915 43178 665921
rect 43126 665857 43178 665863
rect 43222 665693 43274 665699
rect 43222 665635 43274 665641
rect 43124 665510 43180 665519
rect 43124 665445 43180 665454
rect 43030 661697 43082 661703
rect 43030 661639 43082 661645
rect 43028 661514 43084 661523
rect 43028 661449 43084 661458
rect 42934 657997 42986 658003
rect 42934 657939 42986 657945
rect 42166 657479 42218 657485
rect 42166 657421 42218 657427
rect 42838 657479 42890 657485
rect 42838 657421 42890 657427
rect 42178 656898 42206 657421
rect 43042 656819 43070 661449
rect 43138 660297 43166 665445
rect 43126 660291 43178 660297
rect 43126 660233 43178 660239
rect 43234 659409 43262 665635
rect 43222 659403 43274 659409
rect 43222 659345 43274 659351
rect 42166 656813 42218 656819
rect 42166 656755 42218 656761
rect 43030 656813 43082 656819
rect 43030 656755 43082 656761
rect 42178 656277 42206 656755
rect 42166 656147 42218 656153
rect 42166 656089 42218 656095
rect 42178 655714 42206 656089
rect 41588 644938 41644 644947
rect 41588 644873 41590 644882
rect 41642 644873 41644 644882
rect 41590 644841 41642 644847
rect 41588 644346 41644 644355
rect 41588 644281 41590 644290
rect 41642 644281 41644 644290
rect 41590 644249 41642 644255
rect 41780 644050 41836 644059
rect 41780 643985 41782 643994
rect 41834 643985 41836 643994
rect 41782 643953 41834 643959
rect 41590 643789 41642 643795
rect 41588 643754 41590 643763
rect 41642 643754 41644 643763
rect 41588 643689 41644 643698
rect 41588 642866 41644 642875
rect 41588 642801 41590 642810
rect 41642 642801 41644 642810
rect 43222 642827 43274 642833
rect 41590 642769 41642 642775
rect 43222 642769 43274 642775
rect 43126 642531 43178 642537
rect 43126 642473 43178 642479
rect 43138 642283 43166 642473
rect 43124 642274 43180 642283
rect 43124 642209 43180 642218
rect 41588 641386 41644 641395
rect 41588 641321 41590 641330
rect 41642 641321 41644 641330
rect 41590 641289 41642 641295
rect 41588 639906 41644 639915
rect 41588 639841 41644 639850
rect 41602 639725 41630 639841
rect 41590 639719 41642 639725
rect 41590 639661 41642 639667
rect 43030 639719 43082 639725
rect 43030 639661 43082 639667
rect 41876 637982 41932 637991
rect 41876 637917 41932 637926
rect 41780 636132 41836 636141
rect 41780 636067 41836 636076
rect 41794 634249 41822 636067
rect 41782 634243 41834 634249
rect 41782 634185 41834 634191
rect 41780 634134 41836 634143
rect 41780 634069 41836 634078
rect 41794 633953 41822 634069
rect 41782 633947 41834 633953
rect 41782 633889 41834 633895
rect 41780 633542 41836 633551
rect 41780 633477 41836 633486
rect 28820 632802 28876 632811
rect 28820 632737 28876 632746
rect 28834 632367 28862 632737
rect 41794 632589 41822 633477
rect 41780 632580 41836 632589
rect 41780 632515 41782 632524
rect 41834 632515 41836 632524
rect 41782 632483 41834 632489
rect 28820 632358 28876 632367
rect 28820 632293 28876 632302
rect 41890 628033 41918 637917
rect 42934 633947 42986 633953
rect 42934 633889 42986 633895
rect 41878 628027 41930 628033
rect 41878 627969 41930 627975
rect 42838 627879 42890 627885
rect 42838 627821 42890 627827
rect 41878 627805 41930 627811
rect 41878 627747 41930 627753
rect 41890 627224 41918 627747
rect 42166 625955 42218 625961
rect 42166 625897 42218 625903
rect 42178 625405 42206 625897
rect 42850 625295 42878 627821
rect 42946 626553 42974 633889
rect 42934 626547 42986 626553
rect 42934 626489 42986 626495
rect 42932 625994 42988 626003
rect 43042 625961 43070 639661
rect 43126 634243 43178 634249
rect 43126 634185 43178 634191
rect 43138 626701 43166 634185
rect 43126 626695 43178 626701
rect 43126 626637 43178 626643
rect 43126 626547 43178 626553
rect 43126 626489 43178 626495
rect 42932 625929 42988 625938
rect 43030 625955 43082 625961
rect 42070 625289 42122 625295
rect 42070 625231 42122 625237
rect 42838 625289 42890 625295
rect 42838 625231 42890 625237
rect 42082 624782 42110 625231
rect 42836 625106 42892 625115
rect 42836 625041 42892 625050
rect 42166 624105 42218 624111
rect 42166 624047 42218 624053
rect 42178 623565 42206 624047
rect 42070 622699 42122 622705
rect 42070 622641 42122 622647
rect 42082 622369 42110 622641
rect 42178 622557 42206 622932
rect 42166 622551 42218 622557
rect 42166 622493 42218 622499
rect 42850 622261 42878 625041
rect 42070 622255 42122 622261
rect 42070 622197 42122 622203
rect 42838 622255 42890 622261
rect 42838 622197 42890 622203
rect 42082 621748 42110 622197
rect 42836 622146 42892 622155
rect 42836 622081 42892 622090
rect 42166 621515 42218 621521
rect 42166 621457 42218 621463
rect 42178 621082 42206 621457
rect 42164 620814 42220 620823
rect 42164 620749 42220 620758
rect 42178 620529 42206 620749
rect 42850 618487 42878 622081
rect 42946 621521 42974 625929
rect 43030 625897 43082 625903
rect 43030 625807 43082 625813
rect 43030 625749 43082 625755
rect 43042 624111 43070 625749
rect 43030 624105 43082 624111
rect 43030 624047 43082 624053
rect 43028 623922 43084 623931
rect 43028 623857 43084 623866
rect 42934 621515 42986 621521
rect 42934 621457 42986 621463
rect 42932 621406 42988 621415
rect 42932 621341 42988 621350
rect 42166 618481 42218 618487
rect 42166 618423 42218 618429
rect 42838 618481 42890 618487
rect 42838 618423 42890 618429
rect 42178 618048 42206 618423
rect 42166 617815 42218 617821
rect 42166 617757 42218 617763
rect 42178 617382 42206 617757
rect 42164 617262 42220 617271
rect 42164 617197 42220 617206
rect 42178 616757 42206 617197
rect 41780 616670 41836 616679
rect 41780 616605 41836 616614
rect 41794 616198 41822 616605
rect 42838 616409 42890 616415
rect 42838 616351 42890 616357
rect 42166 614855 42218 614861
rect 42166 614797 42218 614803
rect 42178 614348 42206 614797
rect 42166 614263 42218 614269
rect 42166 614205 42218 614211
rect 42178 613721 42206 614205
rect 42070 613523 42122 613529
rect 42070 613465 42122 613471
rect 42082 613090 42110 613465
rect 42850 613011 42878 616351
rect 42946 614861 42974 621341
rect 43042 617821 43070 623857
rect 43138 622705 43166 626489
rect 43126 622699 43178 622705
rect 43126 622641 43178 622647
rect 43124 621998 43180 622007
rect 43124 621933 43180 621942
rect 43030 617815 43082 617821
rect 43030 617757 43082 617763
rect 43028 617706 43084 617715
rect 43028 617641 43084 617650
rect 42934 614855 42986 614861
rect 42934 614797 42986 614803
rect 43042 613529 43070 617641
rect 43138 614269 43166 621933
rect 43126 614263 43178 614269
rect 43126 614205 43178 614211
rect 43030 613523 43082 613529
rect 43030 613465 43082 613471
rect 42166 613005 42218 613011
rect 42166 612947 42218 612953
rect 42838 613005 42890 613011
rect 42838 612947 42890 612953
rect 42178 612498 42206 612947
rect 40340 601722 40396 601731
rect 40340 601657 40396 601666
rect 39766 599463 39818 599469
rect 39766 599405 39818 599411
rect 39778 598031 39806 599405
rect 40354 599247 40382 601657
rect 41588 601574 41644 601583
rect 41588 601509 41644 601518
rect 40342 599241 40394 599247
rect 40342 599183 40394 599189
rect 40354 598771 40382 599183
rect 41602 599099 41630 601509
rect 41780 601426 41836 601435
rect 41780 601361 41782 601370
rect 41834 601361 41836 601370
rect 41782 601329 41834 601335
rect 41780 600834 41836 600843
rect 41780 600769 41782 600778
rect 41834 600769 41836 600778
rect 41782 600737 41834 600743
rect 43234 600431 43262 642769
rect 43426 642315 43454 679666
rect 43522 643795 43550 685985
rect 43510 643789 43562 643795
rect 43510 643731 43562 643737
rect 43414 642309 43466 642315
rect 43414 642251 43466 642257
rect 43318 641347 43370 641353
rect 43318 641289 43370 641295
rect 43330 600505 43358 641289
rect 43426 641099 43454 642251
rect 43412 641090 43468 641099
rect 43412 641025 43468 641034
rect 43414 622551 43466 622557
rect 43414 622493 43466 622499
rect 43426 616267 43454 622493
rect 43414 616261 43466 616267
rect 43414 616203 43466 616209
rect 43318 600499 43370 600505
rect 43318 600441 43370 600447
rect 41782 600425 41834 600431
rect 41780 600390 41782 600399
rect 43222 600425 43274 600431
rect 41834 600390 41836 600399
rect 43222 600367 43274 600373
rect 41780 600325 41836 600334
rect 41780 599872 41836 599881
rect 41780 599807 41782 599816
rect 41834 599807 41836 599816
rect 43222 599833 43274 599839
rect 41782 599775 41834 599781
rect 43222 599775 43274 599781
rect 41780 599354 41836 599363
rect 41780 599289 41782 599298
rect 41834 599289 41836 599298
rect 41782 599257 41834 599263
rect 41590 599093 41642 599099
rect 41590 599035 41642 599041
rect 40340 598762 40396 598771
rect 40340 598697 40396 598706
rect 41780 598392 41836 598401
rect 41780 598327 41782 598336
rect 41834 598327 41836 598336
rect 41782 598295 41834 598301
rect 39764 598022 39820 598031
rect 39764 597957 39820 597966
rect 41588 596690 41644 596699
rect 41588 596625 41590 596634
rect 41642 596625 41644 596634
rect 43126 596651 43178 596657
rect 41590 596593 41642 596599
rect 43126 596593 43178 596599
rect 41876 594840 41932 594849
rect 41876 594775 41932 594784
rect 41780 592990 41836 592999
rect 41780 592925 41836 592934
rect 41794 591033 41822 592925
rect 41782 591027 41834 591033
rect 41782 590969 41834 590975
rect 41780 590918 41836 590927
rect 41780 590853 41782 590862
rect 41834 590853 41836 590862
rect 41782 590821 41834 590827
rect 28820 589586 28876 589595
rect 28820 589521 28876 589530
rect 28834 589151 28862 589521
rect 28820 589142 28876 589151
rect 28820 589077 28876 589086
rect 41588 589142 41644 589151
rect 41588 589077 41644 589086
rect 41602 587555 41630 589077
rect 41590 587549 41642 587555
rect 41590 587491 41642 587497
rect 41890 584817 41918 594775
rect 43030 591027 43082 591033
rect 43030 590969 43082 590975
rect 42934 590879 42986 590885
rect 42934 590821 42986 590827
rect 41878 584811 41930 584817
rect 41878 584753 41930 584759
rect 42838 584737 42890 584743
rect 42838 584679 42890 584685
rect 41878 584589 41930 584595
rect 41878 584531 41930 584537
rect 41890 584045 41918 584531
rect 42452 583074 42508 583083
rect 42452 583009 42508 583018
rect 42070 582739 42122 582745
rect 42070 582681 42122 582687
rect 42082 582232 42110 582681
rect 42070 582073 42122 582079
rect 42070 582015 42122 582021
rect 42082 581566 42110 582015
rect 42070 580889 42122 580895
rect 42070 580831 42122 580837
rect 42082 580382 42110 580831
rect 42082 579489 42110 579716
rect 42166 579631 42218 579637
rect 42166 579573 42218 579579
rect 42070 579483 42122 579489
rect 42070 579425 42122 579431
rect 42178 579169 42206 579573
rect 42466 579045 42494 583009
rect 42850 582079 42878 584679
rect 42838 582073 42890 582079
rect 42838 582015 42890 582021
rect 42836 581742 42892 581751
rect 42836 581677 42892 581686
rect 42070 579039 42122 579045
rect 42070 578981 42122 578987
rect 42454 579039 42506 579045
rect 42454 578981 42506 578987
rect 42082 578532 42110 578981
rect 42452 578930 42508 578939
rect 42452 578865 42508 578874
rect 42166 578299 42218 578305
rect 42166 578241 42218 578247
rect 42178 577866 42206 578241
rect 42070 577559 42122 577565
rect 42070 577501 42122 577507
rect 42082 577348 42110 577501
rect 42356 576118 42412 576127
rect 42356 576053 42412 576062
rect 42166 575265 42218 575271
rect 42166 575207 42218 575213
rect 42178 574832 42206 575207
rect 42166 574747 42218 574753
rect 42166 574689 42218 574695
rect 42178 574201 42206 574689
rect 42070 574081 42122 574087
rect 42070 574023 42122 574029
rect 42082 573574 42110 574023
rect 42370 573347 42398 576053
rect 42466 575271 42494 578865
rect 42454 575265 42506 575271
rect 42454 575207 42506 575213
rect 42850 574087 42878 581677
rect 42946 579637 42974 590821
rect 43042 580895 43070 590969
rect 43138 582745 43166 596593
rect 43126 582739 43178 582745
rect 43126 582681 43178 582687
rect 43124 582630 43180 582639
rect 43124 582565 43180 582574
rect 43030 580889 43082 580895
rect 43030 580831 43082 580837
rect 43138 580692 43166 582565
rect 43042 580664 43166 580692
rect 42934 579631 42986 579637
rect 42934 579573 42986 579579
rect 42932 579522 42988 579531
rect 42932 579457 42988 579466
rect 42946 577565 42974 579457
rect 43042 578305 43070 580664
rect 43124 580558 43180 580567
rect 43124 580493 43180 580502
rect 43030 578299 43082 578305
rect 43030 578241 43082 578247
rect 42934 577559 42986 577565
rect 42934 577501 42986 577507
rect 43028 576414 43084 576423
rect 43028 576349 43084 576358
rect 42932 576266 42988 576275
rect 42932 576201 42988 576210
rect 42838 574081 42890 574087
rect 42838 574023 42890 574029
rect 42836 573898 42892 573907
rect 42836 573833 42892 573842
rect 42358 573341 42410 573347
rect 42358 573283 42410 573289
rect 42166 573267 42218 573273
rect 42166 573209 42218 573215
rect 42178 572982 42206 573209
rect 42070 571047 42122 571053
rect 42070 570989 42122 570995
rect 42082 570540 42110 570989
rect 42178 570979 42206 571165
rect 42166 570973 42218 570979
rect 42166 570915 42218 570921
rect 42850 570313 42878 573833
rect 42946 571053 42974 576201
rect 42934 571047 42986 571053
rect 42934 570989 42986 570995
rect 43042 570979 43070 576349
rect 43138 574753 43166 580493
rect 43126 574747 43178 574753
rect 43126 574689 43178 574695
rect 43030 570973 43082 570979
rect 43030 570915 43082 570921
rect 42166 570307 42218 570313
rect 42166 570249 42218 570255
rect 42838 570307 42890 570313
rect 42838 570249 42890 570255
rect 42178 569874 42206 570249
rect 42166 569789 42218 569795
rect 42166 569731 42218 569737
rect 42178 569325 42206 569731
rect 42934 541595 42986 541601
rect 42934 541537 42986 541543
rect 42838 541521 42890 541527
rect 42838 541463 42890 541469
rect 41794 540459 41822 540866
rect 41780 540450 41836 540459
rect 41780 540385 41836 540394
rect 41794 538831 41822 539016
rect 41780 538822 41836 538831
rect 41780 538757 41836 538766
rect 42166 538487 42218 538493
rect 42166 538429 42218 538435
rect 42178 538350 42206 538429
rect 41794 536907 41822 537166
rect 42850 537087 42878 541463
rect 42946 538493 42974 541537
rect 42934 538487 42986 538493
rect 42934 538429 42986 538435
rect 42166 537081 42218 537087
rect 42166 537023 42218 537029
rect 42838 537081 42890 537087
rect 42838 537023 42890 537029
rect 41780 536898 41836 536907
rect 41780 536833 41836 536842
rect 42178 536500 42206 537023
rect 42178 535755 42206 535982
rect 42166 535749 42218 535755
rect 42166 535691 42218 535697
rect 41794 534835 41822 535316
rect 41780 534826 41836 534835
rect 41780 534761 41836 534770
rect 41794 534539 41822 534681
rect 41780 534530 41836 534539
rect 41780 534465 41836 534474
rect 41890 533651 41918 534132
rect 41876 533642 41932 533651
rect 41876 533577 41932 533586
rect 41794 531431 41822 531645
rect 41780 531422 41836 531431
rect 41780 531357 41836 531366
rect 41794 530691 41822 531024
rect 41780 530682 41836 530691
rect 41780 530617 41836 530626
rect 41794 530099 41822 530358
rect 41780 530090 41836 530099
rect 41780 530025 41836 530034
rect 42178 529359 42206 529805
rect 42164 529350 42220 529359
rect 42164 529285 42220 529294
rect 42178 527731 42206 527990
rect 42164 527722 42220 527731
rect 42164 527657 42220 527666
rect 42082 527139 42110 527324
rect 42068 527130 42124 527139
rect 42068 527065 42124 527074
rect 42082 526547 42110 526658
rect 42068 526538 42124 526547
rect 42068 526473 42124 526482
rect 42070 526425 42122 526431
rect 42070 526367 42122 526373
rect 42082 526140 42110 526367
rect 41782 476105 41834 476111
rect 41780 476070 41782 476079
rect 41834 476070 41836 476079
rect 41780 476005 41836 476014
rect 41782 475587 41834 475593
rect 41780 475552 41782 475561
rect 41834 475552 41836 475561
rect 41780 475487 41836 475496
rect 41780 475034 41836 475043
rect 41780 474969 41836 474978
rect 40340 473850 40396 473859
rect 40340 473785 40396 473794
rect 39668 472370 39724 472379
rect 39668 472305 39724 472314
rect 34484 464378 34540 464387
rect 34484 464313 34540 464322
rect 23060 463786 23116 463795
rect 23060 463721 23116 463730
rect 23074 463351 23102 463721
rect 23060 463342 23116 463351
rect 23060 463277 23116 463286
rect 34498 463161 34526 464313
rect 34486 463155 34538 463161
rect 34486 463097 34538 463103
rect 39682 426309 39710 472305
rect 40354 427979 40382 473785
rect 41684 473258 41740 473267
rect 41684 473193 41740 473202
rect 41590 465301 41642 465307
rect 41588 465266 41590 465275
rect 41642 465266 41644 465275
rect 41588 465201 41644 465210
rect 41698 432081 41726 473193
rect 41794 472411 41822 474969
rect 43234 474631 43262 599775
rect 43330 599469 43358 600441
rect 43318 599463 43370 599469
rect 43318 599405 43370 599411
rect 43318 599315 43370 599321
rect 43318 599257 43370 599263
rect 41878 474625 41930 474631
rect 41876 474590 41878 474599
rect 43222 474625 43274 474631
rect 41930 474590 41932 474599
rect 43222 474567 43274 474573
rect 41876 474525 41932 474534
rect 43330 473119 43358 599257
rect 43414 535749 43466 535755
rect 43414 535691 43466 535697
rect 43316 473110 43372 473119
rect 43316 473045 43372 473054
rect 41782 472405 41834 472411
rect 41782 472347 41834 472353
rect 41780 472074 41836 472083
rect 41780 472009 41782 472018
rect 41834 472009 41836 472018
rect 41782 471977 41834 471983
rect 43426 465307 43454 535691
rect 43414 465301 43466 465307
rect 43414 465243 43466 465249
rect 41780 463638 41836 463647
rect 41780 463573 41782 463582
rect 41834 463573 41836 463582
rect 41782 463541 41834 463547
rect 41794 463161 41822 463541
rect 41782 463155 41834 463161
rect 41782 463097 41834 463103
rect 41686 432075 41738 432081
rect 41686 432017 41738 432023
rect 41588 428562 41644 428571
rect 41588 428497 41590 428506
rect 41642 428497 41644 428506
rect 41590 428465 41642 428471
rect 40340 427970 40396 427979
rect 40340 427905 40396 427914
rect 41588 427082 41644 427091
rect 41588 427017 41590 427026
rect 41642 427017 41644 427026
rect 41590 426985 41642 426991
rect 41698 426499 41726 432017
rect 41780 429302 41836 429311
rect 41780 429237 41782 429246
rect 41834 429237 41836 429246
rect 41782 429205 41834 429211
rect 41780 428266 41836 428275
rect 41780 428201 41782 428210
rect 41834 428201 41836 428210
rect 41782 428169 41834 428175
rect 43318 427043 43370 427049
rect 43318 426985 43370 426991
rect 41780 426712 41836 426721
rect 41780 426647 41782 426656
rect 41834 426647 41836 426656
rect 43222 426673 43274 426679
rect 41782 426615 41834 426621
rect 43222 426615 43274 426621
rect 41684 426490 41740 426499
rect 41684 426425 41740 426434
rect 39670 426303 39722 426309
rect 39670 426245 39722 426251
rect 41686 426303 41738 426309
rect 41686 426245 41738 426251
rect 41588 425602 41644 425611
rect 41588 425537 41644 425546
rect 41602 420463 41630 425537
rect 41698 425019 41726 426245
rect 41684 425010 41740 425019
rect 41684 424945 41740 424954
rect 41590 420457 41642 420463
rect 41590 420399 41642 420405
rect 41588 420126 41644 420135
rect 41588 420061 41644 420070
rect 41602 417873 41630 420061
rect 41590 417867 41642 417873
rect 41590 417809 41642 417815
rect 28916 417018 28972 417027
rect 28916 416953 28972 416962
rect 28930 416583 28958 416953
rect 28916 416574 28972 416583
rect 28916 416509 28972 416518
rect 41588 416574 41644 416583
rect 41588 416509 41590 416518
rect 41642 416509 41644 416518
rect 41590 416477 41642 416483
rect 41698 414691 41726 424945
rect 41780 422198 41836 422207
rect 41780 422133 41836 422142
rect 41686 414685 41738 414691
rect 41686 414627 41738 414633
rect 41794 413877 41822 422133
rect 42838 417867 42890 417873
rect 42838 417809 42890 417815
rect 41782 413871 41834 413877
rect 41782 413813 41834 413819
rect 41782 413575 41834 413581
rect 41782 413517 41834 413523
rect 41794 413068 41822 413517
rect 41876 411690 41932 411699
rect 41876 411625 41932 411634
rect 41890 411218 41918 411625
rect 42082 410177 42110 410552
rect 42070 410171 42122 410177
rect 42070 410113 42122 410119
rect 42742 410171 42794 410177
rect 42742 410113 42794 410119
rect 42166 409875 42218 409881
rect 42166 409817 42218 409823
rect 42178 409368 42206 409817
rect 41780 408434 41836 408443
rect 41780 408369 41836 408378
rect 41794 408184 41822 408369
rect 42082 408327 42110 408702
rect 42070 408321 42122 408327
rect 42070 408263 42122 408269
rect 41780 407990 41836 407999
rect 41780 407925 41836 407934
rect 41794 407518 41822 407925
rect 42164 407398 42220 407407
rect 42164 407333 42220 407342
rect 42178 406881 42206 407333
rect 42068 406510 42124 406519
rect 42068 406445 42124 406454
rect 42082 406334 42110 406445
rect 42754 406107 42782 410113
rect 42850 409881 42878 417809
rect 42838 409875 42890 409881
rect 42838 409817 42890 409823
rect 42838 408321 42890 408327
rect 42838 408263 42890 408269
rect 42742 406101 42794 406107
rect 42742 406043 42794 406049
rect 41780 404290 41836 404299
rect 41780 404225 41836 404234
rect 41794 403818 41822 404225
rect 41780 403698 41836 403707
rect 41780 403633 41836 403642
rect 41794 403226 41822 403633
rect 41780 402958 41836 402967
rect 41780 402893 41836 402902
rect 41794 402560 41822 402893
rect 42850 402851 42878 408263
rect 42838 402845 42890 402851
rect 42838 402787 42890 402793
rect 41780 402366 41836 402375
rect 41780 402301 41836 402310
rect 41794 402005 41822 402301
rect 41876 400294 41932 400303
rect 41876 400229 41932 400238
rect 41890 400192 41918 400229
rect 41780 399850 41836 399859
rect 41780 399785 41836 399794
rect 41794 399526 41822 399785
rect 42164 399406 42220 399415
rect 42164 399341 42220 399350
rect 42178 398860 42206 399341
rect 42178 394563 42206 398342
rect 42166 394557 42218 394563
rect 42166 394499 42218 394505
rect 41780 386086 41836 386095
rect 41780 386021 41782 386030
rect 41834 386021 41836 386030
rect 41782 385989 41834 385995
rect 41588 385346 41644 385355
rect 41588 385281 41590 385290
rect 41642 385281 41644 385290
rect 41590 385249 41642 385255
rect 41780 385050 41836 385059
rect 41780 384985 41782 384994
rect 41834 384985 41836 384994
rect 41782 384953 41834 384959
rect 41590 384789 41642 384795
rect 41588 384754 41590 384763
rect 41642 384754 41644 384763
rect 41588 384689 41644 384698
rect 41588 383866 41644 383875
rect 41588 383801 41590 383810
rect 41642 383801 41644 383810
rect 41590 383769 41642 383775
rect 41780 383570 41836 383579
rect 41780 383505 41782 383514
rect 41834 383505 41836 383514
rect 41782 383473 41834 383479
rect 43234 383315 43262 426615
rect 43330 384795 43358 426985
rect 43414 420457 43466 420463
rect 43414 420399 43466 420405
rect 43318 384789 43370 384795
rect 43318 384731 43370 384737
rect 43318 383827 43370 383833
rect 43318 383769 43370 383775
rect 41590 383309 41642 383315
rect 41588 383274 41590 383283
rect 43222 383309 43274 383315
rect 41642 383274 41644 383283
rect 43222 383251 43274 383257
rect 41588 383209 41644 383218
rect 39956 382238 40012 382247
rect 39956 382173 40012 382182
rect 39970 377247 39998 382173
rect 41782 382051 41834 382057
rect 41780 382016 41782 382025
rect 41834 382016 41836 382025
rect 41780 381951 41836 381960
rect 41780 378982 41836 378991
rect 41780 378917 41836 378926
rect 39958 377241 40010 377247
rect 39958 377183 40010 377189
rect 41588 376910 41644 376919
rect 41588 376845 41644 376854
rect 41602 374509 41630 376845
rect 41590 374503 41642 374509
rect 41590 374445 41642 374451
rect 28820 373802 28876 373811
rect 28820 373737 28876 373746
rect 28834 373367 28862 373737
rect 28820 373358 28876 373367
rect 28820 373293 28876 373302
rect 41588 373358 41644 373367
rect 41588 373293 41590 373302
rect 41642 373293 41644 373302
rect 41590 373261 41642 373267
rect 41794 370661 41822 378917
rect 42838 374503 42890 374509
rect 42838 374445 42890 374451
rect 41782 370655 41834 370661
rect 41782 370597 41834 370603
rect 41782 370359 41834 370365
rect 41782 370301 41834 370307
rect 41794 369852 41822 370301
rect 42068 368474 42124 368483
rect 42068 368409 42124 368418
rect 42082 368002 42110 368409
rect 42082 366961 42110 367336
rect 42070 366955 42122 366961
rect 42070 366897 42122 366903
rect 42742 366955 42794 366961
rect 42742 366897 42794 366903
rect 42166 366733 42218 366739
rect 42166 366675 42218 366681
rect 42178 366152 42206 366675
rect 41780 365218 41836 365227
rect 41780 365153 41836 365162
rect 41794 364968 41822 365153
rect 42178 365111 42206 365521
rect 42166 365105 42218 365111
rect 42166 365047 42218 365053
rect 41972 364626 42028 364635
rect 41972 364561 42028 364570
rect 41986 364302 42014 364561
rect 41780 364182 41836 364191
rect 41780 364117 41836 364126
rect 41794 363681 41822 364117
rect 42164 363590 42220 363599
rect 42164 363525 42220 363534
rect 42178 363118 42206 363525
rect 42754 362595 42782 366897
rect 42850 366739 42878 374445
rect 42838 366733 42890 366739
rect 42838 366675 42890 366681
rect 42838 365105 42890 365111
rect 42838 365047 42890 365053
rect 42742 362589 42794 362595
rect 42742 362531 42794 362537
rect 41780 361074 41836 361083
rect 41780 361009 41836 361018
rect 41794 360645 41822 361009
rect 41780 360482 41836 360491
rect 41780 360417 41836 360426
rect 41794 360010 41822 360417
rect 42850 360005 42878 365047
rect 42838 359999 42890 360005
rect 42838 359941 42890 359947
rect 41780 359742 41836 359751
rect 41780 359677 41836 359686
rect 41794 359344 41822 359677
rect 42068 359002 42124 359011
rect 42068 358937 42124 358946
rect 42082 358826 42110 358937
rect 41780 357226 41836 357235
rect 41780 357161 41836 357170
rect 41794 356976 41822 357161
rect 41780 356634 41836 356643
rect 41780 356569 41836 356578
rect 41794 356310 41822 356569
rect 42164 356190 42220 356199
rect 42164 356125 42220 356134
rect 42178 355677 42206 356125
rect 42178 351347 42206 355126
rect 42166 351341 42218 351347
rect 42166 351283 42218 351289
rect 41780 342870 41836 342879
rect 41780 342805 41782 342814
rect 41834 342805 41836 342814
rect 41782 342773 41834 342779
rect 41780 342352 41836 342361
rect 41780 342287 41782 342296
rect 41834 342287 41836 342296
rect 41782 342255 41834 342261
rect 41780 341834 41836 341843
rect 41780 341769 41782 341778
rect 41834 341769 41836 341778
rect 41782 341737 41834 341743
rect 43330 341431 43358 383769
rect 43426 382057 43454 420399
rect 43510 383531 43562 383537
rect 43510 383473 43562 383479
rect 43414 382051 43466 382057
rect 43414 381993 43466 381999
rect 43414 377241 43466 377247
rect 43414 377183 43466 377189
rect 41782 341425 41834 341431
rect 41780 341390 41782 341399
rect 43318 341425 43370 341431
rect 41834 341390 41836 341399
rect 43318 341367 43370 341373
rect 41780 341325 41836 341334
rect 41588 340650 41644 340659
rect 41588 340585 41590 340594
rect 41642 340585 41644 340594
rect 43222 340611 43274 340617
rect 41590 340553 41642 340559
rect 43222 340553 43274 340559
rect 41780 340354 41836 340363
rect 41780 340289 41782 340298
rect 41834 340289 41836 340298
rect 41782 340257 41834 340263
rect 41590 340093 41642 340099
rect 41588 340058 41590 340067
rect 41642 340058 41644 340067
rect 41588 339993 41644 340002
rect 41588 339170 41644 339179
rect 41588 339105 41590 339114
rect 41642 339105 41644 339114
rect 41590 339073 41642 339079
rect 41782 338909 41834 338915
rect 41780 338874 41782 338883
rect 41834 338874 41836 338883
rect 41780 338809 41836 338818
rect 34484 335618 34540 335627
rect 34484 335553 34540 335562
rect 28820 330586 28876 330595
rect 28820 330521 28876 330530
rect 28834 330151 28862 330521
rect 28820 330142 28876 330151
rect 28820 330077 28876 330086
rect 34498 329813 34526 335553
rect 41780 330438 41836 330447
rect 41780 330373 41782 330382
rect 41834 330373 41836 330382
rect 41782 330341 41834 330347
rect 34486 329807 34538 329813
rect 34486 329749 34538 329755
rect 41782 329807 41834 329813
rect 41782 329749 41834 329755
rect 41794 327223 41822 329749
rect 41782 327217 41834 327223
rect 41782 327159 41834 327165
rect 41782 326995 41834 327001
rect 41782 326937 41834 326943
rect 41794 326445 41822 326937
rect 41780 325110 41836 325119
rect 41780 325045 41836 325054
rect 41794 324605 41822 325045
rect 42178 323597 42206 323972
rect 42166 323591 42218 323597
rect 42166 323533 42218 323539
rect 42454 323591 42506 323597
rect 42454 323533 42506 323539
rect 41780 323334 41836 323343
rect 41780 323269 41836 323278
rect 41794 322788 41822 323269
rect 41780 321854 41836 321863
rect 41780 321789 41836 321798
rect 41794 321569 41822 321789
rect 42178 321747 42206 322122
rect 42166 321741 42218 321747
rect 42166 321683 42218 321689
rect 42068 321262 42124 321271
rect 42068 321197 42124 321206
rect 42082 320938 42110 321197
rect 41876 320818 41932 320827
rect 41876 320753 41932 320762
rect 41890 320272 41918 320753
rect 42068 319930 42124 319939
rect 42068 319865 42124 319874
rect 42082 319754 42110 319865
rect 42466 319675 42494 323533
rect 42838 321741 42890 321747
rect 42838 321683 42890 321689
rect 42454 319669 42506 319675
rect 42454 319611 42506 319617
rect 41876 317710 41932 317719
rect 41876 317645 41932 317654
rect 41890 317238 41918 317645
rect 41780 316822 41836 316831
rect 42850 316789 42878 321683
rect 41780 316757 41836 316766
rect 42838 316783 42890 316789
rect 41794 316601 41822 316757
rect 42838 316725 42890 316731
rect 41780 316230 41836 316239
rect 41780 316165 41836 316174
rect 41794 315980 41822 316165
rect 41780 315638 41836 315647
rect 41780 315573 41836 315582
rect 41794 315388 41822 315573
rect 42164 313862 42220 313871
rect 42164 313797 42220 313806
rect 42178 313538 42206 313797
rect 41780 313270 41836 313279
rect 41780 313205 41836 313214
rect 41794 312946 41822 313205
rect 41780 312678 41836 312687
rect 41780 312613 41836 312622
rect 41794 312280 41822 312613
rect 42178 308131 42206 311725
rect 42166 308125 42218 308131
rect 42166 308067 42218 308073
rect 39670 299689 39722 299695
rect 39670 299631 39722 299637
rect 41780 299654 41836 299663
rect 39682 296555 39710 299631
rect 41780 299589 41782 299598
rect 41834 299589 41836 299598
rect 41782 299557 41834 299563
rect 41588 298766 41644 298775
rect 41588 298701 41644 298710
rect 39862 296803 39914 296809
rect 39862 296745 39914 296751
rect 39668 296546 39724 296555
rect 39668 296481 39724 296490
rect 39874 295963 39902 296745
rect 41602 296735 41630 298701
rect 41780 298618 41836 298627
rect 41780 298553 41782 298562
rect 41834 298553 41836 298562
rect 41782 298521 41834 298527
rect 43234 298215 43262 340553
rect 43426 338915 43454 377183
rect 43522 340099 43550 383473
rect 43510 340093 43562 340099
rect 43510 340035 43562 340041
rect 44374 340093 44426 340099
rect 44374 340035 44426 340041
rect 43414 338909 43466 338915
rect 43414 338851 43466 338857
rect 41782 298209 41834 298215
rect 41780 298174 41782 298183
rect 43222 298209 43274 298215
rect 41834 298174 41836 298183
rect 43222 298151 43274 298157
rect 41780 298109 41836 298118
rect 41780 297656 41836 297665
rect 41780 297591 41782 297600
rect 41834 297591 41836 297600
rect 43222 297617 43274 297623
rect 41782 297559 41834 297565
rect 43222 297559 43274 297565
rect 41780 297138 41836 297147
rect 41780 297073 41782 297082
rect 41834 297073 41836 297082
rect 41782 297041 41834 297047
rect 41590 296729 41642 296735
rect 41590 296671 41642 296677
rect 39860 295954 39916 295963
rect 39860 295889 39916 295898
rect 41588 295954 41644 295963
rect 41588 295889 41590 295898
rect 41642 295889 41644 295898
rect 41590 295857 41642 295863
rect 34484 292402 34540 292411
rect 34484 292337 34540 292346
rect 28820 287370 28876 287379
rect 28820 287305 28876 287314
rect 28834 286935 28862 287305
rect 28820 286926 28876 286935
rect 28820 286861 28876 286870
rect 34498 286597 34526 292337
rect 41780 287222 41836 287231
rect 41780 287157 41782 287166
rect 41834 287157 41836 287166
rect 41782 287125 41834 287131
rect 34486 286591 34538 286597
rect 34486 286533 34538 286539
rect 41782 286591 41834 286597
rect 41782 286533 41834 286539
rect 41794 284081 41822 286533
rect 41782 284075 41834 284081
rect 41782 284017 41834 284023
rect 41782 283779 41834 283785
rect 41782 283721 41834 283727
rect 41794 283272 41822 283721
rect 42068 281894 42124 281903
rect 42068 281829 42124 281838
rect 42082 281422 42110 281829
rect 42166 281337 42218 281343
rect 42166 281279 42218 281285
rect 42178 280756 42206 281279
rect 41780 280118 41836 280127
rect 41780 280053 41836 280062
rect 41794 279572 41822 280053
rect 42166 279339 42218 279345
rect 42166 279281 42218 279287
rect 42178 278906 42206 279281
rect 41780 278786 41836 278795
rect 41780 278721 41836 278730
rect 41794 278388 41822 278721
rect 42068 278046 42124 278055
rect 42068 277981 42124 277990
rect 42082 277722 42110 277981
rect 41876 277602 41932 277611
rect 41876 277537 41932 277546
rect 41890 277056 41918 277537
rect 42068 276714 42124 276723
rect 42068 276649 42124 276658
rect 42082 276538 42110 276649
rect 41780 274494 41836 274503
rect 41780 274429 41836 274438
rect 41794 274022 41822 274429
rect 41780 273606 41836 273615
rect 41780 273541 41836 273550
rect 41794 273401 41822 273541
rect 41780 273310 41836 273319
rect 41780 273245 41836 273254
rect 41794 272764 41822 273245
rect 41780 272422 41836 272431
rect 41780 272357 41836 272366
rect 41794 272205 41822 272357
rect 41876 270646 41932 270655
rect 41876 270581 41932 270590
rect 41890 270365 41918 270581
rect 41780 270054 41836 270063
rect 41780 269989 41836 269998
rect 41794 269730 41822 269989
rect 42164 269610 42220 269619
rect 42164 269545 42220 269554
rect 42178 269064 42206 269545
rect 42070 268831 42122 268837
rect 42070 268773 42122 268779
rect 42082 268546 42110 268773
rect 23062 265057 23114 265063
rect 23062 264999 23114 265005
rect 23074 253339 23102 264999
rect 23350 263651 23402 263657
rect 23350 263593 23402 263599
rect 23254 263577 23306 263583
rect 23254 263519 23306 263525
rect 23158 262171 23210 262177
rect 23158 262113 23210 262119
rect 23170 254227 23198 262113
rect 23156 254218 23212 254227
rect 23156 254153 23212 254162
rect 23060 253330 23116 253339
rect 23060 253265 23116 253274
rect 23266 252747 23294 263519
rect 23362 253339 23390 263593
rect 40246 256399 40298 256405
rect 40246 256341 40298 256347
rect 40258 256299 40286 256341
rect 40244 256290 40300 256299
rect 40244 256225 40300 256234
rect 41588 255698 41644 255707
rect 41588 255633 41644 255642
rect 41602 253519 41630 255633
rect 41782 255437 41834 255443
rect 41780 255402 41782 255411
rect 41834 255402 41836 255411
rect 41780 255337 41836 255346
rect 43234 254999 43262 297559
rect 44182 290957 44234 290963
rect 44182 290899 44234 290905
rect 44194 268837 44222 290899
rect 44278 287183 44330 287189
rect 44278 287125 44330 287131
rect 44182 268831 44234 268837
rect 44182 268773 44234 268779
rect 41782 254993 41834 254999
rect 41780 254958 41782 254967
rect 43222 254993 43274 254999
rect 41834 254958 41836 254967
rect 43222 254935 43274 254941
rect 41780 254893 41836 254902
rect 41780 254514 41836 254523
rect 41780 254449 41782 254458
rect 41834 254449 41836 254458
rect 43222 254475 43274 254481
rect 41782 254417 41834 254423
rect 43222 254417 43274 254423
rect 41590 253513 41642 253519
rect 41590 253455 41642 253461
rect 23348 253330 23404 253339
rect 23348 253265 23404 253274
rect 23252 252738 23308 252747
rect 23252 252673 23308 252682
rect 41684 249186 41740 249195
rect 41684 249121 41740 249130
rect 41590 245003 41642 245009
rect 41590 244945 41642 244951
rect 41602 244755 41630 244945
rect 41588 244746 41644 244755
rect 41698 244732 41726 249121
rect 41780 244894 41836 244903
rect 41780 244829 41782 244838
rect 41834 244829 41836 244838
rect 41782 244797 41834 244803
rect 41698 244704 41822 244732
rect 41588 244681 41644 244690
rect 41588 243710 41644 243719
rect 41588 243645 41644 243654
rect 41602 242641 41630 243645
rect 41590 242635 41642 242641
rect 41590 242577 41642 242583
rect 41794 240865 41822 244704
rect 41782 240859 41834 240865
rect 41782 240801 41834 240807
rect 41782 240563 41834 240569
rect 41782 240505 41834 240511
rect 41794 240056 41822 240505
rect 42068 238678 42124 238687
rect 42068 238613 42124 238622
rect 42082 238206 42110 238613
rect 41876 236902 41932 236911
rect 41876 236837 41932 236846
rect 41890 236356 41918 236837
rect 41780 235570 41836 235579
rect 41780 235505 41836 235514
rect 41794 235172 41822 235505
rect 42164 234830 42220 234839
rect 42164 234765 42220 234774
rect 42178 234506 42206 234765
rect 42164 234386 42220 234395
rect 42164 234321 42220 234330
rect 42178 233881 42206 234321
rect 42164 233646 42220 233655
rect 42164 233581 42220 233590
rect 42178 233322 42206 233581
rect 41780 231278 41836 231287
rect 41780 231213 41836 231222
rect 41794 230845 41822 231213
rect 41780 230390 41836 230399
rect 41780 230325 41836 230334
rect 41794 230214 41822 230325
rect 41780 230094 41836 230103
rect 41780 230029 41836 230038
rect 41794 229548 41822 230029
rect 41780 229354 41836 229363
rect 41780 229289 41836 229298
rect 41794 229030 41822 229289
rect 41876 227430 41932 227439
rect 41876 227365 41932 227374
rect 41890 227180 41918 227365
rect 41780 226838 41836 226847
rect 41780 226773 41836 226782
rect 41794 226514 41822 226773
rect 42164 226394 42220 226403
rect 42164 226329 42220 226338
rect 42178 225877 42206 226329
rect 42262 226207 42314 226213
rect 42262 226149 42314 226155
rect 42274 225344 42302 226149
rect 42192 225316 42302 225344
rect 41782 213331 41834 213337
rect 41780 213296 41782 213305
rect 41834 213296 41836 213305
rect 41780 213231 41836 213240
rect 41590 212961 41642 212967
rect 41588 212926 41590 212935
rect 41642 212926 41644 212935
rect 41588 212861 41644 212870
rect 41782 212221 41834 212227
rect 41780 212186 41782 212195
rect 41834 212186 41836 212195
rect 41780 212121 41836 212130
rect 43234 211783 43262 254417
rect 44290 246267 44318 287125
rect 44386 276279 44414 340035
rect 44470 338909 44522 338915
rect 44470 338851 44522 338857
rect 44482 278499 44510 338851
rect 44468 278490 44524 278499
rect 44468 278425 44524 278434
rect 44372 276270 44428 276279
rect 44372 276205 44428 276214
rect 44578 275539 44606 813561
rect 44674 277315 44702 814819
rect 44770 785653 44798 817261
rect 44854 816579 44906 816585
rect 44854 816521 44906 816527
rect 44866 789131 44894 816521
rect 47446 805183 47498 805189
rect 47446 805125 47498 805131
rect 44854 789125 44906 789131
rect 44854 789067 44906 789073
rect 44758 785647 44810 785653
rect 44758 785589 44810 785595
rect 44758 773955 44810 773961
rect 44758 773897 44810 773903
rect 44770 742955 44798 773897
rect 44950 773511 45002 773517
rect 44950 773453 45002 773459
rect 44854 746131 44906 746137
rect 44854 746073 44906 746079
rect 44758 742949 44810 742955
rect 44758 742891 44810 742897
rect 44758 730369 44810 730375
rect 44758 730311 44810 730317
rect 44770 702625 44798 730311
rect 44758 702619 44810 702625
rect 44758 702561 44810 702567
rect 44758 685377 44810 685383
rect 44758 685319 44810 685325
rect 44660 277306 44716 277315
rect 44660 277241 44716 277250
rect 44564 275530 44620 275539
rect 44564 275465 44620 275474
rect 44770 266363 44798 685319
rect 44866 277907 44894 746073
rect 44962 745397 44990 773453
rect 44950 745391 45002 745397
rect 44950 745333 45002 745339
rect 44950 684193 45002 684199
rect 44950 684135 45002 684141
rect 44852 277898 44908 277907
rect 44852 277833 44908 277842
rect 44962 275095 44990 684135
rect 45044 658850 45100 658859
rect 45044 658785 45100 658794
rect 45058 656153 45086 658785
rect 45046 656147 45098 656153
rect 45046 656089 45098 656095
rect 45142 642309 45194 642315
rect 45142 642251 45194 642257
rect 45044 572418 45100 572427
rect 45044 572353 45100 572362
rect 45058 569795 45086 572353
rect 45046 569789 45098 569795
rect 45046 569731 45098 569737
rect 45044 529350 45100 529359
rect 45044 529285 45100 529294
rect 45058 526431 45086 529285
rect 45046 526425 45098 526431
rect 45046 526367 45098 526373
rect 45044 473110 45100 473119
rect 45044 473045 45100 473054
rect 45058 278647 45086 473045
rect 45044 278638 45100 278647
rect 45044 278573 45100 278582
rect 45154 276427 45182 642251
rect 46102 598353 46154 598359
rect 46102 598295 46154 598301
rect 46114 472060 46142 598295
rect 46018 472041 46142 472060
rect 46006 472035 46142 472041
rect 46058 472032 46142 472035
rect 46006 471977 46058 471983
rect 45334 414685 45386 414691
rect 45334 414627 45386 414633
rect 45238 383309 45290 383315
rect 45238 383251 45290 383257
rect 45140 276418 45196 276427
rect 45140 276353 45196 276362
rect 44948 275086 45004 275095
rect 44948 275021 45004 275030
rect 45250 270655 45278 383251
rect 45346 302359 45374 414627
rect 45430 382051 45482 382057
rect 45430 381993 45482 381999
rect 45334 302353 45386 302359
rect 45334 302295 45386 302301
rect 45334 282595 45386 282601
rect 45334 282537 45386 282543
rect 45236 270646 45292 270655
rect 45236 270581 45292 270590
rect 44756 266354 44812 266363
rect 44756 266289 44812 266298
rect 44278 246261 44330 246267
rect 44278 246203 44330 246209
rect 44758 244929 44810 244935
rect 44758 244871 44810 244877
rect 44662 242857 44714 242863
rect 44662 242799 44714 242805
rect 44566 242783 44618 242789
rect 44566 242725 44618 242731
rect 41782 211777 41834 211783
rect 41780 211742 41782 211751
rect 43222 211777 43274 211783
rect 41834 211742 41836 211751
rect 43222 211719 43274 211725
rect 41780 211677 41836 211686
rect 41590 211481 41642 211487
rect 41588 211446 41590 211455
rect 41642 211446 41644 211455
rect 41588 211381 41644 211390
rect 41782 210741 41834 210747
rect 41780 210706 41782 210715
rect 41834 210706 41836 210715
rect 41780 210641 41836 210650
rect 41780 210262 41836 210271
rect 41780 210197 41782 210206
rect 41834 210197 41836 210206
rect 41782 210165 41834 210171
rect 41590 210001 41642 210007
rect 41588 209966 41590 209975
rect 41642 209966 41644 209975
rect 41588 209901 41644 209910
rect 41590 209409 41642 209415
rect 41588 209374 41590 209383
rect 41642 209374 41644 209383
rect 41588 209309 41644 209318
rect 41780 206266 41836 206275
rect 41780 206201 41836 206210
rect 41590 201565 41642 201571
rect 41588 201530 41590 201539
rect 41642 201530 41644 201539
rect 41588 201465 41644 201474
rect 41590 200973 41642 200979
rect 41588 200938 41590 200947
rect 41642 200938 41644 200947
rect 41588 200873 41644 200882
rect 41794 197649 41822 206201
rect 41878 201713 41930 201719
rect 41876 201678 41878 201687
rect 41930 201678 41932 201687
rect 41876 201613 41932 201622
rect 44578 200979 44606 242725
rect 44674 201571 44702 242799
rect 44770 201719 44798 244871
rect 44854 242709 44906 242715
rect 44854 242651 44906 242657
rect 44866 211487 44894 242651
rect 44854 211481 44906 211487
rect 44854 211423 44906 211429
rect 44758 201713 44810 201719
rect 44758 201655 44810 201661
rect 44662 201565 44714 201571
rect 44662 201507 44714 201513
rect 44566 200973 44618 200979
rect 44566 200915 44618 200921
rect 41782 197643 41834 197649
rect 41782 197585 41834 197591
rect 41782 197421 41834 197427
rect 41782 197363 41834 197369
rect 41794 196840 41822 197363
rect 41876 195462 41932 195471
rect 41876 195397 41932 195406
rect 41890 194990 41918 195397
rect 41780 193686 41836 193695
rect 41780 193621 41836 193630
rect 41794 193140 41822 193621
rect 42164 192354 42220 192363
rect 42164 192289 42220 192298
rect 42178 191956 42206 192289
rect 42164 191762 42220 191771
rect 42164 191697 42220 191706
rect 42178 191325 42206 191697
rect 41780 191170 41836 191179
rect 41780 191105 41836 191114
rect 41794 190698 41822 191105
rect 41780 190430 41836 190439
rect 41780 190365 41836 190374
rect 41794 190106 41822 190365
rect 42068 188062 42124 188071
rect 42068 187997 42124 188006
rect 42082 187664 42110 187997
rect 41780 187174 41836 187183
rect 41780 187109 41836 187118
rect 41794 186998 41822 187109
rect 41780 186878 41836 186887
rect 41780 186813 41836 186822
rect 41794 186332 41822 186813
rect 41780 185990 41836 185999
rect 41780 185925 41836 185934
rect 41794 185814 41822 185925
rect 42164 184214 42220 184223
rect 42164 184149 42220 184158
rect 42178 183964 42206 184149
rect 41780 183622 41836 183631
rect 41780 183557 41836 183566
rect 41794 183298 41822 183557
rect 41876 183178 41932 183187
rect 41876 183113 41932 183122
rect 41890 182677 41918 183113
rect 45346 182405 45374 282537
rect 45442 278351 45470 381993
rect 45526 330399 45578 330405
rect 45526 330341 45578 330347
rect 45428 278342 45484 278351
rect 45428 278277 45484 278286
rect 45538 246341 45566 330341
rect 45814 288071 45866 288077
rect 45814 288013 45866 288019
rect 45622 282373 45674 282379
rect 45622 282315 45674 282321
rect 45526 246335 45578 246341
rect 45526 246277 45578 246283
rect 45634 212227 45662 282315
rect 45718 279487 45770 279493
rect 45718 279429 45770 279435
rect 45730 212967 45758 279429
rect 45826 226213 45854 288013
rect 45910 279413 45962 279419
rect 45910 279355 45962 279361
rect 45814 226207 45866 226213
rect 45814 226149 45866 226155
rect 45922 213337 45950 279355
rect 46018 278203 46046 471977
rect 46198 340315 46250 340321
rect 46198 340257 46250 340263
rect 46102 339131 46154 339137
rect 46102 339073 46154 339079
rect 46114 298141 46142 339073
rect 46210 300953 46238 340257
rect 46486 302353 46538 302359
rect 46486 302295 46538 302301
rect 46198 300947 46250 300953
rect 46198 300889 46250 300895
rect 46498 299547 46526 302295
rect 46870 300947 46922 300953
rect 46870 300889 46922 300895
rect 46882 299695 46910 300889
rect 46870 299689 46922 299695
rect 46870 299631 46922 299637
rect 46486 299541 46538 299547
rect 46486 299483 46538 299489
rect 46102 298135 46154 298141
rect 46102 298077 46154 298083
rect 46870 298135 46922 298141
rect 46870 298077 46922 298083
rect 46198 297099 46250 297105
rect 46198 297041 46250 297047
rect 46102 293917 46154 293923
rect 46102 293859 46154 293865
rect 46114 281343 46142 293859
rect 46102 281337 46154 281343
rect 46102 281279 46154 281285
rect 46004 278194 46060 278203
rect 46004 278129 46060 278138
rect 46102 266389 46154 266395
rect 46102 266331 46154 266337
rect 46114 265063 46142 266331
rect 46102 265057 46154 265063
rect 46102 264999 46154 265005
rect 45910 213331 45962 213337
rect 45910 213273 45962 213279
rect 45718 212961 45770 212967
rect 45718 212903 45770 212909
rect 45622 212221 45674 212227
rect 45622 212163 45674 212169
rect 46114 209415 46142 264999
rect 46210 264989 46238 297041
rect 46882 296809 46910 298077
rect 46870 296803 46922 296809
rect 46870 296745 46922 296751
rect 46294 295915 46346 295921
rect 46294 295857 46346 295863
rect 46198 264983 46250 264989
rect 46198 264925 46250 264931
rect 46210 263657 46238 264925
rect 46198 263651 46250 263657
rect 46198 263593 46250 263599
rect 46306 263583 46334 295857
rect 46294 263577 46346 263583
rect 46292 263542 46294 263551
rect 46346 263542 46348 263551
rect 46292 263477 46348 263486
rect 46196 263394 46252 263403
rect 46196 263329 46252 263338
rect 46210 262177 46238 263329
rect 46198 262171 46250 262177
rect 46198 262113 46250 262119
rect 46210 210229 46238 262113
rect 47458 246489 47486 805125
rect 47554 785283 47582 817927
rect 57622 800669 57674 800675
rect 57622 800611 57674 800617
rect 57634 789691 57662 800611
rect 58004 789830 58060 789839
rect 58004 789765 58006 789774
rect 58058 789765 58060 789774
rect 58006 789733 58058 789739
rect 57620 789682 57676 789691
rect 57620 789617 57676 789626
rect 58198 789199 58250 789205
rect 58198 789141 58250 789147
rect 58210 788507 58238 789141
rect 58390 789125 58442 789131
rect 58390 789067 58442 789073
rect 58196 788498 58252 788507
rect 58196 788433 58252 788442
rect 58402 787323 58430 789067
rect 58388 787314 58444 787323
rect 58388 787249 58444 787258
rect 58678 785647 58730 785653
rect 58678 785589 58730 785595
rect 47542 785277 47594 785283
rect 47542 785219 47594 785225
rect 58690 784955 58718 785589
rect 59636 785390 59692 785399
rect 59636 785325 59692 785334
rect 59650 785283 59678 785325
rect 59638 785277 59690 785283
rect 59638 785219 59690 785225
rect 58676 784946 58732 784955
rect 58676 784881 58732 784890
rect 47638 774695 47690 774701
rect 47638 774637 47690 774643
rect 47542 762115 47594 762121
rect 47542 762057 47594 762063
rect 47554 254999 47582 762057
rect 47650 743029 47678 774637
rect 62038 772179 62090 772185
rect 62038 772121 62090 772127
rect 61846 771957 61898 771963
rect 61846 771899 61898 771905
rect 57910 748795 57962 748801
rect 57910 748737 57962 748743
rect 57922 747659 57950 748737
rect 57908 747650 57964 747659
rect 57908 747585 57964 747594
rect 54740 746022 54796 746031
rect 54646 745983 54698 745989
rect 54740 745957 54742 745966
rect 54646 745925 54698 745931
rect 54794 745957 54796 745966
rect 57622 745983 57674 745989
rect 54742 745925 54794 745931
rect 57622 745925 57674 745931
rect 54658 745883 54686 745925
rect 54644 745874 54700 745883
rect 54644 745809 54700 745818
rect 57634 745291 57662 745925
rect 59636 745430 59692 745439
rect 59254 745391 59306 745397
rect 59636 745365 59692 745374
rect 59254 745333 59306 745339
rect 57620 745282 57676 745291
rect 57620 745217 57676 745226
rect 59266 744107 59294 745333
rect 59650 745323 59678 745365
rect 59638 745317 59690 745323
rect 59638 745259 59690 745265
rect 59252 744098 59308 744107
rect 59252 744033 59308 744042
rect 47638 743023 47690 743029
rect 47638 742965 47690 742971
rect 59638 743023 59690 743029
rect 59638 742965 59690 742971
rect 59650 742923 59678 742965
rect 59734 742949 59786 742955
rect 59636 742914 59692 742923
rect 59734 742891 59786 742897
rect 59636 742849 59692 742858
rect 59746 741739 59774 742891
rect 59732 741730 59788 741739
rect 59732 741665 59788 741674
rect 50326 731479 50378 731485
rect 50326 731421 50378 731427
rect 47734 730739 47786 730745
rect 47734 730681 47786 730687
rect 47638 718751 47690 718757
rect 47638 718693 47690 718699
rect 47542 254993 47594 254999
rect 47542 254935 47594 254941
rect 47650 246637 47678 718693
rect 47746 699739 47774 730681
rect 50338 699813 50366 731421
rect 58390 704913 58442 704919
rect 58390 704855 58442 704861
rect 58402 704443 58430 704855
rect 58388 704434 58444 704443
rect 58388 704369 58444 704378
rect 58774 702693 58826 702699
rect 58772 702658 58774 702667
rect 58826 702658 58828 702667
rect 58678 702619 58730 702625
rect 58772 702593 58828 702602
rect 58678 702561 58730 702567
rect 58690 700891 58718 702561
rect 58676 700882 58732 700891
rect 58676 700817 58732 700826
rect 50326 699807 50378 699813
rect 50326 699749 50378 699755
rect 59254 699807 59306 699813
rect 59254 699749 59306 699755
rect 47734 699733 47786 699739
rect 47734 699675 47786 699681
rect 58870 699733 58922 699739
rect 59266 699707 59294 699749
rect 58870 699675 58922 699681
rect 59252 699698 59308 699707
rect 58882 698523 58910 699675
rect 59252 699633 59308 699642
rect 58868 698514 58924 698523
rect 58868 698449 58924 698458
rect 53206 688263 53258 688269
rect 53206 688205 53258 688211
rect 50326 687523 50378 687529
rect 50326 687465 50378 687471
rect 47830 687227 47882 687233
rect 47830 687169 47882 687175
rect 47734 675757 47786 675763
rect 47734 675699 47786 675705
rect 47638 246631 47690 246637
rect 47638 246573 47690 246579
rect 47746 246563 47774 675699
rect 47842 659483 47870 687169
rect 47830 659477 47882 659483
rect 47830 659419 47882 659425
rect 50338 656597 50366 687465
rect 53218 656671 53246 688205
rect 59638 671095 59690 671101
rect 59638 671037 59690 671043
rect 59650 661227 59678 671037
rect 59636 661218 59692 661227
rect 59636 661153 59692 661162
rect 59158 659477 59210 659483
rect 58772 659442 58828 659451
rect 59158 659419 59210 659425
rect 58772 659377 58774 659386
rect 58826 659377 58828 659386
rect 58774 659345 58826 659351
rect 59170 657675 59198 659419
rect 59156 657666 59212 657675
rect 59156 657601 59212 657610
rect 53206 656665 53258 656671
rect 53206 656607 53258 656613
rect 58198 656665 58250 656671
rect 58198 656607 58250 656613
rect 50326 656591 50378 656597
rect 50326 656533 50378 656539
rect 58210 656491 58238 656607
rect 58390 656591 58442 656597
rect 58390 656533 58442 656539
rect 58196 656482 58252 656491
rect 58196 656417 58252 656426
rect 58402 655307 58430 656533
rect 58388 655298 58444 655307
rect 58388 655233 58444 655242
rect 53206 644899 53258 644905
rect 53206 644841 53258 644847
rect 50326 644307 50378 644313
rect 50326 644249 50378 644255
rect 47926 644011 47978 644017
rect 47926 643953 47978 643959
rect 47830 632541 47882 632547
rect 47830 632483 47882 632489
rect 47734 246557 47786 246563
rect 47734 246499 47786 246505
rect 47446 246483 47498 246489
rect 47446 246425 47498 246431
rect 47842 246415 47870 632483
rect 47938 616341 47966 643953
rect 47926 616335 47978 616341
rect 47926 616277 47978 616283
rect 50338 613381 50366 644249
rect 53218 613455 53246 644841
rect 54646 627879 54698 627885
rect 54646 627821 54698 627827
rect 54658 624851 54686 627821
rect 54646 624845 54698 624851
rect 54646 624787 54698 624793
rect 58966 624845 59018 624851
rect 58966 624787 59018 624793
rect 58978 618011 59006 624787
rect 58964 618002 59020 618011
rect 58964 617937 59020 617946
rect 58198 616409 58250 616415
rect 58198 616351 58250 616357
rect 58210 615643 58238 616351
rect 58966 616335 59018 616341
rect 58966 616277 59018 616283
rect 58196 615634 58252 615643
rect 58196 615569 58252 615578
rect 58978 614459 59006 616277
rect 59638 616261 59690 616267
rect 59636 616226 59638 616235
rect 59690 616226 59692 616235
rect 59636 616161 59692 616170
rect 58964 614450 59020 614459
rect 58964 614385 59020 614394
rect 53206 613449 53258 613455
rect 53206 613391 53258 613397
rect 59638 613449 59690 613455
rect 59638 613391 59690 613397
rect 50326 613375 50378 613381
rect 50326 613317 50378 613323
rect 59542 613375 59594 613381
rect 59542 613317 59594 613323
rect 59554 612091 59582 613317
rect 59650 613275 59678 613391
rect 59636 613266 59692 613275
rect 59636 613201 59692 613210
rect 59540 612082 59596 612091
rect 59540 612017 59596 612026
rect 53206 601387 53258 601393
rect 53206 601329 53258 601335
rect 50326 600795 50378 600801
rect 50326 600737 50378 600743
rect 47926 579483 47978 579489
rect 47926 579425 47978 579431
rect 47938 573051 47966 579425
rect 50338 573125 50366 600737
rect 50326 573119 50378 573125
rect 50326 573061 50378 573067
rect 47926 573045 47978 573051
rect 47926 572987 47978 572993
rect 53218 570165 53246 601329
rect 56182 599093 56234 599099
rect 56182 599035 56234 599041
rect 56086 587549 56138 587555
rect 56086 587491 56138 587497
rect 53206 570159 53258 570165
rect 53206 570101 53258 570107
rect 50326 524353 50378 524359
rect 50326 524295 50378 524301
rect 47926 524279 47978 524285
rect 47926 524221 47978 524227
rect 47938 475593 47966 524221
rect 50338 476111 50366 524295
rect 50326 476105 50378 476111
rect 50326 476047 50378 476053
rect 47926 475587 47978 475593
rect 47926 475529 47978 475535
rect 47926 463599 47978 463605
rect 47926 463541 47978 463547
rect 47938 249153 47966 463541
rect 53206 429263 53258 429269
rect 53206 429205 53258 429211
rect 50326 428523 50378 428529
rect 50326 428465 50378 428471
rect 48118 428227 48170 428233
rect 48118 428169 48170 428175
rect 48022 416535 48074 416541
rect 48022 416477 48074 416483
rect 48034 255073 48062 416477
rect 48130 400187 48158 428169
rect 50338 400261 50366 428465
rect 53218 400335 53246 429205
rect 53206 400329 53258 400335
rect 53206 400271 53258 400277
rect 50326 400255 50378 400261
rect 50326 400197 50378 400203
rect 48118 400181 48170 400187
rect 48118 400123 48170 400129
rect 53206 386047 53258 386053
rect 53206 385989 53258 385995
rect 50326 385307 50378 385313
rect 50326 385249 50378 385255
rect 48214 385011 48266 385017
rect 48214 384953 48266 384959
rect 48118 373319 48170 373325
rect 48118 373261 48170 373267
rect 48022 255067 48074 255073
rect 48022 255009 48074 255015
rect 48130 254925 48158 373261
rect 48226 357045 48254 384953
rect 48214 357039 48266 357045
rect 48214 356981 48266 356987
rect 50338 356971 50366 385249
rect 53218 357119 53246 385989
rect 53206 357113 53258 357119
rect 53206 357055 53258 357061
rect 50326 356965 50378 356971
rect 50326 356907 50378 356913
rect 53206 342831 53258 342837
rect 53206 342773 53258 342779
rect 50326 342313 50378 342319
rect 50326 342255 50378 342261
rect 48214 341795 48266 341801
rect 48214 341737 48266 341743
rect 48226 313755 48254 341737
rect 50338 313829 50366 342255
rect 53218 313903 53246 342773
rect 53206 313897 53258 313903
rect 53206 313839 53258 313845
rect 50326 313823 50378 313829
rect 50326 313765 50378 313771
rect 48214 313749 48266 313755
rect 48214 313691 48266 313697
rect 54550 299541 54602 299547
rect 54550 299483 54602 299489
rect 52822 298579 52874 298585
rect 52822 298521 52874 298527
rect 48982 293843 49034 293849
rect 48982 293785 49034 293791
rect 48214 285259 48266 285265
rect 48214 285201 48266 285207
rect 48226 256405 48254 285201
rect 48994 279345 49022 293785
rect 52834 291333 52862 298521
rect 52822 291327 52874 291333
rect 52822 291269 52874 291275
rect 54562 291037 54590 299483
rect 54550 291031 54602 291037
rect 54550 290973 54602 290979
rect 53206 285185 53258 285191
rect 53206 285127 53258 285133
rect 48982 279339 49034 279345
rect 48982 279281 49034 279287
rect 50516 275382 50572 275391
rect 50516 275317 50572 275326
rect 50324 275234 50380 275243
rect 50324 275169 50380 275178
rect 48214 256399 48266 256405
rect 48214 256341 48266 256347
rect 48118 254919 48170 254925
rect 48118 254861 48170 254867
rect 47926 249147 47978 249153
rect 47926 249089 47978 249095
rect 47830 246409 47882 246415
rect 47830 246351 47882 246357
rect 46198 210223 46250 210229
rect 46198 210165 46250 210171
rect 50338 210007 50366 275169
rect 50530 210747 50558 275317
rect 53218 255443 53246 285127
rect 53206 255437 53258 255443
rect 53206 255379 53258 255385
rect 56098 252039 56126 587491
rect 56194 570239 56222 599035
rect 58966 584737 59018 584743
rect 58966 584679 59018 584685
rect 58978 574795 59006 584679
rect 58964 574786 59020 574795
rect 58964 574721 59020 574730
rect 58966 573119 59018 573125
rect 58966 573061 59018 573067
rect 58978 571243 59006 573061
rect 59638 573045 59690 573051
rect 59636 573010 59638 573019
rect 59690 573010 59692 573019
rect 59636 572945 59692 572954
rect 58964 571234 59020 571243
rect 58964 571169 59020 571178
rect 56182 570233 56234 570239
rect 56182 570175 56234 570181
rect 60406 570233 60458 570239
rect 60406 570175 60458 570181
rect 59158 570159 59210 570165
rect 59158 570101 59210 570107
rect 59170 568875 59198 570101
rect 60418 570059 60446 570175
rect 60404 570050 60460 570059
rect 60404 569985 60460 569994
rect 59156 568866 59212 568875
rect 59156 568801 59212 568810
rect 57718 541595 57770 541601
rect 57718 541537 57770 541543
rect 57622 541521 57674 541527
rect 57622 541463 57674 541469
rect 57634 530543 57662 541463
rect 57730 531727 57758 541537
rect 57716 531718 57772 531727
rect 57716 531653 57772 531662
rect 57620 530534 57676 530543
rect 57620 530469 57676 530478
rect 58964 527130 59020 527139
rect 58964 527065 59020 527074
rect 58580 525946 58636 525955
rect 58580 525881 58636 525890
rect 58594 524359 58622 525881
rect 58582 524353 58634 524359
rect 58582 524295 58634 524301
rect 58978 472411 59006 527065
rect 59348 524762 59404 524771
rect 59348 524697 59404 524706
rect 59362 524285 59390 524697
rect 59350 524279 59402 524285
rect 59350 524221 59402 524227
rect 58966 472405 59018 472411
rect 58966 472347 59018 472353
rect 58486 406101 58538 406107
rect 58486 406043 58538 406049
rect 58498 404151 58526 406043
rect 58484 404142 58540 404151
rect 58484 404077 58540 404086
rect 59638 402845 59690 402851
rect 59636 402810 59638 402819
rect 59690 402810 59692 402819
rect 59636 402745 59692 402754
rect 57620 400590 57676 400599
rect 57620 400525 57676 400534
rect 57634 394563 57662 400525
rect 59734 400329 59786 400335
rect 59734 400271 59786 400277
rect 59542 400255 59594 400261
rect 59542 400197 59594 400203
rect 59554 398231 59582 400197
rect 59638 400181 59690 400187
rect 59638 400123 59690 400129
rect 59650 400007 59678 400123
rect 59636 399998 59692 400007
rect 59636 399933 59692 399942
rect 59746 399415 59774 400271
rect 59732 399406 59788 399415
rect 59732 399341 59788 399350
rect 59540 398222 59596 398231
rect 59540 398157 59596 398166
rect 57622 394557 57674 394563
rect 57622 394499 57674 394505
rect 58294 362589 58346 362595
rect 58294 362531 58346 362537
rect 58306 360935 58334 362531
rect 58292 360926 58348 360935
rect 58292 360861 58348 360870
rect 59158 359999 59210 360005
rect 59158 359941 59210 359947
rect 59170 359751 59198 359941
rect 59156 359742 59212 359751
rect 59156 359677 59212 359686
rect 57620 357522 57676 357531
rect 57620 357457 57676 357466
rect 57634 351347 57662 357457
rect 58198 357113 58250 357119
rect 58198 357055 58250 357061
rect 58210 356199 58238 357055
rect 59638 357039 59690 357045
rect 59638 356981 59690 356987
rect 58582 356965 58634 356971
rect 58582 356907 58634 356913
rect 58196 356190 58252 356199
rect 58196 356125 58252 356134
rect 58594 355015 58622 356907
rect 59650 356791 59678 356981
rect 59636 356782 59692 356791
rect 59636 356717 59692 356726
rect 58580 355006 58636 355015
rect 58580 354941 58636 354950
rect 57622 351341 57674 351347
rect 57622 351283 57674 351289
rect 58486 319669 58538 319675
rect 58486 319611 58538 319617
rect 58498 317719 58526 319611
rect 58484 317710 58540 317719
rect 58484 317645 58540 317654
rect 59158 316783 59210 316789
rect 59158 316725 59210 316731
rect 59170 316535 59198 316725
rect 59156 316526 59212 316535
rect 59156 316461 59212 316470
rect 59060 314158 59116 314167
rect 59060 314093 59116 314102
rect 59074 308131 59102 314093
rect 59734 313897 59786 313903
rect 59734 313839 59786 313845
rect 59542 313823 59594 313829
rect 59542 313765 59594 313771
rect 59554 311799 59582 313765
rect 59638 313749 59690 313755
rect 59638 313691 59690 313697
rect 59650 313575 59678 313691
rect 59636 313566 59692 313575
rect 59636 313501 59692 313510
rect 59746 312983 59774 313839
rect 59732 312974 59788 312983
rect 59732 312909 59788 312918
rect 59540 311790 59596 311799
rect 59540 311725 59596 311734
rect 59062 308125 59114 308131
rect 59062 308067 59114 308073
rect 60214 299615 60266 299621
rect 60214 299557 60266 299563
rect 57526 296729 57578 296735
rect 57526 296671 57578 296677
rect 57538 290339 57566 296671
rect 59636 295214 59692 295223
rect 59636 295149 59692 295158
rect 58196 294030 58252 294039
rect 58196 293965 58252 293974
rect 58210 293849 58238 293965
rect 59650 293923 59678 295149
rect 59638 293917 59690 293923
rect 59638 293859 59690 293865
rect 58198 293843 58250 293849
rect 58198 293785 58250 293791
rect 59060 292846 59116 292855
rect 59060 292781 59116 292790
rect 59074 290963 59102 292781
rect 59636 291662 59692 291671
rect 59636 291597 59692 291606
rect 59650 291333 59678 291597
rect 60226 291523 60254 299557
rect 60212 291514 60268 291523
rect 60212 291449 60268 291458
rect 59638 291327 59690 291333
rect 59638 291269 59690 291275
rect 59062 290957 59114 290963
rect 59062 290899 59114 290905
rect 57524 290330 57580 290339
rect 57524 290265 57580 290274
rect 59636 288110 59692 288119
rect 59636 288045 59638 288054
rect 59690 288045 59692 288054
rect 59638 288013 59690 288019
rect 58100 286926 58156 286935
rect 58100 286861 58156 286870
rect 58114 285191 58142 286861
rect 59540 285742 59596 285751
rect 59540 285677 59596 285686
rect 59554 285265 59582 285677
rect 59542 285259 59594 285265
rect 59542 285201 59594 285207
rect 58102 285185 58154 285191
rect 58102 285127 58154 285133
rect 57620 284558 57676 284567
rect 57620 284493 57676 284502
rect 57634 282305 57662 284493
rect 59636 283374 59692 283383
rect 59636 283309 59692 283318
rect 59650 282601 59678 283309
rect 59638 282595 59690 282601
rect 59638 282537 59690 282543
rect 58964 282486 59020 282495
rect 58964 282421 59020 282430
rect 58978 282379 59006 282421
rect 58966 282373 59018 282379
rect 58966 282315 59018 282321
rect 56182 282299 56234 282305
rect 56182 282241 56234 282247
rect 57622 282299 57674 282305
rect 57622 282241 57674 282247
rect 56194 253519 56222 282241
rect 58196 281006 58252 281015
rect 58196 280941 58252 280950
rect 58210 279419 58238 280941
rect 59636 279822 59692 279831
rect 59636 279757 59692 279766
rect 59650 279493 59678 279757
rect 59638 279487 59690 279493
rect 59638 279429 59690 279435
rect 58198 279413 58250 279419
rect 58198 279355 58250 279361
rect 61858 266955 61886 771899
rect 61942 642531 61994 642537
rect 61942 642473 61994 642479
rect 61954 276131 61982 642473
rect 61940 276122 61996 276131
rect 61940 276057 61996 276066
rect 61844 266946 61900 266955
rect 61844 266881 61900 266890
rect 62050 266807 62078 772121
rect 62230 728889 62282 728895
rect 62230 728831 62282 728837
rect 62134 599241 62186 599247
rect 62134 599183 62186 599189
rect 62146 278055 62174 599183
rect 62242 286745 62270 728831
rect 62422 728815 62474 728821
rect 62422 728757 62474 728763
rect 62326 600499 62378 600505
rect 62326 600441 62378 600447
rect 62230 286739 62282 286745
rect 62230 286681 62282 286687
rect 62132 278046 62188 278055
rect 62132 277981 62188 277990
rect 62338 277759 62366 600441
rect 62324 277750 62380 277759
rect 62324 277685 62380 277694
rect 62434 277588 62462 728757
rect 62518 432075 62570 432081
rect 62518 432017 62570 432023
rect 62242 277560 62462 277588
rect 62036 266798 62092 266807
rect 62036 266733 62092 266742
rect 62242 266659 62270 277560
rect 62530 271543 62558 432017
rect 62710 300947 62762 300953
rect 62710 300889 62762 300895
rect 62722 277611 62750 300889
rect 62806 298135 62858 298141
rect 62806 298077 62858 298083
rect 62708 277602 62764 277611
rect 62708 277537 62764 277546
rect 62818 277463 62846 298077
rect 63286 290883 63338 290889
rect 63286 290825 63338 290831
rect 62902 286739 62954 286745
rect 62902 286681 62954 286687
rect 62804 277454 62860 277463
rect 62804 277389 62860 277398
rect 62516 271534 62572 271543
rect 62516 271469 62572 271478
rect 62228 266650 62284 266659
rect 62228 266585 62284 266594
rect 62914 266511 62942 286681
rect 63298 282176 63326 290825
rect 63298 282148 63422 282176
rect 63394 277939 63422 282148
rect 313558 278377 313610 278383
rect 313558 278319 313610 278325
rect 404758 278377 404810 278383
rect 404810 278325 405072 278328
rect 404758 278319 405072 278325
rect 63382 277933 63434 277939
rect 63382 277875 63434 277881
rect 65890 269323 65918 278018
rect 65876 269314 65932 269323
rect 67042 269281 67070 278018
rect 68290 273277 68318 278018
rect 68278 273271 68330 273277
rect 68278 273213 68330 273219
rect 69442 269619 69470 278018
rect 70594 272135 70622 278018
rect 70580 272126 70636 272135
rect 70580 272061 70636 272070
rect 69428 269610 69484 269619
rect 69428 269545 69484 269554
rect 71746 269471 71774 278018
rect 72994 272283 73022 278018
rect 72980 272274 73036 272283
rect 72980 272209 73036 272218
rect 71732 269462 71788 269471
rect 71732 269397 71788 269406
rect 74146 269355 74174 278018
rect 75298 271649 75326 278018
rect 76546 272167 76574 278018
rect 77698 276494 77726 278018
rect 77602 276466 77726 276494
rect 76534 272161 76586 272167
rect 76534 272103 76586 272109
rect 75286 271643 75338 271649
rect 75286 271585 75338 271591
rect 77602 269767 77630 276466
rect 78850 272431 78878 278018
rect 80112 278004 80606 278032
rect 78836 272422 78892 272431
rect 78836 272357 78892 272366
rect 77686 271643 77738 271649
rect 77686 271585 77738 271591
rect 77588 269758 77644 269767
rect 77588 269693 77644 269702
rect 74134 269349 74186 269355
rect 74134 269291 74186 269297
rect 65876 269249 65932 269258
rect 67030 269275 67082 269281
rect 67030 269217 67082 269223
rect 62900 266502 62956 266511
rect 62900 266437 62956 266446
rect 56182 253513 56234 253519
rect 56182 253455 56234 253461
rect 56086 252033 56138 252039
rect 56086 251975 56138 251981
rect 77698 249375 77726 271585
rect 77686 249369 77738 249375
rect 77686 249311 77738 249317
rect 80578 249227 80606 278004
rect 81250 269503 81278 278018
rect 81238 269497 81290 269503
rect 81238 269439 81290 269445
rect 82402 269429 82430 278018
rect 83650 269651 83678 278018
rect 84802 272241 84830 278018
rect 84790 272235 84842 272241
rect 84790 272177 84842 272183
rect 85954 271131 85982 278018
rect 86326 272235 86378 272241
rect 86326 272177 86378 272183
rect 85942 271125 85994 271131
rect 85942 271067 85994 271073
rect 83638 269645 83690 269651
rect 83638 269587 83690 269593
rect 82390 269423 82442 269429
rect 82390 269365 82442 269371
rect 86338 249301 86366 272177
rect 87202 269577 87230 278018
rect 88354 272579 88382 278018
rect 88340 272570 88396 272579
rect 88340 272505 88396 272514
rect 89506 271575 89534 278018
rect 89494 271569 89546 271575
rect 89494 271511 89546 271517
rect 90658 269725 90686 278018
rect 91906 272727 91934 278018
rect 91892 272718 91948 272727
rect 91892 272653 91948 272662
rect 92086 271569 92138 271575
rect 92086 271511 92138 271517
rect 90646 269719 90698 269725
rect 90646 269661 90698 269667
rect 87190 269571 87242 269577
rect 87190 269513 87242 269519
rect 92098 249449 92126 271511
rect 93058 269799 93086 278018
rect 94210 270761 94238 278018
rect 94198 270755 94250 270761
rect 94198 270697 94250 270703
rect 94966 270755 95018 270761
rect 94966 270697 95018 270703
rect 93046 269793 93098 269799
rect 93046 269735 93098 269741
rect 94978 252335 95006 270697
rect 95458 269873 95486 278018
rect 96610 272315 96638 278018
rect 97776 278004 97886 278032
rect 96598 272309 96650 272315
rect 96598 272251 96650 272257
rect 95446 269867 95498 269873
rect 95446 269809 95498 269815
rect 97858 252409 97886 278004
rect 99010 272389 99038 278018
rect 98998 272383 99050 272389
rect 98998 272325 99050 272331
rect 100162 269947 100190 278018
rect 101314 271797 101342 278018
rect 101302 271791 101354 271797
rect 101302 271733 101354 271739
rect 102562 270095 102590 278018
rect 103714 272463 103742 278018
rect 103702 272457 103754 272463
rect 103702 272399 103754 272405
rect 104866 272241 104894 278018
rect 106114 272537 106142 278018
rect 106102 272531 106154 272537
rect 106102 272473 106154 272479
rect 104854 272235 104906 272241
rect 104854 272177 104906 272183
rect 106486 272235 106538 272241
rect 106486 272177 106538 272183
rect 103606 271791 103658 271797
rect 103606 271733 103658 271739
rect 102550 270089 102602 270095
rect 102550 270031 102602 270037
rect 100150 269941 100202 269947
rect 100150 269883 100202 269889
rect 97846 252403 97898 252409
rect 97846 252345 97898 252351
rect 94966 252329 95018 252335
rect 94966 252271 95018 252277
rect 103618 252261 103646 271733
rect 103606 252255 103658 252261
rect 103606 252197 103658 252203
rect 106498 252187 106526 272177
rect 107266 270021 107294 278018
rect 108418 273499 108446 278018
rect 108406 273493 108458 273499
rect 108406 273435 108458 273441
rect 109366 273493 109418 273499
rect 109366 273435 109418 273441
rect 107254 270015 107306 270021
rect 107254 269957 107306 269963
rect 106486 252181 106538 252187
rect 106486 252123 106538 252129
rect 109378 252113 109406 273435
rect 109570 270169 109598 278018
rect 110818 272611 110846 278018
rect 111984 278004 112286 278032
rect 110806 272605 110858 272611
rect 110806 272547 110858 272553
rect 109558 270163 109610 270169
rect 109558 270105 109610 270111
rect 109366 252107 109418 252113
rect 109366 252049 109418 252055
rect 92086 249443 92138 249449
rect 92086 249385 92138 249391
rect 86326 249295 86378 249301
rect 86326 249237 86378 249243
rect 80566 249221 80618 249227
rect 80566 249163 80618 249169
rect 112258 246711 112286 278004
rect 113122 272685 113150 278018
rect 113110 272679 113162 272685
rect 113110 272621 113162 272627
rect 114370 270243 114398 278018
rect 115522 270761 115550 278018
rect 116674 272833 116702 278018
rect 116662 272827 116714 272833
rect 116662 272769 116714 272775
rect 115510 270755 115562 270761
rect 115510 270697 115562 270703
rect 117922 270317 117950 278018
rect 119074 270761 119102 278018
rect 120226 272759 120254 278018
rect 120214 272753 120266 272759
rect 120214 272695 120266 272701
rect 118006 270755 118058 270761
rect 118006 270697 118058 270703
rect 119062 270755 119114 270761
rect 119062 270697 119114 270703
rect 120886 270755 120938 270761
rect 120886 270697 120938 270703
rect 117910 270311 117962 270317
rect 117910 270253 117962 270259
rect 114358 270237 114410 270243
rect 114358 270179 114410 270185
rect 118018 249819 118046 270697
rect 118006 249813 118058 249819
rect 118006 249755 118058 249761
rect 120898 249597 120926 270697
rect 121474 270391 121502 278018
rect 122626 273425 122654 278018
rect 123778 276494 123806 278018
rect 123682 276466 123806 276494
rect 122614 273419 122666 273425
rect 122614 273361 122666 273367
rect 123682 272907 123710 276466
rect 123766 273419 123818 273425
rect 123766 273361 123818 273367
rect 123670 272901 123722 272907
rect 123670 272843 123722 272849
rect 121462 270385 121514 270391
rect 121462 270327 121514 270333
rect 123778 249745 123806 273361
rect 125026 273055 125054 278018
rect 126192 278004 126686 278032
rect 125014 273049 125066 273055
rect 125014 272991 125066 272997
rect 123766 249739 123818 249745
rect 123766 249681 123818 249687
rect 126658 249671 126686 278004
rect 127330 273129 127358 278018
rect 127318 273123 127370 273129
rect 127318 273065 127370 273071
rect 128482 272981 128510 278018
rect 128470 272975 128522 272981
rect 128470 272917 128522 272923
rect 129730 271649 129758 278018
rect 130882 273499 130910 278018
rect 130870 273493 130922 273499
rect 130870 273435 130922 273441
rect 132034 273203 132062 278018
rect 132022 273197 132074 273203
rect 132022 273139 132074 273145
rect 129718 271643 129770 271649
rect 129718 271585 129770 271591
rect 132406 271643 132458 271649
rect 132406 271585 132458 271591
rect 126646 249665 126698 249671
rect 126646 249607 126698 249613
rect 120886 249591 120938 249597
rect 120886 249533 120938 249539
rect 132418 249523 132446 271585
rect 133282 270761 133310 278018
rect 133270 270755 133322 270761
rect 133270 270697 133322 270703
rect 134434 270465 134462 278018
rect 135586 273351 135614 278018
rect 135574 273345 135626 273351
rect 135574 273287 135626 273293
rect 136834 270761 136862 278018
rect 135286 270755 135338 270761
rect 135286 270697 135338 270703
rect 136822 270755 136874 270761
rect 136822 270697 136874 270703
rect 134422 270459 134474 270465
rect 134422 270401 134474 270407
rect 135298 249967 135326 270697
rect 137986 270613 138014 278018
rect 138166 270755 138218 270761
rect 138166 270697 138218 270703
rect 137974 270607 138026 270613
rect 137974 270549 138026 270555
rect 135286 249961 135338 249967
rect 135286 249903 135338 249909
rect 138178 249893 138206 270697
rect 139138 269915 139166 278018
rect 140400 278004 141086 278032
rect 139124 269906 139180 269915
rect 139124 269841 139180 269850
rect 141058 252483 141086 278004
rect 141538 270539 141566 278018
rect 142690 273425 142718 278018
rect 142678 273419 142730 273425
rect 142678 273361 142730 273367
rect 142486 273271 142538 273277
rect 142486 273213 142538 273219
rect 141526 270533 141578 270539
rect 141526 270475 141578 270481
rect 141046 252477 141098 252483
rect 141046 252419 141098 252425
rect 138166 249887 138218 249893
rect 138166 249829 138218 249835
rect 132406 249517 132458 249523
rect 132406 249459 132458 249465
rect 112246 246705 112298 246711
rect 112246 246647 112298 246653
rect 142498 216014 142526 273213
rect 142582 242635 142634 242641
rect 142582 242577 142634 242583
rect 142594 236174 142622 242577
rect 142594 236146 143102 236174
rect 143074 218887 143102 236146
rect 143062 218881 143114 218887
rect 143062 218823 143114 218829
rect 142498 215986 143102 216014
rect 50518 210741 50570 210747
rect 50518 210683 50570 210689
rect 50326 210001 50378 210007
rect 50326 209943 50378 209949
rect 46102 209409 46154 209415
rect 46102 209351 46154 209357
rect 143074 201571 143102 215986
rect 143062 201565 143114 201571
rect 143062 201507 143114 201513
rect 143938 190101 143966 278018
rect 145090 269207 145118 278018
rect 146242 270687 146270 278018
rect 147394 271797 147422 278018
rect 147382 271791 147434 271797
rect 147382 271733 147434 271739
rect 146230 270681 146282 270687
rect 146230 270623 146282 270629
rect 145078 269201 145130 269207
rect 145078 269143 145130 269149
rect 148642 268985 148670 278018
rect 149686 271791 149738 271797
rect 149686 271733 149738 271739
rect 148630 268979 148682 268985
rect 148630 268921 148682 268927
rect 145558 249961 145610 249967
rect 145558 249903 145610 249909
rect 145366 249369 145418 249375
rect 145366 249311 145418 249317
rect 143926 190095 143978 190101
rect 143926 190037 143978 190043
rect 42166 182399 42218 182405
rect 42166 182341 42218 182347
rect 45334 182399 45386 182405
rect 45334 182341 45386 182347
rect 42178 182114 42206 182341
rect 145378 175597 145406 249311
rect 145462 245003 145514 245009
rect 145462 244945 145514 244951
rect 145474 175671 145502 244945
rect 145570 187215 145598 249903
rect 145654 244855 145706 244861
rect 145654 244797 145706 244803
rect 145666 221773 145694 244797
rect 148340 244598 148396 244607
rect 148340 244533 148396 244542
rect 148244 239714 148300 239723
rect 148244 239649 148300 239658
rect 146996 236014 147052 236023
rect 146996 235949 146998 235958
rect 147050 235949 147052 235958
rect 146998 235917 147050 235923
rect 147476 231130 147532 231139
rect 147476 231065 147532 231074
rect 147490 230505 147518 231065
rect 147478 230499 147530 230505
rect 147478 230441 147530 230447
rect 147092 229946 147148 229955
rect 147092 229881 147148 229890
rect 147106 229839 147134 229881
rect 147094 229833 147146 229839
rect 147094 229775 147146 229781
rect 147092 226394 147148 226403
rect 147092 226329 147148 226338
rect 147106 226287 147134 226329
rect 147094 226281 147146 226287
rect 147094 226223 147146 226229
rect 145654 221767 145706 221773
rect 145654 221709 145706 221715
rect 147284 217810 147340 217819
rect 147284 217745 147286 217754
rect 147338 217745 147340 217754
rect 147286 217713 147338 217719
rect 146900 212926 146956 212935
rect 146900 212861 146956 212870
rect 146914 212819 146942 212861
rect 146902 212813 146954 212819
rect 146902 212755 146954 212761
rect 147092 211742 147148 211751
rect 147092 211677 147148 211686
rect 147106 211043 147134 211677
rect 147094 211037 147146 211043
rect 147094 210979 147146 210985
rect 147476 210410 147532 210419
rect 147476 210345 147478 210354
rect 147530 210345 147532 210354
rect 147478 210313 147530 210319
rect 146900 209226 146956 209235
rect 146900 209161 146956 209170
rect 146914 207417 146942 209161
rect 147188 208042 147244 208051
rect 147188 207977 147244 207986
rect 147202 207935 147230 207977
rect 147190 207929 147242 207935
rect 147190 207871 147242 207877
rect 146902 207411 146954 207417
rect 146902 207353 146954 207359
rect 146900 206414 146956 206423
rect 146900 206349 146956 206358
rect 146914 206307 146942 206349
rect 146902 206301 146954 206307
rect 146902 206243 146954 206249
rect 147860 203306 147916 203315
rect 147860 203241 147916 203250
rect 147874 202903 147902 203241
rect 147862 202897 147914 202903
rect 147862 202839 147914 202845
rect 147572 199606 147628 199615
rect 147572 199541 147628 199550
rect 147586 199351 147614 199541
rect 147574 199345 147626 199351
rect 147574 199287 147626 199293
rect 147286 196015 147338 196021
rect 147286 195957 147338 195963
rect 147298 195915 147326 195957
rect 147284 195906 147340 195915
rect 147284 195841 147340 195850
rect 147668 189838 147724 189847
rect 147668 189773 147724 189782
rect 147682 189583 147710 189773
rect 147670 189577 147722 189583
rect 147670 189519 147722 189525
rect 145558 187209 145610 187215
rect 145558 187151 145610 187157
rect 145462 175665 145514 175671
rect 145462 175607 145514 175613
rect 145366 175591 145418 175597
rect 145366 175533 145418 175539
rect 147764 175186 147820 175195
rect 147764 175121 147820 175130
rect 147778 174413 147806 175121
rect 147766 174407 147818 174413
rect 147766 174349 147818 174355
rect 148258 169751 148286 239649
rect 148354 172711 148382 244533
rect 148724 243414 148780 243423
rect 148724 243349 148780 243358
rect 148532 242082 148588 242091
rect 148532 242017 148588 242026
rect 148436 238530 148492 238539
rect 148436 238465 148492 238474
rect 148342 172705 148394 172711
rect 148342 172647 148394 172653
rect 148450 169899 148478 238465
rect 148546 172563 148574 242017
rect 148628 236754 148684 236763
rect 148628 236689 148684 236698
rect 148534 172557 148586 172563
rect 148534 172499 148586 172505
rect 148438 169893 148490 169899
rect 148438 169835 148490 169841
rect 148642 169825 148670 236689
rect 148738 172785 148766 243349
rect 148916 240898 148972 240907
rect 148916 240833 148972 240842
rect 148820 234830 148876 234839
rect 148820 234765 148876 234774
rect 148726 172779 148778 172785
rect 148726 172721 148778 172727
rect 148630 169819 148682 169825
rect 148630 169761 148682 169767
rect 148246 169745 148298 169751
rect 148246 169687 148298 169693
rect 148724 169118 148780 169127
rect 148724 169053 148780 169062
rect 148532 168082 148588 168091
rect 148532 168017 148588 168026
rect 148436 165566 148492 165575
rect 148436 165501 148492 165510
rect 148244 164382 148300 164391
rect 148244 164317 148300 164326
rect 147092 159498 147148 159507
rect 147092 159433 147148 159442
rect 147106 158503 147134 159433
rect 147094 158497 147146 158503
rect 147094 158439 147146 158445
rect 147092 156982 147148 156991
rect 147092 156917 147148 156926
rect 147106 156209 147134 156917
rect 147094 156203 147146 156209
rect 147094 156145 147146 156151
rect 147092 141294 147148 141303
rect 147092 141229 147094 141238
rect 147146 141229 147148 141238
rect 147094 141197 147146 141203
rect 146902 141107 146954 141113
rect 146902 141049 146954 141055
rect 146914 139971 146942 141049
rect 146900 139962 146956 139971
rect 146900 139897 146956 139906
rect 148258 123871 148286 164317
rect 148340 161866 148396 161875
rect 148340 161801 148396 161810
rect 148246 123865 148298 123871
rect 148246 123807 148298 123813
rect 148354 120985 148382 161801
rect 148450 124408 148478 165501
rect 148546 126683 148574 168017
rect 148628 166306 148684 166315
rect 148628 166241 148684 166250
rect 148534 126677 148586 126683
rect 148534 126619 148586 126625
rect 148450 124380 148574 124408
rect 148436 124274 148492 124283
rect 148436 124209 148492 124218
rect 148450 123945 148478 124209
rect 148438 123939 148490 123945
rect 148438 123881 148490 123887
rect 148546 123797 148574 124380
rect 148534 123791 148586 123797
rect 148534 123733 148586 123739
rect 148642 123723 148670 166241
rect 148738 126609 148766 169053
rect 148834 166939 148862 234765
rect 148930 172637 148958 240833
rect 149012 233646 149068 233655
rect 149012 233581 149068 233590
rect 148918 172631 148970 172637
rect 148918 172573 148970 172579
rect 149026 167013 149054 233581
rect 149108 232314 149164 232323
rect 149108 232249 149164 232258
rect 149122 174136 149150 232249
rect 149396 228170 149452 228179
rect 149396 228105 149452 228114
rect 149410 227619 149438 228105
rect 149398 227613 149450 227619
rect 149398 227555 149450 227561
rect 149492 227430 149548 227439
rect 149492 227365 149548 227374
rect 149396 225210 149452 225219
rect 149396 225145 149452 225154
rect 149410 224807 149438 225145
rect 149506 224881 149534 227365
rect 149494 224875 149546 224881
rect 149494 224817 149546 224823
rect 149398 224801 149450 224807
rect 149398 224743 149450 224749
rect 149492 223878 149548 223887
rect 149492 223813 149548 223822
rect 149396 222694 149452 222703
rect 149396 222629 149452 222638
rect 149410 221921 149438 222629
rect 149398 221915 149450 221921
rect 149398 221857 149450 221863
rect 149506 221847 149534 223813
rect 149494 221841 149546 221847
rect 149494 221783 149546 221789
rect 149492 221510 149548 221519
rect 149492 221445 149548 221454
rect 149396 219734 149452 219743
rect 149396 219669 149452 219678
rect 149410 219109 149438 219669
rect 149398 219103 149450 219109
rect 149398 219045 149450 219051
rect 149506 219035 149534 221445
rect 149494 219029 149546 219035
rect 149396 218994 149452 219003
rect 149494 218971 149546 218977
rect 149396 218929 149398 218938
rect 149450 218929 149452 218938
rect 149398 218897 149450 218903
rect 149396 216626 149452 216635
rect 149396 216561 149452 216570
rect 149410 216075 149438 216561
rect 149398 216069 149450 216075
rect 149398 216011 149450 216017
rect 149492 214850 149548 214859
rect 149492 214785 149548 214794
rect 149396 214110 149452 214119
rect 149396 214045 149452 214054
rect 149410 213189 149438 214045
rect 149506 213263 149534 214785
rect 149494 213257 149546 213263
rect 149494 213199 149546 213205
rect 149398 213183 149450 213189
rect 149398 213125 149450 213131
rect 149492 205674 149548 205683
rect 149492 205609 149548 205618
rect 149506 204531 149534 205609
rect 149494 204525 149546 204531
rect 149396 204490 149452 204499
rect 149494 204467 149546 204473
rect 149396 204425 149452 204434
rect 149410 204235 149438 204425
rect 149398 204229 149450 204235
rect 149398 204171 149450 204177
rect 149396 201678 149452 201687
rect 149396 201613 149398 201622
rect 149450 201613 149452 201622
rect 149398 201581 149450 201587
rect 149396 200790 149452 200799
rect 149396 200725 149452 200734
rect 149410 200535 149438 200725
rect 149398 200529 149450 200535
rect 149398 200471 149450 200477
rect 149300 198422 149356 198431
rect 149300 198357 149356 198366
rect 149314 195873 149342 198357
rect 149396 197090 149452 197099
rect 149396 197025 149452 197034
rect 149410 195947 149438 197025
rect 149398 195941 149450 195947
rect 149398 195883 149450 195889
rect 149302 195867 149354 195873
rect 149302 195809 149354 195815
rect 149492 194722 149548 194731
rect 149492 194657 149548 194666
rect 149396 193242 149452 193251
rect 149396 193177 149452 193186
rect 149410 193135 149438 193177
rect 149398 193129 149450 193135
rect 149398 193071 149450 193077
rect 149506 193061 149534 194657
rect 149494 193055 149546 193061
rect 149494 192997 149546 193003
rect 149492 192206 149548 192215
rect 149492 192141 149548 192150
rect 149396 191022 149452 191031
rect 149396 190957 149452 190966
rect 149410 190249 149438 190957
rect 149398 190243 149450 190249
rect 149398 190185 149450 190191
rect 149506 190175 149534 192141
rect 149494 190169 149546 190175
rect 149494 190111 149546 190117
rect 149698 190027 149726 271733
rect 149794 269059 149822 278018
rect 150946 271575 150974 278018
rect 150934 271569 150986 271575
rect 150934 271511 150986 271517
rect 152194 269133 152222 278018
rect 153346 273277 153374 278018
rect 153334 273271 153386 273277
rect 153334 273213 153386 273219
rect 152374 271569 152426 271575
rect 152374 271511 152426 271517
rect 152182 269127 152234 269133
rect 152182 269069 152234 269075
rect 149782 269053 149834 269059
rect 149782 268995 149834 269001
rect 151222 235975 151274 235981
rect 151222 235917 151274 235923
rect 151126 226133 151178 226139
rect 151126 226075 151178 226081
rect 149686 190021 149738 190027
rect 149686 189963 149738 189969
rect 149300 188062 149356 188071
rect 149300 187997 149356 188006
rect 149204 184510 149260 184519
rect 149204 184445 149260 184454
rect 149218 174265 149246 184445
rect 149314 182923 149342 187997
rect 149396 187470 149452 187479
rect 149396 187405 149452 187414
rect 149410 182997 149438 187405
rect 149588 186286 149644 186295
rect 149588 186221 149644 186230
rect 149492 183770 149548 183779
rect 149492 183705 149548 183714
rect 149398 182991 149450 182997
rect 149398 182933 149450 182939
rect 149302 182917 149354 182923
rect 149302 182859 149354 182865
rect 149396 182586 149452 182595
rect 149396 182521 149452 182530
rect 149410 181517 149438 182521
rect 149506 181591 149534 183705
rect 149494 181585 149546 181591
rect 149494 181527 149546 181533
rect 149398 181511 149450 181517
rect 149398 181453 149450 181459
rect 149492 181402 149548 181411
rect 149492 181337 149548 181346
rect 149300 179626 149356 179635
rect 149300 179561 149356 179570
rect 149314 178631 149342 179561
rect 149396 178886 149452 178895
rect 149396 178821 149452 178830
rect 149410 178705 149438 178821
rect 149506 178779 149534 181337
rect 149602 180037 149630 186221
rect 149590 180031 149642 180037
rect 149590 179973 149642 179979
rect 149494 178773 149546 178779
rect 149494 178715 149546 178721
rect 149398 178699 149450 178705
rect 149398 178641 149450 178647
rect 149302 178625 149354 178631
rect 149302 178567 149354 178573
rect 149492 177702 149548 177711
rect 149492 177637 149548 177646
rect 149396 176518 149452 176527
rect 149396 176453 149452 176462
rect 149410 175819 149438 176453
rect 149398 175813 149450 175819
rect 149398 175755 149450 175761
rect 149506 175745 149534 177637
rect 149494 175739 149546 175745
rect 149494 175681 149546 175687
rect 149206 174259 149258 174265
rect 149206 174201 149258 174207
rect 149122 174108 149438 174136
rect 149108 174002 149164 174011
rect 149108 173937 149164 173946
rect 149014 167007 149066 167013
rect 149014 166949 149066 166955
rect 148822 166933 148874 166939
rect 148822 166875 148874 166881
rect 148916 163198 148972 163207
rect 148916 163133 148972 163142
rect 148820 160682 148876 160691
rect 148820 160617 148876 160626
rect 148834 134009 148862 160617
rect 148822 134003 148874 134009
rect 148822 133945 148874 133951
rect 148820 133894 148876 133903
rect 148820 133829 148876 133838
rect 148726 126603 148778 126609
rect 148726 126545 148778 126551
rect 148630 123717 148682 123723
rect 148630 123659 148682 123665
rect 148532 122498 148588 122507
rect 148532 122433 148588 122442
rect 148342 120979 148394 120985
rect 148342 120921 148394 120927
rect 148340 110954 148396 110963
rect 148340 110889 148396 110898
rect 147860 108438 147916 108447
rect 147860 108373 147862 108382
rect 147914 108373 147916 108382
rect 147862 108341 147914 108347
rect 147188 107254 147244 107263
rect 147188 107189 147190 107198
rect 147242 107189 147244 107198
rect 147190 107157 147242 107163
rect 148244 104738 148300 104747
rect 148244 104673 148300 104682
rect 148258 86353 148286 104673
rect 148354 92125 148382 110889
rect 148436 103554 148492 103563
rect 148436 103489 148492 103498
rect 148342 92119 148394 92125
rect 148342 92061 148394 92067
rect 148450 86427 148478 103489
rect 148546 97897 148574 122433
rect 148724 121758 148780 121767
rect 148724 121693 148780 121702
rect 148738 115214 148766 121693
rect 148834 115255 148862 133829
rect 148930 132973 148958 163133
rect 149014 147915 149066 147921
rect 149014 147857 149066 147863
rect 148918 132967 148970 132973
rect 148918 132909 148970 132915
rect 149026 132844 149054 147857
rect 149122 147792 149150 173937
rect 149300 171042 149356 171051
rect 149300 170977 149356 170986
rect 149204 170302 149260 170311
rect 149204 170237 149260 170246
rect 149218 147921 149246 170237
rect 149314 155636 149342 170977
rect 149410 166865 149438 174108
rect 149588 172818 149644 172827
rect 149588 172753 149644 172762
rect 149398 166859 149450 166865
rect 149398 166801 149450 166807
rect 149396 158018 149452 158027
rect 149396 157953 149452 157962
rect 149410 157689 149438 157953
rect 149398 157683 149450 157689
rect 149398 157625 149450 157631
rect 149396 155798 149452 155807
rect 149396 155733 149398 155742
rect 149450 155733 149452 155742
rect 149398 155701 149450 155707
rect 149314 155608 149438 155636
rect 149410 155534 149438 155608
rect 149314 155506 149438 155534
rect 149314 147940 149342 155506
rect 149492 154614 149548 154623
rect 149492 154549 149548 154558
rect 149396 152986 149452 152995
rect 149396 152921 149452 152930
rect 149410 152731 149438 152921
rect 149506 152805 149534 154549
rect 149494 152799 149546 152805
rect 149494 152741 149546 152747
rect 149398 152725 149450 152731
rect 149398 152667 149450 152673
rect 149492 150914 149548 150923
rect 149492 150849 149548 150858
rect 149398 149987 149450 149993
rect 149398 149929 149450 149935
rect 149410 149887 149438 149929
rect 149506 149919 149534 150849
rect 149494 149913 149546 149919
rect 149396 149878 149452 149887
rect 149494 149855 149546 149861
rect 149396 149813 149452 149822
rect 149492 148546 149548 148555
rect 149492 148481 149548 148490
rect 149206 147915 149258 147921
rect 149314 147912 149438 147940
rect 149206 147857 149258 147863
rect 149122 147764 149342 147792
rect 149206 147471 149258 147477
rect 149206 147413 149258 147419
rect 148930 132816 149054 132844
rect 148930 126535 148958 132816
rect 149012 132710 149068 132719
rect 149012 132645 149068 132654
rect 148918 126529 148970 126535
rect 148918 126471 148970 126477
rect 148642 115186 148766 115214
rect 148820 115246 148876 115255
rect 148534 97891 148586 97897
rect 148534 97833 148586 97839
rect 148642 97823 148670 115186
rect 148820 115181 148876 115190
rect 148724 111990 148780 111999
rect 148724 111925 148780 111934
rect 148630 97817 148682 97823
rect 148630 97759 148682 97765
rect 148738 92051 148766 111925
rect 148820 106070 148876 106079
rect 148820 106005 148876 106014
rect 148726 92045 148778 92051
rect 148726 91987 148778 91993
rect 148834 89239 148862 106005
rect 149026 103595 149054 132645
rect 149218 131216 149246 147413
rect 149122 131188 149246 131216
rect 149122 129421 149150 131188
rect 149314 131068 149342 147764
rect 149410 147477 149438 147912
rect 149398 147471 149450 147477
rect 149398 147413 149450 147419
rect 149396 147362 149452 147371
rect 149396 147297 149452 147306
rect 149410 147033 149438 147297
rect 149398 147027 149450 147033
rect 149398 146969 149450 146975
rect 149506 146959 149534 148481
rect 149494 146953 149546 146959
rect 149494 146895 149546 146901
rect 149492 146178 149548 146187
rect 149492 146113 149548 146122
rect 149396 144550 149452 144559
rect 149396 144485 149452 144494
rect 149410 144147 149438 144485
rect 149398 144141 149450 144147
rect 149398 144083 149450 144089
rect 149506 144073 149534 146113
rect 149494 144067 149546 144073
rect 149494 144009 149546 144015
rect 149492 143662 149548 143671
rect 149492 143597 149548 143606
rect 149396 142478 149452 142487
rect 149396 142413 149452 142422
rect 149410 141853 149438 142413
rect 149506 142371 149534 143597
rect 149494 142365 149546 142371
rect 149494 142307 149546 142313
rect 149398 141847 149450 141853
rect 149398 141789 149450 141795
rect 149396 138778 149452 138787
rect 149396 138713 149452 138722
rect 149410 138301 149438 138713
rect 149398 138295 149450 138301
rect 149398 138237 149450 138243
rect 149396 135966 149452 135975
rect 149396 135901 149452 135910
rect 149410 135489 149438 135901
rect 149398 135483 149450 135489
rect 149398 135425 149450 135431
rect 149602 135374 149630 172753
rect 149684 152098 149740 152107
rect 149684 152033 149740 152042
rect 149698 149845 149726 152033
rect 149686 149839 149738 149845
rect 149686 149781 149738 149787
rect 151138 141113 151166 226075
rect 151234 169677 151262 235917
rect 151414 229833 151466 229839
rect 151414 229775 151466 229781
rect 151318 226281 151370 226287
rect 151318 226223 151370 226229
rect 151222 169671 151274 169677
rect 151222 169613 151274 169619
rect 151330 161019 151358 226223
rect 151426 164127 151454 229775
rect 151798 217771 151850 217777
rect 151798 217713 151850 217719
rect 151702 211037 151754 211043
rect 151702 210979 151754 210985
rect 151606 210371 151658 210377
rect 151606 210313 151658 210319
rect 151510 207929 151562 207935
rect 151510 207871 151562 207877
rect 151414 164121 151466 164127
rect 151414 164063 151466 164069
rect 151318 161013 151370 161019
rect 151318 160955 151370 160961
rect 151414 158497 151466 158503
rect 151414 158439 151466 158445
rect 151222 156203 151274 156209
rect 151222 156145 151274 156151
rect 151126 141107 151178 141113
rect 151126 141049 151178 141055
rect 149684 137594 149740 137603
rect 149684 137529 149740 137538
rect 149698 135415 149726 137529
rect 149506 135346 149630 135374
rect 149686 135409 149738 135415
rect 149686 135351 149738 135357
rect 149396 135078 149452 135087
rect 149396 135013 149452 135022
rect 149410 132529 149438 135013
rect 149398 132523 149450 132529
rect 149398 132465 149450 132471
rect 149218 131040 149342 131068
rect 149218 129569 149246 131040
rect 149300 130934 149356 130943
rect 149300 130869 149356 130878
rect 149314 129643 149342 130869
rect 149396 130342 149452 130351
rect 149396 130277 149452 130286
rect 149410 129717 149438 130277
rect 149398 129711 149450 129717
rect 149398 129653 149450 129659
rect 149302 129637 149354 129643
rect 149302 129579 149354 129585
rect 149206 129563 149258 129569
rect 149206 129505 149258 129511
rect 149506 129495 149534 135346
rect 149590 134003 149642 134009
rect 149590 133945 149642 133951
rect 149494 129489 149546 129495
rect 149494 129431 149546 129437
rect 149110 129415 149162 129421
rect 149110 129357 149162 129363
rect 149108 129158 149164 129167
rect 149108 129093 149164 129102
rect 149122 103669 149150 129093
rect 149396 127974 149452 127983
rect 149396 127909 149452 127918
rect 149410 126757 149438 127909
rect 149398 126751 149450 126757
rect 149398 126693 149450 126699
rect 149300 126642 149356 126651
rect 149300 126577 149356 126586
rect 149110 103663 149162 103669
rect 149110 103605 149162 103611
rect 149014 103589 149066 103595
rect 149014 103531 149066 103537
rect 148916 102370 148972 102379
rect 148916 102305 148972 102314
rect 148822 89233 148874 89239
rect 148822 89175 148874 89181
rect 148724 86534 148780 86543
rect 148724 86469 148726 86478
rect 148778 86469 148780 86478
rect 148726 86437 148778 86443
rect 148438 86421 148490 86427
rect 148438 86363 148490 86369
rect 148246 86347 148298 86353
rect 148246 86289 148298 86295
rect 148930 86279 148958 102305
rect 149314 100709 149342 126577
rect 149602 125592 149630 133945
rect 149686 132967 149738 132973
rect 149686 132909 149738 132915
rect 149506 125564 149630 125592
rect 149506 120911 149534 125564
rect 149588 125458 149644 125467
rect 149588 125393 149644 125402
rect 149494 120905 149546 120911
rect 149494 120847 149546 120853
rect 149396 120574 149452 120583
rect 149396 120509 149452 120518
rect 149410 118321 149438 120509
rect 149492 119390 149548 119399
rect 149492 119325 149548 119334
rect 149398 118315 149450 118321
rect 149398 118257 149450 118263
rect 149506 118247 149534 119325
rect 149494 118241 149546 118247
rect 149396 118206 149452 118215
rect 149494 118183 149546 118189
rect 149396 118141 149398 118150
rect 149450 118141 149452 118150
rect 149398 118109 149450 118115
rect 149492 116874 149548 116883
rect 149492 116809 149548 116818
rect 149396 115690 149452 115699
rect 149396 115625 149452 115634
rect 149410 115361 149438 115625
rect 149398 115355 149450 115361
rect 149398 115297 149450 115303
rect 149506 115287 149534 116809
rect 149494 115281 149546 115287
rect 149396 115246 149452 115255
rect 149494 115223 149546 115229
rect 149396 115181 149452 115190
rect 149602 115214 149630 125393
rect 149698 123649 149726 132909
rect 149686 123643 149738 123649
rect 149686 123585 149738 123591
rect 149602 115186 149726 115214
rect 149410 114640 149438 115181
rect 149410 114612 149630 114640
rect 149492 114506 149548 114515
rect 149492 114441 149548 114450
rect 149396 113174 149452 113183
rect 149396 113109 149452 113118
rect 149410 112401 149438 113109
rect 149506 112771 149534 114441
rect 149494 112765 149546 112771
rect 149494 112707 149546 112713
rect 149398 112395 149450 112401
rect 149398 112337 149450 112343
rect 149396 109622 149452 109631
rect 149396 109557 149398 109566
rect 149450 109557 149452 109566
rect 149398 109525 149450 109531
rect 149602 106333 149630 114612
rect 149590 106327 149642 106333
rect 149590 106269 149642 106275
rect 149396 100890 149452 100899
rect 149396 100825 149398 100834
rect 149450 100825 149452 100834
rect 149398 100793 149450 100799
rect 149698 100783 149726 115186
rect 151234 112327 151262 156145
rect 151426 115213 151454 158439
rect 151522 149771 151550 207871
rect 151618 152583 151646 210313
rect 151606 152577 151658 152583
rect 151606 152519 151658 152525
rect 151714 152509 151742 210979
rect 151810 158429 151838 217713
rect 151990 212813 152042 212819
rect 151990 212755 152042 212761
rect 151894 207411 151946 207417
rect 151894 207353 151946 207359
rect 151798 158423 151850 158429
rect 151798 158365 151850 158371
rect 151906 152657 151934 207353
rect 152002 155543 152030 212755
rect 152086 206301 152138 206307
rect 152086 206243 152138 206249
rect 151990 155537 152042 155543
rect 151990 155479 152042 155485
rect 151894 152651 151946 152657
rect 151894 152593 151946 152599
rect 151702 152503 151754 152509
rect 151702 152445 151754 152451
rect 151510 149765 151562 149771
rect 151510 149707 151562 149713
rect 152098 149697 152126 206243
rect 152182 199345 152234 199351
rect 152182 199287 152234 199293
rect 152086 149691 152138 149697
rect 152086 149633 152138 149639
rect 152194 146663 152222 199287
rect 152386 192987 152414 271511
rect 154498 270761 154526 278018
rect 154486 270755 154538 270761
rect 154486 270697 154538 270703
rect 155446 270755 155498 270761
rect 155446 270697 155498 270703
rect 154006 252329 154058 252335
rect 154006 252271 154058 252277
rect 152374 192981 152426 192987
rect 152374 192923 152426 192929
rect 154018 181443 154046 252271
rect 154102 230499 154154 230505
rect 154102 230441 154154 230447
rect 154006 181437 154058 181443
rect 154006 181379 154058 181385
rect 154006 174407 154058 174413
rect 154006 174349 154058 174355
rect 152182 146657 152234 146663
rect 152182 146599 152234 146605
rect 154018 129347 154046 174349
rect 154114 164053 154142 230441
rect 154198 202897 154250 202903
rect 154198 202839 154250 202845
rect 154102 164047 154154 164053
rect 154102 163989 154154 163995
rect 154210 146811 154238 202839
rect 155458 192913 155486 270697
rect 155746 268911 155774 278018
rect 155734 268905 155786 268911
rect 155734 268847 155786 268853
rect 156898 268837 156926 278018
rect 158050 276494 158078 278018
rect 158050 276466 158174 276494
rect 156886 268831 156938 268837
rect 156886 268773 156938 268779
rect 156886 252403 156938 252409
rect 156886 252345 156938 252351
rect 155446 192907 155498 192913
rect 155446 192849 155498 192855
rect 154294 189577 154346 189583
rect 154294 189519 154346 189525
rect 154198 146805 154250 146811
rect 154198 146747 154250 146753
rect 154102 141255 154154 141261
rect 154102 141197 154154 141203
rect 154006 129341 154058 129347
rect 154006 129283 154058 129289
rect 151414 115207 151466 115213
rect 151414 115149 151466 115155
rect 154114 115139 154142 141197
rect 154306 141113 154334 189519
rect 156898 181369 156926 252345
rect 156982 249813 157034 249819
rect 156982 249755 157034 249761
rect 156994 184329 157022 249755
rect 157078 204229 157130 204235
rect 157078 204171 157130 204177
rect 156982 184323 157034 184329
rect 156982 184265 157034 184271
rect 156886 181363 156938 181369
rect 156886 181305 156938 181311
rect 156886 175813 156938 175819
rect 156886 175755 156938 175761
rect 154294 141107 154346 141113
rect 154294 141049 154346 141055
rect 156898 132455 156926 175755
rect 157090 149623 157118 204171
rect 158146 192839 158174 276466
rect 159298 271945 159326 278018
rect 160450 273573 160478 278018
rect 160438 273567 160490 273573
rect 160438 273509 160490 273515
rect 159286 271939 159338 271945
rect 159286 271881 159338 271887
rect 161602 271279 161630 278018
rect 161590 271273 161642 271279
rect 161590 271215 161642 271221
rect 162850 268763 162878 278018
rect 163894 271273 163946 271279
rect 163894 271215 163946 271221
rect 162838 268757 162890 268763
rect 162838 268699 162890 268705
rect 162742 249739 162794 249745
rect 162742 249681 162794 249687
rect 159766 249443 159818 249449
rect 159766 249385 159818 249391
rect 158134 192833 158186 192839
rect 158134 192775 158186 192781
rect 157174 190243 157226 190249
rect 157174 190185 157226 190191
rect 157078 149617 157130 149623
rect 157078 149559 157130 149565
rect 156982 141847 157034 141853
rect 156982 141789 157034 141795
rect 156886 132449 156938 132455
rect 156886 132391 156938 132397
rect 156886 126751 156938 126757
rect 156886 126693 156938 126699
rect 154198 123939 154250 123945
rect 154198 123881 154250 123887
rect 154102 115133 154154 115139
rect 154102 115075 154154 115081
rect 151222 112321 151274 112327
rect 151222 112263 151274 112269
rect 154006 108399 154058 108405
rect 154006 108341 154058 108347
rect 151126 107215 151178 107221
rect 151126 107157 151178 107163
rect 149686 100777 149738 100783
rect 149686 100719 149738 100725
rect 149302 100703 149354 100709
rect 149302 100645 149354 100651
rect 149492 99854 149548 99863
rect 149492 99789 149548 99798
rect 149396 98670 149452 98679
rect 149396 98605 149452 98614
rect 149410 98045 149438 98605
rect 149398 98039 149450 98045
rect 149398 97981 149450 97987
rect 149506 97971 149534 99789
rect 149494 97965 149546 97971
rect 149494 97907 149546 97913
rect 149492 97486 149548 97495
rect 149492 97421 149548 97430
rect 149396 95710 149452 95719
rect 149396 95645 149452 95654
rect 149410 95085 149438 95645
rect 149506 95159 149534 97421
rect 149494 95153 149546 95159
rect 149494 95095 149546 95101
rect 149398 95079 149450 95085
rect 149398 95021 149450 95027
rect 149588 94970 149644 94979
rect 149588 94905 149644 94914
rect 149492 93786 149548 93795
rect 149492 93721 149548 93730
rect 149396 92602 149452 92611
rect 149396 92537 149452 92546
rect 149410 92421 149438 92537
rect 149398 92415 149450 92421
rect 149398 92357 149450 92363
rect 149506 92199 149534 93721
rect 149494 92193 149546 92199
rect 149494 92135 149546 92141
rect 149300 91418 149356 91427
rect 149300 91353 149356 91362
rect 149204 90234 149260 90243
rect 149204 90169 149260 90178
rect 148918 86273 148970 86279
rect 148918 86215 148970 86221
rect 148628 85350 148684 85359
rect 148628 85285 148684 85294
rect 146996 84166 147052 84175
rect 146996 84101 147052 84110
rect 147010 83615 147038 84101
rect 146998 83609 147050 83615
rect 146998 83551 147050 83557
rect 148244 81650 148300 81659
rect 148244 81585 148300 81594
rect 148258 71997 148286 81585
rect 148642 74883 148670 85285
rect 148916 82390 148972 82399
rect 148916 82325 148972 82334
rect 148820 77950 148876 77959
rect 148820 77885 148876 77894
rect 148630 74877 148682 74883
rect 148630 74819 148682 74825
rect 148246 71991 148298 71997
rect 148246 71933 148298 71939
rect 148834 69111 148862 77885
rect 148930 74809 148958 82325
rect 149218 77621 149246 90169
rect 149314 77769 149342 91353
rect 149396 89050 149452 89059
rect 149396 88985 149452 88994
rect 149302 77763 149354 77769
rect 149302 77705 149354 77711
rect 149410 77695 149438 88985
rect 149492 87274 149548 87283
rect 149492 87209 149548 87218
rect 149506 86797 149534 87209
rect 149494 86791 149546 86797
rect 149494 86733 149546 86739
rect 149602 80655 149630 94905
rect 151138 89165 151166 107157
rect 151126 89159 151178 89165
rect 151126 89101 151178 89107
rect 154018 89091 154046 108341
rect 154210 108035 154238 123881
rect 154198 108029 154250 108035
rect 154198 107971 154250 107977
rect 156898 100635 156926 126693
rect 156994 115065 157022 141789
rect 157186 141039 157214 190185
rect 159778 178557 159806 249385
rect 159862 224801 159914 224807
rect 159862 224743 159914 224749
rect 159766 178551 159818 178557
rect 159766 178493 159818 178499
rect 159874 161167 159902 224743
rect 162646 219103 162698 219109
rect 162646 219045 162698 219051
rect 159958 213257 160010 213263
rect 159958 213199 160010 213205
rect 159862 161161 159914 161167
rect 159862 161103 159914 161109
rect 159766 157683 159818 157689
rect 159766 157625 159818 157631
rect 157174 141033 157226 141039
rect 157174 140975 157226 140981
rect 156982 115059 157034 115065
rect 156982 115001 157034 115007
rect 159778 114991 159806 157625
rect 159970 155469 159998 213199
rect 160054 200529 160106 200535
rect 160054 200471 160106 200477
rect 159958 155463 160010 155469
rect 159958 155405 160010 155411
rect 160066 146737 160094 200471
rect 162658 158355 162686 219045
rect 162754 187141 162782 249681
rect 163906 192765 163934 271215
rect 164002 268689 164030 278018
rect 165154 270761 165182 278018
rect 166306 271723 166334 278018
rect 167554 272093 167582 278018
rect 167542 272087 167594 272093
rect 167542 272029 167594 272035
rect 166294 271717 166346 271723
rect 166294 271659 166346 271665
rect 168706 270761 168734 278018
rect 169762 278004 169872 278032
rect 165142 270755 165194 270761
rect 165142 270697 165194 270703
rect 166966 270755 167018 270761
rect 166966 270697 167018 270703
rect 168694 270755 168746 270761
rect 168694 270697 168746 270703
rect 163990 268683 164042 268689
rect 163990 268625 164042 268631
rect 165526 252255 165578 252261
rect 165526 252197 165578 252203
rect 163894 192759 163946 192765
rect 163894 192701 163946 192707
rect 162838 190169 162890 190175
rect 162838 190111 162890 190117
rect 162742 187135 162794 187141
rect 162742 187077 162794 187083
rect 162742 178773 162794 178779
rect 162742 178715 162794 178721
rect 162646 158349 162698 158355
rect 162646 158291 162698 158297
rect 160054 146731 160106 146737
rect 160054 146673 160106 146679
rect 159862 142365 159914 142371
rect 159862 142307 159914 142313
rect 159874 118099 159902 142307
rect 162646 138295 162698 138301
rect 162646 138237 162698 138243
rect 159862 118093 159914 118099
rect 159862 118035 159914 118041
rect 159766 114985 159818 114991
rect 159766 114927 159818 114933
rect 159862 112765 159914 112771
rect 159862 112707 159914 112713
rect 156982 109583 157034 109589
rect 156982 109525 157034 109531
rect 156886 100629 156938 100635
rect 156886 100571 156938 100577
rect 154006 89085 154058 89091
rect 154006 89027 154058 89033
rect 156994 89017 157022 109525
rect 159574 92415 159626 92421
rect 159574 92357 159626 92363
rect 156982 89011 157034 89017
rect 156982 88953 157034 88959
rect 156406 86791 156458 86797
rect 156406 86733 156458 86739
rect 154102 86495 154154 86501
rect 154102 86437 154154 86443
rect 151126 83609 151178 83615
rect 151126 83551 151178 83557
rect 149590 80649 149642 80655
rect 149590 80591 149642 80597
rect 149588 80466 149644 80475
rect 149588 80401 149644 80410
rect 149398 77689 149450 77695
rect 149398 77631 149450 77637
rect 149206 77615 149258 77621
rect 149206 77557 149258 77563
rect 149396 76766 149452 76775
rect 149396 76701 149452 76710
rect 149204 75582 149260 75591
rect 149204 75517 149260 75526
rect 148918 74803 148970 74809
rect 148918 74745 148970 74751
rect 149012 73066 149068 73075
rect 149012 73001 149068 73010
rect 148822 69105 148874 69111
rect 148822 69047 148874 69053
rect 149026 66003 149054 73001
rect 149108 72030 149164 72039
rect 149108 71965 149164 71974
rect 149122 66225 149150 71965
rect 149218 68889 149246 75517
rect 149410 74894 149438 76701
rect 149410 74866 149534 74894
rect 149300 73806 149356 73815
rect 149300 73741 149356 73750
rect 149314 68963 149342 73741
rect 149506 70980 149534 74866
rect 149602 71923 149630 80401
rect 149684 79282 149740 79291
rect 149684 79217 149740 79226
rect 149590 71917 149642 71923
rect 149590 71859 149642 71865
rect 149698 71849 149726 79217
rect 151138 74735 151166 83551
rect 151126 74729 151178 74735
rect 151126 74671 151178 74677
rect 154114 74661 154142 86437
rect 156418 77547 156446 86733
rect 159586 80581 159614 92357
rect 159874 91977 159902 112707
rect 162658 109441 162686 138237
rect 162754 135341 162782 178715
rect 162850 140965 162878 190111
rect 165538 181295 165566 252197
rect 165622 249591 165674 249597
rect 165622 249533 165674 249539
rect 165634 184255 165662 249533
rect 165718 204525 165770 204531
rect 165718 204467 165770 204473
rect 165622 184249 165674 184255
rect 165622 184191 165674 184197
rect 165526 181289 165578 181295
rect 165526 181231 165578 181237
rect 165526 175739 165578 175745
rect 165526 175681 165578 175687
rect 162934 144141 162986 144147
rect 162934 144083 162986 144089
rect 162838 140959 162890 140965
rect 162838 140901 162890 140907
rect 162742 135335 162794 135341
rect 162742 135277 162794 135283
rect 162946 118025 162974 144083
rect 165538 132381 165566 175681
rect 165730 149549 165758 204467
rect 166978 195799 167006 270697
rect 169762 268615 169790 278004
rect 169846 270755 169898 270761
rect 169846 270697 169898 270703
rect 169750 268609 169802 268615
rect 169750 268551 169802 268557
rect 168502 249665 168554 249671
rect 168502 249607 168554 249613
rect 168406 219029 168458 219035
rect 168406 218971 168458 218977
rect 166966 195793 167018 195799
rect 166966 195735 167018 195741
rect 165814 193129 165866 193135
rect 165814 193071 165866 193077
rect 165718 149543 165770 149549
rect 165718 149485 165770 149491
rect 165718 144067 165770 144073
rect 165718 144009 165770 144015
rect 165526 132375 165578 132381
rect 165526 132317 165578 132323
rect 165622 129711 165674 129717
rect 165622 129653 165674 129659
rect 162934 118019 162986 118025
rect 162934 117961 162986 117967
rect 162742 115355 162794 115361
rect 162742 115297 162794 115303
rect 162646 109435 162698 109441
rect 162646 109377 162698 109383
rect 162754 95011 162782 115297
rect 165526 115281 165578 115287
rect 165526 115223 165578 115229
rect 162742 95005 162794 95011
rect 162742 94947 162794 94953
rect 165538 94937 165566 115223
rect 165634 103521 165662 129653
rect 165730 117951 165758 144009
rect 165826 140891 165854 193071
rect 168418 158281 168446 218971
rect 168514 187067 168542 249607
rect 169858 195725 169886 270697
rect 171106 268541 171134 278018
rect 172272 278004 172766 278032
rect 171094 268535 171146 268541
rect 171094 268477 171146 268483
rect 171286 252181 171338 252187
rect 171286 252123 171338 252129
rect 169846 195719 169898 195725
rect 169846 195661 169898 195667
rect 168598 193055 168650 193061
rect 168598 192997 168650 193003
rect 168502 187061 168554 187067
rect 168502 187003 168554 187009
rect 168502 178699 168554 178705
rect 168502 178641 168554 178647
rect 168406 158275 168458 158281
rect 168406 158217 168458 158223
rect 168406 147027 168458 147033
rect 168406 146969 168458 146975
rect 165814 140885 165866 140891
rect 165814 140827 165866 140833
rect 165718 117945 165770 117951
rect 165718 117887 165770 117893
rect 168418 117877 168446 146969
rect 168514 132307 168542 178641
rect 168610 143999 168638 192997
rect 171298 181221 171326 252123
rect 171478 249887 171530 249893
rect 171478 249829 171530 249835
rect 171382 221915 171434 221921
rect 171382 221857 171434 221863
rect 171286 181215 171338 181221
rect 171286 181157 171338 181163
rect 171394 161093 171422 221857
rect 171490 189953 171518 249829
rect 171574 196015 171626 196021
rect 171574 195957 171626 195963
rect 171478 189947 171530 189953
rect 171478 189889 171530 189895
rect 171478 178625 171530 178631
rect 171478 178567 171530 178573
rect 171382 161087 171434 161093
rect 171382 161029 171434 161035
rect 171382 146953 171434 146959
rect 171382 146895 171434 146901
rect 168598 143993 168650 143999
rect 168598 143935 168650 143941
rect 171286 132523 171338 132529
rect 171286 132465 171338 132471
rect 168502 132301 168554 132307
rect 168502 132243 168554 132249
rect 168502 118315 168554 118321
rect 168502 118257 168554 118263
rect 168406 117871 168458 117877
rect 168406 117813 168458 117819
rect 165622 103515 165674 103521
rect 165622 103457 165674 103463
rect 168406 100851 168458 100857
rect 168406 100793 168458 100799
rect 166678 95153 166730 95159
rect 166678 95095 166730 95101
rect 165526 94931 165578 94937
rect 165526 94873 165578 94879
rect 162358 92193 162410 92199
rect 162358 92135 162410 92141
rect 159862 91971 159914 91977
rect 159862 91913 159914 91919
rect 159574 80575 159626 80581
rect 159574 80517 159626 80523
rect 162370 80507 162398 92135
rect 166690 83541 166718 95095
rect 166678 83535 166730 83541
rect 166678 83477 166730 83483
rect 168418 83467 168446 100793
rect 168514 97749 168542 118257
rect 171298 106481 171326 132465
rect 171394 120837 171422 146895
rect 171490 132233 171518 178567
rect 171586 143925 171614 195957
rect 172738 195651 172766 278004
rect 173410 271501 173438 278018
rect 174658 272019 174686 278018
rect 174646 272013 174698 272019
rect 174646 271955 174698 271961
rect 173398 271495 173450 271501
rect 173398 271437 173450 271443
rect 175810 271205 175838 278018
rect 175798 271199 175850 271205
rect 175798 271141 175850 271147
rect 176962 268467 176990 278018
rect 176950 268461 177002 268467
rect 176950 268403 177002 268409
rect 178210 268393 178238 278018
rect 178294 271199 178346 271205
rect 178294 271141 178346 271147
rect 178198 268387 178250 268393
rect 178198 268329 178250 268335
rect 174262 252477 174314 252483
rect 174262 252419 174314 252425
rect 174166 224875 174218 224881
rect 174166 224817 174218 224823
rect 172726 195645 172778 195651
rect 172726 195587 172778 195593
rect 174178 163979 174206 224817
rect 174274 189879 174302 252419
rect 177046 249295 177098 249301
rect 177046 249237 177098 249243
rect 174358 213183 174410 213189
rect 174358 213125 174410 213131
rect 174262 189873 174314 189879
rect 174262 189815 174314 189821
rect 174166 163973 174218 163979
rect 174166 163915 174218 163921
rect 174370 155395 174398 213125
rect 174454 195941 174506 195947
rect 174454 195883 174506 195889
rect 174358 155389 174410 155395
rect 174358 155331 174410 155337
rect 172822 152799 172874 152805
rect 172822 152741 172874 152747
rect 171574 143919 171626 143925
rect 171574 143861 171626 143867
rect 172834 136821 172862 152741
rect 174262 149987 174314 149993
rect 174262 149929 174314 149935
rect 172822 136815 172874 136821
rect 172822 136757 172874 136763
rect 174166 135483 174218 135489
rect 174166 135425 174218 135431
rect 171478 132227 171530 132233
rect 171478 132169 171530 132175
rect 171382 120831 171434 120837
rect 171382 120773 171434 120779
rect 171286 106475 171338 106481
rect 171286 106417 171338 106423
rect 174178 106407 174206 135425
rect 174274 120763 174302 149929
rect 174466 143851 174494 195883
rect 177058 178409 177086 249237
rect 177142 227613 177194 227619
rect 177142 227555 177194 227561
rect 177046 178403 177098 178409
rect 177046 178345 177098 178351
rect 177154 163905 177182 227555
rect 177238 216069 177290 216075
rect 177238 216011 177290 216017
rect 177142 163899 177194 163905
rect 177142 163841 177194 163847
rect 177250 155321 177278 216011
rect 178306 198611 178334 271141
rect 179362 270761 179390 278018
rect 180514 271575 180542 278018
rect 181762 271649 181790 278018
rect 181750 271643 181802 271649
rect 181750 271585 181802 271591
rect 180502 271569 180554 271575
rect 180502 271511 180554 271517
rect 182914 270761 182942 278018
rect 184066 271353 184094 278018
rect 185218 271427 185246 278018
rect 185206 271421 185258 271427
rect 185206 271363 185258 271369
rect 184054 271347 184106 271353
rect 184054 271289 184106 271295
rect 186466 270761 186494 278018
rect 187618 271205 187646 278018
rect 188770 271279 188798 278018
rect 189730 278004 190032 278032
rect 188758 271273 188810 271279
rect 188758 271215 188810 271221
rect 187606 271199 187658 271205
rect 187606 271141 187658 271147
rect 179350 270755 179402 270761
rect 179350 270697 179402 270703
rect 181366 270755 181418 270761
rect 181366 270697 181418 270703
rect 182902 270755 182954 270761
rect 182902 270697 182954 270703
rect 184246 270755 184298 270761
rect 184246 270697 184298 270703
rect 185494 270755 185546 270761
rect 185494 270697 185546 270703
rect 186454 270755 186506 270761
rect 186454 270697 186506 270703
rect 179926 252107 179978 252113
rect 179926 252049 179978 252055
rect 178294 198605 178346 198611
rect 178294 198547 178346 198553
rect 179938 184181 179966 252049
rect 180118 249517 180170 249523
rect 180118 249459 180170 249465
rect 180022 218955 180074 218961
rect 180022 218897 180074 218903
rect 179926 184175 179978 184181
rect 179926 184117 179978 184123
rect 177334 181585 177386 181591
rect 177334 181527 177386 181533
rect 177238 155315 177290 155321
rect 177238 155257 177290 155263
rect 177046 149913 177098 149919
rect 177046 149855 177098 149861
rect 174454 143845 174506 143851
rect 174454 143787 174506 143793
rect 174262 120757 174314 120763
rect 174262 120699 174314 120705
rect 174358 118241 174410 118247
rect 174358 118183 174410 118189
rect 174166 106401 174218 106407
rect 174166 106343 174218 106349
rect 168502 97743 168554 97749
rect 168502 97685 168554 97691
rect 174370 94863 174398 118183
rect 177058 109293 177086 149855
rect 177346 134897 177374 181527
rect 180034 158207 180062 218897
rect 180130 186993 180158 249459
rect 181378 198685 181406 270697
rect 182806 249221 182858 249227
rect 182806 249163 182858 249169
rect 181366 198679 181418 198685
rect 181366 198621 181418 198627
rect 180214 195867 180266 195873
rect 180214 195809 180266 195815
rect 180118 186987 180170 186993
rect 180118 186929 180170 186935
rect 180022 158201 180074 158207
rect 180022 158143 180074 158149
rect 179926 152725 179978 152731
rect 179926 152667 179978 152673
rect 177334 134891 177386 134897
rect 177334 134833 177386 134839
rect 177238 129637 177290 129643
rect 177238 129579 177290 129585
rect 177250 113955 177278 129579
rect 177238 113949 177290 113955
rect 177238 113891 177290 113897
rect 177142 112395 177194 112401
rect 177142 112337 177194 112343
rect 177046 109287 177098 109293
rect 177046 109229 177098 109235
rect 174358 94857 174410 94863
rect 174358 94799 174410 94805
rect 177154 91903 177182 112337
rect 179938 109367 179966 152667
rect 180022 149839 180074 149845
rect 180022 149781 180074 149787
rect 180034 120689 180062 149781
rect 180226 143777 180254 195809
rect 182818 178483 182846 249163
rect 182902 221841 182954 221847
rect 182902 221783 182954 221789
rect 182806 178477 182858 178483
rect 182806 178419 182858 178425
rect 182914 161241 182942 221783
rect 182998 201639 183050 201645
rect 182998 201581 183050 201587
rect 182902 161235 182954 161241
rect 182902 161177 182954 161183
rect 182806 155759 182858 155765
rect 182806 155701 182858 155707
rect 180214 143771 180266 143777
rect 180214 143713 180266 143719
rect 180022 120683 180074 120689
rect 180022 120625 180074 120631
rect 180118 118167 180170 118173
rect 180118 118109 180170 118115
rect 179926 109361 179978 109367
rect 179926 109303 179978 109309
rect 179926 95079 179978 95085
rect 179926 95021 179978 95027
rect 177142 91897 177194 91903
rect 177142 91839 177194 91845
rect 168406 83461 168458 83467
rect 168406 83403 168458 83409
rect 162358 80501 162410 80507
rect 162358 80443 162410 80449
rect 179938 80433 179966 95021
rect 180130 94641 180158 118109
rect 182818 112253 182846 155701
rect 183010 146885 183038 201581
rect 184258 197691 184286 270697
rect 184342 221767 184394 221773
rect 184342 221709 184394 221715
rect 184354 219595 184382 221709
rect 184340 219586 184396 219595
rect 184340 219521 184396 219530
rect 184342 218881 184394 218887
rect 184340 218846 184342 218855
rect 184394 218846 184396 218855
rect 184340 218781 184396 218790
rect 184342 201565 184394 201571
rect 184342 201507 184394 201513
rect 184354 199763 184382 201507
rect 184340 199754 184396 199763
rect 184340 199689 184396 199698
rect 184342 198679 184394 198685
rect 184342 198621 184394 198627
rect 184244 197682 184300 197691
rect 184244 197617 184300 197626
rect 184354 196803 184382 198621
rect 184438 198605 184490 198611
rect 184438 198547 184490 198553
rect 184340 196794 184396 196803
rect 184340 196729 184396 196738
rect 184450 196063 184478 198547
rect 185506 198283 185534 270697
rect 185686 269867 185738 269873
rect 185686 269809 185738 269815
rect 185698 268319 185726 269809
rect 185686 268313 185738 268319
rect 185686 268255 185738 268261
rect 189730 266469 189758 278004
rect 190102 273493 190154 273499
rect 190102 273435 190154 273441
rect 190114 268171 190142 273435
rect 191170 271871 191198 278018
rect 191158 271865 191210 271871
rect 191158 271807 191210 271813
rect 192322 271797 192350 278018
rect 193570 273499 193598 278018
rect 193558 273493 193610 273499
rect 193558 273435 193610 273441
rect 194420 272274 194476 272283
rect 194420 272209 194476 272218
rect 193748 272126 193804 272135
rect 193748 272061 193804 272070
rect 192982 271939 193034 271945
rect 192982 271881 193034 271887
rect 192310 271791 192362 271797
rect 192310 271733 192362 271739
rect 192404 269314 192460 269323
rect 192404 269249 192460 269258
rect 192598 269275 192650 269281
rect 190102 268165 190154 268171
rect 190102 268107 190154 268113
rect 187222 266463 187274 266469
rect 187222 266405 187274 266411
rect 189718 266463 189770 266469
rect 189718 266405 189770 266411
rect 186358 255067 186410 255073
rect 186358 255009 186410 255015
rect 185974 254993 186026 254999
rect 185974 254935 186026 254941
rect 185782 246705 185834 246711
rect 185782 246647 185834 246653
rect 185686 242857 185738 242863
rect 185686 242799 185738 242805
rect 185590 242783 185642 242789
rect 185590 242725 185642 242731
rect 185602 220335 185630 242725
rect 185588 220326 185644 220335
rect 185588 220261 185644 220270
rect 185492 198274 185548 198283
rect 185492 198209 185548 198218
rect 184436 196054 184492 196063
rect 184436 195989 184492 195998
rect 184534 195793 184586 195799
rect 184534 195735 184586 195741
rect 184438 195719 184490 195725
rect 184438 195661 184490 195667
rect 184342 195645 184394 195651
rect 184342 195587 184394 195593
rect 184354 195323 184382 195587
rect 184340 195314 184396 195323
rect 184340 195249 184396 195258
rect 184450 194435 184478 195661
rect 184436 194426 184492 194435
rect 184436 194361 184492 194370
rect 184546 193843 184574 195735
rect 184532 193834 184588 193843
rect 184532 193769 184588 193778
rect 184630 192981 184682 192987
rect 184436 192946 184492 192955
rect 184630 192923 184682 192929
rect 184436 192881 184492 192890
rect 184534 192907 184586 192913
rect 184342 192833 184394 192839
rect 184342 192775 184394 192781
rect 184354 192363 184382 192775
rect 184450 192765 184478 192881
rect 184534 192849 184586 192855
rect 184438 192759 184490 192765
rect 184438 192701 184490 192707
rect 184340 192354 184396 192363
rect 184340 192289 184396 192298
rect 184546 191475 184574 192849
rect 184532 191466 184588 191475
rect 184532 191401 184588 191410
rect 184642 190735 184670 192923
rect 184628 190726 184684 190735
rect 184628 190661 184684 190670
rect 184534 190095 184586 190101
rect 184534 190037 184586 190043
rect 184342 190021 184394 190027
rect 184340 189986 184342 189995
rect 184394 189986 184396 189995
rect 184340 189921 184396 189930
rect 184438 189947 184490 189953
rect 184438 189889 184490 189895
rect 184342 189873 184394 189879
rect 184342 189815 184394 189821
rect 184354 188515 184382 189815
rect 184340 188506 184396 188515
rect 184340 188441 184396 188450
rect 184450 187627 184478 189889
rect 184546 189255 184574 190037
rect 184532 189246 184588 189255
rect 184532 189181 184588 189190
rect 184436 187618 184492 187627
rect 184436 187553 184492 187562
rect 184342 187209 184394 187215
rect 184342 187151 184394 187157
rect 184354 186887 184382 187151
rect 184534 187135 184586 187141
rect 184534 187077 184586 187083
rect 184438 187061 184490 187067
rect 184438 187003 184490 187009
rect 184340 186878 184396 186887
rect 184340 186813 184396 186822
rect 184450 185407 184478 187003
rect 184436 185398 184492 185407
rect 184436 185333 184492 185342
rect 184546 184667 184574 187077
rect 185398 186987 185450 186993
rect 185398 186929 185450 186935
rect 185410 186147 185438 186929
rect 185396 186138 185452 186147
rect 185396 186073 185452 186082
rect 184532 184658 184588 184667
rect 184532 184593 184588 184602
rect 184438 184323 184490 184329
rect 184438 184265 184490 184271
rect 184342 184249 184394 184255
rect 184342 184191 184394 184197
rect 184354 183927 184382 184191
rect 184340 183918 184396 183927
rect 184340 183853 184396 183862
rect 184450 183187 184478 184265
rect 184534 184175 184586 184181
rect 184534 184117 184586 184123
rect 184436 183178 184492 183187
rect 184436 183113 184492 183122
rect 184546 181559 184574 184117
rect 184532 181550 184588 181559
rect 183094 181511 183146 181517
rect 184532 181485 184588 181494
rect 183094 181453 183146 181459
rect 182998 146879 183050 146885
rect 182998 146821 183050 146827
rect 182902 135409 182954 135415
rect 182902 135351 182954 135357
rect 182806 112247 182858 112253
rect 182806 112189 182858 112195
rect 182914 106555 182942 135351
rect 183106 134971 183134 181453
rect 184630 181437 184682 181443
rect 184630 181379 184682 181385
rect 184534 181363 184586 181369
rect 184534 181305 184586 181311
rect 184438 181289 184490 181295
rect 184438 181231 184490 181237
rect 184342 181215 184394 181221
rect 184342 181157 184394 181163
rect 184354 180819 184382 181157
rect 184340 180810 184396 180819
rect 184340 180745 184396 180754
rect 184450 180079 184478 181231
rect 184436 180070 184492 180079
rect 184436 180005 184492 180014
rect 184546 179339 184574 181305
rect 184532 179330 184588 179339
rect 184532 179265 184588 179274
rect 184642 178599 184670 181379
rect 185398 180031 185450 180037
rect 185398 179973 185450 179979
rect 184628 178590 184684 178599
rect 184342 178551 184394 178557
rect 184628 178525 184684 178534
rect 184342 178493 184394 178499
rect 184354 177711 184382 178493
rect 184534 178477 184586 178483
rect 184534 178419 184586 178425
rect 184438 178403 184490 178409
rect 184438 178345 184490 178351
rect 184340 177702 184396 177711
rect 184340 177637 184396 177646
rect 184450 177119 184478 178345
rect 184436 177110 184492 177119
rect 184436 177045 184492 177054
rect 184546 176231 184574 178419
rect 184532 176222 184588 176231
rect 184532 176157 184588 176166
rect 184438 175665 184490 175671
rect 184340 175630 184396 175639
rect 184438 175607 184490 175613
rect 184340 175565 184342 175574
rect 184394 175565 184396 175574
rect 184342 175533 184394 175539
rect 184450 174011 184478 175607
rect 184436 174002 184492 174011
rect 184436 173937 184492 173946
rect 184534 172779 184586 172785
rect 184534 172721 184586 172727
rect 184342 172705 184394 172711
rect 184342 172647 184394 172653
rect 184354 172531 184382 172647
rect 184438 172557 184490 172563
rect 184340 172522 184396 172531
rect 184438 172499 184490 172505
rect 184340 172457 184396 172466
rect 184450 170903 184478 172499
rect 184546 171791 184574 172721
rect 184630 172631 184682 172637
rect 184630 172573 184682 172579
rect 184532 171782 184588 171791
rect 184532 171717 184588 171726
rect 184436 170894 184492 170903
rect 184436 170829 184492 170838
rect 184642 170311 184670 172573
rect 184628 170302 184684 170311
rect 184628 170237 184684 170246
rect 184534 169893 184586 169899
rect 184534 169835 184586 169841
rect 184342 169745 184394 169751
rect 184342 169687 184394 169693
rect 184354 169423 184382 169687
rect 184438 169671 184490 169677
rect 184438 169613 184490 169619
rect 184340 169414 184396 169423
rect 184340 169349 184396 169358
rect 184450 167203 184478 169613
rect 184546 168683 184574 169835
rect 184630 169819 184682 169825
rect 184630 169761 184682 169767
rect 184532 168674 184588 168683
rect 184532 168609 184588 168618
rect 184642 167943 184670 169761
rect 184628 167934 184684 167943
rect 184628 167869 184684 167878
rect 184436 167194 184492 167203
rect 184436 167129 184492 167138
rect 184534 167007 184586 167013
rect 184534 166949 184586 166955
rect 184342 166933 184394 166939
rect 184342 166875 184394 166881
rect 184354 166463 184382 166875
rect 184438 166859 184490 166865
rect 184438 166801 184490 166807
rect 184340 166454 184396 166463
rect 184340 166389 184396 166398
rect 184450 164835 184478 166801
rect 184546 165723 184574 166949
rect 184532 165714 184588 165723
rect 184532 165649 184588 165658
rect 185410 165626 185438 179973
rect 185698 173271 185726 242799
rect 185794 205937 185822 246647
rect 185878 242709 185930 242715
rect 185878 242651 185930 242657
rect 185782 205931 185834 205937
rect 185782 205873 185834 205879
rect 185890 174751 185918 242651
rect 185986 204351 186014 254935
rect 186070 246631 186122 246637
rect 186070 246573 186122 246579
rect 186082 205979 186110 246573
rect 186262 246557 186314 246563
rect 186262 246499 186314 246505
rect 186166 246483 186218 246489
rect 186166 246425 186218 246431
rect 186068 205970 186124 205979
rect 186068 205905 186124 205914
rect 185972 204342 186028 204351
rect 185972 204277 186028 204286
rect 186178 202871 186206 246425
rect 186274 207311 186302 246499
rect 186370 213527 186398 255009
rect 186550 254919 186602 254925
rect 186550 254861 186602 254867
rect 186454 252033 186506 252039
rect 186454 251975 186506 251981
rect 186356 213518 186412 213527
rect 186356 213453 186412 213462
rect 186466 210567 186494 251975
rect 186562 215007 186590 254861
rect 186742 249147 186794 249153
rect 186742 249089 186794 249095
rect 186646 246409 186698 246415
rect 186646 246351 186698 246357
rect 186548 214998 186604 215007
rect 186548 214933 186604 214942
rect 186452 210558 186508 210567
rect 186452 210493 186508 210502
rect 186658 209087 186686 246351
rect 186754 212047 186782 249089
rect 186838 246335 186890 246341
rect 186838 246277 186890 246283
rect 186850 216487 186878 246277
rect 187030 246261 187082 246267
rect 187030 246203 187082 246209
rect 186934 244929 186986 244935
rect 186934 244871 186986 244877
rect 186946 221075 186974 244871
rect 186932 221066 186988 221075
rect 186932 221001 186988 221010
rect 187042 218115 187070 246203
rect 187124 243414 187180 243423
rect 187124 243349 187180 243358
rect 187138 227545 187166 243349
rect 187126 227539 187178 227545
rect 187126 227481 187178 227487
rect 187138 226139 187166 227481
rect 187126 226133 187178 226139
rect 187126 226075 187178 226081
rect 187028 218106 187084 218115
rect 187028 218041 187084 218050
rect 186836 216478 186892 216487
rect 186836 216413 186892 216422
rect 186740 212038 186796 212047
rect 186740 211973 186796 211982
rect 186644 209078 186700 209087
rect 186644 209013 186700 209022
rect 186260 207302 186316 207311
rect 186260 207237 186316 207246
rect 186262 205931 186314 205937
rect 186262 205873 186314 205879
rect 186164 202862 186220 202871
rect 186164 202797 186220 202806
rect 185974 182991 186026 182997
rect 185974 182933 186026 182939
rect 185876 174742 185932 174751
rect 185876 174677 185932 174686
rect 185684 173262 185740 173271
rect 185684 173197 185740 173206
rect 185410 165598 185726 165626
rect 184436 164826 184492 164835
rect 184436 164761 184492 164770
rect 184534 164121 184586 164127
rect 184340 164086 184396 164095
rect 184534 164063 184586 164069
rect 184340 164021 184342 164030
rect 184394 164021 184396 164030
rect 184342 163989 184394 163995
rect 184438 163973 184490 163979
rect 184438 163915 184490 163921
rect 184342 163899 184394 163905
rect 184342 163841 184394 163847
rect 184354 162615 184382 163841
rect 184340 162606 184396 162615
rect 184340 162541 184396 162550
rect 184450 161875 184478 163915
rect 184546 163355 184574 164063
rect 184532 163346 184588 163355
rect 184532 163281 184588 163290
rect 184436 161866 184492 161875
rect 184436 161801 184492 161810
rect 184630 161235 184682 161241
rect 184630 161177 184682 161183
rect 184438 161161 184490 161167
rect 184438 161103 184490 161109
rect 184342 161013 184394 161019
rect 184340 160978 184342 160987
rect 184394 160978 184396 160987
rect 184340 160913 184396 160922
rect 184450 160395 184478 161103
rect 184534 161087 184586 161093
rect 184534 161029 184586 161035
rect 184436 160386 184492 160395
rect 184436 160321 184492 160330
rect 184546 158915 184574 161029
rect 184642 159507 184670 161177
rect 184628 159498 184684 159507
rect 184628 159433 184684 159442
rect 184532 158906 184588 158915
rect 184532 158841 184588 158850
rect 184534 158423 184586 158429
rect 184534 158365 184586 158371
rect 184438 158349 184490 158355
rect 184438 158291 184490 158297
rect 184342 158275 184394 158281
rect 184342 158217 184394 158223
rect 184354 158027 184382 158217
rect 184340 158018 184396 158027
rect 184340 157953 184396 157962
rect 184450 157435 184478 158291
rect 184436 157426 184492 157435
rect 184436 157361 184492 157370
rect 184546 155659 184574 158365
rect 184630 158201 184682 158207
rect 184630 158143 184682 158149
rect 184642 156547 184670 158143
rect 184628 156538 184684 156547
rect 184628 156473 184684 156482
rect 184532 155650 184588 155659
rect 184532 155585 184588 155594
rect 184630 155537 184682 155543
rect 185698 155534 185726 165598
rect 185698 155506 185822 155534
rect 184630 155479 184682 155485
rect 184342 155463 184394 155469
rect 184342 155405 184394 155411
rect 184354 154179 184382 155405
rect 184438 155389 184490 155395
rect 184438 155331 184490 155337
rect 184340 154170 184396 154179
rect 184340 154105 184396 154114
rect 184450 153587 184478 155331
rect 184534 155315 184586 155321
rect 184534 155257 184586 155263
rect 184546 155067 184574 155257
rect 184532 155058 184588 155067
rect 184532 154993 184588 155002
rect 184436 153578 184492 153587
rect 184436 153513 184492 153522
rect 184642 152699 184670 155479
rect 184628 152690 184684 152699
rect 184534 152651 184586 152657
rect 184628 152625 184684 152634
rect 184534 152593 184586 152599
rect 184438 152577 184490 152583
rect 184438 152519 184490 152525
rect 184342 152503 184394 152509
rect 184342 152445 184394 152451
rect 184354 151959 184382 152445
rect 184340 151950 184396 151959
rect 184340 151885 184396 151894
rect 184450 151219 184478 152519
rect 184436 151210 184492 151219
rect 184436 151145 184492 151154
rect 184546 150479 184574 152593
rect 184532 150470 184588 150479
rect 184532 150405 184588 150414
rect 184342 149765 184394 149771
rect 184340 149730 184342 149739
rect 184394 149730 184396 149739
rect 184340 149665 184396 149674
rect 184438 149691 184490 149697
rect 184438 149633 184490 149639
rect 184342 149543 184394 149549
rect 184342 149485 184394 149491
rect 184354 148111 184382 149485
rect 184450 148999 184478 149633
rect 184534 149617 184586 149623
rect 184534 149559 184586 149565
rect 184436 148990 184492 148999
rect 184436 148925 184492 148934
rect 184340 148102 184396 148111
rect 184340 148037 184396 148046
rect 184546 147371 184574 149559
rect 184532 147362 184588 147371
rect 184532 147297 184588 147306
rect 184342 146805 184394 146811
rect 184342 146747 184394 146753
rect 184354 146631 184382 146747
rect 184438 146731 184490 146737
rect 184438 146673 184490 146679
rect 184340 146622 184396 146631
rect 184340 146557 184396 146566
rect 184450 145151 184478 146673
rect 184534 146657 184586 146663
rect 184534 146599 184586 146605
rect 184436 145142 184492 145151
rect 184436 145077 184492 145086
rect 184546 144411 184574 146599
rect 184532 144402 184588 144411
rect 184532 144337 184588 144346
rect 184534 143993 184586 143999
rect 184534 143935 184586 143941
rect 184438 143919 184490 143925
rect 184438 143861 184490 143867
rect 184342 143845 184394 143851
rect 184342 143787 184394 143793
rect 184354 142783 184382 143787
rect 184340 142774 184396 142783
rect 184340 142709 184396 142718
rect 184450 142191 184478 143861
rect 184436 142182 184492 142191
rect 184436 142117 184492 142126
rect 184546 141303 184574 143935
rect 185398 143771 185450 143777
rect 185398 143713 185450 143719
rect 185410 143671 185438 143713
rect 185396 143662 185452 143671
rect 185396 143597 185452 143606
rect 184532 141294 184588 141303
rect 184532 141229 184588 141238
rect 184630 141107 184682 141113
rect 184630 141049 184682 141055
rect 184534 141033 184586 141039
rect 184534 140975 184586 140981
rect 184438 140959 184490 140965
rect 184438 140901 184490 140907
rect 184342 140885 184394 140891
rect 184342 140827 184394 140833
rect 184354 140563 184382 140827
rect 184340 140554 184396 140563
rect 184340 140489 184396 140498
rect 184450 139823 184478 140901
rect 184436 139814 184492 139823
rect 184436 139749 184492 139758
rect 184546 138935 184574 140975
rect 184532 138926 184588 138935
rect 184532 138861 184588 138870
rect 184642 138343 184670 141049
rect 184628 138334 184684 138343
rect 184628 138269 184684 138278
rect 185686 136815 185738 136821
rect 185686 136757 185738 136763
rect 184342 135335 184394 135341
rect 184342 135277 184394 135283
rect 183094 134965 183146 134971
rect 183094 134907 183146 134913
rect 184354 133015 184382 135277
rect 184534 134965 184586 134971
rect 184534 134907 184586 134913
rect 184438 134891 184490 134897
rect 184438 134833 184490 134839
rect 184450 134495 184478 134833
rect 184436 134486 184492 134495
rect 184436 134421 184492 134430
rect 184546 133755 184574 134907
rect 184532 133746 184588 133755
rect 184532 133681 184588 133690
rect 184340 133006 184396 133015
rect 184340 132941 184396 132950
rect 184630 132449 184682 132455
rect 184630 132391 184682 132397
rect 184534 132375 184586 132381
rect 184534 132317 184586 132323
rect 184438 132301 184490 132307
rect 184340 132266 184396 132275
rect 184438 132243 184490 132249
rect 184340 132201 184342 132210
rect 184394 132201 184396 132210
rect 184342 132169 184394 132175
rect 184450 131535 184478 132243
rect 184436 131526 184492 131535
rect 184436 131461 184492 131470
rect 184546 130647 184574 132317
rect 184532 130638 184588 130647
rect 184532 130573 184588 130582
rect 184642 129907 184670 132391
rect 184628 129898 184684 129907
rect 184628 129833 184684 129842
rect 184438 129563 184490 129569
rect 184438 129505 184490 129511
rect 184342 129341 184394 129347
rect 184342 129283 184394 129289
rect 184354 129167 184382 129283
rect 184340 129158 184396 129167
rect 184340 129093 184396 129102
rect 184450 128427 184478 129505
rect 184534 129489 184586 129495
rect 184534 129431 184586 129437
rect 184436 128418 184492 128427
rect 184436 128353 184492 128362
rect 184546 127687 184574 129431
rect 184630 129415 184682 129421
rect 184630 129357 184682 129363
rect 184532 127678 184588 127687
rect 184532 127613 184588 127622
rect 184642 126947 184670 129357
rect 184628 126938 184684 126947
rect 184628 126873 184684 126882
rect 184534 126677 184586 126683
rect 184534 126619 184586 126625
rect 184438 126603 184490 126609
rect 184438 126545 184490 126551
rect 184342 126529 184394 126535
rect 184342 126471 184394 126477
rect 184354 126059 184382 126471
rect 184340 126050 184396 126059
rect 184340 125985 184396 125994
rect 184450 125467 184478 126545
rect 184436 125458 184492 125467
rect 184436 125393 184492 125402
rect 184546 124579 184574 126619
rect 184532 124570 184588 124579
rect 184532 124505 184588 124514
rect 184630 123865 184682 123871
rect 184340 123830 184396 123839
rect 184630 123807 184682 123813
rect 184340 123765 184396 123774
rect 184438 123791 184490 123797
rect 184354 123723 184382 123765
rect 184438 123733 184490 123739
rect 184342 123717 184394 123723
rect 184342 123659 184394 123665
rect 184450 123099 184478 123733
rect 184534 123643 184586 123649
rect 184534 123585 184586 123591
rect 184436 123090 184492 123099
rect 184436 123025 184492 123034
rect 184546 121619 184574 123585
rect 184642 122211 184670 123807
rect 184628 122202 184684 122211
rect 184628 122137 184684 122146
rect 184532 121610 184588 121619
rect 184532 121545 184588 121554
rect 184438 120979 184490 120985
rect 184438 120921 184490 120927
rect 184342 120757 184394 120763
rect 184450 120731 184478 120921
rect 184534 120905 184586 120911
rect 184534 120847 184586 120853
rect 184342 120699 184394 120705
rect 184436 120722 184492 120731
rect 184354 119251 184382 120699
rect 184436 120657 184492 120666
rect 184546 120139 184574 120847
rect 184630 120831 184682 120837
rect 184630 120773 184682 120779
rect 184532 120130 184588 120139
rect 184532 120065 184588 120074
rect 184340 119242 184396 119251
rect 184340 119177 184396 119186
rect 184642 118659 184670 120773
rect 184628 118650 184684 118659
rect 184628 118585 184684 118594
rect 184630 118093 184682 118099
rect 184630 118035 184682 118041
rect 184534 118019 184586 118025
rect 184534 117961 184586 117967
rect 184438 117945 184490 117951
rect 184438 117887 184490 117893
rect 184342 117871 184394 117877
rect 184342 117813 184394 117819
rect 184354 117771 184382 117813
rect 184340 117762 184396 117771
rect 184340 117697 184396 117706
rect 184450 117031 184478 117887
rect 184436 117022 184492 117031
rect 184436 116957 184492 116966
rect 184546 116291 184574 117961
rect 184532 116282 184588 116291
rect 184532 116217 184588 116226
rect 184642 115403 184670 118035
rect 184628 115394 184684 115403
rect 184628 115329 184684 115338
rect 184630 115207 184682 115213
rect 184630 115149 184682 115155
rect 184438 115133 184490 115139
rect 184438 115075 184490 115081
rect 184342 115059 184394 115065
rect 184342 115001 184394 115007
rect 184354 114811 184382 115001
rect 184340 114802 184396 114811
rect 184340 114737 184396 114746
rect 184450 113923 184478 115075
rect 184534 114985 184586 114991
rect 184534 114927 184586 114933
rect 184436 113914 184492 113923
rect 184436 113849 184492 113858
rect 184546 112443 184574 114927
rect 184642 113183 184670 115149
rect 184726 113949 184778 113955
rect 184726 113891 184778 113897
rect 184628 113174 184684 113183
rect 184628 113109 184684 113118
rect 184532 112434 184588 112443
rect 184532 112369 184588 112378
rect 184342 112321 184394 112327
rect 184342 112263 184394 112269
rect 184354 111703 184382 112263
rect 184534 112247 184586 112253
rect 184534 112189 184586 112195
rect 184340 111694 184396 111703
rect 184340 111629 184396 111638
rect 184546 110963 184574 112189
rect 184532 110954 184588 110963
rect 184532 110889 184588 110898
rect 184342 109435 184394 109441
rect 184342 109377 184394 109383
rect 184354 107115 184382 109377
rect 184438 109287 184490 109293
rect 184438 109229 184490 109235
rect 184450 107855 184478 109229
rect 184630 108029 184682 108035
rect 184630 107971 184682 107977
rect 184436 107846 184492 107855
rect 184436 107781 184492 107790
rect 184340 107106 184396 107115
rect 184340 107041 184396 107050
rect 182902 106549 182954 106555
rect 182902 106491 182954 106497
rect 184534 106475 184586 106481
rect 184534 106417 184586 106423
rect 184342 106401 184394 106407
rect 184342 106343 184394 106349
rect 184354 105635 184382 106343
rect 184438 106327 184490 106333
rect 184438 106269 184490 106275
rect 184340 105626 184396 105635
rect 184340 105561 184396 105570
rect 184450 104007 184478 106269
rect 184546 104895 184574 106417
rect 184532 104886 184588 104895
rect 184532 104821 184588 104830
rect 184436 103998 184492 104007
rect 184436 103933 184492 103942
rect 184534 103663 184586 103669
rect 184534 103605 184586 103611
rect 184342 103589 184394 103595
rect 184342 103531 184394 103537
rect 184354 103415 184382 103531
rect 184438 103515 184490 103521
rect 184438 103457 184490 103463
rect 184340 103406 184396 103415
rect 184340 103341 184396 103350
rect 184450 101935 184478 103457
rect 184436 101926 184492 101935
rect 184436 101861 184492 101870
rect 184546 101047 184574 103605
rect 184532 101038 184588 101047
rect 184532 100973 184588 100982
rect 184534 100777 184586 100783
rect 184534 100719 184586 100725
rect 184438 100703 184490 100709
rect 184438 100645 184490 100651
rect 184342 100629 184394 100635
rect 184342 100571 184394 100577
rect 184354 100307 184382 100571
rect 184340 100298 184396 100307
rect 184340 100233 184396 100242
rect 184450 99567 184478 100645
rect 184436 99558 184492 99567
rect 184436 99493 184492 99502
rect 184546 98679 184574 100719
rect 184532 98670 184588 98679
rect 184532 98605 184588 98614
rect 184642 98087 184670 107971
rect 184738 102527 184766 113891
rect 185698 110223 185726 136757
rect 185794 135975 185822 155506
rect 185986 136863 186014 182933
rect 186166 182917 186218 182923
rect 186166 182859 186218 182865
rect 186070 174259 186122 174265
rect 186070 174201 186122 174207
rect 185972 136854 186028 136863
rect 185972 136789 186028 136798
rect 185780 135966 185836 135975
rect 185780 135901 185836 135910
rect 186082 135374 186110 174201
rect 186178 137455 186206 182859
rect 186274 182447 186302 205873
rect 187234 199171 187262 266405
rect 192418 263810 192446 269249
rect 192598 269217 192650 269223
rect 192610 263824 192638 269217
rect 192994 268245 193022 271881
rect 193076 269610 193132 269619
rect 193076 269545 193132 269554
rect 192982 268239 193034 268245
rect 192982 268181 193034 268187
rect 193090 263824 193118 269545
rect 192610 263796 192864 263824
rect 193090 263796 193344 263824
rect 193762 263810 193790 272061
rect 194228 269462 194284 269471
rect 194228 269397 194284 269406
rect 194242 263810 194270 269397
rect 194434 263824 194462 272209
rect 194722 272167 194750 278018
rect 195670 272235 195722 272241
rect 195670 272177 195722 272183
rect 194710 272161 194762 272167
rect 194710 272103 194762 272109
rect 194998 269349 195050 269355
rect 194998 269291 195050 269297
rect 195010 263824 195038 269291
rect 194434 263796 194736 263824
rect 195010 263796 195264 263824
rect 195682 263810 195710 272177
rect 195874 271945 195902 278018
rect 196628 272422 196684 272431
rect 196628 272357 196684 272366
rect 195862 271939 195914 271945
rect 195862 271881 195914 271887
rect 196148 269758 196204 269767
rect 196148 269693 196204 269702
rect 196162 263810 196190 269693
rect 196642 263810 196670 272357
rect 196822 269497 196874 269503
rect 196822 269439 196874 269445
rect 196834 263824 196862 269439
rect 197122 269281 197150 278018
rect 198274 272241 198302 278018
rect 199220 272570 199276 272579
rect 199220 272505 199276 272514
rect 199126 272383 199178 272389
rect 199126 272325 199178 272331
rect 198262 272235 198314 272241
rect 198262 272177 198314 272183
rect 198646 271717 198698 271723
rect 198646 271659 198698 271665
rect 198550 271125 198602 271131
rect 198550 271067 198602 271073
rect 198070 269645 198122 269651
rect 198070 269587 198122 269593
rect 197398 269423 197450 269429
rect 197398 269365 197450 269371
rect 197110 269275 197162 269281
rect 197110 269217 197162 269223
rect 197410 263824 197438 269365
rect 196834 263796 197088 263824
rect 197410 263796 197664 263824
rect 198082 263810 198110 269587
rect 198562 263810 198590 271067
rect 198658 269651 198686 271659
rect 198646 269645 198698 269651
rect 198646 269587 198698 269593
rect 199030 269571 199082 269577
rect 199030 269513 199082 269519
rect 199042 263810 199070 269513
rect 199138 267875 199166 272325
rect 199126 267869 199178 267875
rect 199126 267811 199178 267817
rect 199234 263824 199262 272505
rect 199426 271723 199454 278018
rect 200468 272718 200524 272727
rect 200468 272653 200524 272662
rect 199414 271717 199466 271723
rect 199414 271659 199466 271665
rect 199702 269719 199754 269725
rect 199702 269661 199754 269667
rect 199714 263824 199742 269661
rect 199234 263796 199488 263824
rect 199714 263796 199968 263824
rect 200482 263810 200510 272653
rect 200674 269355 200702 278018
rect 201622 272309 201674 272315
rect 201622 272251 201674 272257
rect 201526 271495 201578 271501
rect 201526 271437 201578 271443
rect 200950 269793 201002 269799
rect 200950 269735 201002 269741
rect 200662 269349 200714 269355
rect 200662 269291 200714 269297
rect 200962 263810 200990 269735
rect 201538 269725 201566 271437
rect 201526 269719 201578 269725
rect 201526 269661 201578 269667
rect 201142 268313 201194 268319
rect 201142 268255 201194 268261
rect 201154 263824 201182 268255
rect 201634 263824 201662 272251
rect 201826 271501 201854 278018
rect 201814 271495 201866 271501
rect 201814 271437 201866 271443
rect 202870 269941 202922 269947
rect 202870 269883 202922 269889
rect 202294 267869 202346 267875
rect 202294 267811 202346 267817
rect 201154 263796 201408 263824
rect 201634 263796 201888 263824
rect 202306 263810 202334 267811
rect 202882 263810 202910 269883
rect 202978 269503 203006 278018
rect 204022 272531 204074 272537
rect 204022 272473 204074 272479
rect 203542 272457 203594 272463
rect 203542 272399 203594 272405
rect 203350 270089 203402 270095
rect 203350 270031 203402 270037
rect 202966 269497 203018 269503
rect 202966 269439 203018 269445
rect 203362 263810 203390 270031
rect 203554 263824 203582 272399
rect 204034 263824 204062 272473
rect 204130 269429 204158 278018
rect 205174 271569 205226 271575
rect 205174 271511 205226 271517
rect 204694 270015 204746 270021
rect 204694 269957 204746 269963
rect 204118 269423 204170 269429
rect 204118 269365 204170 269371
rect 203554 263796 203808 263824
rect 204034 263796 204288 263824
rect 204706 263810 204734 269957
rect 205186 269947 205214 271511
rect 205378 271131 205406 278018
rect 206038 272679 206090 272685
rect 206038 272621 206090 272627
rect 205750 272605 205802 272611
rect 205750 272547 205802 272553
rect 205366 271125 205418 271131
rect 205366 271067 205418 271073
rect 205270 270163 205322 270169
rect 205270 270105 205322 270111
rect 205174 269941 205226 269947
rect 205174 269883 205226 269889
rect 205282 263810 205310 270105
rect 205762 263810 205790 272547
rect 205942 271347 205994 271353
rect 205942 271289 205994 271295
rect 205846 271199 205898 271205
rect 205846 271141 205898 271147
rect 205858 269799 205886 271141
rect 205954 269873 205982 271289
rect 205942 269867 205994 269873
rect 205942 269809 205994 269815
rect 205846 269793 205898 269799
rect 205846 269735 205898 269741
rect 206050 263824 206078 272621
rect 206422 270237 206474 270243
rect 206422 270179 206474 270185
rect 206434 263824 206462 270179
rect 206530 269577 206558 278018
rect 207478 273567 207530 273573
rect 207478 273509 207530 273515
rect 207382 273271 207434 273277
rect 207382 273213 207434 273219
rect 207286 273049 207338 273055
rect 207286 272991 207338 272997
rect 207094 272827 207146 272833
rect 207094 272769 207146 272775
rect 206518 269571 206570 269577
rect 206518 269513 206570 269519
rect 206050 263796 206208 263824
rect 206434 263796 206688 263824
rect 207106 263810 207134 272769
rect 207298 267949 207326 272991
rect 207394 268097 207422 273213
rect 207490 268319 207518 273509
rect 207682 272389 207710 278018
rect 207862 272753 207914 272759
rect 207862 272695 207914 272701
rect 207670 272383 207722 272389
rect 207670 272325 207722 272331
rect 207574 270311 207626 270317
rect 207574 270253 207626 270259
rect 207478 268313 207530 268319
rect 207478 268255 207530 268261
rect 207382 268091 207434 268097
rect 207382 268033 207434 268039
rect 207286 267943 207338 267949
rect 207286 267885 207338 267891
rect 207586 263810 207614 270253
rect 207874 263824 207902 272695
rect 208930 272537 208958 278018
rect 209590 273419 209642 273425
rect 209590 273361 209642 273367
rect 209014 272901 209066 272907
rect 209014 272843 209066 272849
rect 208918 272531 208970 272537
rect 208918 272473 208970 272479
rect 208342 270385 208394 270391
rect 208342 270327 208394 270333
rect 208354 263824 208382 270327
rect 207874 263796 208128 263824
rect 208354 263796 208608 263824
rect 209026 263810 209054 272843
rect 209602 268139 209630 273361
rect 209878 273345 209930 273351
rect 209878 273287 209930 273293
rect 209686 273197 209738 273203
rect 209686 273139 209738 273145
rect 209588 268130 209644 268139
rect 209588 268065 209644 268074
rect 209494 267943 209546 267949
rect 209494 267885 209546 267891
rect 209506 263810 209534 267885
rect 209698 267875 209726 273139
rect 209890 268023 209918 273287
rect 209974 273123 210026 273129
rect 209974 273065 210026 273071
rect 209878 268017 209930 268023
rect 209878 267959 209930 267965
rect 209686 267869 209738 267875
rect 209686 267811 209738 267817
rect 209986 263810 210014 273065
rect 210082 272463 210110 278018
rect 210166 272975 210218 272981
rect 210166 272917 210218 272923
rect 210070 272457 210122 272463
rect 210070 272399 210122 272405
rect 210178 267968 210206 272917
rect 211234 272611 211262 278018
rect 212482 272759 212510 278018
rect 212470 272753 212522 272759
rect 212470 272695 212522 272701
rect 213634 272685 213662 278018
rect 214786 272833 214814 278018
rect 216034 272981 216062 278018
rect 217186 273055 217214 278018
rect 217174 273049 217226 273055
rect 217174 272991 217226 272997
rect 216022 272975 216074 272981
rect 216022 272917 216074 272923
rect 218338 272907 218366 278018
rect 219586 273351 219614 278018
rect 219574 273345 219626 273351
rect 219574 273287 219626 273293
rect 220738 273129 220766 278018
rect 221494 273493 221546 273499
rect 221494 273435 221546 273441
rect 220726 273123 220778 273129
rect 220726 273065 220778 273071
rect 218326 272901 218378 272907
rect 218326 272843 218378 272849
rect 214774 272827 214826 272833
rect 214774 272769 214826 272775
rect 213622 272679 213674 272685
rect 213622 272621 213674 272627
rect 211222 272605 211274 272611
rect 211222 272547 211274 272553
rect 210646 272087 210698 272093
rect 210646 272029 210698 272035
rect 210550 272013 210602 272019
rect 210550 271955 210602 271961
rect 210454 271643 210506 271649
rect 210454 271585 210506 271591
rect 210358 271421 210410 271427
rect 210358 271363 210410 271369
rect 210262 271273 210314 271279
rect 210262 271215 210314 271221
rect 210274 270169 210302 271215
rect 210262 270163 210314 270169
rect 210262 270105 210314 270111
rect 210370 270095 210398 271363
rect 210358 270089 210410 270095
rect 210358 270031 210410 270037
rect 210466 270021 210494 271585
rect 210562 270243 210590 271955
rect 210550 270237 210602 270243
rect 210550 270179 210602 270185
rect 210454 270015 210506 270021
rect 210454 269957 210506 269963
rect 210178 267940 210302 267968
rect 210658 267949 210686 272029
rect 214966 270681 215018 270687
rect 214966 270623 215018 270629
rect 212662 270607 212714 270613
rect 212662 270549 212714 270555
rect 211894 270459 211946 270465
rect 211894 270401 211946 270407
rect 211030 268313 211082 268319
rect 210850 268261 211030 268264
rect 210850 268255 211082 268261
rect 210850 268245 211070 268255
rect 210838 268239 211070 268245
rect 210890 268236 211070 268239
rect 210838 268181 210890 268187
rect 210742 268165 210794 268171
rect 210742 268107 210794 268113
rect 210274 263824 210302 267940
rect 210646 267943 210698 267949
rect 210646 267885 210698 267891
rect 210754 263824 210782 268107
rect 211414 267869 211466 267875
rect 211414 267811 211466 267817
rect 210274 263796 210528 263824
rect 210754 263796 211008 263824
rect 211426 263810 211454 267811
rect 211906 263810 211934 270401
rect 212374 268017 212426 268023
rect 212374 267959 212426 267965
rect 212386 263810 212414 267959
rect 212674 263824 212702 270549
rect 213814 270533 213866 270539
rect 213814 270475 213866 270481
rect 213332 269906 213388 269915
rect 213332 269841 213388 269850
rect 212674 263796 212928 263824
rect 213346 263810 213374 269841
rect 213826 263810 213854 270475
rect 214486 269201 214538 269207
rect 214486 269143 214538 269149
rect 214292 268130 214348 268139
rect 214292 268065 214348 268074
rect 214306 263810 214334 268065
rect 214498 263824 214526 269143
rect 214978 263824 215006 270623
rect 220534 269645 220586 269651
rect 220534 269587 220586 269593
rect 216694 269127 216746 269133
rect 216694 269069 216746 269075
rect 216214 269053 216266 269059
rect 216214 268995 216266 269001
rect 215734 268979 215786 268985
rect 215734 268921 215786 268927
rect 214498 263796 214752 263824
rect 214978 263796 215232 263824
rect 215746 263810 215774 268921
rect 216226 263810 216254 268995
rect 216706 263810 216734 269069
rect 217366 268905 217418 268911
rect 217366 268847 217418 268853
rect 216886 268091 216938 268097
rect 216886 268033 216938 268039
rect 216898 263824 216926 268033
rect 217378 263824 217406 268847
rect 218134 268831 218186 268837
rect 218134 268773 218186 268779
rect 216898 263796 217152 263824
rect 217378 263796 217632 263824
rect 218146 263810 218174 268773
rect 219286 268757 219338 268763
rect 219286 268699 219338 268705
rect 218614 268313 218666 268319
rect 218614 268255 218666 268261
rect 218626 263810 218654 268255
rect 218902 268165 218954 268171
rect 218902 268107 218954 268113
rect 218914 263824 218942 268107
rect 219298 263824 219326 268699
rect 219958 268683 220010 268689
rect 219958 268625 220010 268631
rect 218914 263796 219072 263824
rect 219298 263796 219552 263824
rect 219970 263810 219998 268625
rect 220546 263810 220574 269587
rect 221206 268609 221258 268615
rect 221206 268551 221258 268557
rect 221014 267943 221066 267949
rect 221014 267885 221066 267891
rect 221026 263810 221054 267885
rect 221218 263824 221246 268551
rect 221506 268319 221534 273435
rect 221686 271939 221738 271945
rect 221686 271881 221738 271887
rect 221590 271717 221642 271723
rect 221590 271659 221642 271665
rect 221494 268313 221546 268319
rect 221494 268255 221546 268261
rect 221602 268097 221630 271659
rect 221590 268091 221642 268097
rect 221590 268033 221642 268039
rect 221698 268023 221726 271881
rect 221890 271057 221918 278018
rect 221878 271051 221930 271057
rect 221878 270993 221930 270999
rect 223042 270983 223070 278018
rect 223702 271495 223754 271501
rect 223702 271437 223754 271443
rect 223030 270977 223082 270983
rect 223030 270919 223082 270925
rect 222838 270237 222890 270243
rect 222838 270179 222890 270185
rect 222358 269719 222410 269725
rect 222358 269661 222410 269667
rect 221782 268535 221834 268541
rect 221782 268477 221834 268483
rect 221686 268017 221738 268023
rect 221686 267959 221738 267965
rect 221794 263824 221822 268477
rect 221218 263796 221472 263824
rect 221794 263796 221952 263824
rect 222370 263810 222398 269661
rect 222850 263810 222878 270179
rect 223414 268461 223466 268467
rect 223414 268403 223466 268409
rect 223426 263810 223454 268403
rect 223606 268387 223658 268393
rect 223606 268329 223658 268335
rect 223618 263824 223646 268329
rect 223714 268171 223742 271437
rect 224290 270909 224318 278018
rect 224374 272235 224426 272241
rect 224374 272177 224426 272183
rect 224278 270903 224330 270909
rect 224278 270845 224330 270851
rect 224086 269941 224138 269947
rect 224086 269883 224138 269889
rect 223702 268165 223754 268171
rect 223702 268107 223754 268113
rect 224098 263824 224126 269883
rect 224386 268245 224414 272177
rect 224470 272161 224522 272167
rect 224470 272103 224522 272109
rect 224374 268239 224426 268245
rect 224374 268181 224426 268187
rect 224482 267949 224510 272103
rect 224566 271791 224618 271797
rect 224566 271733 224618 271739
rect 224470 267943 224522 267949
rect 224470 267885 224522 267891
rect 224578 267875 224606 271733
rect 225442 270835 225470 278018
rect 225430 270829 225482 270835
rect 225430 270771 225482 270777
rect 226594 270761 226622 278018
rect 227842 272241 227870 278018
rect 227830 272235 227882 272241
rect 227830 272177 227882 272183
rect 228994 272167 229022 278018
rect 230146 273499 230174 278018
rect 230134 273493 230186 273499
rect 230134 273435 230186 273441
rect 228982 272161 229034 272167
rect 228982 272103 229034 272109
rect 231394 272019 231422 278018
rect 232546 272315 232574 278018
rect 232534 272309 232586 272315
rect 232534 272251 232586 272257
rect 231382 272013 231434 272019
rect 231382 271955 231434 271961
rect 233698 271945 233726 278018
rect 234358 272531 234410 272537
rect 234358 272473 234410 272479
rect 233878 272383 233930 272389
rect 233878 272325 233930 272331
rect 233686 271939 233738 271945
rect 233686 271881 233738 271887
rect 227158 271865 227210 271871
rect 227158 271807 227210 271813
rect 226582 270755 226634 270761
rect 226582 270697 226634 270703
rect 226678 270163 226730 270169
rect 226678 270105 226730 270111
rect 225526 270089 225578 270095
rect 225526 270031 225578 270037
rect 224758 270015 224810 270021
rect 224758 269957 224810 269963
rect 224566 267869 224618 267875
rect 224566 267811 224618 267817
rect 223618 263796 223872 263824
rect 224098 263796 224352 263824
rect 224770 263810 224798 269957
rect 225238 269867 225290 269873
rect 225238 269809 225290 269815
rect 225250 263810 225278 269809
rect 225538 263824 225566 270031
rect 226006 269793 226058 269799
rect 226006 269735 226058 269741
rect 226018 263824 226046 269735
rect 225538 263796 225792 263824
rect 226018 263796 226272 263824
rect 226690 263810 226718 270105
rect 227170 263810 227198 271807
rect 232630 271125 232682 271131
rect 232630 271067 232682 271073
rect 231958 269497 232010 269503
rect 231958 269439 232010 269445
rect 230998 269349 231050 269355
rect 230998 269291 231050 269297
rect 229558 269275 229610 269281
rect 229558 269217 229610 269223
rect 227830 268313 227882 268319
rect 227830 268255 227882 268261
rect 227638 267869 227690 267875
rect 227638 267811 227690 267817
rect 227650 263810 227678 267811
rect 227842 263824 227870 268255
rect 229078 268017 229130 268023
rect 229078 267959 229130 267965
rect 228406 267943 228458 267949
rect 228406 267885 228458 267891
rect 228418 263824 228446 267885
rect 227842 263796 228096 263824
rect 228418 263796 228672 263824
rect 229090 263810 229118 267959
rect 229570 263810 229598 269217
rect 230038 268239 230090 268245
rect 230038 268181 230090 268187
rect 230050 263810 230078 268181
rect 230518 268091 230570 268097
rect 230518 268033 230570 268039
rect 230530 264120 230558 268033
rect 230482 264092 230558 264120
rect 230482 263810 230510 264092
rect 231010 263810 231038 269291
rect 231478 268165 231530 268171
rect 231478 268107 231530 268113
rect 231490 263810 231518 268107
rect 231970 263810 231998 269439
rect 232150 269423 232202 269429
rect 232150 269365 232202 269371
rect 232162 263824 232190 269365
rect 232642 263824 232670 271067
rect 233398 269571 233450 269577
rect 233398 269513 233450 269519
rect 232162 263796 232416 263824
rect 232642 263796 232896 263824
rect 233410 263810 233438 269513
rect 233890 263810 233918 272325
rect 234370 263810 234398 272473
rect 234550 272457 234602 272463
rect 234550 272399 234602 272405
rect 234562 263824 234590 272399
rect 234946 272389 234974 278018
rect 235702 272753 235754 272759
rect 235702 272695 235754 272701
rect 235030 272605 235082 272611
rect 235030 272547 235082 272553
rect 234934 272383 234986 272389
rect 234934 272325 234986 272331
rect 235042 263824 235070 272547
rect 234562 263796 234816 263824
rect 235042 263796 235296 263824
rect 235714 263810 235742 272695
rect 236098 272463 236126 278018
rect 236950 272975 237002 272981
rect 236950 272917 237002 272923
rect 236470 272827 236522 272833
rect 236470 272769 236522 272775
rect 236278 272679 236330 272685
rect 236278 272621 236330 272627
rect 236086 272457 236138 272463
rect 236086 272399 236138 272405
rect 236290 263810 236318 272621
rect 236482 263824 236510 272769
rect 236962 263824 236990 272917
rect 237250 271279 237278 278018
rect 237622 273049 237674 273055
rect 237622 272991 237674 272997
rect 237238 271273 237290 271279
rect 237238 271215 237290 271221
rect 236482 263796 236736 263824
rect 236962 263796 237216 263824
rect 237634 263810 237662 272991
rect 238102 272901 238154 272907
rect 238102 272843 238154 272849
rect 238114 263810 238142 272843
rect 238498 271205 238526 278018
rect 238678 273345 238730 273351
rect 238678 273287 238730 273293
rect 238486 271199 238538 271205
rect 238486 271141 238538 271147
rect 238690 263810 238718 273287
rect 239158 273123 239210 273129
rect 239158 273065 239210 273071
rect 239170 263824 239198 273065
rect 239350 271051 239402 271057
rect 239350 270993 239402 270999
rect 239542 271051 239594 271057
rect 239542 270993 239594 270999
rect 239136 263796 239198 263824
rect 239362 263824 239390 270993
rect 239554 270761 239582 270993
rect 239650 270761 239678 278018
rect 240802 271131 240830 278018
rect 240790 271125 240842 271131
rect 240790 271067 240842 271073
rect 241954 271057 241982 278018
rect 242902 273493 242954 273499
rect 242902 273435 242954 273441
rect 242134 272235 242186 272241
rect 242134 272177 242186 272183
rect 241270 271051 241322 271057
rect 241270 270993 241322 270999
rect 241942 271051 241994 271057
rect 241942 270993 241994 270999
rect 240022 270977 240074 270983
rect 240022 270919 240074 270925
rect 239542 270755 239594 270761
rect 239542 270697 239594 270703
rect 239638 270755 239690 270761
rect 239638 270697 239690 270703
rect 239362 263796 239616 263824
rect 240034 263810 240062 270919
rect 240502 270903 240554 270909
rect 240502 270845 240554 270851
rect 240514 263810 240542 270845
rect 241078 270829 241130 270835
rect 241078 270771 241130 270777
rect 241090 263810 241118 270771
rect 241282 263824 241310 270993
rect 242146 263824 242174 272177
rect 242422 272161 242474 272167
rect 242422 272103 242474 272109
rect 241282 263796 241536 263824
rect 242016 263796 242174 263824
rect 242434 263810 242462 272103
rect 242914 263810 242942 273435
rect 243094 272013 243146 272019
rect 243094 271955 243146 271961
rect 243106 263824 243134 271955
rect 243202 270983 243230 278018
rect 243670 272309 243722 272315
rect 243670 272251 243722 272257
rect 243190 270977 243242 270983
rect 243190 270919 243242 270925
rect 243682 263824 243710 272251
rect 244054 271939 244106 271945
rect 244054 271881 244106 271887
rect 244066 263824 244094 271881
rect 244354 270909 244382 278018
rect 245302 272457 245354 272463
rect 245302 272399 245354 272405
rect 244822 272383 244874 272389
rect 244822 272325 244874 272331
rect 244342 270903 244394 270909
rect 244342 270845 244394 270851
rect 243106 263796 243360 263824
rect 243682 263796 243936 263824
rect 244066 263796 244368 263824
rect 244834 263810 244862 272325
rect 245314 263810 245342 272399
rect 245506 270835 245534 278018
rect 245590 271273 245642 271279
rect 245590 271215 245642 271221
rect 245494 270829 245546 270835
rect 245494 270771 245546 270777
rect 245602 263824 245630 271215
rect 246070 271199 246122 271205
rect 246070 271141 246122 271147
rect 246082 263824 246110 271141
rect 246754 270761 246782 278018
rect 247222 271125 247274 271131
rect 247222 271067 247274 271073
rect 246454 270755 246506 270761
rect 246454 270697 246506 270703
rect 246742 270755 246794 270761
rect 246742 270697 246794 270703
rect 246466 263824 246494 270697
rect 245602 263796 245760 263824
rect 246082 263796 246336 263824
rect 246466 263796 246768 263824
rect 247234 263810 247262 271067
rect 247702 271051 247754 271057
rect 247702 270993 247754 270999
rect 247714 263810 247742 270993
rect 247906 268393 247934 278018
rect 247990 270977 248042 270983
rect 247990 270919 248042 270925
rect 247894 268387 247946 268393
rect 247894 268329 247946 268335
rect 248002 263824 248030 270919
rect 248662 270903 248714 270909
rect 248662 270845 248714 270851
rect 248002 263796 248160 263824
rect 248674 263810 248702 270845
rect 249058 269651 249086 278018
rect 250320 278004 250526 278032
rect 249142 270829 249194 270835
rect 249142 270771 249194 270777
rect 250498 270780 250526 278004
rect 249046 269645 249098 269651
rect 249046 269587 249098 269593
rect 249154 263810 249182 270771
rect 249622 270755 249674 270761
rect 250498 270752 250718 270780
rect 249622 270697 249674 270703
rect 249634 263810 249662 270697
rect 250294 269645 250346 269651
rect 250294 269587 250346 269593
rect 249814 268387 249866 268393
rect 249814 268329 249866 268335
rect 249826 263824 249854 268329
rect 250306 263824 250334 269587
rect 250690 263824 250718 270752
rect 251458 263824 251486 278018
rect 252322 278004 252624 278032
rect 252322 263824 252350 278004
rect 253366 269127 253418 269133
rect 253366 269069 253418 269075
rect 253174 268979 253226 268985
rect 253174 268921 253226 268927
rect 252694 268091 252746 268097
rect 252694 268033 252746 268039
rect 252706 263824 252734 268033
rect 253186 263824 253214 268921
rect 249826 263796 250080 263824
rect 250306 263796 250560 263824
rect 250690 263796 250992 263824
rect 251458 263796 251568 263824
rect 252048 263796 252350 263824
rect 252480 263796 252734 263824
rect 252960 263796 253214 263824
rect 253378 263810 253406 269069
rect 253762 268097 253790 278018
rect 253942 270459 253994 270465
rect 253942 270401 253994 270407
rect 253750 268091 253802 268097
rect 253750 268033 253802 268039
rect 253954 263810 253982 270401
rect 255010 268985 255038 278018
rect 255286 270311 255338 270317
rect 255286 270253 255338 270259
rect 254998 268979 255050 268985
rect 254998 268921 255050 268927
rect 254614 268683 254666 268689
rect 254614 268625 254666 268631
rect 254626 263824 254654 268625
rect 255094 268387 255146 268393
rect 255094 268329 255146 268335
rect 255106 263824 255134 268329
rect 254400 263796 254654 263824
rect 254880 263796 255134 263824
rect 255298 263810 255326 270253
rect 255766 269867 255818 269873
rect 255766 269809 255818 269815
rect 255778 263810 255806 269809
rect 256162 269133 256190 278018
rect 257314 270465 257342 278018
rect 257302 270459 257354 270465
rect 257302 270401 257354 270407
rect 256246 269941 256298 269947
rect 256246 269883 256298 269889
rect 256150 269127 256202 269133
rect 256150 269069 256202 269075
rect 256258 263810 256286 269883
rect 257686 269645 257738 269651
rect 257686 269587 257738 269593
rect 257494 269275 257546 269281
rect 257494 269217 257546 269223
rect 257014 268239 257066 268245
rect 257014 268181 257066 268187
rect 257026 263824 257054 268181
rect 257506 263824 257534 269217
rect 256800 263796 257054 263824
rect 257280 263796 257534 263824
rect 257698 263810 257726 269587
rect 258166 268831 258218 268837
rect 258166 268773 258218 268779
rect 258178 263810 258206 268773
rect 258562 268689 258590 278018
rect 258646 269349 258698 269355
rect 258646 269291 258698 269297
rect 258550 268683 258602 268689
rect 258550 268625 258602 268631
rect 258658 263810 258686 269291
rect 259414 269127 259466 269133
rect 259414 269069 259466 269075
rect 259426 263824 259454 269069
rect 259714 268393 259742 278018
rect 260866 270317 260894 278018
rect 260854 270311 260906 270317
rect 260854 270253 260906 270259
rect 262114 269873 262142 278018
rect 262486 270385 262538 270391
rect 262486 270327 262538 270333
rect 262102 269867 262154 269873
rect 262102 269809 262154 269815
rect 259894 269719 259946 269725
rect 259894 269661 259946 269667
rect 259702 268387 259754 268393
rect 259702 268329 259754 268335
rect 259906 263824 259934 269661
rect 260086 269497 260138 269503
rect 260086 269439 260138 269445
rect 259200 263796 259454 263824
rect 259680 263796 259934 263824
rect 260098 263810 260126 269439
rect 262006 269201 262058 269207
rect 262006 269143 262058 269149
rect 261814 269053 261866 269059
rect 261814 268995 261866 269001
rect 261238 268979 261290 268985
rect 261238 268921 261290 268927
rect 260566 268683 260618 268689
rect 260566 268625 260618 268631
rect 260578 263810 260606 268625
rect 261250 263824 261278 268921
rect 261826 263824 261854 268995
rect 261024 263796 261278 263824
rect 261600 263796 261854 263824
rect 262018 263810 262046 269143
rect 262498 263810 262526 270327
rect 263266 269947 263294 278018
rect 263254 269941 263306 269947
rect 263254 269883 263306 269889
rect 264118 268905 264170 268911
rect 264118 268847 264170 268853
rect 263638 268535 263690 268541
rect 263638 268477 263690 268483
rect 262966 268387 263018 268393
rect 262966 268329 263018 268335
rect 262978 263810 263006 268329
rect 263650 263824 263678 268477
rect 264130 263824 264158 268847
rect 264418 268245 264446 278018
rect 264694 270533 264746 270539
rect 264694 270475 264746 270481
rect 264406 268239 264458 268245
rect 264406 268181 264458 268187
rect 264706 263824 264734 270475
rect 264886 270459 264938 270465
rect 264886 270401 264938 270407
rect 263424 263796 263678 263824
rect 263904 263796 264158 263824
rect 264432 263796 264734 263824
rect 264898 263810 264926 270401
rect 265366 270237 265418 270243
rect 265366 270179 265418 270185
rect 265378 263810 265406 270179
rect 265666 269281 265694 278018
rect 266038 270311 266090 270317
rect 266038 270253 266090 270259
rect 265654 269275 265706 269281
rect 265654 269217 265706 269223
rect 266050 263824 266078 270253
rect 266518 270163 266570 270169
rect 266518 270105 266570 270111
rect 266530 263824 266558 270105
rect 266818 269651 266846 278018
rect 267286 270089 267338 270095
rect 267286 270031 267338 270037
rect 267094 270015 267146 270021
rect 267094 269957 267146 269963
rect 266806 269645 266858 269651
rect 266806 269587 266858 269593
rect 267106 263824 267134 269957
rect 265824 263796 266078 263824
rect 266304 263796 266558 263824
rect 266832 263796 267134 263824
rect 267298 263810 267326 270031
rect 267766 269941 267818 269947
rect 267766 269883 267818 269889
rect 267778 263824 267806 269883
rect 267970 268837 267998 278018
rect 269122 269355 269150 278018
rect 270262 272605 270314 272611
rect 270262 272547 270314 272553
rect 269206 269867 269258 269873
rect 269206 269809 269258 269815
rect 269110 269349 269162 269355
rect 269110 269291 269162 269297
rect 268630 269275 268682 269281
rect 268630 269217 268682 269223
rect 267958 268831 268010 268837
rect 267958 268773 268010 268779
rect 268438 268757 268490 268763
rect 268438 268699 268490 268705
rect 268450 263824 268478 268699
rect 267744 263796 267806 263824
rect 268224 263796 268478 263824
rect 268642 263810 268670 269217
rect 269218 263810 269246 269809
rect 269686 269645 269738 269651
rect 269686 269587 269738 269593
rect 269698 263810 269726 269587
rect 270274 263824 270302 272547
rect 270370 269133 270398 278018
rect 271030 272975 271082 272981
rect 271030 272917 271082 272923
rect 270550 272531 270602 272537
rect 270550 272473 270602 272479
rect 270358 269127 270410 269133
rect 270358 269069 270410 269075
rect 270144 263796 270302 263824
rect 270562 263824 270590 272473
rect 270562 263796 270624 263824
rect 271042 263810 271070 272917
rect 271522 269725 271550 278018
rect 272278 271939 272330 271945
rect 272278 271881 272330 271887
rect 271510 269719 271562 269725
rect 271510 269661 271562 269667
rect 271606 269719 271658 269725
rect 271606 269661 271658 269667
rect 271510 269571 271562 269577
rect 271510 269513 271562 269519
rect 271522 263810 271550 269513
rect 271618 269281 271646 269661
rect 271606 269275 271658 269281
rect 271606 269217 271658 269223
rect 272290 263824 272318 271881
rect 272674 269503 272702 278018
rect 272758 272383 272810 272389
rect 272758 272325 272810 272331
rect 272662 269497 272714 269503
rect 272662 269439 272714 269445
rect 272770 263824 272798 272325
rect 273430 272235 273482 272241
rect 273430 272177 273482 272183
rect 272950 269497 273002 269503
rect 272950 269439 273002 269445
rect 272064 263796 272318 263824
rect 272544 263796 272798 263824
rect 272962 263810 272990 269439
rect 273442 263810 273470 272177
rect 273922 268689 273950 278018
rect 274198 272457 274250 272463
rect 274198 272399 274250 272405
rect 273910 268683 273962 268689
rect 273910 268625 273962 268631
rect 274210 263824 274238 272399
rect 274678 269423 274730 269429
rect 274678 269365 274730 269371
rect 274690 263824 274718 269365
rect 275074 268985 275102 278018
rect 275350 273493 275402 273499
rect 275350 273435 275402 273441
rect 275158 272309 275210 272315
rect 275158 272251 275210 272257
rect 275062 268979 275114 268985
rect 275062 268921 275114 268927
rect 275170 263824 275198 272251
rect 273936 263796 274238 263824
rect 274464 263796 274718 263824
rect 274944 263796 275198 263824
rect 275362 263810 275390 273435
rect 275830 269275 275882 269281
rect 275830 269217 275882 269223
rect 275842 263810 275870 269217
rect 276226 269059 276254 278018
rect 277078 273419 277130 273425
rect 277078 273361 277130 273367
rect 276310 272161 276362 272167
rect 276310 272103 276362 272109
rect 276214 269053 276266 269059
rect 276214 268995 276266 269001
rect 276322 263810 276350 272103
rect 276406 270459 276458 270465
rect 276406 270401 276458 270407
rect 276418 270243 276446 270401
rect 276406 270237 276458 270243
rect 276406 270179 276458 270185
rect 277090 263824 277118 273361
rect 277474 269207 277502 278018
rect 277750 273567 277802 273573
rect 277750 273509 277802 273515
rect 277462 269201 277514 269207
rect 277462 269143 277514 269149
rect 277558 269201 277610 269207
rect 277558 269143 277610 269149
rect 277570 263824 277598 269143
rect 276864 263796 277118 263824
rect 277344 263796 277598 263824
rect 277762 263810 277790 273509
rect 278230 273271 278282 273277
rect 278230 273213 278282 273219
rect 278242 263810 278270 273213
rect 278626 270391 278654 278018
rect 279670 273345 279722 273351
rect 279670 273287 279722 273293
rect 279286 270459 279338 270465
rect 279286 270401 279338 270407
rect 278614 270385 278666 270391
rect 278614 270327 278666 270333
rect 278902 269349 278954 269355
rect 278902 269291 278954 269297
rect 278914 263824 278942 269291
rect 279298 263824 279326 270401
rect 278688 263796 278942 263824
rect 279168 263796 279326 263824
rect 279682 263810 279710 273287
rect 279778 268393 279806 278018
rect 280150 270681 280202 270687
rect 280150 270623 280202 270629
rect 279766 268387 279818 268393
rect 279766 268329 279818 268335
rect 280162 263810 280190 270623
rect 280630 270607 280682 270613
rect 280630 270549 280682 270555
rect 280642 263810 280670 270549
rect 281026 268541 281054 278018
rect 281782 274899 281834 274905
rect 281782 274841 281834 274847
rect 281302 269053 281354 269059
rect 281302 268995 281354 269001
rect 281014 268535 281066 268541
rect 281014 268477 281066 268483
rect 281314 263824 281342 268995
rect 281794 263824 281822 274841
rect 282070 268979 282122 268985
rect 282070 268921 282122 268927
rect 281088 263796 281342 263824
rect 281568 263796 281822 263824
rect 282082 263810 282110 268921
rect 282178 268911 282206 278018
rect 283030 274973 283082 274979
rect 283030 274915 283082 274921
rect 282166 268905 282218 268911
rect 282166 268847 282218 268853
rect 282550 267869 282602 267875
rect 282550 267811 282602 267817
rect 282562 263810 282590 267811
rect 283042 263810 283070 274915
rect 283330 270539 283358 278018
rect 284470 276453 284522 276459
rect 284470 276395 284522 276401
rect 283318 270533 283370 270539
rect 283318 270475 283370 270481
rect 283702 270459 283754 270465
rect 283702 270401 283754 270407
rect 283714 263824 283742 270401
rect 284182 270385 284234 270391
rect 284182 270327 284234 270333
rect 284194 263824 284222 270327
rect 283488 263796 283742 263824
rect 283968 263796 284222 263824
rect 284482 263810 284510 276395
rect 284578 270243 284606 278018
rect 285622 273197 285674 273203
rect 285622 273139 285674 273145
rect 284950 273049 285002 273055
rect 284950 272991 285002 272997
rect 284566 270237 284618 270243
rect 284566 270179 284618 270185
rect 284962 263810 284990 272991
rect 285634 263824 285662 273139
rect 285730 270169 285758 278018
rect 286102 276379 286154 276385
rect 286102 276321 286154 276327
rect 285718 270163 285770 270169
rect 285718 270105 285770 270111
rect 286114 263824 286142 276321
rect 286774 273123 286826 273129
rect 286774 273065 286826 273071
rect 286294 270237 286346 270243
rect 286294 270179 286346 270185
rect 285408 263796 285662 263824
rect 285888 263796 286142 263824
rect 286306 263810 286334 270179
rect 286786 263810 286814 273065
rect 286882 270317 286910 278018
rect 287350 276231 287402 276237
rect 287350 276173 287402 276179
rect 286870 270311 286922 270317
rect 286870 270253 286922 270259
rect 287362 263810 287390 276173
rect 287926 270163 287978 270169
rect 287926 270105 287978 270111
rect 287938 263824 287966 270105
rect 288034 270095 288062 278018
rect 288694 276305 288746 276311
rect 288694 276247 288746 276253
rect 288502 270237 288554 270243
rect 288502 270179 288554 270185
rect 288022 270089 288074 270095
rect 288022 270031 288074 270037
rect 288514 263824 288542 270179
rect 287808 263796 287966 263824
rect 288288 263796 288542 263824
rect 288706 263810 288734 276247
rect 289282 269947 289310 278018
rect 290326 276083 290378 276089
rect 290326 276025 290378 276031
rect 289942 272901 289994 272907
rect 289942 272843 289994 272849
rect 289270 269941 289322 269947
rect 289270 269883 289322 269889
rect 289174 268831 289226 268837
rect 289174 268773 289226 268779
rect 289186 263810 289214 268773
rect 289954 263824 289982 272843
rect 290338 263824 290366 276025
rect 290434 270021 290462 278018
rect 290614 270089 290666 270095
rect 290614 270031 290666 270037
rect 290422 270015 290474 270021
rect 290422 269957 290474 269963
rect 289728 263796 289982 263824
rect 290208 263796 290366 263824
rect 290626 263810 290654 270031
rect 291094 270015 291146 270021
rect 291094 269957 291146 269963
rect 291106 263810 291134 269957
rect 291586 269873 291614 278018
rect 291862 276157 291914 276163
rect 291862 276099 291914 276105
rect 291574 269867 291626 269873
rect 291574 269809 291626 269815
rect 291874 263824 291902 276099
rect 292246 272827 292298 272833
rect 292246 272769 292298 272775
rect 292258 263824 292286 272769
rect 292726 272753 292778 272759
rect 292726 272695 292778 272701
rect 292738 263824 292766 272695
rect 292834 268763 292862 278018
rect 293794 278004 294000 278032
rect 293014 276009 293066 276015
rect 293014 275951 293066 275957
rect 292822 268757 292874 268763
rect 292822 268699 292874 268705
rect 291600 263796 291902 263824
rect 292032 263796 292286 263824
rect 292608 263796 292766 263824
rect 293026 263810 293054 275951
rect 293494 269867 293546 269873
rect 293494 269809 293546 269815
rect 293506 263810 293534 269809
rect 293794 269725 293822 278004
rect 294646 275935 294698 275941
rect 294646 275877 294698 275883
rect 293974 269941 294026 269947
rect 293974 269883 294026 269889
rect 293782 269719 293834 269725
rect 293782 269661 293834 269667
rect 293986 263810 294014 269883
rect 294658 263824 294686 275877
rect 295138 269799 295166 278018
rect 295894 275861 295946 275867
rect 295894 275803 295946 275809
rect 295414 272679 295466 272685
rect 295414 272621 295466 272627
rect 295126 269793 295178 269799
rect 295126 269735 295178 269741
rect 295222 269127 295274 269133
rect 295222 269069 295274 269075
rect 295234 263824 295262 269069
rect 294432 263796 294686 263824
rect 295008 263796 295262 263824
rect 295426 263810 295454 272621
rect 295906 263810 295934 275803
rect 296386 269651 296414 278018
rect 297334 275787 297386 275793
rect 297334 275729 297386 275735
rect 297046 269793 297098 269799
rect 297046 269735 297098 269741
rect 296374 269645 296426 269651
rect 296374 269587 296426 269593
rect 296470 267129 296522 267135
rect 296470 267071 296522 267077
rect 296482 263824 296510 267071
rect 297058 263824 297086 269735
rect 296352 263796 296510 263824
rect 296832 263796 297086 263824
rect 297346 263810 297374 275729
rect 297538 272611 297566 278018
rect 297814 275639 297866 275645
rect 297814 275581 297866 275587
rect 297526 272605 297578 272611
rect 297526 272547 297578 272553
rect 297826 263810 297854 275581
rect 298294 272605 298346 272611
rect 298294 272547 298346 272553
rect 298006 272087 298058 272093
rect 298006 272029 298058 272035
rect 298018 268985 298046 272029
rect 298006 268979 298058 268985
rect 298006 268921 298058 268927
rect 298306 263810 298334 272547
rect 298690 272537 298718 278018
rect 298966 275713 299018 275719
rect 298966 275655 299018 275661
rect 298678 272531 298730 272537
rect 298678 272473 298730 272479
rect 298978 263824 299006 275655
rect 299350 275565 299402 275571
rect 299350 275507 299402 275513
rect 299362 263824 299390 275507
rect 299938 272981 299966 278018
rect 299926 272975 299978 272981
rect 299926 272917 299978 272923
rect 299446 272013 299498 272019
rect 299446 271955 299498 271961
rect 299458 267875 299486 271955
rect 299638 269719 299690 269725
rect 299638 269661 299690 269667
rect 299446 267869 299498 267875
rect 299446 267811 299498 267817
rect 298752 263796 299006 263824
rect 299232 263796 299390 263824
rect 299650 263810 299678 269661
rect 301090 269577 301118 278018
rect 301954 278004 302256 278032
rect 301846 275491 301898 275497
rect 301846 275433 301898 275439
rect 301366 272531 301418 272537
rect 301366 272473 301418 272479
rect 301078 269571 301130 269577
rect 301078 269513 301130 269519
rect 300694 268979 300746 268985
rect 300694 268921 300746 268927
rect 300214 267055 300266 267061
rect 300214 266997 300266 267003
rect 300226 263810 300254 266997
rect 300706 263810 300734 268921
rect 301378 263824 301406 272473
rect 301858 263824 301886 275433
rect 301954 271945 301982 278004
rect 303286 275417 303338 275423
rect 303286 275359 303338 275365
rect 301942 271939 301994 271945
rect 301942 271881 301994 271887
rect 302326 271939 302378 271945
rect 302326 271881 302378 271887
rect 302338 269059 302366 271881
rect 302614 269645 302666 269651
rect 302614 269587 302666 269593
rect 302326 269053 302378 269059
rect 302326 268995 302378 269001
rect 302038 266981 302090 266987
rect 302038 266923 302090 266929
rect 301152 263796 301406 263824
rect 301632 263796 301886 263824
rect 302050 263810 302078 266923
rect 302626 263810 302654 269587
rect 303298 263824 303326 275359
rect 303490 272389 303518 278018
rect 303478 272383 303530 272389
rect 303478 272325 303530 272331
rect 303958 272383 304010 272389
rect 303958 272325 304010 272331
rect 303766 268905 303818 268911
rect 303766 268847 303818 268853
rect 303778 263824 303806 268847
rect 303072 263796 303326 263824
rect 303552 263796 303806 263824
rect 303970 263810 303998 272325
rect 304642 269503 304670 278018
rect 305398 272975 305450 272981
rect 305398 272917 305450 272923
rect 304630 269497 304682 269503
rect 304630 269439 304682 269445
rect 305410 269133 305438 272917
rect 305794 272241 305822 278018
rect 306166 275343 306218 275349
rect 306166 275285 306218 275291
rect 305782 272235 305834 272241
rect 305782 272177 305834 272183
rect 305686 269571 305738 269577
rect 305686 269513 305738 269519
rect 305398 269127 305450 269133
rect 305398 269069 305450 269075
rect 304438 266907 304490 266913
rect 304438 266849 304490 266855
rect 304450 263810 304478 266849
rect 305014 266833 305066 266839
rect 305014 266775 305066 266781
rect 305026 263810 305054 266775
rect 305698 263824 305726 269513
rect 306178 263824 306206 275285
rect 306946 272463 306974 278018
rect 306934 272457 306986 272463
rect 306934 272399 306986 272405
rect 307126 272457 307178 272463
rect 307126 272399 307178 272405
rect 306358 269053 306410 269059
rect 306358 268995 306410 269001
rect 305472 263796 305726 263824
rect 305952 263796 306206 263824
rect 306370 263810 306398 268995
rect 307138 263824 307166 272399
rect 308194 269429 308222 278018
rect 308758 275269 308810 275275
rect 308758 275211 308810 275217
rect 308278 269497 308330 269503
rect 308278 269439 308330 269445
rect 308182 269423 308234 269429
rect 308182 269365 308234 269371
rect 308086 266759 308138 266765
rect 308086 266701 308138 266707
rect 307318 266685 307370 266691
rect 307318 266627 307370 266633
rect 306864 263796 307166 263824
rect 307330 263810 307358 266627
rect 308098 263824 308126 266701
rect 307872 263796 308126 263824
rect 308290 263810 308318 269439
rect 308770 263810 308798 275211
rect 309346 272315 309374 278018
rect 310390 275195 310442 275201
rect 310390 275137 310442 275143
rect 309334 272309 309386 272315
rect 309334 272251 309386 272257
rect 309910 272309 309962 272315
rect 309910 272251 309962 272257
rect 309238 269127 309290 269133
rect 309238 269069 309290 269075
rect 309250 263810 309278 269069
rect 309922 263824 309950 272251
rect 310402 263824 310430 275137
rect 310498 273499 310526 278018
rect 310486 273493 310538 273499
rect 310486 273435 310538 273441
rect 310582 273493 310634 273499
rect 310582 273435 310634 273441
rect 310594 268837 310622 273435
rect 311158 269423 311210 269429
rect 311158 269365 311210 269371
rect 310582 268831 310634 268837
rect 310582 268773 310634 268779
rect 310678 266611 310730 266617
rect 310678 266553 310730 266559
rect 309696 263796 309950 263824
rect 310272 263796 310430 263824
rect 310690 263810 310718 266553
rect 311170 263810 311198 269365
rect 311746 269281 311774 278018
rect 312790 272235 312842 272241
rect 312790 272177 312842 272183
rect 311734 269275 311786 269281
rect 311734 269217 311786 269223
rect 312310 268313 312362 268319
rect 312310 268255 312362 268261
rect 311638 266463 311690 266469
rect 311638 266405 311690 266411
rect 311650 263810 311678 266405
rect 312322 263824 312350 268255
rect 312802 263824 312830 272177
rect 312898 272167 312926 278018
rect 313078 275121 313130 275127
rect 313078 275063 313130 275069
rect 312886 272161 312938 272167
rect 312886 272103 312938 272109
rect 312096 263796 312350 263824
rect 312672 263796 312830 263824
rect 313090 263810 313118 275063
rect 313570 263810 313598 278319
rect 314902 278303 314954 278309
rect 404770 278300 405072 278319
rect 408322 278309 408624 278328
rect 408310 278303 408624 278309
rect 314902 278245 314954 278251
rect 408362 278300 408624 278303
rect 408310 278245 408362 278251
rect 314050 273425 314078 278018
rect 314710 275047 314762 275053
rect 314710 274989 314762 274995
rect 314038 273419 314090 273425
rect 314038 273361 314090 273367
rect 314230 269275 314282 269281
rect 314230 269217 314282 269223
rect 314242 263824 314270 269217
rect 314722 263824 314750 274989
rect 314016 263796 314270 263824
rect 314496 263796 314750 263824
rect 314914 263810 314942 278245
rect 316630 278229 316682 278235
rect 316630 278171 316682 278177
rect 411862 278229 411914 278235
rect 411914 278177 412176 278180
rect 411862 278171 412176 278177
rect 315298 269207 315326 278018
rect 316450 273573 316478 278018
rect 316438 273567 316490 273573
rect 316438 273509 316490 273515
rect 315478 272161 315530 272167
rect 315478 272103 315530 272109
rect 315286 269201 315338 269207
rect 315286 269143 315338 269149
rect 315490 263810 315518 272103
rect 315958 266537 316010 266543
rect 315958 266479 316010 266485
rect 315970 263810 315998 266479
rect 316642 263824 316670 278171
rect 319510 278155 319562 278161
rect 411874 278152 412176 278171
rect 418978 278161 419280 278180
rect 418966 278155 419280 278161
rect 319510 278097 319562 278103
rect 419018 278152 419280 278155
rect 418966 278097 419018 278103
rect 317302 274159 317354 274165
rect 317302 274101 317354 274107
rect 317110 267869 317162 267875
rect 317110 267811 317162 267817
rect 317122 263824 317150 267811
rect 316416 263796 316670 263824
rect 316896 263796 317150 263824
rect 317314 263810 317342 274101
rect 317602 273277 317630 278018
rect 317878 277711 317930 277717
rect 317878 277653 317930 277659
rect 317590 273271 317642 273277
rect 317590 273213 317642 273219
rect 317890 263810 317918 277653
rect 318358 271273 318410 271279
rect 318358 271215 318410 271221
rect 318370 263810 318398 271215
rect 318850 269355 318878 278018
rect 318934 274233 318986 274239
rect 318934 274175 318986 274181
rect 318838 269349 318890 269355
rect 318838 269291 318890 269297
rect 318946 263824 318974 274175
rect 319030 269349 319082 269355
rect 319030 269291 319082 269297
rect 319042 267875 319070 269291
rect 319030 267869 319082 267875
rect 319030 267811 319082 267817
rect 319522 263824 319550 278097
rect 320950 278081 321002 278087
rect 320950 278023 321002 278029
rect 422518 278081 422570 278087
rect 422570 278029 422832 278032
rect 422518 278023 422832 278029
rect 320002 270539 320030 278018
rect 319990 270533 320042 270539
rect 319990 270475 320042 270481
rect 319702 268387 319754 268393
rect 319702 268329 319754 268335
rect 318816 263796 318974 263824
rect 319296 263796 319550 263824
rect 319714 263810 319742 268329
rect 320182 265575 320234 265581
rect 320182 265517 320234 265523
rect 320194 263810 320222 265517
rect 320962 263824 320990 278023
rect 321154 273351 321182 278018
rect 322102 278007 322154 278013
rect 322102 277949 322154 277955
rect 321622 274381 321674 274387
rect 321622 274323 321674 274329
rect 321142 273345 321194 273351
rect 321142 273287 321194 273293
rect 321430 271347 321482 271353
rect 321430 271289 321482 271295
rect 321442 263824 321470 271289
rect 320736 263796 320990 263824
rect 321216 263796 321470 263824
rect 321634 263810 321662 274323
rect 322114 263810 322142 277949
rect 322402 270687 322430 278018
rect 323350 274307 323402 274313
rect 323350 274249 323402 274255
rect 322390 270681 322442 270687
rect 322390 270623 322442 270629
rect 322582 268461 322634 268467
rect 322582 268403 322634 268409
rect 322594 263810 322622 268403
rect 323362 263824 323390 274249
rect 323554 270613 323582 278018
rect 323830 277859 323882 277865
rect 323830 277801 323882 277807
rect 323542 270607 323594 270613
rect 323542 270549 323594 270555
rect 323842 263824 323870 277801
rect 324706 271945 324734 278018
rect 325858 274905 325886 278018
rect 326422 277785 326474 277791
rect 326422 277727 326474 277733
rect 325846 274899 325898 274905
rect 325846 274841 325898 274847
rect 325942 274455 325994 274461
rect 325942 274397 325994 274403
rect 324694 271939 324746 271945
rect 324694 271881 324746 271887
rect 324022 271199 324074 271205
rect 324022 271141 324074 271147
rect 323136 263796 323390 263824
rect 323616 263796 323870 263824
rect 324034 263810 324062 271141
rect 325750 268535 325802 268541
rect 325750 268477 325802 268483
rect 324502 265649 324554 265655
rect 324502 265591 324554 265597
rect 324514 263810 324542 265591
rect 324982 264095 325034 264101
rect 324982 264037 325034 264043
rect 324994 263810 325022 264037
rect 325762 263824 325790 268477
rect 325536 263796 325790 263824
rect 325954 263810 325982 274397
rect 326434 263810 326462 277727
rect 326806 273789 326858 273795
rect 326806 273731 326858 273737
rect 326818 268985 326846 273731
rect 327106 272093 327134 278018
rect 327094 272087 327146 272093
rect 327094 272029 327146 272035
rect 328258 272019 328286 278018
rect 329302 277637 329354 277643
rect 329302 277579 329354 277585
rect 328822 274529 328874 274535
rect 328822 274471 328874 274477
rect 328342 273937 328394 273943
rect 328342 273879 328394 273885
rect 328246 272013 328298 272019
rect 328246 271955 328298 271961
rect 326902 271495 326954 271501
rect 326902 271437 326954 271443
rect 326806 268979 326858 268985
rect 326806 268921 326858 268927
rect 326914 263810 326942 271437
rect 328354 268911 328382 273879
rect 328342 268905 328394 268911
rect 328342 268847 328394 268853
rect 328342 268609 328394 268615
rect 328342 268551 328394 268557
rect 327574 265723 327626 265729
rect 327574 265665 327626 265671
rect 327586 263824 327614 265665
rect 328054 264465 328106 264471
rect 328054 264407 328106 264413
rect 328066 263824 328094 264407
rect 327360 263796 327614 263824
rect 327840 263796 328094 263824
rect 328354 263810 328382 268551
rect 328834 263810 328862 274471
rect 329314 263810 329342 277579
rect 329410 274979 329438 278018
rect 329398 274973 329450 274979
rect 329398 274915 329450 274921
rect 329974 271569 330026 271575
rect 329974 271511 330026 271517
rect 329986 263824 330014 271511
rect 330658 270465 330686 278018
rect 330646 270459 330698 270465
rect 330646 270401 330698 270407
rect 331810 270391 331838 278018
rect 332962 276459 332990 278018
rect 333622 277563 333674 277569
rect 333622 277505 333674 277511
rect 332950 276453 333002 276459
rect 332950 276395 333002 276401
rect 333142 274677 333194 274683
rect 333142 274619 333194 274625
rect 331894 274603 331946 274609
rect 331894 274545 331946 274551
rect 331798 270385 331850 270391
rect 331798 270327 331850 270333
rect 331222 268683 331274 268689
rect 331222 268625 331274 268631
rect 330454 265797 330506 265803
rect 330454 265739 330506 265745
rect 330466 263824 330494 265739
rect 331126 264613 331178 264619
rect 331126 264555 331178 264561
rect 331138 263824 331166 264555
rect 329760 263796 330014 263824
rect 330240 263796 330494 263824
rect 330768 263796 331166 263824
rect 331234 263810 331262 268625
rect 331906 263824 331934 274545
rect 332566 271643 332618 271649
rect 332566 271585 332618 271591
rect 332374 268239 332426 268245
rect 332374 268181 332426 268187
rect 332386 263824 332414 268181
rect 331680 263796 331934 263824
rect 332160 263796 332414 263824
rect 332578 263810 332606 271585
rect 333154 263810 333182 274619
rect 333634 263810 333662 277505
rect 334210 273055 334238 278018
rect 334294 274011 334346 274017
rect 334294 273953 334346 273959
rect 334198 273049 334250 273055
rect 334198 272991 334250 272997
rect 334102 271421 334154 271427
rect 334102 271363 334154 271369
rect 334114 270317 334142 271363
rect 334102 270311 334154 270317
rect 334102 270253 334154 270259
rect 334306 269059 334334 273953
rect 335362 273203 335390 278018
rect 336514 276385 336542 278018
rect 336694 277489 336746 277495
rect 336694 277431 336746 277437
rect 336502 276379 336554 276385
rect 336502 276321 336554 276327
rect 336022 274751 336074 274757
rect 336022 274693 336074 274699
rect 335350 273197 335402 273203
rect 335350 273139 335402 273145
rect 335446 271717 335498 271723
rect 335446 271659 335498 271665
rect 334294 269053 334346 269059
rect 334294 268995 334346 269001
rect 334294 268757 334346 268763
rect 334294 268699 334346 268705
rect 334306 263824 334334 268699
rect 334966 268165 335018 268171
rect 334966 268107 335018 268113
rect 334774 265871 334826 265877
rect 334774 265813 334826 265819
rect 334786 263824 334814 265813
rect 334080 263796 334334 263824
rect 334560 263796 334814 263824
rect 334978 263810 335006 268107
rect 335458 263810 335486 271659
rect 336034 263810 336062 274693
rect 336706 263824 336734 277431
rect 337762 271427 337790 278018
rect 337942 273419 337994 273425
rect 337942 273361 337994 273367
rect 337750 271421 337802 271427
rect 337750 271363 337802 271369
rect 337954 270169 337982 273361
rect 338914 273129 338942 278018
rect 339286 277415 339338 277421
rect 339286 277357 339338 277363
rect 339094 274825 339146 274831
rect 339094 274767 339146 274773
rect 338902 273123 338954 273129
rect 338902 273065 338954 273071
rect 338614 271791 338666 271797
rect 338614 271733 338666 271739
rect 337942 270163 337994 270169
rect 337942 270105 337994 270111
rect 336886 268831 336938 268837
rect 336886 268773 336938 268779
rect 336480 263796 336734 263824
rect 336898 263824 336926 268773
rect 337846 268017 337898 268023
rect 337846 267959 337898 267965
rect 337366 265945 337418 265951
rect 337366 265887 337418 265893
rect 336898 263796 336960 263824
rect 337378 263810 337406 265887
rect 337858 263810 337886 267959
rect 338626 263824 338654 271733
rect 339106 263824 339134 274767
rect 338400 263796 338654 263824
rect 338880 263796 339134 263824
rect 339298 263810 339326 277357
rect 340066 276237 340094 278018
rect 340054 276231 340106 276237
rect 340054 276173 340106 276179
rect 341314 273425 341342 278018
rect 342166 277341 342218 277347
rect 342166 277283 342218 277289
rect 341686 274899 341738 274905
rect 341686 274841 341738 274847
rect 341302 273419 341354 273425
rect 341302 273361 341354 273367
rect 341494 271865 341546 271871
rect 341494 271807 341546 271813
rect 339766 268905 339818 268911
rect 339766 268847 339818 268853
rect 339778 263810 339806 268847
rect 341014 268091 341066 268097
rect 341014 268033 341066 268039
rect 340246 266019 340298 266025
rect 340246 265961 340298 265967
rect 340258 263810 340286 265961
rect 341026 263824 341054 268033
rect 341506 263824 341534 271807
rect 340800 263796 341054 263824
rect 341280 263796 341534 263824
rect 341698 263810 341726 274841
rect 342178 263810 342206 277283
rect 342466 270243 342494 278018
rect 343618 276311 343646 278018
rect 343606 276305 343658 276311
rect 343606 276247 343658 276253
rect 344566 274973 344618 274979
rect 344566 274915 344618 274921
rect 343606 273863 343658 273869
rect 343606 273805 343658 273811
rect 342742 271051 342794 271057
rect 342742 270993 342794 270999
rect 342454 270237 342506 270243
rect 342454 270179 342506 270185
rect 342754 270095 342782 270993
rect 342742 270089 342794 270095
rect 342742 270031 342794 270037
rect 343618 269133 343646 273805
rect 344086 271939 344138 271945
rect 344086 271881 344138 271887
rect 343606 269127 343658 269133
rect 343606 269069 343658 269075
rect 342646 268979 342698 268985
rect 342646 268921 342698 268927
rect 342658 263810 342686 268921
rect 343606 267943 343658 267949
rect 343606 267885 343658 267891
rect 343318 266093 343370 266099
rect 343318 266035 343370 266041
rect 343330 263824 343358 266035
rect 343104 263796 343358 263824
rect 343618 263810 343646 267885
rect 344098 263810 344126 271881
rect 344578 263810 344606 274915
rect 344770 273499 344798 278018
rect 344758 273493 344810 273499
rect 344758 273435 344810 273441
rect 346018 272907 346046 278018
rect 347170 276089 347198 278018
rect 347158 276083 347210 276089
rect 347158 276025 347210 276031
rect 347636 274346 347692 274355
rect 347636 274281 347692 274290
rect 347062 274085 347114 274091
rect 347062 274027 347114 274033
rect 346006 272901 346058 272907
rect 346006 272843 346058 272849
rect 346486 272013 346538 272019
rect 346486 271955 346538 271961
rect 345430 269053 345482 269059
rect 345430 268995 345482 269001
rect 344854 268239 344906 268245
rect 344854 268181 344906 268187
rect 345238 268239 345290 268245
rect 345238 268181 345290 268187
rect 344866 264545 344894 268181
rect 344854 264539 344906 264545
rect 344854 264481 344906 264487
rect 345250 263824 345278 268181
rect 345024 263796 345278 263824
rect 345442 263676 345470 268995
rect 346006 266167 346058 266173
rect 346006 266109 346058 266115
rect 346018 263810 346046 266109
rect 346498 263810 346526 271955
rect 346966 271421 347018 271427
rect 346966 271363 347018 271369
rect 346978 271205 347006 271363
rect 346966 271199 347018 271205
rect 346966 271141 347018 271147
rect 347074 268319 347102 274027
rect 347254 272087 347306 272093
rect 347254 272029 347306 272035
rect 347062 268313 347114 268319
rect 347062 268255 347114 268261
rect 347266 263824 347294 272029
rect 347650 263824 347678 274281
rect 348322 271057 348350 278018
rect 349462 273567 349514 273573
rect 349462 273509 349514 273515
rect 348310 271051 348362 271057
rect 348310 270993 348362 270999
rect 348118 269201 348170 269207
rect 348118 269143 348170 269149
rect 348130 263824 348158 269143
rect 348406 269127 348458 269133
rect 348406 269069 348458 269075
rect 346992 263796 347294 263824
rect 347424 263796 347678 263824
rect 347904 263796 348158 263824
rect 348418 263810 348446 269069
rect 348502 268165 348554 268171
rect 348502 268107 348554 268113
rect 348514 264693 348542 268107
rect 348886 266241 348938 266247
rect 348886 266183 348938 266189
rect 348502 264687 348554 264693
rect 348502 264629 348554 264635
rect 348898 263810 348926 266183
rect 349474 263824 349502 273509
rect 349570 270021 349598 278018
rect 350230 276453 350282 276459
rect 350230 276395 350282 276401
rect 350038 273493 350090 273499
rect 350038 273435 350090 273441
rect 349558 270015 349610 270021
rect 349558 269957 349610 269963
rect 350050 263824 350078 273435
rect 349344 263796 349502 263824
rect 349824 263796 350078 263824
rect 350242 263810 350270 276395
rect 350722 276163 350750 278018
rect 350710 276157 350762 276163
rect 350710 276099 350762 276105
rect 351874 272833 351902 278018
rect 352438 273419 352490 273425
rect 352438 273361 352490 273367
rect 351862 272827 351914 272833
rect 351862 272769 351914 272775
rect 351382 270755 351434 270761
rect 351382 270697 351434 270703
rect 350710 270681 350762 270687
rect 350710 270623 350762 270629
rect 350722 263810 350750 270623
rect 351286 270607 351338 270613
rect 351286 270549 351338 270555
rect 351298 263810 351326 270549
rect 351394 269873 351422 270697
rect 351382 269867 351434 269873
rect 351382 269809 351434 269815
rect 351958 266315 352010 266321
rect 351958 266257 352010 266263
rect 351970 263824 351998 266257
rect 352450 263824 352478 273361
rect 352630 273345 352682 273351
rect 352630 273287 352682 273293
rect 351744 263796 351998 263824
rect 352224 263796 352478 263824
rect 352642 263810 352670 273287
rect 353122 272759 353150 278018
rect 354274 276015 354302 278018
rect 354262 276009 354314 276015
rect 354262 275951 354314 275957
rect 353396 274494 353452 274503
rect 353396 274429 353452 274438
rect 353110 272753 353162 272759
rect 353110 272695 353162 272701
rect 353410 263824 353438 274429
rect 355030 273197 355082 273203
rect 355030 273139 355082 273145
rect 353686 270533 353738 270539
rect 353686 270475 353738 270481
rect 353136 263796 353438 263824
rect 353698 263810 353726 270475
rect 354070 270459 354122 270465
rect 354070 270401 354122 270407
rect 354082 264120 354110 270401
rect 354550 268239 354602 268245
rect 354550 268181 354602 268187
rect 354262 268017 354314 268023
rect 354262 267959 354314 267965
rect 354274 264767 354302 267959
rect 354562 267949 354590 268181
rect 354550 267943 354602 267949
rect 354550 267885 354602 267891
rect 354838 267795 354890 267801
rect 354838 267737 354890 267743
rect 354262 264761 354314 264767
rect 354262 264703 354314 264709
rect 354082 264092 354158 264120
rect 354130 263810 354158 264092
rect 354850 263824 354878 267737
rect 354624 263796 354878 263824
rect 355042 263810 355070 273139
rect 355426 270761 355454 278018
rect 356182 276379 356234 276385
rect 356182 276321 356234 276327
rect 355510 273271 355562 273277
rect 355510 273213 355562 273219
rect 355414 270755 355466 270761
rect 355414 270697 355466 270703
rect 355522 263810 355550 273213
rect 356194 263824 356222 276321
rect 356674 269947 356702 278018
rect 357826 275941 357854 278018
rect 357814 275935 357866 275941
rect 357814 275877 357866 275883
rect 358582 273123 358634 273129
rect 358582 273065 358634 273071
rect 357910 271199 357962 271205
rect 357910 271141 357962 271147
rect 356758 270385 356810 270391
rect 356758 270327 356810 270333
rect 356662 269941 356714 269947
rect 356662 269883 356714 269889
rect 356770 263824 356798 270327
rect 356950 270311 357002 270317
rect 356950 270253 357002 270259
rect 355968 263796 356222 263824
rect 356544 263796 356798 263824
rect 356962 263810 356990 270253
rect 357526 268017 357578 268023
rect 357526 267959 357578 267965
rect 357430 267721 357482 267727
rect 357430 267663 357482 267669
rect 357442 263810 357470 267663
rect 357538 264841 357566 267959
rect 357526 264835 357578 264841
rect 357526 264777 357578 264783
rect 357922 263810 357950 271141
rect 358594 263824 358622 273065
rect 358978 272981 359006 278018
rect 359158 276305 359210 276311
rect 359158 276247 359210 276253
rect 358966 272975 359018 272981
rect 358966 272917 359018 272923
rect 359170 263824 359198 276247
rect 360226 272685 360254 278018
rect 361378 275867 361406 278018
rect 361750 276231 361802 276237
rect 361750 276173 361802 276179
rect 361366 275861 361418 275867
rect 361366 275803 361418 275809
rect 360982 273049 361034 273055
rect 360982 272991 361034 272997
rect 360214 272679 360266 272685
rect 360214 272621 360266 272627
rect 359830 270237 359882 270243
rect 359830 270179 359882 270185
rect 359350 270163 359402 270169
rect 359350 270105 359402 270111
rect 358368 263796 358622 263824
rect 358944 263796 359198 263824
rect 359362 263810 359390 270105
rect 359842 263810 359870 270179
rect 360694 267869 360746 267875
rect 360694 267811 360746 267817
rect 360310 267647 360362 267653
rect 360310 267589 360362 267595
rect 360322 263810 360350 267589
rect 360706 264915 360734 267811
rect 360694 264909 360746 264915
rect 360694 264851 360746 264857
rect 360994 263824 361022 272991
rect 361270 272975 361322 272981
rect 361270 272917 361322 272923
rect 360768 263796 361022 263824
rect 361282 263810 361310 272917
rect 361762 263810 361790 276173
rect 362230 270089 362282 270095
rect 362230 270031 362282 270037
rect 362242 263810 362270 270031
rect 362530 267135 362558 278018
rect 363574 272901 363626 272907
rect 363574 272843 363626 272849
rect 362806 270015 362858 270021
rect 362806 269957 362858 269963
rect 362518 267129 362570 267135
rect 362518 267071 362570 267077
rect 362818 263824 362846 269957
rect 363382 267573 363434 267579
rect 363382 267515 363434 267521
rect 363394 263824 363422 267515
rect 362688 263796 362846 263824
rect 363168 263796 363422 263824
rect 363586 263810 363614 272843
rect 363682 269799 363710 278018
rect 364630 276157 364682 276163
rect 364630 276099 364682 276105
rect 364150 272827 364202 272833
rect 364150 272769 364202 272775
rect 363670 269793 363722 269799
rect 363670 269735 363722 269741
rect 364162 263810 364190 272769
rect 364642 263810 364670 276099
rect 364930 275793 364958 278018
rect 364918 275787 364970 275793
rect 364918 275729 364970 275735
rect 366082 275645 366110 278018
rect 366070 275639 366122 275645
rect 366070 275581 366122 275587
rect 366550 272753 366602 272759
rect 366550 272695 366602 272701
rect 365302 269941 365354 269947
rect 365302 269883 365354 269889
rect 365314 263824 365342 269883
rect 365686 269867 365738 269873
rect 365686 269809 365738 269815
rect 365698 263824 365726 269809
rect 365974 267499 366026 267505
rect 365974 267441 366026 267447
rect 365088 263796 365342 263824
rect 365568 263796 365726 263824
rect 365986 263810 366014 267441
rect 366562 263810 366590 272695
rect 367126 272679 367178 272685
rect 367126 272621 367178 272627
rect 367138 263824 367166 272621
rect 367234 272611 367262 278018
rect 367702 276083 367754 276089
rect 367702 276025 367754 276031
rect 367222 272605 367274 272611
rect 367222 272547 367274 272553
rect 367714 263824 367742 276025
rect 368482 275719 368510 278018
rect 368470 275713 368522 275719
rect 368470 275655 368522 275661
rect 369634 275571 369662 278018
rect 370294 275935 370346 275941
rect 370294 275877 370346 275883
rect 369622 275565 369674 275571
rect 369622 275507 369674 275513
rect 370100 271830 370156 271839
rect 370100 271765 370156 271774
rect 369620 271682 369676 271691
rect 369620 271617 369676 271626
rect 368372 269018 368428 269027
rect 368372 268953 368428 268962
rect 367892 268870 367948 268879
rect 367892 268805 367948 268814
rect 367008 263796 367166 263824
rect 367488 263796 367742 263824
rect 367906 263810 367934 268805
rect 368386 263810 368414 268953
rect 368950 267425 369002 267431
rect 368950 267367 369002 267373
rect 368962 263810 368990 267367
rect 369634 263824 369662 271617
rect 370114 263824 370142 271765
rect 369408 263796 369662 263824
rect 369888 263796 370142 263824
rect 370306 263810 370334 275877
rect 370786 269725 370814 278018
rect 371062 276009 371114 276015
rect 371062 275951 371114 275957
rect 370774 269719 370826 269725
rect 370774 269661 370826 269667
rect 371074 263824 371102 275951
rect 371926 275861 371978 275867
rect 371926 275803 371978 275809
rect 371254 269793 371306 269799
rect 371254 269735 371306 269741
rect 370800 263796 371102 263824
rect 371266 263810 371294 269735
rect 371938 263824 371966 275803
rect 372034 267061 372062 278018
rect 372502 277267 372554 277273
rect 372502 277209 372554 277215
rect 372022 267055 372074 267061
rect 372022 266997 372074 267003
rect 372514 263824 372542 277209
rect 373186 273795 373214 278018
rect 373846 277193 373898 277199
rect 373846 277135 373898 277141
rect 373460 274642 373516 274651
rect 373460 274577 373516 274586
rect 373174 273789 373226 273795
rect 373174 273731 373226 273737
rect 372694 272605 372746 272611
rect 372694 272547 372746 272553
rect 371808 263796 371966 263824
rect 372288 263796 372542 263824
rect 372706 263810 372734 272547
rect 373474 263824 373502 274577
rect 373858 263824 373886 277135
rect 374338 272537 374366 278018
rect 374614 275787 374666 275793
rect 374614 275729 374666 275735
rect 374326 272531 374378 272537
rect 374326 272473 374378 272479
rect 374324 269166 374380 269175
rect 374324 269101 374380 269110
rect 374338 263824 374366 269101
rect 373200 263796 373502 263824
rect 373632 263796 373886 263824
rect 374208 263796 374366 263824
rect 374626 263810 374654 275729
rect 375586 275497 375614 278018
rect 375574 275491 375626 275497
rect 375574 275433 375626 275439
rect 376244 274790 376300 274799
rect 376244 274725 376300 274734
rect 375190 273123 375242 273129
rect 375190 273065 375242 273071
rect 375202 271205 375230 273065
rect 375572 271978 375628 271987
rect 375572 271913 375628 271922
rect 375190 271199 375242 271205
rect 375190 271141 375242 271147
rect 375094 267351 375146 267357
rect 375094 267293 375146 267299
rect 375106 263810 375134 267293
rect 375586 263810 375614 271913
rect 376258 263824 376286 274725
rect 376738 266987 376766 278018
rect 376822 277119 376874 277125
rect 376822 277061 376874 277067
rect 376726 266981 376778 266987
rect 376726 266923 376778 266929
rect 376834 263824 376862 277061
rect 377494 275713 377546 275719
rect 377494 275655 377546 275661
rect 377012 270498 377068 270507
rect 377012 270433 377068 270442
rect 376032 263796 376286 263824
rect 376608 263796 376862 263824
rect 377026 263810 377054 270433
rect 377506 263810 377534 275655
rect 377890 269651 377918 278018
rect 377974 277045 378026 277051
rect 377974 276987 378026 276993
rect 377878 269645 377930 269651
rect 377878 269587 377930 269593
rect 377986 263810 378014 276987
rect 379138 275423 379166 278018
rect 379414 276897 379466 276903
rect 379414 276839 379466 276845
rect 379126 275417 379178 275423
rect 379126 275359 379178 275365
rect 379124 274938 379180 274947
rect 379124 274873 379180 274882
rect 378644 273458 378700 273467
rect 378644 273393 378700 273402
rect 378658 263824 378686 273393
rect 379138 263824 379166 274873
rect 378432 263796 378686 263824
rect 378912 263796 379166 263824
rect 379426 263810 379454 276839
rect 380290 273943 380318 278018
rect 381238 277933 381290 277939
rect 381238 277875 381290 277881
rect 381046 276971 381098 276977
rect 381046 276913 381098 276919
rect 380566 275639 380618 275645
rect 380566 275581 380618 275587
rect 380278 273937 380330 273943
rect 380278 273879 380330 273885
rect 379894 269719 379946 269725
rect 379894 269661 379946 269667
rect 379906 263810 379934 269661
rect 380578 263824 380606 275581
rect 381058 263824 381086 276913
rect 381250 273615 381278 277875
rect 381236 273606 381292 273615
rect 381236 273541 381292 273550
rect 381442 272389 381470 278018
rect 382294 276749 382346 276755
rect 382294 276691 382346 276697
rect 381812 275974 381868 275983
rect 381812 275909 381868 275918
rect 381430 272383 381482 272389
rect 381430 272325 381482 272331
rect 381236 267982 381292 267991
rect 381236 267917 381292 267926
rect 380352 263796 380606 263824
rect 380832 263796 381086 263824
rect 381250 263810 381278 267917
rect 381826 263810 381854 275909
rect 382306 263810 382334 276691
rect 382594 266913 382622 278018
rect 383638 276823 383690 276829
rect 383638 276765 383690 276771
rect 382964 273310 383020 273319
rect 382964 273245 383020 273254
rect 382582 266907 382634 266913
rect 382582 266849 382634 266855
rect 382978 263824 383006 273245
rect 383446 272383 383498 272389
rect 383446 272325 383498 272331
rect 383458 263824 383486 272325
rect 382752 263796 383006 263824
rect 383232 263796 383486 263824
rect 383650 263810 383678 276765
rect 383842 266839 383870 278018
rect 384118 269645 384170 269651
rect 384118 269587 384170 269593
rect 383830 266833 383882 266839
rect 383830 266775 383882 266781
rect 384130 263810 384158 269587
rect 384994 269577 385022 278018
rect 386146 275349 386174 278018
rect 386518 276675 386570 276681
rect 386518 276617 386570 276623
rect 386134 275343 386186 275349
rect 386134 275285 386186 275291
rect 385556 270350 385612 270359
rect 385556 270285 385612 270294
rect 384982 269571 385034 269577
rect 384982 269513 385034 269519
rect 385366 269571 385418 269577
rect 385366 269513 385418 269519
rect 384886 267277 384938 267283
rect 384886 267219 384938 267225
rect 384898 263824 384926 267219
rect 385378 263824 385406 269513
rect 385462 267943 385514 267949
rect 385462 267885 385514 267891
rect 385474 265359 385502 267885
rect 385462 265353 385514 265359
rect 385462 265295 385514 265301
rect 384672 263796 384926 263824
rect 385152 263796 385406 263824
rect 385570 263810 385598 270285
rect 386038 267203 386090 267209
rect 386038 267145 386090 267151
rect 386050 263810 386078 267145
rect 386530 263810 386558 276617
rect 387394 274017 387422 278018
rect 387766 275491 387818 275497
rect 387766 275433 387818 275439
rect 387382 274011 387434 274017
rect 387382 273953 387434 273959
rect 387284 273162 387340 273171
rect 387284 273097 387340 273106
rect 387298 263824 387326 273097
rect 387778 263824 387806 275433
rect 388546 272463 388574 278018
rect 388918 275565 388970 275571
rect 388918 275507 388970 275513
rect 388534 272457 388586 272463
rect 388534 272399 388586 272405
rect 388630 272457 388682 272463
rect 388630 272399 388682 272405
rect 388436 270202 388492 270211
rect 388436 270137 388492 270146
rect 387958 267129 388010 267135
rect 387958 267071 388010 267077
rect 387072 263796 387326 263824
rect 387552 263796 387806 263824
rect 387970 263810 387998 267071
rect 388450 263810 388478 270137
rect 388642 267991 388670 272399
rect 388628 267982 388684 267991
rect 388628 267917 388684 267926
rect 388930 263810 388958 275507
rect 389698 266691 389726 278018
rect 390838 276601 390890 276607
rect 390838 276543 390890 276549
rect 390356 275826 390412 275835
rect 390356 275761 390412 275770
rect 390164 273014 390220 273023
rect 390164 272949 390220 272958
rect 389686 266685 389738 266691
rect 389686 266627 389738 266633
rect 389446 264021 389498 264027
rect 389446 263963 389498 263969
rect 389458 263810 389486 263963
rect 390178 263824 390206 272949
rect 389952 263796 390206 263824
rect 390370 263810 390398 275761
rect 390850 263810 390878 276543
rect 390946 266765 390974 278018
rect 391508 270054 391564 270063
rect 391508 269989 391564 269998
rect 390934 266759 390986 266765
rect 390934 266701 390986 266707
rect 391522 263824 391550 269989
rect 392098 269503 392126 278018
rect 393250 275275 393278 278018
rect 393910 276527 393962 276533
rect 393910 276469 393962 276475
rect 393238 275269 393290 275275
rect 393238 275211 393290 275217
rect 392756 272866 392812 272875
rect 392756 272801 392812 272810
rect 392086 269497 392138 269503
rect 392086 269439 392138 269445
rect 391990 267055 392042 267061
rect 391990 266997 392042 267003
rect 392002 263824 392030 266997
rect 392278 263947 392330 263953
rect 392278 263889 392330 263895
rect 391296 263796 391550 263824
rect 391776 263796 392030 263824
rect 392290 263810 392318 263889
rect 392770 263810 392798 272801
rect 393238 266981 393290 266987
rect 393238 266923 393290 266929
rect 393250 263810 393278 266923
rect 393922 263824 393950 276469
rect 394498 273869 394526 278018
rect 394678 275417 394730 275423
rect 394678 275359 394730 275365
rect 394486 273863 394538 273869
rect 394486 273805 394538 273811
rect 394390 268239 394442 268245
rect 394390 268181 394442 268187
rect 394402 263824 394430 268181
rect 393696 263796 393950 263824
rect 394176 263796 394430 263824
rect 394690 263810 394718 275359
rect 395650 272315 395678 278018
rect 396692 276566 396748 276575
rect 396692 276501 396748 276510
rect 395638 272309 395690 272315
rect 395638 272251 395690 272257
rect 395926 272309 395978 272315
rect 395926 272251 395978 272257
rect 395446 263873 395498 263879
rect 395184 263821 395446 263824
rect 395938 263824 395966 272251
rect 396310 266907 396362 266913
rect 396310 266849 396362 266855
rect 396322 263824 396350 266849
rect 396706 263824 396734 276501
rect 396802 275201 396830 278018
rect 396790 275195 396842 275201
rect 396790 275137 396842 275143
rect 397558 274011 397610 274017
rect 397558 273953 397610 273959
rect 397076 269906 397132 269915
rect 397076 269841 397132 269850
rect 395184 263815 395498 263821
rect 395184 263796 395486 263815
rect 395664 263796 395966 263824
rect 396096 263796 396350 263824
rect 396576 263796 396734 263824
rect 397090 263810 397118 269841
rect 397570 263810 397598 273953
rect 398050 266617 398078 278018
rect 398230 275343 398282 275349
rect 398230 275285 398282 275291
rect 398038 266611 398090 266617
rect 398038 266553 398090 266559
rect 398242 263824 398270 275285
rect 398708 272718 398764 272727
rect 398708 272653 398764 272662
rect 398722 263824 398750 272653
rect 399202 269429 399230 278018
rect 399190 269423 399242 269429
rect 399190 269365 399242 269371
rect 399958 269423 400010 269429
rect 399958 269365 400010 269371
rect 398902 266833 398954 266839
rect 398902 266775 398954 266781
rect 398016 263796 398270 263824
rect 398496 263796 398750 263824
rect 398914 263810 398942 266775
rect 399408 263805 399710 263824
rect 399970 263810 399998 269365
rect 400354 266469 400382 278018
rect 400630 275269 400682 275275
rect 400630 275211 400682 275217
rect 400342 266463 400394 266469
rect 400342 266405 400394 266411
rect 400642 263824 400670 275211
rect 401506 274091 401534 278018
rect 402548 276714 402604 276723
rect 402548 276649 402604 276658
rect 401494 274085 401546 274091
rect 401494 274027 401546 274033
rect 401300 272570 401356 272579
rect 401300 272505 401356 272514
rect 399408 263799 399722 263805
rect 399408 263796 399670 263799
rect 400416 263796 400670 263824
rect 401314 263810 401342 272505
rect 401782 266759 401834 266765
rect 401782 266701 401834 266707
rect 401794 263810 401822 266701
rect 402562 263824 402590 276649
rect 402754 272241 402782 278018
rect 403222 275195 403274 275201
rect 403222 275137 403274 275143
rect 402742 272235 402794 272241
rect 402742 272177 402794 272183
rect 403028 269758 403084 269767
rect 403028 269693 403084 269702
rect 403042 263824 403070 269693
rect 402336 263796 402590 263824
rect 402816 263796 403070 263824
rect 403234 263810 403262 275137
rect 403906 275127 403934 278018
rect 403894 275121 403946 275127
rect 403894 275063 403946 275069
rect 404180 272422 404236 272431
rect 404180 272357 404236 272366
rect 403702 266685 403754 266691
rect 403702 266627 403754 266633
rect 403714 263810 403742 266627
rect 404194 263810 404222 272357
rect 406102 272235 406154 272241
rect 406102 272177 406154 272183
rect 405620 269610 405676 269619
rect 405620 269545 405676 269554
rect 404950 266611 405002 266617
rect 404950 266553 405002 266559
rect 404962 263824 404990 266553
rect 404736 263796 404990 263824
rect 405634 263810 405662 269545
rect 406114 269355 406142 272177
rect 406102 269349 406154 269355
rect 406102 269291 406154 269297
rect 406306 269281 406334 278018
rect 406390 275121 406442 275127
rect 406390 275063 406442 275069
rect 406294 269275 406346 269281
rect 406294 269217 406346 269223
rect 406402 263824 406430 275063
rect 407458 275053 407486 278018
rect 408980 275678 409036 275687
rect 408980 275613 409036 275622
rect 407926 275343 407978 275349
rect 407926 275285 407978 275291
rect 407446 275047 407498 275053
rect 407446 274989 407498 274995
rect 407938 274017 407966 275285
rect 407926 274011 407978 274017
rect 407926 273953 407978 273959
rect 408994 273615 409022 275613
rect 408980 273606 409036 273615
rect 408980 273541 409036 273550
rect 409858 272167 409886 278018
rect 410900 272274 410956 272283
rect 410900 272209 410956 272218
rect 409846 272161 409898 272167
rect 409846 272103 409898 272109
rect 409846 271199 409898 271205
rect 409846 271141 409898 271147
rect 409654 269349 409706 269355
rect 409654 269291 409706 269297
rect 408502 269275 408554 269281
rect 408502 269217 408554 269223
rect 407254 267869 407306 267875
rect 407254 267811 407306 267817
rect 407266 263824 407294 267811
rect 407830 266463 407882 266469
rect 407830 266405 407882 266411
rect 407842 263824 407870 266405
rect 408022 264169 408074 264175
rect 408022 264111 408074 264117
rect 406128 263796 406430 263824
rect 407040 263796 407294 263824
rect 407616 263796 407870 263824
rect 408034 263810 408062 264111
rect 408514 263810 408542 269217
rect 408982 266537 409034 266543
rect 408982 266479 409034 266485
rect 409174 266537 409226 266543
rect 409174 266479 409226 266485
rect 408994 265581 409022 266479
rect 408982 265575 409034 265581
rect 408982 265517 409034 265523
rect 409186 263824 409214 266479
rect 409666 263824 409694 269291
rect 409858 267875 409886 271141
rect 410420 269462 410476 269471
rect 410420 269397 410476 269406
rect 409846 267869 409898 267875
rect 409846 267811 409898 267817
rect 409942 267869 409994 267875
rect 409942 267811 409994 267817
rect 408960 263796 409214 263824
rect 409440 263796 409694 263824
rect 409954 263810 409982 267811
rect 410434 263810 410462 269397
rect 410914 263810 410942 272209
rect 411010 265581 411038 278018
rect 413410 272241 413438 278018
rect 414562 274165 414590 278018
rect 415714 277717 415742 278018
rect 415702 277711 415754 277717
rect 415702 277653 415754 277659
rect 414550 274159 414602 274165
rect 414550 274101 414602 274107
rect 413398 272235 413450 272241
rect 413398 272177 413450 272183
rect 413494 272235 413546 272241
rect 413494 272177 413546 272183
rect 411862 272161 411914 272167
rect 411764 272126 411820 272135
rect 411862 272103 411914 272109
rect 411764 272061 411820 272070
rect 411572 269314 411628 269323
rect 411572 269249 411628 269258
rect 410998 265575 411050 265581
rect 410998 265517 411050 265523
rect 411586 263824 411614 269249
rect 411360 263796 411614 263824
rect 411778 263824 411806 272061
rect 411874 267875 411902 272103
rect 413506 271205 413534 272177
rect 416962 271279 416990 278018
rect 418114 274239 418142 278018
rect 418102 274233 418154 274239
rect 418102 274175 418154 274181
rect 416950 271273 417002 271279
rect 416950 271215 417002 271221
rect 413494 271199 413546 271205
rect 413494 271141 413546 271147
rect 420514 268393 420542 278018
rect 420502 268387 420554 268393
rect 420502 268329 420554 268335
rect 411862 267869 411914 267875
rect 411862 267811 411914 267817
rect 421666 265433 421694 278018
rect 422530 278004 422832 278023
rect 423970 271353 423998 278018
rect 425218 274387 425246 278018
rect 426274 278013 426384 278032
rect 426262 278007 426384 278013
rect 426314 278004 426384 278007
rect 426262 277949 426314 277955
rect 425206 274381 425258 274387
rect 425206 274323 425258 274329
rect 423958 271347 424010 271353
rect 423958 271289 424010 271295
rect 427522 268467 427550 278018
rect 428770 274313 428798 278018
rect 429922 277865 429950 278018
rect 429910 277859 429962 277865
rect 429910 277801 429962 277807
rect 428758 274307 428810 274313
rect 428758 274249 428810 274255
rect 431074 271427 431102 278018
rect 431062 271421 431114 271427
rect 431062 271363 431114 271369
rect 427510 268461 427562 268467
rect 427510 268403 427562 268409
rect 432322 265655 432350 278018
rect 432310 265649 432362 265655
rect 432310 265591 432362 265597
rect 421654 265427 421706 265433
rect 421654 265369 421706 265375
rect 412822 264169 412874 264175
rect 412822 264111 412874 264117
rect 411778 263796 411840 263824
rect 399670 263741 399722 263747
rect 401110 263725 401162 263731
rect 345442 263648 345504 263676
rect 400896 263673 401110 263676
rect 400896 263667 401162 263673
rect 400896 263648 401150 263667
rect 406608 263657 406910 263676
rect 406608 263651 406922 263657
rect 406608 263648 406870 263651
rect 406870 263593 406922 263599
rect 405430 263577 405482 263583
rect 405216 263525 405430 263528
rect 405216 263519 405482 263525
rect 405216 263500 405470 263519
rect 412834 263509 412862 264111
rect 433474 264101 433502 278018
rect 434626 268541 434654 278018
rect 435874 274461 435902 278018
rect 437026 277791 437054 278018
rect 437014 277785 437066 277791
rect 437014 277727 437066 277733
rect 435862 274455 435914 274461
rect 435862 274397 435914 274403
rect 438178 271501 438206 278018
rect 438166 271495 438218 271501
rect 438166 271437 438218 271443
rect 434614 268535 434666 268541
rect 434614 268477 434666 268483
rect 439330 265729 439358 278018
rect 439318 265723 439370 265729
rect 439318 265665 439370 265671
rect 440578 264471 440606 278018
rect 441730 268615 441758 278018
rect 442882 274535 442910 278018
rect 444130 277643 444158 278018
rect 444118 277637 444170 277643
rect 444118 277579 444170 277585
rect 442870 274529 442922 274535
rect 442870 274471 442922 274477
rect 445282 271575 445310 278018
rect 445270 271569 445322 271575
rect 445270 271511 445322 271517
rect 441718 268609 441770 268615
rect 441718 268551 441770 268557
rect 446434 265803 446462 278018
rect 446422 265797 446474 265803
rect 446422 265739 446474 265745
rect 447682 264619 447710 278018
rect 448834 268689 448862 278018
rect 449986 274609 450014 278018
rect 449974 274603 450026 274609
rect 449974 274545 450026 274551
rect 448822 268683 448874 268689
rect 448822 268625 448874 268631
rect 447670 264613 447722 264619
rect 447670 264555 447722 264561
rect 451234 264545 451262 278018
rect 452386 271649 452414 278018
rect 453538 274683 453566 278018
rect 454786 277569 454814 278018
rect 454774 277563 454826 277569
rect 454774 277505 454826 277511
rect 453526 274677 453578 274683
rect 453526 274619 453578 274625
rect 452374 271643 452426 271649
rect 452374 271585 452426 271591
rect 455938 268763 455966 278018
rect 455926 268757 455978 268763
rect 455926 268699 455978 268705
rect 457090 265877 457118 278018
rect 457078 265871 457130 265877
rect 457078 265813 457130 265819
rect 458242 264693 458270 278018
rect 459490 271723 459518 278018
rect 460642 274757 460670 278018
rect 461794 277495 461822 278018
rect 461782 277489 461834 277495
rect 461782 277431 461834 277437
rect 460630 274751 460682 274757
rect 460630 274693 460682 274699
rect 459478 271717 459530 271723
rect 459478 271659 459530 271665
rect 463042 268837 463070 278018
rect 463030 268831 463082 268837
rect 463030 268773 463082 268779
rect 464194 265951 464222 278018
rect 464182 265945 464234 265951
rect 464182 265887 464234 265893
rect 465346 264767 465374 278018
rect 466594 271797 466622 278018
rect 467746 274831 467774 278018
rect 468898 277421 468926 278018
rect 468886 277415 468938 277421
rect 468886 277357 468938 277363
rect 467734 274825 467786 274831
rect 467734 274767 467786 274773
rect 466582 271791 466634 271797
rect 466582 271733 466634 271739
rect 470146 268911 470174 278018
rect 470134 268905 470186 268911
rect 470134 268847 470186 268853
rect 471298 266025 471326 278018
rect 471286 266019 471338 266025
rect 471286 265961 471338 265967
rect 472450 264841 472478 278018
rect 473698 271871 473726 278018
rect 474850 274905 474878 278018
rect 476002 277347 476030 278018
rect 475990 277341 476042 277347
rect 475990 277283 476042 277289
rect 474838 274899 474890 274905
rect 474838 274841 474890 274847
rect 473686 271865 473738 271871
rect 473686 271807 473738 271813
rect 477154 268985 477182 278018
rect 477142 268979 477194 268985
rect 477142 268921 477194 268927
rect 478402 266099 478430 278018
rect 478390 266093 478442 266099
rect 478390 266035 478442 266041
rect 479554 264915 479582 278018
rect 480706 271945 480734 278018
rect 481954 274979 481982 278018
rect 481942 274973 481994 274979
rect 481942 274915 481994 274921
rect 480694 271939 480746 271945
rect 480694 271881 480746 271887
rect 483106 265507 483134 278018
rect 484258 269059 484286 278018
rect 484246 269053 484298 269059
rect 484246 268995 484298 269001
rect 485506 266173 485534 278018
rect 486658 272019 486686 278018
rect 487810 272093 487838 278018
rect 489058 274355 489086 278018
rect 489044 274346 489100 274355
rect 489044 274281 489100 274290
rect 487798 272087 487850 272093
rect 487798 272029 487850 272035
rect 486646 272013 486698 272019
rect 486646 271955 486698 271961
rect 490210 269207 490238 278018
rect 490198 269201 490250 269207
rect 490198 269143 490250 269149
rect 491362 269133 491390 278018
rect 491350 269127 491402 269133
rect 491350 269069 491402 269075
rect 492610 266247 492638 278018
rect 493762 273573 493790 278018
rect 493750 273567 493802 273573
rect 493750 273509 493802 273515
rect 494914 273499 494942 278018
rect 496066 276459 496094 278018
rect 496054 276453 496106 276459
rect 496054 276395 496106 276401
rect 494902 273493 494954 273499
rect 494902 273435 494954 273441
rect 497314 270687 497342 278018
rect 497302 270681 497354 270687
rect 497302 270623 497354 270629
rect 498466 270613 498494 278018
rect 498454 270607 498506 270613
rect 498454 270549 498506 270555
rect 499618 266321 499646 278018
rect 500866 273425 500894 278018
rect 500854 273419 500906 273425
rect 500854 273361 500906 273367
rect 502018 273351 502046 278018
rect 503170 274503 503198 278018
rect 503156 274494 503212 274503
rect 503156 274429 503212 274438
rect 502006 273345 502058 273351
rect 502006 273287 502058 273293
rect 504418 270539 504446 278018
rect 504406 270533 504458 270539
rect 504406 270475 504458 270481
rect 505570 270465 505598 278018
rect 505558 270459 505610 270465
rect 505558 270401 505610 270407
rect 506722 267801 506750 278018
rect 507970 273203 507998 278018
rect 509122 273277 509150 278018
rect 510274 276385 510302 278018
rect 510262 276379 510314 276385
rect 510262 276321 510314 276327
rect 509110 273271 509162 273277
rect 509110 273213 509162 273219
rect 507958 273197 508010 273203
rect 507958 273139 508010 273145
rect 511522 270391 511550 278018
rect 511510 270385 511562 270391
rect 511510 270327 511562 270333
rect 512674 270317 512702 278018
rect 512662 270311 512714 270317
rect 512662 270253 512714 270259
rect 506710 267795 506762 267801
rect 506710 267737 506762 267743
rect 513826 267727 513854 278018
rect 514978 273129 515006 278018
rect 514966 273123 515018 273129
rect 514966 273065 515018 273071
rect 516226 273055 516254 278018
rect 517378 276311 517406 278018
rect 517366 276305 517418 276311
rect 517366 276247 517418 276253
rect 516214 273049 516266 273055
rect 516214 272991 516266 272997
rect 518530 270169 518558 278018
rect 519778 270243 519806 278018
rect 519766 270237 519818 270243
rect 519766 270179 519818 270185
rect 518518 270163 518570 270169
rect 518518 270105 518570 270111
rect 513814 267721 513866 267727
rect 513814 267663 513866 267669
rect 520930 267653 520958 278018
rect 522082 272981 522110 278018
rect 522070 272975 522122 272981
rect 522070 272917 522122 272923
rect 523330 272907 523358 278018
rect 524482 276237 524510 278018
rect 524470 276231 524522 276237
rect 524470 276173 524522 276179
rect 523318 272901 523370 272907
rect 523318 272843 523370 272849
rect 525634 270095 525662 278018
rect 525622 270089 525674 270095
rect 525622 270031 525674 270037
rect 526882 270021 526910 278018
rect 526870 270015 526922 270021
rect 526870 269957 526922 269963
rect 520918 267647 520970 267653
rect 520918 267589 520970 267595
rect 528034 267579 528062 278018
rect 529186 272833 529214 278018
rect 529844 276714 529900 276723
rect 529844 276649 529900 276658
rect 529858 273573 529886 276649
rect 529846 273567 529898 273573
rect 529846 273509 529898 273515
rect 529174 272827 529226 272833
rect 529174 272769 529226 272775
rect 530434 272759 530462 278018
rect 531586 276163 531614 278018
rect 531574 276157 531626 276163
rect 531574 276099 531626 276105
rect 530422 272753 530474 272759
rect 530422 272695 530474 272701
rect 532738 269947 532766 278018
rect 532726 269941 532778 269947
rect 532726 269883 532778 269889
rect 533890 269873 533918 278018
rect 533878 269867 533930 269873
rect 533878 269809 533930 269815
rect 528022 267573 528074 267579
rect 528022 267515 528074 267521
rect 535138 267505 535166 278018
rect 536290 272685 536318 278018
rect 536278 272679 536330 272685
rect 536278 272621 536330 272627
rect 537442 272611 537470 278018
rect 538690 276089 538718 278018
rect 538678 276083 538730 276089
rect 538678 276025 538730 276031
rect 537430 272605 537482 272611
rect 537430 272547 537482 272553
rect 539842 268879 539870 278018
rect 540994 269027 541022 278018
rect 540980 269018 541036 269027
rect 540980 268953 541036 268962
rect 539828 268870 539884 268879
rect 539828 268805 539884 268814
rect 535126 267499 535178 267505
rect 535126 267441 535178 267447
rect 542242 267431 542270 278018
rect 543394 271691 543422 278018
rect 544546 271839 544574 278018
rect 545794 275941 545822 278018
rect 546946 276015 546974 278018
rect 546934 276009 546986 276015
rect 546934 275951 546986 275957
rect 545782 275935 545834 275941
rect 545782 275877 545834 275883
rect 544532 271830 544588 271839
rect 544532 271765 544588 271774
rect 543380 271682 543436 271691
rect 543380 271617 543436 271626
rect 548098 269799 548126 278018
rect 549346 275867 549374 278018
rect 550498 277273 550526 278018
rect 550486 277267 550538 277273
rect 550486 277209 550538 277215
rect 549334 275861 549386 275867
rect 549334 275803 549386 275809
rect 551650 272537 551678 278018
rect 552802 274651 552830 278018
rect 554050 277199 554078 278018
rect 554038 277193 554090 277199
rect 554038 277135 554090 277141
rect 552788 274642 552844 274651
rect 552788 274577 552844 274586
rect 551638 272531 551690 272537
rect 551638 272473 551690 272479
rect 548086 269793 548138 269799
rect 548086 269735 548138 269741
rect 555202 269175 555230 278018
rect 556354 275793 556382 278018
rect 556342 275787 556394 275793
rect 556342 275729 556394 275735
rect 555188 269166 555244 269175
rect 555188 269101 555244 269110
rect 542230 267425 542282 267431
rect 542230 267367 542282 267373
rect 557602 267357 557630 278018
rect 558754 271987 558782 278018
rect 559906 274799 559934 278018
rect 561154 277125 561182 278018
rect 561142 277119 561194 277125
rect 561142 277061 561194 277067
rect 559892 274790 559948 274799
rect 559892 274725 559948 274734
rect 558740 271978 558796 271987
rect 558740 271913 558796 271922
rect 562306 270507 562334 278018
rect 563458 275719 563486 278018
rect 564706 277051 564734 278018
rect 564694 277045 564746 277051
rect 564694 276987 564746 276993
rect 563446 275713 563498 275719
rect 563446 275655 563498 275661
rect 565858 273467 565886 278018
rect 567010 274947 567038 278018
rect 568258 276903 568286 278018
rect 568246 276897 568298 276903
rect 568246 276839 568298 276845
rect 566996 274938 567052 274947
rect 566996 274873 567052 274882
rect 565844 273458 565900 273467
rect 565844 273393 565900 273402
rect 562292 270498 562348 270507
rect 562292 270433 562348 270442
rect 569410 269725 569438 278018
rect 570562 275645 570590 278018
rect 571714 276977 571742 278018
rect 571702 276971 571754 276977
rect 571702 276913 571754 276919
rect 570550 275639 570602 275645
rect 570550 275581 570602 275587
rect 572962 272463 572990 278018
rect 574114 275983 574142 278018
rect 575266 276755 575294 278018
rect 575254 276749 575306 276755
rect 575254 276691 575306 276697
rect 574100 275974 574156 275983
rect 574100 275909 574156 275918
rect 576514 273319 576542 278018
rect 576500 273310 576556 273319
rect 576500 273245 576556 273254
rect 572950 272457 573002 272463
rect 572950 272399 573002 272405
rect 577666 272389 577694 278018
rect 578818 276829 578846 278018
rect 578806 276823 578858 276829
rect 578806 276765 578858 276771
rect 577654 272383 577706 272389
rect 577654 272325 577706 272331
rect 569398 269719 569450 269725
rect 569398 269661 569450 269667
rect 580066 269651 580094 278018
rect 580054 269645 580106 269651
rect 580054 269587 580106 269593
rect 557590 267351 557642 267357
rect 557590 267293 557642 267299
rect 581218 267283 581246 278018
rect 582370 269577 582398 278018
rect 583618 270359 583646 278018
rect 583604 270350 583660 270359
rect 583604 270285 583660 270294
rect 582358 269571 582410 269577
rect 582358 269513 582410 269519
rect 581206 267277 581258 267283
rect 581206 267219 581258 267225
rect 584770 267209 584798 278018
rect 585922 276681 585950 278018
rect 585910 276675 585962 276681
rect 585910 276617 585962 276623
rect 587170 273171 587198 278018
rect 588322 275497 588350 278018
rect 588310 275491 588362 275497
rect 588310 275433 588362 275439
rect 587156 273162 587212 273171
rect 587156 273097 587212 273106
rect 584758 267203 584810 267209
rect 584758 267145 584810 267151
rect 589474 267135 589502 278018
rect 590626 270211 590654 278018
rect 591874 275571 591902 278018
rect 591862 275565 591914 275571
rect 591862 275507 591914 275513
rect 590612 270202 590668 270211
rect 590612 270137 590668 270146
rect 589462 267129 589514 267135
rect 589462 267071 589514 267077
rect 499606 266315 499658 266321
rect 499606 266257 499658 266263
rect 492598 266241 492650 266247
rect 492598 266183 492650 266189
rect 485494 266167 485546 266173
rect 485494 266109 485546 266115
rect 483094 265501 483146 265507
rect 483094 265443 483146 265449
rect 479542 264909 479594 264915
rect 479542 264851 479594 264857
rect 472438 264835 472490 264841
rect 472438 264777 472490 264783
rect 465334 264761 465386 264767
rect 465334 264703 465386 264709
rect 458230 264687 458282 264693
rect 458230 264629 458282 264635
rect 451222 264539 451274 264545
rect 451222 264481 451274 264487
rect 440566 264465 440618 264471
rect 440566 264407 440618 264413
rect 433462 264095 433514 264101
rect 433462 264037 433514 264043
rect 593026 264027 593054 278018
rect 594178 273023 594206 278018
rect 595426 275835 595454 278018
rect 596578 276607 596606 278018
rect 596566 276601 596618 276607
rect 596566 276543 596618 276549
rect 595412 275826 595468 275835
rect 595412 275761 595468 275770
rect 594164 273014 594220 273023
rect 594164 272949 594220 272958
rect 597730 270063 597758 278018
rect 597716 270054 597772 270063
rect 597716 269989 597772 269998
rect 598978 267061 599006 278018
rect 598966 267055 599018 267061
rect 598966 266997 599018 267003
rect 593014 264021 593066 264027
rect 593014 263963 593066 263969
rect 600130 263953 600158 278018
rect 601282 272875 601310 278018
rect 601268 272866 601324 272875
rect 601268 272801 601324 272810
rect 602530 266987 602558 278018
rect 603682 276533 603710 278018
rect 603670 276527 603722 276533
rect 603670 276469 603722 276475
rect 604834 268245 604862 278018
rect 606082 275423 606110 278018
rect 606070 275417 606122 275423
rect 606070 275359 606122 275365
rect 604822 268239 604874 268245
rect 604822 268181 604874 268187
rect 602518 266981 602570 266987
rect 602518 266923 602570 266929
rect 600118 263947 600170 263953
rect 600118 263889 600170 263895
rect 607234 263879 607262 278018
rect 608386 272315 608414 278018
rect 608374 272309 608426 272315
rect 608374 272251 608426 272257
rect 609538 266913 609566 278018
rect 610786 276575 610814 278018
rect 610772 276566 610828 276575
rect 610772 276501 610828 276510
rect 611938 269915 611966 278018
rect 613090 275349 613118 278018
rect 613078 275343 613130 275349
rect 613078 275285 613130 275291
rect 614338 275275 614366 278018
rect 614326 275269 614378 275275
rect 614326 275211 614378 275217
rect 615490 272727 615518 278018
rect 615476 272718 615532 272727
rect 615476 272653 615532 272662
rect 611924 269906 611980 269915
rect 611924 269841 611980 269850
rect 609526 266907 609578 266913
rect 609526 266849 609578 266855
rect 616642 266839 616670 278018
rect 616630 266833 616682 266839
rect 616630 266775 616682 266781
rect 607222 263873 607274 263879
rect 607222 263815 607274 263821
rect 617890 263805 617918 278018
rect 619042 269429 619070 278018
rect 620194 275201 620222 278018
rect 620182 275195 620234 275201
rect 620182 275137 620234 275143
rect 619030 269423 619082 269429
rect 619030 269365 619082 269371
rect 617878 263799 617930 263805
rect 617878 263741 617930 263747
rect 621442 263731 621470 278018
rect 622594 272579 622622 278018
rect 622580 272570 622636 272579
rect 622580 272505 622636 272514
rect 623746 266765 623774 278018
rect 624994 273573 625022 278018
rect 624982 273567 625034 273573
rect 624982 273509 625034 273515
rect 626146 269767 626174 278018
rect 627298 275127 627326 278018
rect 627286 275121 627338 275127
rect 627286 275063 627338 275069
rect 626132 269758 626188 269767
rect 626132 269693 626188 269702
rect 623734 266759 623786 266765
rect 623734 266701 623786 266707
rect 628450 266691 628478 278018
rect 629698 272431 629726 278018
rect 629684 272422 629740 272431
rect 629684 272357 629740 272366
rect 628438 266685 628490 266691
rect 628438 266627 628490 266633
rect 630850 266617 630878 278018
rect 630838 266611 630890 266617
rect 630838 266553 630890 266559
rect 621430 263725 621482 263731
rect 621430 263667 621482 263673
rect 632002 263657 632030 278018
rect 633250 269619 633278 278018
rect 634402 275053 634430 278018
rect 634390 275047 634442 275053
rect 634390 274989 634442 274995
rect 633236 269610 633292 269619
rect 633236 269545 633292 269554
rect 427606 263651 427658 263657
rect 427606 263593 427658 263599
rect 631990 263651 632042 263657
rect 631990 263593 632042 263599
rect 427618 263528 427646 263593
rect 635554 263583 635582 278018
rect 636802 272241 636830 278018
rect 636790 272235 636842 272241
rect 636790 272177 636842 272183
rect 637954 266469 637982 278018
rect 637942 266463 637994 266469
rect 637942 266405 637994 266411
rect 427894 263577 427946 263583
rect 427618 263525 427894 263528
rect 427618 263519 427946 263525
rect 635542 263577 635594 263583
rect 635542 263519 635594 263525
rect 412822 263503 412874 263509
rect 427618 263500 427934 263519
rect 639106 263509 639134 278018
rect 640354 269281 640382 278018
rect 640342 269275 640394 269281
rect 640342 269217 640394 269223
rect 641506 266543 641534 278018
rect 642658 269355 642686 278018
rect 643906 272167 643934 278018
rect 643894 272161 643946 272167
rect 643894 272103 643946 272109
rect 645058 269471 645086 278018
rect 646210 272283 646238 278018
rect 646580 277306 646636 277315
rect 646580 277241 646636 277250
rect 646484 275530 646540 275539
rect 646484 275465 646540 275474
rect 646196 272274 646252 272283
rect 646196 272209 646252 272218
rect 645044 269462 645100 269471
rect 645044 269397 645100 269406
rect 642646 269349 642698 269355
rect 642646 269291 642698 269297
rect 641494 266537 641546 266543
rect 641494 266479 641546 266485
rect 639094 263503 639146 263509
rect 412822 263445 412874 263451
rect 639094 263445 639146 263451
rect 420404 262210 420460 262219
rect 420404 262145 420406 262154
rect 420458 262145 420460 262154
rect 606166 262171 606218 262177
rect 420406 262113 420458 262119
rect 606166 262113 606218 262119
rect 420404 259842 420460 259851
rect 420404 259777 420460 259786
rect 191540 259398 191596 259407
rect 191540 259333 191596 259342
rect 190196 251702 190252 251711
rect 190196 251637 190252 251646
rect 190210 228581 190238 251637
rect 190198 228575 190250 228581
rect 190198 228517 190250 228523
rect 190774 227539 190826 227545
rect 190774 227481 190826 227487
rect 190786 221792 190814 227481
rect 190786 221764 190862 221792
rect 190834 221482 190862 221764
rect 191554 221482 191582 259333
rect 420418 259291 420446 259777
rect 420406 259285 420458 259291
rect 420406 259227 420458 259233
rect 420404 257030 420460 257039
rect 420404 256965 420460 256974
rect 420418 256405 420446 256965
rect 420406 256399 420458 256405
rect 420406 256341 420458 256347
rect 420404 255254 420460 255263
rect 420404 255189 420460 255198
rect 420418 253519 420446 255189
rect 420406 253513 420458 253519
rect 420406 253455 420458 253461
rect 603286 253513 603338 253519
rect 603286 253455 603338 253461
rect 420404 252886 420460 252895
rect 420404 252821 420460 252830
rect 420418 250633 420446 252821
rect 420406 250627 420458 250633
rect 420406 250569 420458 250575
rect 420308 250518 420364 250527
rect 420308 250453 420364 250462
rect 420322 247821 420350 250453
rect 420404 248150 420460 248159
rect 420404 248085 420460 248094
rect 420310 247815 420362 247821
rect 420310 247757 420362 247763
rect 420418 247747 420446 248085
rect 420406 247741 420458 247747
rect 420406 247683 420458 247689
rect 420404 245338 420460 245347
rect 420404 245273 420460 245282
rect 420418 244861 420446 245273
rect 420406 244855 420458 244861
rect 420406 244797 420458 244803
rect 420404 243562 420460 243571
rect 420404 243497 420460 243506
rect 420418 241975 420446 243497
rect 420406 241969 420458 241975
rect 420406 241911 420458 241917
rect 600406 241969 600458 241975
rect 600406 241911 600458 241917
rect 420404 241194 420460 241203
rect 420404 241129 420460 241138
rect 412148 240158 412204 240167
rect 412148 240093 412204 240102
rect 412052 240010 412108 240019
rect 380640 239977 380894 239996
rect 380640 239971 380906 239977
rect 380640 239968 380854 239971
rect 412052 239945 412054 239954
rect 380854 239913 380906 239919
rect 412106 239945 412108 239954
rect 412054 239913 412106 239919
rect 412162 239903 412190 240093
rect 409558 239897 409610 239903
rect 409344 239845 409558 239848
rect 409344 239839 409610 239845
rect 412150 239897 412202 239903
rect 412150 239839 412202 239845
rect 357142 239823 357194 239829
rect 409344 239820 409598 239839
rect 357142 239765 357194 239771
rect 192418 233391 192446 239686
rect 192768 239672 192926 239700
rect 192898 233613 192926 239672
rect 192994 239672 193152 239700
rect 192886 233607 192938 233613
rect 192886 233549 192938 233555
rect 192406 233385 192458 233391
rect 192406 233327 192458 233333
rect 192310 228575 192362 228581
rect 192310 228517 192362 228523
rect 192322 221482 192350 228517
rect 192994 221792 193022 239672
rect 193474 233317 193502 239686
rect 193858 233391 193886 239686
rect 194242 233539 194270 239686
rect 194230 233533 194282 233539
rect 194230 233475 194282 233481
rect 194626 233465 194654 239686
rect 194976 239672 195230 239700
rect 195360 239672 195614 239700
rect 194614 233459 194666 233465
rect 194614 233401 194666 233407
rect 193750 233385 193802 233391
rect 193750 233327 193802 233333
rect 193846 233385 193898 233391
rect 193846 233327 193898 233333
rect 193462 233311 193514 233317
rect 193462 233253 193514 233259
rect 192994 221764 193070 221792
rect 193042 221482 193070 221764
rect 193762 221482 193790 233327
rect 195202 233317 195230 239672
rect 195586 233613 195614 239672
rect 195682 233687 195710 239686
rect 195670 233681 195722 233687
rect 195670 233623 195722 233629
rect 195286 233607 195338 233613
rect 195286 233549 195338 233555
rect 195574 233607 195626 233613
rect 195574 233549 195626 233555
rect 194614 233311 194666 233317
rect 194614 233253 194666 233259
rect 195190 233311 195242 233317
rect 195190 233253 195242 233259
rect 194626 221482 194654 233253
rect 195298 221792 195326 233549
rect 196162 233465 196190 239686
rect 196546 233761 196574 239686
rect 196930 233835 196958 239686
rect 197280 239672 197534 239700
rect 197664 239672 197918 239700
rect 197506 233983 197534 239672
rect 197494 233977 197546 233983
rect 197494 233919 197546 233925
rect 196918 233829 196970 233835
rect 196918 233771 196970 233777
rect 196534 233755 196586 233761
rect 196534 233697 196586 233703
rect 196054 233459 196106 233465
rect 196054 233401 196106 233407
rect 196150 233459 196202 233465
rect 196150 233401 196202 233407
rect 195298 221764 195374 221792
rect 195346 221482 195374 221764
rect 196066 221482 196094 233401
rect 196822 233385 196874 233391
rect 196822 233327 196874 233333
rect 196834 221482 196862 233327
rect 197890 233317 197918 239672
rect 197986 233391 198014 239686
rect 198370 234057 198398 239686
rect 198754 234131 198782 239686
rect 198742 234125 198794 234131
rect 198742 234067 198794 234073
rect 198358 234051 198410 234057
rect 198358 233993 198410 233999
rect 199138 233909 199166 239686
rect 199488 239672 199742 239700
rect 199968 239672 200222 239700
rect 199126 233903 199178 233909
rect 199126 233845 199178 233851
rect 198358 233533 198410 233539
rect 198358 233475 198410 233481
rect 197974 233385 198026 233391
rect 197974 233327 198026 233333
rect 197494 233311 197546 233317
rect 197494 233253 197546 233259
rect 197878 233311 197930 233317
rect 197878 233253 197930 233259
rect 197506 221792 197534 233253
rect 197506 221764 197582 221792
rect 197554 221482 197582 221764
rect 198370 221482 198398 233475
rect 199714 233465 199742 239672
rect 200194 234205 200222 239672
rect 200290 234279 200318 239686
rect 200278 234273 200330 234279
rect 200278 234215 200330 234221
rect 200182 234199 200234 234205
rect 200182 234141 200234 234147
rect 200566 233755 200618 233761
rect 200566 233697 200618 233703
rect 199798 233607 199850 233613
rect 199798 233549 199850 233555
rect 199126 233459 199178 233465
rect 199126 233401 199178 233407
rect 199702 233459 199754 233465
rect 199702 233401 199754 233407
rect 199138 221482 199166 233401
rect 199810 221792 199838 233549
rect 199810 221764 199886 221792
rect 199858 221482 199886 221764
rect 200578 221482 200606 233697
rect 200674 233539 200702 239686
rect 201058 233613 201086 239686
rect 201408 239672 201566 239700
rect 201792 239672 202046 239700
rect 202176 239672 202430 239700
rect 201538 233761 201566 239672
rect 202018 234575 202046 239672
rect 202006 234569 202058 234575
rect 202006 234511 202058 234517
rect 201526 233755 201578 233761
rect 201526 233697 201578 233703
rect 201334 233681 201386 233687
rect 201334 233623 201386 233629
rect 201046 233607 201098 233613
rect 201046 233549 201098 233555
rect 200662 233533 200714 233539
rect 200662 233475 200714 233481
rect 201346 221482 201374 233623
rect 202402 233317 202430 239672
rect 202498 233687 202526 239686
rect 202882 234723 202910 239686
rect 202870 234717 202922 234723
rect 202870 234659 202922 234665
rect 203266 234501 203294 239686
rect 203712 239672 203966 239700
rect 204096 239672 204254 239700
rect 203254 234495 203306 234501
rect 203254 234437 203306 234443
rect 202870 233829 202922 233835
rect 202870 233771 202922 233777
rect 202486 233681 202538 233687
rect 202486 233623 202538 233629
rect 202102 233311 202154 233317
rect 202102 233253 202154 233259
rect 202390 233311 202442 233317
rect 202390 233253 202442 233259
rect 202114 221792 202142 233253
rect 202114 221764 202190 221792
rect 202162 221482 202190 221764
rect 202882 221482 202910 233771
rect 203938 233391 203966 239672
rect 204226 233835 204254 239672
rect 204418 239672 204480 239700
rect 204418 234797 204446 239672
rect 204406 234791 204458 234797
rect 204406 234733 204458 234739
rect 204802 234649 204830 239686
rect 204790 234643 204842 234649
rect 204790 234585 204842 234591
rect 204310 233977 204362 233983
rect 204310 233919 204362 233925
rect 204214 233829 204266 233835
rect 204214 233771 204266 233777
rect 203638 233385 203690 233391
rect 203638 233327 203690 233333
rect 203926 233385 203978 233391
rect 203926 233327 203978 233333
rect 203650 221482 203678 233327
rect 204322 221792 204350 233919
rect 205186 233909 205214 239686
rect 205570 233983 205598 239686
rect 205920 239672 206174 239700
rect 206304 239672 206558 239700
rect 206688 239672 206942 239700
rect 206146 234427 206174 239672
rect 206134 234421 206186 234427
rect 206134 234363 206186 234369
rect 206530 234353 206558 239672
rect 206518 234347 206570 234353
rect 206518 234289 206570 234295
rect 205942 234051 205994 234057
rect 205942 233993 205994 233999
rect 205558 233977 205610 233983
rect 205558 233919 205610 233925
rect 205078 233903 205130 233909
rect 205078 233845 205130 233851
rect 205174 233903 205226 233909
rect 205174 233845 205226 233851
rect 204322 221764 204398 221792
rect 204370 221482 204398 221764
rect 205090 221482 205118 233845
rect 205954 221496 205982 233993
rect 206914 233983 206942 239672
rect 207010 235389 207038 239686
rect 207490 235981 207518 239686
rect 207478 235975 207530 235981
rect 207478 235917 207530 235923
rect 206998 235383 207050 235389
rect 206998 235325 207050 235331
rect 207874 235093 207902 239686
rect 208224 239672 208478 239700
rect 208608 239672 208766 239700
rect 208450 236055 208478 239672
rect 208438 236049 208490 236055
rect 208438 235991 208490 235997
rect 207862 235087 207914 235093
rect 207862 235029 207914 235035
rect 208738 234871 208766 239672
rect 208930 235833 208958 239686
rect 208918 235827 208970 235833
rect 208918 235769 208970 235775
rect 209314 235241 209342 239686
rect 209698 235907 209726 239686
rect 209686 235901 209738 235907
rect 209686 235843 209738 235849
rect 210082 235611 210110 239686
rect 210432 239672 210686 239700
rect 210816 239672 211070 239700
rect 210658 235685 210686 239672
rect 210646 235679 210698 235685
rect 210646 235621 210698 235627
rect 210070 235605 210122 235611
rect 210070 235547 210122 235553
rect 209302 235235 209354 235241
rect 209302 235177 209354 235183
rect 211042 235019 211070 239672
rect 211234 235759 211262 239686
rect 211222 235753 211274 235759
rect 211222 235695 211274 235701
rect 211618 235167 211646 239686
rect 212002 235463 212030 239686
rect 211990 235457 212042 235463
rect 211990 235399 212042 235405
rect 211606 235161 211658 235167
rect 211606 235103 211658 235109
rect 211030 235013 211082 235019
rect 211030 234955 211082 234961
rect 208726 234865 208778 234871
rect 208726 234807 208778 234813
rect 207766 234495 207818 234501
rect 207766 234437 207818 234443
rect 207778 234131 207806 234437
rect 210358 234273 210410 234279
rect 210358 234215 210410 234221
rect 208822 234199 208874 234205
rect 208822 234141 208874 234147
rect 207382 234125 207434 234131
rect 207382 234067 207434 234073
rect 207766 234125 207818 234131
rect 207766 234067 207818 234073
rect 206902 233977 206954 233983
rect 206902 233919 206954 233925
rect 206614 233459 206666 233465
rect 206614 233401 206666 233407
rect 205920 221468 205982 221496
rect 206626 221496 206654 233401
rect 206626 221468 206688 221496
rect 207394 221482 207422 234067
rect 208150 233533 208202 233539
rect 208150 233475 208202 233481
rect 208162 221496 208190 233475
rect 208128 221468 208190 221496
rect 208834 221496 208862 234141
rect 209686 233607 209738 233613
rect 209686 233549 209738 233555
rect 208834 221468 208896 221496
rect 209698 221482 209726 233549
rect 210370 221792 210398 234215
rect 211894 233755 211946 233761
rect 211894 233697 211946 233703
rect 211126 233311 211178 233317
rect 211126 233253 211178 233259
rect 210370 221764 210446 221792
rect 210418 221482 210446 221764
rect 211138 221482 211166 233253
rect 211906 221482 211934 233697
rect 212386 225991 212414 239686
rect 212736 239672 212990 239700
rect 212962 235537 212990 239672
rect 213058 239672 213120 239700
rect 212950 235531 213002 235537
rect 212950 235473 213002 235479
rect 212566 233681 212618 233687
rect 212566 233623 212618 233629
rect 212374 225985 212426 225991
rect 212374 225927 212426 225933
rect 212578 221792 212606 233623
rect 213058 227471 213086 239672
rect 213442 234945 213470 239686
rect 213430 234939 213482 234945
rect 213430 234881 213482 234887
rect 213430 234569 213482 234575
rect 213430 234511 213482 234517
rect 213046 227465 213098 227471
rect 213046 227407 213098 227413
rect 212578 221764 212654 221792
rect 212626 221482 212654 221764
rect 213442 221482 213470 234511
rect 213826 226361 213854 239686
rect 214210 235315 214238 239686
rect 214198 235309 214250 235315
rect 214198 235251 214250 235257
rect 214198 233385 214250 233391
rect 214198 233327 214250 233333
rect 213814 226355 213866 226361
rect 213814 226297 213866 226303
rect 214210 221482 214238 233327
rect 214594 226065 214622 239686
rect 215040 239672 215294 239700
rect 215424 239672 215678 239700
rect 214870 234717 214922 234723
rect 214870 234659 214922 234665
rect 214582 226059 214634 226065
rect 214582 226001 214634 226007
rect 214882 221792 214910 234659
rect 215266 229691 215294 239672
rect 215542 233829 215594 233835
rect 215542 233771 215594 233777
rect 215254 229685 215306 229691
rect 215254 229627 215306 229633
rect 215554 226084 215582 233771
rect 215650 226213 215678 239672
rect 215746 227101 215774 239686
rect 215926 235087 215978 235093
rect 215926 235029 215978 235035
rect 215830 234791 215882 234797
rect 215830 234733 215882 234739
rect 215842 233835 215870 234733
rect 215938 234501 215966 235029
rect 215926 234495 215978 234501
rect 215926 234437 215978 234443
rect 215830 233829 215882 233835
rect 215830 233771 215882 233777
rect 216130 227545 216158 239686
rect 216514 236174 216542 239686
rect 216864 239672 217118 239700
rect 217248 239672 217502 239700
rect 217632 239672 217886 239700
rect 216514 236146 216638 236174
rect 216502 234125 216554 234131
rect 216502 234067 216554 234073
rect 216118 227539 216170 227545
rect 216118 227481 216170 227487
rect 215734 227095 215786 227101
rect 215734 227037 215786 227043
rect 215638 226207 215690 226213
rect 215638 226149 215690 226155
rect 215554 226056 215678 226084
rect 214882 221764 214958 221792
rect 214930 221482 214958 221764
rect 215650 221482 215678 226056
rect 216514 221482 216542 234067
rect 216610 232799 216638 236146
rect 216598 232793 216650 232799
rect 216598 232735 216650 232741
rect 217090 226287 217118 239672
rect 217174 233681 217226 233687
rect 217174 233623 217226 233629
rect 217078 226281 217130 226287
rect 217078 226223 217130 226229
rect 217186 221792 217214 233623
rect 217474 227397 217502 239672
rect 217462 227391 217514 227397
rect 217462 227333 217514 227339
rect 217858 227249 217886 239672
rect 217954 236174 217982 239686
rect 217954 236146 218078 236174
rect 217942 233829 217994 233835
rect 217942 233771 217994 233777
rect 217846 227243 217898 227249
rect 217846 227185 217898 227191
rect 217186 221764 217262 221792
rect 217234 221482 217262 221764
rect 217954 221482 217982 233771
rect 218050 232651 218078 236146
rect 218038 232645 218090 232651
rect 218038 232587 218090 232593
rect 218338 226139 218366 239686
rect 218710 234051 218762 234057
rect 218710 233993 218762 233999
rect 218326 226133 218378 226139
rect 218326 226075 218378 226081
rect 218722 221482 218750 233993
rect 218818 225917 218846 239686
rect 219168 239672 219422 239700
rect 219552 239672 219806 239700
rect 219936 239672 220190 239700
rect 219394 236174 219422 239672
rect 219394 236146 219518 236174
rect 219382 234421 219434 234427
rect 219382 234363 219434 234369
rect 218806 225911 218858 225917
rect 218806 225853 218858 225859
rect 219394 221792 219422 234363
rect 219490 227323 219518 236146
rect 219778 232577 219806 239672
rect 219766 232571 219818 232577
rect 219766 232513 219818 232519
rect 220162 229617 220190 239672
rect 220258 236174 220286 239686
rect 220258 236146 220382 236174
rect 220246 233977 220298 233983
rect 220246 233919 220298 233925
rect 220150 229611 220202 229617
rect 220150 229553 220202 229559
rect 219478 227317 219530 227323
rect 219478 227259 219530 227265
rect 219394 221764 219470 221792
rect 219442 221482 219470 221764
rect 220258 221482 220286 233919
rect 220354 227175 220382 236146
rect 220642 235093 220670 239686
rect 221026 236174 221054 239686
rect 221376 239672 221630 239700
rect 221026 236146 221150 236174
rect 220630 235087 220682 235093
rect 220630 235029 220682 235035
rect 221014 234347 221066 234353
rect 221014 234289 221066 234295
rect 220342 227169 220394 227175
rect 220342 227111 220394 227117
rect 221026 221482 221054 234289
rect 221122 232503 221150 236146
rect 221110 232497 221162 232503
rect 221110 232439 221162 232445
rect 221602 229543 221630 239672
rect 221746 239404 221774 239686
rect 222144 239672 222398 239700
rect 221698 239376 221774 239404
rect 221590 229537 221642 229543
rect 221590 229479 221642 229485
rect 221698 226953 221726 239376
rect 221782 235383 221834 235389
rect 221782 235325 221834 235331
rect 221686 226947 221738 226953
rect 221686 226889 221738 226895
rect 221794 221792 221822 235325
rect 222370 234649 222398 239672
rect 222358 234643 222410 234649
rect 222358 234585 222410 234591
rect 222454 234273 222506 234279
rect 222454 234215 222506 234221
rect 221746 221764 221822 221792
rect 221746 221482 221774 221764
rect 222466 221482 222494 234215
rect 222562 232429 222590 239686
rect 222550 232423 222602 232429
rect 222550 232365 222602 232371
rect 222946 232355 222974 239686
rect 223222 236049 223274 236055
rect 223222 235991 223274 235997
rect 222934 232349 222986 232355
rect 222934 232291 222986 232297
rect 223234 221482 223262 235991
rect 223330 226805 223358 239686
rect 223680 239672 223934 239700
rect 224064 239672 224318 239700
rect 223906 235389 223934 239672
rect 223990 235975 224042 235981
rect 223990 235917 224042 235923
rect 223894 235383 223946 235389
rect 223894 235325 223946 235331
rect 223318 226799 223370 226805
rect 223318 226741 223370 226747
rect 224002 221792 224030 235917
rect 224290 232281 224318 239672
rect 224278 232275 224330 232281
rect 224278 232217 224330 232223
rect 224386 228507 224414 239686
rect 224784 239672 224990 239700
rect 224758 234865 224810 234871
rect 224758 234807 224810 234813
rect 224374 228501 224426 228507
rect 224374 228443 224426 228449
rect 224002 221764 224078 221792
rect 224050 221482 224078 221764
rect 224770 221482 224798 234807
rect 224962 226879 224990 239672
rect 225154 234723 225182 239686
rect 225538 234871 225566 239686
rect 225984 239672 226238 239700
rect 226368 239672 226622 239700
rect 226210 236174 226238 239672
rect 226210 236146 226334 236174
rect 226198 235901 226250 235907
rect 226198 235843 226250 235849
rect 225526 234865 225578 234871
rect 225526 234807 225578 234813
rect 225142 234717 225194 234723
rect 225142 234659 225194 234665
rect 225526 234495 225578 234501
rect 225526 234437 225578 234443
rect 224950 226873 225002 226879
rect 224950 226815 225002 226821
rect 225538 221482 225566 234437
rect 226210 221792 226238 235843
rect 226306 232207 226334 236146
rect 226294 232201 226346 232207
rect 226294 232143 226346 232149
rect 226594 226731 226622 239672
rect 226690 233391 226718 239686
rect 226966 235827 227018 235833
rect 226966 235769 227018 235775
rect 226678 233385 226730 233391
rect 226678 233327 226730 233333
rect 226582 226725 226634 226731
rect 226582 226667 226634 226673
rect 226210 221764 226286 221792
rect 226258 221482 226286 221764
rect 226978 221482 227006 235769
rect 227074 232133 227102 239686
rect 227062 232127 227114 232133
rect 227062 232069 227114 232075
rect 227458 229987 227486 239686
rect 227856 239672 227966 239700
rect 228192 239672 228446 239700
rect 228576 239672 228830 239700
rect 227830 235605 227882 235611
rect 227830 235547 227882 235553
rect 227446 229981 227498 229987
rect 227446 229923 227498 229929
rect 227842 221482 227870 235547
rect 227938 226657 227966 239672
rect 228418 233613 228446 239672
rect 228502 235235 228554 235241
rect 228502 235177 228554 235183
rect 228406 233607 228458 233613
rect 228406 233549 228458 233555
rect 227926 226651 227978 226657
rect 227926 226593 227978 226599
rect 228514 221792 228542 235177
rect 228802 228581 228830 239672
rect 228898 228729 228926 239686
rect 229296 239672 229598 239700
rect 229270 235753 229322 235759
rect 229270 235695 229322 235701
rect 228886 228723 228938 228729
rect 228886 228665 228938 228671
rect 228790 228575 228842 228581
rect 228790 228517 228842 228523
rect 228514 221764 228590 221792
rect 228562 221482 228590 221764
rect 229282 221482 229310 235695
rect 229570 226583 229598 239672
rect 229762 235241 229790 239686
rect 230112 239672 230366 239700
rect 230496 239672 230654 239700
rect 230880 239672 231134 239700
rect 230038 235679 230090 235685
rect 230038 235621 230090 235627
rect 229750 235235 229802 235241
rect 229750 235177 229802 235183
rect 229558 226577 229610 226583
rect 229558 226519 229610 226525
rect 230050 221482 230078 235621
rect 230338 229395 230366 239672
rect 230326 229389 230378 229395
rect 230326 229331 230378 229337
rect 230626 228655 230654 239672
rect 230710 235161 230762 235167
rect 230710 235103 230762 235109
rect 230614 228649 230666 228655
rect 230614 228591 230666 228597
rect 230722 221792 230750 235103
rect 231106 226509 231134 239672
rect 231202 235759 231230 239686
rect 231600 239672 231902 239700
rect 231190 235753 231242 235759
rect 231190 235695 231242 235701
rect 231574 235013 231626 235019
rect 231574 234955 231626 234961
rect 231094 226503 231146 226509
rect 231094 226445 231146 226451
rect 230722 221764 230798 221792
rect 230770 221482 230798 221764
rect 231586 221482 231614 234955
rect 231874 229321 231902 239672
rect 231862 229315 231914 229321
rect 231862 229257 231914 229263
rect 231970 229173 231998 239686
rect 232320 239672 232574 239700
rect 232704 239672 232958 239700
rect 233088 239672 233246 239700
rect 232342 235531 232394 235537
rect 232342 235473 232394 235479
rect 231958 229167 232010 229173
rect 231958 229109 232010 229115
rect 232354 221482 232382 235473
rect 232546 226435 232574 239672
rect 232930 235167 232958 239672
rect 233014 235457 233066 235463
rect 233014 235399 233066 235405
rect 232918 235161 232970 235167
rect 232918 235103 232970 235109
rect 232534 226429 232586 226435
rect 232534 226371 232586 226377
rect 233026 221792 233054 235399
rect 233218 231911 233246 239672
rect 233206 231905 233258 231911
rect 233206 231847 233258 231853
rect 233506 229247 233534 239686
rect 233890 232059 233918 239686
rect 234274 235907 234302 239686
rect 234624 239672 234878 239700
rect 235008 239672 235262 239700
rect 235392 239672 235646 239700
rect 234262 235901 234314 235907
rect 234262 235843 234314 235849
rect 233878 232053 233930 232059
rect 233878 231995 233930 232001
rect 234850 231985 234878 239672
rect 234838 231979 234890 231985
rect 234838 231921 234890 231927
rect 233494 229241 233546 229247
rect 233494 229183 233546 229189
rect 235234 229025 235262 239672
rect 235318 235309 235370 235315
rect 235318 235251 235370 235257
rect 235222 229019 235274 229025
rect 235222 228961 235274 228967
rect 233782 227465 233834 227471
rect 233782 227407 233834 227413
rect 233026 221764 233102 221792
rect 233074 221482 233102 221764
rect 233794 221482 233822 227407
rect 234550 225985 234602 225991
rect 234550 225927 234602 225933
rect 234562 221482 234590 225927
rect 235330 221496 235358 235251
rect 235618 234501 235646 239672
rect 235714 234945 235742 239686
rect 236002 239672 236112 239700
rect 235702 234939 235754 234945
rect 235702 234881 235754 234887
rect 235606 234495 235658 234501
rect 235606 234437 235658 234443
rect 236002 231837 236030 239672
rect 236482 235611 236510 239686
rect 236832 239672 237086 239700
rect 237312 239672 237566 239700
rect 236470 235605 236522 235611
rect 236470 235547 236522 235553
rect 236086 234791 236138 234797
rect 236086 234733 236138 234739
rect 235990 231831 236042 231837
rect 235990 231773 236042 231779
rect 235330 221468 235392 221496
rect 236098 221482 236126 234733
rect 237058 234427 237086 239672
rect 237538 235833 237566 239672
rect 237526 235827 237578 235833
rect 237526 235769 237578 235775
rect 237046 234421 237098 234427
rect 237046 234363 237098 234369
rect 236758 233385 236810 233391
rect 236758 233327 236810 233333
rect 236770 225991 236798 233327
rect 237634 232725 237662 239686
rect 238018 235537 238046 239686
rect 238006 235531 238058 235537
rect 238006 235473 238058 235479
rect 238102 233607 238154 233613
rect 238102 233549 238154 233555
rect 237622 232719 237674 232725
rect 237622 232661 237674 232667
rect 238114 227027 238142 233549
rect 238402 229099 238430 239686
rect 238390 229093 238442 229099
rect 238390 229035 238442 229041
rect 238786 227471 238814 239686
rect 239136 239672 239390 239700
rect 239520 239672 239774 239700
rect 239362 235685 239390 239672
rect 239350 235679 239402 235685
rect 239350 235621 239402 235627
rect 239062 229685 239114 229691
rect 239062 229627 239114 229633
rect 238774 227465 238826 227471
rect 238774 227407 238826 227413
rect 238390 227095 238442 227101
rect 238390 227037 238442 227043
rect 238102 227021 238154 227027
rect 238102 226963 238154 226969
rect 237526 226355 237578 226361
rect 237526 226297 237578 226303
rect 236854 226059 236906 226065
rect 236854 226001 236906 226007
rect 236758 225985 236810 225991
rect 236758 225927 236810 225933
rect 236866 221496 236894 226001
rect 236832 221468 236894 221496
rect 237538 221496 237566 226297
rect 237538 221468 237600 221496
rect 238402 221482 238430 227037
rect 239074 221792 239102 229627
rect 239746 228803 239774 239672
rect 239842 234353 239870 239686
rect 240226 234649 240254 239686
rect 240214 234643 240266 234649
rect 240214 234585 240266 234591
rect 239830 234347 239882 234353
rect 239830 234289 239882 234295
rect 240610 233539 240638 239686
rect 240598 233533 240650 233539
rect 240598 233475 240650 233481
rect 241090 230357 241118 239686
rect 241440 239672 241694 239700
rect 241078 230351 241130 230357
rect 241078 230293 241130 230299
rect 241666 228877 241694 239672
rect 241762 239672 241824 239700
rect 241654 228871 241706 228877
rect 241654 228813 241706 228819
rect 239734 228797 239786 228803
rect 239734 228739 239786 228745
rect 239830 227539 239882 227545
rect 239830 227481 239882 227487
rect 239074 221764 239150 221792
rect 239122 221482 239150 221764
rect 239842 221482 239870 227481
rect 241270 227391 241322 227397
rect 241270 227333 241322 227339
rect 240598 226207 240650 226213
rect 240598 226149 240650 226155
rect 240610 221482 240638 226149
rect 241282 221792 241310 227333
rect 241762 225843 241790 239672
rect 242146 235463 242174 239686
rect 242134 235457 242186 235463
rect 242134 235399 242186 235405
rect 241846 235087 241898 235093
rect 241846 235029 241898 235035
rect 241858 226065 241886 235029
rect 242134 232793 242186 232799
rect 242134 232735 242186 232741
rect 241846 226059 241898 226065
rect 241846 226001 241898 226007
rect 241750 225837 241802 225843
rect 241750 225779 241802 225785
rect 241282 221764 241358 221792
rect 241330 221482 241358 221764
rect 242146 221482 242174 232735
rect 242530 228951 242558 239686
rect 242914 234279 242942 239686
rect 243298 235981 243326 239686
rect 243648 239672 243902 239700
rect 244032 239672 244286 239700
rect 243286 235975 243338 235981
rect 243286 235917 243338 235923
rect 243874 235019 243902 239672
rect 243862 235013 243914 235019
rect 243862 234955 243914 234961
rect 243958 234569 244010 234575
rect 243958 234511 244010 234517
rect 242902 234273 242954 234279
rect 242902 234215 242954 234221
rect 242518 228945 242570 228951
rect 242518 228887 242570 228893
rect 242902 227243 242954 227249
rect 242902 227185 242954 227191
rect 242914 221482 242942 227185
rect 243574 226281 243626 226287
rect 243574 226223 243626 226229
rect 243586 221792 243614 226223
rect 243970 226213 243998 234511
rect 244258 229691 244286 239672
rect 244354 234131 244382 239686
rect 244726 235383 244778 235389
rect 244726 235325 244778 235331
rect 244342 234125 244394 234131
rect 244342 234067 244394 234073
rect 244246 229685 244298 229691
rect 244246 229627 244298 229633
rect 244738 227397 244766 235325
rect 244726 227391 244778 227397
rect 244726 227333 244778 227339
rect 244834 226361 244862 239686
rect 245110 232645 245162 232651
rect 245110 232587 245162 232593
rect 244822 226355 244874 226361
rect 244822 226297 244874 226303
rect 243958 226207 244010 226213
rect 243958 226149 244010 226155
rect 244342 225911 244394 225917
rect 244342 225853 244394 225859
rect 243586 221764 243662 221792
rect 243634 221482 243662 221764
rect 244354 221482 244382 225853
rect 245122 221482 245150 232587
rect 245218 231319 245246 239686
rect 245568 239672 245822 239700
rect 245952 239672 246206 239700
rect 246336 239672 246590 239700
rect 245206 231313 245258 231319
rect 245206 231255 245258 231261
rect 245794 230283 245822 239672
rect 246178 230431 246206 239672
rect 246166 230425 246218 230431
rect 246166 230367 246218 230373
rect 245782 230277 245834 230283
rect 245782 230219 245834 230225
rect 245878 227317 245930 227323
rect 245878 227259 245930 227265
rect 245890 221792 245918 227259
rect 246562 226287 246590 239672
rect 246658 235093 246686 239686
rect 246646 235087 246698 235093
rect 246646 235029 246698 235035
rect 247042 227767 247070 239686
rect 247426 234057 247454 239686
rect 247776 239672 248030 239700
rect 248160 239672 248414 239700
rect 248640 239672 248798 239700
rect 248002 236055 248030 239672
rect 247990 236049 248042 236055
rect 247990 235991 248042 235997
rect 247702 234717 247754 234723
rect 247702 234659 247754 234665
rect 247414 234051 247466 234057
rect 247414 233993 247466 233999
rect 247030 227761 247082 227767
rect 247030 227703 247082 227709
rect 247414 227169 247466 227175
rect 247414 227111 247466 227117
rect 246550 226281 246602 226287
rect 246550 226223 246602 226229
rect 246646 226133 246698 226139
rect 246646 226075 246698 226081
rect 245890 221764 245966 221792
rect 245938 221482 245966 221764
rect 246658 221482 246686 226075
rect 247426 221482 247454 227111
rect 247714 225769 247742 234659
rect 248086 232571 248138 232577
rect 248086 232513 248138 232519
rect 247702 225763 247754 225769
rect 247702 225705 247754 225711
rect 248098 221792 248126 232513
rect 248386 231541 248414 239672
rect 248374 231535 248426 231541
rect 248374 231477 248426 231483
rect 248770 230061 248798 239672
rect 248962 230209 248990 239686
rect 248950 230203 249002 230209
rect 248950 230145 249002 230151
rect 248758 230055 248810 230061
rect 248758 229997 248810 230003
rect 249346 227545 249374 239686
rect 249730 235389 249758 239686
rect 250080 239672 250238 239700
rect 249718 235383 249770 235389
rect 249718 235325 249770 235331
rect 250210 229913 250238 239672
rect 250450 239404 250478 239686
rect 250848 239672 251102 239700
rect 250450 239376 250526 239404
rect 250498 234501 250526 239376
rect 251074 236129 251102 239672
rect 251062 236123 251114 236129
rect 251062 236065 251114 236071
rect 251170 234723 251198 239686
rect 251158 234717 251210 234723
rect 251158 234659 251210 234665
rect 250582 234569 250634 234575
rect 250582 234511 250634 234517
rect 250486 234495 250538 234501
rect 250486 234437 250538 234443
rect 250198 229907 250250 229913
rect 250198 229849 250250 229855
rect 249718 229611 249770 229617
rect 249718 229553 249770 229559
rect 249334 227539 249386 227545
rect 249334 227481 249386 227487
rect 248854 226059 248906 226065
rect 248854 226001 248906 226007
rect 248098 221764 248174 221792
rect 248146 221482 248174 221764
rect 248866 221482 248894 226001
rect 249730 221482 249758 229553
rect 250594 228433 250622 234511
rect 251158 232497 251210 232503
rect 251158 232439 251210 232445
rect 250582 228427 250634 228433
rect 250582 228369 250634 228375
rect 250390 226947 250442 226953
rect 250390 226889 250442 226895
rect 250402 221792 250430 226889
rect 250402 221764 250478 221792
rect 250450 221482 250478 221764
rect 251170 221482 251198 232439
rect 251554 229839 251582 239686
rect 251938 230135 251966 239686
rect 252384 239672 252638 239700
rect 252768 239672 253022 239700
rect 252610 236174 252638 239672
rect 252610 236146 252734 236174
rect 251926 230129 251978 230135
rect 251926 230071 251978 230077
rect 251542 229833 251594 229839
rect 251542 229775 251594 229781
rect 252598 229537 252650 229543
rect 252598 229479 252650 229485
rect 252214 227465 252266 227471
rect 252214 227407 252266 227413
rect 252226 226361 252254 227407
rect 252214 226355 252266 226361
rect 252214 226297 252266 226303
rect 251926 226207 251978 226213
rect 251926 226149 251978 226155
rect 252118 226207 252170 226213
rect 252118 226149 252170 226155
rect 251938 221482 251966 226149
rect 252130 225843 252158 226149
rect 252118 225837 252170 225843
rect 252118 225779 252170 225785
rect 252610 221792 252638 229479
rect 252706 225103 252734 236146
rect 252994 231097 253022 239672
rect 252982 231091 253034 231097
rect 252982 231033 253034 231039
rect 253090 229617 253118 239686
rect 253474 233835 253502 239686
rect 253558 235235 253610 235241
rect 253558 235177 253610 235183
rect 253462 233829 253514 233835
rect 253462 233771 253514 233777
rect 253078 229611 253130 229617
rect 253078 229553 253130 229559
rect 253570 226953 253598 235177
rect 253858 227471 253886 239686
rect 254242 234797 254270 239686
rect 254592 239672 254846 239700
rect 254976 239672 255230 239700
rect 254230 234791 254282 234797
rect 254230 234733 254282 234739
rect 254230 232423 254282 232429
rect 254230 232365 254282 232371
rect 253846 227465 253898 227471
rect 253846 227407 253898 227413
rect 253558 226947 253610 226953
rect 253558 226889 253610 226895
rect 253462 226799 253514 226805
rect 253462 226741 253514 226747
rect 252694 225097 252746 225103
rect 252694 225039 252746 225045
rect 252610 221764 252686 221792
rect 252658 221482 252686 221764
rect 253474 221482 253502 226741
rect 254242 221482 254270 232365
rect 254818 229765 254846 239672
rect 254806 229759 254858 229765
rect 254806 229701 254858 229707
rect 255202 229543 255230 239672
rect 255298 234575 255326 239686
rect 255286 234569 255338 234575
rect 255286 234511 255338 234517
rect 255670 232349 255722 232355
rect 255670 232291 255722 232297
rect 255190 229537 255242 229543
rect 255190 229479 255242 229485
rect 254902 227391 254954 227397
rect 254902 227333 254954 227339
rect 254914 221792 254942 227333
rect 254914 221764 254990 221792
rect 254962 221482 254990 221764
rect 255682 221482 255710 232291
rect 255778 231689 255806 239686
rect 255766 231683 255818 231689
rect 255766 231625 255818 231631
rect 256162 231171 256190 239686
rect 256546 234205 256574 239686
rect 256896 239672 257150 239700
rect 257280 239672 257534 239700
rect 256534 234199 256586 234205
rect 256534 234141 256586 234147
rect 256150 231165 256202 231171
rect 256150 231107 256202 231113
rect 256438 226873 256490 226879
rect 256438 226815 256490 226821
rect 256450 221482 256478 226815
rect 257122 226065 257150 239672
rect 257506 235241 257534 239672
rect 257494 235235 257546 235241
rect 257494 235177 257546 235183
rect 257206 232275 257258 232281
rect 257206 232217 257258 232223
rect 257110 226059 257162 226065
rect 257110 226001 257162 226007
rect 257218 221792 257246 232217
rect 257602 231615 257630 239686
rect 257986 233317 258014 239686
rect 258070 234421 258122 234427
rect 258070 234363 258122 234369
rect 257974 233311 258026 233317
rect 257974 233253 258026 233259
rect 257590 231609 257642 231615
rect 257590 231551 257642 231557
rect 258082 228063 258110 234363
rect 258370 233909 258398 239686
rect 258358 233903 258410 233909
rect 258358 233845 258410 233851
rect 258754 231763 258782 239686
rect 259104 239672 259166 239700
rect 259584 239672 259838 239700
rect 259030 235753 259082 235759
rect 259030 235695 259082 235701
rect 258742 231757 258794 231763
rect 258742 231699 258794 231705
rect 258742 228501 258794 228507
rect 258742 228443 258794 228449
rect 258070 228057 258122 228063
rect 258070 227999 258122 228005
rect 257974 225763 258026 225769
rect 257974 225705 258026 225711
rect 257218 221764 257294 221792
rect 257266 221482 257294 221764
rect 257986 221482 258014 225705
rect 258754 221482 258782 228443
rect 259042 225473 259070 235695
rect 259138 233243 259166 239672
rect 259810 233983 259838 239672
rect 259798 233977 259850 233983
rect 259798 233919 259850 233925
rect 259906 233613 259934 239686
rect 260290 234871 260318 239686
rect 260182 234865 260234 234871
rect 260182 234807 260234 234813
rect 260278 234865 260330 234871
rect 260278 234807 260330 234813
rect 259894 233607 259946 233613
rect 259894 233549 259946 233555
rect 259126 233237 259178 233243
rect 259126 233179 259178 233185
rect 259414 226725 259466 226731
rect 259414 226667 259466 226673
rect 259030 225467 259082 225473
rect 259030 225409 259082 225415
rect 259426 221792 259454 226667
rect 259426 221764 259502 221792
rect 259474 221482 259502 221764
rect 260194 221482 260222 234807
rect 260470 234347 260522 234353
rect 260470 234289 260522 234295
rect 260482 228507 260510 234289
rect 260674 233021 260702 239686
rect 261024 239672 261278 239700
rect 261408 239672 261662 239700
rect 261792 239672 261950 239700
rect 261250 234279 261278 239672
rect 260758 234273 260810 234279
rect 260758 234215 260810 234221
rect 261238 234273 261290 234279
rect 261238 234215 261290 234221
rect 260662 233015 260714 233021
rect 260662 232957 260714 232963
rect 260470 228501 260522 228507
rect 260470 228443 260522 228449
rect 260770 228359 260798 234215
rect 261634 233391 261662 239672
rect 261622 233385 261674 233391
rect 261622 233327 261674 233333
rect 261718 232201 261770 232207
rect 261718 232143 261770 232149
rect 260758 228353 260810 228359
rect 260758 228295 260810 228301
rect 261046 225985 261098 225991
rect 261046 225927 261098 225933
rect 261058 221482 261086 225927
rect 261730 221792 261758 232143
rect 261922 223771 261950 239672
rect 262006 235161 262058 235167
rect 262006 235103 262058 235109
rect 262018 225917 262046 235103
rect 262114 233169 262142 239686
rect 262498 234427 262526 239686
rect 262882 235759 262910 239686
rect 263328 239672 263582 239700
rect 263712 239672 263966 239700
rect 264096 239672 264350 239700
rect 262870 235753 262922 235759
rect 262870 235695 262922 235701
rect 262486 234421 262538 234427
rect 262486 234363 262538 234369
rect 262102 233163 262154 233169
rect 262102 233105 262154 233111
rect 263254 232127 263306 232133
rect 263254 232069 263306 232075
rect 262486 226651 262538 226657
rect 262486 226593 262538 226599
rect 262006 225911 262058 225917
rect 262006 225853 262058 225859
rect 261910 223765 261962 223771
rect 261910 223707 261962 223713
rect 261730 221764 261806 221792
rect 261778 221482 261806 221764
rect 262498 221482 262526 226593
rect 263266 221482 263294 232069
rect 263554 223697 263582 239672
rect 263830 234125 263882 234131
rect 263830 234067 263882 234073
rect 263842 227989 263870 234067
rect 263938 232873 263966 239672
rect 263926 232867 263978 232873
rect 263926 232809 263978 232815
rect 264322 229469 264350 239672
rect 264418 233465 264446 239686
rect 264610 239672 264816 239700
rect 264406 233459 264458 233465
rect 264406 233401 264458 233407
rect 264310 229463 264362 229469
rect 264310 229405 264362 229411
rect 263830 227983 263882 227989
rect 263830 227925 263882 227931
rect 264022 227021 264074 227027
rect 264022 226963 264074 226969
rect 263542 223691 263594 223697
rect 263542 223633 263594 223639
rect 264034 221496 264062 226963
rect 264610 223475 264638 239672
rect 264886 235901 264938 235907
rect 264886 235843 264938 235849
rect 264694 234643 264746 234649
rect 264694 234585 264746 234591
rect 264706 227175 264734 234585
rect 264790 229981 264842 229987
rect 264790 229923 264842 229929
rect 264694 227169 264746 227175
rect 264694 227111 264746 227117
rect 264598 223469 264650 223475
rect 264598 223411 264650 223417
rect 264034 221468 264096 221496
rect 264802 221482 264830 229923
rect 264898 226657 264926 235843
rect 265186 232799 265214 239686
rect 265536 239672 265790 239700
rect 265920 239672 266174 239700
rect 266304 239672 266558 239700
rect 265762 233095 265790 239672
rect 266146 235167 266174 239672
rect 266134 235161 266186 235167
rect 266134 235103 266186 235109
rect 266326 234051 266378 234057
rect 266326 233993 266378 233999
rect 265750 233089 265802 233095
rect 265750 233031 265802 233037
rect 265174 232793 265226 232799
rect 265174 232735 265226 232741
rect 266338 228581 266366 233993
rect 266230 228575 266282 228581
rect 266230 228517 266282 228523
rect 266326 228575 266378 228581
rect 266326 228517 266378 228523
rect 264886 226651 264938 226657
rect 264886 226593 264938 226599
rect 265558 226577 265610 226583
rect 265558 226519 265610 226525
rect 265570 221496 265598 226519
rect 265536 221468 265598 221496
rect 266242 221496 266270 228517
rect 266530 223549 266558 239672
rect 266626 232577 266654 239686
rect 266902 234939 266954 234945
rect 266902 234881 266954 234887
rect 266614 232571 266666 232577
rect 266614 232513 266666 232519
rect 266914 226065 266942 234881
rect 267106 234057 267134 239686
rect 267490 234649 267518 239686
rect 267840 239672 268094 239700
rect 268224 239672 268478 239700
rect 267478 234643 267530 234649
rect 267478 234585 267530 234591
rect 267958 234495 268010 234501
rect 267958 234437 268010 234443
rect 267094 234051 267146 234057
rect 267094 233993 267146 233999
rect 267766 233607 267818 233613
rect 267766 233549 267818 233555
rect 266998 226947 267050 226953
rect 266998 226889 267050 226895
rect 266902 226059 266954 226065
rect 266902 226001 266954 226007
rect 266518 223543 266570 223549
rect 266518 223485 266570 223491
rect 266242 221468 266304 221496
rect 267010 221482 267038 226889
rect 267778 225843 267806 233549
rect 267862 228723 267914 228729
rect 267862 228665 267914 228671
rect 267766 225837 267818 225843
rect 267766 225779 267818 225785
rect 267874 221792 267902 228665
rect 267970 228211 267998 234437
rect 267958 228205 268010 228211
rect 267958 228147 268010 228153
rect 268066 223623 268094 239672
rect 268450 232651 268478 239672
rect 268546 234131 268574 239686
rect 268630 235827 268682 235833
rect 268630 235769 268682 235775
rect 268534 234125 268586 234131
rect 268534 234067 268586 234073
rect 268438 232645 268490 232651
rect 268438 232587 268490 232593
rect 268534 226503 268586 226509
rect 268534 226445 268586 226451
rect 268054 223617 268106 223623
rect 268054 223559 268106 223565
rect 267826 221764 267902 221792
rect 267826 221482 267854 221764
rect 268546 221482 268574 226445
rect 268642 224733 268670 235769
rect 268930 234945 268958 239686
rect 269314 236174 269342 239686
rect 269314 236146 269438 236174
rect 268918 234939 268970 234945
rect 268918 234881 268970 234887
rect 269014 233385 269066 233391
rect 269014 233327 269066 233333
rect 269026 225769 269054 233327
rect 269302 229389 269354 229395
rect 269302 229331 269354 229337
rect 269014 225763 269066 225769
rect 269014 225705 269066 225711
rect 268630 224727 268682 224733
rect 268630 224669 268682 224675
rect 269314 221482 269342 229331
rect 269410 223327 269438 236146
rect 269494 233311 269546 233317
rect 269494 233253 269546 233259
rect 269506 228137 269534 233253
rect 269698 232355 269726 239686
rect 270048 239672 270302 239700
rect 270274 233317 270302 239672
rect 270418 239404 270446 239686
rect 270418 239376 270494 239404
rect 270466 233391 270494 239376
rect 270850 236174 270878 239686
rect 270850 236146 270974 236174
rect 270838 233829 270890 233835
rect 270838 233771 270890 233777
rect 270454 233385 270506 233391
rect 270454 233327 270506 233333
rect 270262 233311 270314 233317
rect 270262 233253 270314 233259
rect 269686 232349 269738 232355
rect 269686 232291 269738 232297
rect 270742 228649 270794 228655
rect 270742 228591 270794 228597
rect 269494 228131 269546 228137
rect 269494 228073 269546 228079
rect 269974 225467 270026 225473
rect 269974 225409 270026 225415
rect 269398 223321 269450 223327
rect 269398 223263 269450 223269
rect 269986 221792 270014 225409
rect 269986 221764 270062 221792
rect 270034 221482 270062 221764
rect 270754 221482 270782 228591
rect 270850 228285 270878 233771
rect 270838 228279 270890 228285
rect 270838 228221 270890 228227
rect 270946 223401 270974 236146
rect 271030 235975 271082 235981
rect 271030 235917 271082 235923
rect 271042 226583 271070 235917
rect 271234 232503 271262 239686
rect 271618 234353 271646 239686
rect 271606 234347 271658 234353
rect 271606 234289 271658 234295
rect 271222 232497 271274 232503
rect 271222 232439 271274 232445
rect 272002 227249 272030 239686
rect 272352 239672 272606 239700
rect 272736 239672 272990 239700
rect 272278 229315 272330 229321
rect 272278 229257 272330 229263
rect 271990 227243 272042 227249
rect 271990 227185 272042 227191
rect 271030 226577 271082 226583
rect 271030 226519 271082 226525
rect 271606 226429 271658 226435
rect 271606 226371 271658 226377
rect 270934 223395 270986 223401
rect 270934 223337 270986 223343
rect 271618 221482 271646 226371
rect 272290 221792 272318 229257
rect 272578 223253 272606 239672
rect 272854 233459 272906 233465
rect 272854 233401 272906 233407
rect 272866 226435 272894 233401
rect 272962 232207 272990 239672
rect 273058 234501 273086 239686
rect 273046 234495 273098 234501
rect 273046 234437 273098 234443
rect 272950 232201 273002 232207
rect 272950 232143 273002 232149
rect 273442 226953 273470 239686
rect 273840 239672 274142 239700
rect 273718 236123 273770 236129
rect 273718 236065 273770 236071
rect 273622 236049 273674 236055
rect 273622 235991 273674 235997
rect 273526 233311 273578 233317
rect 273526 233253 273578 233259
rect 273538 229395 273566 233253
rect 273526 229389 273578 229395
rect 273526 229331 273578 229337
rect 273430 226947 273482 226953
rect 273430 226889 273482 226895
rect 272854 226429 272906 226435
rect 272854 226371 272906 226377
rect 273046 225911 273098 225917
rect 273046 225853 273098 225859
rect 272566 223247 272618 223253
rect 272566 223189 272618 223195
rect 272290 221764 272366 221792
rect 272338 221482 272366 221764
rect 273058 221482 273086 225853
rect 273634 225547 273662 235991
rect 273730 225621 273758 236065
rect 273814 229167 273866 229173
rect 273814 229109 273866 229115
rect 273718 225615 273770 225621
rect 273718 225557 273770 225563
rect 273622 225541 273674 225547
rect 273622 225483 273674 225489
rect 273826 221482 273854 229109
rect 274114 222365 274142 239672
rect 274210 232281 274238 239686
rect 274656 239672 274910 239700
rect 275040 239672 275294 239700
rect 274882 232429 274910 239672
rect 275062 233385 275114 233391
rect 275062 233327 275114 233333
rect 274870 232423 274922 232429
rect 274870 232365 274922 232371
rect 274198 232275 274250 232281
rect 274198 232217 274250 232223
rect 274486 232053 274538 232059
rect 274486 231995 274538 232001
rect 274102 222359 274154 222365
rect 274102 222301 274154 222307
rect 274498 221792 274526 231995
rect 275074 227323 275102 233327
rect 275062 227317 275114 227323
rect 275062 227259 275114 227265
rect 275266 227027 275294 239672
rect 275362 237757 275390 239686
rect 275350 237751 275402 237757
rect 275350 237693 275402 237699
rect 275746 232059 275774 239686
rect 276130 236055 276158 239686
rect 276480 239672 276734 239700
rect 276864 239672 277118 239700
rect 277248 239672 277502 239700
rect 276118 236049 276170 236055
rect 276118 235991 276170 235997
rect 275734 232053 275786 232059
rect 275734 231995 275786 232001
rect 275350 231905 275402 231911
rect 275350 231847 275402 231853
rect 275254 227021 275306 227027
rect 275254 226963 275306 226969
rect 274498 221764 274574 221792
rect 274546 221482 274574 221764
rect 275362 221482 275390 231847
rect 276706 227101 276734 239672
rect 277090 237683 277118 239672
rect 277078 237677 277130 237683
rect 277078 237619 277130 237625
rect 277474 232133 277502 239672
rect 277570 236129 277598 239686
rect 277558 236123 277610 236129
rect 277558 236065 277610 236071
rect 277462 232127 277514 232133
rect 277462 232069 277514 232075
rect 276790 229241 276842 229247
rect 276790 229183 276842 229189
rect 276694 227095 276746 227101
rect 276694 227037 276746 227043
rect 276118 226651 276170 226657
rect 276118 226593 276170 226599
rect 276130 221482 276158 226593
rect 276802 221792 276830 229183
rect 277558 228427 277610 228433
rect 277558 228369 277610 228375
rect 276802 221764 276878 221792
rect 276850 221482 276878 221764
rect 277570 221482 277598 228369
rect 277954 224807 277982 239686
rect 278434 236795 278462 239686
rect 278784 239672 279038 239700
rect 279168 239672 279326 239700
rect 279552 239672 279806 239700
rect 278422 236789 278474 236795
rect 278422 236731 278474 236737
rect 278230 234569 278282 234575
rect 278230 234511 278282 234517
rect 278038 234199 278090 234205
rect 278038 234141 278090 234147
rect 278050 227619 278078 234141
rect 278038 227613 278090 227619
rect 278038 227555 278090 227561
rect 278242 225695 278270 234511
rect 278710 233903 278762 233909
rect 278710 233845 278762 233851
rect 278326 231979 278378 231985
rect 278326 231921 278378 231927
rect 278230 225689 278282 225695
rect 278230 225631 278282 225637
rect 277942 224801 277994 224807
rect 277942 224743 277994 224749
rect 278338 221482 278366 231921
rect 278422 225837 278474 225843
rect 278614 225837 278666 225843
rect 278474 225797 278614 225825
rect 278422 225779 278474 225785
rect 278614 225779 278666 225785
rect 278722 225251 278750 233845
rect 279010 231985 279038 239672
rect 279298 235907 279326 239672
rect 279286 235901 279338 235907
rect 279286 235843 279338 235849
rect 278998 231979 279050 231985
rect 278998 231921 279050 231927
rect 279778 226805 279806 239672
rect 279874 236869 279902 239686
rect 279862 236863 279914 236869
rect 279862 236805 279914 236811
rect 280258 231911 280286 239686
rect 280642 235981 280670 239686
rect 280992 239672 281246 239700
rect 281376 239672 281630 239700
rect 281760 239672 282014 239700
rect 280630 235975 280682 235981
rect 280630 235917 280682 235923
rect 280246 231905 280298 231911
rect 280246 231847 280298 231853
rect 281218 231467 281246 239672
rect 281494 233977 281546 233983
rect 281494 233919 281546 233925
rect 281302 231831 281354 231837
rect 281302 231773 281354 231779
rect 281206 231461 281258 231467
rect 281206 231403 281258 231409
rect 279862 229019 279914 229025
rect 279862 228961 279914 228967
rect 279766 226799 279818 226805
rect 279766 226741 279818 226747
rect 279094 226059 279146 226065
rect 279094 226001 279146 226007
rect 278710 225245 278762 225251
rect 278710 225187 278762 225193
rect 279106 221792 279134 226001
rect 279106 221764 279182 221792
rect 279154 221482 279182 221764
rect 279874 221482 279902 228961
rect 280630 228057 280682 228063
rect 280630 227999 280682 228005
rect 280642 221482 280670 227999
rect 281314 221792 281342 231773
rect 281506 227693 281534 233919
rect 281494 227687 281546 227693
rect 281494 227629 281546 227635
rect 281602 222513 281630 239672
rect 281986 231837 282014 239672
rect 281974 231831 282026 231837
rect 281974 231773 282026 231779
rect 282178 229247 282206 239686
rect 282562 230875 282590 239686
rect 282960 239672 283166 239700
rect 283296 239672 283550 239700
rect 283680 239672 283934 239700
rect 282934 235605 282986 235611
rect 282934 235547 282986 235553
rect 282550 230869 282602 230875
rect 282550 230811 282602 230817
rect 282166 229241 282218 229247
rect 282166 229183 282218 229189
rect 282550 226429 282602 226435
rect 282550 226371 282602 226377
rect 282562 226065 282590 226371
rect 282550 226059 282602 226065
rect 282550 226001 282602 226007
rect 282070 224727 282122 224733
rect 282070 224669 282122 224675
rect 281590 222507 281642 222513
rect 281590 222449 281642 222455
rect 281314 221764 281390 221792
rect 281362 221482 281390 221764
rect 282082 221482 282110 224669
rect 282946 221482 282974 235547
rect 283138 222439 283166 239672
rect 283522 229321 283550 239672
rect 283906 234575 283934 239672
rect 283894 234569 283946 234575
rect 283894 234511 283946 234517
rect 284002 234205 284030 239686
rect 284400 239672 284702 239700
rect 283990 234199 284042 234205
rect 283990 234141 284042 234147
rect 284374 232719 284426 232725
rect 284374 232661 284426 232667
rect 283510 229315 283562 229321
rect 283510 229257 283562 229263
rect 283606 229093 283658 229099
rect 283606 229035 283658 229041
rect 283126 222433 283178 222439
rect 283126 222375 283178 222381
rect 283618 221792 283646 229035
rect 283618 221764 283694 221792
rect 283666 221482 283694 221764
rect 284386 221482 284414 232661
rect 284674 226731 284702 239672
rect 284770 229099 284798 239686
rect 285046 234643 285098 234649
rect 285046 234585 285098 234591
rect 284758 229093 284810 229099
rect 284758 229035 284810 229041
rect 284662 226725 284714 226731
rect 284662 226667 284714 226673
rect 285058 225769 285086 234585
rect 285154 233761 285182 239686
rect 285504 239672 285758 239700
rect 285984 239672 286238 239700
rect 285142 233755 285194 233761
rect 285142 233697 285194 233703
rect 285730 226657 285758 239672
rect 285910 235531 285962 235537
rect 285910 235473 285962 235479
rect 285718 226651 285770 226657
rect 285718 226593 285770 226599
rect 285142 226355 285194 226361
rect 285142 226297 285194 226303
rect 285046 225763 285098 225769
rect 285046 225705 285098 225711
rect 285154 221482 285182 226297
rect 285922 221792 285950 235473
rect 286210 222735 286238 239672
rect 286306 229025 286334 239686
rect 286690 234649 286718 239686
rect 287074 235611 287102 239686
rect 287350 235679 287402 235685
rect 287350 235621 287402 235627
rect 287062 235605 287114 235611
rect 287062 235547 287114 235553
rect 286678 234643 286730 234649
rect 286678 234585 286730 234591
rect 286294 229019 286346 229025
rect 286294 228961 286346 228967
rect 286678 228501 286730 228507
rect 286678 228443 286730 228449
rect 286198 222729 286250 222735
rect 286198 222671 286250 222677
rect 285922 221764 285998 221792
rect 285970 221482 285998 221764
rect 286690 221482 286718 228443
rect 287362 228304 287390 235621
rect 287458 233465 287486 239686
rect 287808 239672 287966 239700
rect 288192 239672 288446 239700
rect 287446 233459 287498 233465
rect 287446 233401 287498 233407
rect 287938 229173 287966 239672
rect 288022 234273 288074 234279
rect 288022 234215 288074 234221
rect 287926 229167 287978 229173
rect 287926 229109 287978 229115
rect 288034 228433 288062 234215
rect 288418 233391 288446 239672
rect 288406 233385 288458 233391
rect 288406 233327 288458 233333
rect 288022 228427 288074 228433
rect 288022 228369 288074 228375
rect 287362 228276 287486 228304
rect 287458 221482 287486 228276
rect 288118 227169 288170 227175
rect 288118 227111 288170 227117
rect 288130 221792 288158 227111
rect 288514 226509 288542 239686
rect 288898 235315 288926 239686
rect 288886 235309 288938 235315
rect 288886 235251 288938 235257
rect 288886 228797 288938 228803
rect 288886 228739 288938 228745
rect 288502 226503 288554 226509
rect 288502 226445 288554 226451
rect 288130 221764 288206 221792
rect 288178 221482 288206 221764
rect 288898 221482 288926 228739
rect 289378 228507 289406 239686
rect 289728 239672 289982 239700
rect 290112 239672 290366 239700
rect 290496 239672 290654 239700
rect 289954 232947 289982 239672
rect 290338 235833 290366 239672
rect 290326 235827 290378 235833
rect 290326 235769 290378 235775
rect 290422 233533 290474 233539
rect 290422 233475 290474 233481
rect 289942 232941 289994 232947
rect 289942 232883 289994 232889
rect 289654 231461 289706 231467
rect 289654 231403 289706 231409
rect 289366 228501 289418 228507
rect 289366 228443 289418 228449
rect 289666 227175 289694 231403
rect 289750 228871 289802 228877
rect 289750 228813 289802 228819
rect 289654 227169 289706 227175
rect 289654 227111 289706 227117
rect 289762 221482 289790 228813
rect 290434 221792 290462 233475
rect 290626 231023 290654 239672
rect 290818 231467 290846 239686
rect 291216 239672 291518 239700
rect 290902 234421 290954 234427
rect 290902 234363 290954 234369
rect 290806 231461 290858 231467
rect 290806 231403 290858 231409
rect 290614 231017 290666 231023
rect 290614 230959 290666 230965
rect 290914 229987 290942 234363
rect 290998 234051 291050 234057
rect 290998 233993 291050 233999
rect 290902 229981 290954 229987
rect 290902 229923 290954 229929
rect 291010 228063 291038 233993
rect 291490 228655 291518 239672
rect 291478 228649 291530 228655
rect 291478 228591 291530 228597
rect 290998 228057 291050 228063
rect 290998 227999 291050 228005
rect 291586 226361 291614 239686
rect 291936 239672 292190 239700
rect 292320 239672 292574 239700
rect 292704 239672 292958 239700
rect 291958 230351 292010 230357
rect 291958 230293 292010 230299
rect 291574 226355 291626 226361
rect 291574 226297 291626 226303
rect 291190 226207 291242 226213
rect 291190 226149 291242 226155
rect 290434 221764 290510 221792
rect 290482 221482 290510 221764
rect 291202 221482 291230 226149
rect 291970 221482 291998 230293
rect 292162 229067 292190 239672
rect 292546 231393 292574 239672
rect 292930 234427 292958 239672
rect 292918 234421 292970 234427
rect 292918 234363 292970 234369
rect 292534 231387 292586 231393
rect 292534 231329 292586 231335
rect 292148 229058 292204 229067
rect 292148 228993 292204 229002
rect 293122 228919 293150 239686
rect 293398 235457 293450 235463
rect 293398 235399 293450 235405
rect 293108 228910 293164 228919
rect 293108 228845 293164 228854
rect 292630 228353 292682 228359
rect 292630 228295 292682 228301
rect 292642 221792 292670 228295
rect 293410 228156 293438 235399
rect 293506 231245 293534 239686
rect 293782 234125 293834 234131
rect 293782 234067 293834 234073
rect 293494 231239 293546 231245
rect 293494 231181 293546 231187
rect 293410 228128 293534 228156
rect 292642 221764 292718 221792
rect 292690 221482 292718 221764
rect 293506 221482 293534 228128
rect 293794 227915 293822 234067
rect 293890 228359 293918 239686
rect 294240 239672 294494 239700
rect 294624 239672 294878 239700
rect 295008 239672 295262 239700
rect 294466 233835 294494 239672
rect 294850 235463 294878 239672
rect 294838 235457 294890 235463
rect 294838 235399 294890 235405
rect 295234 234279 295262 239672
rect 295222 234273 295274 234279
rect 295222 234215 295274 234221
rect 294454 233829 294506 233835
rect 294454 233771 294506 233777
rect 295330 232725 295358 239686
rect 295714 234131 295742 239686
rect 295702 234125 295754 234131
rect 295702 234067 295754 234073
rect 296098 233909 296126 239686
rect 296448 239672 296606 239700
rect 296928 239672 297182 239700
rect 296470 235013 296522 235019
rect 296470 234955 296522 234961
rect 296086 233903 296138 233909
rect 296086 233845 296138 233851
rect 295318 232719 295370 232725
rect 295318 232661 295370 232667
rect 294934 228945 294986 228951
rect 294934 228887 294986 228893
rect 293878 228353 293930 228359
rect 293878 228295 293930 228301
rect 293782 227909 293834 227915
rect 293782 227851 293834 227857
rect 294262 226577 294314 226583
rect 294262 226519 294314 226525
rect 294274 221496 294302 226519
rect 294240 221468 294302 221496
rect 294946 221496 294974 228887
rect 295702 227983 295754 227989
rect 295702 227925 295754 227931
rect 294946 221468 295008 221496
rect 295714 221482 295742 227925
rect 296482 221496 296510 234955
rect 296578 229215 296606 239672
rect 297154 233317 297182 239672
rect 297250 233539 297278 239686
rect 297238 233533 297290 233539
rect 297238 233475 297290 233481
rect 297142 233311 297194 233317
rect 297142 233253 297194 233259
rect 297430 231017 297482 231023
rect 297430 230959 297482 230965
rect 296564 229206 296620 229215
rect 296564 229141 296620 229150
rect 297442 226583 297470 230959
rect 297430 226577 297482 226583
rect 297430 226519 297482 226525
rect 297634 226287 297662 239686
rect 298018 235019 298046 239686
rect 298006 235013 298058 235019
rect 298006 234955 298058 234961
rect 298402 229691 298430 239686
rect 298752 239672 299006 239700
rect 299136 239672 299390 239700
rect 298978 236943 299006 239672
rect 298966 236937 299018 236943
rect 298966 236879 299018 236885
rect 299254 235087 299306 235093
rect 299254 235029 299306 235035
rect 299266 230505 299294 235029
rect 299362 234691 299390 239672
rect 299458 234987 299486 239686
rect 299842 235537 299870 239686
rect 299830 235531 299882 235537
rect 299830 235473 299882 235479
rect 299444 234978 299500 234987
rect 299444 234913 299500 234922
rect 299348 234682 299404 234691
rect 299348 234617 299404 234626
rect 300226 231319 300254 239686
rect 299446 231313 299498 231319
rect 299446 231255 299498 231261
rect 300214 231313 300266 231319
rect 300214 231255 300266 231261
rect 299254 230499 299306 230505
rect 299254 230441 299306 230447
rect 298678 230425 298730 230431
rect 298678 230367 298730 230373
rect 298006 229685 298058 229691
rect 298006 229627 298058 229633
rect 298390 229685 298442 229691
rect 298390 229627 298442 229633
rect 297238 226281 297290 226287
rect 297238 226223 297290 226229
rect 297622 226281 297674 226287
rect 297622 226223 297674 226229
rect 296448 221468 296510 221496
rect 297250 221482 297278 226223
rect 298018 221482 298046 229627
rect 298210 226805 298430 226824
rect 298198 226799 298442 226805
rect 298250 226796 298390 226799
rect 298198 226741 298250 226747
rect 298390 226741 298442 226747
rect 298102 226725 298154 226731
rect 298102 226667 298154 226673
rect 298114 226435 298142 226667
rect 298102 226429 298154 226435
rect 298102 226371 298154 226377
rect 298690 221792 298718 230367
rect 298690 221764 298766 221792
rect 298738 221482 298766 221764
rect 299458 221482 299486 231255
rect 300598 230869 300650 230875
rect 300598 230811 300650 230817
rect 300610 226731 300638 230811
rect 300598 226725 300650 226731
rect 300598 226667 300650 226673
rect 300706 226139 300734 239686
rect 301056 239672 301310 239700
rect 301440 239672 301694 239700
rect 301776 239672 302078 239700
rect 300982 230277 301034 230283
rect 300982 230219 301034 230225
rect 300214 226133 300266 226139
rect 300214 226075 300266 226081
rect 300694 226133 300746 226139
rect 300694 226075 300746 226081
rect 300226 221482 300254 226075
rect 300994 221792 301022 230219
rect 301282 226213 301310 239672
rect 301666 234057 301694 239672
rect 302050 236174 302078 239672
rect 301954 236146 302078 236174
rect 301654 234051 301706 234057
rect 301654 233993 301706 233999
rect 301750 228575 301802 228581
rect 301750 228517 301802 228523
rect 301270 226207 301322 226213
rect 301270 226149 301322 226155
rect 300994 221764 301070 221792
rect 301042 221482 301070 221764
rect 301762 221482 301790 228517
rect 301954 222587 301982 236146
rect 302146 225325 302174 239686
rect 302544 239672 302846 239700
rect 302326 235383 302378 235389
rect 302326 235325 302378 235331
rect 302230 234347 302282 234353
rect 302230 234289 302282 234295
rect 302242 227841 302270 234289
rect 302338 230653 302366 235325
rect 302326 230647 302378 230653
rect 302326 230589 302378 230595
rect 302518 230499 302570 230505
rect 302518 230441 302570 230447
rect 302230 227835 302282 227841
rect 302230 227777 302282 227783
rect 302134 225319 302186 225325
rect 302134 225261 302186 225267
rect 301942 222581 301994 222587
rect 301942 222523 301994 222529
rect 302530 221482 302558 230441
rect 302818 222661 302846 239672
rect 302914 233613 302942 239686
rect 303264 239672 303518 239700
rect 303648 239672 303902 239700
rect 303984 239672 304286 239700
rect 302902 233607 302954 233613
rect 302902 233549 302954 233555
rect 303490 228581 303518 239672
rect 303478 228575 303530 228581
rect 303478 228517 303530 228523
rect 303190 225541 303242 225547
rect 303190 225483 303242 225489
rect 302806 222655 302858 222661
rect 302806 222597 302858 222603
rect 303202 221792 303230 225483
rect 303874 225399 303902 239672
rect 304150 234717 304202 234723
rect 304150 234659 304202 234665
rect 304162 230505 304190 234659
rect 304150 230499 304202 230505
rect 304150 230441 304202 230447
rect 303958 227761 304010 227767
rect 303958 227703 304010 227709
rect 303862 225393 303914 225399
rect 303862 225335 303914 225341
rect 303202 221764 303278 221792
rect 303250 221482 303278 221764
rect 303970 221482 303998 227703
rect 304258 222809 304286 239672
rect 304450 228729 304478 239686
rect 304834 235389 304862 239686
rect 305184 239672 305246 239700
rect 305568 239672 305822 239700
rect 305952 239672 306206 239700
rect 305110 235753 305162 235759
rect 305110 235695 305162 235701
rect 304822 235383 304874 235389
rect 304822 235325 304874 235331
rect 304726 234495 304778 234501
rect 304726 234437 304778 234443
rect 304438 228723 304490 228729
rect 304438 228665 304490 228671
rect 304738 227767 304766 234437
rect 304822 230203 304874 230209
rect 304822 230145 304874 230151
rect 304726 227761 304778 227767
rect 304726 227703 304778 227709
rect 304246 222803 304298 222809
rect 304246 222745 304298 222751
rect 304834 221482 304862 230145
rect 305122 225177 305150 235695
rect 305218 233983 305246 239672
rect 305794 237017 305822 239672
rect 305782 237011 305834 237017
rect 305782 236953 305834 236959
rect 305206 233977 305258 233983
rect 305206 233919 305258 233925
rect 305494 231535 305546 231541
rect 305494 231477 305546 231483
rect 305110 225171 305162 225177
rect 305110 225113 305162 225119
rect 305506 221792 305534 231477
rect 306178 228803 306206 239672
rect 306274 233687 306302 239686
rect 306658 236174 306686 239686
rect 307056 239672 307262 239700
rect 307392 239672 307646 239700
rect 307776 239672 308030 239700
rect 308256 239672 308510 239700
rect 306658 236146 306782 236174
rect 306646 234791 306698 234797
rect 306646 234733 306698 234739
rect 306262 233681 306314 233687
rect 306262 233623 306314 233629
rect 306658 230579 306686 234733
rect 306646 230573 306698 230579
rect 306646 230515 306698 230521
rect 306166 228797 306218 228803
rect 306166 228739 306218 228745
rect 306262 227539 306314 227545
rect 306262 227481 306314 227487
rect 305506 221764 305582 221792
rect 305554 221482 305582 221764
rect 306274 221482 306302 227481
rect 306754 225473 306782 236146
rect 307030 230055 307082 230061
rect 307030 229997 307082 230003
rect 306742 225467 306794 225473
rect 306742 225409 306794 225415
rect 307042 221482 307070 229997
rect 307234 223031 307262 239672
rect 307618 231139 307646 239672
rect 307604 231130 307660 231139
rect 307604 231065 307660 231074
rect 307702 228205 307754 228211
rect 307702 228147 307754 228153
rect 307222 223025 307274 223031
rect 307222 222967 307274 222973
rect 307714 221792 307742 228147
rect 308002 222883 308030 239672
rect 308278 236049 308330 236055
rect 308278 235991 308330 235997
rect 308182 235235 308234 235241
rect 308182 235177 308234 235183
rect 308194 231023 308222 235177
rect 308182 231017 308234 231023
rect 308182 230959 308234 230965
rect 308290 227989 308318 235991
rect 308482 234353 308510 239672
rect 308578 237165 308606 239686
rect 308566 237159 308618 237165
rect 308566 237101 308618 237107
rect 308470 234347 308522 234353
rect 308470 234289 308522 234295
rect 308566 230647 308618 230653
rect 308566 230589 308618 230595
rect 308278 227983 308330 227989
rect 308278 227925 308330 227931
rect 307990 222877 308042 222883
rect 307990 222819 308042 222825
rect 307714 221764 307790 221792
rect 307762 221482 307790 221764
rect 308578 221482 308606 230589
rect 308962 228951 308990 239686
rect 309346 235093 309374 239686
rect 309696 239672 309950 239700
rect 310080 239672 310334 239700
rect 310464 239672 310718 239700
rect 309334 235087 309386 235093
rect 309334 235029 309386 235035
rect 308950 228945 309002 228951
rect 308950 228887 309002 228893
rect 309334 225615 309386 225621
rect 309334 225557 309386 225563
rect 309346 221482 309374 225557
rect 309922 225547 309950 239672
rect 310006 229907 310058 229913
rect 310006 229849 310058 229855
rect 309910 225541 309962 225547
rect 309910 225483 309962 225489
rect 310018 221792 310046 229849
rect 310306 223105 310334 239672
rect 310690 228877 310718 239672
rect 310786 237091 310814 239686
rect 310774 237085 310826 237091
rect 310774 237027 310826 237033
rect 311170 235685 311198 239686
rect 311554 237239 311582 239686
rect 312000 239672 312254 239700
rect 312384 239672 312638 239700
rect 311542 237233 311594 237239
rect 311542 237175 311594 237181
rect 311158 235679 311210 235685
rect 311158 235621 311210 235627
rect 311254 234199 311306 234205
rect 311254 234141 311306 234147
rect 311158 233459 311210 233465
rect 311158 233401 311210 233407
rect 311062 233385 311114 233391
rect 311062 233327 311114 233333
rect 310774 230129 310826 230135
rect 310774 230071 310826 230077
rect 310678 228871 310730 228877
rect 310678 228813 310730 228819
rect 310294 223099 310346 223105
rect 310294 223041 310346 223047
rect 310018 221764 310094 221792
rect 310066 221482 310094 221764
rect 310786 221482 310814 230071
rect 311074 228211 311102 233327
rect 311062 228205 311114 228211
rect 311062 228147 311114 228153
rect 311170 227397 311198 233401
rect 311266 227545 311294 234141
rect 312226 231541 312254 239672
rect 312214 231535 312266 231541
rect 312214 231477 312266 231483
rect 311638 230499 311690 230505
rect 311638 230441 311690 230447
rect 311254 227539 311306 227545
rect 311254 227481 311306 227487
rect 311158 227391 311210 227397
rect 311158 227333 311210 227339
rect 311650 221482 311678 230441
rect 312310 225097 312362 225103
rect 312310 225039 312362 225045
rect 312322 221792 312350 225039
rect 312610 222957 312638 239672
rect 312706 234427 312734 239686
rect 313104 239672 313406 239700
rect 312694 234421 312746 234427
rect 312694 234363 312746 234369
rect 313078 229833 313130 229839
rect 313078 229775 313130 229781
rect 312598 222951 312650 222957
rect 312598 222893 312650 222899
rect 312322 221764 312398 221792
rect 312370 221482 312398 221764
rect 313090 221482 313118 229775
rect 313378 223179 313406 239672
rect 313474 230431 313502 239686
rect 313858 236055 313886 239686
rect 314208 239672 314462 239700
rect 314592 239672 314846 239700
rect 313942 236123 313994 236129
rect 313942 236065 313994 236071
rect 313846 236049 313898 236055
rect 313846 235991 313898 235997
rect 313846 234495 313898 234501
rect 313846 234437 313898 234443
rect 313462 230425 313514 230431
rect 313462 230367 313514 230373
rect 313858 228452 313886 234437
rect 313954 230727 313982 236065
rect 314434 234501 314462 239672
rect 314818 237313 314846 239672
rect 314806 237307 314858 237313
rect 314806 237249 314858 237255
rect 314422 234495 314474 234501
rect 314422 234437 314474 234443
rect 314518 231091 314570 231097
rect 314518 231033 314570 231039
rect 313942 230721 313994 230727
rect 313942 230663 313994 230669
rect 313858 228424 313982 228452
rect 313954 228285 313982 228424
rect 313846 228279 313898 228285
rect 313846 228221 313898 228227
rect 313942 228279 313994 228285
rect 313942 228221 313994 228227
rect 313366 223173 313418 223179
rect 313366 223115 313418 223121
rect 313858 221482 313886 228221
rect 314530 221792 314558 231033
rect 314914 230357 314942 239686
rect 315298 234723 315326 239686
rect 315286 234717 315338 234723
rect 315286 234659 315338 234665
rect 314902 230351 314954 230357
rect 314902 230293 314954 230299
rect 315382 227465 315434 227471
rect 315382 227407 315434 227413
rect 314530 221764 314606 221792
rect 314578 221482 314606 221764
rect 315394 221482 315422 227407
rect 315778 225621 315806 239686
rect 316176 239672 316382 239700
rect 316512 239672 316766 239700
rect 316896 239672 317150 239700
rect 316150 229611 316202 229617
rect 316150 229553 316202 229559
rect 315766 225615 315818 225621
rect 315766 225557 315818 225563
rect 316162 221482 316190 229553
rect 316354 224659 316382 239672
rect 316738 231287 316766 239672
rect 317122 237387 317150 239672
rect 317110 237381 317162 237387
rect 317110 237323 317162 237329
rect 317218 235759 317246 239686
rect 317602 237461 317630 239686
rect 317590 237455 317642 237461
rect 317590 237397 317642 237403
rect 317206 235753 317258 235759
rect 317206 235695 317258 235701
rect 316724 231278 316780 231287
rect 316724 231213 316780 231222
rect 317590 230573 317642 230579
rect 317590 230515 317642 230521
rect 316822 229537 316874 229543
rect 316822 229479 316874 229485
rect 316342 224653 316394 224659
rect 316342 224595 316394 224601
rect 316834 221792 316862 229479
rect 316834 221764 316910 221792
rect 316882 221482 316910 221764
rect 317602 221482 317630 230515
rect 317986 230283 318014 239686
rect 318166 235605 318218 235611
rect 318166 235547 318218 235553
rect 317974 230277 318026 230283
rect 317974 230219 318026 230225
rect 318178 227471 318206 235547
rect 318370 234205 318398 239686
rect 318720 239672 318974 239700
rect 319200 239672 319454 239700
rect 318358 234199 318410 234205
rect 318358 234141 318410 234147
rect 318166 227465 318218 227471
rect 318166 227407 318218 227413
rect 318358 225689 318410 225695
rect 318358 225631 318410 225637
rect 318370 221482 318398 225631
rect 318946 225367 318974 239672
rect 319426 236174 319454 239672
rect 319330 236146 319454 236174
rect 319126 229759 319178 229765
rect 319126 229701 319178 229707
rect 318932 225358 318988 225367
rect 318932 225293 318988 225302
rect 319138 221792 319166 229701
rect 319330 224585 319358 236146
rect 319414 233311 319466 233317
rect 319414 233253 319466 233259
rect 319426 227712 319454 233253
rect 319522 231435 319550 239686
rect 319606 235901 319658 235907
rect 319606 235843 319658 235849
rect 319508 231426 319564 231435
rect 319508 231361 319564 231370
rect 319618 230801 319646 235843
rect 319906 233317 319934 239686
rect 320290 233465 320318 239686
rect 320640 239672 320894 239700
rect 321024 239672 321278 239700
rect 321408 239672 321662 239700
rect 320866 237535 320894 239672
rect 320854 237529 320906 237535
rect 320854 237471 320906 237477
rect 320854 235975 320906 235981
rect 320854 235917 320906 235923
rect 320662 234569 320714 234575
rect 320662 234511 320714 234517
rect 320278 233459 320330 233465
rect 320278 233401 320330 233407
rect 319894 233311 319946 233317
rect 319894 233253 319946 233259
rect 320566 231683 320618 231689
rect 320566 231625 320618 231631
rect 319606 230795 319658 230801
rect 319606 230737 319658 230743
rect 319426 227684 320030 227712
rect 320002 227619 320030 227684
rect 319894 227613 319946 227619
rect 319894 227555 319946 227561
rect 319990 227613 320042 227619
rect 319990 227555 320042 227561
rect 319318 224579 319370 224585
rect 319318 224521 319370 224527
rect 319138 221764 319214 221792
rect 319186 221482 319214 221764
rect 319906 221482 319934 227555
rect 320578 226232 320606 231625
rect 320674 230653 320702 234511
rect 320662 230647 320714 230653
rect 320662 230589 320714 230595
rect 320866 230505 320894 235917
rect 320854 230499 320906 230505
rect 320854 230441 320906 230447
rect 321250 230209 321278 239672
rect 321634 234797 321662 239672
rect 321622 234791 321674 234797
rect 321622 234733 321674 234739
rect 321238 230203 321290 230209
rect 321238 230145 321290 230151
rect 320578 226204 320702 226232
rect 320674 221482 320702 226204
rect 321334 225985 321386 225991
rect 321334 225927 321386 225933
rect 321346 221792 321374 225927
rect 321730 225695 321758 239686
rect 322128 239672 322334 239700
rect 322102 231165 322154 231171
rect 322102 231107 322154 231113
rect 321718 225689 321770 225695
rect 321718 225631 321770 225637
rect 321346 221764 321422 221792
rect 321394 221482 321422 221764
rect 322114 221482 322142 231107
rect 322306 224437 322334 239672
rect 322498 231583 322526 239686
rect 322944 239672 323198 239700
rect 323328 239672 323582 239700
rect 323712 239672 323966 239700
rect 323170 236174 323198 239672
rect 323170 236146 323294 236174
rect 323062 234865 323114 234871
rect 323062 234807 323114 234813
rect 322484 231574 322540 231583
rect 322484 231509 322540 231518
rect 323074 230949 323102 234807
rect 323158 233755 323210 233761
rect 323158 233697 323210 233703
rect 323062 230943 323114 230949
rect 323062 230885 323114 230891
rect 323170 230579 323198 233697
rect 323158 230573 323210 230579
rect 323158 230515 323210 230521
rect 322966 228131 323018 228137
rect 322966 228073 323018 228079
rect 322294 224431 322346 224437
rect 322294 224373 322346 224379
rect 322978 221496 323006 228073
rect 323266 224511 323294 236146
rect 323554 234575 323582 239672
rect 323938 238941 323966 239672
rect 323926 238935 323978 238941
rect 323926 238877 323978 238883
rect 323542 234569 323594 234575
rect 323542 234511 323594 234517
rect 323638 231017 323690 231023
rect 323638 230959 323690 230965
rect 323254 224505 323306 224511
rect 323254 224447 323306 224453
rect 322944 221468 323006 221496
rect 323650 221496 323678 230959
rect 324034 230061 324062 239686
rect 324418 239015 324446 239686
rect 324406 239009 324458 239015
rect 324406 238951 324458 238957
rect 324214 235161 324266 235167
rect 324214 235103 324266 235109
rect 324022 230055 324074 230061
rect 324022 229997 324074 230003
rect 324226 226879 324254 235103
rect 324802 233391 324830 239686
rect 325152 239672 325214 239700
rect 325536 239672 325790 239700
rect 325920 239672 326174 239700
rect 325186 236174 325214 239672
rect 325186 236146 325310 236174
rect 324790 233385 324842 233391
rect 324790 233327 324842 233333
rect 325174 231609 325226 231615
rect 325174 231551 325226 231557
rect 324214 226873 324266 226879
rect 324214 226815 324266 226821
rect 324406 225245 324458 225251
rect 324406 225187 324458 225193
rect 323650 221468 323712 221496
rect 324418 221482 324446 225187
rect 325186 221496 325214 231551
rect 325282 224363 325310 236146
rect 325762 230135 325790 239672
rect 326146 236129 326174 239672
rect 326134 236123 326186 236129
rect 326134 236065 326186 236071
rect 326242 235907 326270 239686
rect 326722 238867 326750 239686
rect 326710 238861 326762 238867
rect 326710 238803 326762 238809
rect 326230 235901 326282 235907
rect 326230 235843 326282 235849
rect 326806 234643 326858 234649
rect 326806 234585 326858 234591
rect 326710 231757 326762 231763
rect 326710 231699 326762 231705
rect 325750 230129 325802 230135
rect 325750 230071 325802 230077
rect 325846 227687 325898 227693
rect 325846 227629 325898 227635
rect 325270 224357 325322 224363
rect 325270 224299 325322 224305
rect 325152 221468 325214 221496
rect 325858 221496 325886 227629
rect 325858 221468 325920 221496
rect 326722 221482 326750 231699
rect 326818 230875 326846 234585
rect 327106 231615 327134 239686
rect 327456 239672 327710 239700
rect 327840 239672 328094 239700
rect 327682 234871 327710 239672
rect 327670 234865 327722 234871
rect 327670 234807 327722 234813
rect 327766 233385 327818 233391
rect 327766 233327 327818 233333
rect 327094 231609 327146 231615
rect 327094 231551 327146 231557
rect 326806 230869 326858 230875
rect 326806 230811 326858 230817
rect 327382 225837 327434 225843
rect 327382 225779 327434 225785
rect 327394 221792 327422 225779
rect 327778 225515 327806 233327
rect 328066 225663 328094 239672
rect 328162 236174 328190 239686
rect 328162 236146 328286 236174
rect 328150 233237 328202 233243
rect 328150 233179 328202 233185
rect 328052 225654 328108 225663
rect 328052 225589 328108 225598
rect 327764 225506 327820 225515
rect 327764 225441 327820 225450
rect 327394 221764 327470 221792
rect 327442 221482 327470 221764
rect 328162 221482 328190 233179
rect 328258 224289 328286 236146
rect 328342 233533 328394 233539
rect 328342 233475 328394 233481
rect 328354 231023 328382 233475
rect 328546 233391 328574 239686
rect 328930 238793 328958 239686
rect 328918 238787 328970 238793
rect 328918 238729 328970 238735
rect 329314 234649 329342 239686
rect 329664 239672 329918 239700
rect 330048 239672 330302 239700
rect 330480 239672 330782 239700
rect 329890 238719 329918 239672
rect 329878 238713 329930 238719
rect 329878 238655 329930 238661
rect 329302 234643 329354 234649
rect 329302 234585 329354 234591
rect 328534 233385 328586 233391
rect 328534 233327 328586 233333
rect 330274 231731 330302 239672
rect 330260 231722 330316 231731
rect 330260 231657 330316 231666
rect 328342 231017 328394 231023
rect 328342 230959 328394 230965
rect 329590 230943 329642 230949
rect 329590 230885 329642 230891
rect 328918 228427 328970 228433
rect 328918 228369 328970 228375
rect 328246 224283 328298 224289
rect 328246 224225 328298 224231
rect 328930 221482 328958 228369
rect 329602 221792 329630 230885
rect 330454 225911 330506 225917
rect 330454 225853 330506 225859
rect 329602 221764 329678 221792
rect 329650 221482 329678 221764
rect 330466 221482 330494 225853
rect 330754 224141 330782 239672
rect 330850 225811 330878 239686
rect 331248 239672 331550 239700
rect 331414 234939 331466 234945
rect 331414 234881 331466 234887
rect 331222 233829 331274 233835
rect 331222 233771 331274 233777
rect 331126 233385 331178 233391
rect 331126 233327 331178 233333
rect 331138 228433 331166 233327
rect 331234 230949 331262 233771
rect 331318 233015 331370 233021
rect 331318 232957 331370 232963
rect 331222 230943 331274 230949
rect 331222 230885 331274 230891
rect 331126 228427 331178 228433
rect 331126 228369 331178 228375
rect 331330 226972 331358 232957
rect 331234 226944 331358 226972
rect 330836 225802 330892 225811
rect 330836 225737 330892 225746
rect 330742 224135 330794 224141
rect 330742 224077 330794 224083
rect 331234 221482 331262 226944
rect 331426 225917 331454 234881
rect 331414 225911 331466 225917
rect 331414 225853 331466 225859
rect 331522 224215 331550 239672
rect 331618 229913 331646 239686
rect 331968 239672 332222 239700
rect 332352 239672 332606 239700
rect 332194 235167 332222 239672
rect 332182 235161 332234 235167
rect 332182 235103 332234 235109
rect 332578 234099 332606 239672
rect 332674 238645 332702 239686
rect 332662 238639 332714 238645
rect 332662 238581 332714 238587
rect 332564 234090 332620 234099
rect 332564 234025 332620 234034
rect 331894 229981 331946 229987
rect 331894 229923 331946 229929
rect 331606 229907 331658 229913
rect 331606 229849 331658 229855
rect 331510 224209 331562 224215
rect 331510 224151 331562 224157
rect 331906 221792 331934 229923
rect 333058 228179 333086 239686
rect 333442 234945 333470 239686
rect 333430 234939 333482 234945
rect 333430 234881 333482 234887
rect 333826 231879 333854 239686
rect 334272 239672 334526 239700
rect 334656 239672 334910 239700
rect 334294 239527 334346 239533
rect 334294 239469 334346 239475
rect 334306 236129 334334 239469
rect 334294 236123 334346 236129
rect 334294 236065 334346 236071
rect 334102 235827 334154 235833
rect 334102 235769 334154 235775
rect 333812 231870 333868 231879
rect 333812 231805 333868 231814
rect 333044 228170 333100 228179
rect 333044 228105 333100 228114
rect 334114 225991 334142 235769
rect 334198 233163 334250 233169
rect 334198 233105 334250 233111
rect 334102 225985 334154 225991
rect 334102 225927 334154 225933
rect 333526 225171 333578 225177
rect 333526 225113 333578 225119
rect 332662 223765 332714 223771
rect 332662 223707 332714 223713
rect 331906 221764 331982 221792
rect 331954 221482 331982 221764
rect 332674 221482 332702 223707
rect 333538 221482 333566 225113
rect 334210 221792 334238 233105
rect 334498 224067 334526 239672
rect 334882 231689 334910 239672
rect 334978 235241 335006 239686
rect 334966 235235 335018 235241
rect 334966 235177 335018 235183
rect 335362 233391 335390 239686
rect 335746 238571 335774 239686
rect 336096 239672 336350 239700
rect 336480 239672 336734 239700
rect 335734 238565 335786 238571
rect 335734 238507 335786 238513
rect 335350 233385 335402 233391
rect 335350 233327 335402 233333
rect 334870 231683 334922 231689
rect 334870 231625 334922 231631
rect 336322 229839 336350 239672
rect 336706 238497 336734 239672
rect 336850 239404 336878 239686
rect 336850 239376 336926 239404
rect 336694 238491 336746 238497
rect 336694 238433 336746 238439
rect 336310 229833 336362 229839
rect 336310 229775 336362 229781
rect 334966 229463 335018 229469
rect 334966 229405 335018 229411
rect 334486 224061 334538 224067
rect 334486 224003 334538 224009
rect 334210 221764 334286 221792
rect 334258 221482 334286 221764
rect 334978 221482 335006 229405
rect 336898 227439 336926 239376
rect 336884 227430 336940 227439
rect 336884 227365 336940 227374
rect 336406 226059 336458 226065
rect 336406 226001 336458 226007
rect 335734 223691 335786 223697
rect 335734 223633 335786 223639
rect 335746 221482 335774 223633
rect 336418 221792 336446 226001
rect 337186 223993 337214 239686
rect 337366 233607 337418 233613
rect 337366 233549 337418 233555
rect 337270 232867 337322 232873
rect 337270 232809 337322 232815
rect 337174 223987 337226 223993
rect 337174 223929 337226 223935
rect 336418 221764 336494 221792
rect 336466 221482 336494 221764
rect 337282 221482 337310 232809
rect 337378 231171 337406 233549
rect 337570 231763 337598 239686
rect 337654 235457 337706 235463
rect 337654 235399 337706 235405
rect 337558 231757 337610 231763
rect 337558 231699 337610 231705
rect 337366 231165 337418 231171
rect 337366 231107 337418 231113
rect 337666 225103 337694 235399
rect 338050 233761 338078 239686
rect 338400 239672 338654 239700
rect 338784 239672 339038 239700
rect 339168 239672 339422 239700
rect 338038 233755 338090 233761
rect 338038 233697 338090 233703
rect 338626 233539 338654 239672
rect 339010 238423 339038 239672
rect 338998 238417 339050 238423
rect 338998 238359 339050 238365
rect 338614 233533 338666 233539
rect 338614 233475 338666 233481
rect 338038 233089 338090 233095
rect 338038 233031 338090 233037
rect 337654 225097 337706 225103
rect 337654 225039 337706 225045
rect 338050 221482 338078 233031
rect 339394 228327 339422 239672
rect 339490 235463 339518 239686
rect 339888 239672 340190 239700
rect 340272 239672 340478 239700
rect 340608 239672 340862 239700
rect 340992 239672 341246 239700
rect 341376 239672 341630 239700
rect 339478 235457 339530 235463
rect 339478 235399 339530 235405
rect 339766 233903 339818 233909
rect 339766 233845 339818 233851
rect 339380 228318 339436 228327
rect 339380 228253 339436 228262
rect 339478 226873 339530 226879
rect 339478 226815 339530 226821
rect 338710 223469 338762 223475
rect 338710 223411 338762 223417
rect 338722 221792 338750 223411
rect 338722 221764 338798 221792
rect 338770 221482 338798 221764
rect 339490 221482 339518 226815
rect 339778 225177 339806 233845
rect 340162 225959 340190 239672
rect 340246 232793 340298 232799
rect 340246 232735 340298 232741
rect 340148 225950 340204 225959
rect 340148 225885 340204 225894
rect 339766 225171 339818 225177
rect 339766 225113 339818 225119
rect 340258 221482 340286 232735
rect 340450 223919 340478 239672
rect 340834 233243 340862 239672
rect 341218 236129 341246 239672
rect 341206 236123 341258 236129
rect 341206 236065 341258 236071
rect 341602 234247 341630 239672
rect 341794 238349 341822 239686
rect 341782 238343 341834 238349
rect 341782 238285 341834 238291
rect 341588 234238 341644 234247
rect 341588 234173 341644 234182
rect 341206 234125 341258 234131
rect 341206 234067 341258 234073
rect 340822 233237 340874 233243
rect 340822 233179 340874 233185
rect 341218 228063 341246 234067
rect 342178 228623 342206 239686
rect 342562 235727 342590 239686
rect 342912 239672 343166 239700
rect 343296 239672 343550 239700
rect 342548 235718 342604 235727
rect 342548 235653 342604 235662
rect 342164 228614 342220 228623
rect 342164 228549 342220 228558
rect 341014 228057 341066 228063
rect 341014 227999 341066 228005
rect 341206 228057 341258 228063
rect 341206 227999 341258 228005
rect 340438 223913 340490 223919
rect 340438 223855 340490 223861
rect 341026 221792 341054 227999
rect 343138 227291 343166 239672
rect 343522 235833 343550 239672
rect 343510 235827 343562 235833
rect 343510 235769 343562 235775
rect 343222 232571 343274 232577
rect 343222 232513 343274 232519
rect 343124 227282 343180 227291
rect 343124 227217 343180 227226
rect 342550 225763 342602 225769
rect 342550 225705 342602 225711
rect 341782 223543 341834 223549
rect 341782 223485 341834 223491
rect 341026 221764 341102 221792
rect 341074 221482 341102 221764
rect 341794 221482 341822 223485
rect 342562 221482 342590 225705
rect 343234 221792 343262 232513
rect 343618 223845 343646 239686
rect 344002 233211 344030 239686
rect 344386 234057 344414 239686
rect 344086 234051 344138 234057
rect 344086 233993 344138 233999
rect 344374 234051 344426 234057
rect 344374 233993 344426 233999
rect 343988 233202 344044 233211
rect 343988 233137 344044 233146
rect 344098 228137 344126 233993
rect 344470 233681 344522 233687
rect 344470 233623 344522 233629
rect 344482 231097 344510 233623
rect 344470 231091 344522 231097
rect 344470 231033 344522 231039
rect 344086 228131 344138 228137
rect 344086 228073 344138 228079
rect 343990 227909 344042 227915
rect 343990 227851 344042 227857
rect 343606 223839 343658 223845
rect 343606 223781 343658 223787
rect 343234 221764 343310 221792
rect 343282 221482 343310 221764
rect 344002 221482 344030 227851
rect 344770 227143 344798 239686
rect 345120 239672 345374 239700
rect 345346 238275 345374 239672
rect 345442 239672 345600 239700
rect 345334 238269 345386 238275
rect 345334 238211 345386 238217
rect 345442 228475 345470 239672
rect 345922 234131 345950 239686
rect 346320 239672 346622 239700
rect 345910 234125 345962 234131
rect 345910 234067 345962 234073
rect 346294 232645 346346 232651
rect 346294 232587 346346 232593
rect 345428 228466 345484 228475
rect 345428 228401 345484 228410
rect 344756 227134 344812 227143
rect 344756 227069 344812 227078
rect 345526 225911 345578 225917
rect 345526 225853 345578 225859
rect 344854 223617 344906 223623
rect 344854 223559 344906 223565
rect 344866 221482 344894 223559
rect 345538 221792 345566 225853
rect 345538 221764 345614 221792
rect 345586 221482 345614 221764
rect 346306 221482 346334 232587
rect 346594 223771 346622 239672
rect 346690 238201 346718 239686
rect 346678 238195 346730 238201
rect 346678 238137 346730 238143
rect 346870 235309 346922 235315
rect 346870 235251 346922 235257
rect 346882 225917 346910 235251
rect 347074 233169 347102 239686
rect 347424 239672 347678 239700
rect 347808 239672 348062 239700
rect 347650 234839 347678 239672
rect 347636 234830 347692 234839
rect 347636 234765 347692 234774
rect 347062 233163 347114 233169
rect 347062 233105 347114 233111
rect 346966 232349 347018 232355
rect 346966 232291 347018 232297
rect 346978 232059 347006 232291
rect 346966 232053 347018 232059
rect 346966 231995 347018 232001
rect 347062 229389 347114 229395
rect 347062 229331 347114 229337
rect 346870 225911 346922 225917
rect 346870 225853 346922 225859
rect 346582 223765 346634 223771
rect 346582 223707 346634 223713
rect 347074 221482 347102 229331
rect 348034 223623 348062 239672
rect 348022 223617 348074 223623
rect 348022 223559 348074 223565
rect 348130 223549 348158 239686
rect 348514 229765 348542 239686
rect 348694 234273 348746 234279
rect 348694 234215 348746 234221
rect 348502 229759 348554 229765
rect 348502 229701 348554 229707
rect 348598 227317 348650 227323
rect 348598 227259 348650 227265
rect 348118 223543 348170 223549
rect 348118 223485 348170 223491
rect 347734 223321 347786 223327
rect 347734 223263 347786 223269
rect 347746 221792 347774 223263
rect 347746 221764 347822 221792
rect 347794 221482 347822 221764
rect 348610 221482 348638 227259
rect 348706 225029 348734 234215
rect 348898 233613 348926 239686
rect 349344 239672 349598 239700
rect 349728 239672 349982 239700
rect 350112 239672 350366 239700
rect 348886 233607 348938 233613
rect 348886 233549 348938 233555
rect 349366 232423 349418 232429
rect 349366 232365 349418 232371
rect 348694 225023 348746 225029
rect 348694 224965 348746 224971
rect 349378 221482 349406 232365
rect 349570 223697 349598 239672
rect 349954 238127 349982 239672
rect 349942 238121 349994 238127
rect 349942 238063 349994 238069
rect 350338 233095 350366 239672
rect 350434 239163 350462 239686
rect 350832 239672 351134 239700
rect 350422 239157 350474 239163
rect 350422 239099 350474 239105
rect 350326 233089 350378 233095
rect 350326 233031 350378 233037
rect 350038 227835 350090 227841
rect 350038 227777 350090 227783
rect 349558 223691 349610 223697
rect 349558 223633 349610 223639
rect 350050 221792 350078 227777
rect 351106 223475 351134 239672
rect 351094 223469 351146 223475
rect 351094 223411 351146 223417
rect 350806 223395 350858 223401
rect 350806 223337 350858 223343
rect 350050 221764 350126 221792
rect 350098 221482 350126 221764
rect 350818 221482 350846 223337
rect 351202 223327 351230 239686
rect 351552 239672 351806 239700
rect 351936 239672 352190 239700
rect 352320 239672 352574 239700
rect 351382 233977 351434 233983
rect 351382 233919 351434 233925
rect 351394 225251 351422 233919
rect 351778 229617 351806 239672
rect 352162 234279 352190 239672
rect 352150 234273 352202 234279
rect 352150 234215 352202 234221
rect 352342 232645 352394 232651
rect 352342 232587 352394 232593
rect 351766 229611 351818 229617
rect 351766 229553 351818 229559
rect 351574 227243 351626 227249
rect 351574 227185 351626 227191
rect 351382 225245 351434 225251
rect 351382 225187 351434 225193
rect 351190 223321 351242 223327
rect 351190 223263 351242 223269
rect 351586 221482 351614 227185
rect 352354 221496 352382 232587
rect 352546 223401 352574 239672
rect 352738 237979 352766 239686
rect 352726 237973 352778 237979
rect 352726 237915 352778 237921
rect 353122 233021 353150 239686
rect 353506 238053 353534 239686
rect 353856 239672 354110 239700
rect 353494 238047 353546 238053
rect 353494 237989 353546 237995
rect 353110 233015 353162 233021
rect 353110 232957 353162 232963
rect 353110 227761 353162 227767
rect 353110 227703 353162 227709
rect 352534 223395 352586 223401
rect 352534 223337 352586 223343
rect 352354 221468 352416 221496
rect 353122 221482 353150 227703
rect 354082 223253 354110 239672
rect 354226 239404 354254 239686
rect 354624 239672 354878 239700
rect 354178 239376 354254 239404
rect 353878 223247 353930 223253
rect 353878 223189 353930 223195
rect 354070 223247 354122 223253
rect 354070 223189 354122 223195
rect 353890 221496 353918 223189
rect 354178 222999 354206 239376
rect 354262 235531 354314 235537
rect 354262 235473 354314 235479
rect 354274 232059 354302 235473
rect 354644 234978 354700 234987
rect 354644 234913 354700 234922
rect 354262 232053 354314 232059
rect 354262 231995 354314 232001
rect 354658 226953 354686 234913
rect 354850 229543 354878 239672
rect 354946 233835 354974 239686
rect 355344 239672 355646 239700
rect 354934 233829 354986 233835
rect 354934 233771 354986 233777
rect 355318 232201 355370 232207
rect 355318 232143 355370 232149
rect 354838 229537 354890 229543
rect 354838 229479 354890 229485
rect 354550 226947 354602 226953
rect 354550 226889 354602 226895
rect 354646 226947 354698 226953
rect 354646 226889 354698 226895
rect 354164 222990 354220 222999
rect 354164 222925 354220 222934
rect 353856 221468 353918 221496
rect 354562 221496 354590 226889
rect 354562 221468 354624 221496
rect 355330 221482 355358 232143
rect 355618 222703 355646 239672
rect 355714 237905 355742 239686
rect 356064 239672 356318 239700
rect 356544 239672 356798 239700
rect 355702 237899 355754 237905
rect 355702 237841 355754 237847
rect 356290 232873 356318 239672
rect 356770 234987 356798 239672
rect 356866 236171 356894 239686
rect 356852 236162 356908 236171
rect 356852 236097 356908 236106
rect 357154 236055 357182 239765
rect 377302 239749 377354 239755
rect 357142 236049 357194 236055
rect 357142 235991 357194 235997
rect 356756 234978 356812 234987
rect 356756 234913 356812 234922
rect 356278 232867 356330 232873
rect 356278 232809 356330 232815
rect 356086 232571 356138 232577
rect 356086 232513 356138 232519
rect 355604 222694 355660 222703
rect 355604 222629 355660 222638
rect 356098 221792 356126 232513
rect 357250 222851 357278 239686
rect 357526 237751 357578 237757
rect 357526 237693 357578 237699
rect 357430 229315 357482 229321
rect 357430 229257 357482 229263
rect 357442 229025 357470 229257
rect 357538 229025 357566 237693
rect 357634 229469 357662 239686
rect 358018 235611 358046 239686
rect 358368 239672 358622 239700
rect 358752 239672 359006 239700
rect 358006 235605 358058 235611
rect 358006 235547 358058 235553
rect 358294 232275 358346 232281
rect 358294 232217 358346 232223
rect 357622 229463 357674 229469
rect 357622 229405 357674 229411
rect 357430 229019 357482 229025
rect 357430 228961 357482 228967
rect 357526 229019 357578 229025
rect 357526 228961 357578 228967
rect 357622 227021 357674 227027
rect 357622 226963 357674 226969
rect 357236 222842 357292 222851
rect 357236 222777 357292 222786
rect 356854 222359 356906 222365
rect 356854 222301 356906 222307
rect 356098 221764 356174 221792
rect 356146 221482 356174 221764
rect 356866 221482 356894 222301
rect 357634 221482 357662 226963
rect 358306 221792 358334 232217
rect 358594 224627 358622 239672
rect 358978 230103 359006 239672
rect 359074 232799 359102 239686
rect 359062 232793 359114 232799
rect 359062 232735 359114 232741
rect 358964 230094 359020 230103
rect 358964 230029 359020 230038
rect 359158 227983 359210 227989
rect 359158 227925 359210 227931
rect 358580 224618 358636 224627
rect 358580 224553 358636 224562
rect 358306 221764 358382 221792
rect 358354 221482 358382 221764
rect 359170 221482 359198 227925
rect 359458 224479 359486 239686
rect 359842 236174 359870 239686
rect 359746 236146 359870 236174
rect 359444 224470 359500 224479
rect 359444 224405 359500 224414
rect 359746 224331 359774 236146
rect 359828 229058 359884 229067
rect 359828 228993 359884 229002
rect 359926 229019 359978 229025
rect 359842 227027 359870 228993
rect 359926 228961 359978 228967
rect 359830 227021 359882 227027
rect 359830 226963 359882 226969
rect 359732 224322 359788 224331
rect 359732 224257 359788 224266
rect 359938 221482 359966 228961
rect 360322 224183 360350 239686
rect 360672 239672 360926 239700
rect 361056 239672 361310 239700
rect 360898 228771 360926 239672
rect 361282 233983 361310 239672
rect 361378 236174 361406 239686
rect 361762 237757 361790 239686
rect 361750 237751 361802 237757
rect 361750 237693 361802 237699
rect 361378 236146 361502 236174
rect 361270 233977 361322 233983
rect 361270 233919 361322 233925
rect 361366 232349 361418 232355
rect 361366 232291 361418 232297
rect 360884 228762 360940 228771
rect 360884 228697 360940 228706
rect 360598 227095 360650 227101
rect 360598 227037 360650 227043
rect 360308 224174 360364 224183
rect 360308 224109 360364 224118
rect 360610 221792 360638 227037
rect 360610 221764 360686 221792
rect 360658 221482 360686 221764
rect 361378 221482 361406 232291
rect 361474 224035 361502 236146
rect 362146 232651 362174 239686
rect 362530 235019 362558 239686
rect 362880 239672 363134 239700
rect 363264 239672 363518 239700
rect 363106 237831 363134 239672
rect 363094 237825 363146 237831
rect 363094 237767 363146 237773
rect 362614 235383 362666 235389
rect 362614 235325 362666 235331
rect 362422 235013 362474 235019
rect 362422 234955 362474 234961
rect 362518 235013 362570 235019
rect 362518 234955 362570 234961
rect 362134 232645 362186 232651
rect 362134 232587 362186 232593
rect 362134 230721 362186 230727
rect 362134 230663 362186 230669
rect 361460 224026 361516 224035
rect 361460 223961 361516 223970
rect 362146 221482 362174 230663
rect 362434 224733 362462 234955
rect 362626 230727 362654 235325
rect 363490 233687 363518 239672
rect 363478 233681 363530 233687
rect 363478 233623 363530 233629
rect 362614 230721 362666 230727
rect 362614 230663 362666 230669
rect 363586 230251 363614 239686
rect 363670 237677 363722 237683
rect 363670 237619 363722 237625
rect 363572 230242 363628 230251
rect 363572 230177 363628 230186
rect 362804 229206 362860 229215
rect 362804 229141 362860 229150
rect 362818 224881 362846 229141
rect 363682 227268 363710 237619
rect 364066 233803 364094 239686
rect 364450 237683 364478 239686
rect 364800 239672 365054 239700
rect 365184 239672 365438 239700
rect 365568 239672 365726 239700
rect 364438 237677 364490 237683
rect 364438 237619 364490 237625
rect 364052 233794 364108 233803
rect 364052 233729 364108 233738
rect 364150 233681 364202 233687
rect 364150 233623 364202 233629
rect 363010 227240 363710 227268
rect 362806 224875 362858 224881
rect 362806 224817 362858 224823
rect 362422 224727 362474 224733
rect 362422 224669 362474 224675
rect 363010 221792 363038 227240
rect 363670 224801 363722 224807
rect 363670 224743 363722 224749
rect 362962 221764 363038 221792
rect 362962 221482 362990 221764
rect 363682 221482 363710 224743
rect 364162 223887 364190 233623
rect 365026 232429 365054 239672
rect 365410 232577 365438 239672
rect 365698 233359 365726 239672
rect 365890 237609 365918 239686
rect 365878 237603 365930 237609
rect 365878 237545 365930 237551
rect 365684 233350 365740 233359
rect 365684 233285 365740 233294
rect 365398 232571 365450 232577
rect 365398 232513 365450 232519
rect 366274 232503 366302 239686
rect 366262 232497 366314 232503
rect 366262 232439 366314 232445
rect 365014 232423 365066 232429
rect 365014 232365 365066 232371
rect 364438 232127 364490 232133
rect 364438 232069 364490 232075
rect 364148 223878 364204 223887
rect 364148 223813 364204 223822
rect 364450 221482 364478 232069
rect 365110 231239 365162 231245
rect 365110 231181 365162 231187
rect 365014 230795 365066 230801
rect 365014 230737 365066 230743
rect 365026 221792 365054 230737
rect 365122 226879 365150 231181
rect 366658 229955 366686 239686
rect 367008 239672 367262 239700
rect 367392 239672 367646 239700
rect 367872 239672 368126 239700
rect 366742 236789 366794 236795
rect 366742 236731 366794 236737
rect 366644 229946 366700 229955
rect 366644 229881 366700 229890
rect 365684 228910 365740 228919
rect 365684 228845 365740 228854
rect 365110 226873 365162 226879
rect 365110 226815 365162 226821
rect 365698 225769 365726 228845
rect 366754 228489 366782 236731
rect 367234 235579 367262 239672
rect 367220 235570 367276 235579
rect 367220 235505 367276 235514
rect 367126 232053 367178 232059
rect 367126 231995 367178 232001
rect 367138 230801 367166 231995
rect 367414 231979 367466 231985
rect 367414 231921 367466 231927
rect 367126 230795 367178 230801
rect 367126 230737 367178 230743
rect 365890 228461 366782 228489
rect 365686 225763 365738 225769
rect 365686 225705 365738 225711
rect 365026 221764 365198 221792
rect 365170 221482 365198 221764
rect 365890 221482 365918 228461
rect 366742 226799 366794 226805
rect 366742 226741 366794 226747
rect 366754 221482 366782 226741
rect 367426 221792 367454 231921
rect 367618 223739 367646 239672
rect 368098 232207 368126 239672
rect 368194 232355 368222 239686
rect 368578 239089 368606 239686
rect 368566 239083 368618 239089
rect 368566 239025 368618 239031
rect 368962 236467 368990 239686
rect 369312 239672 369566 239700
rect 369696 239672 369950 239700
rect 370080 239672 370334 239700
rect 368948 236458 369004 236467
rect 368948 236393 369004 236402
rect 368854 235087 368906 235093
rect 368854 235029 368906 235035
rect 368182 232349 368234 232355
rect 368182 232291 368234 232297
rect 368086 232201 368138 232207
rect 368086 232143 368138 232149
rect 368660 231870 368716 231879
rect 368660 231805 368716 231814
rect 368182 230499 368234 230505
rect 368182 230441 368234 230447
rect 367604 223730 367660 223739
rect 367604 223665 367660 223674
rect 367426 221764 367502 221792
rect 367474 221482 367502 221764
rect 368194 221482 368222 230441
rect 368674 225219 368702 231805
rect 368866 227989 368894 235029
rect 369538 232281 369566 239672
rect 369526 232275 369578 232281
rect 369526 232217 369578 232223
rect 369922 229395 369950 239672
rect 370306 233909 370334 239672
rect 370402 236763 370430 239686
rect 370486 236863 370538 236869
rect 370486 236805 370538 236811
rect 370388 236754 370444 236763
rect 370388 236689 370444 236698
rect 370294 233903 370346 233909
rect 370294 233845 370346 233851
rect 370390 231905 370442 231911
rect 370390 231847 370442 231853
rect 369526 229389 369578 229395
rect 369526 229331 369578 229337
rect 369910 229389 369962 229395
rect 369910 229331 369962 229337
rect 368950 229019 369002 229025
rect 368950 228961 369002 228967
rect 368854 227983 368906 227989
rect 368854 227925 368906 227931
rect 368660 225210 368716 225219
rect 368660 225145 368716 225154
rect 368962 221482 368990 228961
rect 369430 224949 369482 224955
rect 369430 224891 369482 224897
rect 369442 224733 369470 224891
rect 369538 224733 369566 229331
rect 370402 227534 370430 231847
rect 370498 229025 370526 236805
rect 370786 232915 370814 239686
rect 371170 233063 371198 239686
rect 371616 239672 371870 239700
rect 372000 239672 372254 239700
rect 371842 236055 371870 239672
rect 372226 237059 372254 239672
rect 372212 237050 372268 237059
rect 372212 236985 372268 236994
rect 371830 236049 371882 236055
rect 371830 235991 371882 235997
rect 371638 234199 371690 234205
rect 371638 234141 371690 234147
rect 371156 233054 371212 233063
rect 371156 232989 371212 232998
rect 370772 232906 370828 232915
rect 370772 232841 370828 232850
rect 371254 229241 371306 229247
rect 371254 229183 371306 229189
rect 370486 229019 370538 229025
rect 370486 228961 370538 228967
rect 370402 227506 370526 227534
rect 369622 227169 369674 227175
rect 369622 227111 369674 227117
rect 369430 224727 369482 224733
rect 369430 224669 369482 224675
rect 369526 224727 369578 224733
rect 369526 224669 369578 224675
rect 369634 221792 369662 227111
rect 369634 221764 369710 221792
rect 369682 221482 369710 221764
rect 370498 221482 370526 227506
rect 371266 221482 371294 229183
rect 371542 229093 371594 229099
rect 371542 229035 371594 229041
rect 371554 224807 371582 229035
rect 371542 224801 371594 224807
rect 371542 224743 371594 224749
rect 371650 222365 371678 234141
rect 372322 232059 372350 239686
rect 372706 232133 372734 239686
rect 372694 232127 372746 232133
rect 372694 232069 372746 232075
rect 372310 232053 372362 232059
rect 372310 231995 372362 232001
rect 373090 229807 373118 239686
rect 373474 236911 373502 239686
rect 373824 239672 374078 239700
rect 374208 239672 374366 239700
rect 373460 236902 373516 236911
rect 373460 236837 373516 236846
rect 374050 232767 374078 239672
rect 374036 232758 374092 232767
rect 374036 232693 374092 232702
rect 373462 231831 373514 231837
rect 373462 231773 373514 231779
rect 373076 229798 373132 229807
rect 373076 229733 373132 229742
rect 372694 226799 372746 226805
rect 372694 226741 372746 226747
rect 371926 222507 371978 222513
rect 371926 222449 371978 222455
rect 371638 222359 371690 222365
rect 371638 222301 371690 222307
rect 371938 221792 371966 222449
rect 371938 221764 372014 221792
rect 371986 221482 372014 221764
rect 372706 221482 372734 226741
rect 373474 221482 373502 231773
rect 374230 230647 374282 230653
rect 374230 230589 374282 230595
rect 374242 221792 374270 230589
rect 374338 229247 374366 239672
rect 374422 239601 374474 239607
rect 374422 239543 374474 239549
rect 374434 236129 374462 239543
rect 374422 236123 374474 236129
rect 374422 236065 374474 236071
rect 374530 231911 374558 239686
rect 374914 236319 374942 239686
rect 374900 236310 374956 236319
rect 374900 236245 374956 236254
rect 375394 232619 375422 239686
rect 375380 232610 375436 232619
rect 375380 232545 375436 232554
rect 375778 231985 375806 239686
rect 376128 239672 376382 239700
rect 376512 239672 376766 239700
rect 377302 239691 377354 239697
rect 376354 236129 376382 239672
rect 376342 236123 376394 236129
rect 376342 236065 376394 236071
rect 375766 231979 375818 231985
rect 375766 231921 375818 231927
rect 374518 231905 374570 231911
rect 374518 231847 374570 231853
rect 374614 231461 374666 231467
rect 374614 231403 374666 231409
rect 374518 229315 374570 229321
rect 374518 229257 374570 229263
rect 374326 229241 374378 229247
rect 374326 229183 374378 229189
rect 374422 229167 374474 229173
rect 374422 229109 374474 229115
rect 374434 226657 374462 229109
rect 374422 226651 374474 226657
rect 374422 226593 374474 226599
rect 374530 225843 374558 229257
rect 374626 226805 374654 231403
rect 375766 227539 375818 227545
rect 375766 227481 375818 227487
rect 374614 226799 374666 226805
rect 374614 226741 374666 226747
rect 374518 225837 374570 225843
rect 374518 225779 374570 225785
rect 374998 222433 375050 222439
rect 374998 222375 375050 222381
rect 374242 221764 374318 221792
rect 374290 221482 374318 221764
rect 375010 221482 375038 222375
rect 375778 221482 375806 227481
rect 376438 224727 376490 224733
rect 376438 224669 376490 224675
rect 376450 221792 376478 224669
rect 376738 223443 376766 239672
rect 376834 229099 376862 239686
rect 377110 230573 377162 230579
rect 377110 230515 377162 230521
rect 376822 229093 376874 229099
rect 376822 229035 376874 229041
rect 377122 227534 377150 230515
rect 377218 229173 377246 239686
rect 377314 233317 377342 239691
rect 377302 233311 377354 233317
rect 377302 233253 377354 233259
rect 377206 229167 377258 229173
rect 377206 229109 377258 229115
rect 377122 227506 377246 227534
rect 376724 223434 376780 223443
rect 376724 223369 376780 223378
rect 376450 221764 376526 221792
rect 376498 221482 376526 221764
rect 377218 221482 377246 227506
rect 377602 223591 377630 239686
rect 378000 239672 378206 239700
rect 378336 239672 378590 239700
rect 378720 239672 378974 239700
rect 377972 236606 378028 236615
rect 377972 236541 378028 236550
rect 377986 236319 378014 236541
rect 378178 236319 378206 239672
rect 377972 236310 378028 236319
rect 377972 236245 378028 236254
rect 378164 236310 378220 236319
rect 378164 236245 378220 236254
rect 378562 234205 378590 239672
rect 378550 234199 378602 234205
rect 378550 234141 378602 234147
rect 378946 231837 378974 239672
rect 379138 234543 379166 239686
rect 379536 239672 379838 239700
rect 379810 236721 379838 239672
rect 379798 236715 379850 236721
rect 379798 236657 379850 236663
rect 379124 234534 379180 234543
rect 379124 234469 379180 234478
rect 378934 231831 378986 231837
rect 378934 231773 378986 231779
rect 379906 229659 379934 239686
rect 380256 239672 380510 239700
rect 381024 239672 381278 239700
rect 380084 233350 380140 233359
rect 380084 233285 380140 233294
rect 379990 231387 380042 231393
rect 379990 231329 380042 231335
rect 379892 229650 379948 229659
rect 379892 229585 379948 229594
rect 378742 226725 378794 226731
rect 378742 226667 378794 226673
rect 378070 226429 378122 226435
rect 378070 226371 378122 226377
rect 377588 223582 377644 223591
rect 377588 223517 377644 223526
rect 378082 221482 378110 226371
rect 378754 221792 378782 226667
rect 379894 226429 379946 226435
rect 379894 226371 379946 226377
rect 379906 226065 379934 226371
rect 380002 226065 380030 231329
rect 380098 229469 380126 233285
rect 380182 230869 380234 230875
rect 380182 230811 380234 230817
rect 380086 229463 380138 229469
rect 380086 229405 380138 229411
rect 380086 228501 380138 228507
rect 380086 228443 380138 228449
rect 379894 226059 379946 226065
rect 379894 226001 379946 226007
rect 379990 226059 380042 226065
rect 379990 226001 380042 226007
rect 380098 224807 380126 228443
rect 379510 224801 379562 224807
rect 379510 224743 379562 224749
rect 380086 224801 380138 224807
rect 380086 224743 380138 224749
rect 378754 221764 378830 221792
rect 378802 221482 378830 221764
rect 379522 221482 379550 224743
rect 380194 224160 380222 230811
rect 380482 229025 380510 239672
rect 380470 229019 380522 229025
rect 380470 228961 380522 228967
rect 380278 228353 380330 228359
rect 380278 228295 380330 228301
rect 380290 226731 380318 228295
rect 380278 226725 380330 226731
rect 380278 226667 380330 226673
rect 380194 224132 380318 224160
rect 380290 221482 380318 224132
rect 381250 223295 381278 239672
rect 381346 229511 381374 239686
rect 381730 232471 381758 239686
rect 382114 234395 382142 239686
rect 382560 239672 382622 239700
rect 382594 236319 382622 239672
rect 382690 239672 382944 239700
rect 383328 239672 383582 239700
rect 382388 236310 382444 236319
rect 382388 236245 382444 236254
rect 382580 236310 382636 236319
rect 382580 236245 382636 236254
rect 382402 236203 382430 236245
rect 382390 236197 382442 236203
rect 382390 236139 382442 236145
rect 382100 234386 382156 234395
rect 382100 234321 382156 234330
rect 381716 232462 381772 232471
rect 381716 232397 381772 232406
rect 382690 232027 382718 239672
rect 382870 232941 382922 232947
rect 382870 232883 382922 232889
rect 382676 232018 382732 232027
rect 382676 231953 382732 231962
rect 381332 229502 381388 229511
rect 381332 229437 381388 229446
rect 381814 227465 381866 227471
rect 381814 227407 381866 227413
rect 381236 223286 381292 223295
rect 381236 223221 381292 223230
rect 381046 222729 381098 222735
rect 381046 222671 381098 222677
rect 381058 221496 381086 222671
rect 381058 221468 381120 221496
rect 381826 221482 381854 227407
rect 382582 225837 382634 225843
rect 382582 225779 382634 225785
rect 382594 221496 382622 225779
rect 382882 224733 382910 232883
rect 383554 229363 383582 239672
rect 383650 233687 383678 239686
rect 384048 239672 384350 239700
rect 383638 233681 383690 233687
rect 383638 233623 383690 233629
rect 383540 229354 383596 229363
rect 383540 229289 383596 229298
rect 382966 228649 383018 228655
rect 382966 228591 383018 228597
rect 382978 225991 383006 228591
rect 383254 228205 383306 228211
rect 383254 228147 383306 228153
rect 382966 225985 383018 225991
rect 382966 225927 383018 225933
rect 382870 224727 382922 224733
rect 382870 224669 382922 224675
rect 382560 221468 382622 221496
rect 383266 221496 383294 228147
rect 384022 227391 384074 227397
rect 384022 227333 384074 227339
rect 383266 221468 383328 221496
rect 384034 221482 384062 227333
rect 384322 223147 384350 239672
rect 384418 229215 384446 239686
rect 384768 239672 385022 239700
rect 385152 239672 385310 239700
rect 384994 232323 385022 239672
rect 384980 232314 385036 232323
rect 384980 232249 385036 232258
rect 385282 232175 385310 239672
rect 385366 239675 385418 239681
rect 385536 239672 385790 239700
rect 385366 239617 385418 239623
rect 385378 235167 385406 239617
rect 385366 235161 385418 235167
rect 385366 235103 385418 235109
rect 385268 232166 385324 232175
rect 385268 232101 385324 232110
rect 384404 229206 384460 229215
rect 384404 229141 384460 229150
rect 385558 226651 385610 226657
rect 385558 226593 385610 226599
rect 384790 226503 384842 226509
rect 384790 226445 384842 226451
rect 384308 223138 384364 223147
rect 384308 223073 384364 223082
rect 384802 221792 384830 226445
rect 384802 221764 384878 221792
rect 384850 221482 384878 221764
rect 385570 221482 385598 226593
rect 385762 226509 385790 239672
rect 385858 236023 385886 239686
rect 385844 236014 385900 236023
rect 385844 235949 385900 235958
rect 386230 233755 386282 233761
rect 386230 233697 386282 233703
rect 385846 231313 385898 231319
rect 385846 231255 385898 231261
rect 385750 226503 385802 226509
rect 385750 226445 385802 226451
rect 385858 225843 385886 231255
rect 385846 225837 385898 225843
rect 385846 225779 385898 225785
rect 386242 222439 386270 233697
rect 386338 233317 386366 239686
rect 386722 235981 386750 239686
rect 387072 239672 387326 239700
rect 387456 239672 387710 239700
rect 386998 236863 387050 236869
rect 386998 236805 387050 236811
rect 387010 236319 387038 236805
rect 386996 236310 387052 236319
rect 386996 236245 387052 236254
rect 387298 236174 387326 239672
rect 387380 236902 387436 236911
rect 387380 236837 387436 236846
rect 387572 236902 387628 236911
rect 387572 236837 387574 236846
rect 387394 236467 387422 236837
rect 387626 236837 387628 236846
rect 387574 236805 387626 236811
rect 387380 236458 387436 236467
rect 387380 236393 387436 236402
rect 387298 236146 387422 236174
rect 386710 235975 386762 235981
rect 386710 235917 386762 235923
rect 387286 234791 387338 234797
rect 387286 234733 387338 234739
rect 386326 233311 386378 233317
rect 386326 233253 386378 233259
rect 387298 230875 387326 234733
rect 387286 230869 387338 230875
rect 387286 230811 387338 230817
rect 387394 225917 387422 236146
rect 387682 235167 387710 239672
rect 387670 235161 387722 235167
rect 387670 235103 387722 235109
rect 387778 227767 387806 239686
rect 387766 227761 387818 227767
rect 387766 227703 387818 227709
rect 388162 226435 388190 239686
rect 388546 227397 388574 239686
rect 388726 233311 388778 233317
rect 388726 233253 388778 233259
rect 388534 227391 388586 227397
rect 388534 227333 388586 227339
rect 387766 226429 387818 226435
rect 387766 226371 387818 226377
rect 388150 226429 388202 226435
rect 388150 226371 388202 226377
rect 386998 225911 387050 225917
rect 386998 225853 387050 225859
rect 387382 225911 387434 225917
rect 387382 225853 387434 225859
rect 386326 224727 386378 224733
rect 386326 224669 386378 224675
rect 386230 222433 386282 222439
rect 386230 222375 386282 222381
rect 386338 221482 386366 224669
rect 387010 221792 387038 225853
rect 387010 221764 387086 221792
rect 387058 221482 387086 221764
rect 387778 221482 387806 226371
rect 388738 225991 388766 233253
rect 388930 227323 388958 239686
rect 389280 239672 389534 239700
rect 389664 239672 389918 239700
rect 389506 227545 389534 239672
rect 389890 235875 389918 239672
rect 389876 235866 389932 235875
rect 389876 235801 389932 235810
rect 389494 227539 389546 227545
rect 389494 227481 389546 227487
rect 388918 227317 388970 227323
rect 388918 227259 388970 227265
rect 390082 227175 390110 239686
rect 390466 227471 390494 239686
rect 390742 236345 390794 236351
rect 390742 236287 390794 236293
rect 390754 235727 390782 236287
rect 390740 235718 390796 235727
rect 390740 235653 390796 235662
rect 390454 227465 390506 227471
rect 390454 227407 390506 227413
rect 390070 227169 390122 227175
rect 390070 227111 390122 227117
rect 390850 227101 390878 239686
rect 390838 227095 390890 227101
rect 390838 227037 390890 227043
rect 391234 226847 391262 239686
rect 391584 239672 391646 239700
rect 391968 239672 392222 239700
rect 391618 226995 391646 239672
rect 392194 235315 392222 239672
rect 392182 235309 392234 235315
rect 392182 235251 392234 235257
rect 391702 235235 391754 235241
rect 391702 235177 391754 235183
rect 391714 228359 391742 235177
rect 391702 228353 391754 228359
rect 391702 228295 391754 228301
rect 391604 226986 391660 226995
rect 391604 226921 391660 226930
rect 392182 226947 392234 226953
rect 392182 226889 392234 226895
rect 391220 226838 391276 226847
rect 391220 226773 391276 226782
rect 391510 226799 391562 226805
rect 391510 226741 391562 226747
rect 390070 226577 390122 226583
rect 390070 226519 390122 226525
rect 388630 225985 388682 225991
rect 388630 225927 388682 225933
rect 388726 225985 388778 225991
rect 388726 225927 388778 225933
rect 388642 224900 388670 225927
rect 388642 224872 388766 224900
rect 388738 224807 388766 224872
rect 388630 224801 388682 224807
rect 388630 224743 388682 224749
rect 388726 224801 388778 224807
rect 388726 224743 388778 224749
rect 389302 224801 389354 224807
rect 389302 224743 389354 224749
rect 388642 221482 388670 224743
rect 389314 221792 389342 224743
rect 389314 221764 389390 221792
rect 389362 221482 389390 221764
rect 390082 221482 390110 226519
rect 390838 226355 390890 226361
rect 390838 226297 390890 226303
rect 390850 221482 390878 226297
rect 391522 221792 391550 226741
rect 392194 226583 392222 226889
rect 392182 226577 392234 226583
rect 392182 226519 392234 226525
rect 392290 224807 392318 239686
rect 392470 234865 392522 234871
rect 392470 234807 392522 234813
rect 392482 228285 392510 234807
rect 392374 228279 392426 228285
rect 392374 228221 392426 228227
rect 392470 228279 392522 228285
rect 392470 228221 392522 228227
rect 392278 224801 392330 224807
rect 392278 224743 392330 224749
rect 391522 221764 391598 221792
rect 391570 221482 391598 221764
rect 392386 221482 392414 228221
rect 392674 227027 392702 239686
rect 393058 235727 393086 239686
rect 393044 235718 393100 235727
rect 393044 235653 393100 235662
rect 393442 235389 393470 239686
rect 393888 239672 394142 239700
rect 394272 239672 394526 239700
rect 394608 239672 394910 239700
rect 393430 235383 393482 235389
rect 393430 235325 393482 235331
rect 392662 227021 392714 227027
rect 392662 226963 392714 226969
rect 393142 226947 393194 226953
rect 393142 226889 393194 226895
rect 393154 221482 393182 226889
rect 394114 226699 394142 239672
rect 394100 226690 394156 226699
rect 394100 226625 394156 226634
rect 394498 226551 394526 239672
rect 394678 239453 394730 239459
rect 394678 239395 394730 239401
rect 394582 236271 394634 236277
rect 394582 236213 394634 236219
rect 394594 233613 394622 236213
rect 394690 235019 394718 239395
rect 394882 235093 394910 239672
rect 394978 235537 395006 239686
rect 395376 239672 395582 239700
rect 395712 239672 395966 239700
rect 396096 239672 396350 239700
rect 396480 239672 396734 239700
rect 394966 235531 395018 235537
rect 394966 235473 395018 235479
rect 395062 235457 395114 235463
rect 395062 235399 395114 235405
rect 394870 235087 394922 235093
rect 394870 235029 394922 235035
rect 394678 235013 394730 235019
rect 394678 234955 394730 234961
rect 394774 234939 394826 234945
rect 394774 234881 394826 234887
rect 394678 234717 394730 234723
rect 394678 234659 394730 234665
rect 394582 233607 394634 233613
rect 394582 233549 394634 233555
rect 394690 228211 394718 234659
rect 394786 231245 394814 234881
rect 394870 234051 394922 234057
rect 394870 233993 394922 233999
rect 394774 231239 394826 231245
rect 394774 231181 394826 231187
rect 394678 228205 394730 228211
rect 394678 228147 394730 228153
rect 394484 226542 394540 226551
rect 394484 226477 394540 226486
rect 394582 226059 394634 226065
rect 394582 226001 394634 226007
rect 393814 225763 393866 225769
rect 393814 225705 393866 225711
rect 393826 221792 393854 225705
rect 393826 221764 393902 221792
rect 393874 221482 393902 221764
rect 394594 221482 394622 226001
rect 394882 222513 394910 233993
rect 395074 231319 395102 235399
rect 395062 231313 395114 231319
rect 395062 231255 395114 231261
rect 395350 230943 395402 230949
rect 395350 230885 395402 230891
rect 394870 222507 394922 222513
rect 394870 222449 394922 222455
rect 395362 221482 395390 230885
rect 395554 226879 395582 239672
rect 395938 233317 395966 239672
rect 396322 235241 396350 239672
rect 396310 235235 396362 235241
rect 396310 235177 396362 235183
rect 396706 234057 396734 239672
rect 396802 235463 396830 239686
rect 396980 237050 397036 237059
rect 396980 236985 397036 236994
rect 396994 236795 397022 236985
rect 397076 236902 397132 236911
rect 397076 236837 397078 236846
rect 397130 236837 397132 236846
rect 397078 236805 397130 236811
rect 396982 236789 397034 236795
rect 396982 236731 397034 236737
rect 396790 235457 396842 235463
rect 396790 235399 396842 235405
rect 396694 234051 396746 234057
rect 396694 233993 396746 233999
rect 395926 233311 395978 233317
rect 395926 233253 395978 233259
rect 396214 227761 396266 227767
rect 396214 227703 396266 227709
rect 395542 226873 395594 226879
rect 395542 226815 395594 226821
rect 396118 226799 396170 226805
rect 396118 226741 396170 226747
rect 396130 221792 396158 226741
rect 396226 225769 396254 227703
rect 397186 226657 397214 239686
rect 397680 239672 397886 239700
rect 398016 239672 398270 239700
rect 398400 239672 398654 239700
rect 398784 239672 399038 239700
rect 399120 239672 399422 239700
rect 397750 239379 397802 239385
rect 397750 239321 397802 239327
rect 397652 237050 397708 237059
rect 397652 236985 397708 236994
rect 397666 236869 397694 236985
rect 397654 236863 397706 236869
rect 397654 236805 397706 236811
rect 397364 236310 397420 236319
rect 397364 236245 397420 236254
rect 397378 236203 397406 236245
rect 397366 236197 397418 236203
rect 397366 236139 397418 236145
rect 397762 235579 397790 239321
rect 397748 235570 397804 235579
rect 397748 235505 397804 235514
rect 397366 232719 397418 232725
rect 397366 232661 397418 232667
rect 397378 232596 397406 232661
rect 397378 232568 397502 232596
rect 397174 226651 397226 226657
rect 397174 226593 397226 226599
rect 396214 225763 396266 225769
rect 396214 225705 396266 225711
rect 396886 225097 396938 225103
rect 396886 225039 396938 225045
rect 396130 221764 396206 221792
rect 396178 221482 396206 221764
rect 396898 221482 396926 225039
rect 397474 224733 397502 232568
rect 397654 226725 397706 226731
rect 397654 226667 397706 226673
rect 397462 224727 397514 224733
rect 397462 224669 397514 224675
rect 397666 221482 397694 226667
rect 397858 226287 397886 239672
rect 398036 236902 398092 236911
rect 398036 236837 398038 236846
rect 398090 236837 398092 236846
rect 398038 236805 398090 236811
rect 398242 233835 398270 239672
rect 398324 236902 398380 236911
rect 398324 236837 398380 236846
rect 398338 236721 398366 236837
rect 398326 236715 398378 236721
rect 398326 236657 398378 236663
rect 398626 234945 398654 239672
rect 399010 235019 399038 239672
rect 398998 235013 399050 235019
rect 398998 234955 399050 234961
rect 398614 234939 398666 234945
rect 398614 234881 398666 234887
rect 399190 234199 399242 234205
rect 399190 234141 399242 234147
rect 398230 233829 398282 233835
rect 398230 233771 398282 233777
rect 399202 232725 399230 234141
rect 399190 232719 399242 232725
rect 399190 232661 399242 232667
rect 398326 228057 398378 228063
rect 398326 227999 398378 228005
rect 397846 226281 397898 226287
rect 397846 226223 397898 226229
rect 398338 221792 398366 227999
rect 398902 227243 398954 227249
rect 398902 227185 398954 227191
rect 398806 226503 398858 226509
rect 398806 226445 398858 226451
rect 398818 226065 398846 226445
rect 398914 226435 398942 227185
rect 398902 226429 398954 226435
rect 398902 226371 398954 226377
rect 398806 226059 398858 226065
rect 398806 226001 398858 226007
rect 398902 225985 398954 225991
rect 398722 225945 398902 225973
rect 398722 225917 398750 225945
rect 398902 225927 398954 225933
rect 398710 225911 398762 225917
rect 398710 225853 398762 225859
rect 398614 225837 398666 225843
rect 398614 225779 398666 225785
rect 398626 225103 398654 225779
rect 399394 225103 399422 239672
rect 399490 228919 399518 239686
rect 399874 235579 399902 239686
rect 400224 239672 400286 239700
rect 400608 239672 400862 239700
rect 400992 239672 401246 239700
rect 399860 235570 399916 235579
rect 399860 235505 399916 235514
rect 400150 234125 400202 234131
rect 400150 234067 400202 234073
rect 400162 231393 400190 234067
rect 400258 233951 400286 239672
rect 400342 236197 400394 236203
rect 400342 236139 400394 236145
rect 400354 235611 400382 236139
rect 400342 235605 400394 235611
rect 400342 235547 400394 235553
rect 400244 233942 400300 233951
rect 400244 233877 400300 233886
rect 400246 233311 400298 233317
rect 400246 233253 400298 233259
rect 400150 231387 400202 231393
rect 400150 231329 400202 231335
rect 400258 229067 400286 233253
rect 400244 229058 400300 229067
rect 400244 228993 400300 229002
rect 399476 228910 399532 228919
rect 399476 228845 399532 228854
rect 400834 226805 400862 239672
rect 401110 234273 401162 234279
rect 401110 234215 401162 234221
rect 400822 226799 400874 226805
rect 400822 226741 400874 226747
rect 400246 226281 400298 226287
rect 400246 226223 400298 226229
rect 400258 225917 400286 226223
rect 400246 225911 400298 225917
rect 400246 225853 400298 225859
rect 399958 225171 400010 225177
rect 399958 225113 400010 225119
rect 398614 225097 398666 225103
rect 398614 225039 398666 225045
rect 399382 225097 399434 225103
rect 399382 225039 399434 225045
rect 399094 225023 399146 225029
rect 399094 224965 399146 224971
rect 398338 221764 398414 221792
rect 398386 221482 398414 221764
rect 399106 221482 399134 224965
rect 399970 221482 399998 225113
rect 400630 224727 400682 224733
rect 400630 224669 400682 224675
rect 400642 221792 400670 224669
rect 401122 222735 401150 234215
rect 401218 233317 401246 239672
rect 401410 235431 401438 239686
rect 401396 235422 401452 235431
rect 401396 235357 401452 235366
rect 401794 234131 401822 239686
rect 401782 234125 401834 234131
rect 401782 234067 401834 234073
rect 401206 233311 401258 233317
rect 401206 233253 401258 233259
rect 401398 231017 401450 231023
rect 401398 230959 401450 230965
rect 401110 222729 401162 222735
rect 401110 222671 401162 222677
rect 400642 221764 400718 221792
rect 400690 221482 400718 221764
rect 401410 221482 401438 230959
rect 402178 226731 402206 239686
rect 402528 239672 402590 239700
rect 402166 226725 402218 226731
rect 402166 226667 402218 226673
rect 402562 226583 402590 239672
rect 402658 239672 402912 239700
rect 403248 239672 403550 239700
rect 402658 235283 402686 239672
rect 402644 235274 402700 235283
rect 402644 235209 402700 235218
rect 403124 234978 403180 234987
rect 403124 234913 403180 234922
rect 403138 231467 403166 234913
rect 403522 234205 403550 239672
rect 403618 234871 403646 239686
rect 404002 234987 404030 239686
rect 403988 234978 404044 234987
rect 403988 234913 404044 234922
rect 403606 234865 403658 234871
rect 403606 234807 403658 234813
rect 403510 234199 403562 234205
rect 403510 234141 403562 234147
rect 403126 231461 403178 231467
rect 403126 231403 403178 231409
rect 403702 227613 403754 227619
rect 403702 227555 403754 227561
rect 402550 226577 402602 226583
rect 402550 226519 402602 226525
rect 402838 226355 402890 226361
rect 402838 226297 402890 226303
rect 402166 224875 402218 224881
rect 402166 224817 402218 224823
rect 402178 221482 402206 224817
rect 402850 221792 402878 226297
rect 402850 221764 402926 221792
rect 402898 221482 402926 221764
rect 403714 221482 403742 227555
rect 404386 226403 404414 239686
rect 404736 239672 404990 239700
rect 405216 239672 405470 239700
rect 404470 236937 404522 236943
rect 404470 236879 404522 236885
rect 404372 226394 404428 226403
rect 404372 226329 404428 226338
rect 404482 221482 404510 236879
rect 404962 226509 404990 239672
rect 405442 235135 405470 239672
rect 405428 235126 405484 235135
rect 405428 235061 405484 235070
rect 405538 234839 405566 239686
rect 405826 239672 405936 239700
rect 405826 236174 405854 239672
rect 406006 239305 406058 239311
rect 406006 239247 406058 239253
rect 405910 236937 405962 236943
rect 405910 236879 405962 236885
rect 405730 236146 405854 236174
rect 405622 235975 405674 235981
rect 405622 235917 405674 235923
rect 405634 235685 405662 235917
rect 405622 235679 405674 235685
rect 405622 235621 405674 235627
rect 405332 234830 405388 234839
rect 405332 234765 405388 234774
rect 405524 234830 405580 234839
rect 405524 234765 405580 234774
rect 405346 228507 405374 234765
rect 405334 228501 405386 228507
rect 405334 228443 405386 228449
rect 404950 226503 405002 226509
rect 404950 226445 405002 226451
rect 405730 226255 405758 236146
rect 405814 233829 405866 233835
rect 405922 233803 405950 236879
rect 406018 236055 406046 239247
rect 406306 236055 406334 239686
rect 406484 236162 406540 236171
rect 406484 236097 406540 236106
rect 406006 236049 406058 236055
rect 406006 235991 406058 235997
rect 406294 236049 406346 236055
rect 406294 235991 406346 235997
rect 406004 234682 406060 234691
rect 406004 234617 406060 234626
rect 405814 233771 405866 233777
rect 405908 233794 405964 233803
rect 405826 231879 405854 233771
rect 405908 233729 405964 233738
rect 405812 231870 405868 231879
rect 405812 231805 405868 231814
rect 406018 227712 406046 234617
rect 405922 227684 406046 227712
rect 405716 226246 405772 226255
rect 405716 226181 405772 226190
rect 405142 224949 405194 224955
rect 405142 224891 405194 224897
rect 405154 221792 405182 224891
rect 405154 221764 405230 221792
rect 405202 221482 405230 221764
rect 405922 221482 405950 227684
rect 406498 222555 406526 236097
rect 406690 234797 406718 239686
rect 407040 239672 407294 239700
rect 407424 239672 407678 239700
rect 407760 239672 408062 239700
rect 406678 234791 406730 234797
rect 406678 234733 406730 234739
rect 407266 234279 407294 239672
rect 407444 236754 407500 236763
rect 407444 236689 407500 236698
rect 407458 236319 407486 236689
rect 407444 236310 407500 236319
rect 407444 236245 407500 236254
rect 407446 234421 407498 234427
rect 407446 234363 407498 234369
rect 407254 234273 407306 234279
rect 407254 234215 407306 234221
rect 407458 233835 407486 234363
rect 407446 233829 407498 233835
rect 407446 233771 407498 233777
rect 407542 233755 407594 233761
rect 407542 233697 407594 233703
rect 406774 229685 406826 229691
rect 406774 229627 406826 229633
rect 406484 222546 406540 222555
rect 406484 222481 406540 222490
rect 406786 221482 406814 229627
rect 407554 228655 407582 233697
rect 407542 228649 407594 228655
rect 407542 228591 407594 228597
rect 407650 226107 407678 239672
rect 408034 226361 408062 239672
rect 408130 234723 408158 239686
rect 408118 234717 408170 234723
rect 408514 234691 408542 239686
rect 408960 239672 409214 239700
rect 409728 239672 409982 239700
rect 409186 235611 409214 239672
rect 409954 236171 409982 239672
rect 409940 236162 409996 236171
rect 410050 236129 410078 239686
rect 409940 236097 409996 236106
rect 410038 236123 410090 236129
rect 410038 236065 410090 236071
rect 408982 235605 409034 235611
rect 408982 235547 409034 235553
rect 409174 235605 409226 235611
rect 409174 235547 409226 235553
rect 408118 234659 408170 234665
rect 408500 234682 408556 234691
rect 408500 234617 408556 234626
rect 408994 234427 409022 235547
rect 409844 234534 409900 234543
rect 409844 234469 409900 234478
rect 408982 234421 409034 234427
rect 408982 234363 409034 234369
rect 408118 233681 408170 233687
rect 408118 233623 408170 233629
rect 408130 230399 408158 233623
rect 408886 233311 408938 233317
rect 408886 233253 408938 233259
rect 408116 230390 408172 230399
rect 408116 230325 408172 230334
rect 408214 226429 408266 226435
rect 408214 226371 408266 226377
rect 408022 226355 408074 226361
rect 408022 226297 408074 226303
rect 407636 226098 407692 226107
rect 407636 226033 407692 226042
rect 407446 225023 407498 225029
rect 407446 224965 407498 224971
rect 407458 221792 407486 224965
rect 407458 221764 407534 221792
rect 407506 221482 407534 221764
rect 408226 221482 408254 226371
rect 408898 225177 408926 233253
rect 409654 230795 409706 230801
rect 409654 230737 409706 230743
rect 408982 226133 409034 226139
rect 408982 226075 409034 226081
rect 408886 225171 408938 225177
rect 408886 225113 408938 225119
rect 408994 221482 409022 226075
rect 409666 221792 409694 230737
rect 409858 229691 409886 234469
rect 410036 234386 410092 234395
rect 410036 234321 410092 234330
rect 410050 232947 410078 234321
rect 410038 232941 410090 232947
rect 410038 232883 410090 232889
rect 409846 229685 409898 229691
rect 409846 229627 409898 229633
rect 410434 226213 410462 239686
rect 410710 236419 410762 236425
rect 410710 236361 410762 236367
rect 410722 235759 410750 236361
rect 410710 235753 410762 235759
rect 410710 235695 410762 235701
rect 410614 234421 410666 234427
rect 410818 234395 410846 239686
rect 411168 239672 411422 239700
rect 411552 239672 411710 239700
rect 411936 239672 412190 239700
rect 411394 234543 411422 239672
rect 411380 234534 411436 234543
rect 411380 234469 411436 234478
rect 410614 234363 410666 234369
rect 410804 234386 410860 234395
rect 410422 226207 410474 226213
rect 410422 226149 410474 226155
rect 410626 222587 410654 234363
rect 410804 234321 410860 234330
rect 411682 226139 411710 239672
rect 412162 235685 412190 239672
rect 420418 239237 420446 241129
rect 567380 240010 567436 240019
rect 567380 239945 567436 239954
rect 434614 239823 434666 239829
rect 434614 239765 434666 239771
rect 420406 239231 420458 239237
rect 420406 239173 420458 239179
rect 413396 238974 413452 238983
rect 413396 238909 413452 238918
rect 413410 236795 413438 238909
rect 414068 238826 414124 238835
rect 414068 238761 414124 238770
rect 413684 238678 413740 238687
rect 413602 238636 413684 238664
rect 413602 236869 413630 238636
rect 413684 238613 413740 238622
rect 413972 238382 414028 238391
rect 413698 238340 413972 238368
rect 413590 236863 413642 236869
rect 413590 236805 413642 236811
rect 413398 236789 413450 236795
rect 413398 236731 413450 236737
rect 413698 236319 413726 238340
rect 413972 238317 414028 238326
rect 414082 237480 414110 238761
rect 415220 238234 415276 238243
rect 415220 238169 415276 238178
rect 414452 238086 414508 238095
rect 414452 238021 414508 238030
rect 413794 237452 414110 237480
rect 413684 236310 413740 236319
rect 413684 236245 413740 236254
rect 413794 236148 413822 237452
rect 414466 236943 414494 238021
rect 414454 236937 414506 236943
rect 414454 236879 414506 236885
rect 415234 236319 415262 238169
rect 432406 237233 432458 237239
rect 432406 237175 432458 237181
rect 426358 237159 426410 237165
rect 426358 237101 426410 237107
rect 420310 237011 420362 237017
rect 420310 236953 420362 236959
rect 415220 236310 415276 236319
rect 415220 236245 415276 236254
rect 415412 236310 415468 236319
rect 415412 236245 415468 236254
rect 413698 236120 413822 236148
rect 413876 236162 413932 236171
rect 413698 235759 413726 236120
rect 413876 236097 413932 236106
rect 413890 235981 413918 236097
rect 415426 236055 415454 236245
rect 415414 236049 415466 236055
rect 415414 235991 415466 235997
rect 413878 235975 413930 235981
rect 413878 235917 413930 235923
rect 413686 235753 413738 235759
rect 413686 235695 413738 235701
rect 412150 235679 412202 235685
rect 412150 235621 412202 235627
rect 414742 234347 414794 234353
rect 414742 234289 414794 234295
rect 414754 231171 414782 234289
rect 414742 231165 414794 231171
rect 414742 231107 414794 231113
rect 415702 231017 415754 231023
rect 415702 230959 415754 230965
rect 413494 228575 413546 228581
rect 413494 228517 413546 228523
rect 412726 228131 412778 228137
rect 412726 228073 412778 228079
rect 411286 226133 411338 226139
rect 411286 226075 411338 226081
rect 411670 226133 411722 226139
rect 411670 226075 411722 226081
rect 410518 222581 410570 222587
rect 410518 222523 410570 222529
rect 410614 222581 410666 222587
rect 410614 222523 410666 222529
rect 409666 221764 409742 221792
rect 409714 221482 409742 221764
rect 410530 221482 410558 222523
rect 411298 221496 411326 226075
rect 411958 225319 412010 225325
rect 411958 225261 412010 225267
rect 411264 221468 411326 221496
rect 411970 221496 411998 225261
rect 411970 221468 412032 221496
rect 412738 221482 412766 228073
rect 413506 221496 413534 228517
rect 415030 225393 415082 225399
rect 415030 225335 415082 225341
rect 414262 222655 414314 222661
rect 414262 222597 414314 222603
rect 413472 221468 413534 221496
rect 414274 221482 414302 222597
rect 415042 221482 415070 225335
rect 415714 221792 415742 230959
rect 419542 230943 419594 230949
rect 419542 230885 419594 230891
rect 416470 230721 416522 230727
rect 416470 230663 416522 230669
rect 415714 221764 415790 221792
rect 415762 221482 415790 221764
rect 416482 221482 416510 230663
rect 418774 228723 418826 228729
rect 418774 228665 418826 228671
rect 418006 225245 418058 225251
rect 418006 225187 418058 225193
rect 417238 222803 417290 222809
rect 417238 222745 417290 222751
rect 417250 221482 417278 222745
rect 418018 221792 418046 225187
rect 418018 221764 418094 221792
rect 418066 221482 418094 221764
rect 418786 221482 418814 228665
rect 419158 226799 419210 226805
rect 419158 226741 419210 226747
rect 419254 226799 419306 226805
rect 419254 226741 419306 226747
rect 418870 226725 418922 226731
rect 418922 226673 419102 226676
rect 418870 226667 419102 226673
rect 418882 226648 419102 226667
rect 419074 226509 419102 226648
rect 419170 226583 419198 226741
rect 419158 226577 419210 226583
rect 419158 226519 419210 226525
rect 419062 226503 419114 226509
rect 419062 226445 419114 226451
rect 419266 225917 419294 226741
rect 419254 225911 419306 225917
rect 419254 225853 419306 225859
rect 419554 221482 419582 230885
rect 420322 221792 420350 236953
rect 426166 234495 426218 234501
rect 426166 234437 426218 234443
rect 423286 233829 423338 233835
rect 423286 233771 423338 233777
rect 421846 228797 421898 228803
rect 421846 228739 421898 228745
rect 420982 225467 421034 225473
rect 420982 225409 421034 225415
rect 420274 221764 420350 221792
rect 420274 221482 420302 221764
rect 420994 221482 421022 225409
rect 421858 221482 421886 228739
rect 423298 227619 423326 233771
rect 424054 231165 424106 231171
rect 424054 231107 424106 231113
rect 424724 231130 424780 231139
rect 423286 227613 423338 227619
rect 423286 227555 423338 227561
rect 423286 223025 423338 223031
rect 423286 222967 423338 222973
rect 422518 222877 422570 222883
rect 422518 222819 422570 222825
rect 422530 221792 422558 222819
rect 422530 221764 422606 221792
rect 422578 221482 422606 221764
rect 423298 221482 423326 222967
rect 424066 221482 424094 231107
rect 424724 231065 424780 231074
rect 424738 221792 424766 231065
rect 426178 230505 426206 234437
rect 426166 230499 426218 230505
rect 426166 230441 426218 230447
rect 425590 227983 425642 227989
rect 425590 227925 425642 227931
rect 424738 221764 424814 221792
rect 424786 221482 424814 221764
rect 425602 221482 425630 227925
rect 426370 221482 426398 237101
rect 428662 237085 428714 237091
rect 428662 237027 428714 237033
rect 427894 233903 427946 233909
rect 427894 233845 427946 233851
rect 427906 228951 427934 233845
rect 427798 228945 427850 228951
rect 427798 228887 427850 228893
rect 427894 228945 427946 228951
rect 427894 228887 427946 228893
rect 427030 225541 427082 225547
rect 427030 225483 427082 225489
rect 427042 221792 427070 225483
rect 427042 221764 427118 221792
rect 427090 221482 427118 221764
rect 427810 221482 427838 228887
rect 428674 221482 428702 237027
rect 432022 233977 432074 233983
rect 432022 233919 432074 233925
rect 432034 228877 432062 233919
rect 430870 228871 430922 228877
rect 430870 228813 430922 228819
rect 432022 228871 432074 228877
rect 432022 228813 432074 228819
rect 429334 223099 429386 223105
rect 429334 223041 429386 223047
rect 429346 221792 429374 223041
rect 430102 222581 430154 222587
rect 430102 222523 430154 222529
rect 429346 221764 429422 221792
rect 429394 221482 429422 221764
rect 430114 221482 430142 222523
rect 430882 221482 430910 228813
rect 431542 222951 431594 222957
rect 431542 222893 431594 222899
rect 431554 221792 431582 222893
rect 431554 221764 431630 221792
rect 431602 221482 431630 221764
rect 432418 221482 432446 237175
rect 433846 231535 433898 231541
rect 433846 231477 433898 231483
rect 433174 227613 433226 227619
rect 433174 227555 433226 227561
rect 433186 221482 433214 227555
rect 433858 221792 433886 231477
rect 433858 221764 433934 221792
rect 433906 221482 433934 221764
rect 434626 221482 434654 239765
rect 446710 239749 446762 239755
rect 446710 239691 446762 239697
rect 444502 237455 444554 237461
rect 444502 237397 444554 237403
rect 441430 237381 441482 237387
rect 441430 237323 441482 237329
rect 438358 237307 438410 237313
rect 438358 237249 438410 237255
rect 434902 234569 434954 234575
rect 434902 234511 434954 234517
rect 434914 229987 434942 234511
rect 436150 230499 436202 230505
rect 436150 230441 436202 230447
rect 434902 229981 434954 229987
rect 434902 229923 434954 229929
rect 435382 223173 435434 223179
rect 435382 223115 435434 223121
rect 435394 221482 435422 223115
rect 436162 221792 436190 230441
rect 436918 230425 436970 230431
rect 436918 230367 436970 230373
rect 436162 221764 436238 221792
rect 436210 221482 436238 221764
rect 436930 221482 436958 230367
rect 437686 228205 437738 228211
rect 437686 228147 437738 228153
rect 437698 221482 437726 228147
rect 438370 221792 438398 237249
rect 441442 236174 441470 237323
rect 442198 236419 442250 236425
rect 442198 236361 442250 236367
rect 440770 236146 441470 236174
rect 439990 230351 440042 230357
rect 439990 230293 440042 230299
rect 439126 225615 439178 225621
rect 439126 225557 439178 225563
rect 438370 221764 438446 221792
rect 438418 221482 438446 221764
rect 439138 221482 439166 225557
rect 440002 221496 440030 230293
rect 440770 221792 440798 236146
rect 441430 224653 441482 224659
rect 441430 224595 441482 224601
rect 439968 221468 440030 221496
rect 440722 221764 440798 221792
rect 440722 221482 440750 221764
rect 441442 221482 441470 224595
rect 442210 221496 442238 236361
rect 442868 231278 442924 231287
rect 442868 231213 442924 231222
rect 442176 221468 442238 221496
rect 442882 221496 442910 231213
rect 443734 222359 443786 222365
rect 443734 222301 443786 222307
rect 442882 221468 442944 221496
rect 443746 221482 443774 222301
rect 444514 221792 444542 237397
rect 445942 230277 445994 230283
rect 445942 230219 445994 230225
rect 445172 225358 445228 225367
rect 445172 225293 445228 225302
rect 444466 221764 444542 221792
rect 444466 221482 444494 221764
rect 445186 221482 445214 225293
rect 445954 221482 445982 230219
rect 446722 221792 446750 239691
rect 470902 239675 470954 239681
rect 470902 239617 470954 239623
rect 458806 239527 458858 239533
rect 458806 239469 458858 239475
rect 455062 239009 455114 239015
rect 455062 238951 455114 238957
rect 450454 237529 450506 237535
rect 450454 237471 450506 237477
rect 449302 234643 449354 234649
rect 449302 234585 449354 234591
rect 448246 233459 448298 233465
rect 448246 233401 448298 233407
rect 447478 224579 447530 224585
rect 447478 224521 447530 224527
rect 446674 221764 446750 221792
rect 446674 221482 446702 221764
rect 447490 221482 447518 224521
rect 448258 221482 448286 233401
rect 448916 231426 448972 231435
rect 448916 231361 448972 231370
rect 448930 221792 448958 231361
rect 449314 230209 449342 234585
rect 449686 230869 449738 230875
rect 449686 230811 449738 230817
rect 449302 230203 449354 230209
rect 449302 230145 449354 230151
rect 448930 221764 449006 221792
rect 448978 221482 449006 221764
rect 449698 221482 449726 230811
rect 450466 221482 450494 237471
rect 451990 230277 452042 230283
rect 451990 230219 452042 230225
rect 451222 225689 451274 225695
rect 451222 225631 451274 225637
rect 451234 221792 451262 225631
rect 451234 221764 451310 221792
rect 451282 221482 451310 221764
rect 452002 221482 452030 230219
rect 454294 229981 454346 229987
rect 454294 229923 454346 229929
rect 452758 224505 452810 224511
rect 452758 224447 452810 224453
rect 452770 221482 452798 224447
rect 453430 224431 453482 224437
rect 453430 224373 453482 224379
rect 453442 221792 453470 224373
rect 453442 221764 453518 221792
rect 453490 221482 453518 221764
rect 454306 221482 454334 229923
rect 455074 228729 455102 238951
rect 455158 238935 455210 238941
rect 455158 238877 455210 238883
rect 455062 228723 455114 228729
rect 455062 228665 455114 228671
rect 455170 228581 455198 238877
rect 455252 231574 455308 231583
rect 455252 231509 455308 231518
rect 455158 228575 455210 228581
rect 455158 228517 455210 228523
rect 455266 223272 455294 231509
rect 458038 230055 458090 230061
rect 458038 229997 458090 230003
rect 455734 228723 455786 228729
rect 455734 228665 455786 228671
rect 455074 223244 455294 223272
rect 455074 221482 455102 223244
rect 455746 221792 455774 228665
rect 456502 228575 456554 228581
rect 456502 228517 456554 228523
rect 455746 221764 455822 221792
rect 455794 221482 455822 221764
rect 456514 221482 456542 228517
rect 457268 225506 457324 225515
rect 457268 225441 457324 225450
rect 457282 221482 457310 225441
rect 458050 221792 458078 229997
rect 458050 221764 458126 221792
rect 458098 221482 458126 221764
rect 458818 221482 458846 239469
rect 462550 238861 462602 238867
rect 462550 238803 462602 238809
rect 460246 235901 460298 235907
rect 460246 235843 460298 235849
rect 459574 224357 459626 224363
rect 459574 224299 459626 224305
rect 459586 221482 459614 224299
rect 460258 221792 460286 235843
rect 461014 230129 461066 230135
rect 461014 230071 461066 230077
rect 460258 221764 460334 221792
rect 460306 221482 460334 221764
rect 461026 221482 461054 230071
rect 461878 228279 461930 228285
rect 461878 228221 461930 228227
rect 461890 221482 461918 228221
rect 462562 221792 462590 238803
rect 464758 238787 464810 238793
rect 464758 238729 464810 238735
rect 463606 233385 463658 233391
rect 463606 233327 463658 233333
rect 463618 230135 463646 233327
rect 464086 231609 464138 231615
rect 464086 231551 464138 231557
rect 463606 230129 463658 230135
rect 463606 230071 463658 230077
rect 463316 225654 463372 225663
rect 463316 225589 463372 225598
rect 462562 221764 462638 221792
rect 462610 221482 462638 221764
rect 463330 221482 463358 225589
rect 464098 221482 464126 231551
rect 464770 221792 464798 238729
rect 468598 238713 468650 238719
rect 468598 238655 468650 238661
rect 466486 233533 466538 233539
rect 466486 233475 466538 233481
rect 466390 230203 466442 230209
rect 466390 230145 466442 230151
rect 465622 224283 465674 224289
rect 465622 224225 465674 224231
rect 464770 221764 464846 221792
rect 464818 221482 464846 221764
rect 465634 221482 465662 224225
rect 466402 221482 466430 230145
rect 466498 230061 466526 233475
rect 466486 230055 466538 230061
rect 466486 229997 466538 230003
rect 467062 228427 467114 228433
rect 467062 228369 467114 228375
rect 467074 221792 467102 228369
rect 467830 224135 467882 224141
rect 467830 224077 467882 224083
rect 467074 221764 467150 221792
rect 467122 221482 467150 221764
rect 467842 221482 467870 224077
rect 468610 221482 468638 238655
rect 470132 231722 470188 231731
rect 470132 231657 470188 231666
rect 469364 225802 469420 225811
rect 469364 225737 469420 225746
rect 469378 221496 469406 225737
rect 469378 221468 469440 221496
rect 470146 221482 470174 231657
rect 470914 221496 470942 239617
rect 488278 239601 488330 239607
rect 488278 239543 488330 239549
rect 474646 238639 474698 238645
rect 474646 238581 474698 238587
rect 472340 234090 472396 234099
rect 472340 234025 472396 234034
rect 471574 224209 471626 224215
rect 471574 224151 471626 224157
rect 470880 221468 470942 221496
rect 471586 221496 471614 224151
rect 471586 221468 471648 221496
rect 472354 221482 472382 234025
rect 473878 231239 473930 231245
rect 473878 231181 473930 231187
rect 473110 229907 473162 229913
rect 473110 229849 473162 229855
rect 473122 221792 473150 229849
rect 473122 221764 473198 221792
rect 473170 221482 473198 221764
rect 473890 221482 473918 231181
rect 474658 221482 474686 238581
rect 480694 238565 480746 238571
rect 480694 238507 480746 238513
rect 478102 238491 478154 238497
rect 478102 238433 478154 238439
rect 475222 234051 475274 234057
rect 475222 233993 475274 233999
rect 475234 229987 475262 233993
rect 475222 229981 475274 229987
rect 475222 229923 475274 229929
rect 476950 228353 477002 228359
rect 476950 228295 477002 228301
rect 476180 228170 476236 228179
rect 476180 228105 476236 228114
rect 475316 225210 475372 225219
rect 475316 225145 475372 225154
rect 475330 221792 475358 225145
rect 475330 221764 475406 221792
rect 475378 221482 475406 221764
rect 476194 221482 476222 228105
rect 476962 221482 476990 228295
rect 477622 224061 477674 224067
rect 477622 224003 477674 224009
rect 477634 221792 477662 224003
rect 477634 221764 477710 221792
rect 478114 221773 478142 238433
rect 479158 231683 479210 231689
rect 479158 231625 479210 231631
rect 478390 230129 478442 230135
rect 478390 230071 478442 230077
rect 477682 221482 477710 221764
rect 478102 221767 478154 221773
rect 478102 221709 478154 221715
rect 478402 221482 478430 230071
rect 479170 221482 479198 231625
rect 479974 221767 480026 221773
rect 479974 221709 480026 221715
rect 479986 221482 480014 221709
rect 480706 221482 480734 238507
rect 486742 238417 486794 238423
rect 486742 238359 486794 238365
rect 484630 234125 484682 234131
rect 484630 234067 484682 234073
rect 480884 233942 480940 233951
rect 480884 233877 480940 233886
rect 480898 229913 480926 233877
rect 484438 230055 484490 230061
rect 484438 229997 484490 230003
rect 480886 229907 480938 229913
rect 480886 229849 480938 229855
rect 482134 229833 482186 229839
rect 482134 229775 482186 229781
rect 481460 227430 481516 227439
rect 481460 227365 481516 227374
rect 481474 221482 481502 227365
rect 482146 221792 482174 229775
rect 483766 223987 483818 223993
rect 483766 223929 483818 223935
rect 482902 222433 482954 222439
rect 482902 222375 482954 222381
rect 482146 221764 482222 221792
rect 482194 221482 482222 221764
rect 482914 221482 482942 222375
rect 483778 221482 483806 223929
rect 484450 221792 484478 229997
rect 484642 229839 484670 234067
rect 485206 231757 485258 231763
rect 485206 231699 485258 231705
rect 484630 229833 484682 229839
rect 484630 229775 484682 229781
rect 484450 221764 484526 221792
rect 484498 221482 484526 221764
rect 485218 221482 485246 231699
rect 485974 231313 486026 231319
rect 485974 231255 486026 231261
rect 485986 221482 486014 231255
rect 486754 221792 486782 238359
rect 488290 236174 488318 239543
rect 532822 239453 532874 239459
rect 532822 239395 532874 239401
rect 508630 239157 508682 239163
rect 508630 239099 508682 239105
rect 492790 238343 492842 238349
rect 492790 238285 492842 238291
rect 492022 236345 492074 236351
rect 492022 236287 492074 236293
rect 488290 236146 488990 236174
rect 488276 228318 488332 228327
rect 488276 228253 488332 228262
rect 487508 225950 487564 225959
rect 487508 225885 487564 225894
rect 486706 221764 486782 221792
rect 486706 221482 486734 221764
rect 487522 221482 487550 225885
rect 488290 221482 488318 228253
rect 488962 221792 488990 236146
rect 490484 234238 490540 234247
rect 490484 234173 490540 234182
rect 489718 223913 489770 223919
rect 489718 223855 489770 223861
rect 488962 221764 489038 221792
rect 489010 221482 489038 221764
rect 489730 221482 489758 223855
rect 490498 221482 490526 234173
rect 491254 233237 491306 233243
rect 491254 233179 491306 233185
rect 491266 221792 491294 233179
rect 491266 221764 491342 221792
rect 491314 221482 491342 221764
rect 492034 221482 492062 236287
rect 492802 221482 492830 238285
rect 500278 238269 500330 238275
rect 500278 238211 500330 238217
rect 495766 235827 495818 235833
rect 495766 235769 495818 235775
rect 495382 234199 495434 234205
rect 495382 234141 495434 234147
rect 495394 233243 495422 234141
rect 495382 233237 495434 233243
rect 495092 233202 495148 233211
rect 495382 233179 495434 233185
rect 495092 233137 495148 233146
rect 494228 228614 494284 228623
rect 494228 228549 494284 228558
rect 493460 227282 493516 227291
rect 493460 227217 493516 227226
rect 493474 221792 493502 227217
rect 493474 221764 493550 221792
rect 493522 221482 493550 221764
rect 494242 221482 494270 228549
rect 495106 221482 495134 233137
rect 495778 221792 495806 235769
rect 499606 231387 499658 231393
rect 499606 231329 499658 231335
rect 497972 228466 498028 228475
rect 497972 228401 498028 228410
rect 497302 223839 497354 223845
rect 497302 223781 497354 223787
rect 496534 222507 496586 222513
rect 496534 222449 496586 222455
rect 495778 221764 495854 221792
rect 495826 221482 495854 221764
rect 496546 221482 496574 222449
rect 497314 221482 497342 223781
rect 497986 221792 498014 228401
rect 498836 227134 498892 227143
rect 498836 227069 498892 227078
rect 497986 221764 498062 221792
rect 498034 221482 498062 221764
rect 498850 221482 498878 227069
rect 499618 221496 499646 231329
rect 499584 221468 499646 221496
rect 500290 221496 500318 238211
rect 503350 238195 503402 238201
rect 503350 238137 503402 238143
rect 501046 233163 501098 233169
rect 501046 233105 501098 233111
rect 500290 221468 500352 221496
rect 501058 221482 501086 233105
rect 502582 228501 502634 228507
rect 502582 228443 502634 228449
rect 501814 223765 501866 223771
rect 501814 223707 501866 223713
rect 501826 221792 501854 223707
rect 501826 221764 501902 221792
rect 501874 221482 501902 221764
rect 502594 221482 502622 228443
rect 503362 221482 503390 238137
rect 505654 236271 505706 236277
rect 505654 236213 505706 236219
rect 503926 234273 503978 234279
rect 503926 234215 503978 234221
rect 503938 230061 503966 234215
rect 503926 230055 503978 230061
rect 503926 229997 503978 230003
rect 504022 229759 504074 229765
rect 504022 229701 504074 229707
rect 504034 221792 504062 229701
rect 504790 223617 504842 223623
rect 504790 223559 504842 223565
rect 504034 221764 504110 221792
rect 504082 221482 504110 221764
rect 504802 221482 504830 223559
rect 505666 221482 505694 236213
rect 507094 233089 507146 233095
rect 507094 233031 507146 233037
rect 506326 223543 506378 223549
rect 506326 223485 506378 223491
rect 506338 221792 506366 223485
rect 506338 221764 506414 221792
rect 506386 221482 506414 221764
rect 507106 221482 507134 233031
rect 507862 223691 507914 223697
rect 507862 223633 507914 223639
rect 507874 221482 507902 223633
rect 508642 221792 508670 239099
rect 509398 238121 509450 238127
rect 509398 238063 509450 238069
rect 508594 221764 508670 221792
rect 508594 221482 508622 221764
rect 509410 221482 509438 238063
rect 514678 238047 514730 238053
rect 514678 237989 514730 237995
rect 512758 237973 512810 237979
rect 512758 237915 512810 237921
rect 510166 229611 510218 229617
rect 510166 229553 510218 229559
rect 510178 221482 510206 229553
rect 510838 223469 510890 223475
rect 510838 223411 510890 223417
rect 510850 221792 510878 223411
rect 512374 223321 512426 223327
rect 512374 223263 512426 223269
rect 511606 222729 511658 222735
rect 511606 222671 511658 222677
rect 510850 221764 510926 221792
rect 510898 221482 510926 221764
rect 511618 221482 511646 222671
rect 512386 221482 512414 223263
rect 512770 221773 512798 237915
rect 513142 233015 513194 233021
rect 513142 232957 513194 232963
rect 513154 221792 513182 232957
rect 513910 223395 513962 223401
rect 513910 223337 513962 223343
rect 512758 221767 512810 221773
rect 513154 221764 513230 221792
rect 512758 221709 512810 221715
rect 513202 221482 513230 221764
rect 513922 221482 513950 223337
rect 514690 221482 514718 237989
rect 522166 237899 522218 237905
rect 522166 237841 522218 237847
rect 522178 236174 522206 237841
rect 521506 236146 522206 236174
rect 523798 236197 523850 236203
rect 519190 232867 519242 232873
rect 519190 232809 519242 232815
rect 516118 229537 516170 229543
rect 516118 229479 516170 229485
rect 515398 221767 515450 221773
rect 515398 221709 515450 221715
rect 515410 221482 515438 221709
rect 516130 221482 516158 229479
rect 517654 228649 517706 228655
rect 517654 228591 517706 228597
rect 516982 223247 517034 223253
rect 516982 223189 517034 223195
rect 516994 221482 517022 223189
rect 517666 221792 517694 228591
rect 518420 222990 518476 222999
rect 518420 222925 518476 222934
rect 517666 221764 517742 221792
rect 517714 221482 517742 221764
rect 518434 221482 518462 222925
rect 519202 221482 519230 232809
rect 520726 231461 520778 231467
rect 520726 231403 520778 231409
rect 519860 222694 519916 222703
rect 519860 222629 519916 222638
rect 519874 221792 519902 222629
rect 519874 221764 519950 221792
rect 519922 221482 519950 221764
rect 520738 221482 520766 231403
rect 521506 221482 521534 236146
rect 523798 236139 523850 236145
rect 522166 229389 522218 229395
rect 522166 229331 522218 229337
rect 522178 221792 522206 229331
rect 522932 222546 522988 222555
rect 522932 222481 522988 222490
rect 522178 221764 522254 221792
rect 522226 221482 522254 221764
rect 522946 221482 522974 222481
rect 523810 221482 523838 236139
rect 525238 232793 525290 232799
rect 525238 232735 525290 232741
rect 524468 222842 524524 222851
rect 524468 222777 524524 222786
rect 524482 221792 524510 222777
rect 524482 221764 524558 221792
rect 524530 221482 524558 221764
rect 525250 221482 525278 232735
rect 531286 232645 531338 232651
rect 531286 232587 531338 232593
rect 527540 230094 527596 230103
rect 527540 230029 527596 230038
rect 526004 224618 526060 224627
rect 526004 224553 526060 224562
rect 526018 221482 526046 224553
rect 526676 224470 526732 224479
rect 526676 224405 526732 224414
rect 526690 221792 526718 224405
rect 526690 221764 526766 221792
rect 526738 221482 526766 221764
rect 527554 221482 527582 230029
rect 529750 228871 529802 228877
rect 529750 228813 529802 228819
rect 528308 228762 528364 228771
rect 528308 228697 528364 228706
rect 528322 221496 528350 228697
rect 528980 224322 529036 224331
rect 528980 224257 529036 224266
rect 528288 221468 528350 221496
rect 528994 221496 529022 224257
rect 528994 221468 529056 221496
rect 529762 221482 529790 228813
rect 530516 224174 530572 224183
rect 530516 224109 530572 224118
rect 530530 221496 530558 224109
rect 530496 221468 530558 221496
rect 531298 221482 531326 232587
rect 532052 224026 532108 224035
rect 532052 223961 532108 223970
rect 532066 221482 532094 223961
rect 532834 221792 532862 239395
rect 541462 239379 541514 239385
rect 541462 239321 541514 239327
rect 538004 238086 538060 238095
rect 538004 238021 538060 238030
rect 535126 237825 535178 237831
rect 535126 237767 535178 237773
rect 533494 237751 533546 237757
rect 533494 237693 533546 237699
rect 532786 221764 532862 221792
rect 532786 221482 532814 221764
rect 533506 221482 533534 237693
rect 534260 230242 534316 230251
rect 534260 230177 534316 230186
rect 534274 221482 534302 230177
rect 535138 221792 535166 237767
rect 535798 237677 535850 237683
rect 535798 237619 535850 237625
rect 535810 228581 535838 237619
rect 538018 236174 538046 238021
rect 541078 237603 541130 237609
rect 541078 237545 541130 237551
rect 537922 236146 538046 236174
rect 537238 232571 537290 232577
rect 537238 232513 537290 232519
rect 535798 228575 535850 228581
rect 535798 228517 535850 228523
rect 535798 228427 535850 228433
rect 535798 228369 535850 228375
rect 535090 221764 535166 221792
rect 535090 221482 535118 221764
rect 535810 221482 535838 228369
rect 536564 223878 536620 223887
rect 536564 223813 536620 223822
rect 536578 221482 536606 223813
rect 537250 221792 537278 232513
rect 537922 228433 537950 236146
rect 539542 232423 539594 232429
rect 539542 232365 539594 232371
rect 538870 229463 538922 229469
rect 538870 229405 538922 229411
rect 538006 228575 538058 228581
rect 538006 228517 538058 228523
rect 537910 228427 537962 228433
rect 537910 228369 537962 228375
rect 537250 221764 537326 221792
rect 537298 221482 537326 221764
rect 538018 221482 538046 228517
rect 538882 221482 538910 229405
rect 539554 221792 539582 232365
rect 540308 229946 540364 229955
rect 540308 229881 540364 229890
rect 539554 221764 539630 221792
rect 539602 221482 539630 221764
rect 540322 221482 540350 229881
rect 541090 221482 541118 237545
rect 541474 236174 541502 239321
rect 550870 239305 550922 239311
rect 550870 239247 550922 239253
rect 544822 239083 544874 239089
rect 544822 239025 544874 239031
rect 544340 238382 544396 238391
rect 544340 238317 544396 238326
rect 541474 236146 541790 236174
rect 541762 221792 541790 236146
rect 542614 232497 542666 232503
rect 542614 232439 542666 232445
rect 541762 221764 541838 221792
rect 541810 221482 541838 221764
rect 542626 221482 542654 232439
rect 543382 232349 543434 232355
rect 543382 232291 543434 232297
rect 543394 221482 543422 232291
rect 544354 228581 544382 238317
rect 544342 228575 544394 228581
rect 544342 228517 544394 228523
rect 544052 223730 544108 223739
rect 544052 223665 544108 223674
rect 544066 221792 544094 223665
rect 544066 221764 544142 221792
rect 544114 221482 544142 221764
rect 544834 221482 544862 239025
rect 550196 238678 550252 238687
rect 550196 238613 550252 238622
rect 549428 233054 549484 233063
rect 549428 232989 549484 232998
rect 548566 232275 548618 232281
rect 548566 232217 548618 232223
rect 545590 232201 545642 232207
rect 545590 232143 545642 232149
rect 545602 221482 545630 232143
rect 546358 229315 546410 229321
rect 546358 229257 546410 229263
rect 546370 221792 546398 229257
rect 547894 228945 547946 228951
rect 547894 228887 547946 228893
rect 547126 228575 547178 228581
rect 547126 228517 547178 228523
rect 546370 221764 546446 221792
rect 546418 221482 546446 221764
rect 547138 221482 547166 228517
rect 547906 221482 547934 228887
rect 548578 221792 548606 232217
rect 548578 221764 548654 221792
rect 548626 221482 548654 221764
rect 549442 221482 549470 232989
rect 550210 221482 550238 238613
rect 550882 221792 550910 239247
rect 555380 238974 555436 238983
rect 555380 238909 555436 238918
rect 551636 232906 551692 232915
rect 551636 232841 551692 232850
rect 550882 221764 550958 221792
rect 550930 221482 550958 221764
rect 551650 221482 551678 232841
rect 552406 232127 552458 232133
rect 552406 232069 552458 232075
rect 552418 221482 552446 232069
rect 554710 232053 554762 232059
rect 554710 231995 554762 232001
rect 553940 229798 553996 229807
rect 553940 229733 553996 229742
rect 553270 224209 553322 224215
rect 553270 224151 553322 224157
rect 553282 221792 553310 224151
rect 553234 221764 553310 221792
rect 553234 221482 553262 221764
rect 553954 221482 553982 229733
rect 554722 221482 554750 231995
rect 555286 229241 555338 229247
rect 555286 229183 555338 229189
rect 555298 221792 555326 229183
rect 555394 224215 555422 238909
rect 559892 238234 559948 238243
rect 559892 238169 559948 238178
rect 559220 236606 559276 236615
rect 559220 236541 559276 236550
rect 557684 236458 557740 236467
rect 557684 236393 557740 236402
rect 557588 232758 557644 232767
rect 557588 232693 557644 232702
rect 557014 231905 557066 231911
rect 557014 231847 557066 231853
rect 556150 228575 556202 228581
rect 556150 228517 556202 228523
rect 555382 224209 555434 224215
rect 555382 224151 555434 224157
rect 555298 221764 555470 221792
rect 555442 221482 555470 221764
rect 556162 221482 556190 228517
rect 557026 221496 557054 231847
rect 557602 227534 557630 232693
rect 557698 228581 557726 236393
rect 558454 231979 558506 231985
rect 558454 231921 558506 231927
rect 557686 228575 557738 228581
rect 557686 228517 557738 228523
rect 557602 227506 557726 227534
rect 556992 221468 557054 221496
rect 557698 221496 557726 227506
rect 557698 221468 557760 221496
rect 558466 221482 558494 231921
rect 559234 221496 559262 236541
rect 559200 221468 559262 221496
rect 559906 221496 559934 238169
rect 565268 236754 565324 236763
rect 565268 236689 565324 236698
rect 560756 232610 560812 232619
rect 560756 232545 560812 232554
rect 559906 221468 559968 221496
rect 560770 221482 560798 232545
rect 564502 231831 564554 231837
rect 564502 231773 564554 231779
rect 561430 229167 561482 229173
rect 561430 229109 561482 229115
rect 561442 221792 561470 229109
rect 563638 229093 563690 229099
rect 563638 229035 563690 229041
rect 562964 223582 563020 223591
rect 562964 223517 563020 223526
rect 562196 223434 562252 223443
rect 562196 223369 562252 223378
rect 561442 221764 561518 221792
rect 561490 221482 561518 221764
rect 562210 221482 562238 223369
rect 562978 221482 563006 223517
rect 563650 221792 563678 229035
rect 563650 221764 563726 221792
rect 563698 221482 563726 221764
rect 564514 221482 564542 231773
rect 565282 221482 565310 236689
rect 566710 232719 566762 232725
rect 566710 232661 566762 232667
rect 565942 229685 565994 229691
rect 565942 229627 565994 229633
rect 565954 221792 565982 229627
rect 565954 221764 566030 221792
rect 566002 221482 566030 221764
rect 566722 221482 566750 232661
rect 567394 228581 567422 239945
rect 599158 239231 599210 239237
rect 599158 239173 599210 239179
rect 581780 238826 581836 238835
rect 581780 238761 581836 238770
rect 573140 237050 573196 237059
rect 573140 236985 573196 236994
rect 567476 236902 567532 236911
rect 567476 236837 567532 236846
rect 567490 236174 567518 236837
rect 573154 236174 573182 236985
rect 567490 236146 568286 236174
rect 573154 236146 574334 236174
rect 567478 229019 567530 229025
rect 567478 228961 567530 228967
rect 567382 228575 567434 228581
rect 567382 228517 567434 228523
rect 567490 221482 567518 228961
rect 568258 221792 568286 236146
rect 572086 232941 572138 232947
rect 572086 232883 572138 232889
rect 570452 232462 570508 232471
rect 570452 232397 570508 232406
rect 569780 229650 569836 229659
rect 569780 229585 569836 229594
rect 569014 228575 569066 228581
rect 569014 228517 569066 228523
rect 568258 221764 568334 221792
rect 568306 221482 568334 221764
rect 569026 221482 569054 228517
rect 569794 221482 569822 229585
rect 570466 221792 570494 232397
rect 571316 223286 571372 223295
rect 571316 223221 571372 223230
rect 570466 221764 570542 221792
rect 570514 221482 570542 221764
rect 571330 221482 571358 223221
rect 572098 221482 572126 232883
rect 572756 229502 572812 229511
rect 572756 229437 572812 229446
rect 572770 221792 572798 229437
rect 573524 229354 573580 229363
rect 573524 229289 573580 229298
rect 572770 221764 572846 221792
rect 572818 221482 572846 221764
rect 573538 221482 573566 229289
rect 574306 221482 574334 236146
rect 580340 236014 580396 236023
rect 580340 235949 580396 235958
rect 576596 232314 576652 232323
rect 576596 232249 576652 232258
rect 575828 232018 575884 232027
rect 575828 231953 575884 231962
rect 575060 230390 575116 230399
rect 575060 230325 575116 230334
rect 575074 221792 575102 230325
rect 575074 221764 575150 221792
rect 575122 221482 575150 221764
rect 575842 221482 575870 231953
rect 576610 221482 576638 232249
rect 578036 232166 578092 232175
rect 578036 232101 578092 232110
rect 577268 223138 577324 223147
rect 577268 223073 577324 223082
rect 577282 221792 577310 223073
rect 577282 221764 577358 221792
rect 577330 221482 577358 221764
rect 578050 221482 578078 232101
rect 578900 229206 578956 229215
rect 578900 229141 578956 229150
rect 578914 221482 578942 229141
rect 579574 226059 579626 226065
rect 579574 226001 579626 226007
rect 579586 221792 579614 226001
rect 579586 221764 579662 221792
rect 579634 221482 579662 221764
rect 580354 221482 580382 235949
rect 581110 225837 581162 225843
rect 581110 225779 581162 225785
rect 581122 221482 581150 225779
rect 581794 221792 581822 238761
rect 591476 236162 591532 236171
rect 584566 236123 584618 236129
rect 591476 236097 591532 236106
rect 584566 236065 584618 236071
rect 583414 235161 583466 235167
rect 583414 235103 583466 235109
rect 582646 225985 582698 225991
rect 582646 225927 582698 225933
rect 581794 221764 581870 221792
rect 581842 221482 581870 221764
rect 582658 221482 582686 225927
rect 583426 221482 583454 235103
rect 584578 226065 584606 236065
rect 587924 235866 587980 235875
rect 587924 235801 587980 235810
rect 587350 235531 587402 235537
rect 587350 235473 587402 235479
rect 587062 235383 587114 235389
rect 587062 235325 587114 235331
rect 585526 235309 585578 235315
rect 585526 235251 585578 235257
rect 584854 227243 584906 227249
rect 584854 227185 584906 227191
rect 584566 226059 584618 226065
rect 584566 226001 584618 226007
rect 584086 225763 584138 225769
rect 584086 225705 584138 225711
rect 584098 221792 584126 225705
rect 584098 221764 584174 221792
rect 584146 221482 584174 221764
rect 584866 221482 584894 227185
rect 585538 225547 585566 235251
rect 585622 227391 585674 227397
rect 585622 227333 585674 227339
rect 585526 225541 585578 225547
rect 585526 225483 585578 225489
rect 585634 221482 585662 227333
rect 586390 227317 586442 227323
rect 586390 227259 586442 227265
rect 586402 221496 586430 227259
rect 587074 225769 587102 235325
rect 587158 227539 587210 227545
rect 587158 227481 587210 227487
rect 587062 225763 587114 225769
rect 587062 225705 587114 225711
rect 586402 221468 586464 221496
rect 587170 221482 587198 227481
rect 587362 226953 587390 235473
rect 587638 235457 587690 235463
rect 587638 235399 587690 235405
rect 587444 234386 587500 234395
rect 587444 234321 587500 234330
rect 587458 227249 587486 234321
rect 587446 227243 587498 227249
rect 587446 227185 587498 227191
rect 587350 226947 587402 226953
rect 587350 226889 587402 226895
rect 587650 226731 587678 235399
rect 587638 226725 587690 226731
rect 587638 226667 587690 226673
rect 587938 221496 587966 235801
rect 590708 235718 590764 235727
rect 590422 235679 590474 235685
rect 590708 235653 590764 235662
rect 590422 235621 590474 235627
rect 588790 235605 588842 235611
rect 588790 235547 588842 235553
rect 588598 235235 588650 235241
rect 588598 235177 588650 235183
rect 588610 227471 588638 235177
rect 588598 227465 588650 227471
rect 588598 227407 588650 227413
rect 588802 227323 588830 235547
rect 589366 227391 589418 227397
rect 589366 227333 589418 227339
rect 588790 227317 588842 227323
rect 588790 227259 588842 227265
rect 588598 227169 588650 227175
rect 588598 227111 588650 227117
rect 587904 221468 587966 221496
rect 588610 221496 588638 227111
rect 588610 221468 588672 221496
rect 589378 221482 589406 227333
rect 590434 227101 590462 235621
rect 590722 227545 590750 235653
rect 590900 234534 590956 234543
rect 590900 234469 590956 234478
rect 590710 227539 590762 227545
rect 590710 227481 590762 227487
rect 590914 227175 590942 234469
rect 590902 227169 590954 227175
rect 590902 227111 590954 227117
rect 590134 227095 590186 227101
rect 590134 227037 590186 227043
rect 590422 227095 590474 227101
rect 590422 227037 590474 227043
rect 590146 221792 590174 227037
rect 590900 226838 590956 226847
rect 590900 226773 590956 226782
rect 590146 221764 590222 221792
rect 590194 221482 590222 221764
rect 590914 221482 590942 226773
rect 591490 225843 591518 236097
rect 596086 235087 596138 235093
rect 596086 235029 596138 235035
rect 594646 227539 594698 227545
rect 594646 227481 594698 227487
rect 593974 227021 594026 227027
rect 591668 226986 591724 226995
rect 593974 226963 594026 226969
rect 591668 226921 591724 226930
rect 591478 225837 591530 225843
rect 591478 225779 591530 225785
rect 591682 221482 591710 226921
rect 592342 225541 592394 225547
rect 592342 225483 592394 225489
rect 592354 221792 592382 225483
rect 593110 224727 593162 224733
rect 593110 224669 593162 224675
rect 592354 221764 592430 221792
rect 592402 221482 592430 221764
rect 593122 221482 593150 224669
rect 593986 221482 594014 226963
rect 594658 221792 594686 227481
rect 595414 225763 595466 225769
rect 595414 225705 595466 225711
rect 594658 221764 594734 221792
rect 594706 221482 594734 221764
rect 595426 221482 595454 225705
rect 596098 224733 596126 235029
rect 599170 227027 599198 239173
rect 599924 229058 599980 229067
rect 599924 228993 599980 229002
rect 599158 227021 599210 227027
rect 599158 226963 599210 226969
rect 598486 226947 598538 226953
rect 598486 226889 598538 226895
rect 596180 226690 596236 226699
rect 596180 226625 596236 226634
rect 596086 224727 596138 224733
rect 596086 224669 596138 224675
rect 596194 221482 596222 226625
rect 596948 226542 597004 226551
rect 596948 226477 597004 226486
rect 596962 221792 596990 226477
rect 597718 224727 597770 224733
rect 597718 224669 597770 224675
rect 596962 221764 597038 221792
rect 597010 221482 597038 221764
rect 597730 221482 597758 224669
rect 598498 221482 598526 226889
rect 599158 226873 599210 226879
rect 599158 226815 599210 226821
rect 599170 221792 599198 226815
rect 599170 221764 599246 221792
rect 599218 221482 599246 221764
rect 599938 221482 599966 228993
rect 600418 226879 600446 241911
rect 601462 229981 601514 229987
rect 601462 229923 601514 229929
rect 600790 227465 600842 227471
rect 600790 227407 600842 227413
rect 600406 226873 600458 226879
rect 600406 226815 600458 226821
rect 600802 221482 600830 227407
rect 601474 221792 601502 229923
rect 603298 226805 603326 253455
rect 603382 250627 603434 250633
rect 603382 250569 603434 250575
rect 603394 227027 603422 250569
rect 603478 247815 603530 247821
rect 603478 247757 603530 247763
rect 603382 227021 603434 227027
rect 603382 226963 603434 226969
rect 603286 226799 603338 226805
rect 603286 226741 603338 226747
rect 602230 226725 602282 226731
rect 602230 226667 602282 226673
rect 601474 221764 601550 221792
rect 601522 221482 601550 221764
rect 602242 221482 602270 226667
rect 602998 226651 603050 226657
rect 602998 226593 603050 226599
rect 603010 221482 603038 226593
rect 603490 225991 603518 247757
rect 605974 235013 606026 235019
rect 605974 234955 606026 234961
rect 605302 234939 605354 234945
rect 605302 234881 605354 234887
rect 604532 231870 604588 231879
rect 604532 231805 604588 231814
rect 603670 226725 603722 226731
rect 603670 226667 603722 226673
rect 603478 225985 603530 225991
rect 603478 225927 603530 225933
rect 603682 221792 603710 226667
rect 603682 221764 603758 221792
rect 603730 221482 603758 221764
rect 604546 221482 604574 231805
rect 605314 221482 605342 234881
rect 605986 221792 606014 234955
rect 606178 226657 606206 262113
rect 606262 259285 606314 259291
rect 606262 259227 606314 259233
rect 606274 226731 606302 259227
rect 606358 256399 606410 256405
rect 606358 256341 606410 256347
rect 606370 227471 606398 256341
rect 629206 247741 629258 247747
rect 629206 247683 629258 247689
rect 627188 240158 627244 240167
rect 627188 240093 627244 240102
rect 621140 236310 621196 236319
rect 621140 236245 621196 236254
rect 608276 235570 608332 235579
rect 608276 235505 608332 235514
rect 607508 228910 607564 228919
rect 607508 228845 607564 228854
rect 606358 227465 606410 227471
rect 606358 227407 606410 227413
rect 606262 226725 606314 226731
rect 606262 226667 606314 226673
rect 606166 226651 606218 226657
rect 606166 226593 606218 226599
rect 606742 225097 606794 225103
rect 606742 225039 606794 225045
rect 605986 221764 606062 221792
rect 606034 221482 606062 221764
rect 606754 221482 606782 225039
rect 607522 221482 607550 228845
rect 608290 221792 608318 235505
rect 611252 235422 611308 235431
rect 611252 235357 611308 235366
rect 609046 229907 609098 229913
rect 609046 229849 609098 229855
rect 608290 221764 608366 221792
rect 608338 221482 608366 221764
rect 609058 221482 609086 229849
rect 609814 226577 609866 226583
rect 609814 226519 609866 226525
rect 609826 221482 609854 226519
rect 610486 225171 610538 225177
rect 610486 225113 610538 225119
rect 610498 221792 610526 225113
rect 610498 221764 610574 221792
rect 610546 221482 610574 221764
rect 611266 221482 611294 235357
rect 614324 235274 614380 235283
rect 614324 235209 614380 235218
rect 612118 229833 612170 229839
rect 612118 229775 612170 229781
rect 612130 221482 612158 229775
rect 612790 226503 612842 226509
rect 612790 226445 612842 226451
rect 612802 221792 612830 226445
rect 613558 226429 613610 226435
rect 613558 226371 613610 226377
rect 612802 221764 612878 221792
rect 612850 221482 612878 221764
rect 613570 221482 613598 226371
rect 614338 221482 614366 235209
rect 618836 235126 618892 235135
rect 618836 235061 618892 235070
rect 616628 234978 616684 234987
rect 616628 234913 616684 234922
rect 615862 234865 615914 234871
rect 615862 234807 615914 234813
rect 614998 233237 615050 233243
rect 614998 233179 615050 233185
rect 615010 221792 615038 233179
rect 615010 221764 615086 221792
rect 615058 221482 615086 221764
rect 615874 221482 615902 234807
rect 616642 221496 616670 234913
rect 617300 226394 617356 226403
rect 617300 226329 617356 226338
rect 618070 226355 618122 226361
rect 616608 221468 616670 221496
rect 617314 221496 617342 226329
rect 618070 226297 618122 226303
rect 617314 221468 617376 221496
rect 618082 221482 618110 226297
rect 618850 221792 618878 235061
rect 619604 234830 619660 234839
rect 619604 234765 619660 234774
rect 618850 221764 618926 221792
rect 618898 221482 618926 221764
rect 619618 221482 619646 234765
rect 620372 226246 620428 226255
rect 620372 226181 620428 226190
rect 620386 221482 620414 226181
rect 621154 221792 621182 236245
rect 621814 234791 621866 234797
rect 621814 234733 621866 234739
rect 621106 221764 621182 221792
rect 621106 221482 621134 221764
rect 621826 221482 621854 234733
rect 624886 234717 624938 234723
rect 624886 234659 624938 234665
rect 625556 234682 625612 234691
rect 622678 230055 622730 230061
rect 622678 229997 622730 230003
rect 622690 221482 622718 229997
rect 624118 226281 624170 226287
rect 624118 226223 624170 226229
rect 623348 226098 623404 226107
rect 623348 226033 623404 226042
rect 623362 221792 623390 226033
rect 623362 221764 623438 221792
rect 623410 221482 623438 221764
rect 624130 221482 624158 226223
rect 624898 221482 624926 234659
rect 625556 234617 625612 234626
rect 625570 221792 625598 234617
rect 626422 227317 626474 227323
rect 626422 227259 626474 227265
rect 625570 221764 625646 221792
rect 625618 221482 625646 221764
rect 626434 221482 626462 227259
rect 627202 221482 627230 240093
rect 629218 226435 629246 247683
rect 629302 244855 629354 244861
rect 629302 244797 629354 244803
rect 629314 227545 629342 244797
rect 629302 227539 629354 227545
rect 629302 227481 629354 227487
rect 634006 227539 634058 227545
rect 634006 227481 634058 227487
rect 630166 227243 630218 227249
rect 630166 227185 630218 227191
rect 629206 226429 629258 226435
rect 629206 226371 629258 226377
rect 629398 226207 629450 226213
rect 629398 226149 629450 226155
rect 628630 226059 628682 226065
rect 628630 226001 628682 226007
rect 627862 225763 627914 225769
rect 627862 225705 627914 225711
rect 627874 221792 627902 225705
rect 627874 221764 627950 221792
rect 627922 221482 627950 221764
rect 628642 221482 628670 226001
rect 629410 221482 629438 226149
rect 630178 221792 630206 227185
rect 630934 227169 630986 227175
rect 630934 227111 630986 227117
rect 630178 221764 630254 221792
rect 630226 221482 630254 221764
rect 630946 221482 630974 227111
rect 632374 227095 632426 227101
rect 632374 227037 632426 227043
rect 631702 226133 631754 226139
rect 631702 226075 631754 226081
rect 631714 221482 631742 226075
rect 632386 221792 632414 227037
rect 633142 226947 633194 226953
rect 633142 226889 633194 226895
rect 632386 221764 632462 221792
rect 632434 221482 632462 221764
rect 633154 221482 633182 226889
rect 634018 221482 634046 227481
rect 638518 227465 638570 227471
rect 638518 227407 638570 227413
rect 636886 227021 636938 227027
rect 636886 226963 636938 226969
rect 634678 226873 634730 226879
rect 634678 226815 634730 226821
rect 634690 221792 634718 226815
rect 635446 226429 635498 226435
rect 635446 226371 635498 226377
rect 634690 221764 634766 221792
rect 634738 221482 634766 221764
rect 635458 221482 635486 226371
rect 636214 225985 636266 225991
rect 636214 225927 636266 225933
rect 636226 221482 636254 225927
rect 636898 221792 636926 226963
rect 637750 226799 637802 226805
rect 637750 226741 637802 226747
rect 636898 221764 636974 221792
rect 636946 221482 636974 221764
rect 637762 221482 637790 226741
rect 638530 221482 638558 227407
rect 639190 226725 639242 226731
rect 639190 226667 639242 226673
rect 639202 221792 639230 226667
rect 639958 226651 640010 226657
rect 639958 226593 640010 226599
rect 639202 221764 639278 221792
rect 639250 221482 639278 221764
rect 639970 221482 639998 226593
rect 640148 212334 640204 212343
rect 640148 212269 640204 212278
rect 640162 211603 640190 212269
rect 640148 211594 640204 211603
rect 640148 211529 640204 211538
rect 190292 201382 190348 201391
rect 190292 201317 190348 201326
rect 190306 200577 190334 201317
rect 640148 200938 640204 200947
rect 640148 200873 640204 200882
rect 190292 200568 190348 200577
rect 190292 200503 190348 200512
rect 640162 200207 640190 200873
rect 640148 200198 640204 200207
rect 640148 200133 640204 200142
rect 187220 199162 187276 199171
rect 187220 199097 187276 199106
rect 640244 185694 640300 185703
rect 640244 185629 640300 185638
rect 640258 184963 640286 185629
rect 640244 184954 640300 184963
rect 640244 184889 640300 184898
rect 645142 183139 645194 183145
rect 645142 183081 645194 183087
rect 645154 183039 645182 183081
rect 645140 183030 645196 183039
rect 645140 182965 645196 182974
rect 186260 182438 186316 182447
rect 186260 182373 186316 182382
rect 645142 179439 645194 179445
rect 645142 179381 645194 179387
rect 645154 179339 645182 179381
rect 645140 179330 645196 179339
rect 645140 179265 645196 179274
rect 645142 174925 645194 174931
rect 645140 174890 645142 174899
rect 645194 174890 645196 174899
rect 645140 174825 645196 174834
rect 645142 171077 645194 171083
rect 645140 171042 645142 171051
rect 645194 171042 645196 171051
rect 645140 170977 645196 170986
rect 645142 168265 645194 168271
rect 645142 168207 645194 168213
rect 645154 167795 645182 168207
rect 645140 167786 645196 167795
rect 645140 167721 645196 167730
rect 645142 163381 645194 163387
rect 645140 163346 645142 163355
rect 645194 163346 645196 163355
rect 645140 163281 645196 163290
rect 645142 159755 645194 159761
rect 645142 159697 645194 159703
rect 645154 159507 645182 159697
rect 645140 159498 645196 159507
rect 645140 159433 645196 159442
rect 645142 156055 645194 156061
rect 645142 155997 645194 156003
rect 645154 155511 645182 155997
rect 645140 155502 645196 155511
rect 645140 155437 645196 155446
rect 645142 152577 645194 152583
rect 645140 152542 645142 152551
rect 645194 152542 645196 152551
rect 645140 152477 645196 152486
rect 645142 148211 645194 148217
rect 645142 148153 645194 148159
rect 645154 148111 645182 148153
rect 645140 148102 645196 148111
rect 645140 148037 645196 148046
rect 186742 146879 186794 146885
rect 186742 146821 186794 146827
rect 186754 145891 186782 146821
rect 186740 145882 186796 145891
rect 186740 145817 186796 145826
rect 186164 137446 186220 137455
rect 186164 137381 186220 137390
rect 186082 135346 186302 135374
rect 186274 135235 186302 135346
rect 186260 135226 186316 135235
rect 186260 135161 186316 135170
rect 646498 123945 646526 275465
rect 646594 126757 646622 277241
rect 647362 269323 647390 278018
rect 648610 272135 648638 278018
rect 648596 272126 648652 272135
rect 648596 272061 648652 272070
rect 647348 269314 647404 269323
rect 647348 269249 647404 269258
rect 646678 249147 646730 249153
rect 646678 249089 646730 249095
rect 646690 144263 646718 249089
rect 646774 207559 646826 207565
rect 646774 207501 646826 207507
rect 646676 144254 646732 144263
rect 646676 144189 646732 144198
rect 646786 141007 646814 207501
rect 649378 183145 649406 861106
rect 655220 778286 655276 778295
rect 655220 778221 655276 778230
rect 654164 774882 654220 774891
rect 654164 774817 654220 774826
rect 654178 774775 654206 774817
rect 654166 774769 654218 774775
rect 654166 774711 654218 774717
rect 654836 772366 654892 772375
rect 654836 772301 654892 772310
rect 654850 771963 654878 772301
rect 654838 771957 654890 771963
rect 654838 771899 654890 771905
rect 655124 734478 655180 734487
rect 655124 734413 655180 734422
rect 654164 730334 654220 730343
rect 654164 730269 654220 730278
rect 654178 728747 654206 730269
rect 654260 729150 654316 729159
rect 654260 729085 654316 729094
rect 654166 728741 654218 728747
rect 654166 728683 654218 728689
rect 654164 727966 654220 727975
rect 654164 727901 654220 727910
rect 654178 724381 654206 727901
rect 654274 727193 654302 729085
rect 654262 727187 654314 727193
rect 654262 727129 654314 727135
rect 654166 724375 654218 724381
rect 654166 724317 654218 724323
rect 649462 688411 649514 688417
rect 649462 688353 649514 688359
rect 649366 183139 649418 183145
rect 649366 183081 649418 183087
rect 649474 179445 649502 688353
rect 654452 683566 654508 683575
rect 654452 683501 654508 683510
rect 654466 681165 654494 683501
rect 654454 681159 654506 681165
rect 654454 681101 654506 681107
rect 655138 656893 655166 734413
rect 655234 702921 655262 778221
rect 655604 777694 655660 777703
rect 655604 777629 655660 777638
rect 655412 775918 655468 775927
rect 655412 775853 655468 775862
rect 655316 731666 655372 731675
rect 655316 731601 655372 731610
rect 655222 702915 655274 702921
rect 655222 702857 655274 702863
rect 655220 689486 655276 689495
rect 655220 689421 655276 689430
rect 655126 656887 655178 656893
rect 655126 656829 655178 656835
rect 652246 655333 652298 655339
rect 652246 655275 652298 655281
rect 649750 655259 649802 655265
rect 649750 655201 649802 655207
rect 649558 645195 649610 645201
rect 649558 645137 649610 645143
rect 649462 179439 649514 179445
rect 649462 179381 649514 179387
rect 649570 174931 649598 645137
rect 649654 601979 649706 601985
rect 649654 601921 649706 601927
rect 649558 174925 649610 174931
rect 649558 174867 649610 174873
rect 649666 171083 649694 601921
rect 649762 263403 649790 655201
rect 649846 555877 649898 555883
rect 649846 555819 649898 555825
rect 649748 263394 649804 263403
rect 649748 263329 649804 263338
rect 649654 171077 649706 171083
rect 649654 171019 649706 171025
rect 649858 168271 649886 555819
rect 649942 512735 649994 512741
rect 649942 512677 649994 512683
rect 649846 168265 649898 168271
rect 649846 168207 649898 168213
rect 649954 163387 649982 512677
rect 650038 469519 650090 469525
rect 650038 469461 650090 469467
rect 649942 163381 649994 163387
rect 649942 163323 649994 163329
rect 646870 161531 646922 161537
rect 646870 161473 646922 161479
rect 646772 140998 646828 141007
rect 646772 140933 646828 140942
rect 646582 126751 646634 126757
rect 646582 126693 646634 126699
rect 646486 123939 646538 123945
rect 646486 123881 646538 123887
rect 646498 122063 646526 123881
rect 646594 123839 646622 126693
rect 646882 125763 646910 161473
rect 647062 161457 647114 161463
rect 647062 161399 647114 161405
rect 646966 161383 647018 161389
rect 646966 161325 647018 161331
rect 646978 127687 647006 161325
rect 647074 134791 647102 161399
rect 650050 159761 650078 469461
rect 650134 383087 650186 383093
rect 650134 383029 650186 383035
rect 650038 159755 650090 159761
rect 650038 159697 650090 159703
rect 650146 156061 650174 383029
rect 650230 337059 650282 337065
rect 650230 337001 650282 337007
rect 650134 156055 650186 156061
rect 650134 155997 650186 156003
rect 650242 152583 650270 337001
rect 650422 334173 650474 334179
rect 650422 334115 650474 334121
rect 650326 291697 650378 291703
rect 650326 291639 650378 291645
rect 650230 152577 650282 152583
rect 650230 152519 650282 152525
rect 650338 148217 650366 291639
rect 650434 275687 650462 334115
rect 650420 275678 650476 275687
rect 650420 275613 650476 275622
rect 652258 266395 652286 655275
rect 655124 643014 655180 643023
rect 655124 642949 655180 642958
rect 654166 642235 654218 642241
rect 654166 642177 654218 642183
rect 654178 640655 654206 642177
rect 654164 640646 654220 640655
rect 654164 640581 654220 640590
rect 654550 602053 654602 602059
rect 654550 601995 654602 602001
rect 654562 595367 654590 601995
rect 654548 595358 654604 595367
rect 654548 595293 654604 595302
rect 654164 593434 654220 593443
rect 654164 593369 654166 593378
rect 654218 593369 654220 593378
rect 654166 593337 654218 593343
rect 654356 591954 654412 591963
rect 654356 591889 654412 591898
rect 654370 590515 654398 591889
rect 654358 590509 654410 590515
rect 654358 590451 654410 590457
rect 655138 567427 655166 642949
rect 655234 613677 655262 689421
rect 655330 657041 655358 731601
rect 655426 699887 655454 775853
rect 655508 732702 655564 732711
rect 655508 732637 655564 732646
rect 655414 699881 655466 699887
rect 655414 699823 655466 699829
rect 655412 688450 655468 688459
rect 655412 688385 655468 688394
rect 655318 657035 655370 657041
rect 655318 656977 655370 656983
rect 655316 642422 655372 642431
rect 655316 642357 655372 642366
rect 655222 613671 655274 613677
rect 655222 613613 655274 613619
rect 655220 597874 655276 597883
rect 655220 597809 655276 597818
rect 655126 567421 655178 567427
rect 655126 567363 655178 567369
rect 655124 553326 655180 553335
rect 655124 553261 655180 553270
rect 653782 552917 653834 552923
rect 653782 552859 653834 552865
rect 653794 550967 653822 552859
rect 653780 550958 653836 550967
rect 653780 550893 653836 550902
rect 654164 547554 654220 547563
rect 654164 547489 654220 547498
rect 654178 547447 654206 547489
rect 654166 547441 654218 547447
rect 654166 547383 654218 547389
rect 655138 480995 655166 553261
rect 655234 524211 655262 597809
rect 655330 567797 655358 642357
rect 655426 613825 655454 688385
rect 655522 657189 655550 732637
rect 655618 703069 655646 777629
rect 656180 773550 656236 773559
rect 656180 773485 656236 773494
rect 656194 771889 656222 773485
rect 656182 771883 656234 771889
rect 656182 771825 656234 771831
rect 655606 703063 655658 703069
rect 655606 703005 655658 703011
rect 670882 700849 670910 877201
rect 670966 876223 671018 876229
rect 670966 876165 671018 876171
rect 669526 700843 669578 700849
rect 669526 700785 669578 700791
rect 670870 700843 670922 700849
rect 670870 700785 670922 700791
rect 655604 687118 655660 687127
rect 655604 687053 655660 687062
rect 655510 657183 655562 657189
rect 655510 657125 655562 657131
rect 655508 640794 655564 640803
rect 655508 640729 655564 640738
rect 655414 613819 655466 613825
rect 655414 613761 655466 613767
rect 655412 596690 655468 596699
rect 655412 596625 655468 596634
rect 655318 567791 655370 567797
rect 655318 567733 655370 567739
rect 655316 552142 655372 552151
rect 655316 552077 655372 552086
rect 655222 524205 655274 524211
rect 655222 524147 655274 524153
rect 655330 481217 655358 552077
rect 655426 524433 655454 596625
rect 655522 567945 655550 640729
rect 655618 613973 655646 687053
rect 656372 685934 656428 685943
rect 656372 685869 656428 685878
rect 656386 685605 656414 685869
rect 656374 685599 656426 685605
rect 656374 685541 656426 685547
rect 655988 684750 656044 684759
rect 655988 684685 656044 684694
rect 656002 681239 656030 684685
rect 655990 681233 656042 681239
rect 655990 681175 656042 681181
rect 655796 638278 655852 638287
rect 655796 638213 655852 638222
rect 655810 636691 655838 638213
rect 655892 637094 655948 637103
rect 655892 637029 655948 637038
rect 655798 636685 655850 636691
rect 655798 636627 655850 636633
rect 655906 635063 655934 637029
rect 655894 635057 655946 635063
rect 655894 634999 655946 635005
rect 655606 613967 655658 613973
rect 655606 613909 655658 613915
rect 655604 595506 655660 595515
rect 655604 595441 655660 595450
rect 655510 567939 655562 567945
rect 655510 567881 655562 567887
rect 655508 551106 655564 551115
rect 655508 551041 655564 551050
rect 655414 524427 655466 524433
rect 655414 524369 655466 524375
rect 655522 481365 655550 551041
rect 655618 524581 655646 595441
rect 656276 548590 656332 548599
rect 656276 548525 656332 548534
rect 656290 547373 656318 548525
rect 656278 547367 656330 547373
rect 656278 547309 656330 547315
rect 655606 524575 655658 524581
rect 655606 524517 655658 524523
rect 655510 481359 655562 481365
rect 655510 481301 655562 481307
rect 655318 481211 655370 481217
rect 655318 481153 655370 481159
rect 655126 480989 655178 480995
rect 655126 480931 655178 480937
rect 655510 394779 655562 394785
rect 655510 394721 655562 394727
rect 655318 394705 655370 394711
rect 655318 394647 655370 394653
rect 655126 394631 655178 394637
rect 655126 394573 655178 394579
rect 655138 374403 655166 394573
rect 655124 374394 655180 374403
rect 655124 374329 655180 374338
rect 655330 372183 655358 394647
rect 655522 373367 655550 394721
rect 666646 383013 666698 383019
rect 666646 382955 666698 382961
rect 655508 373358 655564 373367
rect 655508 373293 655564 373302
rect 655316 372174 655372 372183
rect 655316 372109 655372 372118
rect 654166 371543 654218 371549
rect 654166 371485 654218 371491
rect 654178 370999 654206 371485
rect 654164 370990 654220 370999
rect 654164 370925 654220 370934
rect 666658 360893 666686 382955
rect 660310 360887 660362 360893
rect 660310 360829 660362 360835
rect 666646 360887 666698 360893
rect 666646 360829 666698 360835
rect 655222 351637 655274 351643
rect 655222 351579 655274 351585
rect 655126 351563 655178 351569
rect 655126 351505 655178 351511
rect 654166 328327 654218 328333
rect 654166 328269 654218 328275
rect 654178 326303 654206 328269
rect 655138 328079 655166 351505
rect 655234 329855 655262 351579
rect 660322 351421 660350 360829
rect 655414 351415 655466 351421
rect 655414 351357 655466 351363
rect 660310 351415 660362 351421
rect 660310 351357 660362 351363
rect 655318 348529 655370 348535
rect 655318 348471 655370 348477
rect 655220 329846 655276 329855
rect 655220 329781 655276 329790
rect 655124 328070 655180 328079
rect 655124 328005 655180 328014
rect 655330 327487 655358 348471
rect 655426 334179 655454 351357
rect 655414 334173 655466 334179
rect 655414 334115 655466 334121
rect 655316 327478 655372 327487
rect 655316 327413 655372 327422
rect 654164 326294 654220 326303
rect 654164 326229 654220 326238
rect 654070 305313 654122 305319
rect 654070 305255 654122 305261
rect 653782 305239 653834 305245
rect 653782 305181 653834 305187
rect 653794 303363 653822 305181
rect 653780 303354 653836 303363
rect 653780 303289 653836 303298
rect 654082 302179 654110 305255
rect 654166 302353 654218 302359
rect 654166 302295 654218 302301
rect 654068 302170 654124 302179
rect 654068 302105 654124 302114
rect 654178 300995 654206 302295
rect 654164 300986 654220 300995
rect 654164 300921 654220 300930
rect 656564 298766 656620 298775
rect 656564 298701 656620 298710
rect 656372 297582 656428 297591
rect 656372 297517 656428 297526
rect 656180 296842 656236 296851
rect 656180 296777 656236 296786
rect 656084 295214 656140 295223
rect 656084 295149 656140 295158
rect 655892 294030 655948 294039
rect 655892 293965 655948 293974
rect 655796 292846 655852 292855
rect 655796 292781 655852 292790
rect 655604 290922 655660 290931
rect 655604 290857 655660 290866
rect 654164 289294 654220 289303
rect 654164 289229 654220 289238
rect 654178 289187 654206 289229
rect 654166 289181 654218 289187
rect 654166 289123 654218 289129
rect 655412 288110 655468 288119
rect 655412 288045 655468 288054
rect 653780 284558 653836 284567
rect 653780 284493 653836 284502
rect 653794 284303 653822 284493
rect 653782 284297 653834 284303
rect 653782 284239 653834 284245
rect 655124 283374 655180 283383
rect 655124 283309 655180 283318
rect 654740 279822 654796 279831
rect 654740 279757 654796 279766
rect 654754 279419 654782 279757
rect 654742 279413 654794 279419
rect 654742 279355 654794 279361
rect 652246 266389 652298 266395
rect 652246 266331 652298 266337
rect 650326 148211 650378 148217
rect 650326 148153 650378 148159
rect 647060 134782 647116 134791
rect 647060 134717 647116 134726
rect 647732 130934 647788 130943
rect 647732 130869 647788 130878
rect 646964 127678 647020 127687
rect 646964 127613 647020 127622
rect 646868 125754 646924 125763
rect 646868 125689 646924 125698
rect 646580 123830 646636 123839
rect 646580 123765 646636 123774
rect 646484 122054 646540 122063
rect 646484 121989 646540 121998
rect 186262 120683 186314 120689
rect 186262 120625 186314 120631
rect 185684 110214 185740 110223
rect 185684 110149 185740 110158
rect 185302 109361 185354 109367
rect 185300 109326 185302 109335
rect 185354 109326 185356 109335
rect 185300 109261 185356 109270
rect 186274 108743 186302 120625
rect 646198 118463 646250 118469
rect 646198 118405 646250 118411
rect 646210 117623 646238 118405
rect 646196 117614 646252 117623
rect 646196 117549 646252 117558
rect 647746 115509 647774 130869
rect 647924 129010 647980 129019
rect 647924 128945 647980 128954
rect 647938 126831 647966 128945
rect 655138 126979 655166 283309
rect 655316 282338 655372 282347
rect 655316 282273 655372 282282
rect 655220 281006 655276 281015
rect 655220 280941 655276 280950
rect 655234 127127 655262 280941
rect 655330 129643 655358 282273
rect 655426 172859 655454 288045
rect 655508 286926 655564 286935
rect 655508 286861 655564 286870
rect 655522 173081 655550 286861
rect 655618 219109 655646 290857
rect 655700 285742 655756 285751
rect 655700 285677 655756 285686
rect 655606 219103 655658 219109
rect 655606 219045 655658 219051
rect 655714 173229 655742 285677
rect 655810 219257 655838 292781
rect 655906 241901 655934 293965
rect 655988 291662 656044 291671
rect 655988 291597 656044 291606
rect 655894 241895 655946 241901
rect 655894 241837 655946 241843
rect 656002 219405 656030 291597
rect 656098 259513 656126 295149
rect 656194 262325 656222 296777
rect 656386 262473 656414 297517
rect 656578 288003 656606 298701
rect 660886 289181 660938 289187
rect 660886 289123 660938 289129
rect 656566 287997 656618 288003
rect 656566 287939 656618 287945
rect 658006 284297 658058 284303
rect 658006 284239 658058 284245
rect 656374 262467 656426 262473
rect 656374 262409 656426 262415
rect 656182 262319 656234 262325
rect 656182 262261 656234 262267
rect 656086 259507 656138 259513
rect 656086 259449 656138 259455
rect 655990 219399 656042 219405
rect 655990 219341 656042 219347
rect 655798 219251 655850 219257
rect 655798 219193 655850 219199
rect 655702 173223 655754 173229
rect 655702 173165 655754 173171
rect 655510 173075 655562 173081
rect 655510 173017 655562 173023
rect 655414 172853 655466 172859
rect 655414 172795 655466 172801
rect 658018 155543 658046 284239
rect 660898 198685 660926 289123
rect 663766 279413 663818 279419
rect 663766 279355 663818 279361
rect 660886 198679 660938 198685
rect 660886 198621 660938 198627
rect 658006 155537 658058 155543
rect 658006 155479 658058 155485
rect 655318 129637 655370 129643
rect 655318 129579 655370 129585
rect 655222 127121 655274 127127
rect 655222 127063 655274 127069
rect 655126 126973 655178 126979
rect 655126 126915 655178 126921
rect 647926 126825 647978 126831
rect 647926 126767 647978 126773
rect 647828 119538 647884 119547
rect 647828 119473 647884 119482
rect 647734 115503 647786 115509
rect 647734 115445 647786 115451
rect 647842 115361 647870 119473
rect 647924 115690 647980 115699
rect 647924 115625 647980 115634
rect 647830 115355 647882 115361
rect 647830 115297 647882 115303
rect 647938 115287 647966 115625
rect 647926 115281 647978 115287
rect 647926 115223 647978 115229
rect 663778 114695 663806 279355
rect 668180 277898 668236 277907
rect 668180 277833 668236 277842
rect 665302 115281 665354 115287
rect 665302 115223 665354 115229
rect 663766 114689 663818 114695
rect 663766 114631 663818 114637
rect 646580 113174 646636 113183
rect 646580 113109 646636 113118
rect 186260 108734 186316 108743
rect 186260 108669 186316 108678
rect 186646 106549 186698 106555
rect 186646 106491 186698 106497
rect 186658 106375 186686 106491
rect 186644 106366 186700 106375
rect 186644 106301 186700 106310
rect 645908 106070 645964 106079
rect 645908 106005 645964 106014
rect 645922 103891 645950 106005
rect 645910 103885 645962 103891
rect 645910 103827 645962 103833
rect 184724 102518 184780 102527
rect 184724 102453 184780 102462
rect 645140 102222 645196 102231
rect 645140 102157 645196 102166
rect 645154 102115 645182 102157
rect 645142 102109 645194 102115
rect 645142 102051 645194 102057
rect 184628 98078 184684 98087
rect 184246 98039 184298 98045
rect 184628 98013 184684 98022
rect 184246 97981 184298 97987
rect 180118 94635 180170 94641
rect 180118 94577 180170 94583
rect 184258 81955 184286 97981
rect 186166 97965 186218 97971
rect 186166 97907 186218 97913
rect 184342 97891 184394 97897
rect 184342 97833 184394 97839
rect 184354 97199 184382 97833
rect 184438 97817 184490 97823
rect 184438 97759 184490 97765
rect 184340 97190 184396 97199
rect 184340 97125 184396 97134
rect 184450 96459 184478 97759
rect 184534 97743 184586 97749
rect 184534 97685 184586 97691
rect 184436 96450 184492 96459
rect 184436 96385 184492 96394
rect 184546 95719 184574 97685
rect 184532 95710 184588 95719
rect 184532 95645 184588 95654
rect 184534 95005 184586 95011
rect 184534 94947 184586 94953
rect 184438 94931 184490 94937
rect 184438 94873 184490 94879
rect 184342 94857 184394 94863
rect 184340 94822 184342 94831
rect 184394 94822 184396 94831
rect 184340 94757 184396 94766
rect 184450 93499 184478 94873
rect 184436 93490 184492 93499
rect 184436 93425 184492 93434
rect 184546 92759 184574 94947
rect 184630 94635 184682 94641
rect 184630 94577 184682 94583
rect 184642 94239 184670 94577
rect 184628 94230 184684 94239
rect 184628 94165 184684 94174
rect 184532 92750 184588 92759
rect 184532 92685 184588 92694
rect 184534 92119 184586 92125
rect 184534 92061 184586 92067
rect 184438 92045 184490 92051
rect 184340 92010 184396 92019
rect 184438 91987 184490 91993
rect 184340 91945 184342 91954
rect 184394 91945 184396 91954
rect 184342 91913 184394 91919
rect 184450 90391 184478 91987
rect 184436 90382 184492 90391
rect 184436 90317 184492 90326
rect 184546 89651 184574 92061
rect 184630 91897 184682 91903
rect 184630 91839 184682 91845
rect 184642 91131 184670 91839
rect 184628 91122 184684 91131
rect 184628 91057 184684 91066
rect 184532 89642 184588 89651
rect 184532 89577 184588 89586
rect 184630 89233 184682 89239
rect 184630 89175 184682 89181
rect 184534 89159 184586 89165
rect 184534 89101 184586 89107
rect 184438 89085 184490 89091
rect 184438 89027 184490 89033
rect 184342 89011 184394 89017
rect 184342 88953 184394 88959
rect 184354 88911 184382 88953
rect 184340 88902 184396 88911
rect 184340 88837 184396 88846
rect 184450 88171 184478 89027
rect 184436 88162 184492 88171
rect 184436 88097 184492 88106
rect 184546 87283 184574 89101
rect 184532 87274 184588 87283
rect 184532 87209 184588 87218
rect 184642 86691 184670 89175
rect 184628 86682 184684 86691
rect 184628 86617 184684 86626
rect 184534 86421 184586 86427
rect 184534 86363 184586 86369
rect 184342 86347 184394 86353
rect 184342 86289 184394 86295
rect 184354 85803 184382 86289
rect 184438 86273 184490 86279
rect 184438 86215 184490 86221
rect 184340 85794 184396 85803
rect 184340 85729 184396 85738
rect 184450 84323 184478 86215
rect 184546 85211 184574 86363
rect 184532 85202 184588 85211
rect 184532 85137 184588 85146
rect 184436 84314 184492 84323
rect 184436 84249 184492 84258
rect 184438 83535 184490 83541
rect 184438 83477 184490 83483
rect 184342 83461 184394 83467
rect 184340 83426 184342 83435
rect 184394 83426 184396 83435
rect 184340 83361 184396 83370
rect 184244 81946 184300 81955
rect 184244 81881 184300 81890
rect 184450 81363 184478 83477
rect 186178 82843 186206 97907
rect 640726 96559 640778 96565
rect 640726 96501 640778 96507
rect 186164 82834 186220 82843
rect 186164 82769 186220 82778
rect 184436 81354 184492 81363
rect 184436 81289 184492 81298
rect 184438 80649 184490 80655
rect 184438 80591 184490 80597
rect 184342 80501 184394 80507
rect 184342 80443 184394 80449
rect 179926 80427 179978 80433
rect 179926 80369 179978 80375
rect 184354 78995 184382 80443
rect 184450 79883 184478 80591
rect 184534 80575 184586 80581
rect 184534 80517 184586 80523
rect 184436 79874 184492 79883
rect 184436 79809 184492 79818
rect 184340 78986 184396 78995
rect 184340 78921 184396 78930
rect 184546 78255 184574 80517
rect 184628 80466 184684 80475
rect 184628 80401 184630 80410
rect 184682 80401 184684 80410
rect 184630 80369 184682 80375
rect 184532 78246 184588 78255
rect 184532 78181 184588 78190
rect 184438 77763 184490 77769
rect 184438 77705 184490 77711
rect 184342 77615 184394 77621
rect 184342 77557 184394 77563
rect 156406 77541 156458 77547
rect 156406 77483 156458 77489
rect 184354 76775 184382 77557
rect 184450 77515 184478 77705
rect 184630 77689 184682 77695
rect 184630 77631 184682 77637
rect 184534 77541 184586 77547
rect 184436 77506 184492 77515
rect 184534 77483 184586 77489
rect 184436 77441 184492 77450
rect 184340 76766 184396 76775
rect 184340 76701 184396 76710
rect 184546 75147 184574 77483
rect 184642 76035 184670 77631
rect 184628 76026 184684 76035
rect 184628 75961 184684 75970
rect 184532 75138 184588 75147
rect 184532 75073 184588 75082
rect 184534 74877 184586 74883
rect 184534 74819 184586 74825
rect 184438 74729 184490 74735
rect 184438 74671 184490 74677
rect 154102 74655 154154 74661
rect 154102 74597 154154 74603
rect 184342 74655 184394 74661
rect 184342 74597 184394 74603
rect 184354 74407 184382 74597
rect 184340 74398 184396 74407
rect 184340 74333 184396 74342
rect 184450 72927 184478 74671
rect 184546 73667 184574 74819
rect 184630 74803 184682 74809
rect 184630 74745 184682 74751
rect 184532 73658 184588 73667
rect 184532 73593 184588 73602
rect 184436 72918 184492 72927
rect 184436 72853 184492 72862
rect 184642 72187 184670 74745
rect 184628 72178 184684 72187
rect 184628 72113 184684 72122
rect 184342 71991 184394 71997
rect 184342 71933 184394 71939
rect 149686 71843 149738 71849
rect 149686 71785 149738 71791
rect 184354 71447 184382 71933
rect 184438 71917 184490 71923
rect 184438 71859 184490 71865
rect 184340 71438 184396 71447
rect 184340 71373 184396 71382
rect 149506 70952 149630 70980
rect 149492 70846 149548 70855
rect 149492 70781 149548 70790
rect 149396 69514 149452 69523
rect 149396 69449 149452 69458
rect 149302 68957 149354 68963
rect 149302 68899 149354 68905
rect 149206 68883 149258 68889
rect 149206 68825 149258 68831
rect 149204 68330 149260 68339
rect 149204 68265 149260 68274
rect 149110 66219 149162 66225
rect 149110 66161 149162 66167
rect 149014 65997 149066 66003
rect 149014 65939 149066 65945
rect 149218 63117 149246 68265
rect 149410 66077 149438 69449
rect 149506 66151 149534 70781
rect 149602 69037 149630 70952
rect 184450 70559 184478 71859
rect 184534 71843 184586 71849
rect 184534 71785 184586 71791
rect 184436 70550 184492 70559
rect 184436 70485 184492 70494
rect 184546 69967 184574 71785
rect 184532 69958 184588 69967
rect 184532 69893 184588 69902
rect 184342 69105 184394 69111
rect 184340 69070 184342 69079
rect 184394 69070 184396 69079
rect 149590 69031 149642 69037
rect 184340 69005 184396 69014
rect 184438 69031 184490 69037
rect 149590 68973 149642 68979
rect 184438 68973 184490 68979
rect 184342 68883 184394 68889
rect 184342 68825 184394 68831
rect 184354 67599 184382 68825
rect 184450 68487 184478 68973
rect 184534 68957 184586 68963
rect 184534 68899 184586 68905
rect 184436 68478 184492 68487
rect 184436 68413 184492 68422
rect 184340 67590 184396 67599
rect 184340 67525 184396 67534
rect 149588 67146 149644 67155
rect 149588 67081 149644 67090
rect 149494 66145 149546 66151
rect 149494 66087 149546 66093
rect 149398 66071 149450 66077
rect 149398 66013 149450 66019
rect 149492 65370 149548 65379
rect 149492 65305 149548 65314
rect 149396 64630 149452 64639
rect 149396 64565 149452 64574
rect 149300 63446 149356 63455
rect 149300 63381 149356 63390
rect 149206 63111 149258 63117
rect 149206 63053 149258 63059
rect 149314 60379 149342 63381
rect 149410 63191 149438 64565
rect 149506 63265 149534 65305
rect 149602 63339 149630 67081
rect 184546 66859 184574 68899
rect 184532 66850 184588 66859
rect 184532 66785 184588 66794
rect 184534 66219 184586 66225
rect 184534 66161 184586 66167
rect 184340 66110 184396 66119
rect 184340 66045 184396 66054
rect 184438 66071 184490 66077
rect 184354 66003 184382 66045
rect 184438 66013 184490 66019
rect 184342 65997 184394 66003
rect 184342 65939 184394 65945
rect 184450 63751 184478 66013
rect 184546 65231 184574 66161
rect 184630 66145 184682 66151
rect 184630 66087 184682 66093
rect 184532 65222 184588 65231
rect 184532 65157 184588 65166
rect 184642 64639 184670 66087
rect 184628 64630 184684 64639
rect 184628 64565 184684 64574
rect 184436 63742 184492 63751
rect 184436 63677 184492 63686
rect 149590 63333 149642 63339
rect 149590 63275 149642 63281
rect 184438 63333 184490 63339
rect 184438 63275 184490 63281
rect 149494 63259 149546 63265
rect 149494 63201 149546 63207
rect 149398 63185 149450 63191
rect 149398 63127 149450 63133
rect 184340 63150 184396 63159
rect 184340 63085 184342 63094
rect 184394 63085 184396 63094
rect 184342 63053 184394 63059
rect 184450 62271 184478 63275
rect 184534 63259 184586 63265
rect 184534 63201 184586 63207
rect 149492 62262 149548 62271
rect 149492 62197 149548 62206
rect 184436 62262 184492 62271
rect 184436 62197 184492 62206
rect 149396 60634 149452 60643
rect 149396 60569 149452 60578
rect 149410 60453 149438 60569
rect 149398 60447 149450 60453
rect 149398 60389 149450 60395
rect 149302 60373 149354 60379
rect 149302 60315 149354 60321
rect 149506 60305 149534 62197
rect 184546 61531 184574 63201
rect 184630 63185 184682 63191
rect 184630 63127 184682 63133
rect 184532 61522 184588 61531
rect 184532 61457 184588 61466
rect 184642 60791 184670 63127
rect 184628 60782 184684 60791
rect 184628 60717 184684 60726
rect 184534 60447 184586 60453
rect 184534 60389 184586 60395
rect 184342 60373 184394 60379
rect 184342 60315 184394 60321
rect 149494 60299 149546 60305
rect 149494 60241 149546 60247
rect 184354 60051 184382 60315
rect 184438 60299 184490 60305
rect 184438 60241 184490 60247
rect 184340 60042 184396 60051
rect 184340 59977 184396 59986
rect 149396 59746 149452 59755
rect 149396 59681 149452 59690
rect 149410 59047 149438 59681
rect 184450 59311 184478 60241
rect 184436 59302 184492 59311
rect 184436 59237 184492 59246
rect 149398 59041 149450 59047
rect 149398 58983 149450 58989
rect 184342 59041 184394 59047
rect 184342 58983 184394 58989
rect 149396 58562 149452 58571
rect 149396 58497 149452 58506
rect 149410 57567 149438 58497
rect 184354 57683 184382 58983
rect 184546 58423 184574 60389
rect 184532 58414 184588 58423
rect 184532 58349 184588 58358
rect 184340 57674 184396 57683
rect 184340 57609 184396 57618
rect 149398 57561 149450 57567
rect 149398 57503 149450 57509
rect 184342 57561 184394 57567
rect 184342 57503 184394 57509
rect 149492 57378 149548 57387
rect 149492 57313 149548 57322
rect 149398 56229 149450 56235
rect 149396 56194 149398 56203
rect 149450 56194 149452 56203
rect 149506 56161 149534 57313
rect 184354 56943 184382 57503
rect 184340 56934 184396 56943
rect 184340 56869 184396 56878
rect 184438 56229 184490 56235
rect 184340 56194 184396 56203
rect 149396 56129 149452 56138
rect 149494 56155 149546 56161
rect 184438 56171 184490 56177
rect 184340 56129 184342 56138
rect 149494 56097 149546 56103
rect 184394 56129 184396 56138
rect 184342 56097 184394 56103
rect 184450 55463 184478 56171
rect 184436 55454 184492 55463
rect 184436 55389 184492 55398
rect 149684 54862 149740 54871
rect 149684 54797 149740 54806
rect 149698 54681 149726 54797
rect 184340 54714 184396 54723
rect 149686 54675 149738 54681
rect 184340 54649 184342 54658
rect 149686 54617 149738 54623
rect 184394 54649 184396 54658
rect 184342 54617 184394 54623
rect 184340 53974 184396 53983
rect 184340 53909 184396 53918
rect 149396 53826 149452 53835
rect 149396 53761 149452 53770
rect 149410 53275 149438 53761
rect 184354 53275 184382 53909
rect 149398 53269 149450 53275
rect 149398 53211 149450 53217
rect 184342 53269 184394 53275
rect 184342 53211 184394 53217
rect 145104 49788 145406 49816
rect 145378 47133 145406 49788
rect 199138 47133 199166 53650
rect 145366 47127 145418 47133
rect 145366 47069 145418 47075
rect 199126 47127 199178 47133
rect 199126 47069 199178 47075
rect 142114 46680 142416 46708
rect 142114 40219 142142 46680
rect 216418 46245 216446 53650
rect 233698 47725 233726 53650
rect 233686 47719 233738 47725
rect 233686 47661 233738 47667
rect 250978 47577 251006 53650
rect 268320 53636 268574 53664
rect 285600 53636 285854 53664
rect 268546 47651 268574 53636
rect 268534 47645 268586 47651
rect 268534 47587 268586 47593
rect 250966 47571 251018 47577
rect 250966 47513 251018 47519
rect 207382 46239 207434 46245
rect 207382 46181 207434 46187
rect 216406 46239 216458 46245
rect 216406 46181 216458 46187
rect 186262 42021 186314 42027
rect 186262 41963 186314 41969
rect 187030 42021 187082 42027
rect 194326 42021 194378 42027
rect 187082 41969 187344 41972
rect 187030 41963 187344 41969
rect 186274 41509 186302 41963
rect 187042 41944 187344 41963
rect 194064 41969 194326 41972
rect 194064 41963 194378 41969
rect 194064 41944 194366 41963
rect 207394 41509 207422 46181
rect 285826 43285 285854 53636
rect 302914 47873 302942 53650
rect 305302 48015 305354 48021
rect 305302 47957 305354 47963
rect 302902 47867 302954 47873
rect 302902 47809 302954 47815
rect 285814 43279 285866 43285
rect 285814 43221 285866 43227
rect 305314 43211 305342 47957
rect 311062 47941 311114 47947
rect 311062 47883 311114 47889
rect 302902 43205 302954 43211
rect 302902 43147 302954 43153
rect 305302 43205 305354 43211
rect 305302 43147 305354 43153
rect 302914 42120 302942 43147
rect 311074 42268 311102 47883
rect 320194 47799 320222 53650
rect 320182 47793 320234 47799
rect 320182 47735 320234 47741
rect 337474 46763 337502 53650
rect 354850 48021 354878 53650
rect 371938 53636 372192 53664
rect 389218 53636 389472 53664
rect 354838 48015 354890 48021
rect 354838 47957 354890 47963
rect 371938 47947 371966 53636
rect 371926 47941 371978 47947
rect 371926 47883 371978 47889
rect 328342 46757 328394 46763
rect 328342 46699 328394 46705
rect 337462 46757 337514 46763
rect 337462 46699 337514 46705
rect 310498 42240 311102 42268
rect 310498 42120 310526 42240
rect 302688 42092 302942 42120
rect 307008 42101 307262 42120
rect 307008 42095 307274 42101
rect 307008 42092 307222 42095
rect 310128 42092 310526 42120
rect 311062 42095 311114 42101
rect 307222 42037 307274 42043
rect 311062 42037 311114 42043
rect 186262 41503 186314 41509
rect 186262 41445 186314 41451
rect 207382 41503 207434 41509
rect 207382 41445 207434 41451
rect 142100 40210 142156 40219
rect 142100 40145 142156 40154
rect 311074 37259 311102 42037
rect 328354 37259 328382 46699
rect 365314 42240 365726 42268
rect 357718 42169 357770 42175
rect 357456 42117 357718 42120
rect 365314 42120 365342 42240
rect 357456 42111 357770 42117
rect 357456 42092 357758 42111
rect 361776 42101 362078 42120
rect 361776 42095 362090 42101
rect 361776 42092 362038 42095
rect 364944 42092 365342 42120
rect 362038 42037 362090 42043
rect 365698 41824 365726 42240
rect 365974 42095 366026 42101
rect 365974 42037 366026 42043
rect 365698 41796 365918 41824
rect 365890 37439 365918 41796
rect 365878 37433 365930 37439
rect 365878 37375 365930 37381
rect 365986 37365 366014 42037
rect 389218 37365 389246 53636
rect 405526 47941 405578 47947
rect 405526 47883 405578 47889
rect 401782 46165 401834 46171
rect 401782 46107 401834 46113
rect 401794 42101 401822 46107
rect 403222 43205 403274 43211
rect 403222 43147 403274 43153
rect 401782 42095 401834 42101
rect 401782 42037 401834 42043
rect 403234 37513 403262 43147
rect 405538 42106 405566 47883
rect 406786 46171 406814 53650
rect 424066 48465 424094 53650
rect 418774 48459 418826 48465
rect 418774 48401 418826 48407
rect 424054 48459 424106 48465
rect 424054 48401 424106 48407
rect 406774 46165 406826 46171
rect 406774 46107 406826 46113
rect 418786 43211 418814 48401
rect 426166 48015 426218 48021
rect 426166 47957 426218 47963
rect 426178 44955 426206 47957
rect 441346 47947 441374 53650
rect 441334 47941 441386 47947
rect 441334 47883 441386 47889
rect 426164 44946 426220 44955
rect 426164 44881 426220 44890
rect 458626 43211 458654 53650
rect 475714 53636 475968 53664
rect 492994 53636 493248 53664
rect 510370 53636 510624 53664
rect 460342 48089 460394 48095
rect 460342 48031 460394 48037
rect 418774 43205 418826 43211
rect 418774 43147 418826 43153
rect 444886 43205 444938 43211
rect 444886 43147 444938 43153
rect 458614 43205 458666 43211
rect 458614 43147 458666 43153
rect 415220 41986 415276 41995
rect 415220 41921 415276 41930
rect 415234 41810 415262 41921
rect 416852 41838 416908 41847
rect 416592 41796 416852 41824
rect 416852 41773 416908 41782
rect 420788 40506 420844 40515
rect 420788 40441 420844 40450
rect 403222 37507 403274 37513
rect 403222 37449 403274 37455
rect 365974 37359 366026 37365
rect 365974 37301 366026 37307
rect 389206 37359 389258 37365
rect 389206 37301 389258 37307
rect 311060 37250 311116 37259
rect 311060 37185 311116 37194
rect 328340 37250 328396 37259
rect 328340 37185 328396 37194
rect 420802 34553 420830 40441
rect 444898 34553 444926 43147
rect 460354 42106 460382 48031
rect 472246 47941 472298 47947
rect 472246 47883 472298 47889
rect 464854 46461 464906 46467
rect 464854 46403 464906 46409
rect 464866 41847 464894 46403
rect 472258 44955 472286 47883
rect 475510 47719 475562 47725
rect 475510 47661 475562 47667
rect 472244 44946 472300 44955
rect 472244 44881 472300 44890
rect 471408 42101 471710 42120
rect 471408 42095 471722 42101
rect 471408 42092 471670 42095
rect 471670 42037 471722 42043
rect 464852 41838 464908 41847
rect 470324 41838 470380 41847
rect 470160 41796 470324 41824
rect 464852 41773 464908 41782
rect 470324 41773 470380 41782
rect 475522 37439 475550 47661
rect 475714 46467 475742 53636
rect 480982 48163 481034 48169
rect 480982 48105 481034 48111
rect 475702 46461 475754 46467
rect 475702 46403 475754 46409
rect 480994 42101 481022 48105
rect 492994 48021 493022 53636
rect 510370 48095 510398 53636
rect 527938 48169 527966 53650
rect 527926 48163 527978 48169
rect 527926 48105 527978 48111
rect 510358 48089 510410 48095
rect 510358 48031 510410 48037
rect 492982 48015 493034 48021
rect 492982 47957 493034 47963
rect 506806 47867 506858 47873
rect 506806 47809 506858 47815
rect 506818 44913 506846 47809
rect 529270 47793 529322 47799
rect 529270 47735 529322 47741
rect 520630 47645 520682 47651
rect 520630 47587 520682 47593
rect 506806 44907 506858 44913
rect 506806 44849 506858 44855
rect 512182 44907 512234 44913
rect 512182 44849 512234 44855
rect 480982 42095 481034 42101
rect 480982 42037 481034 42043
rect 512194 41847 512222 44849
rect 518722 43285 518834 43304
rect 518710 43279 518834 43285
rect 518762 43276 518834 43279
rect 518710 43221 518762 43227
rect 520642 42106 520670 47587
rect 521206 47571 521258 47577
rect 521206 47513 521258 47519
rect 521218 43304 521246 47513
rect 521218 43276 521534 43304
rect 521506 42120 521534 43276
rect 521506 42092 521856 42120
rect 529282 42106 529310 47735
rect 545218 46245 545246 53650
rect 562498 47947 562526 53650
rect 579796 53602 579852 54402
rect 597092 53602 597148 54402
rect 614388 53602 614444 54402
rect 631684 53602 631740 54402
rect 562486 47941 562538 47947
rect 562486 47883 562538 47889
rect 539734 46239 539786 46245
rect 539734 46181 539786 46187
rect 545206 46239 545258 46245
rect 545206 46181 545258 46187
rect 512180 41838 512236 41847
rect 525908 41838 525964 41847
rect 514882 41805 515136 41824
rect 512180 41773 512236 41782
rect 514006 41799 514058 41805
rect 514006 41741 514058 41747
rect 514870 41799 515136 41805
rect 514922 41796 515136 41799
rect 525964 41796 526176 41824
rect 525908 41773 525964 41782
rect 514870 41741 514922 41747
rect 514018 37439 514046 41741
rect 539746 40515 539774 46181
rect 640738 43729 640766 96501
rect 645428 96006 645484 96015
rect 645428 95941 645430 95950
rect 645482 95941 645484 95950
rect 645430 95909 645482 95915
rect 646486 92415 646538 92421
rect 646486 92357 646538 92363
rect 645526 92341 645578 92347
rect 645526 92283 645578 92289
rect 645538 79439 645566 92283
rect 645908 88902 645964 88911
rect 645908 88837 645964 88846
rect 645922 87537 645950 88837
rect 645910 87531 645962 87537
rect 645910 87473 645962 87479
rect 645908 84462 645964 84471
rect 645908 84397 645964 84406
rect 645922 84059 645950 84397
rect 645910 84053 645962 84059
rect 645910 83995 645962 84001
rect 645524 79430 645580 79439
rect 645524 79365 645580 79374
rect 646006 76135 646058 76141
rect 646006 76077 646058 76083
rect 646018 75591 646046 76077
rect 646004 75582 646060 75591
rect 646004 75517 646060 75526
rect 646004 66258 646060 66267
rect 646004 66193 646006 66202
rect 646058 66193 646060 66202
rect 646006 66161 646058 66167
rect 646006 59115 646058 59121
rect 646006 59057 646058 59063
rect 646018 59015 646046 59057
rect 646004 59006 646060 59015
rect 646004 58941 646060 58950
rect 646498 54723 646526 92357
rect 646594 77695 646622 113109
rect 647156 111398 647212 111407
rect 647156 111333 647212 111342
rect 646676 109474 646732 109483
rect 646676 109409 646732 109418
rect 646582 77689 646634 77695
rect 646582 77631 646634 77637
rect 646690 77621 646718 109409
rect 646772 107994 646828 108003
rect 646772 107929 646828 107938
rect 646786 92717 646814 107929
rect 646964 98078 647020 98087
rect 646964 98013 647020 98022
rect 646774 92711 646826 92717
rect 646774 92653 646826 92659
rect 646870 92267 646922 92273
rect 646870 92209 646922 92215
rect 646774 83609 646826 83615
rect 646774 83551 646826 83557
rect 646678 77615 646730 77621
rect 646678 77557 646730 77563
rect 646786 57091 646814 83551
rect 646882 68635 646910 92209
rect 646978 77769 647006 98013
rect 647062 92193 647114 92199
rect 647062 92135 647114 92141
rect 646966 77763 647018 77769
rect 646966 77705 647018 77711
rect 647074 71891 647102 92135
rect 647170 87093 647198 111333
rect 665314 105191 665342 115223
rect 668194 106375 668222 277833
rect 669538 275391 669566 700785
rect 670678 700103 670730 700109
rect 670678 700045 670730 700051
rect 669718 696995 669770 697001
rect 669718 696937 669770 696943
rect 669622 611155 669674 611161
rect 669622 611097 669674 611103
rect 669524 275382 669580 275391
rect 669524 275317 669580 275326
rect 669634 263551 669662 611097
rect 669730 275243 669758 696937
rect 670690 656523 670718 700045
rect 670978 699739 671006 876165
rect 673270 724967 673322 724973
rect 673270 724909 673322 724915
rect 672886 720749 672938 720755
rect 672886 720691 672938 720697
rect 670966 699733 671018 699739
rect 670966 699675 671018 699681
rect 670870 699141 670922 699147
rect 670870 699083 670922 699089
rect 670774 691223 670826 691229
rect 670774 691165 670826 691171
rect 670786 657633 670814 691165
rect 670882 679694 670910 699083
rect 670978 697001 671006 699675
rect 670966 696995 671018 697001
rect 670966 696937 671018 696943
rect 672406 685377 672458 685383
rect 672406 685319 672458 685325
rect 672214 680789 672266 680795
rect 672214 680731 672266 680737
rect 670882 679666 671006 679694
rect 670774 657627 670826 657633
rect 670774 657569 670826 657575
rect 670678 656517 670730 656523
rect 670678 656459 670730 656465
rect 670690 655265 670718 656459
rect 670870 656073 670922 656079
rect 670870 656015 670922 656021
rect 670678 655259 670730 655265
rect 670678 655201 670730 655207
rect 670774 654815 670826 654821
rect 670774 654757 670826 654763
rect 669814 611895 669866 611901
rect 669814 611837 669866 611843
rect 669716 275234 669772 275243
rect 669716 275169 669772 275178
rect 669826 264989 669854 611837
rect 670582 611673 670634 611679
rect 670582 611615 670634 611621
rect 670594 567131 670622 611615
rect 670786 611161 670814 654757
rect 670882 611901 670910 656015
rect 670978 655783 671006 679666
rect 670966 655777 671018 655783
rect 670966 655719 671018 655725
rect 670978 655339 671006 655719
rect 670966 655333 671018 655339
rect 670966 655275 671018 655281
rect 670966 637869 671018 637875
rect 670966 637811 671018 637817
rect 670870 611895 670922 611901
rect 670870 611837 670922 611843
rect 670774 611155 670826 611161
rect 670774 611097 670826 611103
rect 670678 610637 670730 610643
rect 670678 610579 670730 610585
rect 670102 567125 670154 567131
rect 670102 567067 670154 567073
rect 670582 567125 670634 567131
rect 670582 567067 670634 567073
rect 669910 565941 669962 565947
rect 669910 565883 669962 565889
rect 669922 277463 669950 565883
rect 670006 479435 670058 479441
rect 670006 479377 670058 479383
rect 669908 277454 669964 277463
rect 669908 277389 669964 277398
rect 670018 270655 670046 479377
rect 670114 277611 670142 567067
rect 670690 565947 670718 610579
rect 670870 567495 670922 567501
rect 670870 567437 670922 567443
rect 670678 565941 670730 565947
rect 670678 565883 670730 565889
rect 670882 524063 670910 567437
rect 670978 561507 671006 637811
rect 672118 612635 672170 612641
rect 672118 612577 672170 612583
rect 672130 578971 672158 612577
rect 672226 604723 672254 680731
rect 672310 675165 672362 675171
rect 672310 675107 672362 675113
rect 672322 605759 672350 675107
rect 672418 607239 672446 685319
rect 672694 682121 672746 682127
rect 672694 682063 672746 682069
rect 672502 677089 672554 677095
rect 672502 677031 672554 677037
rect 672406 607233 672458 607239
rect 672406 607175 672458 607181
rect 672310 605753 672362 605759
rect 672310 605695 672362 605701
rect 672514 605167 672542 677031
rect 672598 630765 672650 630771
rect 672598 630707 672650 630713
rect 672502 605161 672554 605167
rect 672502 605103 672554 605109
rect 672214 604717 672266 604723
rect 672214 604659 672266 604665
rect 672310 592137 672362 592143
rect 672310 592079 672362 592085
rect 672214 588585 672266 588591
rect 672214 588527 672266 588533
rect 672118 578965 672170 578971
rect 672118 578907 672170 578913
rect 670966 561501 671018 561507
rect 670966 561443 671018 561449
rect 670870 524057 670922 524063
rect 670870 523999 670922 524005
rect 672226 516219 672254 588527
rect 672214 516213 672266 516219
rect 672214 516155 672266 516161
rect 672322 515479 672350 592079
rect 672406 566311 672458 566317
rect 672406 566253 672458 566259
rect 672418 523915 672446 566253
rect 672502 565423 672554 565429
rect 672502 565365 672554 565371
rect 672406 523909 672458 523915
rect 672406 523851 672458 523857
rect 672310 515473 672362 515479
rect 672310 515415 672362 515421
rect 670294 479139 670346 479145
rect 670294 479081 670346 479087
rect 670306 278351 670334 479081
rect 670484 348642 670540 348651
rect 670484 348577 670540 348586
rect 670292 278342 670348 278351
rect 670292 278277 670348 278286
rect 670498 278203 670526 348577
rect 670484 278194 670540 278203
rect 670484 278129 670540 278138
rect 670100 277602 670156 277611
rect 670100 277537 670156 277546
rect 672418 276279 672446 523851
rect 672514 521251 672542 565365
rect 672610 560767 672638 630707
rect 672706 606721 672734 682063
rect 672898 648087 672926 720691
rect 672982 681307 673034 681313
rect 672982 681249 673034 681255
rect 672886 648081 672938 648087
rect 672886 648023 672938 648029
rect 672790 633651 672842 633657
rect 672790 633593 672842 633599
rect 672694 606715 672746 606721
rect 672694 606657 672746 606663
rect 672694 586513 672746 586519
rect 672694 586455 672746 586461
rect 672598 560761 672650 560767
rect 672598 560703 672650 560709
rect 672502 521245 672554 521251
rect 672502 521187 672554 521193
rect 672514 278499 672542 521187
rect 672706 516515 672734 586455
rect 672802 559065 672830 633593
rect 672886 632393 672938 632399
rect 672886 632335 672938 632341
rect 672790 559059 672842 559065
rect 672790 559001 672842 559007
rect 672898 558695 672926 632335
rect 672994 606351 673022 681249
rect 673078 677607 673130 677613
rect 673078 677549 673130 677555
rect 672982 606345 673034 606351
rect 672982 606287 673034 606293
rect 673090 604427 673118 677549
rect 673174 676719 673226 676725
rect 673174 676661 673226 676667
rect 673078 604421 673130 604427
rect 673078 604363 673130 604369
rect 673186 603687 673214 676661
rect 673282 649271 673310 724909
rect 673378 714243 673406 878385
rect 676244 877298 676300 877307
rect 676244 877233 676246 877242
rect 676298 877233 676300 877242
rect 676246 877201 676298 877207
rect 676244 876262 676300 876271
rect 676244 876197 676246 876206
rect 676298 876197 676300 876206
rect 676246 876165 676298 876171
rect 680276 875670 680332 875679
rect 680276 875605 680332 875614
rect 676052 875522 676108 875531
rect 676052 875457 676108 875466
rect 674038 872745 674090 872751
rect 674038 872687 674090 872693
rect 674050 858321 674078 872687
rect 676066 872677 676094 875457
rect 679796 875078 679852 875087
rect 679796 875013 679852 875022
rect 676244 873746 676300 873755
rect 676244 873681 676300 873690
rect 676258 872751 676286 873681
rect 676246 872745 676298 872751
rect 676246 872687 676298 872693
rect 679700 872710 679756 872719
rect 674326 872671 674378 872677
rect 674326 872613 674378 872619
rect 676054 872671 676106 872677
rect 679700 872645 679756 872654
rect 676054 872613 676106 872619
rect 674134 870155 674186 870161
rect 674134 870097 674186 870103
rect 674038 858315 674090 858321
rect 674038 858257 674090 858263
rect 674146 852179 674174 870097
rect 674230 863199 674282 863205
rect 674230 863141 674282 863147
rect 674242 858173 674270 863141
rect 674230 858167 674282 858173
rect 674230 858109 674282 858115
rect 674134 852173 674186 852179
rect 674134 852115 674186 852121
rect 674338 850181 674366 872613
rect 676052 871526 676108 871535
rect 676052 871461 676108 871470
rect 676066 870161 676094 871461
rect 676244 870786 676300 870795
rect 676244 870721 676300 870730
rect 676054 870155 676106 870161
rect 676054 870097 676106 870103
rect 676052 870046 676108 870055
rect 676052 869981 676108 869990
rect 674902 869933 674954 869939
rect 674902 869875 674954 869881
rect 674518 867047 674570 867053
rect 674518 866989 674570 866995
rect 674422 863125 674474 863131
rect 674422 863067 674474 863073
rect 674434 857729 674462 863067
rect 674422 857723 674474 857729
rect 674422 857665 674474 857671
rect 674530 853215 674558 866989
rect 674914 866036 674942 869875
rect 676066 869865 676094 869981
rect 676258 869939 676286 870721
rect 676246 869933 676298 869939
rect 676246 869875 676298 869881
rect 675094 869859 675146 869865
rect 675094 869801 675146 869807
rect 676054 869859 676106 869865
rect 676054 869801 676106 869807
rect 674998 869785 675050 869791
rect 674998 869727 675050 869733
rect 674818 866008 674942 866036
rect 674614 864309 674666 864315
rect 674614 864251 674666 864257
rect 674626 861873 674654 864251
rect 674614 861867 674666 861873
rect 674614 861809 674666 861815
rect 674614 861275 674666 861281
rect 674614 861217 674666 861223
rect 674518 853209 674570 853215
rect 674518 853151 674570 853157
rect 674626 850921 674654 861217
rect 674818 857304 674846 866008
rect 675010 864297 675038 869727
rect 674914 864269 675038 864297
rect 674914 862021 674942 864269
rect 674998 864235 675050 864241
rect 674998 864177 675050 864183
rect 674902 862015 674954 862021
rect 674902 861957 674954 861963
rect 674902 861867 674954 861873
rect 674902 861809 674954 861815
rect 674914 858765 674942 861809
rect 675010 859579 675038 864177
rect 674998 859573 675050 859579
rect 674998 859515 675050 859521
rect 674902 858759 674954 858765
rect 674902 858701 674954 858707
rect 674998 858315 675050 858321
rect 674998 858257 675050 858263
rect 674818 857276 674942 857304
rect 674914 854029 674942 857276
rect 675010 855213 675038 858257
rect 674998 855207 675050 855213
rect 674998 855149 675050 855155
rect 675106 854547 675134 869801
rect 679714 869791 679742 872645
rect 679702 869785 679754 869791
rect 679702 869727 679754 869733
rect 679810 869717 679838 875013
rect 680180 874190 680236 874199
rect 680180 874125 680236 874134
rect 679892 872118 679948 872127
rect 679892 872053 679948 872062
rect 675190 869711 675242 869717
rect 675190 869653 675242 869659
rect 679798 869711 679850 869717
rect 679798 869653 679850 869659
rect 675202 862465 675230 869653
rect 676244 869306 676300 869315
rect 676244 869241 676300 869250
rect 676258 867053 676286 869241
rect 679796 868714 679852 868723
rect 679796 868649 679852 868658
rect 679810 868279 679838 868649
rect 679796 868270 679852 868279
rect 679796 868205 679852 868214
rect 676246 867047 676298 867053
rect 676246 866989 676298 866995
rect 679810 866979 679838 868205
rect 679798 866973 679850 866979
rect 679798 866915 679850 866921
rect 679906 864315 679934 872053
rect 680084 871674 680140 871683
rect 680084 871609 680140 871618
rect 679988 870194 680044 870203
rect 679988 870129 680044 870138
rect 679894 864309 679946 864315
rect 679894 864251 679946 864257
rect 675286 864161 675338 864167
rect 675286 864103 675338 864109
rect 675190 862459 675242 862465
rect 675190 862401 675242 862407
rect 675190 861201 675242 861207
rect 675190 861143 675242 861149
rect 675094 854541 675146 854547
rect 675094 854483 675146 854489
rect 674902 854023 674954 854029
rect 674902 853965 674954 853971
rect 675202 852771 675230 861143
rect 675298 860856 675326 864103
rect 675478 864087 675530 864093
rect 675478 864029 675530 864035
rect 675490 862692 675518 864029
rect 680002 863131 680030 870129
rect 680098 863205 680126 871609
rect 680194 864241 680222 874125
rect 680182 864235 680234 864241
rect 680182 864177 680234 864183
rect 680290 864167 680318 875605
rect 685460 868270 685516 868279
rect 685460 868205 685516 868214
rect 685474 867835 685502 868205
rect 685460 867826 685516 867835
rect 685460 867761 685516 867770
rect 680278 864161 680330 864167
rect 680278 864103 680330 864109
rect 680086 863199 680138 863205
rect 680086 863141 680138 863147
rect 679990 863125 680042 863131
rect 679990 863067 680042 863073
rect 675382 862459 675434 862465
rect 675382 862401 675434 862407
rect 675394 862100 675422 862401
rect 675382 862015 675434 862021
rect 675382 861957 675434 861963
rect 675394 861479 675422 861957
rect 675298 860828 675408 860856
rect 675478 859573 675530 859579
rect 675478 859515 675530 859521
rect 675490 858992 675518 859515
rect 675382 858759 675434 858765
rect 675382 858701 675434 858707
rect 675394 858443 675422 858701
rect 675478 858167 675530 858173
rect 675478 858109 675530 858115
rect 675490 857808 675518 858109
rect 675382 857723 675434 857729
rect 675382 857665 675434 857671
rect 675394 857142 675422 857665
rect 675382 855207 675434 855213
rect 675382 855149 675434 855155
rect 675394 854671 675422 855149
rect 675382 854541 675434 854547
rect 675382 854483 675434 854489
rect 675394 854108 675422 854483
rect 675382 854023 675434 854029
rect 675382 853965 675434 853971
rect 675394 853475 675422 853965
rect 675478 853209 675530 853215
rect 675478 853151 675530 853157
rect 675490 852850 675518 853151
rect 675190 852765 675242 852771
rect 675190 852707 675242 852713
rect 675382 852765 675434 852771
rect 675382 852707 675434 852713
rect 675188 852582 675244 852591
rect 675188 852517 675244 852526
rect 674614 850915 674666 850921
rect 674614 850857 674666 850863
rect 674326 850175 674378 850181
rect 674326 850117 674378 850123
rect 675202 848479 675230 852517
rect 675394 852258 675422 852707
rect 675382 852173 675434 852179
rect 675382 852115 675434 852121
rect 675394 851635 675422 852115
rect 675382 850915 675434 850921
rect 675382 850857 675434 850863
rect 675394 850439 675422 850857
rect 675478 850175 675530 850181
rect 675478 850117 675530 850123
rect 675490 849816 675518 850117
rect 675190 848473 675242 848479
rect 675190 848415 675242 848421
rect 675478 848473 675530 848479
rect 675478 848415 675530 848421
rect 675490 847966 675518 848415
rect 675394 774849 675422 775298
rect 675382 774843 675434 774849
rect 675382 774785 675434 774791
rect 675490 774595 675518 774706
rect 675476 774586 675532 774595
rect 675476 774521 675532 774530
rect 675394 773707 675422 774079
rect 675380 773698 675436 773707
rect 675380 773633 675436 773642
rect 675778 773115 675806 773448
rect 675764 773106 675820 773115
rect 675764 773041 675820 773050
rect 674998 771957 675050 771963
rect 674998 771899 675050 771905
rect 674230 771365 674282 771371
rect 674230 771307 674282 771313
rect 674134 766333 674186 766339
rect 674134 766275 674186 766281
rect 673942 724375 673994 724381
rect 673942 724317 673994 724323
rect 673954 723419 673982 724317
rect 673942 723413 673994 723419
rect 673942 723355 673994 723361
rect 674038 721193 674090 721199
rect 674038 721135 674090 721141
rect 673366 714237 673418 714243
rect 673366 714179 673418 714185
rect 674050 709951 674078 721135
rect 674038 709945 674090 709951
rect 674038 709887 674090 709893
rect 674146 693671 674174 766275
rect 674242 699221 674270 771307
rect 674422 766851 674474 766857
rect 674422 766793 674474 766799
rect 674326 765741 674378 765747
rect 674326 765683 674378 765689
rect 674230 699215 674282 699221
rect 674230 699157 674282 699163
rect 674338 694041 674366 765683
rect 674434 696853 674462 766793
rect 674518 765149 674570 765155
rect 674518 765091 674570 765097
rect 674530 731675 674558 765091
rect 674902 763743 674954 763749
rect 674902 763685 674954 763691
rect 674914 762288 674942 763685
rect 675010 763527 675038 771899
rect 675094 771883 675146 771889
rect 675094 771825 675146 771831
rect 675106 765303 675134 771825
rect 675394 771371 675422 771598
rect 675382 771365 675434 771371
rect 675382 771307 675434 771313
rect 675778 770747 675806 771043
rect 675764 770738 675820 770747
rect 675764 770673 675820 770682
rect 675490 770007 675518 770414
rect 675476 769998 675532 770007
rect 675476 769933 675532 769942
rect 675490 769415 675518 769748
rect 675476 769406 675532 769415
rect 675476 769341 675532 769350
rect 675394 766857 675422 767271
rect 675382 766851 675434 766857
rect 675382 766793 675434 766799
rect 675490 766339 675518 766714
rect 675478 766333 675530 766339
rect 675478 766275 675530 766281
rect 675490 765747 675518 766048
rect 675478 765741 675530 765747
rect 675478 765683 675530 765689
rect 675094 765297 675146 765303
rect 675094 765239 675146 765245
rect 675382 765297 675434 765303
rect 675382 765239 675434 765245
rect 675394 764864 675422 765239
rect 675490 765155 675518 765456
rect 675478 765149 675530 765155
rect 675478 765091 675530 765097
rect 675394 763749 675422 764235
rect 675382 763743 675434 763749
rect 675382 763685 675434 763691
rect 674998 763521 675050 763527
rect 674998 763463 675050 763469
rect 675382 763521 675434 763527
rect 675382 763463 675434 763469
rect 675394 763014 675422 763463
rect 674818 762260 674942 762288
rect 674516 731666 674572 731675
rect 674516 731601 674572 731610
rect 674614 727187 674666 727193
rect 674614 727129 674666 727135
rect 674518 722451 674570 722457
rect 674518 722393 674570 722399
rect 674530 719516 674558 722393
rect 674626 720903 674654 727129
rect 674614 720897 674666 720903
rect 674614 720839 674666 720845
rect 674530 719488 674654 719516
rect 674518 719343 674570 719349
rect 674518 719285 674570 719291
rect 674422 696847 674474 696853
rect 674422 696789 674474 696795
rect 674326 694035 674378 694041
rect 674326 693977 674378 693983
rect 674134 693665 674186 693671
rect 674134 693607 674186 693613
rect 674326 689817 674378 689823
rect 674326 689759 674378 689765
rect 674038 686265 674090 686271
rect 674038 686207 674090 686213
rect 674050 685605 674078 686207
rect 674038 685599 674090 685605
rect 674038 685541 674090 685547
rect 674338 676915 674366 689759
rect 674422 681159 674474 681165
rect 674422 681101 674474 681107
rect 674324 676906 674380 676915
rect 674324 676841 674380 676850
rect 674434 676207 674462 681101
rect 674422 676201 674474 676207
rect 674422 676143 674474 676149
rect 673750 656961 673802 656967
rect 673750 656903 673802 656909
rect 673270 649265 673322 649271
rect 673270 649207 673322 649213
rect 673366 637129 673418 637135
rect 673366 637071 673418 637077
rect 673270 636537 673322 636543
rect 673270 636479 673322 636485
rect 673174 603681 673226 603687
rect 673174 603623 673226 603629
rect 672982 592729 673034 592735
rect 672982 592671 673034 592677
rect 672886 558689 672938 558695
rect 672886 558631 672938 558637
rect 672886 549143 672938 549149
rect 672886 549085 672938 549091
rect 672790 544925 672842 544931
rect 672790 544867 672842 544873
rect 672694 516509 672746 516515
rect 672694 516451 672746 516457
rect 672802 472263 672830 544867
rect 672898 474705 672926 549085
rect 672994 516959 673022 592671
rect 673174 589029 673226 589035
rect 673174 588971 673226 588977
rect 673078 587993 673130 587999
rect 673078 587935 673130 587941
rect 672982 516953 673034 516959
rect 672982 516895 673034 516901
rect 673090 514517 673118 587935
rect 673186 515035 673214 588971
rect 673282 559435 673310 636479
rect 673378 560915 673406 637071
rect 673762 613233 673790 656903
rect 674530 650899 674558 719285
rect 674626 653785 674654 719488
rect 674818 696724 674846 762260
rect 675394 761899 675422 762422
rect 674998 761893 675050 761899
rect 674998 761835 675050 761841
rect 675382 761893 675434 761899
rect 675382 761835 675434 761841
rect 674902 760339 674954 760345
rect 674902 760281 674954 760287
rect 674914 696927 674942 760281
rect 675010 698999 675038 761835
rect 675394 760345 675422 760572
rect 675382 760339 675434 760345
rect 675382 760281 675434 760287
rect 675394 730468 675422 730898
rect 675298 730440 675422 730468
rect 675298 728747 675326 730440
rect 675490 729899 675518 730306
rect 675476 729890 675532 729899
rect 675476 729825 675532 729834
rect 675778 729455 675806 729679
rect 675764 729446 675820 729455
rect 675764 729381 675820 729390
rect 675286 728741 675338 728747
rect 675682 728715 675710 729048
rect 675286 728683 675338 728689
rect 675668 728706 675724 728715
rect 675668 728641 675724 728650
rect 675394 726791 675422 727198
rect 675380 726782 675436 726791
rect 675380 726717 675436 726726
rect 675778 726199 675806 726643
rect 675764 726190 675820 726199
rect 675764 726125 675820 726134
rect 675394 725903 675422 726014
rect 675380 725894 675436 725903
rect 675380 725829 675436 725838
rect 675490 724973 675518 725348
rect 675478 724967 675530 724973
rect 675478 724909 675530 724915
rect 675286 723413 675338 723419
rect 675286 723355 675338 723361
rect 675298 719072 675326 723355
rect 675394 722457 675422 722871
rect 675382 722451 675434 722457
rect 675382 722393 675434 722399
rect 675778 721907 675806 722314
rect 675764 721898 675820 721907
rect 675764 721833 675820 721842
rect 675490 721199 675518 721648
rect 675478 721193 675530 721199
rect 675478 721135 675530 721141
rect 675382 720897 675434 720903
rect 675382 720839 675434 720845
rect 675394 720464 675422 720839
rect 675490 720755 675518 721056
rect 675478 720749 675530 720755
rect 675478 720691 675530 720697
rect 675394 719349 675422 719835
rect 675382 719343 675434 719349
rect 675382 719285 675434 719291
rect 675298 719044 675422 719072
rect 675394 718614 675422 719044
rect 675298 718156 675518 718184
rect 675298 715649 675326 718156
rect 675490 718022 675518 718156
rect 675394 715649 675422 716172
rect 675286 715643 675338 715649
rect 675286 715585 675338 715591
rect 675382 715643 675434 715649
rect 675382 715585 675434 715591
rect 675382 715421 675434 715427
rect 675382 715363 675434 715369
rect 674998 698993 675050 698999
rect 674998 698935 675050 698941
rect 674902 696921 674954 696927
rect 674902 696863 674954 696869
rect 674818 696705 674942 696724
rect 674818 696699 674954 696705
rect 674818 696696 674902 696699
rect 674902 696641 674954 696647
rect 675394 689768 675422 715363
rect 675574 715347 675626 715353
rect 675574 715289 675626 715295
rect 675202 689740 675422 689768
rect 674998 689447 675050 689453
rect 674998 689389 675050 689395
rect 674902 681233 674954 681239
rect 674902 681175 674954 681181
rect 674914 679685 674942 681175
rect 674902 679679 674954 679685
rect 674902 679621 674954 679627
rect 675010 679112 675038 689389
rect 674818 679084 675038 679112
rect 675202 679093 675230 689740
rect 675586 689453 675614 715289
rect 679702 714237 679754 714243
rect 679702 714179 679754 714185
rect 675670 709945 675722 709951
rect 675670 709887 675722 709893
rect 675682 689823 675710 709887
rect 676244 703102 676300 703111
rect 676244 703037 676246 703046
rect 676298 703037 676300 703046
rect 676246 703005 676298 703011
rect 676244 702954 676300 702963
rect 676244 702889 676246 702898
rect 676298 702889 676300 702898
rect 676246 702857 676298 702863
rect 676052 702214 676108 702223
rect 676052 702149 676108 702158
rect 676066 699887 676094 702149
rect 679714 701631 679742 714179
rect 679700 701622 679756 701631
rect 679700 701557 679756 701566
rect 676244 700882 676300 700891
rect 676244 700817 676246 700826
rect 676298 700817 676300 700826
rect 679700 700882 679756 700891
rect 679700 700817 679756 700826
rect 676246 700785 676298 700791
rect 676244 700142 676300 700151
rect 676244 700077 676246 700086
rect 676298 700077 676300 700086
rect 676246 700045 676298 700051
rect 676054 699881 676106 699887
rect 676054 699823 676106 699829
rect 676052 699772 676108 699781
rect 676052 699707 676054 699716
rect 676106 699707 676108 699716
rect 676054 699675 676106 699681
rect 676052 699254 676108 699263
rect 676052 699189 676108 699198
rect 676246 699215 676298 699221
rect 676066 699147 676094 699189
rect 676246 699157 676298 699163
rect 676054 699141 676106 699147
rect 676054 699083 676106 699089
rect 676054 698993 676106 698999
rect 676054 698935 676106 698941
rect 676066 698227 676094 698935
rect 676052 698218 676108 698227
rect 676052 698153 676108 698162
rect 676258 697487 676286 699157
rect 676244 697478 676300 697487
rect 676244 697413 676300 697422
rect 676054 696921 676106 696927
rect 676054 696863 676106 696869
rect 675958 696847 676010 696853
rect 675958 696789 676010 696795
rect 675970 696747 675998 696789
rect 675956 696738 676012 696747
rect 675956 696673 676012 696682
rect 676066 696229 676094 696863
rect 676246 696699 676298 696705
rect 676246 696641 676298 696647
rect 676052 696220 676108 696229
rect 676052 696155 676108 696164
rect 676258 694527 676286 696641
rect 676244 694518 676300 694527
rect 676244 694453 676300 694462
rect 676054 694035 676106 694041
rect 676054 693977 676106 693983
rect 676066 693787 676094 693977
rect 676052 693778 676108 693787
rect 676052 693713 676108 693722
rect 676054 693665 676106 693671
rect 676054 693607 676106 693613
rect 676066 692825 676094 693607
rect 676052 692816 676108 692825
rect 676052 692751 676108 692760
rect 679714 691229 679742 700817
rect 679988 691558 680044 691567
rect 679988 691493 680044 691502
rect 679702 691223 679754 691229
rect 679702 691165 679754 691171
rect 680002 690975 680030 691493
rect 679796 690966 679852 690975
rect 679796 690901 679852 690910
rect 679988 690966 680044 690975
rect 679988 690901 680044 690910
rect 679810 690531 679838 690901
rect 679796 690522 679852 690531
rect 679796 690457 679852 690466
rect 675670 689817 675722 689823
rect 675670 689759 675722 689765
rect 675574 689447 675626 689453
rect 675574 689389 675626 689395
rect 680002 688417 680030 690901
rect 679990 688411 680042 688417
rect 679990 688353 680042 688359
rect 675394 686271 675422 686675
rect 675382 686265 675434 686271
rect 675382 686207 675434 686213
rect 675394 685647 675422 686128
rect 675380 685638 675436 685647
rect 675380 685573 675436 685582
rect 675490 685383 675518 685462
rect 675478 685377 675530 685383
rect 675478 685319 675530 685325
rect 675778 684463 675806 684835
rect 675764 684454 675820 684463
rect 675764 684389 675820 684398
rect 675586 682687 675614 683020
rect 675572 682678 675628 682687
rect 675572 682613 675628 682622
rect 675490 682127 675518 682428
rect 675478 682121 675530 682127
rect 675478 682063 675530 682069
rect 675394 681313 675422 681799
rect 675382 681307 675434 681313
rect 675382 681249 675434 681255
rect 675394 680795 675422 681170
rect 675382 680789 675434 680795
rect 675382 680731 675434 680737
rect 675286 679679 675338 679685
rect 675286 679621 675338 679627
rect 675190 679087 675242 679093
rect 674818 678816 674846 679084
rect 675190 679029 675242 679035
rect 674998 678865 675050 678871
rect 674818 678788 674942 678816
rect 674998 678807 675050 678813
rect 674914 669695 674942 678788
rect 674902 669689 674954 669695
rect 674902 669631 674954 669637
rect 675010 669621 675038 678807
rect 675298 676300 675326 679621
rect 675778 678395 675806 678654
rect 675764 678386 675820 678395
rect 675764 678321 675820 678330
rect 675394 677613 675422 678136
rect 675382 677607 675434 677613
rect 675382 677549 675434 677555
rect 675490 677095 675518 677470
rect 675478 677089 675530 677095
rect 675478 677031 675530 677037
rect 675490 676725 675518 676804
rect 675478 676719 675530 676725
rect 675478 676661 675530 676667
rect 675298 676272 675408 676300
rect 675286 676201 675338 676207
rect 675286 676143 675338 676149
rect 675298 674450 675326 676143
rect 675490 675171 675518 675620
rect 675478 675165 675530 675171
rect 675478 675107 675530 675113
rect 675298 674422 675408 674450
rect 675490 673363 675518 673770
rect 675476 673354 675532 673363
rect 675476 673289 675532 673298
rect 675298 671941 675408 671969
rect 675298 671439 675326 671941
rect 675284 671430 675340 671439
rect 675284 671365 675340 671374
rect 675574 669689 675626 669695
rect 675574 669631 675626 669637
rect 674998 669615 675050 669621
rect 674998 669557 675050 669563
rect 675478 669615 675530 669621
rect 675478 669557 675530 669563
rect 674614 653779 674666 653785
rect 674614 653721 674666 653727
rect 675490 652051 675518 669557
rect 675586 654123 675614 669631
rect 676148 658850 676204 658859
rect 676148 658785 676204 658794
rect 676054 657627 676106 657633
rect 676052 657592 676054 657601
rect 676106 657592 676108 657601
rect 676052 657527 676108 657536
rect 676162 657189 676190 658785
rect 676340 658258 676396 658267
rect 676340 658193 676396 658202
rect 676244 657814 676300 657823
rect 676244 657749 676300 657758
rect 676150 657183 676202 657189
rect 676150 657125 676202 657131
rect 676052 657074 676108 657083
rect 676258 657041 676286 657749
rect 676052 657009 676108 657018
rect 676246 657035 676298 657041
rect 676066 656967 676094 657009
rect 676246 656977 676298 656983
rect 676054 656961 676106 656967
rect 676054 656903 676106 656909
rect 676354 656893 676382 658193
rect 676342 656887 676394 656893
rect 676342 656829 676394 656835
rect 676054 656517 676106 656523
rect 676052 656482 676054 656491
rect 676106 656482 676108 656491
rect 676052 656417 676108 656426
rect 676052 656112 676108 656121
rect 676052 656047 676054 656056
rect 676106 656047 676108 656056
rect 676054 656015 676106 656021
rect 676246 655777 676298 655783
rect 676244 655742 676246 655751
rect 676298 655742 676300 655751
rect 676244 655677 676300 655686
rect 676244 654854 676300 654863
rect 676244 654789 676246 654798
rect 676298 654789 676300 654798
rect 676246 654757 676298 654763
rect 675572 654114 675628 654123
rect 675572 654049 675628 654058
rect 676054 653779 676106 653785
rect 676054 653721 676106 653727
rect 676066 652569 676094 653721
rect 676052 652560 676108 652569
rect 676052 652495 676108 652504
rect 675476 652042 675532 652051
rect 675476 651977 675532 651986
rect 674518 650893 674570 650899
rect 674518 650835 674570 650841
rect 676054 650893 676106 650899
rect 676054 650835 676106 650841
rect 676066 650127 676094 650835
rect 676052 650118 676108 650127
rect 676052 650053 676108 650062
rect 676246 649265 676298 649271
rect 676244 649230 676246 649239
rect 676298 649230 676300 649239
rect 676244 649165 676300 649174
rect 676054 648081 676106 648087
rect 676052 648046 676054 648055
rect 676106 648046 676108 648055
rect 676052 647981 676108 647990
rect 679796 647306 679852 647315
rect 679796 647241 679852 647250
rect 679810 646871 679838 647241
rect 679796 646862 679852 646871
rect 679796 646797 679852 646806
rect 685460 646862 685516 646871
rect 685460 646797 685516 646806
rect 679810 645201 679838 646797
rect 685474 646427 685502 646797
rect 685460 646418 685516 646427
rect 685460 646353 685516 646362
rect 679798 645195 679850 645201
rect 679798 645137 679850 645143
rect 675202 642454 675408 642482
rect 675202 642241 675230 642454
rect 675190 642235 675242 642241
rect 675190 642177 675242 642183
rect 675778 641691 675806 641950
rect 675764 641682 675820 641691
rect 675764 641617 675820 641626
rect 675202 641270 675408 641298
rect 675202 640211 675230 641270
rect 675490 640359 675518 640618
rect 675476 640350 675532 640359
rect 675476 640285 675532 640294
rect 675188 640202 675244 640211
rect 675188 640137 675244 640146
rect 675490 638435 675518 638768
rect 675476 638426 675532 638435
rect 675476 638361 675532 638370
rect 675394 637875 675422 638250
rect 675382 637869 675434 637875
rect 675382 637811 675434 637817
rect 675490 637135 675518 637584
rect 675478 637129 675530 637135
rect 675478 637071 675530 637077
rect 675190 636685 675242 636691
rect 675190 636627 675242 636633
rect 675202 635748 675230 636627
rect 675394 636543 675422 636955
rect 675382 636537 675434 636543
rect 675382 636479 675434 636485
rect 675202 635720 675326 635748
rect 674998 635057 675050 635063
rect 674998 634999 675050 635005
rect 675010 630697 675038 634999
rect 675298 632093 675326 635720
rect 675394 634143 675422 634476
rect 675380 634134 675436 634143
rect 675380 634069 675436 634078
rect 675394 633657 675422 633919
rect 675382 633651 675434 633657
rect 675382 633593 675434 633599
rect 675778 632811 675806 633292
rect 675764 632802 675820 632811
rect 675764 632737 675820 632746
rect 675490 632399 675518 632626
rect 675478 632393 675530 632399
rect 675478 632335 675530 632341
rect 675298 632065 675408 632093
rect 675298 631428 675408 631456
rect 675298 630771 675326 631428
rect 675286 630765 675338 630771
rect 675286 630707 675338 630713
rect 674998 630691 675050 630697
rect 674998 630633 675050 630639
rect 675478 630691 675530 630697
rect 675478 630633 675530 630639
rect 675490 630258 675518 630633
rect 675778 629111 675806 629592
rect 675764 629102 675820 629111
rect 675764 629037 675820 629046
rect 675778 627335 675806 627742
rect 675764 627326 675820 627335
rect 675764 627261 675820 627270
rect 676148 614450 676204 614459
rect 676148 614385 676204 614394
rect 676052 614154 676108 614163
rect 676052 614089 676108 614098
rect 676066 613677 676094 614089
rect 676162 613825 676190 614385
rect 676246 613967 676298 613973
rect 676246 613909 676298 613915
rect 676258 613867 676286 613909
rect 676244 613858 676300 613867
rect 676150 613819 676202 613825
rect 676244 613793 676300 613802
rect 676150 613761 676202 613767
rect 676054 613671 676106 613677
rect 676054 613613 676106 613619
rect 673750 613227 673802 613233
rect 676054 613227 676106 613233
rect 673750 613169 673802 613175
rect 676052 613192 676054 613201
rect 676106 613192 676108 613201
rect 676052 613127 676108 613136
rect 676052 612674 676108 612683
rect 676052 612609 676054 612618
rect 676106 612609 676108 612618
rect 676054 612577 676106 612583
rect 676244 611934 676300 611943
rect 676244 611869 676246 611878
rect 676298 611869 676300 611878
rect 676246 611837 676298 611843
rect 676052 611712 676108 611721
rect 676052 611647 676054 611656
rect 676106 611647 676108 611656
rect 676054 611615 676106 611621
rect 676052 611194 676108 611203
rect 676052 611129 676054 611138
rect 676106 611129 676108 611138
rect 676054 611097 676106 611103
rect 676054 610637 676106 610643
rect 676052 610602 676054 610611
rect 676106 610602 676108 610611
rect 676052 610537 676108 610546
rect 676054 607233 676106 607239
rect 676052 607198 676054 607207
rect 676106 607198 676108 607207
rect 676052 607133 676108 607142
rect 676054 606715 676106 606721
rect 676052 606680 676054 606689
rect 676106 606680 676108 606689
rect 676052 606615 676108 606624
rect 676246 606345 676298 606351
rect 676244 606310 676246 606319
rect 676298 606310 676300 606319
rect 676244 606245 676300 606254
rect 676054 605753 676106 605759
rect 676052 605718 676054 605727
rect 676106 605718 676108 605727
rect 676052 605653 676108 605662
rect 676054 605161 676106 605167
rect 676052 605126 676054 605135
rect 676106 605126 676108 605135
rect 676052 605061 676108 605070
rect 676054 604717 676106 604723
rect 676052 604682 676054 604691
rect 676106 604682 676108 604691
rect 676052 604617 676108 604626
rect 676246 604421 676298 604427
rect 676244 604386 676246 604395
rect 676298 604386 676300 604395
rect 676244 604321 676300 604330
rect 676054 603681 676106 603687
rect 676052 603646 676054 603655
rect 676106 603646 676108 603655
rect 676052 603581 676108 603590
rect 679988 602906 680044 602915
rect 679988 602841 680044 602850
rect 680002 602471 680030 602841
rect 679796 602462 679852 602471
rect 679796 602397 679852 602406
rect 679988 602462 680044 602471
rect 679988 602397 680044 602406
rect 675382 602053 675434 602059
rect 679810 602027 679838 602397
rect 675382 601995 675434 602001
rect 679796 602018 679852 602027
rect 675394 598068 675422 601995
rect 680002 601985 680030 602397
rect 679796 601953 679852 601962
rect 679990 601979 680042 601985
rect 679990 601921 680042 601927
rect 675394 597143 675422 597550
rect 675380 597134 675436 597143
rect 675380 597069 675436 597078
rect 675394 596361 675422 596884
rect 674902 596355 674954 596361
rect 674902 596297 674954 596303
rect 675382 596355 675434 596361
rect 675382 596297 675434 596303
rect 674914 593568 674942 596297
rect 675490 596107 675518 596218
rect 675476 596098 675532 596107
rect 675476 596033 675532 596042
rect 675490 594035 675518 594368
rect 675476 594026 675532 594035
rect 675476 593961 675532 593970
rect 674818 593540 674942 593568
rect 673654 593321 673706 593327
rect 673654 593263 673706 593269
rect 673366 560909 673418 560915
rect 673366 560851 673418 560857
rect 673270 559429 673322 559435
rect 673270 559371 673322 559377
rect 673366 547959 673418 547965
rect 673366 547901 673418 547907
rect 673270 547293 673322 547299
rect 673270 547235 673322 547241
rect 673174 515029 673226 515035
rect 673174 514971 673226 514977
rect 673078 514511 673130 514517
rect 673078 514453 673130 514459
rect 672886 474699 672938 474705
rect 672886 474641 672938 474647
rect 673282 474335 673310 547235
rect 673270 474329 673322 474335
rect 673270 474271 673322 474277
rect 673378 472855 673406 547901
rect 673666 517699 673694 593263
rect 674818 578894 674846 593540
rect 674902 593395 674954 593401
rect 674902 593337 674954 593343
rect 674914 588147 674942 593337
rect 675394 593327 675422 593850
rect 675382 593321 675434 593327
rect 675382 593263 675434 593269
rect 675490 592735 675518 593184
rect 675478 592729 675530 592735
rect 675478 592671 675530 592677
rect 675394 592143 675422 592555
rect 675382 592137 675434 592143
rect 675382 592079 675434 592085
rect 674998 590509 675050 590515
rect 674998 590451 675050 590457
rect 674902 588141 674954 588147
rect 674902 588083 674954 588089
rect 675010 586297 675038 590451
rect 675490 589743 675518 590076
rect 675476 589734 675532 589743
rect 675476 589669 675532 589678
rect 675394 589035 675422 589519
rect 675382 589029 675434 589035
rect 675382 588971 675434 588977
rect 675394 588591 675422 588892
rect 675382 588585 675434 588591
rect 675382 588527 675434 588533
rect 675382 588141 675434 588147
rect 675382 588083 675434 588089
rect 675394 587679 675422 588083
rect 675490 587999 675518 588226
rect 675478 587993 675530 587999
rect 675478 587935 675530 587941
rect 675394 586519 675422 587042
rect 675382 586513 675434 586519
rect 675382 586455 675434 586461
rect 674998 586291 675050 586297
rect 674998 586233 675050 586239
rect 675478 586291 675530 586297
rect 675478 586233 675530 586239
rect 675490 585858 675518 586233
rect 675778 584711 675806 585192
rect 675764 584702 675820 584711
rect 675764 584637 675820 584646
rect 675682 582935 675710 583342
rect 675668 582926 675724 582935
rect 675668 582861 675724 582870
rect 679702 578965 679754 578971
rect 679702 578907 679754 578913
rect 674818 578866 674942 578894
rect 674914 567247 674942 578866
rect 676244 569310 676300 569319
rect 676244 569245 676300 569254
rect 676148 568570 676204 568579
rect 676148 568505 676204 568514
rect 676052 568422 676108 568431
rect 676052 568357 676108 568366
rect 676066 567945 676094 568357
rect 676054 567939 676106 567945
rect 676054 567881 676106 567887
rect 676054 567495 676106 567501
rect 676052 567460 676054 567469
rect 676106 567460 676108 567469
rect 676162 567427 676190 568505
rect 676258 567797 676286 569245
rect 679714 567839 679742 578907
rect 679700 567830 679756 567839
rect 676246 567791 676298 567797
rect 679700 567765 679756 567774
rect 676246 567733 676298 567739
rect 676052 567395 676108 567404
rect 676150 567421 676202 567427
rect 676150 567363 676202 567369
rect 674900 567238 674956 567247
rect 674900 567173 674956 567182
rect 676246 567125 676298 567131
rect 676244 567090 676246 567099
rect 676298 567090 676300 567099
rect 676244 567025 676300 567034
rect 676244 566350 676300 566359
rect 676244 566285 676246 566294
rect 676298 566285 676300 566294
rect 676246 566253 676298 566259
rect 676054 565941 676106 565947
rect 676052 565906 676054 565915
rect 676106 565906 676108 565915
rect 676052 565841 676108 565850
rect 676052 565462 676108 565471
rect 676052 565397 676054 565406
rect 676106 565397 676108 565406
rect 676054 565365 676106 565371
rect 676054 561501 676106 561507
rect 676052 561466 676054 561475
rect 676106 561466 676108 561475
rect 676052 561401 676108 561410
rect 676054 560909 676106 560915
rect 676052 560874 676054 560883
rect 676106 560874 676108 560883
rect 676052 560809 676108 560818
rect 676246 560761 676298 560767
rect 676244 560726 676246 560735
rect 676298 560726 676300 560735
rect 676244 560661 676300 560670
rect 676054 559429 676106 559435
rect 676052 559394 676054 559403
rect 676106 559394 676108 559403
rect 676052 559329 676108 559338
rect 676054 559059 676106 559065
rect 676052 559024 676054 559033
rect 676106 559024 676108 559033
rect 676052 558959 676108 558968
rect 676246 558689 676298 558695
rect 676244 558654 676246 558663
rect 676298 558654 676300 558663
rect 676244 558589 676300 558598
rect 679796 557766 679852 557775
rect 679796 557701 679852 557710
rect 679810 557183 679838 557701
rect 679796 557174 679852 557183
rect 679796 557109 679852 557118
rect 685460 557174 685516 557183
rect 685460 557109 685516 557118
rect 679810 555883 679838 557109
rect 685474 556739 685502 557109
rect 685460 556730 685516 556739
rect 685460 556665 685516 556674
rect 679798 555877 679850 555883
rect 679798 555819 679850 555825
rect 675394 553460 675422 553890
rect 675298 553432 675422 553460
rect 675298 552923 675326 553432
rect 675490 553039 675518 553298
rect 675476 553030 675532 553039
rect 675476 552965 675532 552974
rect 675286 552917 675338 552923
rect 675286 552859 675338 552865
rect 675394 552299 675422 552706
rect 675380 552290 675436 552299
rect 675380 552225 675436 552234
rect 675202 552026 675408 552054
rect 675202 551707 675230 552026
rect 675188 551698 675244 551707
rect 675188 551633 675244 551642
rect 675284 550218 675340 550227
rect 675340 550176 675408 550204
rect 675284 550153 675340 550162
rect 675298 549629 675408 549657
rect 675298 549149 675326 549629
rect 675286 549143 675338 549149
rect 675286 549085 675338 549091
rect 675298 548992 675408 549020
rect 674902 547441 674954 547447
rect 674902 547383 674954 547389
rect 673846 543741 673898 543747
rect 673846 543683 673898 543689
rect 673654 517693 673706 517699
rect 673654 517635 673706 517641
rect 673654 478399 673706 478405
rect 673654 478341 673706 478347
rect 673366 472849 673418 472855
rect 673366 472791 673418 472797
rect 672790 472257 672842 472263
rect 672790 472199 672842 472205
rect 673666 440665 673694 478341
rect 673858 471671 673886 543683
rect 674914 542119 674942 547383
rect 674998 547367 675050 547373
rect 674998 547309 675050 547315
rect 675010 543969 675038 547309
rect 675298 547299 675326 548992
rect 675490 547965 675518 548340
rect 675478 547959 675530 547965
rect 675478 547901 675530 547907
rect 675286 547293 675338 547299
rect 675286 547235 675338 547241
rect 675394 545491 675422 545898
rect 675380 545482 675436 545491
rect 675380 545417 675436 545426
rect 675490 544931 675518 545306
rect 675478 544925 675530 544931
rect 675478 544867 675530 544873
rect 675394 544307 675422 544675
rect 675380 544298 675436 544307
rect 675380 544233 675436 544242
rect 674998 543963 675050 543969
rect 674998 543905 675050 543911
rect 675382 543963 675434 543969
rect 675382 543905 675434 543911
rect 675394 543456 675422 543905
rect 675490 543747 675518 544048
rect 675478 543741 675530 543747
rect 675478 543683 675530 543689
rect 675394 542341 675422 542835
rect 675190 542335 675242 542341
rect 675190 542277 675242 542283
rect 675382 542335 675434 542341
rect 675382 542277 675434 542283
rect 674902 542113 674954 542119
rect 674902 542055 674954 542061
rect 675202 538683 675230 542277
rect 675382 542113 675434 542119
rect 675382 542055 675434 542061
rect 675394 541639 675422 542055
rect 675778 540607 675806 541014
rect 675764 540598 675820 540607
rect 675764 540533 675820 540542
rect 675188 538674 675244 538683
rect 673942 538635 673994 538641
rect 675490 538641 675518 539164
rect 675188 538609 675244 538618
rect 675478 538635 675530 538641
rect 673942 538577 673994 538583
rect 675478 538577 675530 538583
rect 673954 476851 673982 538577
rect 676340 525206 676396 525215
rect 676340 525141 676396 525150
rect 676148 524762 676204 524771
rect 676148 524697 676204 524706
rect 676162 524211 676190 524697
rect 676244 524614 676300 524623
rect 676244 524549 676246 524558
rect 676298 524549 676300 524558
rect 676246 524517 676298 524523
rect 676354 524433 676382 525141
rect 676342 524427 676394 524433
rect 676342 524369 676394 524375
rect 676150 524205 676202 524211
rect 676150 524147 676202 524153
rect 676054 524057 676106 524063
rect 676052 524022 676054 524031
rect 676106 524022 676108 524031
rect 676052 523957 676108 523966
rect 676054 523909 676106 523915
rect 676054 523851 676106 523857
rect 676066 522921 676094 523851
rect 676532 523282 676588 523291
rect 676532 523217 676588 523226
rect 676052 522912 676108 522921
rect 676052 522847 676108 522856
rect 676244 521802 676300 521811
rect 676244 521737 676300 521746
rect 676258 521251 676286 521737
rect 676246 521245 676298 521251
rect 676246 521187 676298 521193
rect 676246 517693 676298 517699
rect 676244 517658 676246 517667
rect 676298 517658 676300 517667
rect 676244 517593 676300 517602
rect 676054 516953 676106 516959
rect 676052 516918 676054 516927
rect 676106 516918 676108 516927
rect 676052 516853 676108 516862
rect 676054 516509 676106 516515
rect 676052 516474 676054 516483
rect 676106 516474 676108 516483
rect 676052 516409 676108 516418
rect 676246 516213 676298 516219
rect 676244 516178 676246 516187
rect 676298 516178 676300 516187
rect 676244 516113 676300 516122
rect 676054 515473 676106 515479
rect 676052 515438 676054 515447
rect 676106 515438 676108 515447
rect 676052 515373 676108 515382
rect 676054 515029 676106 515035
rect 676052 514994 676054 515003
rect 676106 514994 676108 515003
rect 676052 514929 676108 514938
rect 676054 514511 676106 514517
rect 676052 514476 676054 514485
rect 676106 514476 676108 514485
rect 676052 514411 676108 514420
rect 676438 485355 676490 485361
rect 676438 485297 676490 485303
rect 676340 482434 676396 482443
rect 676340 482369 676396 482378
rect 676148 481842 676204 481851
rect 676148 481777 676204 481786
rect 676162 480995 676190 481777
rect 676244 481398 676300 481407
rect 676244 481333 676246 481342
rect 676298 481333 676300 481342
rect 676246 481301 676298 481307
rect 676354 481217 676382 482369
rect 676342 481211 676394 481217
rect 676342 481153 676394 481159
rect 676150 480989 676202 480995
rect 676150 480931 676202 480937
rect 676450 480371 676478 485297
rect 676546 481407 676574 523217
rect 676628 522246 676684 522255
rect 676628 522181 676684 522190
rect 676642 485361 676670 522181
rect 676724 521210 676780 521219
rect 676724 521145 676780 521154
rect 676630 485355 676682 485361
rect 676630 485297 676682 485303
rect 676738 485232 676766 521145
rect 679988 514106 680044 514115
rect 679988 514041 680044 514050
rect 680002 513227 680030 514041
rect 679796 513218 679852 513227
rect 679796 513153 679852 513162
rect 679988 513218 680044 513227
rect 679988 513153 680044 513162
rect 679810 512783 679838 513153
rect 679796 512774 679852 512783
rect 680002 512741 680030 513153
rect 679796 512709 679852 512718
rect 679990 512735 680042 512741
rect 679990 512677 680042 512683
rect 676642 485204 676766 485232
rect 676532 481398 676588 481407
rect 676532 481333 676588 481342
rect 676436 480362 676492 480371
rect 676436 480297 676492 480306
rect 676052 479696 676108 479705
rect 676052 479631 676108 479640
rect 676066 478701 676094 479631
rect 676450 479441 676478 480297
rect 676438 479435 676490 479441
rect 676438 479377 676490 479383
rect 676642 479335 676670 485204
rect 676724 480362 676780 480371
rect 676724 480297 676780 480306
rect 676628 479326 676684 479335
rect 676628 479261 676684 479270
rect 676642 479145 676670 479261
rect 676630 479139 676682 479145
rect 676630 479081 676682 479087
rect 675286 478695 675338 478701
rect 675286 478637 675338 478643
rect 676054 478695 676106 478701
rect 676054 478637 676106 478643
rect 673942 476845 673994 476851
rect 673942 476787 673994 476793
rect 673846 471665 673898 471671
rect 673846 471607 673898 471613
rect 673654 440659 673706 440665
rect 673654 440601 673706 440607
rect 675298 429195 675326 478637
rect 676244 478438 676300 478447
rect 676244 478373 676246 478382
rect 676298 478373 676300 478382
rect 676246 478341 676298 478347
rect 676054 476845 676106 476851
rect 676054 476787 676106 476793
rect 676066 475635 676094 476787
rect 676052 475626 676108 475635
rect 676052 475561 676108 475570
rect 676054 474699 676106 474705
rect 676052 474664 676054 474673
rect 676106 474664 676108 474673
rect 676052 474599 676108 474608
rect 676246 474329 676298 474335
rect 676244 474294 676246 474303
rect 676298 474294 676300 474303
rect 676244 474229 676300 474238
rect 676246 472849 676298 472855
rect 676244 472814 676246 472823
rect 676298 472814 676300 472823
rect 676244 472749 676300 472758
rect 676054 472257 676106 472263
rect 676052 472222 676054 472231
rect 676106 472222 676108 472231
rect 676052 472157 676108 472166
rect 676054 471665 676106 471671
rect 676052 471630 676054 471639
rect 676106 471630 676108 471639
rect 676052 471565 676108 471574
rect 675382 440659 675434 440665
rect 675382 440601 675434 440607
rect 673846 429189 673898 429195
rect 673846 429131 673898 429137
rect 675286 429189 675338 429195
rect 675286 429131 675338 429137
rect 673858 393897 673886 429131
rect 672598 393891 672650 393897
rect 672598 393833 672650 393839
rect 673846 393891 673898 393897
rect 673846 393833 673898 393839
rect 672500 278490 672556 278499
rect 672500 278425 672556 278434
rect 672404 276270 672460 276279
rect 672404 276205 672460 276214
rect 672610 271543 672638 393833
rect 675394 393231 675422 440601
rect 676148 396446 676204 396455
rect 676148 396381 676204 396390
rect 676162 394785 676190 396381
rect 676340 395854 676396 395863
rect 676340 395789 676396 395798
rect 676244 395410 676300 395419
rect 676244 395345 676300 395354
rect 676150 394779 676202 394785
rect 676150 394721 676202 394727
rect 676258 394711 676286 395345
rect 676246 394705 676298 394711
rect 676246 394647 676298 394653
rect 676354 394637 676382 395789
rect 676738 395419 676766 480297
rect 679796 470890 679852 470899
rect 679796 470825 679852 470834
rect 679810 470455 679838 470825
rect 679796 470446 679852 470455
rect 679796 470381 679852 470390
rect 685460 470446 685516 470455
rect 685460 470381 685516 470390
rect 679810 469525 679838 470381
rect 685474 470011 685502 470381
rect 685460 470002 685516 470011
rect 685460 469937 685516 469946
rect 679798 469519 679850 469525
rect 679798 469461 679850 469467
rect 676724 395410 676780 395419
rect 676724 395345 676780 395354
rect 676342 394631 676394 394637
rect 676342 394573 676394 394579
rect 676244 393930 676300 393939
rect 676244 393865 676246 393874
rect 676298 393865 676300 393874
rect 676246 393833 676298 393839
rect 675874 393231 675902 393259
rect 675382 393225 675434 393231
rect 675862 393225 675914 393231
rect 675382 393167 675434 393173
rect 675860 393190 675862 393199
rect 675914 393190 675916 393199
rect 675860 393125 675916 393134
rect 675190 391745 675242 391751
rect 675190 391687 675242 391693
rect 674038 389747 674090 389753
rect 674038 389689 674090 389695
rect 674050 372215 674078 389689
rect 674614 389155 674666 389161
rect 674614 389097 674666 389103
rect 674134 387083 674186 387089
rect 674134 387025 674186 387031
rect 674038 372209 674090 372215
rect 674038 372151 674090 372157
rect 674146 369181 674174 387025
rect 674518 386787 674570 386793
rect 674518 386729 674570 386735
rect 674422 386343 674474 386349
rect 674422 386285 674474 386291
rect 674230 386121 674282 386127
rect 674230 386063 674282 386069
rect 674242 371031 674270 386063
rect 674326 383161 674378 383167
rect 674326 383103 674378 383109
rect 674230 371025 674282 371031
rect 674230 370967 674282 370973
rect 674338 370365 674366 383103
rect 674434 375249 674462 386285
rect 674530 375693 674558 386729
rect 674626 376581 674654 389097
rect 674902 388933 674954 388939
rect 674902 388875 674954 388881
rect 674710 386047 674762 386053
rect 674710 385989 674762 385995
rect 674614 376575 674666 376581
rect 674614 376517 674666 376523
rect 674518 375687 674570 375693
rect 674518 375629 674570 375635
rect 674422 375243 674474 375249
rect 674422 375185 674474 375191
rect 674722 371475 674750 385989
rect 674806 385973 674858 385979
rect 674806 385915 674858 385921
rect 674818 374731 674846 385915
rect 674806 374725 674858 374731
rect 674806 374667 674858 374673
rect 674710 371469 674762 371475
rect 674710 371411 674762 371417
rect 674326 370359 674378 370365
rect 674326 370301 674378 370307
rect 674134 369175 674186 369181
rect 674134 369117 674186 369123
rect 674914 365481 674942 388875
rect 675202 388814 675230 391687
rect 675572 391118 675628 391127
rect 675572 391053 675628 391062
rect 675106 388786 675230 388814
rect 675286 388859 675338 388865
rect 675286 388801 675338 388807
rect 674998 379461 675050 379467
rect 674998 379403 675050 379409
rect 675010 371549 675038 379403
rect 675106 377858 675134 388786
rect 675298 384148 675326 388801
rect 675202 384120 675326 384148
rect 675202 378493 675230 384120
rect 675586 384000 675614 391053
rect 675298 383972 675614 384000
rect 675298 379560 675326 383972
rect 675874 383019 675902 393125
rect 676244 392006 676300 392015
rect 676244 391941 676300 391950
rect 676258 391751 676286 391941
rect 676246 391745 676298 391751
rect 676246 391687 676298 391693
rect 676244 390526 676300 390535
rect 676244 390461 676300 390470
rect 676052 390156 676108 390165
rect 676052 390091 676108 390100
rect 676066 389753 676094 390091
rect 676054 389747 676106 389753
rect 676054 389689 676106 389695
rect 676052 389638 676108 389647
rect 676052 389573 676108 389582
rect 676066 388939 676094 389573
rect 676258 389161 676286 390461
rect 676246 389155 676298 389161
rect 676246 389097 676298 389103
rect 676244 389046 676300 389055
rect 676244 388981 676300 388990
rect 676054 388933 676106 388939
rect 676054 388875 676106 388881
rect 676258 388865 676286 388981
rect 676246 388859 676298 388865
rect 676246 388801 676298 388807
rect 676052 388676 676108 388685
rect 676052 388611 676108 388620
rect 675956 388158 676012 388167
rect 675956 388093 676012 388102
rect 675970 386349 675998 388093
rect 676066 386793 676094 388611
rect 676244 387566 676300 387575
rect 676244 387501 676300 387510
rect 676258 387089 676286 387501
rect 676246 387083 676298 387089
rect 676246 387025 676298 387031
rect 676244 386974 676300 386983
rect 676244 386909 676300 386918
rect 676054 386787 676106 386793
rect 676054 386729 676106 386735
rect 676052 386678 676108 386687
rect 676052 386613 676108 386622
rect 675958 386343 676010 386349
rect 675958 386285 676010 386291
rect 675956 386234 676012 386243
rect 675956 386169 676012 386178
rect 675970 386053 675998 386169
rect 675958 386047 676010 386053
rect 675958 385989 676010 385995
rect 676066 385979 676094 386613
rect 676258 386127 676286 386909
rect 676246 386121 676298 386127
rect 676246 386063 676298 386069
rect 676054 385973 676106 385979
rect 676054 385915 676106 385921
rect 676244 385494 676300 385503
rect 676244 385429 676300 385438
rect 676258 383167 676286 385429
rect 679700 384902 679756 384911
rect 679700 384837 679756 384846
rect 679714 384467 679742 384837
rect 679700 384458 679756 384467
rect 679700 384393 679756 384402
rect 685460 384458 685516 384467
rect 685460 384393 685516 384402
rect 676246 383161 676298 383167
rect 676246 383103 676298 383109
rect 679714 383093 679742 384393
rect 685474 384023 685502 384393
rect 685460 384014 685516 384023
rect 685460 383949 685516 383958
rect 679702 383087 679754 383093
rect 679702 383029 679754 383035
rect 675862 383013 675914 383019
rect 675862 382955 675914 382961
rect 675298 379532 675422 379560
rect 675394 379102 675422 379532
rect 675490 379467 675518 379694
rect 675478 379461 675530 379467
rect 675478 379403 675530 379409
rect 675202 378465 675408 378493
rect 675106 377830 675408 377858
rect 675478 376575 675530 376581
rect 675478 376517 675530 376523
rect 675490 375994 675518 376517
rect 675382 375687 675434 375693
rect 675382 375629 675434 375635
rect 675394 375443 675422 375629
rect 675478 375243 675530 375249
rect 675478 375185 675530 375191
rect 675490 374810 675518 375185
rect 675382 374725 675434 374731
rect 675382 374667 675434 374673
rect 675394 374144 675422 374667
rect 675382 372209 675434 372215
rect 675382 372151 675434 372157
rect 675394 371671 675422 372151
rect 674998 371543 675050 371549
rect 674998 371485 675050 371491
rect 675382 371469 675434 371475
rect 675382 371411 675434 371417
rect 675394 371110 675422 371411
rect 675382 371025 675434 371031
rect 675382 370967 675434 370973
rect 675394 370475 675422 370967
rect 675478 370359 675530 370365
rect 675478 370301 675530 370307
rect 675490 369852 675518 370301
rect 675382 369175 675434 369181
rect 675382 369117 675434 369123
rect 675394 368626 675422 369117
rect 675476 367290 675532 367299
rect 675476 367225 675532 367234
rect 675490 366818 675518 367225
rect 674902 365475 674954 365481
rect 674902 365417 674954 365423
rect 675478 365475 675530 365481
rect 675478 365417 675530 365423
rect 675490 364968 675518 365417
rect 676244 351750 676300 351759
rect 676244 351685 676300 351694
rect 676054 351637 676106 351643
rect 676052 351602 676054 351611
rect 676106 351602 676108 351611
rect 676258 351569 676286 351685
rect 676052 351537 676108 351546
rect 676246 351563 676298 351569
rect 676246 351505 676298 351511
rect 676052 351010 676108 351019
rect 676052 350945 676108 350954
rect 676066 348535 676094 350945
rect 676054 348529 676106 348535
rect 676054 348471 676106 348477
rect 677012 346866 677068 346875
rect 677012 346801 677068 346810
rect 676052 346570 676108 346579
rect 676052 346505 676108 346514
rect 676066 345649 676094 346505
rect 674518 345643 674570 345649
rect 674518 345585 674570 345591
rect 676054 345643 676106 345649
rect 676054 345585 676106 345591
rect 674422 342831 674474 342837
rect 674422 342773 674474 342779
rect 674434 331737 674462 342773
rect 674530 335363 674558 345585
rect 676916 344794 676972 344803
rect 676916 344729 676972 344738
rect 676052 344646 676108 344655
rect 676052 344581 676108 344590
rect 676066 342763 676094 344581
rect 676244 343906 676300 343915
rect 676244 343841 676300 343850
rect 676258 342837 676286 343841
rect 676820 342870 676876 342879
rect 676246 342831 676298 342837
rect 676820 342805 676876 342814
rect 676246 342773 676298 342779
rect 674710 342757 674762 342763
rect 674710 342699 674762 342705
rect 676054 342757 676106 342763
rect 676054 342699 676106 342705
rect 674614 340019 674666 340025
rect 674614 339961 674666 339967
rect 674518 335357 674570 335363
rect 674518 335299 674570 335305
rect 674422 331731 674474 331737
rect 674422 331673 674474 331679
rect 674626 327149 674654 339961
rect 674722 334845 674750 342699
rect 676052 342574 676108 342583
rect 676052 342509 676108 342518
rect 675956 341612 676012 341621
rect 675956 341547 676012 341556
rect 674806 341203 674858 341209
rect 674806 341145 674858 341151
rect 674710 334839 674762 334845
rect 674710 334781 674762 334787
rect 674614 327143 674666 327149
rect 674614 327085 674666 327091
rect 674818 326853 674846 341145
rect 675970 340025 675998 341547
rect 676066 341209 676094 342509
rect 676244 341834 676300 341843
rect 676244 341769 676300 341778
rect 676054 341203 676106 341209
rect 676054 341145 676106 341151
rect 676052 341094 676108 341103
rect 676052 341029 676108 341038
rect 675958 340019 676010 340025
rect 675958 339961 676010 339967
rect 674998 339945 675050 339951
rect 674998 339887 675050 339893
rect 674902 339871 674954 339877
rect 674902 339813 674954 339819
rect 674806 326847 674858 326853
rect 674806 326789 674858 326795
rect 674914 326187 674942 339813
rect 675010 330479 675038 339887
rect 676066 339877 676094 341029
rect 676258 339951 676286 341769
rect 676246 339945 676298 339951
rect 676246 339887 676298 339893
rect 676054 339871 676106 339877
rect 676054 339813 676106 339819
rect 676834 339771 676862 342805
rect 676820 339762 676876 339771
rect 676820 339697 676876 339706
rect 676930 339327 676958 344729
rect 676916 339318 676972 339327
rect 676916 339253 676972 339262
rect 677026 338883 677054 346801
rect 679988 340354 680044 340363
rect 679988 340289 680044 340298
rect 680002 339771 680030 340289
rect 679796 339762 679852 339771
rect 679796 339697 679852 339706
rect 679988 339762 680044 339771
rect 679988 339697 680044 339706
rect 679810 339327 679838 339697
rect 679796 339318 679852 339327
rect 679796 339253 679852 339262
rect 677012 338874 677068 338883
rect 677012 338809 677068 338818
rect 680002 337065 680030 339697
rect 679990 337059 680042 337065
rect 679990 337001 680042 337007
rect 675106 335461 675408 335489
rect 674998 330473 675050 330479
rect 674998 330415 675050 330421
rect 675106 328333 675134 335461
rect 675190 335357 675242 335363
rect 675190 335299 675242 335305
rect 675202 334938 675230 335299
rect 675202 334910 675408 334938
rect 675382 334839 675434 334845
rect 675382 334781 675434 334787
rect 675394 334258 675422 334781
rect 675380 333990 675436 333999
rect 675380 333925 675436 333934
rect 675394 333635 675422 333925
rect 675476 332362 675532 332371
rect 675476 332297 675532 332306
rect 675490 331816 675518 332297
rect 675382 331731 675434 331737
rect 675382 331673 675434 331679
rect 675394 331224 675422 331673
rect 675380 331178 675436 331187
rect 675380 331113 675436 331122
rect 675394 330599 675422 331113
rect 675478 330473 675530 330479
rect 675478 330415 675530 330421
rect 675490 329966 675518 330415
rect 675094 328327 675146 328333
rect 675094 328269 675146 328275
rect 675380 327922 675436 327931
rect 675380 327857 675436 327866
rect 675394 327450 675422 327857
rect 675478 327143 675530 327149
rect 675478 327085 675530 327091
rect 675490 326932 675518 327085
rect 675382 326847 675434 326853
rect 675382 326789 675434 326795
rect 675394 326266 675422 326789
rect 674902 326181 674954 326187
rect 674902 326123 674954 326129
rect 675382 326181 675434 326187
rect 675382 326123 675434 326129
rect 675394 325631 675422 326123
rect 675668 324962 675724 324971
rect 675668 324897 675724 324906
rect 675682 324416 675710 324897
rect 675764 323038 675820 323047
rect 675764 322973 675820 322982
rect 675778 322595 675806 322973
rect 675764 321262 675820 321271
rect 675764 321197 675820 321206
rect 675778 320755 675806 321197
rect 679892 314010 679948 314019
rect 679892 313945 679948 313954
rect 676244 305722 676300 305731
rect 676244 305657 676300 305666
rect 676258 305393 676286 305657
rect 676246 305387 676298 305393
rect 676246 305329 676298 305335
rect 676244 305278 676300 305287
rect 676244 305213 676246 305222
rect 676298 305213 676300 305222
rect 676246 305181 676298 305187
rect 679906 304843 679934 313945
rect 676244 304834 676300 304843
rect 676244 304769 676300 304778
rect 679892 304834 679948 304843
rect 679892 304769 679948 304778
rect 676052 304094 676108 304103
rect 673366 304055 673418 304061
rect 676052 304029 676054 304038
rect 673366 303997 673418 304003
rect 676106 304029 676108 304038
rect 676054 303997 676106 304003
rect 672692 303502 672748 303511
rect 672692 303437 672748 303446
rect 672706 278055 672734 303437
rect 673174 303019 673226 303025
rect 673174 302961 673226 302967
rect 672884 302614 672940 302623
rect 672884 302549 672940 302558
rect 672692 278046 672748 278055
rect 672692 277981 672748 277990
rect 672898 277759 672926 302549
rect 672884 277750 672940 277759
rect 672884 277685 672940 277694
rect 673186 276131 673214 302961
rect 673270 301983 673322 301989
rect 673270 301925 673322 301931
rect 673282 276427 673310 301925
rect 673268 276418 673324 276427
rect 673268 276353 673324 276362
rect 673172 276122 673228 276131
rect 673172 276057 673228 276066
rect 673186 273721 673214 276057
rect 673174 273715 673226 273721
rect 673174 273657 673226 273663
rect 673282 273647 673310 276353
rect 673270 273641 673322 273647
rect 673270 273583 673322 273589
rect 672596 271534 672652 271543
rect 672596 271469 672652 271478
rect 670004 270646 670060 270655
rect 670004 270581 670060 270590
rect 672404 266946 672460 266955
rect 672404 266881 672460 266890
rect 669814 264983 669866 264989
rect 669814 264925 669866 264931
rect 669620 263542 669676 263551
rect 669620 263477 669676 263486
rect 672418 171051 672446 266881
rect 672596 266798 672652 266807
rect 672596 266733 672652 266742
rect 672404 171042 672460 171051
rect 672404 170977 672460 170986
rect 672610 169973 672638 266733
rect 673378 261659 673406 303997
rect 676052 303058 676108 303067
rect 676052 302993 676054 303002
rect 676106 302993 676108 303002
rect 676054 302961 676106 302967
rect 676258 302359 676286 304769
rect 676246 302353 676298 302359
rect 676246 302295 676298 302301
rect 676052 302022 676108 302031
rect 676052 301957 676054 301966
rect 676106 301957 676108 301966
rect 676054 301925 676106 301931
rect 676052 298618 676108 298627
rect 676052 298553 676108 298562
rect 676066 296735 676094 298553
rect 675190 296729 675242 296735
rect 675190 296671 675242 296677
rect 676054 296729 676106 296735
rect 676054 296671 676106 296677
rect 674998 293843 675050 293849
rect 674998 293785 675050 293791
rect 675010 286301 675038 293785
rect 675202 290445 675230 296671
rect 676052 296028 676108 296037
rect 676052 295963 676108 295972
rect 676066 293849 676094 295963
rect 679892 294326 679948 294335
rect 679892 294261 679948 294270
rect 679906 293891 679934 294261
rect 679700 293882 679756 293891
rect 676054 293843 676106 293849
rect 679700 293817 679756 293826
rect 679892 293882 679948 293891
rect 679892 293817 679948 293826
rect 676054 293785 676106 293791
rect 679714 293299 679742 293817
rect 679700 293290 679756 293299
rect 679700 293225 679756 293234
rect 679906 291777 679934 293817
rect 679894 291771 679946 291777
rect 679894 291713 679946 291719
rect 675490 291056 675518 291264
rect 675298 291028 675518 291056
rect 675190 290439 675242 290445
rect 675190 290381 675242 290387
rect 675298 289576 675326 291028
rect 675778 290635 675806 290746
rect 675764 290626 675820 290635
rect 675764 290561 675820 290570
rect 675382 290439 675434 290445
rect 675382 290381 675434 290387
rect 675394 290080 675422 290381
rect 675764 289738 675820 289747
rect 675764 289673 675820 289682
rect 675202 289548 675326 289576
rect 675202 288003 675230 289548
rect 675778 289414 675806 289673
rect 675190 287997 675242 288003
rect 675190 287939 675242 287945
rect 675764 287962 675820 287971
rect 675764 287897 675820 287906
rect 675778 287595 675806 287897
rect 675764 287518 675820 287527
rect 675764 287453 675820 287462
rect 675778 287046 675806 287453
rect 675380 286926 675436 286935
rect 675380 286861 675436 286870
rect 675394 286380 675422 286861
rect 674998 286295 675050 286301
rect 674998 286237 675050 286243
rect 675382 286295 675434 286301
rect 675382 286237 675434 286243
rect 675394 285755 675422 286237
rect 675380 283818 675436 283827
rect 675380 283753 675436 283762
rect 675394 283272 675422 283753
rect 675572 282930 675628 282939
rect 675572 282865 675628 282874
rect 675586 282719 675614 282865
rect 675682 281903 675710 282088
rect 675668 281894 675724 281903
rect 675668 281829 675724 281838
rect 675572 281746 675628 281755
rect 675572 281681 675628 281690
rect 675586 281422 675614 281681
rect 675380 280710 675436 280719
rect 675380 280645 675436 280654
rect 675394 280238 675422 280645
rect 675380 278934 675436 278943
rect 675380 278869 675436 278878
rect 675394 278388 675422 278869
rect 675380 277010 675436 277019
rect 675380 276945 675436 276954
rect 675394 276538 675422 276945
rect 679892 275086 679948 275095
rect 679892 275021 679948 275030
rect 679702 273715 679754 273721
rect 679702 273657 679754 273663
rect 676244 262802 676300 262811
rect 676244 262737 676300 262746
rect 676052 262506 676108 262515
rect 676052 262441 676054 262450
rect 676106 262441 676108 262450
rect 676054 262409 676106 262415
rect 676258 262325 676286 262737
rect 676246 262319 676298 262325
rect 676246 262261 676298 262267
rect 676244 261766 676300 261775
rect 676244 261701 676300 261710
rect 673366 261653 673418 261659
rect 676054 261653 676106 261659
rect 673366 261595 673418 261601
rect 676052 261618 676054 261627
rect 676106 261618 676108 261627
rect 676052 261553 676108 261562
rect 676258 259513 676286 261701
rect 679714 260887 679742 273657
rect 679798 273641 679850 273647
rect 679798 273583 679850 273589
rect 679700 260878 679756 260887
rect 679700 260813 679756 260822
rect 679810 259851 679838 273583
rect 679796 259842 679852 259851
rect 679796 259777 679852 259786
rect 676246 259507 676298 259513
rect 676246 259449 676298 259455
rect 679700 258806 679756 258815
rect 679906 258792 679934 275021
rect 679756 258764 679934 258792
rect 679700 258741 679756 258750
rect 676052 258658 676108 258667
rect 676052 258593 676108 258602
rect 675764 257474 675820 257483
rect 675764 257409 675820 257418
rect 674710 256991 674762 256997
rect 674710 256933 674762 256939
rect 674518 250775 674570 250781
rect 674518 250717 674570 250723
rect 674530 237609 674558 250717
rect 674614 250701 674666 250707
rect 674614 250643 674666 250649
rect 674626 238645 674654 250643
rect 674722 245453 674750 256933
rect 675094 253661 675146 253667
rect 675094 253603 675146 253609
rect 674902 253587 674954 253593
rect 674902 253529 674954 253535
rect 674710 245447 674762 245453
rect 674710 245389 674762 245395
rect 674914 242937 674942 253529
rect 674998 250627 675050 250633
rect 674998 250569 675050 250575
rect 674902 242931 674954 242937
rect 674902 242873 674954 242879
rect 675010 241827 675038 250569
rect 675106 246804 675134 253603
rect 675286 253513 675338 253519
rect 675286 253455 675338 253461
rect 675106 246776 675230 246804
rect 675094 246705 675146 246711
rect 675094 246647 675146 246653
rect 675106 241901 675134 246647
rect 675202 242345 675230 246776
rect 675298 245694 675326 253455
rect 675778 247155 675806 257409
rect 676066 256997 676094 258593
rect 676054 256991 676106 256997
rect 676054 256933 676106 256939
rect 676916 255846 676972 255855
rect 676916 255781 676972 255790
rect 676052 255624 676108 255633
rect 676052 255559 676108 255568
rect 675956 255106 676012 255115
rect 675956 255041 676012 255050
rect 675970 253593 675998 255041
rect 675958 253587 676010 253593
rect 675958 253529 676010 253535
rect 676066 253519 676094 255559
rect 676244 254366 676300 254375
rect 676244 254301 676300 254310
rect 676258 253667 676286 254301
rect 676820 253922 676876 253931
rect 676820 253857 676876 253866
rect 676246 253661 676298 253667
rect 676246 253603 676298 253609
rect 676054 253513 676106 253519
rect 676054 253455 676106 253461
rect 676052 253034 676108 253043
rect 676052 252969 676108 252978
rect 675956 252072 676012 252081
rect 675956 252007 676012 252016
rect 675970 250781 675998 252007
rect 675958 250775 676010 250781
rect 675958 250717 676010 250723
rect 676066 250633 676094 252969
rect 676244 252442 676300 252451
rect 676244 252377 676300 252386
rect 676258 250707 676286 252377
rect 676246 250701 676298 250707
rect 676246 250643 676298 250649
rect 676054 250627 676106 250633
rect 676054 250569 676106 250575
rect 676834 247863 676862 253857
rect 676930 248011 676958 255781
rect 679714 249343 679742 258741
rect 679988 251702 680044 251711
rect 679988 251637 680044 251646
rect 680002 250823 680030 251637
rect 679796 250814 679852 250823
rect 679796 250749 679852 250758
rect 679988 250814 680044 250823
rect 679988 250749 680044 250758
rect 679810 250379 679838 250749
rect 679796 250370 679852 250379
rect 679796 250305 679852 250314
rect 679700 249334 679756 249343
rect 679700 249269 679756 249278
rect 680002 249153 680030 250749
rect 679990 249147 680042 249153
rect 679990 249089 680042 249095
rect 676916 248002 676972 248011
rect 676916 247937 676972 247946
rect 676820 247854 676876 247863
rect 676820 247789 676876 247798
rect 675766 247149 675818 247155
rect 675766 247091 675818 247097
rect 675490 246711 675518 246864
rect 675478 246705 675530 246711
rect 675478 246647 675530 246653
rect 675766 246631 675818 246637
rect 675766 246573 675818 246579
rect 675778 246346 675806 246573
rect 675298 245666 675408 245694
rect 675382 245447 675434 245453
rect 675382 245389 675434 245395
rect 675394 245014 675422 245389
rect 675668 243710 675724 243719
rect 675668 243645 675724 243654
rect 675682 243195 675710 243645
rect 675382 242931 675434 242937
rect 675382 242873 675434 242879
rect 675394 242646 675422 242873
rect 675190 242339 675242 242345
rect 675190 242281 675242 242287
rect 675382 242339 675434 242345
rect 675382 242281 675434 242287
rect 675394 241980 675422 242281
rect 675094 241895 675146 241901
rect 675094 241837 675146 241843
rect 674998 241821 675050 241827
rect 674998 241763 675050 241769
rect 675382 241821 675434 241827
rect 675382 241763 675434 241769
rect 675394 241355 675422 241763
rect 675380 239122 675436 239131
rect 675380 239057 675436 239066
rect 675394 238872 675422 239057
rect 674614 238639 674666 238645
rect 674614 238581 674666 238587
rect 675382 238639 675434 238645
rect 675382 238581 675434 238587
rect 675394 238319 675422 238581
rect 675764 238086 675820 238095
rect 675764 238021 675820 238030
rect 675778 237688 675806 238021
rect 674518 237603 674570 237609
rect 674518 237545 674570 237551
rect 675382 237603 675434 237609
rect 675382 237545 675434 237551
rect 675394 237022 675422 237545
rect 675764 236014 675820 236023
rect 675764 235949 675820 235958
rect 675778 235838 675806 235949
rect 675380 234534 675436 234543
rect 675380 234469 675436 234478
rect 675394 233988 675422 234469
rect 675764 232610 675820 232619
rect 675764 232545 675820 232554
rect 675778 232138 675806 232545
rect 676244 219734 676300 219743
rect 676244 219669 676300 219678
rect 676258 219405 676286 219669
rect 676246 219399 676298 219405
rect 676246 219341 676298 219347
rect 676244 219290 676300 219299
rect 676244 219225 676246 219234
rect 676298 219225 676300 219234
rect 676246 219193 676298 219199
rect 676054 219103 676106 219109
rect 676054 219045 676106 219051
rect 676066 219003 676094 219045
rect 676052 218994 676108 219003
rect 676052 218929 676108 218938
rect 676244 215442 676300 215451
rect 676244 215377 676300 215386
rect 675572 214554 675628 214563
rect 675572 214489 675628 214498
rect 674710 213257 674762 213263
rect 674710 213199 674762 213205
rect 674038 207485 674090 207491
rect 674038 207427 674090 207433
rect 674050 194393 674078 207427
rect 674614 205487 674666 205493
rect 674614 205429 674666 205435
rect 674626 198241 674654 205429
rect 674722 201423 674750 213199
rect 675190 213183 675242 213189
rect 675190 213125 675242 213131
rect 674806 210371 674858 210377
rect 674806 210313 674858 210319
rect 674818 205493 674846 210313
rect 674902 210297 674954 210303
rect 674902 210239 674954 210245
rect 674806 205487 674858 205493
rect 674806 205429 674858 205435
rect 674914 205364 674942 210239
rect 674998 207411 675050 207417
rect 674998 207353 675050 207359
rect 674818 205336 674942 205364
rect 674710 201417 674762 201423
rect 674710 201359 674762 201365
rect 674818 198611 674846 205336
rect 675010 205216 675038 207353
rect 674914 205188 675038 205216
rect 674806 198605 674858 198611
rect 674806 198547 674858 198553
rect 674614 198235 674666 198241
rect 674614 198177 674666 198183
rect 674914 197723 674942 205188
rect 675202 205068 675230 213125
rect 675284 212630 675340 212639
rect 675284 212565 675340 212574
rect 675010 205040 675230 205068
rect 675010 199573 675038 205040
rect 675298 204920 675326 212565
rect 675202 204892 675326 204920
rect 675094 202453 675146 202459
rect 675094 202395 675146 202401
rect 674998 199567 675050 199573
rect 674998 199509 675050 199515
rect 675106 198685 675134 202395
rect 675202 201516 675230 204892
rect 675586 204772 675614 214489
rect 676052 214110 676108 214119
rect 676052 214045 676108 214054
rect 676066 213189 676094 214045
rect 676258 213263 676286 215377
rect 676246 213257 676298 213263
rect 676246 213199 676298 213205
rect 676054 213183 676106 213189
rect 676054 213125 676106 213131
rect 676916 212778 676972 212787
rect 676916 212713 676972 212722
rect 676244 211890 676300 211899
rect 676244 211825 676300 211834
rect 676052 211520 676108 211529
rect 676052 211455 676108 211464
rect 676066 210377 676094 211455
rect 676054 210371 676106 210377
rect 676054 210313 676106 210319
rect 676258 210303 676286 211825
rect 676820 210854 676876 210863
rect 676820 210789 676876 210798
rect 676246 210297 676298 210303
rect 676246 210239 676298 210245
rect 676052 210040 676108 210049
rect 676052 209975 676108 209984
rect 675956 209670 676012 209679
rect 675956 209605 676012 209614
rect 675970 207491 675998 209605
rect 675958 207485 676010 207491
rect 675958 207427 676010 207433
rect 676066 207417 676094 209975
rect 676054 207411 676106 207417
rect 676054 207353 676106 207359
rect 675298 204744 675614 204772
rect 675298 202137 675326 204744
rect 676834 204647 676862 210789
rect 676930 204795 676958 212713
rect 679892 208338 679948 208347
rect 679892 208273 679948 208282
rect 679906 207903 679934 208273
rect 679892 207894 679948 207903
rect 679892 207829 679948 207838
rect 679796 207746 679852 207755
rect 679796 207681 679852 207690
rect 679810 207311 679838 207681
rect 679906 207565 679934 207829
rect 679894 207559 679946 207565
rect 679894 207501 679946 207507
rect 679796 207302 679852 207311
rect 679796 207237 679852 207246
rect 676916 204786 676972 204795
rect 676916 204721 676972 204730
rect 676820 204638 676876 204647
rect 676820 204573 676876 204582
rect 675394 202459 675422 202686
rect 675382 202453 675434 202459
rect 675382 202395 675434 202401
rect 675298 202109 675408 202137
rect 675202 201488 675326 201516
rect 675190 201417 675242 201423
rect 675190 201359 675242 201365
rect 675298 201368 675326 201488
rect 675394 201368 675422 201502
rect 675202 200850 675230 201359
rect 675298 201340 675422 201368
rect 675202 200822 675408 200850
rect 675478 199567 675530 199573
rect 675478 199509 675530 199515
rect 675490 198986 675518 199509
rect 675094 198679 675146 198685
rect 675094 198621 675146 198627
rect 675478 198605 675530 198611
rect 675478 198547 675530 198553
rect 675490 198468 675518 198547
rect 675382 198235 675434 198241
rect 675382 198177 675434 198183
rect 675394 197802 675422 198177
rect 674902 197717 674954 197723
rect 674902 197659 674954 197665
rect 675382 197717 675434 197723
rect 675382 197659 675434 197665
rect 675394 197136 675422 197659
rect 675476 195166 675532 195175
rect 675476 195101 675532 195110
rect 675490 194694 675518 195101
rect 674038 194387 674090 194393
rect 674038 194329 674090 194335
rect 675382 194387 675434 194393
rect 675382 194329 675434 194335
rect 675394 194102 675422 194329
rect 675380 193982 675436 193991
rect 675380 193917 675436 193926
rect 675394 193475 675422 193917
rect 675476 193094 675532 193103
rect 675476 193029 675532 193038
rect 675490 192844 675518 193029
rect 675764 192206 675820 192215
rect 675764 192141 675820 192150
rect 675778 191660 675806 192141
rect 675476 189986 675532 189995
rect 675476 189921 675532 189930
rect 675490 189810 675518 189921
rect 675764 188506 675820 188515
rect 675764 188441 675820 188450
rect 675778 187960 675806 188441
rect 676148 173854 676204 173863
rect 676148 173789 676204 173798
rect 676052 173558 676108 173567
rect 676052 173493 676108 173502
rect 676066 172859 676094 173493
rect 676162 173081 676190 173789
rect 676244 173262 676300 173271
rect 676244 173197 676246 173206
rect 676298 173197 676300 173206
rect 676246 173165 676298 173171
rect 676150 173075 676202 173081
rect 676150 173017 676202 173023
rect 676054 172853 676106 172859
rect 676054 172795 676106 172801
rect 676052 170006 676108 170015
rect 672598 169967 672650 169973
rect 672598 169909 672650 169915
rect 673846 169967 673898 169973
rect 676052 169941 676054 169950
rect 673846 169909 673898 169915
rect 676106 169941 676108 169950
rect 676054 169909 676106 169915
rect 673462 169079 673514 169085
rect 673462 169021 673514 169027
rect 673474 146145 673502 169021
rect 673462 146139 673514 146145
rect 673462 146081 673514 146087
rect 673858 126387 673886 169909
rect 676052 169118 676108 169127
rect 676052 169053 676054 169062
rect 676106 169053 676108 169062
rect 676054 169021 676106 169027
rect 676052 164086 676108 164095
rect 676052 164021 676108 164030
rect 676066 161315 676094 164021
rect 676244 162310 676300 162319
rect 676244 162245 676300 162254
rect 676148 161866 676204 161875
rect 676148 161801 676204 161810
rect 676162 161389 676190 161801
rect 676258 161611 676286 162245
rect 676246 161605 676298 161611
rect 676246 161547 676298 161553
rect 676246 161457 676298 161463
rect 676244 161422 676246 161431
rect 676298 161422 676300 161431
rect 676150 161383 676202 161389
rect 676244 161357 676300 161366
rect 676150 161325 676202 161331
rect 674134 161309 674186 161315
rect 674134 161251 674186 161257
rect 676054 161309 676106 161315
rect 676054 161251 676106 161257
rect 674146 153397 674174 161251
rect 675106 158461 675408 158489
rect 675106 155543 675134 158461
rect 675764 158166 675820 158175
rect 675764 158101 675820 158110
rect 675778 157916 675806 158101
rect 675764 157722 675820 157731
rect 675764 157657 675820 157666
rect 675778 157279 675806 157657
rect 675764 156982 675820 156991
rect 675764 156917 675820 156926
rect 675778 156658 675806 156917
rect 675094 155537 675146 155543
rect 675094 155479 675146 155485
rect 675476 155206 675532 155215
rect 675476 155141 675532 155150
rect 675490 154808 675518 155141
rect 675380 154466 675436 154475
rect 675380 154401 675436 154410
rect 675394 154216 675422 154401
rect 675764 153874 675820 153883
rect 675764 153809 675820 153818
rect 675778 153624 675806 153809
rect 674134 153391 674186 153397
rect 674134 153333 674186 153339
rect 675382 153391 675434 153397
rect 675382 153333 675434 153339
rect 675394 152958 675422 153333
rect 675188 152690 675244 152699
rect 675188 152625 675244 152634
rect 675202 149179 675230 152625
rect 675380 150914 675436 150923
rect 675380 150849 675436 150858
rect 675394 150471 675422 150849
rect 675476 150322 675532 150331
rect 675476 150257 675532 150266
rect 675490 149924 675518 150257
rect 675380 149582 675436 149591
rect 675380 149517 675436 149526
rect 675394 149258 675422 149517
rect 675190 149173 675242 149179
rect 675190 149115 675242 149121
rect 675382 149173 675434 149179
rect 675382 149115 675434 149121
rect 675394 148631 675422 149115
rect 675380 147954 675436 147963
rect 675380 147889 675436 147898
rect 675394 147408 675422 147889
rect 675382 146139 675434 146145
rect 675382 146081 675434 146087
rect 675394 145595 675422 146081
rect 675476 143958 675532 143967
rect 675476 143893 675532 143902
rect 675490 143782 675518 143893
rect 676246 129637 676298 129643
rect 676244 129602 676246 129611
rect 676298 129602 676300 129611
rect 676244 129537 676300 129546
rect 676340 129158 676396 129167
rect 676340 129093 676396 129102
rect 676244 128566 676300 128575
rect 676244 128501 676300 128510
rect 676148 127530 676204 127539
rect 676148 127465 676204 127474
rect 676052 126938 676108 126947
rect 676052 126873 676108 126882
rect 676066 126757 676094 126873
rect 676162 126831 676190 127465
rect 676258 127127 676286 128501
rect 676246 127121 676298 127127
rect 676246 127063 676298 127069
rect 676354 126979 676382 129093
rect 676342 126973 676394 126979
rect 676342 126915 676394 126921
rect 676150 126825 676202 126831
rect 676150 126767 676202 126773
rect 676054 126751 676106 126757
rect 676054 126693 676106 126699
rect 673846 126381 673898 126387
rect 676054 126381 676106 126387
rect 673846 126323 673898 126329
rect 676052 126346 676054 126355
rect 676106 126346 676108 126355
rect 676052 126281 676108 126290
rect 676244 125606 676300 125615
rect 676244 125541 676300 125550
rect 676052 124274 676108 124283
rect 676052 124209 676108 124218
rect 676066 124019 676094 124209
rect 675190 124013 675242 124019
rect 675190 123955 675242 123961
rect 676054 124013 676106 124019
rect 676054 123955 676106 123961
rect 674614 121201 674666 121207
rect 674614 121143 674666 121149
rect 674326 119943 674378 119949
rect 674326 119885 674378 119891
rect 668180 106366 668236 106375
rect 668180 106301 668236 106310
rect 665588 105330 665644 105339
rect 674338 105297 674366 119885
rect 674422 118241 674474 118247
rect 674422 118183 674474 118189
rect 665588 105265 665644 105274
rect 674326 105291 674378 105297
rect 665300 105182 665356 105191
rect 665300 105117 665356 105126
rect 665602 104557 665630 105265
rect 674326 105233 674378 105239
rect 674434 104779 674462 118183
rect 674626 110329 674654 121143
rect 674710 121127 674762 121133
rect 674710 121069 674762 121075
rect 674614 110323 674666 110329
rect 674614 110265 674666 110271
rect 674722 109737 674750 121069
rect 674998 121053 675050 121059
rect 674998 120995 675050 121001
rect 674806 118611 674858 118617
rect 674806 118553 674858 118559
rect 674710 109731 674762 109737
rect 674710 109673 674762 109679
rect 674818 106574 674846 118553
rect 674902 118167 674954 118173
rect 674902 118109 674954 118115
rect 674914 109071 674942 118109
rect 675010 112893 675038 120995
rect 675202 113530 675230 123955
rect 676258 123945 676286 125541
rect 676820 124570 676876 124579
rect 676820 124505 676876 124514
rect 676246 123939 676298 123945
rect 676246 123881 676298 123887
rect 676052 122424 676108 122433
rect 676052 122359 676108 122368
rect 675956 121906 676012 121915
rect 675956 121841 676012 121850
rect 675970 121207 675998 121841
rect 675958 121201 676010 121207
rect 675958 121143 676010 121149
rect 676066 121059 676094 122359
rect 676244 121166 676300 121175
rect 676244 121101 676246 121110
rect 676298 121101 676300 121110
rect 676246 121069 676298 121075
rect 676054 121053 676106 121059
rect 676054 120995 676106 121001
rect 676052 120426 676108 120435
rect 676052 120361 676108 120370
rect 676066 119949 676094 120361
rect 676054 119943 676106 119949
rect 676054 119885 676106 119891
rect 676052 119834 676108 119843
rect 676052 119769 676108 119778
rect 675956 118872 676012 118881
rect 675956 118807 676012 118816
rect 675970 118247 675998 118807
rect 675958 118241 676010 118247
rect 675958 118183 676010 118189
rect 676066 118173 676094 119769
rect 676244 119242 676300 119251
rect 676244 119177 676300 119186
rect 676258 118617 676286 119177
rect 676246 118611 676298 118617
rect 676246 118553 676298 118559
rect 676244 118502 676300 118511
rect 676244 118437 676246 118446
rect 676298 118437 676300 118446
rect 676246 118405 676298 118411
rect 676054 118167 676106 118173
rect 676054 118109 676106 118115
rect 676148 117762 676204 117771
rect 676148 117697 676204 117706
rect 676162 115361 676190 117697
rect 676244 117170 676300 117179
rect 676244 117105 676300 117114
rect 676258 115509 676286 117105
rect 676834 115699 676862 124505
rect 679700 122646 679756 122655
rect 679700 122581 679756 122590
rect 676820 115690 676876 115699
rect 676820 115625 676876 115634
rect 676246 115503 676298 115509
rect 676246 115445 676298 115451
rect 676150 115355 676202 115361
rect 676150 115297 676202 115303
rect 679714 115255 679742 122581
rect 679700 115246 679756 115255
rect 679700 115181 679756 115190
rect 675382 114689 675434 114695
rect 675382 114631 675434 114637
rect 675394 114075 675422 114631
rect 675202 113502 675408 113530
rect 675010 112865 675408 112893
rect 675586 112147 675614 112258
rect 675572 112138 675628 112147
rect 675572 112073 675628 112082
rect 675764 110954 675820 110963
rect 675764 110889 675820 110898
rect 675778 110408 675806 110889
rect 675382 110323 675434 110329
rect 675382 110265 675434 110271
rect 675394 109816 675422 110265
rect 675478 109731 675530 109737
rect 675478 109673 675530 109679
rect 675490 109224 675518 109673
rect 674902 109065 674954 109071
rect 674902 109007 674954 109013
rect 675382 109065 675434 109071
rect 675382 109007 675434 109013
rect 675394 108558 675422 109007
rect 674818 106546 674942 106574
rect 674914 105963 674942 106546
rect 675380 106514 675436 106523
rect 675380 106449 675436 106458
rect 675394 106071 675422 106449
rect 674902 105957 674954 105963
rect 674902 105899 674954 105905
rect 675478 105957 675530 105963
rect 675478 105899 675530 105905
rect 675490 105524 675518 105899
rect 675382 105291 675434 105297
rect 675382 105233 675434 105239
rect 675394 104858 675422 105233
rect 674422 104773 674474 104779
rect 674422 104715 674474 104721
rect 675382 104773 675434 104779
rect 675382 104715 675434 104721
rect 654070 104551 654122 104557
rect 654070 104493 654122 104499
rect 665590 104551 665642 104557
rect 665590 104493 665642 104499
rect 647924 104146 647980 104155
rect 647924 104081 647980 104090
rect 647938 103817 647966 104081
rect 647926 103811 647978 103817
rect 647926 103753 647978 103759
rect 652438 102109 652490 102115
rect 652438 102051 652490 102057
rect 647924 99706 647980 99715
rect 647924 99641 647980 99650
rect 647938 97971 647966 99641
rect 647926 97965 647978 97971
rect 647926 97907 647978 97913
rect 647828 94082 647884 94091
rect 647828 94017 647884 94026
rect 647732 92750 647788 92759
rect 647732 92685 647788 92694
rect 647158 87087 647210 87093
rect 647158 87029 647210 87035
rect 647746 81543 647774 92685
rect 647842 81617 647870 94017
rect 650902 87531 650954 87537
rect 650902 87473 650954 87479
rect 647926 87309 647978 87315
rect 647926 87251 647978 87257
rect 647938 87135 647966 87251
rect 647924 87126 647980 87135
rect 647924 87061 647980 87070
rect 650914 86247 650942 87473
rect 650900 86238 650956 86247
rect 650900 86173 650956 86182
rect 652340 85350 652396 85359
rect 652340 85285 652396 85294
rect 651764 84314 651820 84323
rect 651764 84249 651820 84258
rect 651778 83615 651806 84249
rect 651766 83609 651818 83615
rect 651766 83551 651818 83557
rect 652244 83426 652300 83435
rect 652244 83361 652300 83370
rect 647924 82686 647980 82695
rect 647924 82621 647980 82630
rect 647938 81913 647966 82621
rect 647926 81907 647978 81913
rect 647926 81849 647978 81855
rect 647830 81611 647882 81617
rect 647830 81553 647882 81559
rect 647734 81537 647786 81543
rect 647734 81479 647786 81485
rect 647924 81058 647980 81067
rect 647924 80993 647980 81002
rect 647938 80803 647966 80993
rect 647926 80797 647978 80803
rect 647926 80739 647978 80745
rect 647926 77541 647978 77547
rect 647924 77506 647926 77515
rect 647978 77506 647980 77515
rect 647924 77441 647980 77450
rect 647158 74951 647210 74957
rect 647158 74893 647210 74899
rect 647060 71882 647116 71891
rect 647060 71817 647116 71826
rect 646868 68626 646924 68635
rect 646868 68561 646924 68570
rect 647170 60347 647198 74893
rect 647924 73658 647980 73667
rect 647924 73593 647980 73602
rect 647938 72145 647966 73593
rect 647926 72139 647978 72145
rect 647926 72081 647978 72087
rect 647924 69662 647980 69671
rect 647924 69597 647926 69606
rect 647978 69597 647980 69606
rect 647926 69565 647978 69571
rect 647924 64186 647980 64195
rect 647924 64121 647980 64130
rect 647938 63487 647966 64121
rect 647926 63481 647978 63487
rect 647926 63423 647978 63429
rect 647924 62262 647980 62271
rect 647924 62197 647980 62206
rect 647938 61045 647966 62197
rect 647926 61039 647978 61045
rect 647926 60981 647978 60987
rect 647156 60338 647212 60347
rect 647156 60273 647212 60282
rect 652258 59121 652286 83361
rect 652354 66225 652382 85285
rect 652450 82695 652478 102051
rect 654082 96565 654110 104493
rect 675394 104231 675422 104715
rect 657526 103885 657578 103891
rect 657526 103827 657578 103833
rect 654070 96559 654122 96565
rect 654070 96501 654122 96507
rect 653686 95967 653738 95973
rect 653686 95909 653738 95915
rect 653698 86987 653726 95909
rect 657538 88000 657566 103827
rect 661174 103811 661226 103817
rect 661174 103753 661226 103759
rect 660694 92415 660746 92421
rect 660694 92357 660746 92363
rect 659830 92267 659882 92273
rect 659830 92209 659882 92215
rect 658870 92193 658922 92199
rect 658870 92135 658922 92141
rect 657538 87972 657792 88000
rect 658882 87986 658910 92135
rect 659348 90826 659404 90835
rect 659348 90761 659404 90770
rect 659362 88000 659390 90761
rect 659842 88000 659870 92209
rect 659362 87972 659616 88000
rect 659842 87972 660144 88000
rect 660706 87986 660734 92357
rect 661186 88000 661214 103753
rect 675668 103554 675724 103563
rect 675668 103489 675724 103498
rect 675682 103008 675710 103489
rect 675764 101630 675820 101639
rect 675764 101565 675820 101574
rect 675778 101195 675806 101565
rect 675764 99854 675820 99863
rect 675764 99789 675820 99798
rect 675778 99382 675806 99789
rect 662518 97965 662570 97971
rect 662518 97907 662570 97913
rect 661750 92341 661802 92347
rect 661750 92283 661802 92289
rect 661762 88000 661790 92283
rect 661186 87972 661440 88000
rect 661762 87972 662016 88000
rect 662530 87986 662558 97907
rect 663094 92711 663146 92717
rect 663094 92653 663146 92659
rect 663106 87986 663134 92653
rect 658006 87309 658058 87315
rect 658058 87257 658320 87260
rect 658006 87251 658320 87257
rect 658018 87232 658320 87251
rect 663286 87087 663338 87093
rect 663286 87029 663338 87035
rect 653684 86978 653740 86987
rect 653684 86913 653740 86922
rect 663298 86395 663326 87029
rect 663284 86386 663340 86395
rect 663284 86321 663340 86330
rect 663284 84758 663340 84767
rect 663202 84716 663284 84744
rect 657046 84053 657098 84059
rect 657046 83995 657098 84001
rect 652436 82686 652492 82695
rect 652436 82621 652492 82630
rect 657058 81691 657086 83995
rect 657046 81685 657098 81691
rect 657046 81627 657098 81633
rect 658582 81685 658634 81691
rect 662420 81650 662476 81659
rect 658634 81633 658896 81636
rect 658582 81627 658896 81633
rect 658594 81608 658896 81627
rect 662420 81585 662422 81594
rect 662474 81585 662476 81594
rect 662422 81553 662474 81559
rect 656962 81016 657216 81044
rect 657538 81016 657792 81044
rect 656962 77547 656990 81016
rect 656950 77541 657002 77547
rect 656950 77483 657002 77489
rect 657538 76141 657566 81016
rect 658306 77769 658334 81030
rect 659602 80748 659630 81030
rect 659554 80729 659630 80748
rect 659446 80723 659498 80729
rect 659446 80665 659498 80671
rect 659542 80723 659630 80729
rect 659594 80720 659630 80723
rect 659542 80665 659594 80671
rect 658294 77763 658346 77769
rect 658294 77705 658346 77711
rect 659458 77695 659486 80665
rect 659446 77689 659498 77695
rect 659446 77631 659498 77637
rect 657526 76135 657578 76141
rect 657526 76077 657578 76083
rect 660130 74957 660158 81030
rect 660118 74951 660170 74957
rect 660118 74893 660170 74899
rect 660706 72145 660734 81030
rect 661440 81016 661502 81044
rect 660694 72139 660746 72145
rect 660694 72081 660746 72087
rect 661474 69629 661502 81016
rect 661762 81016 662016 81044
rect 661762 77621 661790 81016
rect 662530 80803 662558 81030
rect 662518 80797 662570 80803
rect 662518 80739 662570 80745
rect 661750 77615 661802 77621
rect 661750 77557 661802 77563
rect 661462 69623 661514 69629
rect 661462 69565 661514 69571
rect 652342 66219 652394 66225
rect 652342 66161 652394 66167
rect 663202 63487 663230 84716
rect 663284 84693 663340 84702
rect 663380 84018 663436 84027
rect 663380 83953 663436 83962
rect 663284 82094 663340 82103
rect 663284 82029 663340 82038
rect 663298 81913 663326 82029
rect 663286 81907 663338 81913
rect 663286 81849 663338 81855
rect 663190 63481 663242 63487
rect 663190 63423 663242 63429
rect 663394 61045 663422 83953
rect 663476 82834 663532 82843
rect 663476 82769 663532 82778
rect 663490 81543 663518 82769
rect 663478 81537 663530 81543
rect 663478 81479 663530 81485
rect 663382 61039 663434 61045
rect 663382 60981 663434 60987
rect 652246 59115 652298 59121
rect 652246 59057 652298 59063
rect 646772 57082 646828 57091
rect 646772 57017 646828 57026
rect 646484 54714 646540 54723
rect 646484 54649 646540 54658
rect 630742 43723 630794 43729
rect 630742 43665 630794 43671
rect 640726 43723 640778 43729
rect 640726 43665 640778 43671
rect 630754 42027 630782 43665
rect 630742 42021 630794 42027
rect 630742 41963 630794 41969
rect 539732 40506 539788 40515
rect 539732 40441 539788 40450
rect 475510 37433 475562 37439
rect 475510 37375 475562 37381
rect 514006 37433 514058 37439
rect 514006 37375 514058 37381
rect 420790 34547 420842 34553
rect 420790 34489 420842 34495
rect 444886 34547 444938 34553
rect 444886 34489 444938 34495
<< via2 >>
rect 175604 997714 175660 997770
rect 80564 997122 80620 997178
rect 129524 997122 129580 997178
rect 80564 982914 80620 982970
rect 132404 982914 132460 982970
rect 238964 997122 239020 997178
rect 238964 983062 239020 983118
rect 486740 997714 486796 997770
rect 538580 997714 538636 997770
rect 639380 997714 639436 997770
rect 293108 997122 293164 997178
rect 432020 997122 432076 997178
rect 287924 983062 287980 983118
rect 184244 982953 184246 982970
rect 184246 982953 184298 982970
rect 184298 982953 184300 982970
rect 184244 982914 184300 982953
rect 233204 982914 233260 982970
rect 239924 982914 239980 982970
rect 285044 982914 285100 982970
rect 293108 982914 293164 982970
rect 392468 982931 392524 982970
rect 392468 982914 392470 982931
rect 392470 982914 392522 982931
rect 392522 982914 392524 982931
rect 394580 982914 394636 982970
rect 399572 982914 399628 982970
rect 486740 982914 486796 982970
rect 538580 982914 538636 982970
rect 639380 982914 639436 982970
rect 40148 961915 40204 961954
rect 40148 961898 40150 961915
rect 40150 961898 40202 961915
rect 40202 961898 40204 961915
rect 60020 961750 60076 961806
rect 653780 959086 653836 959142
rect 676820 944325 676822 944342
rect 676822 944325 676874 944342
rect 676874 944325 676876 944342
rect 676820 944286 676876 944325
rect 676340 880202 676396 880258
rect 676148 879610 676204 879666
rect 654164 868806 654220 868862
rect 654068 867622 654124 867678
rect 676244 879166 676300 879222
rect 676052 878443 676108 878482
rect 676052 878426 676054 878443
rect 676054 878426 676106 878443
rect 676106 878426 676108 878443
rect 654260 866438 654316 866494
rect 654260 864087 654316 864126
rect 654260 864070 654262 864087
rect 654262 864070 654314 864087
rect 654314 864070 654316 864087
rect 654836 862886 654892 862942
rect 656372 861850 656428 861906
rect 41780 817933 41782 817950
rect 41782 817933 41834 817950
rect 41834 817933 41836 817950
rect 41780 817894 41836 817933
rect 41780 817319 41836 817358
rect 41780 817302 41782 817319
rect 41782 817302 41834 817319
rect 41834 817302 41836 817319
rect 41588 816579 41644 816618
rect 41588 816562 41590 816579
rect 41590 816562 41642 816579
rect 41642 816562 41644 816579
rect 41780 815839 41836 815878
rect 41780 815822 41782 815839
rect 41782 815822 41834 815839
rect 41834 815822 41836 815839
rect 41780 814877 41836 814916
rect 41780 814860 41782 814877
rect 41782 814860 41834 814877
rect 41834 814860 41836 814877
rect 41588 813619 41644 813658
rect 41588 813602 41590 813619
rect 41590 813602 41642 813619
rect 41642 813602 41644 813619
rect 42068 812862 42124 812918
rect 34484 812418 34540 812474
rect 34388 810198 34444 810254
rect 28820 805610 28876 805666
rect 28820 805166 28876 805222
rect 37364 811678 37420 811734
rect 41972 811308 42028 811364
rect 41780 810790 41836 810846
rect 40148 809606 40204 809662
rect 34484 805018 34540 805074
rect 40244 809458 40300 809514
rect 41588 808126 41644 808182
rect 41396 807090 41452 807146
rect 41588 806646 41644 806702
rect 41588 806054 41644 806110
rect 41588 805183 41644 805222
rect 41588 805166 41590 805183
rect 41590 805166 41642 805183
rect 41642 805166 41644 805183
rect 41876 808866 41932 808922
rect 41876 807830 41932 807886
rect 41876 801022 41932 801078
rect 42644 800726 42700 800782
rect 42644 798802 42700 798858
rect 43124 800430 43180 800486
rect 42164 790218 42220 790274
rect 41780 786370 41836 786426
rect 43028 793918 43084 793974
rect 41780 774695 41836 774734
rect 41780 774678 41782 774695
rect 41782 774678 41834 774695
rect 41834 774678 41836 774695
rect 41588 773955 41644 773994
rect 41588 773938 41590 773955
rect 41590 773938 41642 773955
rect 41642 773938 41644 773955
rect 41780 773511 41836 773550
rect 41780 773494 41782 773511
rect 41782 773494 41834 773511
rect 41834 773494 41836 773511
rect 43412 800578 43468 800634
rect 41588 773385 41590 773402
rect 41590 773385 41642 773402
rect 41642 773385 41644 773402
rect 41588 773346 41644 773385
rect 41780 772623 41836 772662
rect 41780 772606 41782 772623
rect 41782 772606 41834 772623
rect 41834 772606 41836 772623
rect 41588 772310 41644 772366
rect 43124 771905 43126 771922
rect 43126 771905 43178 771922
rect 43178 771905 43180 771922
rect 43124 771866 43180 771905
rect 41588 770830 41644 770886
rect 41780 769663 41836 769702
rect 41780 769646 41782 769663
rect 41782 769646 41834 769663
rect 41834 769646 41836 769663
rect 37364 768462 37420 768518
rect 28820 762394 28876 762450
rect 28820 761950 28876 762006
rect 42260 768166 42316 768222
rect 41876 767574 41932 767630
rect 40244 766390 40300 766446
rect 40148 766242 40204 766298
rect 41588 765502 41644 765558
rect 41780 765149 41836 765188
rect 41780 765132 41782 765149
rect 41782 765132 41834 765149
rect 41834 765132 41836 765149
rect 41588 763447 41644 763486
rect 41588 763430 41590 763447
rect 41590 763430 41642 763447
rect 41642 763430 41644 763447
rect 41780 762115 41836 762154
rect 41780 762098 41782 762115
rect 41782 762098 41834 762115
rect 41834 762098 41836 762115
rect 41012 760174 41068 760230
rect 41780 757954 41836 758010
rect 42068 767130 42124 767186
rect 41972 764170 42028 764226
rect 42164 764614 42220 764670
rect 42068 757806 42124 757862
rect 42836 752478 42892 752534
rect 42932 751146 42988 751202
rect 42836 747298 42892 747354
rect 41780 747002 41836 747058
rect 43028 748778 43084 748834
rect 41780 731479 41836 731518
rect 41780 731462 41782 731479
rect 41782 731462 41834 731479
rect 41834 731462 41836 731479
rect 41588 730739 41644 730778
rect 41588 730722 41590 730739
rect 41590 730722 41642 730739
rect 41642 730722 41644 730739
rect 41780 730369 41836 730408
rect 41780 730352 41782 730369
rect 41782 730352 41834 730369
rect 41834 730352 41836 730369
rect 41588 730169 41590 730186
rect 41590 730169 41642 730186
rect 41642 730169 41644 730186
rect 41588 730130 41644 730169
rect 41204 729242 41260 729298
rect 41588 729259 41644 729298
rect 41588 729242 41590 729259
rect 41590 729242 41642 729259
rect 41642 729242 41644 729259
rect 40436 728650 40492 728706
rect 41588 728667 41644 728706
rect 41588 728650 41590 728667
rect 41590 728650 41642 728667
rect 41642 728650 41644 728667
rect 41780 727927 41836 727966
rect 41780 727910 41782 727927
rect 41782 727910 41834 727927
rect 41834 727910 41836 727927
rect 34484 726726 34540 726782
rect 28820 719178 28876 719234
rect 28820 718734 28876 718790
rect 41780 726430 41836 726486
rect 37364 725246 37420 725302
rect 41972 724950 42028 725006
rect 41780 724358 41836 724414
rect 40148 723174 40204 723230
rect 37364 718586 37420 718642
rect 34484 717698 34540 717754
rect 40244 723026 40300 723082
rect 41588 722286 41644 722342
rect 41588 720806 41644 720862
rect 41588 720231 41644 720270
rect 41588 720214 41590 720231
rect 41590 720214 41642 720231
rect 41642 720214 41644 720231
rect 41588 718751 41644 718790
rect 41588 718734 41590 718751
rect 41590 718734 41642 718751
rect 41642 718734 41644 718751
rect 40244 716958 40300 717014
rect 40148 716810 40204 716866
rect 41876 721916 41932 721972
rect 42260 721398 42316 721454
rect 42836 708522 42892 708578
rect 42740 705414 42796 705470
rect 41780 701270 41836 701326
rect 43124 708818 43180 708874
rect 43028 708670 43084 708726
rect 42932 705858 42988 705914
rect 42836 702010 42892 702066
rect 41780 688263 41836 688302
rect 41780 688246 41782 688263
rect 41782 688246 41834 688263
rect 41834 688246 41836 688263
rect 41588 687523 41644 687562
rect 41588 687506 41590 687523
rect 41590 687506 41642 687523
rect 41642 687506 41644 687523
rect 41780 687227 41836 687266
rect 41780 687210 41782 687227
rect 41782 687210 41834 687227
rect 41834 687210 41836 687227
rect 41588 686953 41590 686970
rect 41590 686953 41642 686970
rect 41642 686953 41644 686970
rect 41588 686914 41644 686953
rect 41588 686043 41644 686082
rect 41588 686026 41590 686043
rect 41590 686026 41642 686043
rect 41642 686026 41644 686043
rect 41780 685325 41782 685342
rect 41782 685325 41834 685342
rect 41834 685325 41836 685342
rect 41780 685286 41836 685325
rect 41588 684563 41644 684602
rect 41588 684546 41590 684563
rect 41590 684546 41642 684563
rect 41642 684546 41644 684563
rect 41780 684141 41782 684158
rect 41782 684141 41834 684158
rect 41834 684141 41836 684158
rect 41780 684102 41836 684141
rect 41780 683214 41836 683270
rect 42260 681142 42316 681198
rect 41588 679070 41644 679126
rect 41780 677237 41836 677276
rect 41780 677220 41782 677237
rect 41782 677220 41834 677237
rect 41834 677220 41836 677237
rect 41780 676702 41836 676758
rect 28820 675962 28876 676018
rect 41780 675757 41836 675796
rect 41780 675740 41782 675757
rect 41782 675740 41834 675757
rect 41834 675740 41836 675757
rect 28820 675518 28876 675574
rect 42932 668562 42988 668618
rect 42836 668414 42892 668470
rect 42740 668266 42796 668322
rect 42740 665306 42796 665362
rect 42356 662346 42412 662402
rect 43028 666194 43084 666250
rect 42932 664270 42988 664326
rect 42836 663974 42892 664030
rect 43124 665454 43180 665510
rect 43028 661458 43084 661514
rect 41588 644899 41644 644938
rect 41588 644882 41590 644899
rect 41590 644882 41642 644899
rect 41642 644882 41644 644899
rect 41588 644307 41644 644346
rect 41588 644290 41590 644307
rect 41590 644290 41642 644307
rect 41642 644290 41644 644307
rect 41780 644011 41836 644050
rect 41780 643994 41782 644011
rect 41782 643994 41834 644011
rect 41834 643994 41836 644011
rect 41588 643737 41590 643754
rect 41590 643737 41642 643754
rect 41642 643737 41644 643754
rect 41588 643698 41644 643737
rect 41588 642827 41644 642866
rect 41588 642810 41590 642827
rect 41590 642810 41642 642827
rect 41642 642810 41644 642827
rect 43124 642218 43180 642274
rect 41588 641347 41644 641386
rect 41588 641330 41590 641347
rect 41590 641330 41642 641347
rect 41642 641330 41644 641347
rect 41588 639850 41644 639906
rect 41876 637926 41932 637982
rect 41780 636076 41836 636132
rect 41780 634078 41836 634134
rect 41780 633486 41836 633542
rect 28820 632746 28876 632802
rect 41780 632541 41836 632580
rect 41780 632524 41782 632541
rect 41782 632524 41834 632541
rect 41834 632524 41836 632541
rect 28820 632302 28876 632358
rect 42932 625938 42988 625994
rect 42836 625050 42892 625106
rect 42836 622090 42892 622146
rect 42164 620758 42220 620814
rect 43028 623866 43084 623922
rect 42932 621350 42988 621406
rect 42164 617206 42220 617262
rect 41780 616614 41836 616670
rect 43124 621942 43180 621998
rect 43028 617650 43084 617706
rect 40340 601666 40396 601722
rect 41588 601518 41644 601574
rect 41780 601387 41836 601426
rect 41780 601370 41782 601387
rect 41782 601370 41834 601387
rect 41834 601370 41836 601387
rect 41780 600795 41836 600834
rect 41780 600778 41782 600795
rect 41782 600778 41834 600795
rect 41834 600778 41836 600795
rect 43412 641034 43468 641090
rect 41780 600373 41782 600390
rect 41782 600373 41834 600390
rect 41834 600373 41836 600390
rect 41780 600334 41836 600373
rect 41780 599833 41836 599872
rect 41780 599816 41782 599833
rect 41782 599816 41834 599833
rect 41834 599816 41836 599833
rect 41780 599315 41836 599354
rect 41780 599298 41782 599315
rect 41782 599298 41834 599315
rect 41834 599298 41836 599315
rect 40340 598706 40396 598762
rect 41780 598353 41836 598392
rect 41780 598336 41782 598353
rect 41782 598336 41834 598353
rect 41834 598336 41836 598353
rect 39764 597966 39820 598022
rect 41588 596651 41644 596690
rect 41588 596634 41590 596651
rect 41590 596634 41642 596651
rect 41642 596634 41644 596651
rect 41876 594784 41932 594840
rect 41780 592934 41836 592990
rect 41780 590879 41836 590918
rect 41780 590862 41782 590879
rect 41782 590862 41834 590879
rect 41834 590862 41836 590879
rect 28820 589530 28876 589586
rect 28820 589086 28876 589142
rect 41588 589086 41644 589142
rect 42452 583018 42508 583074
rect 42836 581686 42892 581742
rect 42452 578874 42508 578930
rect 42356 576062 42412 576118
rect 43124 582574 43180 582630
rect 42932 579466 42988 579522
rect 43124 580502 43180 580558
rect 43028 576358 43084 576414
rect 42932 576210 42988 576266
rect 42836 573842 42892 573898
rect 41780 540394 41836 540450
rect 41780 538766 41836 538822
rect 41780 536842 41836 536898
rect 41780 534770 41836 534826
rect 41780 534474 41836 534530
rect 41876 533586 41932 533642
rect 41780 531366 41836 531422
rect 41780 530626 41836 530682
rect 41780 530034 41836 530090
rect 42164 529294 42220 529350
rect 42164 527666 42220 527722
rect 42068 527074 42124 527130
rect 42068 526482 42124 526538
rect 41780 476053 41782 476070
rect 41782 476053 41834 476070
rect 41834 476053 41836 476070
rect 41780 476014 41836 476053
rect 41780 475535 41782 475552
rect 41782 475535 41834 475552
rect 41834 475535 41836 475552
rect 41780 475496 41836 475535
rect 41780 474978 41836 475034
rect 40340 473794 40396 473850
rect 39668 472314 39724 472370
rect 34484 464322 34540 464378
rect 23060 463730 23116 463786
rect 23060 463286 23116 463342
rect 41684 473202 41740 473258
rect 41588 465249 41590 465266
rect 41590 465249 41642 465266
rect 41642 465249 41644 465266
rect 41588 465210 41644 465249
rect 41876 474573 41878 474590
rect 41878 474573 41930 474590
rect 41930 474573 41932 474590
rect 41876 474534 41932 474573
rect 43316 473054 43372 473110
rect 41780 472035 41836 472074
rect 41780 472018 41782 472035
rect 41782 472018 41834 472035
rect 41834 472018 41836 472035
rect 41780 463599 41836 463638
rect 41780 463582 41782 463599
rect 41782 463582 41834 463599
rect 41834 463582 41836 463599
rect 41588 428523 41644 428562
rect 41588 428506 41590 428523
rect 41590 428506 41642 428523
rect 41642 428506 41644 428523
rect 40340 427914 40396 427970
rect 41588 427043 41644 427082
rect 41588 427026 41590 427043
rect 41590 427026 41642 427043
rect 41642 427026 41644 427043
rect 41780 429263 41836 429302
rect 41780 429246 41782 429263
rect 41782 429246 41834 429263
rect 41834 429246 41836 429263
rect 41780 428227 41836 428266
rect 41780 428210 41782 428227
rect 41782 428210 41834 428227
rect 41834 428210 41836 428227
rect 41780 426673 41836 426712
rect 41780 426656 41782 426673
rect 41782 426656 41834 426673
rect 41834 426656 41836 426673
rect 41684 426434 41740 426490
rect 41588 425546 41644 425602
rect 41684 424954 41740 425010
rect 41588 420070 41644 420126
rect 28916 416962 28972 417018
rect 28916 416518 28972 416574
rect 41588 416535 41644 416574
rect 41588 416518 41590 416535
rect 41590 416518 41642 416535
rect 41642 416518 41644 416535
rect 41780 422142 41836 422198
rect 41876 411634 41932 411690
rect 41780 408378 41836 408434
rect 41780 407934 41836 407990
rect 42164 407342 42220 407398
rect 42068 406454 42124 406510
rect 41780 404234 41836 404290
rect 41780 403642 41836 403698
rect 41780 402902 41836 402958
rect 41780 402310 41836 402366
rect 41876 400238 41932 400294
rect 41780 399794 41836 399850
rect 42164 399350 42220 399406
rect 41780 386047 41836 386086
rect 41780 386030 41782 386047
rect 41782 386030 41834 386047
rect 41834 386030 41836 386047
rect 41588 385307 41644 385346
rect 41588 385290 41590 385307
rect 41590 385290 41642 385307
rect 41642 385290 41644 385307
rect 41780 385011 41836 385050
rect 41780 384994 41782 385011
rect 41782 384994 41834 385011
rect 41834 384994 41836 385011
rect 41588 384737 41590 384754
rect 41590 384737 41642 384754
rect 41642 384737 41644 384754
rect 41588 384698 41644 384737
rect 41588 383827 41644 383866
rect 41588 383810 41590 383827
rect 41590 383810 41642 383827
rect 41642 383810 41644 383827
rect 41780 383531 41836 383570
rect 41780 383514 41782 383531
rect 41782 383514 41834 383531
rect 41834 383514 41836 383531
rect 41588 383257 41590 383274
rect 41590 383257 41642 383274
rect 41642 383257 41644 383274
rect 41588 383218 41644 383257
rect 39956 382182 40012 382238
rect 41780 381999 41782 382016
rect 41782 381999 41834 382016
rect 41834 381999 41836 382016
rect 41780 381960 41836 381999
rect 41780 378926 41836 378982
rect 41588 376854 41644 376910
rect 28820 373746 28876 373802
rect 28820 373302 28876 373358
rect 41588 373319 41644 373358
rect 41588 373302 41590 373319
rect 41590 373302 41642 373319
rect 41642 373302 41644 373319
rect 42068 368418 42124 368474
rect 41780 365162 41836 365218
rect 41972 364570 42028 364626
rect 41780 364126 41836 364182
rect 42164 363534 42220 363590
rect 41780 361018 41836 361074
rect 41780 360426 41836 360482
rect 41780 359686 41836 359742
rect 42068 358946 42124 359002
rect 41780 357170 41836 357226
rect 41780 356578 41836 356634
rect 42164 356134 42220 356190
rect 41780 342831 41836 342870
rect 41780 342814 41782 342831
rect 41782 342814 41834 342831
rect 41834 342814 41836 342831
rect 41780 342313 41836 342352
rect 41780 342296 41782 342313
rect 41782 342296 41834 342313
rect 41834 342296 41836 342313
rect 41780 341795 41836 341834
rect 41780 341778 41782 341795
rect 41782 341778 41834 341795
rect 41834 341778 41836 341795
rect 41780 341373 41782 341390
rect 41782 341373 41834 341390
rect 41834 341373 41836 341390
rect 41780 341334 41836 341373
rect 41588 340611 41644 340650
rect 41588 340594 41590 340611
rect 41590 340594 41642 340611
rect 41642 340594 41644 340611
rect 41780 340315 41836 340354
rect 41780 340298 41782 340315
rect 41782 340298 41834 340315
rect 41834 340298 41836 340315
rect 41588 340041 41590 340058
rect 41590 340041 41642 340058
rect 41642 340041 41644 340058
rect 41588 340002 41644 340041
rect 41588 339131 41644 339170
rect 41588 339114 41590 339131
rect 41590 339114 41642 339131
rect 41642 339114 41644 339131
rect 41780 338857 41782 338874
rect 41782 338857 41834 338874
rect 41834 338857 41836 338874
rect 41780 338818 41836 338857
rect 34484 335562 34540 335618
rect 28820 330530 28876 330586
rect 28820 330086 28876 330142
rect 41780 330399 41836 330438
rect 41780 330382 41782 330399
rect 41782 330382 41834 330399
rect 41834 330382 41836 330399
rect 41780 325054 41836 325110
rect 41780 323278 41836 323334
rect 41780 321798 41836 321854
rect 42068 321206 42124 321262
rect 41876 320762 41932 320818
rect 42068 319874 42124 319930
rect 41876 317654 41932 317710
rect 41780 316766 41836 316822
rect 41780 316174 41836 316230
rect 41780 315582 41836 315638
rect 42164 313806 42220 313862
rect 41780 313214 41836 313270
rect 41780 312622 41836 312678
rect 41780 299615 41836 299654
rect 41780 299598 41782 299615
rect 41782 299598 41834 299615
rect 41834 299598 41836 299615
rect 41588 298710 41644 298766
rect 39668 296490 39724 296546
rect 41780 298579 41836 298618
rect 41780 298562 41782 298579
rect 41782 298562 41834 298579
rect 41834 298562 41836 298579
rect 41780 298157 41782 298174
rect 41782 298157 41834 298174
rect 41834 298157 41836 298174
rect 41780 298118 41836 298157
rect 41780 297617 41836 297656
rect 41780 297600 41782 297617
rect 41782 297600 41834 297617
rect 41834 297600 41836 297617
rect 41780 297099 41836 297138
rect 41780 297082 41782 297099
rect 41782 297082 41834 297099
rect 41834 297082 41836 297099
rect 39860 295898 39916 295954
rect 41588 295915 41644 295954
rect 41588 295898 41590 295915
rect 41590 295898 41642 295915
rect 41642 295898 41644 295915
rect 34484 292346 34540 292402
rect 28820 287314 28876 287370
rect 28820 286870 28876 286926
rect 41780 287183 41836 287222
rect 41780 287166 41782 287183
rect 41782 287166 41834 287183
rect 41834 287166 41836 287183
rect 42068 281838 42124 281894
rect 41780 280062 41836 280118
rect 41780 278730 41836 278786
rect 42068 277990 42124 278046
rect 41876 277546 41932 277602
rect 42068 276658 42124 276714
rect 41780 274438 41836 274494
rect 41780 273550 41836 273606
rect 41780 273254 41836 273310
rect 41780 272366 41836 272422
rect 41876 270590 41932 270646
rect 41780 269998 41836 270054
rect 42164 269554 42220 269610
rect 23156 254162 23212 254218
rect 23060 253274 23116 253330
rect 40244 256234 40300 256290
rect 41588 255642 41644 255698
rect 41780 255385 41782 255402
rect 41782 255385 41834 255402
rect 41834 255385 41836 255402
rect 41780 255346 41836 255385
rect 41780 254941 41782 254958
rect 41782 254941 41834 254958
rect 41834 254941 41836 254958
rect 41780 254902 41836 254941
rect 41780 254475 41836 254514
rect 41780 254458 41782 254475
rect 41782 254458 41834 254475
rect 41834 254458 41836 254475
rect 23348 253274 23404 253330
rect 23252 252682 23308 252738
rect 41684 249130 41740 249186
rect 41588 244690 41644 244746
rect 41780 244855 41836 244894
rect 41780 244838 41782 244855
rect 41782 244838 41834 244855
rect 41834 244838 41836 244855
rect 41588 243654 41644 243710
rect 42068 238622 42124 238678
rect 41876 236846 41932 236902
rect 41780 235514 41836 235570
rect 42164 234774 42220 234830
rect 42164 234330 42220 234386
rect 42164 233590 42220 233646
rect 41780 231222 41836 231278
rect 41780 230334 41836 230390
rect 41780 230038 41836 230094
rect 41780 229298 41836 229354
rect 41876 227374 41932 227430
rect 41780 226782 41836 226838
rect 42164 226338 42220 226394
rect 41780 213279 41782 213296
rect 41782 213279 41834 213296
rect 41834 213279 41836 213296
rect 41780 213240 41836 213279
rect 41588 212909 41590 212926
rect 41590 212909 41642 212926
rect 41642 212909 41644 212926
rect 41588 212870 41644 212909
rect 41780 212169 41782 212186
rect 41782 212169 41834 212186
rect 41834 212169 41836 212186
rect 41780 212130 41836 212169
rect 44468 278434 44524 278490
rect 44372 276214 44428 276270
rect 44660 277250 44716 277306
rect 44564 275474 44620 275530
rect 44852 277842 44908 277898
rect 45044 658794 45100 658850
rect 45044 572362 45100 572418
rect 45044 529294 45100 529350
rect 45044 473054 45100 473110
rect 45044 278582 45100 278638
rect 45140 276362 45196 276418
rect 44948 275030 45004 275086
rect 45236 270590 45292 270646
rect 44756 266298 44812 266354
rect 41780 211725 41782 211742
rect 41782 211725 41834 211742
rect 41834 211725 41836 211742
rect 41780 211686 41836 211725
rect 41588 211429 41590 211446
rect 41590 211429 41642 211446
rect 41642 211429 41644 211446
rect 41588 211390 41644 211429
rect 41780 210689 41782 210706
rect 41782 210689 41834 210706
rect 41834 210689 41836 210706
rect 41780 210650 41836 210689
rect 41780 210223 41836 210262
rect 41780 210206 41782 210223
rect 41782 210206 41834 210223
rect 41834 210206 41836 210223
rect 41588 209949 41590 209966
rect 41590 209949 41642 209966
rect 41642 209949 41644 209966
rect 41588 209910 41644 209949
rect 41588 209357 41590 209374
rect 41590 209357 41642 209374
rect 41642 209357 41644 209374
rect 41588 209318 41644 209357
rect 41780 206210 41836 206266
rect 41588 201513 41590 201530
rect 41590 201513 41642 201530
rect 41642 201513 41644 201530
rect 41588 201474 41644 201513
rect 41588 200921 41590 200938
rect 41590 200921 41642 200938
rect 41642 200921 41644 200938
rect 41588 200882 41644 200921
rect 41876 201661 41878 201678
rect 41878 201661 41930 201678
rect 41930 201661 41932 201678
rect 41876 201622 41932 201661
rect 41876 195406 41932 195462
rect 41780 193630 41836 193686
rect 42164 192298 42220 192354
rect 42164 191706 42220 191762
rect 41780 191114 41836 191170
rect 41780 190374 41836 190430
rect 42068 188006 42124 188062
rect 41780 187118 41836 187174
rect 41780 186822 41836 186878
rect 41780 185934 41836 185990
rect 42164 184158 42220 184214
rect 41780 183566 41836 183622
rect 41876 183122 41932 183178
rect 45428 278286 45484 278342
rect 46004 278138 46060 278194
rect 46292 263525 46294 263542
rect 46294 263525 46346 263542
rect 46346 263525 46348 263542
rect 46292 263486 46348 263525
rect 46196 263338 46252 263394
rect 58004 789791 58060 789830
rect 58004 789774 58006 789791
rect 58006 789774 58058 789791
rect 58058 789774 58060 789791
rect 57620 789626 57676 789682
rect 58196 788442 58252 788498
rect 58388 787258 58444 787314
rect 59636 785334 59692 785390
rect 58676 784890 58732 784946
rect 57908 747594 57964 747650
rect 54740 745983 54796 746022
rect 54740 745966 54742 745983
rect 54742 745966 54794 745983
rect 54794 745966 54796 745983
rect 54644 745818 54700 745874
rect 59636 745374 59692 745430
rect 57620 745226 57676 745282
rect 59252 744042 59308 744098
rect 59636 742858 59692 742914
rect 59732 741674 59788 741730
rect 58388 704378 58444 704434
rect 58772 702641 58774 702658
rect 58774 702641 58826 702658
rect 58826 702641 58828 702658
rect 58772 702602 58828 702641
rect 58676 700826 58732 700882
rect 59252 699642 59308 699698
rect 58868 698458 58924 698514
rect 59636 661162 59692 661218
rect 58772 659403 58828 659442
rect 58772 659386 58774 659403
rect 58774 659386 58826 659403
rect 58826 659386 58828 659403
rect 59156 657610 59212 657666
rect 58196 656426 58252 656482
rect 58388 655242 58444 655298
rect 58964 617946 59020 618002
rect 58196 615578 58252 615634
rect 59636 616209 59638 616226
rect 59638 616209 59690 616226
rect 59690 616209 59692 616226
rect 59636 616170 59692 616209
rect 58964 614394 59020 614450
rect 59636 613210 59692 613266
rect 59540 612026 59596 612082
rect 50516 275326 50572 275382
rect 50324 275178 50380 275234
rect 58964 574730 59020 574786
rect 59636 572993 59638 573010
rect 59638 572993 59690 573010
rect 59690 572993 59692 573010
rect 59636 572954 59692 572993
rect 58964 571178 59020 571234
rect 60404 569994 60460 570050
rect 59156 568810 59212 568866
rect 57716 531662 57772 531718
rect 57620 530478 57676 530534
rect 58964 527074 59020 527130
rect 58580 525890 58636 525946
rect 59348 524706 59404 524762
rect 58484 404086 58540 404142
rect 59636 402793 59638 402810
rect 59638 402793 59690 402810
rect 59690 402793 59692 402810
rect 59636 402754 59692 402793
rect 57620 400534 57676 400590
rect 59636 399942 59692 399998
rect 59732 399350 59788 399406
rect 59540 398166 59596 398222
rect 58292 360870 58348 360926
rect 59156 359686 59212 359742
rect 57620 357466 57676 357522
rect 58196 356134 58252 356190
rect 59636 356726 59692 356782
rect 58580 354950 58636 355006
rect 58484 317654 58540 317710
rect 59156 316470 59212 316526
rect 59060 314102 59116 314158
rect 59636 313510 59692 313566
rect 59732 312918 59788 312974
rect 59540 311734 59596 311790
rect 59636 295158 59692 295214
rect 58196 293974 58252 294030
rect 59060 292790 59116 292846
rect 59636 291606 59692 291662
rect 60212 291458 60268 291514
rect 57524 290274 57580 290330
rect 59636 288071 59692 288110
rect 59636 288054 59638 288071
rect 59638 288054 59690 288071
rect 59690 288054 59692 288071
rect 58100 286870 58156 286926
rect 59540 285686 59596 285742
rect 57620 284502 57676 284558
rect 59636 283318 59692 283374
rect 58964 282430 59020 282486
rect 58196 280950 58252 281006
rect 59636 279766 59692 279822
rect 61940 276066 61996 276122
rect 61844 266890 61900 266946
rect 62132 277990 62188 278046
rect 62324 277694 62380 277750
rect 62036 266742 62092 266798
rect 62708 277546 62764 277602
rect 62804 277398 62860 277454
rect 62516 271478 62572 271534
rect 62228 266594 62284 266650
rect 65876 269258 65932 269314
rect 70580 272070 70636 272126
rect 69428 269554 69484 269610
rect 72980 272218 73036 272274
rect 71732 269406 71788 269462
rect 78836 272366 78892 272422
rect 77588 269702 77644 269758
rect 62900 266446 62956 266502
rect 88340 272514 88396 272570
rect 91892 272662 91948 272718
rect 139124 269850 139180 269906
rect 148340 244542 148396 244598
rect 148244 239658 148300 239714
rect 146996 235975 147052 236014
rect 146996 235958 146998 235975
rect 146998 235958 147050 235975
rect 147050 235958 147052 235975
rect 147476 231074 147532 231130
rect 147092 229890 147148 229946
rect 147092 226338 147148 226394
rect 147284 217771 147340 217810
rect 147284 217754 147286 217771
rect 147286 217754 147338 217771
rect 147338 217754 147340 217771
rect 146900 212870 146956 212926
rect 147092 211686 147148 211742
rect 147476 210371 147532 210410
rect 147476 210354 147478 210371
rect 147478 210354 147530 210371
rect 147530 210354 147532 210371
rect 146900 209170 146956 209226
rect 147188 207986 147244 208042
rect 146900 206358 146956 206414
rect 147860 203250 147916 203306
rect 147572 199550 147628 199606
rect 147284 195850 147340 195906
rect 147668 189782 147724 189838
rect 147764 175130 147820 175186
rect 148724 243358 148780 243414
rect 148532 242026 148588 242082
rect 148436 238474 148492 238530
rect 148628 236698 148684 236754
rect 148916 240842 148972 240898
rect 148820 234774 148876 234830
rect 148724 169062 148780 169118
rect 148532 168026 148588 168082
rect 148436 165510 148492 165566
rect 148244 164326 148300 164382
rect 147092 159442 147148 159498
rect 147092 156926 147148 156982
rect 147092 141255 147148 141294
rect 147092 141238 147094 141255
rect 147094 141238 147146 141255
rect 147146 141238 147148 141255
rect 146900 139906 146956 139962
rect 148340 161810 148396 161866
rect 148628 166250 148684 166306
rect 148436 124218 148492 124274
rect 149012 233590 149068 233646
rect 149108 232258 149164 232314
rect 149396 228114 149452 228170
rect 149492 227374 149548 227430
rect 149396 225154 149452 225210
rect 149492 223822 149548 223878
rect 149396 222638 149452 222694
rect 149492 221454 149548 221510
rect 149396 219678 149452 219734
rect 149396 218955 149452 218994
rect 149396 218938 149398 218955
rect 149398 218938 149450 218955
rect 149450 218938 149452 218955
rect 149396 216570 149452 216626
rect 149492 214794 149548 214850
rect 149396 214054 149452 214110
rect 149492 205618 149548 205674
rect 149396 204434 149452 204490
rect 149396 201639 149452 201678
rect 149396 201622 149398 201639
rect 149398 201622 149450 201639
rect 149450 201622 149452 201639
rect 149396 200734 149452 200790
rect 149300 198366 149356 198422
rect 149396 197034 149452 197090
rect 149492 194666 149548 194722
rect 149396 193186 149452 193242
rect 149492 192150 149548 192206
rect 149396 190966 149452 191022
rect 149300 188006 149356 188062
rect 149204 184454 149260 184510
rect 149396 187414 149452 187470
rect 149588 186230 149644 186286
rect 149492 183714 149548 183770
rect 149396 182530 149452 182586
rect 149492 181346 149548 181402
rect 149300 179570 149356 179626
rect 149396 178830 149452 178886
rect 149492 177646 149548 177702
rect 149396 176462 149452 176518
rect 149108 173946 149164 174002
rect 148916 163142 148972 163198
rect 148820 160626 148876 160682
rect 148820 133838 148876 133894
rect 148532 122442 148588 122498
rect 148340 110898 148396 110954
rect 147860 108399 147916 108438
rect 147860 108382 147862 108399
rect 147862 108382 147914 108399
rect 147914 108382 147916 108399
rect 147188 107215 147244 107254
rect 147188 107198 147190 107215
rect 147190 107198 147242 107215
rect 147242 107198 147244 107215
rect 148244 104682 148300 104738
rect 148436 103498 148492 103554
rect 148724 121702 148780 121758
rect 149300 170986 149356 171042
rect 149204 170246 149260 170302
rect 149588 172762 149644 172818
rect 149396 157962 149452 158018
rect 149396 155759 149452 155798
rect 149396 155742 149398 155759
rect 149398 155742 149450 155759
rect 149450 155742 149452 155759
rect 149492 154558 149548 154614
rect 149396 152930 149452 152986
rect 149492 150858 149548 150914
rect 149396 149822 149452 149878
rect 149492 148490 149548 148546
rect 149012 132654 149068 132710
rect 148820 115190 148876 115246
rect 148724 111934 148780 111990
rect 148820 106014 148876 106070
rect 149396 147306 149452 147362
rect 149492 146122 149548 146178
rect 149396 144494 149452 144550
rect 149492 143606 149548 143662
rect 149396 142422 149452 142478
rect 149396 138722 149452 138778
rect 149396 135910 149452 135966
rect 149684 152042 149740 152098
rect 149684 137538 149740 137594
rect 149396 135022 149452 135078
rect 149300 130878 149356 130934
rect 149396 130286 149452 130342
rect 149108 129102 149164 129158
rect 149396 127918 149452 127974
rect 149300 126586 149356 126642
rect 148916 102314 148972 102370
rect 148724 86495 148780 86534
rect 148724 86478 148726 86495
rect 148726 86478 148778 86495
rect 148778 86478 148780 86495
rect 149588 125402 149644 125458
rect 149396 120518 149452 120574
rect 149492 119334 149548 119390
rect 149396 118167 149452 118206
rect 149396 118150 149398 118167
rect 149398 118150 149450 118167
rect 149450 118150 149452 118167
rect 149492 116818 149548 116874
rect 149396 115634 149452 115690
rect 149396 115190 149452 115246
rect 149492 114450 149548 114506
rect 149396 113118 149452 113174
rect 149396 109583 149452 109622
rect 149396 109566 149398 109583
rect 149398 109566 149450 109583
rect 149450 109566 149452 109583
rect 149396 100851 149452 100890
rect 149396 100834 149398 100851
rect 149398 100834 149450 100851
rect 149450 100834 149452 100851
rect 149492 99798 149548 99854
rect 149396 98614 149452 98670
rect 149492 97430 149548 97486
rect 149396 95654 149452 95710
rect 149588 94914 149644 94970
rect 149492 93730 149548 93786
rect 149396 92546 149452 92602
rect 149300 91362 149356 91418
rect 149204 90178 149260 90234
rect 148628 85294 148684 85350
rect 146996 84110 147052 84166
rect 148244 81594 148300 81650
rect 148916 82334 148972 82390
rect 148820 77894 148876 77950
rect 149396 88994 149452 89050
rect 149492 87218 149548 87274
rect 149588 80410 149644 80466
rect 149396 76710 149452 76766
rect 149204 75526 149260 75582
rect 149012 73010 149068 73066
rect 149108 71974 149164 72030
rect 149300 73750 149356 73806
rect 149684 79226 149740 79282
rect 184340 219530 184396 219586
rect 184340 218829 184342 218846
rect 184342 218829 184394 218846
rect 184394 218829 184396 218846
rect 184340 218790 184396 218829
rect 184340 199698 184396 199754
rect 184244 197626 184300 197682
rect 184340 196738 184396 196794
rect 194420 272218 194476 272274
rect 193748 272070 193804 272126
rect 192404 269258 192460 269314
rect 185588 220270 185644 220326
rect 185492 198218 185548 198274
rect 184436 195998 184492 196054
rect 184340 195258 184396 195314
rect 184436 194370 184492 194426
rect 184532 193778 184588 193834
rect 184436 192890 184492 192946
rect 184340 192298 184396 192354
rect 184532 191410 184588 191466
rect 184628 190670 184684 190726
rect 184340 189969 184342 189986
rect 184342 189969 184394 189986
rect 184394 189969 184396 189986
rect 184340 189930 184396 189969
rect 184340 188450 184396 188506
rect 184532 189190 184588 189246
rect 184436 187562 184492 187618
rect 184340 186822 184396 186878
rect 184436 185342 184492 185398
rect 185396 186082 185452 186138
rect 184532 184602 184588 184658
rect 184340 183862 184396 183918
rect 184436 183122 184492 183178
rect 184532 181494 184588 181550
rect 184340 180754 184396 180810
rect 184436 180014 184492 180070
rect 184532 179274 184588 179330
rect 184628 178534 184684 178590
rect 184340 177646 184396 177702
rect 184436 177054 184492 177110
rect 184532 176166 184588 176222
rect 184340 175591 184396 175630
rect 184340 175574 184342 175591
rect 184342 175574 184394 175591
rect 184394 175574 184396 175591
rect 184436 173946 184492 174002
rect 184340 172466 184396 172522
rect 184532 171726 184588 171782
rect 184436 170838 184492 170894
rect 184628 170246 184684 170302
rect 184340 169358 184396 169414
rect 184532 168618 184588 168674
rect 184628 167878 184684 167934
rect 184436 167138 184492 167194
rect 184340 166398 184396 166454
rect 184532 165658 184588 165714
rect 186068 205914 186124 205970
rect 185972 204286 186028 204342
rect 186356 213462 186412 213518
rect 186548 214942 186604 214998
rect 186452 210502 186508 210558
rect 186932 221010 186988 221066
rect 187124 243358 187180 243414
rect 187028 218050 187084 218106
rect 186836 216422 186892 216478
rect 186740 211982 186796 212038
rect 186644 209022 186700 209078
rect 186260 207246 186316 207302
rect 186164 202806 186220 202862
rect 185876 174686 185932 174742
rect 185684 173206 185740 173262
rect 184436 164770 184492 164826
rect 184340 164047 184396 164086
rect 184340 164030 184342 164047
rect 184342 164030 184394 164047
rect 184394 164030 184396 164047
rect 184340 162550 184396 162606
rect 184532 163290 184588 163346
rect 184436 161810 184492 161866
rect 184340 160961 184342 160978
rect 184342 160961 184394 160978
rect 184394 160961 184396 160978
rect 184340 160922 184396 160961
rect 184436 160330 184492 160386
rect 184628 159442 184684 159498
rect 184532 158850 184588 158906
rect 184340 157962 184396 158018
rect 184436 157370 184492 157426
rect 184628 156482 184684 156538
rect 184532 155594 184588 155650
rect 184340 154114 184396 154170
rect 184532 155002 184588 155058
rect 184436 153522 184492 153578
rect 184628 152634 184684 152690
rect 184340 151894 184396 151950
rect 184436 151154 184492 151210
rect 184532 150414 184588 150470
rect 184340 149713 184342 149730
rect 184342 149713 184394 149730
rect 184394 149713 184396 149730
rect 184340 149674 184396 149713
rect 184436 148934 184492 148990
rect 184340 148046 184396 148102
rect 184532 147306 184588 147362
rect 184340 146566 184396 146622
rect 184436 145086 184492 145142
rect 184532 144346 184588 144402
rect 184340 142718 184396 142774
rect 184436 142126 184492 142182
rect 185396 143606 185452 143662
rect 184532 141238 184588 141294
rect 184340 140498 184396 140554
rect 184436 139758 184492 139814
rect 184532 138870 184588 138926
rect 184628 138278 184684 138334
rect 184436 134430 184492 134486
rect 184532 133690 184588 133746
rect 184340 132950 184396 133006
rect 184340 132227 184396 132266
rect 184340 132210 184342 132227
rect 184342 132210 184394 132227
rect 184394 132210 184396 132227
rect 184436 131470 184492 131526
rect 184532 130582 184588 130638
rect 184628 129842 184684 129898
rect 184340 129102 184396 129158
rect 184436 128362 184492 128418
rect 184532 127622 184588 127678
rect 184628 126882 184684 126938
rect 184340 125994 184396 126050
rect 184436 125402 184492 125458
rect 184532 124514 184588 124570
rect 184340 123774 184396 123830
rect 184436 123034 184492 123090
rect 184628 122146 184684 122202
rect 184532 121554 184588 121610
rect 184436 120666 184492 120722
rect 184532 120074 184588 120130
rect 184340 119186 184396 119242
rect 184628 118594 184684 118650
rect 184340 117706 184396 117762
rect 184436 116966 184492 117022
rect 184532 116226 184588 116282
rect 184628 115338 184684 115394
rect 184340 114746 184396 114802
rect 184436 113858 184492 113914
rect 184628 113118 184684 113174
rect 184532 112378 184588 112434
rect 184340 111638 184396 111694
rect 184532 110898 184588 110954
rect 184436 107790 184492 107846
rect 184340 107050 184396 107106
rect 184340 105570 184396 105626
rect 184532 104830 184588 104886
rect 184436 103942 184492 103998
rect 184340 103350 184396 103406
rect 184436 101870 184492 101926
rect 184532 100982 184588 101038
rect 184340 100242 184396 100298
rect 184436 99502 184492 99558
rect 184532 98614 184588 98670
rect 185972 136798 186028 136854
rect 185780 135910 185836 135966
rect 193076 269554 193132 269610
rect 194228 269406 194284 269462
rect 196628 272366 196684 272422
rect 196148 269702 196204 269758
rect 199220 272514 199276 272570
rect 200468 272662 200524 272718
rect 209588 268074 209644 268130
rect 213332 269850 213388 269906
rect 214292 268074 214348 268130
rect 347636 274290 347692 274346
rect 353396 274438 353452 274494
rect 370100 271774 370156 271830
rect 369620 271626 369676 271682
rect 368372 268962 368428 269018
rect 367892 268814 367948 268870
rect 373460 274586 373516 274642
rect 374324 269110 374380 269166
rect 376244 274734 376300 274790
rect 375572 271922 375628 271978
rect 377012 270442 377068 270498
rect 379124 274882 379180 274938
rect 378644 273402 378700 273458
rect 381236 273550 381292 273606
rect 381812 275918 381868 275974
rect 381236 267926 381292 267982
rect 382964 273254 383020 273310
rect 385556 270294 385612 270350
rect 387284 273106 387340 273162
rect 388436 270146 388492 270202
rect 388628 267926 388684 267982
rect 390356 275770 390412 275826
rect 390164 272958 390220 273014
rect 391508 269998 391564 270054
rect 392756 272810 392812 272866
rect 396692 276510 396748 276566
rect 397076 269850 397132 269906
rect 398708 272662 398764 272718
rect 402548 276658 402604 276714
rect 401300 272514 401356 272570
rect 403028 269702 403084 269758
rect 404180 272366 404236 272422
rect 405620 269554 405676 269610
rect 408980 275622 409036 275678
rect 408980 273550 409036 273606
rect 410900 272218 410956 272274
rect 410420 269406 410476 269462
rect 411764 272070 411820 272126
rect 411572 269258 411628 269314
rect 489044 274290 489100 274346
rect 503156 274438 503212 274494
rect 529844 276658 529900 276714
rect 540980 268962 541036 269018
rect 539828 268814 539884 268870
rect 544532 271774 544588 271830
rect 543380 271626 543436 271682
rect 552788 274586 552844 274642
rect 555188 269110 555244 269166
rect 559892 274734 559948 274790
rect 558740 271922 558796 271978
rect 566996 274882 567052 274938
rect 565844 273402 565900 273458
rect 562292 270442 562348 270498
rect 574100 275918 574156 275974
rect 576500 273254 576556 273310
rect 583604 270294 583660 270350
rect 587156 273106 587212 273162
rect 590612 270146 590668 270202
rect 595412 275770 595468 275826
rect 594164 272958 594220 273014
rect 597716 269998 597772 270054
rect 601268 272810 601324 272866
rect 610772 276510 610828 276566
rect 615476 272662 615532 272718
rect 611924 269850 611980 269906
rect 622580 272514 622636 272570
rect 626132 269702 626188 269758
rect 629684 272366 629740 272422
rect 633236 269554 633292 269610
rect 646580 277250 646636 277306
rect 646484 275474 646540 275530
rect 646196 272218 646252 272274
rect 645044 269406 645100 269462
rect 420404 262171 420460 262210
rect 420404 262154 420406 262171
rect 420406 262154 420458 262171
rect 420458 262154 420460 262171
rect 420404 259786 420460 259842
rect 191540 259342 191596 259398
rect 190196 251646 190252 251702
rect 420404 256974 420460 257030
rect 420404 255198 420460 255254
rect 420404 252830 420460 252886
rect 420308 250462 420364 250518
rect 420404 248094 420460 248150
rect 420404 245282 420460 245338
rect 420404 243506 420460 243562
rect 420404 241138 420460 241194
rect 412148 240102 412204 240158
rect 412052 239971 412108 240010
rect 412052 239954 412054 239971
rect 412054 239954 412106 239971
rect 412106 239954 412108 239971
rect 292148 229002 292204 229058
rect 293108 228854 293164 228910
rect 296564 229150 296620 229206
rect 299444 234922 299500 234978
rect 299348 234626 299404 234682
rect 307604 231074 307660 231130
rect 316724 231222 316780 231278
rect 318932 225302 318988 225358
rect 319508 231370 319564 231426
rect 322484 231518 322540 231574
rect 328052 225598 328108 225654
rect 327764 225450 327820 225506
rect 330260 231666 330316 231722
rect 330836 225746 330892 225802
rect 332564 234034 332620 234090
rect 333812 231814 333868 231870
rect 333044 228114 333100 228170
rect 336884 227374 336940 227430
rect 339380 228262 339436 228318
rect 340148 225894 340204 225950
rect 341588 234182 341644 234238
rect 342548 235662 342604 235718
rect 342164 228558 342220 228614
rect 343124 227226 343180 227282
rect 343988 233146 344044 233202
rect 345428 228410 345484 228466
rect 344756 227078 344812 227134
rect 347636 234774 347692 234830
rect 354644 234922 354700 234978
rect 354164 222934 354220 222990
rect 356852 236106 356908 236162
rect 356756 234922 356812 234978
rect 355604 222638 355660 222694
rect 357236 222786 357292 222842
rect 358964 230038 359020 230094
rect 358580 224562 358636 224618
rect 359444 224414 359500 224470
rect 359828 229002 359884 229058
rect 359732 224266 359788 224322
rect 360884 228706 360940 228762
rect 360308 224118 360364 224174
rect 361460 223970 361516 224026
rect 363572 230186 363628 230242
rect 362804 229150 362860 229206
rect 364052 233738 364108 233794
rect 365684 233294 365740 233350
rect 364148 223822 364204 223878
rect 366644 229890 366700 229946
rect 365684 228854 365740 228910
rect 367220 235514 367276 235570
rect 368948 236402 369004 236458
rect 368660 231814 368716 231870
rect 367604 223674 367660 223730
rect 370388 236698 370444 236754
rect 368660 225154 368716 225210
rect 372212 236994 372268 237050
rect 371156 232998 371212 233054
rect 370772 232850 370828 232906
rect 373460 236846 373516 236902
rect 374036 232702 374092 232758
rect 373076 229742 373132 229798
rect 374900 236254 374956 236310
rect 375380 232554 375436 232610
rect 376724 223378 376780 223434
rect 377972 236550 378028 236606
rect 377972 236254 378028 236310
rect 378164 236254 378220 236310
rect 379124 234478 379180 234534
rect 380084 233294 380140 233350
rect 379892 229594 379948 229650
rect 377588 223526 377644 223582
rect 382388 236254 382444 236310
rect 382580 236254 382636 236310
rect 382100 234330 382156 234386
rect 381716 232406 381772 232462
rect 382676 231962 382732 232018
rect 381332 229446 381388 229502
rect 381236 223230 381292 223286
rect 383540 229298 383596 229354
rect 384980 232258 385036 232314
rect 385268 232110 385324 232166
rect 384404 229150 384460 229206
rect 384308 223082 384364 223138
rect 385844 235958 385900 236014
rect 386996 236254 387052 236310
rect 387380 236846 387436 236902
rect 387572 236863 387628 236902
rect 387572 236846 387574 236863
rect 387574 236846 387626 236863
rect 387626 236846 387628 236863
rect 387380 236402 387436 236458
rect 389876 235810 389932 235866
rect 390740 235662 390796 235718
rect 391604 226930 391660 226986
rect 391220 226782 391276 226838
rect 393044 235662 393100 235718
rect 394100 226634 394156 226690
rect 394484 226486 394540 226542
rect 396980 236994 397036 237050
rect 397076 236863 397132 236902
rect 397076 236846 397078 236863
rect 397078 236846 397130 236863
rect 397130 236846 397132 236863
rect 397652 236994 397708 237050
rect 397364 236254 397420 236310
rect 397748 235514 397804 235570
rect 398036 236863 398092 236902
rect 398036 236846 398038 236863
rect 398038 236846 398090 236863
rect 398090 236846 398092 236863
rect 398324 236846 398380 236902
rect 399860 235514 399916 235570
rect 400244 233886 400300 233942
rect 400244 229002 400300 229058
rect 399476 228854 399532 228910
rect 401396 235366 401452 235422
rect 402644 235218 402700 235274
rect 403124 234922 403180 234978
rect 403988 234922 404044 234978
rect 404372 226338 404428 226394
rect 405428 235070 405484 235126
rect 405332 234774 405388 234830
rect 405524 234774 405580 234830
rect 406484 236106 406540 236162
rect 406004 234626 406060 234682
rect 405908 233738 405964 233794
rect 405812 231814 405868 231870
rect 405716 226190 405772 226246
rect 407444 236698 407500 236754
rect 407444 236254 407500 236310
rect 406484 222490 406540 222546
rect 409940 236106 409996 236162
rect 408500 234626 408556 234682
rect 409844 234478 409900 234534
rect 408116 230334 408172 230390
rect 407636 226042 407692 226098
rect 410036 234330 410092 234386
rect 411380 234478 411436 234534
rect 410804 234330 410860 234386
rect 567380 239954 567436 240010
rect 413396 238918 413452 238974
rect 414068 238770 414124 238826
rect 413684 238622 413740 238678
rect 413972 238326 414028 238382
rect 415220 238178 415276 238234
rect 414452 238030 414508 238086
rect 413684 236254 413740 236310
rect 415220 236254 415276 236310
rect 415412 236254 415468 236310
rect 413876 236106 413932 236162
rect 424724 231074 424780 231130
rect 442868 231222 442924 231278
rect 445172 225302 445228 225358
rect 448916 231370 448972 231426
rect 455252 231518 455308 231574
rect 457268 225450 457324 225506
rect 463316 225598 463372 225654
rect 470132 231666 470188 231722
rect 469364 225746 469420 225802
rect 472340 234034 472396 234090
rect 476180 228114 476236 228170
rect 475316 225154 475372 225210
rect 480884 233886 480940 233942
rect 481460 227374 481516 227430
rect 488276 228262 488332 228318
rect 487508 225894 487564 225950
rect 490484 234182 490540 234238
rect 495092 233146 495148 233202
rect 494228 228558 494284 228614
rect 493460 227226 493516 227282
rect 497972 228410 498028 228466
rect 498836 227078 498892 227134
rect 518420 222934 518476 222990
rect 519860 222638 519916 222694
rect 522932 222490 522988 222546
rect 524468 222786 524524 222842
rect 527540 230038 527596 230094
rect 526004 224562 526060 224618
rect 526676 224414 526732 224470
rect 528308 228706 528364 228762
rect 528980 224266 529036 224322
rect 530516 224118 530572 224174
rect 532052 223970 532108 224026
rect 538004 238030 538060 238086
rect 534260 230186 534316 230242
rect 536564 223822 536620 223878
rect 540308 229890 540364 229946
rect 544340 238326 544396 238382
rect 544052 223674 544108 223730
rect 550196 238622 550252 238678
rect 549428 232998 549484 233054
rect 555380 238918 555436 238974
rect 551636 232850 551692 232906
rect 553940 229742 553996 229798
rect 559892 238178 559948 238234
rect 559220 236550 559276 236606
rect 557684 236402 557740 236458
rect 557588 232702 557644 232758
rect 565268 236698 565324 236754
rect 560756 232554 560812 232610
rect 562964 223526 563020 223582
rect 562196 223378 562252 223434
rect 581780 238770 581836 238826
rect 573140 236994 573196 237050
rect 567476 236846 567532 236902
rect 570452 232406 570508 232462
rect 569780 229594 569836 229650
rect 571316 223230 571372 223286
rect 572756 229446 572812 229502
rect 573524 229298 573580 229354
rect 580340 235958 580396 236014
rect 576596 232258 576652 232314
rect 575828 231962 575884 232018
rect 575060 230334 575116 230390
rect 578036 232110 578092 232166
rect 577268 223082 577324 223138
rect 578900 229150 578956 229206
rect 591476 236106 591532 236162
rect 587924 235810 587980 235866
rect 587444 234330 587500 234386
rect 590708 235662 590764 235718
rect 590900 234478 590956 234534
rect 590900 226782 590956 226838
rect 591668 226930 591724 226986
rect 599924 229002 599980 229058
rect 596180 226634 596236 226690
rect 596948 226486 597004 226542
rect 604532 231814 604588 231870
rect 627188 240102 627244 240158
rect 621140 236254 621196 236310
rect 608276 235514 608332 235570
rect 607508 228854 607564 228910
rect 611252 235366 611308 235422
rect 614324 235218 614380 235274
rect 618836 235070 618892 235126
rect 616628 234922 616684 234978
rect 617300 226338 617356 226394
rect 619604 234774 619660 234830
rect 620372 226190 620428 226246
rect 623348 226042 623404 226098
rect 625556 234626 625612 234682
rect 640148 212278 640204 212334
rect 640148 211538 640204 211594
rect 190292 201326 190348 201382
rect 640148 200882 640204 200938
rect 190292 200512 190348 200568
rect 640148 200142 640204 200198
rect 187220 199106 187276 199162
rect 640244 185638 640300 185694
rect 640244 184898 640300 184954
rect 645140 182974 645196 183030
rect 186260 182382 186316 182438
rect 645140 179274 645196 179330
rect 645140 174873 645142 174890
rect 645142 174873 645194 174890
rect 645194 174873 645196 174890
rect 645140 174834 645196 174873
rect 645140 171025 645142 171042
rect 645142 171025 645194 171042
rect 645194 171025 645196 171042
rect 645140 170986 645196 171025
rect 645140 167730 645196 167786
rect 645140 163329 645142 163346
rect 645142 163329 645194 163346
rect 645194 163329 645196 163346
rect 645140 163290 645196 163329
rect 645140 159442 645196 159498
rect 645140 155446 645196 155502
rect 645140 152525 645142 152542
rect 645142 152525 645194 152542
rect 645194 152525 645196 152542
rect 645140 152486 645196 152525
rect 645140 148046 645196 148102
rect 186740 145826 186796 145882
rect 186164 137390 186220 137446
rect 186260 135170 186316 135226
rect 648596 272070 648652 272126
rect 647348 269258 647404 269314
rect 646676 144198 646732 144254
rect 655220 778230 655276 778286
rect 654164 774826 654220 774882
rect 654836 772310 654892 772366
rect 655124 734422 655180 734478
rect 654164 730278 654220 730334
rect 654260 729094 654316 729150
rect 654164 727910 654220 727966
rect 654452 683510 654508 683566
rect 655604 777638 655660 777694
rect 655412 775862 655468 775918
rect 655316 731610 655372 731666
rect 655220 689430 655276 689486
rect 649748 263338 649804 263394
rect 646772 140942 646828 140998
rect 650420 275622 650476 275678
rect 655124 642958 655180 643014
rect 654164 640590 654220 640646
rect 654548 595302 654604 595358
rect 654164 593395 654220 593434
rect 654164 593378 654166 593395
rect 654166 593378 654218 593395
rect 654218 593378 654220 593395
rect 654356 591898 654412 591954
rect 655508 732646 655564 732702
rect 655412 688394 655468 688450
rect 655316 642366 655372 642422
rect 655220 597818 655276 597874
rect 655124 553270 655180 553326
rect 653780 550902 653836 550958
rect 654164 547498 654220 547554
rect 656180 773494 656236 773550
rect 655604 687062 655660 687118
rect 655508 640738 655564 640794
rect 655412 596634 655468 596690
rect 655316 552086 655372 552142
rect 656372 685878 656428 685934
rect 655988 684694 656044 684750
rect 655796 638222 655852 638278
rect 655892 637038 655948 637094
rect 655604 595450 655660 595506
rect 655508 551050 655564 551106
rect 656276 548534 656332 548590
rect 655124 374338 655180 374394
rect 655508 373302 655564 373358
rect 655316 372118 655372 372174
rect 654164 370934 654220 370990
rect 655220 329790 655276 329846
rect 655124 328014 655180 328070
rect 655316 327422 655372 327478
rect 654164 326238 654220 326294
rect 653780 303298 653836 303354
rect 654068 302114 654124 302170
rect 654164 300930 654220 300986
rect 656564 298710 656620 298766
rect 656372 297526 656428 297582
rect 656180 296786 656236 296842
rect 656084 295158 656140 295214
rect 655892 293974 655948 294030
rect 655796 292790 655852 292846
rect 655604 290866 655660 290922
rect 654164 289238 654220 289294
rect 655412 288054 655468 288110
rect 653780 284502 653836 284558
rect 655124 283318 655180 283374
rect 654740 279766 654796 279822
rect 647060 134726 647116 134782
rect 647732 130878 647788 130934
rect 646964 127622 647020 127678
rect 646868 125698 646924 125754
rect 646580 123774 646636 123830
rect 646484 121998 646540 122054
rect 185684 110158 185740 110214
rect 185300 109309 185302 109326
rect 185302 109309 185354 109326
rect 185354 109309 185356 109326
rect 185300 109270 185356 109309
rect 646196 117558 646252 117614
rect 647924 128954 647980 129010
rect 655316 282282 655372 282338
rect 655220 280950 655276 281006
rect 655508 286870 655564 286926
rect 655700 285686 655756 285742
rect 655988 291606 656044 291662
rect 647828 119482 647884 119538
rect 647924 115634 647980 115690
rect 668180 277842 668236 277898
rect 646580 113118 646636 113174
rect 186260 108678 186316 108734
rect 186644 106310 186700 106366
rect 645908 106014 645964 106070
rect 184724 102462 184780 102518
rect 645140 102166 645196 102222
rect 184628 98022 184684 98078
rect 184340 97134 184396 97190
rect 184436 96394 184492 96450
rect 184532 95654 184588 95710
rect 184340 94805 184342 94822
rect 184342 94805 184394 94822
rect 184394 94805 184396 94822
rect 184340 94766 184396 94805
rect 184436 93434 184492 93490
rect 184628 94174 184684 94230
rect 184532 92694 184588 92750
rect 184340 91971 184396 92010
rect 184340 91954 184342 91971
rect 184342 91954 184394 91971
rect 184394 91954 184396 91971
rect 184436 90326 184492 90382
rect 184628 91066 184684 91122
rect 184532 89586 184588 89642
rect 184340 88846 184396 88902
rect 184436 88106 184492 88162
rect 184532 87218 184588 87274
rect 184628 86626 184684 86682
rect 184340 85738 184396 85794
rect 184532 85146 184588 85202
rect 184436 84258 184492 84314
rect 184340 83409 184342 83426
rect 184342 83409 184394 83426
rect 184394 83409 184396 83426
rect 184340 83370 184396 83409
rect 184244 81890 184300 81946
rect 186164 82778 186220 82834
rect 184436 81298 184492 81354
rect 184436 79818 184492 79874
rect 184340 78930 184396 78986
rect 184628 80427 184684 80466
rect 184628 80410 184630 80427
rect 184630 80410 184682 80427
rect 184682 80410 184684 80427
rect 184532 78190 184588 78246
rect 184436 77450 184492 77506
rect 184340 76710 184396 76766
rect 184628 75970 184684 76026
rect 184532 75082 184588 75138
rect 184340 74342 184396 74398
rect 184532 73602 184588 73658
rect 184436 72862 184492 72918
rect 184628 72122 184684 72178
rect 184340 71382 184396 71438
rect 149492 70790 149548 70846
rect 149396 69458 149452 69514
rect 149204 68274 149260 68330
rect 184436 70494 184492 70550
rect 184532 69902 184588 69958
rect 184340 69053 184342 69070
rect 184342 69053 184394 69070
rect 184394 69053 184396 69070
rect 184340 69014 184396 69053
rect 184436 68422 184492 68478
rect 184340 67534 184396 67590
rect 149588 67090 149644 67146
rect 149492 65314 149548 65370
rect 149396 64574 149452 64630
rect 149300 63390 149356 63446
rect 184532 66794 184588 66850
rect 184340 66054 184396 66110
rect 184532 65166 184588 65222
rect 184628 64574 184684 64630
rect 184436 63686 184492 63742
rect 184340 63111 184396 63150
rect 184340 63094 184342 63111
rect 184342 63094 184394 63111
rect 184394 63094 184396 63111
rect 149492 62206 149548 62262
rect 184436 62206 184492 62262
rect 149396 60578 149452 60634
rect 184532 61466 184588 61522
rect 184628 60726 184684 60782
rect 184340 59986 184396 60042
rect 149396 59690 149452 59746
rect 184436 59246 184492 59302
rect 149396 58506 149452 58562
rect 184532 58358 184588 58414
rect 184340 57618 184396 57674
rect 149492 57322 149548 57378
rect 149396 56177 149398 56194
rect 149398 56177 149450 56194
rect 149450 56177 149452 56194
rect 149396 56138 149452 56177
rect 184340 56878 184396 56934
rect 184340 56155 184396 56194
rect 184340 56138 184342 56155
rect 184342 56138 184394 56155
rect 184394 56138 184396 56155
rect 184436 55398 184492 55454
rect 149684 54806 149740 54862
rect 184340 54675 184396 54714
rect 184340 54658 184342 54675
rect 184342 54658 184394 54675
rect 184394 54658 184396 54675
rect 184340 53918 184396 53974
rect 149396 53770 149452 53826
rect 142100 40154 142156 40210
rect 426164 44890 426220 44946
rect 415220 41930 415276 41986
rect 416852 41782 416908 41838
rect 420788 40450 420844 40506
rect 311060 37194 311116 37250
rect 328340 37194 328396 37250
rect 472244 44890 472300 44946
rect 464852 41782 464908 41838
rect 470324 41782 470380 41838
rect 512180 41782 512236 41838
rect 525908 41782 525964 41838
rect 645428 95967 645484 96006
rect 645428 95950 645430 95967
rect 645430 95950 645482 95967
rect 645482 95950 645484 95967
rect 645908 88846 645964 88902
rect 645908 84406 645964 84462
rect 645524 79374 645580 79430
rect 646004 75526 646060 75582
rect 646004 66219 646060 66258
rect 646004 66202 646006 66219
rect 646006 66202 646058 66219
rect 646058 66202 646060 66219
rect 646004 58950 646060 59006
rect 647156 111342 647212 111398
rect 646676 109418 646732 109474
rect 646772 107938 646828 107994
rect 646964 98022 647020 98078
rect 669524 275326 669580 275382
rect 669716 275178 669772 275234
rect 669908 277398 669964 277454
rect 670484 348586 670540 348642
rect 670292 278286 670348 278342
rect 670484 278138 670540 278194
rect 670100 277546 670156 277602
rect 676244 877259 676300 877298
rect 676244 877242 676246 877259
rect 676246 877242 676298 877259
rect 676298 877242 676300 877259
rect 676244 876223 676300 876262
rect 676244 876206 676246 876223
rect 676246 876206 676298 876223
rect 676298 876206 676300 876223
rect 680276 875614 680332 875670
rect 676052 875466 676108 875522
rect 679796 875022 679852 875078
rect 676244 873690 676300 873746
rect 679700 872654 679756 872710
rect 676052 871470 676108 871526
rect 676244 870730 676300 870786
rect 676052 869990 676108 870046
rect 680180 874134 680236 874190
rect 679892 872062 679948 872118
rect 676244 869250 676300 869306
rect 679796 868658 679852 868714
rect 679796 868214 679852 868270
rect 680084 871618 680140 871674
rect 679988 870138 680044 870194
rect 685460 868214 685516 868270
rect 685460 867770 685516 867826
rect 675188 852526 675244 852582
rect 675476 774530 675532 774586
rect 675380 773642 675436 773698
rect 675764 773050 675820 773106
rect 675764 770682 675820 770738
rect 675476 769942 675532 769998
rect 675476 769350 675532 769406
rect 674516 731610 674572 731666
rect 674324 676850 674380 676906
rect 675476 729834 675532 729890
rect 675764 729390 675820 729446
rect 675668 728650 675724 728706
rect 675380 726726 675436 726782
rect 675764 726134 675820 726190
rect 675380 725838 675436 725894
rect 675764 721842 675820 721898
rect 676244 703063 676300 703102
rect 676244 703046 676246 703063
rect 676246 703046 676298 703063
rect 676298 703046 676300 703063
rect 676244 702915 676300 702954
rect 676244 702898 676246 702915
rect 676246 702898 676298 702915
rect 676298 702898 676300 702915
rect 676052 702158 676108 702214
rect 679700 701566 679756 701622
rect 676244 700843 676300 700882
rect 676244 700826 676246 700843
rect 676246 700826 676298 700843
rect 676298 700826 676300 700843
rect 679700 700826 679756 700882
rect 676244 700103 676300 700142
rect 676244 700086 676246 700103
rect 676246 700086 676298 700103
rect 676298 700086 676300 700103
rect 676052 699733 676108 699772
rect 676052 699716 676054 699733
rect 676054 699716 676106 699733
rect 676106 699716 676108 699733
rect 676052 699198 676108 699254
rect 676052 698162 676108 698218
rect 676244 697422 676300 697478
rect 675956 696682 676012 696738
rect 676052 696164 676108 696220
rect 676244 694462 676300 694518
rect 676052 693722 676108 693778
rect 676052 692760 676108 692816
rect 679988 691502 680044 691558
rect 679796 690910 679852 690966
rect 679988 690910 680044 690966
rect 679796 690466 679852 690522
rect 675380 685582 675436 685638
rect 675764 684398 675820 684454
rect 675572 682622 675628 682678
rect 675764 678330 675820 678386
rect 675476 673298 675532 673354
rect 675284 671374 675340 671430
rect 676148 658794 676204 658850
rect 676052 657575 676054 657592
rect 676054 657575 676106 657592
rect 676106 657575 676108 657592
rect 676052 657536 676108 657575
rect 676340 658202 676396 658258
rect 676244 657758 676300 657814
rect 676052 657018 676108 657074
rect 676052 656465 676054 656482
rect 676054 656465 676106 656482
rect 676106 656465 676108 656482
rect 676052 656426 676108 656465
rect 676052 656073 676108 656112
rect 676052 656056 676054 656073
rect 676054 656056 676106 656073
rect 676106 656056 676108 656073
rect 676244 655725 676246 655742
rect 676246 655725 676298 655742
rect 676298 655725 676300 655742
rect 676244 655686 676300 655725
rect 676244 654815 676300 654854
rect 676244 654798 676246 654815
rect 676246 654798 676298 654815
rect 676298 654798 676300 654815
rect 675572 654058 675628 654114
rect 676052 652504 676108 652560
rect 675476 651986 675532 652042
rect 676052 650062 676108 650118
rect 676244 649213 676246 649230
rect 676246 649213 676298 649230
rect 676298 649213 676300 649230
rect 676244 649174 676300 649213
rect 676052 648029 676054 648046
rect 676054 648029 676106 648046
rect 676106 648029 676108 648046
rect 676052 647990 676108 648029
rect 679796 647250 679852 647306
rect 679796 646806 679852 646862
rect 685460 646806 685516 646862
rect 685460 646362 685516 646418
rect 675764 641626 675820 641682
rect 675476 640294 675532 640350
rect 675188 640146 675244 640202
rect 675476 638370 675532 638426
rect 675380 634078 675436 634134
rect 675764 632746 675820 632802
rect 675764 629046 675820 629102
rect 675764 627270 675820 627326
rect 676148 614394 676204 614450
rect 676052 614098 676108 614154
rect 676244 613802 676300 613858
rect 676052 613175 676054 613192
rect 676054 613175 676106 613192
rect 676106 613175 676108 613192
rect 676052 613136 676108 613175
rect 676052 612635 676108 612674
rect 676052 612618 676054 612635
rect 676054 612618 676106 612635
rect 676106 612618 676108 612635
rect 676244 611895 676300 611934
rect 676244 611878 676246 611895
rect 676246 611878 676298 611895
rect 676298 611878 676300 611895
rect 676052 611673 676108 611712
rect 676052 611656 676054 611673
rect 676054 611656 676106 611673
rect 676106 611656 676108 611673
rect 676052 611155 676108 611194
rect 676052 611138 676054 611155
rect 676054 611138 676106 611155
rect 676106 611138 676108 611155
rect 676052 610585 676054 610602
rect 676054 610585 676106 610602
rect 676106 610585 676108 610602
rect 676052 610546 676108 610585
rect 676052 607181 676054 607198
rect 676054 607181 676106 607198
rect 676106 607181 676108 607198
rect 676052 607142 676108 607181
rect 676052 606663 676054 606680
rect 676054 606663 676106 606680
rect 676106 606663 676108 606680
rect 676052 606624 676108 606663
rect 676244 606293 676246 606310
rect 676246 606293 676298 606310
rect 676298 606293 676300 606310
rect 676244 606254 676300 606293
rect 676052 605701 676054 605718
rect 676054 605701 676106 605718
rect 676106 605701 676108 605718
rect 676052 605662 676108 605701
rect 676052 605109 676054 605126
rect 676054 605109 676106 605126
rect 676106 605109 676108 605126
rect 676052 605070 676108 605109
rect 676052 604665 676054 604682
rect 676054 604665 676106 604682
rect 676106 604665 676108 604682
rect 676052 604626 676108 604665
rect 676244 604369 676246 604386
rect 676246 604369 676298 604386
rect 676298 604369 676300 604386
rect 676244 604330 676300 604369
rect 676052 603629 676054 603646
rect 676054 603629 676106 603646
rect 676106 603629 676108 603646
rect 676052 603590 676108 603629
rect 679988 602850 680044 602906
rect 679796 602406 679852 602462
rect 679988 602406 680044 602462
rect 679796 601962 679852 602018
rect 675380 597078 675436 597134
rect 675476 596042 675532 596098
rect 675476 593970 675532 594026
rect 675476 589678 675532 589734
rect 675764 584646 675820 584702
rect 675668 582870 675724 582926
rect 676244 569254 676300 569310
rect 676148 568514 676204 568570
rect 676052 568366 676108 568422
rect 676052 567443 676054 567460
rect 676054 567443 676106 567460
rect 676106 567443 676108 567460
rect 676052 567404 676108 567443
rect 679700 567774 679756 567830
rect 674900 567182 674956 567238
rect 676244 567073 676246 567090
rect 676246 567073 676298 567090
rect 676298 567073 676300 567090
rect 676244 567034 676300 567073
rect 676244 566311 676300 566350
rect 676244 566294 676246 566311
rect 676246 566294 676298 566311
rect 676298 566294 676300 566311
rect 676052 565889 676054 565906
rect 676054 565889 676106 565906
rect 676106 565889 676108 565906
rect 676052 565850 676108 565889
rect 676052 565423 676108 565462
rect 676052 565406 676054 565423
rect 676054 565406 676106 565423
rect 676106 565406 676108 565423
rect 676052 561449 676054 561466
rect 676054 561449 676106 561466
rect 676106 561449 676108 561466
rect 676052 561410 676108 561449
rect 676052 560857 676054 560874
rect 676054 560857 676106 560874
rect 676106 560857 676108 560874
rect 676052 560818 676108 560857
rect 676244 560709 676246 560726
rect 676246 560709 676298 560726
rect 676298 560709 676300 560726
rect 676244 560670 676300 560709
rect 676052 559377 676054 559394
rect 676054 559377 676106 559394
rect 676106 559377 676108 559394
rect 676052 559338 676108 559377
rect 676052 559007 676054 559024
rect 676054 559007 676106 559024
rect 676106 559007 676108 559024
rect 676052 558968 676108 559007
rect 676244 558637 676246 558654
rect 676246 558637 676298 558654
rect 676298 558637 676300 558654
rect 676244 558598 676300 558637
rect 679796 557710 679852 557766
rect 679796 557118 679852 557174
rect 685460 557118 685516 557174
rect 685460 556674 685516 556730
rect 675476 552974 675532 553030
rect 675380 552234 675436 552290
rect 675188 551642 675244 551698
rect 675284 550162 675340 550218
rect 675380 545426 675436 545482
rect 675380 544242 675436 544298
rect 675764 540542 675820 540598
rect 675188 538618 675244 538674
rect 676340 525150 676396 525206
rect 676148 524706 676204 524762
rect 676244 524575 676300 524614
rect 676244 524558 676246 524575
rect 676246 524558 676298 524575
rect 676298 524558 676300 524575
rect 676052 524005 676054 524022
rect 676054 524005 676106 524022
rect 676106 524005 676108 524022
rect 676052 523966 676108 524005
rect 676532 523226 676588 523282
rect 676052 522856 676108 522912
rect 676244 521746 676300 521802
rect 676244 517641 676246 517658
rect 676246 517641 676298 517658
rect 676298 517641 676300 517658
rect 676244 517602 676300 517641
rect 676052 516901 676054 516918
rect 676054 516901 676106 516918
rect 676106 516901 676108 516918
rect 676052 516862 676108 516901
rect 676052 516457 676054 516474
rect 676054 516457 676106 516474
rect 676106 516457 676108 516474
rect 676052 516418 676108 516457
rect 676244 516161 676246 516178
rect 676246 516161 676298 516178
rect 676298 516161 676300 516178
rect 676244 516122 676300 516161
rect 676052 515421 676054 515438
rect 676054 515421 676106 515438
rect 676106 515421 676108 515438
rect 676052 515382 676108 515421
rect 676052 514977 676054 514994
rect 676054 514977 676106 514994
rect 676106 514977 676108 514994
rect 676052 514938 676108 514977
rect 676052 514459 676054 514476
rect 676054 514459 676106 514476
rect 676106 514459 676108 514476
rect 676052 514420 676108 514459
rect 676340 482378 676396 482434
rect 676148 481786 676204 481842
rect 676244 481359 676300 481398
rect 676244 481342 676246 481359
rect 676246 481342 676298 481359
rect 676298 481342 676300 481359
rect 676628 522190 676684 522246
rect 676724 521154 676780 521210
rect 679988 514050 680044 514106
rect 679796 513162 679852 513218
rect 679988 513162 680044 513218
rect 679796 512718 679852 512774
rect 676532 481342 676588 481398
rect 676436 480306 676492 480362
rect 676052 479640 676108 479696
rect 676724 480306 676780 480362
rect 676628 479270 676684 479326
rect 676244 478399 676300 478438
rect 676244 478382 676246 478399
rect 676246 478382 676298 478399
rect 676298 478382 676300 478399
rect 676052 475570 676108 475626
rect 676052 474647 676054 474664
rect 676054 474647 676106 474664
rect 676106 474647 676108 474664
rect 676052 474608 676108 474647
rect 676244 474277 676246 474294
rect 676246 474277 676298 474294
rect 676298 474277 676300 474294
rect 676244 474238 676300 474277
rect 676244 472797 676246 472814
rect 676246 472797 676298 472814
rect 676298 472797 676300 472814
rect 676244 472758 676300 472797
rect 676052 472205 676054 472222
rect 676054 472205 676106 472222
rect 676106 472205 676108 472222
rect 676052 472166 676108 472205
rect 676052 471613 676054 471630
rect 676054 471613 676106 471630
rect 676106 471613 676108 471630
rect 676052 471574 676108 471613
rect 672500 278434 672556 278490
rect 672404 276214 672460 276270
rect 676148 396390 676204 396446
rect 676340 395798 676396 395854
rect 676244 395354 676300 395410
rect 679796 470834 679852 470890
rect 679796 470390 679852 470446
rect 685460 470390 685516 470446
rect 685460 469946 685516 470002
rect 676724 395354 676780 395410
rect 676244 393891 676300 393930
rect 676244 393874 676246 393891
rect 676246 393874 676298 393891
rect 676298 393874 676300 393891
rect 675860 393173 675862 393190
rect 675862 393173 675914 393190
rect 675914 393173 675916 393190
rect 675860 393134 675916 393173
rect 675572 391062 675628 391118
rect 676244 391950 676300 392006
rect 676244 390470 676300 390526
rect 676052 390100 676108 390156
rect 676052 389582 676108 389638
rect 676244 388990 676300 389046
rect 676052 388620 676108 388676
rect 675956 388102 676012 388158
rect 676244 387510 676300 387566
rect 676244 386918 676300 386974
rect 676052 386622 676108 386678
rect 675956 386178 676012 386234
rect 676244 385438 676300 385494
rect 679700 384846 679756 384902
rect 679700 384402 679756 384458
rect 685460 384402 685516 384458
rect 685460 383958 685516 384014
rect 675476 367234 675532 367290
rect 676244 351694 676300 351750
rect 676052 351585 676054 351602
rect 676054 351585 676106 351602
rect 676106 351585 676108 351602
rect 676052 351546 676108 351585
rect 676052 350954 676108 351010
rect 677012 346810 677068 346866
rect 676052 346514 676108 346570
rect 676916 344738 676972 344794
rect 676052 344590 676108 344646
rect 676244 343850 676300 343906
rect 676820 342814 676876 342870
rect 676052 342518 676108 342574
rect 675956 341556 676012 341612
rect 676244 341778 676300 341834
rect 676052 341038 676108 341094
rect 676820 339706 676876 339762
rect 676916 339262 676972 339318
rect 679988 340298 680044 340354
rect 679796 339706 679852 339762
rect 679988 339706 680044 339762
rect 679796 339262 679852 339318
rect 677012 338818 677068 338874
rect 675380 333934 675436 333990
rect 675476 332306 675532 332362
rect 675380 331122 675436 331178
rect 675380 327866 675436 327922
rect 675668 324906 675724 324962
rect 675764 322982 675820 323038
rect 675764 321206 675820 321262
rect 679892 313954 679948 314010
rect 676244 305666 676300 305722
rect 676244 305239 676300 305278
rect 676244 305222 676246 305239
rect 676246 305222 676298 305239
rect 676298 305222 676300 305239
rect 676244 304778 676300 304834
rect 679892 304778 679948 304834
rect 676052 304055 676108 304094
rect 676052 304038 676054 304055
rect 676054 304038 676106 304055
rect 676106 304038 676108 304055
rect 672692 303446 672748 303502
rect 672884 302558 672940 302614
rect 672692 277990 672748 278046
rect 672884 277694 672940 277750
rect 673268 276362 673324 276418
rect 673172 276066 673228 276122
rect 672596 271478 672652 271534
rect 670004 270590 670060 270646
rect 672404 266890 672460 266946
rect 669620 263486 669676 263542
rect 672596 266742 672652 266798
rect 672404 170986 672460 171042
rect 676052 303019 676108 303058
rect 676052 303002 676054 303019
rect 676054 303002 676106 303019
rect 676106 303002 676108 303019
rect 676052 301983 676108 302022
rect 676052 301966 676054 301983
rect 676054 301966 676106 301983
rect 676106 301966 676108 301983
rect 676052 298562 676108 298618
rect 676052 295972 676108 296028
rect 679892 294270 679948 294326
rect 679700 293826 679756 293882
rect 679892 293826 679948 293882
rect 679700 293234 679756 293290
rect 675764 290570 675820 290626
rect 675764 289682 675820 289738
rect 675764 287906 675820 287962
rect 675764 287462 675820 287518
rect 675380 286870 675436 286926
rect 675380 283762 675436 283818
rect 675572 282874 675628 282930
rect 675668 281838 675724 281894
rect 675572 281690 675628 281746
rect 675380 280654 675436 280710
rect 675380 278878 675436 278934
rect 675380 276954 675436 277010
rect 679892 275030 679948 275086
rect 676244 262746 676300 262802
rect 676052 262467 676108 262506
rect 676052 262450 676054 262467
rect 676054 262450 676106 262467
rect 676106 262450 676108 262467
rect 676244 261710 676300 261766
rect 676052 261601 676054 261618
rect 676054 261601 676106 261618
rect 676106 261601 676108 261618
rect 676052 261562 676108 261601
rect 679700 260822 679756 260878
rect 679796 259786 679852 259842
rect 679700 258750 679756 258806
rect 676052 258602 676108 258658
rect 675764 257418 675820 257474
rect 676916 255790 676972 255846
rect 676052 255568 676108 255624
rect 675956 255050 676012 255106
rect 676244 254310 676300 254366
rect 676820 253866 676876 253922
rect 676052 252978 676108 253034
rect 675956 252016 676012 252072
rect 676244 252386 676300 252442
rect 679988 251646 680044 251702
rect 679796 250758 679852 250814
rect 679988 250758 680044 250814
rect 679796 250314 679852 250370
rect 679700 249278 679756 249334
rect 676916 247946 676972 248002
rect 676820 247798 676876 247854
rect 675668 243654 675724 243710
rect 675380 239066 675436 239122
rect 675764 238030 675820 238086
rect 675764 235958 675820 236014
rect 675380 234478 675436 234534
rect 675764 232554 675820 232610
rect 676244 219678 676300 219734
rect 676244 219251 676300 219290
rect 676244 219234 676246 219251
rect 676246 219234 676298 219251
rect 676298 219234 676300 219251
rect 676052 218938 676108 218994
rect 676244 215386 676300 215442
rect 675572 214498 675628 214554
rect 675284 212574 675340 212630
rect 676052 214054 676108 214110
rect 676916 212722 676972 212778
rect 676244 211834 676300 211890
rect 676052 211464 676108 211520
rect 676820 210798 676876 210854
rect 676052 209984 676108 210040
rect 675956 209614 676012 209670
rect 679892 208282 679948 208338
rect 679892 207838 679948 207894
rect 679796 207690 679852 207746
rect 679796 207246 679852 207302
rect 676916 204730 676972 204786
rect 676820 204582 676876 204638
rect 675476 195110 675532 195166
rect 675380 193926 675436 193982
rect 675476 193038 675532 193094
rect 675764 192150 675820 192206
rect 675476 189930 675532 189986
rect 675764 188450 675820 188506
rect 676148 173798 676204 173854
rect 676052 173502 676108 173558
rect 676244 173223 676300 173262
rect 676244 173206 676246 173223
rect 676246 173206 676298 173223
rect 676298 173206 676300 173223
rect 676052 169967 676108 170006
rect 676052 169950 676054 169967
rect 676054 169950 676106 169967
rect 676106 169950 676108 169967
rect 676052 169079 676108 169118
rect 676052 169062 676054 169079
rect 676054 169062 676106 169079
rect 676106 169062 676108 169079
rect 676052 164030 676108 164086
rect 676244 162254 676300 162310
rect 676148 161810 676204 161866
rect 676244 161405 676246 161422
rect 676246 161405 676298 161422
rect 676298 161405 676300 161422
rect 676244 161366 676300 161405
rect 675764 158110 675820 158166
rect 675764 157666 675820 157722
rect 675764 156926 675820 156982
rect 675476 155150 675532 155206
rect 675380 154410 675436 154466
rect 675764 153818 675820 153874
rect 675188 152634 675244 152690
rect 675380 150858 675436 150914
rect 675476 150266 675532 150322
rect 675380 149526 675436 149582
rect 675380 147898 675436 147954
rect 675476 143902 675532 143958
rect 676244 129585 676246 129602
rect 676246 129585 676298 129602
rect 676298 129585 676300 129602
rect 676244 129546 676300 129585
rect 676340 129102 676396 129158
rect 676244 128510 676300 128566
rect 676148 127474 676204 127530
rect 676052 126882 676108 126938
rect 676052 126329 676054 126346
rect 676054 126329 676106 126346
rect 676106 126329 676108 126346
rect 676052 126290 676108 126329
rect 676244 125550 676300 125606
rect 676052 124218 676108 124274
rect 668180 106310 668236 106366
rect 665588 105274 665644 105330
rect 665300 105126 665356 105182
rect 676820 124514 676876 124570
rect 676052 122368 676108 122424
rect 675956 121850 676012 121906
rect 676244 121127 676300 121166
rect 676244 121110 676246 121127
rect 676246 121110 676298 121127
rect 676298 121110 676300 121127
rect 676052 120370 676108 120426
rect 676052 119778 676108 119834
rect 675956 118816 676012 118872
rect 676244 119186 676300 119242
rect 676244 118463 676300 118502
rect 676244 118446 676246 118463
rect 676246 118446 676298 118463
rect 676298 118446 676300 118463
rect 676148 117706 676204 117762
rect 676244 117114 676300 117170
rect 679700 122590 679756 122646
rect 676820 115634 676876 115690
rect 679700 115190 679756 115246
rect 675572 112082 675628 112138
rect 675764 110898 675820 110954
rect 675380 106458 675436 106514
rect 647924 104090 647980 104146
rect 647924 99650 647980 99706
rect 647828 94026 647884 94082
rect 647732 92694 647788 92750
rect 647924 87070 647980 87126
rect 650900 86182 650956 86238
rect 652340 85294 652396 85350
rect 651764 84258 651820 84314
rect 652244 83370 652300 83426
rect 647924 82630 647980 82686
rect 647924 81002 647980 81058
rect 647924 77489 647926 77506
rect 647926 77489 647978 77506
rect 647978 77489 647980 77506
rect 647924 77450 647980 77489
rect 647060 71826 647116 71882
rect 646868 68570 646924 68626
rect 647924 73602 647980 73658
rect 647924 69623 647980 69662
rect 647924 69606 647926 69623
rect 647926 69606 647978 69623
rect 647978 69606 647980 69623
rect 647924 64130 647980 64186
rect 647924 62206 647980 62262
rect 647156 60282 647212 60338
rect 659348 90770 659404 90826
rect 675668 103498 675724 103554
rect 675764 101574 675820 101630
rect 675764 99798 675820 99854
rect 653684 86922 653740 86978
rect 663284 86330 663340 86386
rect 652436 82630 652492 82686
rect 662420 81611 662476 81650
rect 662420 81594 662422 81611
rect 662422 81594 662474 81611
rect 662474 81594 662476 81611
rect 663284 84702 663340 84758
rect 663380 83962 663436 84018
rect 663284 82038 663340 82094
rect 663476 82778 663532 82834
rect 646772 57026 646828 57082
rect 646484 54658 646540 54714
rect 539732 40450 539788 40506
<< metal3 >>
rect 175599 997772 175665 997775
rect 486735 997772 486801 997775
rect 538575 997772 538641 997775
rect 639375 997772 639441 997775
rect 175599 997770 176352 997772
rect 80514 997183 80574 997742
rect 129474 997183 129534 997742
rect 175599 997714 175604 997770
rect 175660 997714 176352 997770
rect 485856 997770 486801 997772
rect 175599 997712 176352 997714
rect 175599 997709 175665 997712
rect 80514 997178 80625 997183
rect 80514 997122 80564 997178
rect 80620 997122 80625 997178
rect 80514 997120 80625 997122
rect 129474 997178 129585 997183
rect 129474 997122 129524 997178
rect 129580 997122 129585 997178
rect 129474 997120 129585 997122
rect 80559 997117 80625 997120
rect 129519 997117 129585 997120
rect 238959 997180 239025 997183
rect 239874 997180 239934 997742
rect 238959 997178 239934 997180
rect 238959 997122 238964 997178
rect 239020 997122 239934 997178
rect 238959 997120 239934 997122
rect 293058 997183 293118 997742
rect 432066 997183 432126 997742
rect 485856 997714 486740 997770
rect 486796 997714 486801 997770
rect 485856 997712 486801 997714
rect 535584 997770 538641 997772
rect 535584 997714 538580 997770
rect 538636 997714 538641 997770
rect 535584 997712 538641 997714
rect 636768 997770 639441 997772
rect 636768 997714 639380 997770
rect 639436 997714 639441 997770
rect 636768 997712 639441 997714
rect 486735 997709 486801 997712
rect 538575 997709 538641 997712
rect 639375 997709 639441 997712
rect 293058 997178 293169 997183
rect 293058 997122 293108 997178
rect 293164 997122 293169 997178
rect 293058 997120 293169 997122
rect 238959 997117 239025 997120
rect 293103 997117 293169 997120
rect 432015 997178 432126 997183
rect 432015 997122 432020 997178
rect 432076 997122 432126 997178
rect 432015 997120 432126 997122
rect 432015 997117 432081 997120
rect 238959 983120 239025 983123
rect 287919 983120 287985 983123
rect 238959 983118 241278 983120
rect 238959 983062 238964 983118
rect 239020 983062 241278 983118
rect 238959 983060 241278 983062
rect 238959 983057 239025 983060
rect 80559 982972 80625 982975
rect 132399 982972 132465 982975
rect 184239 982972 184305 982975
rect 233199 982972 233265 982975
rect 239919 982972 239985 982975
rect 80559 982970 81726 982972
rect 80559 982914 80564 982970
rect 80620 982914 81726 982970
rect 80559 982912 81726 982914
rect 80559 982909 80625 982912
rect 81666 982646 81726 982912
rect 132399 982970 133566 982972
rect 132399 982914 132404 982970
rect 132460 982914 133566 982970
rect 132399 982912 133566 982914
rect 132399 982909 132465 982912
rect 133506 982646 133566 982912
rect 184239 982970 185598 982972
rect 184239 982914 184244 982970
rect 184300 982914 185598 982970
rect 184239 982912 185598 982914
rect 184239 982909 184305 982912
rect 185538 982646 185598 982912
rect 233199 982970 236286 982972
rect 233199 982914 233204 982970
rect 233260 982914 236286 982970
rect 233199 982912 236286 982914
rect 233199 982909 233265 982912
rect 236226 982646 236286 982912
rect 239874 982970 239985 982972
rect 239874 982914 239924 982970
rect 239980 982914 239985 982970
rect 239874 982909 239985 982914
rect 239874 982646 239934 982909
rect 241218 982646 241278 983060
rect 287919 983118 290622 983120
rect 287919 983062 287924 983118
rect 287980 983062 290622 983118
rect 287919 983060 290622 983062
rect 287919 983057 287985 983060
rect 285039 982972 285105 982975
rect 285039 982970 288126 982972
rect 285039 982914 285044 982970
rect 285100 982914 288126 982970
rect 285039 982912 288126 982914
rect 285039 982909 285105 982912
rect 288066 982646 288126 982912
rect 290562 982646 290622 983060
rect 293103 982972 293169 982975
rect 392463 982972 392529 982975
rect 394575 982972 394641 982975
rect 399567 982972 399633 982975
rect 486735 982972 486801 982975
rect 538575 982972 538641 982975
rect 639375 982972 639441 982975
rect 293058 982970 293169 982972
rect 293058 982914 293108 982970
rect 293164 982914 293169 982970
rect 293058 982909 293169 982914
rect 391554 982970 392529 982972
rect 391554 982914 392468 982970
rect 392524 982914 392529 982970
rect 391554 982912 392529 982914
rect 293058 982646 293118 982909
rect 391554 982646 391614 982912
rect 392463 982909 392529 982912
rect 394242 982970 394641 982972
rect 394242 982914 394580 982970
rect 394636 982914 394641 982970
rect 394242 982912 394641 982914
rect 394242 982646 394302 982912
rect 394575 982909 394641 982912
rect 399426 982970 399633 982972
rect 399426 982914 399572 982970
rect 399628 982914 399633 982970
rect 399426 982912 399633 982914
rect 399426 982646 399486 982912
rect 399567 982909 399633 982912
rect 483522 982970 486801 982972
rect 483522 982914 486740 982970
rect 486796 982914 486801 982970
rect 483522 982912 486801 982914
rect 483522 982646 483582 982912
rect 486735 982909 486801 982912
rect 535554 982970 538641 982972
rect 535554 982914 538580 982970
rect 538636 982914 538641 982970
rect 535554 982912 538641 982914
rect 535554 982646 535614 982912
rect 538575 982909 538641 982912
rect 636738 982970 639441 982972
rect 636738 982914 639380 982970
rect 639436 982914 639441 982970
rect 636738 982912 639441 982914
rect 636738 982646 636798 982912
rect 639375 982909 639441 982912
rect 40143 961956 40209 961959
rect 39840 961954 40209 961956
rect 39840 961898 40148 961954
rect 40204 961898 40209 961954
rect 39840 961896 40209 961898
rect 40143 961893 40209 961896
rect 60015 961808 60081 961811
rect 60015 961806 65376 961808
rect 60015 961750 60020 961806
rect 60076 961750 65376 961806
rect 60015 961748 65376 961750
rect 60015 961745 60081 961748
rect 653775 959144 653841 959147
rect 649248 959142 653841 959144
rect 649248 959086 653780 959142
rect 653836 959086 653841 959142
rect 649248 959084 653841 959086
rect 653775 959081 653841 959084
rect 676815 944344 676881 944347
rect 676815 944342 677664 944344
rect 676815 944286 676820 944342
rect 676876 944286 677664 944342
rect 676815 944284 677664 944286
rect 676815 944281 676881 944284
rect 676290 880263 676350 880526
rect 676290 880258 676401 880263
rect 676290 880202 676340 880258
rect 676396 880202 676401 880258
rect 676290 880200 676401 880202
rect 676335 880197 676401 880200
rect 676143 879668 676209 879671
rect 676290 879668 676350 879934
rect 676143 879666 676350 879668
rect 676143 879610 676148 879666
rect 676204 879610 676350 879666
rect 676143 879608 676350 879610
rect 676143 879605 676209 879608
rect 676290 879227 676350 879342
rect 676239 879222 676350 879227
rect 676239 879166 676244 879222
rect 676300 879166 676350 879222
rect 676239 879164 676350 879166
rect 676239 879161 676305 879164
rect 676047 878484 676113 878487
rect 676047 878482 676320 878484
rect 676047 878426 676052 878482
rect 676108 878426 676320 878482
rect 676047 878424 676320 878426
rect 676047 878421 676113 878424
rect 676290 877303 676350 877418
rect 676239 877298 676350 877303
rect 676239 877242 676244 877298
rect 676300 877242 676350 877298
rect 676239 877240 676350 877242
rect 676239 877237 676305 877240
rect 676290 876267 676350 876382
rect 676239 876262 676350 876267
rect 676239 876206 676244 876262
rect 676300 876206 676350 876262
rect 676239 876204 676350 876206
rect 676239 876201 676305 876204
rect 680322 875675 680382 875938
rect 680271 875670 680382 875675
rect 680271 875614 680276 875670
rect 680332 875614 680382 875670
rect 680271 875612 680382 875614
rect 680271 875609 680337 875612
rect 676047 875524 676113 875527
rect 676047 875522 676320 875524
rect 676047 875466 676052 875522
rect 676108 875466 676320 875522
rect 676047 875464 676320 875466
rect 676047 875461 676113 875464
rect 679791 875080 679857 875083
rect 679746 875078 679857 875080
rect 679746 875022 679796 875078
rect 679852 875022 679857 875078
rect 679746 875017 679857 875022
rect 679746 874902 679806 875017
rect 680130 874195 680190 874458
rect 680130 874190 680241 874195
rect 680130 874134 680180 874190
rect 680236 874134 680241 874190
rect 680130 874132 680241 874134
rect 680175 874129 680241 874132
rect 676290 873751 676350 873940
rect 676239 873746 676350 873751
rect 676239 873690 676244 873746
rect 676300 873690 676350 873746
rect 676239 873688 676350 873690
rect 676239 873685 676305 873688
rect 673978 873390 673984 873454
rect 674048 873452 674054 873454
rect 674048 873392 676320 873452
rect 674048 873390 674054 873392
rect 679746 872715 679806 872978
rect 679695 872710 679806 872715
rect 679695 872654 679700 872710
rect 679756 872654 679806 872710
rect 679695 872652 679806 872654
rect 679695 872649 679761 872652
rect 679938 872123 679998 872386
rect 679887 872118 679998 872123
rect 679887 872062 679892 872118
rect 679948 872062 679998 872118
rect 679887 872060 679998 872062
rect 679887 872057 679953 872060
rect 680130 871679 680190 871942
rect 680079 871674 680190 871679
rect 680079 871618 680084 871674
rect 680140 871618 680190 871674
rect 680079 871616 680190 871618
rect 680079 871613 680145 871616
rect 676047 871528 676113 871531
rect 676047 871526 676320 871528
rect 676047 871470 676052 871526
rect 676108 871470 676320 871526
rect 676047 871468 676320 871470
rect 676047 871465 676113 871468
rect 676290 870791 676350 870906
rect 676239 870786 676350 870791
rect 676239 870730 676244 870786
rect 676300 870730 676350 870786
rect 676239 870728 676350 870730
rect 676239 870725 676305 870728
rect 679938 870199 679998 870462
rect 679938 870194 680049 870199
rect 679938 870138 679988 870194
rect 680044 870138 680049 870194
rect 679938 870136 680049 870138
rect 679983 870133 680049 870136
rect 676047 870048 676113 870051
rect 676047 870046 676320 870048
rect 676047 869990 676052 870046
rect 676108 869990 676320 870046
rect 676047 869988 676320 869990
rect 676047 869985 676113 869988
rect 676290 869311 676350 869426
rect 676239 869306 676350 869311
rect 676239 869250 676244 869306
rect 676300 869250 676350 869306
rect 676239 869248 676350 869250
rect 676239 869245 676305 869248
rect 654159 868864 654225 868867
rect 649986 868862 654225 868864
rect 649986 868806 654164 868862
rect 654220 868806 654225 868862
rect 649986 868804 654225 868806
rect 649986 868246 650046 868804
rect 654159 868801 654225 868804
rect 679746 868719 679806 868908
rect 679746 868714 679857 868719
rect 679746 868658 679796 868714
rect 679852 868658 679857 868714
rect 679746 868656 679857 868658
rect 679791 868653 679857 868656
rect 685506 868275 685566 868538
rect 679791 868272 679857 868275
rect 679746 868270 679857 868272
rect 679746 868214 679796 868270
rect 679852 868214 679857 868270
rect 679746 868209 679857 868214
rect 685455 868270 685566 868275
rect 685455 868214 685460 868270
rect 685516 868214 685566 868270
rect 685455 868212 685566 868214
rect 685455 868209 685521 868212
rect 679746 867946 679806 868209
rect 685455 867828 685521 867831
rect 685455 867826 685566 867828
rect 685455 867770 685460 867826
rect 685516 867770 685566 867826
rect 685455 867765 685566 867770
rect 654063 867680 654129 867683
rect 649986 867678 654129 867680
rect 649986 867622 654068 867678
rect 654124 867622 654129 867678
rect 649986 867620 654129 867622
rect 649986 867064 650046 867620
rect 654063 867617 654129 867620
rect 685506 867354 685566 867765
rect 654255 866496 654321 866499
rect 649986 866494 654321 866496
rect 649986 866438 654260 866494
rect 654316 866438 654321 866494
rect 649986 866436 654321 866438
rect 649986 865882 650046 866436
rect 654255 866433 654321 866436
rect 649986 864128 650046 864700
rect 654255 864128 654321 864131
rect 649986 864126 654321 864128
rect 649986 864070 654260 864126
rect 654316 864070 654321 864126
rect 649986 864068 654321 864070
rect 654255 864065 654321 864068
rect 649986 862944 650046 863518
rect 654831 862944 654897 862947
rect 649986 862942 654897 862944
rect 649986 862886 654836 862942
rect 654892 862886 654897 862942
rect 649986 862884 654897 862886
rect 654831 862881 654897 862884
rect 649986 861908 650046 862336
rect 656367 861908 656433 861911
rect 649986 861906 656433 861908
rect 649986 861850 656372 861906
rect 656428 861850 656433 861906
rect 649986 861848 656433 861850
rect 656367 861845 656433 861848
rect 673978 852522 673984 852586
rect 674048 852584 674054 852586
rect 675183 852584 675249 852587
rect 674048 852582 675249 852584
rect 674048 852526 675188 852582
rect 675244 852526 675249 852582
rect 674048 852524 675249 852526
rect 674048 852522 674054 852524
rect 675183 852521 675249 852524
rect 41775 817952 41841 817955
rect 41568 817950 41841 817952
rect 41568 817894 41780 817950
rect 41836 817894 41841 817950
rect 41568 817892 41841 817894
rect 41775 817889 41841 817892
rect 41775 817360 41841 817363
rect 41568 817358 41841 817360
rect 41568 817302 41780 817358
rect 41836 817302 41841 817358
rect 41568 817300 41841 817302
rect 41775 817297 41841 817300
rect 41538 816623 41598 816738
rect 41538 816618 41649 816623
rect 41538 816562 41588 816618
rect 41644 816562 41649 816618
rect 41538 816560 41649 816562
rect 41583 816557 41649 816560
rect 41775 815880 41841 815883
rect 41568 815878 41841 815880
rect 41568 815822 41780 815878
rect 41836 815822 41841 815878
rect 41568 815820 41841 815822
rect 41775 815817 41841 815820
rect 40386 815142 40446 815258
rect 40378 815078 40384 815142
rect 40448 815078 40454 815142
rect 41775 814918 41841 814921
rect 41568 814916 41841 814918
rect 41568 814860 41780 814916
rect 41836 814860 41841 814916
rect 41568 814858 41841 814860
rect 41775 814855 41841 814858
rect 40578 814106 40638 814370
rect 40570 814042 40576 814106
rect 40640 814042 40646 814106
rect 41538 813663 41598 813778
rect 41538 813658 41649 813663
rect 41538 813602 41588 813658
rect 41644 813602 41649 813658
rect 41538 813600 41649 813602
rect 41583 813597 41649 813600
rect 40770 813070 40830 813334
rect 40762 813006 40768 813070
rect 40832 813006 40838 813070
rect 42063 812920 42129 812923
rect 41568 812918 42129 812920
rect 41568 812862 42068 812918
rect 42124 812862 42129 812918
rect 41568 812860 42129 812862
rect 42063 812857 42129 812860
rect 34479 812476 34545 812479
rect 34434 812474 34545 812476
rect 34434 812418 34484 812474
rect 34540 812418 34545 812474
rect 34434 812413 34545 812418
rect 34434 812298 34494 812413
rect 37314 811739 37374 811854
rect 37314 811734 37425 811739
rect 37314 811678 37364 811734
rect 37420 811678 37425 811734
rect 37314 811676 37425 811678
rect 37359 811673 37425 811676
rect 41967 811366 42033 811369
rect 41568 811364 42033 811366
rect 41568 811308 41972 811364
rect 42028 811308 42033 811364
rect 41568 811306 42033 811308
rect 41967 811303 42033 811306
rect 41775 810848 41841 810851
rect 41568 810846 41841 810848
rect 41568 810790 41780 810846
rect 41836 810790 41841 810846
rect 41568 810788 41841 810790
rect 41775 810785 41841 810788
rect 34434 810259 34494 810374
rect 34383 810254 34494 810259
rect 34383 810198 34388 810254
rect 34444 810198 34494 810254
rect 34383 810196 34494 810198
rect 34383 810193 34449 810196
rect 40194 809667 40254 809856
rect 40143 809662 40254 809667
rect 40143 809606 40148 809662
rect 40204 809606 40254 809662
rect 40143 809604 40254 809606
rect 40143 809601 40209 809604
rect 40239 809516 40305 809519
rect 40194 809514 40305 809516
rect 40194 809458 40244 809514
rect 40300 809458 40305 809514
rect 40194 809453 40305 809458
rect 40194 809338 40254 809453
rect 41871 808924 41937 808927
rect 41568 808922 41937 808924
rect 41568 808866 41876 808922
rect 41932 808866 41937 808922
rect 41568 808864 41937 808866
rect 41871 808861 41937 808864
rect 41538 808187 41598 808302
rect 41538 808182 41649 808187
rect 41538 808126 41588 808182
rect 41644 808126 41649 808182
rect 41538 808124 41649 808126
rect 41583 808121 41649 808124
rect 41871 807888 41937 807891
rect 41568 807886 41937 807888
rect 41568 807830 41876 807886
rect 41932 807830 41937 807886
rect 41568 807828 41937 807830
rect 41871 807825 41937 807828
rect 41346 807151 41406 807414
rect 41346 807146 41457 807151
rect 41346 807090 41396 807146
rect 41452 807090 41457 807146
rect 41346 807088 41457 807090
rect 41391 807085 41457 807088
rect 41538 806707 41598 806822
rect 41538 806702 41649 806707
rect 41538 806646 41588 806702
rect 41644 806646 41649 806702
rect 41538 806644 41649 806646
rect 41583 806641 41649 806644
rect 41538 806115 41598 806304
rect 41538 806110 41649 806115
rect 41538 806054 41588 806110
rect 41644 806054 41649 806110
rect 41538 806052 41649 806054
rect 41583 806049 41649 806052
rect 28866 805671 28926 805934
rect 28815 805666 28926 805671
rect 28815 805610 28820 805666
rect 28876 805610 28926 805666
rect 28815 805608 28926 805610
rect 28815 805605 28881 805608
rect 41538 805227 41598 805342
rect 28815 805224 28881 805227
rect 28815 805222 28926 805224
rect 28815 805166 28820 805222
rect 28876 805166 28926 805222
rect 28815 805161 28926 805166
rect 41538 805222 41649 805227
rect 41538 805166 41588 805222
rect 41644 805166 41649 805222
rect 41538 805164 41649 805166
rect 41583 805161 41649 805164
rect 28866 804824 28926 805161
rect 34479 805076 34545 805079
rect 41530 805076 41536 805078
rect 34479 805074 41536 805076
rect 34479 805018 34484 805074
rect 34540 805018 41536 805074
rect 34479 805016 41536 805018
rect 34479 805013 34545 805016
rect 41530 805014 41536 805016
rect 41600 805014 41606 805078
rect 41871 801082 41937 801083
rect 41871 801078 41920 801082
rect 41984 801080 41990 801082
rect 41871 801022 41876 801078
rect 41871 801018 41920 801022
rect 41984 801020 42028 801080
rect 41984 801018 41990 801020
rect 41871 801017 41937 801018
rect 42490 800722 42496 800786
rect 42560 800784 42566 800786
rect 42639 800784 42705 800787
rect 42560 800782 42705 800784
rect 42560 800726 42644 800782
rect 42700 800726 42705 800782
rect 42560 800724 42705 800726
rect 42560 800722 42566 800724
rect 42639 800721 42705 800724
rect 42298 800574 42304 800638
rect 42368 800636 42374 800638
rect 43407 800636 43473 800639
rect 42368 800634 43473 800636
rect 42368 800578 43412 800634
rect 43468 800578 43473 800634
rect 42368 800576 43473 800578
rect 42368 800574 42374 800576
rect 43407 800573 43473 800576
rect 42490 800426 42496 800490
rect 42560 800488 42566 800490
rect 43119 800488 43185 800491
rect 42560 800486 43185 800488
rect 42560 800430 43124 800486
rect 43180 800430 43185 800486
rect 42560 800428 43185 800430
rect 42560 800426 42566 800428
rect 43119 800425 43185 800428
rect 41914 798798 41920 798862
rect 41984 798860 41990 798862
rect 42639 798860 42705 798863
rect 41984 798858 42705 798860
rect 41984 798802 42644 798858
rect 42700 798802 42705 798858
rect 41984 798800 42705 798802
rect 41984 798798 41990 798800
rect 42639 798797 42705 798800
rect 40762 793914 40768 793978
rect 40832 793976 40838 793978
rect 43023 793976 43089 793979
rect 40832 793974 43089 793976
rect 40832 793918 43028 793974
rect 43084 793918 43089 793974
rect 40832 793916 43089 793918
rect 40832 793914 40838 793916
rect 43023 793913 43089 793916
rect 42159 790276 42225 790279
rect 42298 790276 42304 790278
rect 42159 790274 42304 790276
rect 42159 790218 42164 790274
rect 42220 790218 42304 790274
rect 42159 790216 42304 790218
rect 42159 790213 42225 790216
rect 42298 790214 42304 790216
rect 42368 790214 42374 790278
rect 57999 789832 58065 789835
rect 64578 789832 64638 790304
rect 57999 789830 64638 789832
rect 57999 789774 58004 789830
rect 58060 789774 64638 789830
rect 57999 789772 64638 789774
rect 57999 789769 58065 789772
rect 57615 789684 57681 789687
rect 57615 789682 64638 789684
rect 57615 789626 57620 789682
rect 57676 789626 64638 789682
rect 57615 789624 64638 789626
rect 57615 789621 57681 789624
rect 64578 789122 64638 789624
rect 58191 788500 58257 788503
rect 58191 788498 64638 788500
rect 58191 788442 58196 788498
rect 58252 788442 64638 788498
rect 58191 788440 64638 788442
rect 58191 788437 58257 788440
rect 64578 787940 64638 788440
rect 58383 787316 58449 787319
rect 58383 787314 64638 787316
rect 58383 787258 58388 787314
rect 58444 787258 64638 787314
rect 58383 787256 64638 787258
rect 58383 787253 58449 787256
rect 64578 786758 64638 787256
rect 41530 786366 41536 786430
rect 41600 786428 41606 786430
rect 41775 786428 41841 786431
rect 41600 786426 41841 786428
rect 41600 786370 41780 786426
rect 41836 786370 41841 786426
rect 41600 786368 41841 786370
rect 41600 786366 41606 786368
rect 41775 786365 41841 786368
rect 59631 785392 59697 785395
rect 64578 785392 64638 785576
rect 59631 785390 64638 785392
rect 59631 785334 59636 785390
rect 59692 785334 64638 785390
rect 59631 785332 64638 785334
rect 59631 785329 59697 785332
rect 58671 784948 58737 784951
rect 58671 784946 64638 784948
rect 58671 784890 58676 784946
rect 58732 784890 64638 784946
rect 58671 784888 64638 784890
rect 58671 784885 58737 784888
rect 64578 784394 64638 784888
rect 649986 778288 650046 778824
rect 655215 778288 655281 778291
rect 649986 778286 655281 778288
rect 649986 778230 655220 778286
rect 655276 778230 655281 778286
rect 649986 778228 655281 778230
rect 655215 778225 655281 778228
rect 655599 777696 655665 777699
rect 649986 777694 655665 777696
rect 649986 777638 655604 777694
rect 655660 777638 655665 777694
rect 649986 777636 655665 777638
rect 655599 777633 655665 777636
rect 649986 775920 650046 776460
rect 655407 775920 655473 775923
rect 649986 775918 655473 775920
rect 649986 775862 655412 775918
rect 655468 775862 655473 775918
rect 649986 775860 655473 775862
rect 655407 775857 655473 775860
rect 649986 774884 650046 775278
rect 654159 774884 654225 774887
rect 649986 774882 654225 774884
rect 649986 774826 654164 774882
rect 654220 774826 654225 774882
rect 649986 774824 654225 774826
rect 654159 774821 654225 774824
rect 41775 774736 41841 774739
rect 41568 774734 41841 774736
rect 41568 774678 41780 774734
rect 41836 774678 41841 774734
rect 41568 774676 41841 774678
rect 41775 774673 41841 774676
rect 674746 774526 674752 774590
rect 674816 774588 674822 774590
rect 675471 774588 675537 774591
rect 674816 774586 675537 774588
rect 674816 774530 675476 774586
rect 675532 774530 675537 774586
rect 674816 774528 675537 774530
rect 674816 774526 674822 774528
rect 675471 774525 675537 774528
rect 41538 773999 41598 774114
rect 41538 773994 41649 773999
rect 41538 773938 41588 773994
rect 41644 773938 41649 773994
rect 41538 773936 41649 773938
rect 41583 773933 41649 773936
rect 41775 773552 41841 773555
rect 41568 773550 41841 773552
rect 41568 773494 41780 773550
rect 41836 773494 41841 773550
rect 41568 773492 41841 773494
rect 649986 773552 650046 774096
rect 674554 773638 674560 773702
rect 674624 773700 674630 773702
rect 675375 773700 675441 773703
rect 674624 773698 675441 773700
rect 674624 773642 675380 773698
rect 675436 773642 675441 773698
rect 674624 773640 675441 773642
rect 674624 773638 674630 773640
rect 675375 773637 675441 773640
rect 656175 773552 656241 773555
rect 649986 773550 656241 773552
rect 649986 773494 656180 773550
rect 656236 773494 656241 773550
rect 649986 773492 656241 773494
rect 41775 773489 41841 773492
rect 656175 773489 656241 773492
rect 41583 773404 41649 773407
rect 41538 773402 41649 773404
rect 41538 773346 41588 773402
rect 41644 773346 41649 773402
rect 41538 773341 41649 773346
rect 41538 773226 41598 773341
rect 675759 773108 675825 773111
rect 676090 773108 676096 773110
rect 675759 773106 676096 773108
rect 675759 773050 675764 773106
rect 675820 773050 676096 773106
rect 675759 773048 676096 773050
rect 675759 773045 675825 773048
rect 676090 773046 676096 773048
rect 676160 773046 676166 773110
rect 41775 772664 41841 772667
rect 41568 772662 41841 772664
rect 41568 772606 41780 772662
rect 41836 772606 41841 772662
rect 41568 772604 41841 772606
rect 41775 772601 41841 772604
rect 40570 772306 40576 772370
rect 40640 772368 40646 772370
rect 41583 772368 41649 772371
rect 40640 772366 41649 772368
rect 40640 772310 41588 772366
rect 41644 772310 41649 772366
rect 40640 772308 41649 772310
rect 649986 772368 650046 772914
rect 654831 772368 654897 772371
rect 649986 772366 654897 772368
rect 649986 772310 654836 772366
rect 654892 772310 654897 772366
rect 649986 772308 654897 772310
rect 40640 772306 40646 772308
rect 41583 772305 41649 772308
rect 654831 772305 654897 772308
rect 40194 771926 40254 772042
rect 40186 771862 40192 771926
rect 40256 771862 40262 771926
rect 40378 771862 40384 771926
rect 40448 771924 40454 771926
rect 43119 771924 43185 771927
rect 40448 771922 43185 771924
rect 40448 771866 43124 771922
rect 43180 771866 43185 771922
rect 40448 771864 43185 771866
rect 40448 771862 40454 771864
rect 41538 771672 41598 771864
rect 43119 771861 43185 771864
rect 40578 770890 40638 771154
rect 40570 770826 40576 770890
rect 40640 770826 40646 770890
rect 41583 770888 41649 770891
rect 41538 770886 41649 770888
rect 41538 770830 41588 770886
rect 41644 770830 41649 770886
rect 41538 770825 41649 770830
rect 41538 770562 41598 770825
rect 675759 770740 675825 770743
rect 675898 770740 675904 770742
rect 675759 770738 675904 770740
rect 675759 770682 675764 770738
rect 675820 770682 675904 770738
rect 675759 770680 675904 770682
rect 675759 770677 675825 770680
rect 675898 770678 675904 770680
rect 675968 770678 675974 770742
rect 40770 769854 40830 770192
rect 675471 770002 675537 770003
rect 675471 769998 675520 770002
rect 675584 770000 675590 770002
rect 675471 769942 675476 769998
rect 675471 769938 675520 769942
rect 675584 769940 675628 770000
rect 675584 769938 675590 769940
rect 675471 769937 675537 769938
rect 40762 769790 40768 769854
rect 40832 769790 40838 769854
rect 41775 769704 41841 769707
rect 41568 769702 41841 769704
rect 41568 769646 41780 769702
rect 41836 769646 41841 769702
rect 41568 769644 41841 769646
rect 41775 769641 41841 769644
rect 674362 769346 674368 769410
rect 674432 769408 674438 769410
rect 675471 769408 675537 769411
rect 674432 769406 675537 769408
rect 674432 769350 675476 769406
rect 675532 769350 675537 769406
rect 674432 769348 675537 769350
rect 674432 769346 674438 769348
rect 675471 769345 675537 769348
rect 41346 768966 41406 769082
rect 41338 768902 41344 768966
rect 41408 768902 41414 768966
rect 37314 768523 37374 768638
rect 37314 768518 37425 768523
rect 37314 768462 37364 768518
rect 37420 768462 37425 768518
rect 37314 768460 37425 768462
rect 37359 768457 37425 768460
rect 42255 768224 42321 768227
rect 41568 768222 42321 768224
rect 41568 768166 42260 768222
rect 42316 768166 42321 768222
rect 41568 768164 42321 768166
rect 42255 768161 42321 768164
rect 41871 767632 41937 767635
rect 41568 767630 41937 767632
rect 41568 767574 41876 767630
rect 41932 767574 41937 767630
rect 41568 767572 41937 767574
rect 41871 767569 41937 767572
rect 42063 767188 42129 767191
rect 41568 767186 42129 767188
rect 41568 767130 42068 767186
rect 42124 767130 42129 767186
rect 41568 767128 42129 767130
rect 42063 767125 42129 767128
rect 40194 766451 40254 766640
rect 40194 766446 40305 766451
rect 40194 766390 40244 766446
rect 40300 766390 40305 766446
rect 40194 766388 40305 766390
rect 40239 766385 40305 766388
rect 40143 766300 40209 766303
rect 40143 766298 40254 766300
rect 40143 766242 40148 766298
rect 40204 766242 40254 766298
rect 40143 766237 40254 766242
rect 40194 766122 40254 766237
rect 41538 765563 41598 765678
rect 41538 765558 41649 765563
rect 41538 765502 41588 765558
rect 41644 765502 41649 765558
rect 41538 765500 41649 765502
rect 41583 765497 41649 765500
rect 41775 765190 41841 765193
rect 41568 765188 41841 765190
rect 41568 765132 41780 765188
rect 41836 765132 41841 765188
rect 41568 765130 41841 765132
rect 41775 765127 41841 765130
rect 42159 764672 42225 764675
rect 41568 764670 42225 764672
rect 41568 764614 42164 764670
rect 42220 764614 42225 764670
rect 41568 764612 42225 764614
rect 42159 764609 42225 764612
rect 41967 764228 42033 764231
rect 41568 764226 42033 764228
rect 41568 764170 41972 764226
rect 42028 764170 42033 764226
rect 41568 764168 42033 764170
rect 41967 764165 42033 764168
rect 41538 763491 41598 763606
rect 41538 763486 41649 763491
rect 41538 763430 41588 763486
rect 41644 763430 41649 763486
rect 41538 763428 41649 763430
rect 41583 763425 41649 763428
rect 41538 762896 41598 763162
rect 41538 762836 41790 762896
rect 28866 762455 28926 762718
rect 28815 762450 28926 762455
rect 41730 762452 41790 762836
rect 28815 762394 28820 762450
rect 28876 762394 28926 762450
rect 28815 762392 28926 762394
rect 41538 762392 41790 762452
rect 28815 762389 28881 762392
rect 41538 762156 41598 762392
rect 41775 762156 41841 762159
rect 41538 762154 41841 762156
rect 41538 762126 41780 762154
rect 41568 762098 41780 762126
rect 41836 762098 41841 762154
rect 41568 762096 41841 762098
rect 41775 762093 41841 762096
rect 28815 762008 28881 762011
rect 28815 762006 28926 762008
rect 28815 761950 28820 762006
rect 28876 761950 28926 762006
rect 28815 761945 28926 761950
rect 28866 761608 28926 761945
rect 41007 760232 41073 760235
rect 41146 760232 41152 760234
rect 41007 760230 41152 760232
rect 41007 760174 41012 760230
rect 41068 760174 41152 760230
rect 41007 760172 41152 760174
rect 41007 760169 41073 760172
rect 41146 760170 41152 760172
rect 41216 760170 41222 760234
rect 41775 758012 41841 758015
rect 42106 758012 42112 758014
rect 41775 758010 42112 758012
rect 41775 757954 41780 758010
rect 41836 757954 42112 758010
rect 41775 757952 42112 757954
rect 41775 757949 41841 757952
rect 42106 757950 42112 757952
rect 42176 757950 42182 758014
rect 42063 757864 42129 757867
rect 42298 757864 42304 757866
rect 42063 757862 42304 757864
rect 42063 757806 42068 757862
rect 42124 757806 42304 757862
rect 42063 757804 42304 757806
rect 42063 757801 42129 757804
rect 42298 757802 42304 757804
rect 42368 757802 42374 757866
rect 42298 752474 42304 752538
rect 42368 752536 42374 752538
rect 42831 752536 42897 752539
rect 42368 752534 42897 752536
rect 42368 752478 42836 752534
rect 42892 752478 42897 752534
rect 42368 752476 42897 752478
rect 42368 752474 42374 752476
rect 42831 752473 42897 752476
rect 42106 751142 42112 751206
rect 42176 751204 42182 751206
rect 42927 751204 42993 751207
rect 42176 751202 42993 751204
rect 42176 751146 42932 751202
rect 42988 751146 42993 751202
rect 42176 751144 42993 751146
rect 42176 751142 42182 751144
rect 42927 751141 42993 751144
rect 40762 748774 40768 748838
rect 40832 748836 40838 748838
rect 43023 748836 43089 748839
rect 40832 748834 43089 748836
rect 40832 748778 43028 748834
rect 43084 748778 43089 748834
rect 40832 748776 43089 748778
rect 40832 748774 40838 748776
rect 43023 748773 43089 748776
rect 57903 747652 57969 747655
rect 57903 747650 64638 747652
rect 57903 747594 57908 747650
rect 57964 747594 64638 747650
rect 57903 747592 64638 747594
rect 57903 747589 57969 747592
rect 41338 747294 41344 747358
rect 41408 747356 41414 747358
rect 42831 747356 42897 747359
rect 41408 747354 42897 747356
rect 41408 747298 42836 747354
rect 42892 747298 42897 747354
rect 41408 747296 42897 747298
rect 41408 747294 41414 747296
rect 42831 747293 42897 747296
rect 64578 747082 64638 747592
rect 41146 746998 41152 747062
rect 41216 747060 41222 747062
rect 41775 747060 41841 747063
rect 41216 747058 41841 747060
rect 41216 747002 41780 747058
rect 41836 747002 41841 747058
rect 41216 747000 41841 747002
rect 41216 746998 41222 747000
rect 41775 746997 41841 747000
rect 54735 746024 54801 746027
rect 54690 746022 54801 746024
rect 54690 745966 54740 746022
rect 54796 745966 54801 746022
rect 54690 745961 54801 745966
rect 54690 745879 54750 745961
rect 54639 745874 54750 745879
rect 54639 745818 54644 745874
rect 54700 745818 54750 745874
rect 54639 745816 54750 745818
rect 54639 745813 54705 745816
rect 59631 745432 59697 745435
rect 64578 745432 64638 745900
rect 59631 745430 64638 745432
rect 59631 745374 59636 745430
rect 59692 745374 64638 745430
rect 59631 745372 64638 745374
rect 59631 745369 59697 745372
rect 57615 745284 57681 745287
rect 57615 745282 64638 745284
rect 57615 745226 57620 745282
rect 57676 745226 64638 745282
rect 57615 745224 64638 745226
rect 57615 745221 57681 745224
rect 64578 744718 64638 745224
rect 59247 744100 59313 744103
rect 59247 744098 64638 744100
rect 59247 744042 59252 744098
rect 59308 744042 64638 744098
rect 59247 744040 64638 744042
rect 59247 744037 59313 744040
rect 64578 743536 64638 744040
rect 59631 742916 59697 742919
rect 59631 742914 64638 742916
rect 59631 742858 59636 742914
rect 59692 742858 64638 742914
rect 59631 742856 64638 742858
rect 59631 742853 59697 742856
rect 64578 742354 64638 742856
rect 59727 741732 59793 741735
rect 59727 741730 64638 741732
rect 59727 741674 59732 741730
rect 59788 741674 64638 741730
rect 59727 741672 64638 741674
rect 59727 741669 59793 741672
rect 64578 741172 64638 741672
rect 655119 734480 655185 734483
rect 649986 734478 655185 734480
rect 649986 734422 655124 734478
rect 655180 734422 655185 734478
rect 649986 734420 655185 734422
rect 649986 734402 650046 734420
rect 655119 734417 655185 734420
rect 649986 732704 650046 733220
rect 655503 732704 655569 732707
rect 649986 732702 655569 732704
rect 649986 732646 655508 732702
rect 655564 732646 655569 732702
rect 649986 732644 655569 732646
rect 655503 732641 655569 732644
rect 649986 731668 650046 732038
rect 655311 731668 655377 731671
rect 649986 731666 655377 731668
rect 649986 731610 655316 731666
rect 655372 731610 655377 731666
rect 649986 731608 655377 731610
rect 655311 731605 655377 731608
rect 674511 731668 674577 731671
rect 677050 731668 677056 731670
rect 674511 731666 677056 731668
rect 674511 731610 674516 731666
rect 674572 731610 677056 731666
rect 674511 731608 677056 731610
rect 674511 731605 674577 731608
rect 677050 731606 677056 731608
rect 677120 731606 677126 731670
rect 41775 731520 41841 731523
rect 41568 731518 41841 731520
rect 41568 731462 41780 731518
rect 41836 731462 41841 731518
rect 41568 731460 41841 731462
rect 41775 731457 41841 731460
rect 41538 730783 41598 730898
rect 41538 730778 41649 730783
rect 41538 730722 41588 730778
rect 41644 730722 41649 730778
rect 41538 730720 41649 730722
rect 41583 730717 41649 730720
rect 41775 730410 41841 730413
rect 41568 730408 41841 730410
rect 41568 730352 41780 730408
rect 41836 730352 41841 730408
rect 41568 730350 41841 730352
rect 41775 730347 41841 730350
rect 649986 730336 650046 730856
rect 654159 730336 654225 730339
rect 649986 730334 654225 730336
rect 649986 730278 654164 730334
rect 654220 730278 654225 730334
rect 649986 730276 654225 730278
rect 654159 730273 654225 730276
rect 41583 730188 41649 730191
rect 41538 730186 41649 730188
rect 41538 730130 41588 730186
rect 41644 730130 41649 730186
rect 41538 730125 41649 730130
rect 41538 730010 41598 730125
rect 674938 729830 674944 729894
rect 675008 729892 675014 729894
rect 675471 729892 675537 729895
rect 675008 729890 675537 729892
rect 675008 729834 675476 729890
rect 675532 729834 675537 729890
rect 675008 729832 675537 729834
rect 675008 729830 675014 729832
rect 675471 729829 675537 729832
rect 41538 729303 41598 729418
rect 40570 729238 40576 729302
rect 40640 729300 40646 729302
rect 41199 729300 41265 729303
rect 40640 729298 41265 729300
rect 40640 729242 41204 729298
rect 41260 729242 41265 729298
rect 40640 729240 41265 729242
rect 41538 729298 41649 729303
rect 41538 729242 41588 729298
rect 41644 729242 41649 729298
rect 41538 729240 41649 729242
rect 40640 729238 40646 729240
rect 41199 729237 41265 729240
rect 41583 729237 41649 729240
rect 649986 729152 650046 729674
rect 675759 729448 675825 729451
rect 676282 729448 676288 729450
rect 675759 729446 676288 729448
rect 675759 729390 675764 729446
rect 675820 729390 676288 729446
rect 675759 729388 676288 729390
rect 675759 729385 675825 729388
rect 676282 729386 676288 729388
rect 676352 729386 676358 729450
rect 654255 729152 654321 729155
rect 649986 729150 654321 729152
rect 649986 729094 654260 729150
rect 654316 729094 654321 729150
rect 649986 729092 654321 729094
rect 654255 729089 654321 729092
rect 41538 728711 41598 728826
rect 40431 728710 40497 728711
rect 40378 728646 40384 728710
rect 40448 728708 40497 728710
rect 40448 728706 40576 728708
rect 40492 728650 40576 728706
rect 40448 728648 40576 728650
rect 41538 728706 41649 728711
rect 41538 728650 41588 728706
rect 41644 728650 41649 728706
rect 41538 728648 41649 728650
rect 40448 728646 40497 728648
rect 40386 728645 40497 728646
rect 41583 728645 41649 728648
rect 675663 728710 675729 728711
rect 675663 728706 675712 728710
rect 675776 728708 675782 728710
rect 675663 728650 675668 728706
rect 675663 728646 675712 728650
rect 675776 728648 675820 728708
rect 675776 728646 675782 728648
rect 675663 728645 675729 728646
rect 40386 728530 40446 728645
rect 41775 727968 41841 727971
rect 41568 727966 41841 727968
rect 41568 727910 41780 727966
rect 41836 727910 41841 727966
rect 41568 727908 41841 727910
rect 649986 727968 650046 728492
rect 654159 727968 654225 727971
rect 649986 727966 654225 727968
rect 649986 727910 654164 727966
rect 654220 727910 654225 727966
rect 649986 727908 654225 727910
rect 41775 727905 41841 727908
rect 654159 727905 654225 727908
rect 40570 727610 40576 727674
rect 40640 727610 40646 727674
rect 40578 727346 40638 727610
rect 34434 726787 34494 726976
rect 34434 726782 34545 726787
rect 675375 726786 675441 726787
rect 675322 726784 675328 726786
rect 34434 726726 34484 726782
rect 34540 726726 34545 726782
rect 34434 726724 34545 726726
rect 675284 726724 675328 726784
rect 675392 726782 675441 726786
rect 675436 726726 675441 726782
rect 34479 726721 34545 726724
rect 675322 726722 675328 726724
rect 675392 726722 675441 726726
rect 675375 726721 675441 726722
rect 41775 726488 41841 726491
rect 41568 726486 41841 726488
rect 41568 726430 41780 726486
rect 41836 726430 41841 726486
rect 41568 726428 41841 726430
rect 41775 726425 41841 726428
rect 675759 726192 675825 726195
rect 676474 726192 676480 726194
rect 675759 726190 676480 726192
rect 675759 726134 675764 726190
rect 675820 726134 676480 726190
rect 675759 726132 676480 726134
rect 675759 726129 675825 726132
rect 676474 726130 676480 726132
rect 676544 726130 676550 726194
rect 41154 725750 41214 725866
rect 673978 725834 673984 725898
rect 674048 725896 674054 725898
rect 675375 725896 675441 725899
rect 674048 725894 675441 725896
rect 674048 725838 675380 725894
rect 675436 725838 675441 725894
rect 674048 725836 675441 725838
rect 674048 725834 674054 725836
rect 675375 725833 675441 725836
rect 41146 725686 41152 725750
rect 41216 725686 41222 725750
rect 37314 725307 37374 725496
rect 37314 725302 37425 725307
rect 37314 725246 37364 725302
rect 37420 725246 37425 725302
rect 37314 725244 37425 725246
rect 37359 725241 37425 725244
rect 41967 725008 42033 725011
rect 41568 725006 42033 725008
rect 41568 724950 41972 725006
rect 42028 724950 42033 725006
rect 41568 724948 42033 724950
rect 41967 724945 42033 724948
rect 41775 724416 41841 724419
rect 41568 724414 41841 724416
rect 41568 724358 41780 724414
rect 41836 724358 41841 724414
rect 41568 724356 41841 724358
rect 41775 724353 41841 724356
rect 40962 723826 41022 723942
rect 40954 723762 40960 723826
rect 41024 723762 41030 723826
rect 40194 723235 40254 723498
rect 40143 723230 40254 723235
rect 40143 723174 40148 723230
rect 40204 723174 40254 723230
rect 40143 723172 40254 723174
rect 40143 723169 40209 723172
rect 40239 723084 40305 723087
rect 40194 723082 40305 723084
rect 40194 723026 40244 723082
rect 40300 723026 40305 723082
rect 40194 723021 40305 723026
rect 40194 722906 40254 723021
rect 41538 722347 41598 722462
rect 41538 722342 41649 722347
rect 41538 722286 41588 722342
rect 41644 722286 41649 722342
rect 41538 722284 41649 722286
rect 41583 722281 41649 722284
rect 41871 721974 41937 721977
rect 41568 721972 41937 721974
rect 41568 721916 41876 721972
rect 41932 721916 41937 721972
rect 41568 721914 41937 721916
rect 41871 721911 41937 721914
rect 675759 721900 675825 721903
rect 676858 721900 676864 721902
rect 675759 721898 676864 721900
rect 675759 721842 675764 721898
rect 675820 721842 676864 721898
rect 675759 721840 676864 721842
rect 675759 721837 675825 721840
rect 676858 721838 676864 721840
rect 676928 721838 676934 721902
rect 42255 721456 42321 721459
rect 41568 721454 42321 721456
rect 41568 721398 42260 721454
rect 42316 721398 42321 721454
rect 41568 721396 42321 721398
rect 42255 721393 42321 721396
rect 41538 720867 41598 720982
rect 41538 720862 41649 720867
rect 41538 720806 41588 720862
rect 41644 720806 41649 720862
rect 41538 720804 41649 720806
rect 41583 720801 41649 720804
rect 41538 720275 41598 720464
rect 41538 720270 41649 720275
rect 41538 720214 41588 720270
rect 41644 720214 41649 720270
rect 41538 720212 41649 720214
rect 41583 720209 41649 720212
rect 41538 719680 41598 719946
rect 41538 719620 41790 719680
rect 28866 719239 28926 719502
rect 28815 719234 28926 719239
rect 41730 719236 41790 719620
rect 28815 719178 28820 719234
rect 28876 719178 28926 719234
rect 28815 719176 28926 719178
rect 41538 719176 41790 719236
rect 28815 719173 28881 719176
rect 41538 718795 41598 719176
rect 28815 718792 28881 718795
rect 28815 718790 28926 718792
rect 28815 718734 28820 718790
rect 28876 718734 28926 718790
rect 28815 718729 28926 718734
rect 41538 718790 41649 718795
rect 41538 718734 41588 718790
rect 41644 718734 41649 718790
rect 41538 718732 41649 718734
rect 41583 718729 41649 718732
rect 28866 718466 28926 718729
rect 37359 718644 37425 718647
rect 42298 718644 42304 718646
rect 37359 718642 42304 718644
rect 37359 718586 37364 718642
rect 37420 718586 42304 718642
rect 37359 718584 42304 718586
rect 37359 718581 37425 718584
rect 42298 718582 42304 718584
rect 42368 718582 42374 718646
rect 34479 717756 34545 717759
rect 40378 717756 40384 717758
rect 34479 717754 40384 717756
rect 34479 717698 34484 717754
rect 34540 717698 40384 717754
rect 34479 717696 40384 717698
rect 34479 717693 34545 717696
rect 40378 717694 40384 717696
rect 40448 717694 40454 717758
rect 40239 717016 40305 717019
rect 40762 717016 40768 717018
rect 40239 717014 40768 717016
rect 40239 716958 40244 717014
rect 40300 716958 40768 717014
rect 40239 716956 40768 716958
rect 40239 716953 40305 716956
rect 40762 716954 40768 716956
rect 40832 716954 40838 717018
rect 40143 716868 40209 716871
rect 40570 716868 40576 716870
rect 40143 716866 40576 716868
rect 40143 716810 40148 716866
rect 40204 716810 40576 716866
rect 40143 716808 40576 716810
rect 40143 716805 40209 716808
rect 40570 716806 40576 716808
rect 40640 716806 40646 716870
rect 40570 708814 40576 708878
rect 40640 708876 40646 708878
rect 43119 708876 43185 708879
rect 40640 708874 43185 708876
rect 40640 708818 43124 708874
rect 43180 708818 43185 708874
rect 40640 708816 43185 708818
rect 40640 708814 40646 708816
rect 43119 708813 43185 708816
rect 42298 708666 42304 708730
rect 42368 708728 42374 708730
rect 43023 708728 43089 708731
rect 42368 708726 43089 708728
rect 42368 708670 43028 708726
rect 43084 708670 43089 708726
rect 42368 708668 43089 708670
rect 42368 708666 42374 708668
rect 43023 708665 43089 708668
rect 40762 708518 40768 708582
rect 40832 708580 40838 708582
rect 42831 708580 42897 708583
rect 40832 708578 42897 708580
rect 40832 708522 42836 708578
rect 42892 708522 42897 708578
rect 40832 708520 42897 708522
rect 40832 708518 40838 708520
rect 42831 708517 42897 708520
rect 40954 705854 40960 705918
rect 41024 705916 41030 705918
rect 42927 705916 42993 705919
rect 41024 705914 42993 705916
rect 41024 705858 42932 705914
rect 42988 705858 42993 705914
rect 41024 705856 42993 705858
rect 41024 705854 41030 705856
rect 42927 705853 42993 705856
rect 41146 705410 41152 705474
rect 41216 705472 41222 705474
rect 42735 705472 42801 705475
rect 41216 705470 42801 705472
rect 41216 705414 42740 705470
rect 42796 705414 42801 705470
rect 41216 705412 42801 705414
rect 41216 705410 41222 705412
rect 42735 705409 42801 705412
rect 58383 704436 58449 704439
rect 58383 704434 64638 704436
rect 58383 704378 58388 704434
rect 58444 704378 64638 704434
rect 58383 704376 64638 704378
rect 58383 704373 58449 704376
rect 64578 703860 64638 704376
rect 676290 703107 676350 703222
rect 676239 703102 676350 703107
rect 676239 703046 676244 703102
rect 676300 703046 676350 703102
rect 676239 703044 676350 703046
rect 676239 703041 676305 703044
rect 676239 702956 676305 702959
rect 676239 702954 676350 702956
rect 676239 702898 676244 702954
rect 676300 702898 676350 702954
rect 676239 702893 676350 702898
rect 676290 702778 676350 702893
rect 58767 702660 58833 702663
rect 64578 702660 64638 702678
rect 58767 702658 64638 702660
rect 58767 702602 58772 702658
rect 58828 702602 64638 702658
rect 58767 702600 64638 702602
rect 58767 702597 58833 702600
rect 676047 702216 676113 702219
rect 676047 702214 676320 702216
rect 676047 702158 676052 702214
rect 676108 702158 676320 702214
rect 676047 702156 676320 702158
rect 676047 702153 676113 702156
rect 42831 702068 42897 702071
rect 42831 702066 64638 702068
rect 42831 702010 42836 702066
rect 42892 702010 64638 702066
rect 42831 702008 64638 702010
rect 42831 702005 42897 702008
rect 64578 701496 64638 702008
rect 679746 701627 679806 701742
rect 679695 701622 679806 701627
rect 679695 701566 679700 701622
rect 679756 701566 679806 701622
rect 679695 701564 679806 701566
rect 679695 701561 679761 701564
rect 40378 701266 40384 701330
rect 40448 701328 40454 701330
rect 41775 701328 41841 701331
rect 40448 701326 41841 701328
rect 40448 701270 41780 701326
rect 41836 701270 41841 701326
rect 40448 701268 41841 701270
rect 40448 701266 40454 701268
rect 41775 701265 41841 701268
rect 679746 700887 679806 701224
rect 58671 700884 58737 700887
rect 676239 700884 676305 700887
rect 58671 700882 64638 700884
rect 58671 700826 58676 700882
rect 58732 700826 64638 700882
rect 58671 700824 64638 700826
rect 58671 700821 58737 700824
rect 64578 700314 64638 700824
rect 676239 700882 676350 700884
rect 676239 700826 676244 700882
rect 676300 700826 676350 700882
rect 676239 700821 676350 700826
rect 679695 700882 679806 700887
rect 679695 700826 679700 700882
rect 679756 700826 679806 700882
rect 679695 700824 679806 700826
rect 679695 700821 679761 700824
rect 676290 700706 676350 700821
rect 676290 700147 676350 700262
rect 676239 700142 676350 700147
rect 676239 700086 676244 700142
rect 676300 700086 676350 700142
rect 676239 700084 676350 700086
rect 676239 700081 676305 700084
rect 676047 699774 676113 699777
rect 676047 699772 676320 699774
rect 676047 699716 676052 699772
rect 676108 699716 676320 699772
rect 676047 699714 676320 699716
rect 676047 699711 676113 699714
rect 59247 699700 59313 699703
rect 59247 699698 64638 699700
rect 59247 699642 59252 699698
rect 59308 699642 64638 699698
rect 59247 699640 64638 699642
rect 59247 699637 59313 699640
rect 64578 699132 64638 699640
rect 676047 699256 676113 699259
rect 676047 699254 676320 699256
rect 676047 699198 676052 699254
rect 676108 699198 676320 699254
rect 676047 699196 676320 699198
rect 676047 699193 676113 699196
rect 676090 698898 676096 698962
rect 676160 698960 676166 698962
rect 676160 698900 676350 698960
rect 676160 698898 676166 698900
rect 676290 698782 676350 698900
rect 58863 698516 58929 698519
rect 58863 698514 64638 698516
rect 58863 698458 58868 698514
rect 58924 698458 64638 698514
rect 58863 698456 64638 698458
rect 58863 698453 58929 698456
rect 64578 697950 64638 698456
rect 676047 698220 676113 698223
rect 676047 698218 676320 698220
rect 676047 698162 676052 698218
rect 676108 698162 676320 698218
rect 676047 698160 676320 698162
rect 676047 698157 676113 698160
rect 674746 697714 674752 697778
rect 674816 697776 674822 697778
rect 674816 697716 676320 697776
rect 674816 697714 674822 697716
rect 676239 697480 676305 697483
rect 676239 697478 676350 697480
rect 676239 697422 676244 697478
rect 676300 697422 676350 697478
rect 676239 697417 676350 697422
rect 676290 697302 676350 697417
rect 675951 696740 676017 696743
rect 675951 696738 676320 696740
rect 675951 696682 675956 696738
rect 676012 696682 676320 696738
rect 675951 696680 676320 696682
rect 675951 696677 676017 696680
rect 676047 696222 676113 696225
rect 676047 696220 676320 696222
rect 676047 696164 676052 696220
rect 676108 696164 676320 696220
rect 676047 696162 676320 696164
rect 676047 696159 676113 696162
rect 674554 695790 674560 695854
rect 674624 695852 674630 695854
rect 674624 695792 676320 695852
rect 674624 695790 674630 695792
rect 675898 695198 675904 695262
rect 675968 695260 675974 695262
rect 675968 695200 676320 695260
rect 675968 695198 675974 695200
rect 675514 695050 675520 695114
rect 675584 695112 675590 695114
rect 675584 695052 676350 695112
rect 675584 695050 675590 695052
rect 676290 694712 676350 695052
rect 676239 694520 676305 694523
rect 676239 694518 676350 694520
rect 676239 694462 676244 694518
rect 676300 694462 676350 694518
rect 676239 694457 676350 694462
rect 676290 694342 676350 694457
rect 676047 693780 676113 693783
rect 676047 693778 676320 693780
rect 676047 693722 676052 693778
rect 676108 693722 676320 693778
rect 676047 693720 676320 693722
rect 676047 693717 676113 693720
rect 674362 693126 674368 693190
rect 674432 693188 674438 693190
rect 674432 693128 676320 693188
rect 674432 693126 674438 693128
rect 676047 692818 676113 692821
rect 676047 692816 676320 692818
rect 676047 692760 676052 692816
rect 676108 692760 676320 692816
rect 676047 692758 676320 692760
rect 676047 692755 676113 692758
rect 677050 692534 677056 692598
rect 677120 692534 677126 692598
rect 677058 692270 677118 692534
rect 679938 691563 679998 691678
rect 679938 691558 680049 691563
rect 679938 691502 679988 691558
rect 680044 691502 680049 691558
rect 679938 691500 680049 691502
rect 679983 691497 680049 691500
rect 679746 690971 679806 691308
rect 679746 690966 679857 690971
rect 679983 690968 680049 690971
rect 679746 690910 679796 690966
rect 679852 690910 679857 690966
rect 679746 690908 679857 690910
rect 679791 690905 679857 690908
rect 679938 690966 680049 690968
rect 679938 690910 679988 690966
rect 680044 690910 680049 690966
rect 679938 690905 680049 690910
rect 679938 690790 679998 690905
rect 679791 690524 679857 690527
rect 679746 690522 679857 690524
rect 679746 690466 679796 690522
rect 679852 690466 679857 690522
rect 679746 690461 679857 690466
rect 679746 690198 679806 690461
rect 649986 689488 650046 689980
rect 655215 689488 655281 689491
rect 649986 689486 655281 689488
rect 649986 689430 655220 689486
rect 655276 689430 655281 689486
rect 649986 689428 655281 689430
rect 655215 689425 655281 689428
rect 649986 688452 650046 688798
rect 655407 688452 655473 688455
rect 649986 688450 655473 688452
rect 649986 688394 655412 688450
rect 655468 688394 655473 688450
rect 649986 688392 655473 688394
rect 655407 688389 655473 688392
rect 41775 688304 41841 688307
rect 41568 688302 41841 688304
rect 41568 688246 41780 688302
rect 41836 688246 41841 688302
rect 41568 688244 41841 688246
rect 41775 688241 41841 688244
rect 41538 687567 41598 687682
rect 41538 687562 41649 687567
rect 41538 687506 41588 687562
rect 41644 687506 41649 687562
rect 41538 687504 41649 687506
rect 41583 687501 41649 687504
rect 41775 687268 41841 687271
rect 41568 687266 41841 687268
rect 41568 687210 41780 687266
rect 41836 687210 41841 687266
rect 41568 687208 41841 687210
rect 41775 687205 41841 687208
rect 649986 687120 650046 687616
rect 655599 687120 655665 687123
rect 649986 687118 655665 687120
rect 649986 687062 655604 687118
rect 655660 687062 655665 687118
rect 649986 687060 655665 687062
rect 655599 687057 655665 687060
rect 41583 686972 41649 686975
rect 41538 686970 41649 686972
rect 41538 686914 41588 686970
rect 41644 686914 41649 686970
rect 41538 686909 41649 686914
rect 41538 686794 41598 686909
rect 41538 686087 41598 686202
rect 41538 686082 41649 686087
rect 41538 686026 41588 686082
rect 41644 686026 41649 686082
rect 41538 686024 41649 686026
rect 41583 686021 41649 686024
rect 649986 685936 650046 686434
rect 656367 685936 656433 685939
rect 649986 685934 656433 685936
rect 649986 685878 656372 685934
rect 656428 685878 656433 685934
rect 649986 685876 656433 685878
rect 656367 685873 656433 685876
rect 40386 685494 40446 685684
rect 674170 685578 674176 685642
rect 674240 685640 674246 685642
rect 675375 685640 675441 685643
rect 674240 685638 675441 685640
rect 674240 685582 675380 685638
rect 675436 685582 675441 685638
rect 674240 685580 675441 685582
rect 674240 685578 674246 685580
rect 675375 685577 675441 685580
rect 40378 685430 40384 685494
rect 40448 685430 40454 685494
rect 41775 685344 41841 685347
rect 41568 685342 41841 685344
rect 41568 685286 41780 685342
rect 41836 685286 41841 685342
rect 41568 685284 41841 685286
rect 41775 685281 41841 685284
rect 649986 684752 650046 685252
rect 655983 684752 656049 684755
rect 649986 684750 656049 684752
rect 41538 684607 41598 684722
rect 649986 684694 655988 684750
rect 656044 684694 656049 684750
rect 649986 684692 656049 684694
rect 655983 684689 656049 684692
rect 41538 684602 41649 684607
rect 41538 684546 41588 684602
rect 41644 684546 41649 684602
rect 41538 684544 41649 684546
rect 41583 684541 41649 684544
rect 675759 684456 675825 684459
rect 675898 684456 675904 684458
rect 675759 684454 675904 684456
rect 675759 684398 675764 684454
rect 675820 684398 675904 684454
rect 675759 684396 675904 684398
rect 675759 684393 675825 684396
rect 675898 684394 675904 684396
rect 675968 684394 675974 684458
rect 41775 684160 41841 684163
rect 41568 684158 41841 684160
rect 41568 684102 41780 684158
rect 41836 684102 41841 684158
rect 41568 684100 41841 684102
rect 41775 684097 41841 684100
rect 40770 683422 40830 683834
rect 649986 683568 650046 684070
rect 654447 683568 654513 683571
rect 649986 683566 654513 683568
rect 649986 683510 654452 683566
rect 654508 683510 654513 683566
rect 649986 683508 654513 683510
rect 654447 683505 654513 683508
rect 40762 683358 40768 683422
rect 40832 683358 40838 683422
rect 41775 683272 41841 683275
rect 41568 683270 41841 683272
rect 41568 683214 41780 683270
rect 41836 683214 41841 683270
rect 41568 683212 41841 683214
rect 41775 683209 41841 683212
rect 675567 682682 675633 682683
rect 675514 682680 675520 682682
rect 40578 682534 40638 682650
rect 675476 682620 675520 682680
rect 675584 682678 675633 682682
rect 675628 682622 675633 682678
rect 675514 682618 675520 682620
rect 675584 682618 675633 682622
rect 675567 682617 675633 682618
rect 40570 682470 40576 682534
rect 40640 682470 40646 682534
rect 41154 681942 41214 682280
rect 41146 681878 41152 681942
rect 41216 681878 41222 681942
rect 41914 681792 41920 681794
rect 41568 681732 41920 681792
rect 41914 681730 41920 681732
rect 41984 681730 41990 681794
rect 42255 681200 42321 681203
rect 41568 681198 42321 681200
rect 41568 681142 42260 681198
rect 42316 681142 42321 681198
rect 41568 681140 42321 681142
rect 42255 681137 42321 681140
rect 40962 680462 41022 680800
rect 40954 680398 40960 680462
rect 41024 680398 41030 680462
rect 42298 680312 42304 680314
rect 41568 680252 42304 680312
rect 42298 680250 42304 680252
rect 42368 680250 42374 680314
rect 42106 679720 42112 679722
rect 41568 679660 42112 679720
rect 42106 679658 42112 679660
rect 42176 679658 42182 679722
rect 41538 679131 41598 679246
rect 41538 679126 41649 679131
rect 41538 679070 41588 679126
rect 41644 679070 41649 679126
rect 41538 679068 41649 679070
rect 41583 679065 41649 679068
rect 41722 678832 41728 678834
rect 41568 678772 41728 678832
rect 41722 678770 41728 678772
rect 41792 678770 41798 678834
rect 675759 678388 675825 678391
rect 676090 678388 676096 678390
rect 675759 678386 676096 678388
rect 675759 678330 675764 678386
rect 675820 678330 676096 678386
rect 675759 678328 676096 678330
rect 675759 678325 675825 678328
rect 676090 678326 676096 678328
rect 676160 678326 676166 678390
rect 42298 678240 42304 678242
rect 41568 678180 42304 678240
rect 42298 678178 42304 678180
rect 42368 678178 42374 678242
rect 41538 677502 41598 677766
rect 41530 677438 41536 677502
rect 41600 677438 41606 677502
rect 41775 677278 41841 677281
rect 41568 677276 41841 677278
rect 41568 677220 41780 677276
rect 41836 677220 41841 677276
rect 41568 677218 41841 677220
rect 41775 677215 41841 677218
rect 674319 676908 674385 676911
rect 677050 676908 677056 676910
rect 674319 676906 677056 676908
rect 674319 676850 674324 676906
rect 674380 676850 677056 676906
rect 674319 676848 677056 676850
rect 674319 676845 674385 676848
rect 677050 676846 677056 676848
rect 677120 676846 677126 676910
rect 41775 676760 41841 676763
rect 41568 676758 41841 676760
rect 41568 676702 41780 676758
rect 41836 676702 41841 676758
rect 41568 676700 41841 676702
rect 41775 676697 41841 676700
rect 28866 676023 28926 676286
rect 28815 676018 28926 676023
rect 28815 675962 28820 676018
rect 28876 675962 28926 676018
rect 28815 675960 28926 675962
rect 28815 675957 28881 675960
rect 41775 675798 41841 675801
rect 41568 675796 41841 675798
rect 41568 675740 41780 675796
rect 41836 675740 41841 675796
rect 41568 675738 41841 675740
rect 41775 675735 41841 675738
rect 28815 675576 28881 675579
rect 28815 675574 28926 675576
rect 28815 675518 28820 675574
rect 28876 675518 28926 675574
rect 28815 675513 28926 675518
rect 28866 675250 28926 675513
rect 674362 673294 674368 673358
rect 674432 673356 674438 673358
rect 675471 673356 675537 673359
rect 674432 673354 675537 673356
rect 674432 673298 675476 673354
rect 675532 673298 675537 673354
rect 674432 673296 675537 673298
rect 674432 673294 674438 673296
rect 675471 673293 675537 673296
rect 674554 671370 674560 671434
rect 674624 671432 674630 671434
rect 675279 671432 675345 671435
rect 674624 671430 675345 671432
rect 674624 671374 675284 671430
rect 675340 671374 675345 671430
rect 674624 671372 675345 671374
rect 674624 671370 674630 671372
rect 675279 671369 675345 671372
rect 41530 668558 41536 668622
rect 41600 668620 41606 668622
rect 42927 668620 42993 668623
rect 41600 668618 42993 668620
rect 41600 668562 42932 668618
rect 42988 668562 42993 668618
rect 41600 668560 42993 668562
rect 41600 668558 41606 668560
rect 42927 668557 42993 668560
rect 41914 668410 41920 668474
rect 41984 668472 41990 668474
rect 42831 668472 42897 668475
rect 41984 668470 42897 668472
rect 41984 668414 42836 668470
rect 42892 668414 42897 668470
rect 41984 668412 42897 668414
rect 41984 668410 41990 668412
rect 42831 668409 42897 668412
rect 41722 668262 41728 668326
rect 41792 668324 41798 668326
rect 42735 668324 42801 668327
rect 41792 668322 42801 668324
rect 41792 668266 42740 668322
rect 42796 668266 42801 668322
rect 41792 668264 42801 668266
rect 41792 668262 41798 668264
rect 42735 668261 42801 668264
rect 42298 666190 42304 666254
rect 42368 666252 42374 666254
rect 43023 666252 43089 666255
rect 42368 666250 43089 666252
rect 42368 666194 43028 666250
rect 43084 666194 43089 666250
rect 42368 666192 43089 666194
rect 42368 666190 42374 666192
rect 43023 666189 43089 666192
rect 42490 665450 42496 665514
rect 42560 665512 42566 665514
rect 43119 665512 43185 665515
rect 42560 665510 43185 665512
rect 42560 665454 43124 665510
rect 43180 665454 43185 665510
rect 42560 665452 43185 665454
rect 42560 665450 42566 665452
rect 43119 665449 43185 665452
rect 42106 665302 42112 665366
rect 42176 665364 42182 665366
rect 42735 665364 42801 665367
rect 42176 665362 42801 665364
rect 42176 665306 42740 665362
rect 42796 665306 42801 665362
rect 42176 665304 42801 665306
rect 42176 665302 42182 665304
rect 42735 665301 42801 665304
rect 40762 664266 40768 664330
rect 40832 664328 40838 664330
rect 42927 664328 42993 664331
rect 40832 664326 42993 664328
rect 40832 664270 42932 664326
rect 42988 664270 42993 664326
rect 40832 664268 42993 664270
rect 40832 664266 40838 664268
rect 42927 664265 42993 664268
rect 40954 663970 40960 664034
rect 41024 664032 41030 664034
rect 42831 664032 42897 664035
rect 41024 664030 42897 664032
rect 41024 663974 42836 664030
rect 42892 663974 42897 664030
rect 41024 663972 42897 663974
rect 41024 663970 41030 663972
rect 42831 663969 42897 663972
rect 41146 662490 41152 662554
rect 41216 662552 41222 662554
rect 41216 662492 42366 662552
rect 41216 662490 41222 662492
rect 42306 662407 42366 662492
rect 42306 662402 42417 662407
rect 42306 662346 42356 662402
rect 42412 662346 42417 662402
rect 42306 662344 42417 662346
rect 42351 662341 42417 662344
rect 40570 661454 40576 661518
rect 40640 661516 40646 661518
rect 43023 661516 43089 661519
rect 40640 661514 43089 661516
rect 40640 661458 43028 661514
rect 43084 661458 43089 661514
rect 40640 661456 43089 661458
rect 40640 661454 40646 661456
rect 43023 661453 43089 661456
rect 59631 661220 59697 661223
rect 59631 661218 64638 661220
rect 59631 661162 59636 661218
rect 59692 661162 64638 661218
rect 59631 661160 64638 661162
rect 59631 661157 59697 661160
rect 64578 660638 64638 661160
rect 58767 659444 58833 659447
rect 64578 659444 64638 659456
rect 58767 659442 64638 659444
rect 58767 659386 58772 659442
rect 58828 659386 64638 659442
rect 58767 659384 64638 659386
rect 58767 659381 58833 659384
rect 45039 658852 45105 658855
rect 676143 658852 676209 658855
rect 676290 658852 676350 659118
rect 45039 658850 64638 658852
rect 45039 658794 45044 658850
rect 45100 658794 64638 658850
rect 45039 658792 64638 658794
rect 45039 658789 45105 658792
rect 64578 658274 64638 658792
rect 676143 658850 676350 658852
rect 676143 658794 676148 658850
rect 676204 658794 676350 658850
rect 676143 658792 676350 658794
rect 676143 658789 676209 658792
rect 676290 658263 676350 658526
rect 676290 658258 676401 658263
rect 676290 658202 676340 658258
rect 676396 658202 676401 658258
rect 676290 658200 676401 658202
rect 676335 658197 676401 658200
rect 676290 657819 676350 657934
rect 676239 657814 676350 657819
rect 676239 657758 676244 657814
rect 676300 657758 676350 657814
rect 676239 657756 676350 657758
rect 676239 657753 676305 657756
rect 59151 657668 59217 657671
rect 59151 657666 64638 657668
rect 59151 657610 59156 657666
rect 59212 657610 64638 657666
rect 59151 657608 64638 657610
rect 59151 657605 59217 657608
rect 64578 657092 64638 657608
rect 676047 657594 676113 657597
rect 676047 657592 676320 657594
rect 676047 657536 676052 657592
rect 676108 657536 676320 657592
rect 676047 657534 676320 657536
rect 676047 657531 676113 657534
rect 676047 657076 676113 657079
rect 676047 657074 676320 657076
rect 676047 657018 676052 657074
rect 676108 657018 676320 657074
rect 676047 657016 676320 657018
rect 676047 657013 676113 657016
rect 58191 656484 58257 656487
rect 676047 656484 676113 656487
rect 58191 656482 64638 656484
rect 58191 656426 58196 656482
rect 58252 656426 64638 656482
rect 58191 656424 64638 656426
rect 58191 656421 58257 656424
rect 64578 655910 64638 656424
rect 676047 656482 676320 656484
rect 676047 656426 676052 656482
rect 676108 656426 676320 656482
rect 676047 656424 676320 656426
rect 676047 656421 676113 656424
rect 676047 656114 676113 656117
rect 676047 656112 676320 656114
rect 676047 656056 676052 656112
rect 676108 656056 676320 656112
rect 676047 656054 676320 656056
rect 676047 656051 676113 656054
rect 676239 655744 676305 655747
rect 676239 655742 676350 655744
rect 676239 655686 676244 655742
rect 676300 655686 676350 655742
rect 676239 655681 676350 655686
rect 676290 655566 676350 655681
rect 58383 655300 58449 655303
rect 58383 655298 64638 655300
rect 58383 655242 58388 655298
rect 58444 655242 64638 655298
rect 58383 655240 64638 655242
rect 58383 655237 58449 655240
rect 64578 654728 64638 655240
rect 676290 654859 676350 654974
rect 676239 654854 676350 654859
rect 676239 654798 676244 654854
rect 676300 654798 676350 654854
rect 676239 654796 676350 654798
rect 676239 654793 676305 654796
rect 675706 654498 675712 654562
rect 675776 654560 675782 654562
rect 675776 654500 676320 654560
rect 675776 654498 675782 654500
rect 675567 654116 675633 654119
rect 675567 654114 676320 654116
rect 675567 654058 675572 654114
rect 675628 654058 676320 654114
rect 675567 654056 676320 654058
rect 675567 654053 675633 654056
rect 674938 653462 674944 653526
rect 675008 653524 675014 653526
rect 675008 653464 676320 653524
rect 675008 653462 675014 653464
rect 675322 653018 675328 653082
rect 675392 653080 675398 653082
rect 675392 653020 676320 653080
rect 675392 653018 675398 653020
rect 676047 652562 676113 652565
rect 676047 652560 676320 652562
rect 676047 652504 676052 652560
rect 676108 652504 676320 652560
rect 676047 652502 676320 652504
rect 676047 652499 676113 652502
rect 675471 652044 675537 652047
rect 675471 652042 676320 652044
rect 675471 651986 675476 652042
rect 675532 651986 676320 652042
rect 675471 651984 676320 651986
rect 675471 651981 675537 651984
rect 676290 651454 676350 651570
rect 676282 651390 676288 651454
rect 676352 651390 676358 651454
rect 676474 651390 676480 651454
rect 676544 651390 676550 651454
rect 676482 651052 676542 651390
rect 673978 650502 673984 650566
rect 674048 650564 674054 650566
rect 674048 650504 676320 650564
rect 674048 650502 674054 650504
rect 676047 650120 676113 650123
rect 676047 650118 676320 650120
rect 676047 650062 676052 650118
rect 676108 650062 676320 650118
rect 676047 650060 676320 650062
rect 676047 650057 676113 650060
rect 677050 649762 677056 649826
rect 677120 649762 677126 649826
rect 677058 649498 677118 649762
rect 676239 649232 676305 649235
rect 676239 649230 676350 649232
rect 676239 649174 676244 649230
rect 676300 649174 676350 649230
rect 676239 649169 676350 649174
rect 676290 649054 676350 649169
rect 676858 648726 676864 648790
rect 676928 648726 676934 648790
rect 676866 648610 676926 648726
rect 676047 648048 676113 648051
rect 676047 648046 676320 648048
rect 676047 647990 676052 648046
rect 676108 647990 676320 648046
rect 676047 647988 676320 647990
rect 676047 647985 676113 647988
rect 679746 647311 679806 647500
rect 679746 647306 679857 647311
rect 679746 647250 679796 647306
rect 679852 647250 679857 647306
rect 679746 647248 679857 647250
rect 679791 647245 679857 647248
rect 685506 646867 685566 647130
rect 679791 646864 679857 646867
rect 679746 646862 679857 646864
rect 679746 646806 679796 646862
rect 679852 646806 679857 646862
rect 679746 646801 679857 646806
rect 685455 646862 685566 646867
rect 685455 646806 685460 646862
rect 685516 646806 685566 646862
rect 685455 646804 685566 646806
rect 685455 646801 685521 646804
rect 679746 646538 679806 646801
rect 685455 646420 685521 646423
rect 685455 646418 685566 646420
rect 685455 646362 685460 646418
rect 685516 646362 685566 646418
rect 685455 646357 685566 646362
rect 685506 646020 685566 646357
rect 41538 644943 41598 645058
rect 41538 644938 41649 644943
rect 41538 644882 41588 644938
rect 41644 644882 41649 644938
rect 41538 644880 41649 644882
rect 41583 644877 41649 644880
rect 41538 644351 41598 644466
rect 41538 644346 41649 644351
rect 41538 644290 41588 644346
rect 41644 644290 41649 644346
rect 41538 644288 41649 644290
rect 41583 644285 41649 644288
rect 41775 644052 41841 644055
rect 41568 644050 41841 644052
rect 41568 643994 41780 644050
rect 41836 643994 41841 644050
rect 41568 643992 41841 643994
rect 41775 643989 41841 643992
rect 41583 643756 41649 643759
rect 41538 643754 41649 643756
rect 41538 643698 41588 643754
rect 41644 643698 41649 643754
rect 41538 643693 41649 643698
rect 41538 643578 41598 643693
rect 649986 643016 650046 643558
rect 655119 643016 655185 643019
rect 649986 643014 655185 643016
rect 41538 642871 41598 642986
rect 649986 642958 655124 643014
rect 655180 642958 655185 643014
rect 649986 642956 655185 642958
rect 655119 642953 655185 642956
rect 41538 642866 41649 642871
rect 41538 642810 41588 642866
rect 41644 642810 41649 642866
rect 41538 642808 41649 642810
rect 41583 642805 41649 642808
rect 40386 642278 40446 642542
rect 655311 642424 655377 642427
rect 649986 642422 655377 642424
rect 649986 642366 655316 642422
rect 655372 642366 655377 642422
rect 649986 642364 655377 642366
rect 655311 642361 655377 642364
rect 40378 642214 40384 642278
rect 40448 642214 40454 642278
rect 40570 642214 40576 642278
rect 40640 642276 40646 642278
rect 43119 642276 43185 642279
rect 40640 642274 43185 642276
rect 40640 642218 43124 642274
rect 43180 642218 43185 642274
rect 40640 642216 43185 642218
rect 40640 642214 40646 642216
rect 41538 642098 41598 642216
rect 43119 642213 43185 642216
rect 675759 641684 675825 641687
rect 676666 641684 676672 641686
rect 675759 641682 676672 641684
rect 675759 641626 675764 641682
rect 675820 641626 676672 641682
rect 675759 641624 676672 641626
rect 675759 641621 675825 641624
rect 676666 641622 676672 641624
rect 676736 641622 676742 641686
rect 41538 641391 41598 641506
rect 41538 641386 41649 641391
rect 41538 641330 41588 641386
rect 41644 641330 41649 641386
rect 41538 641328 41649 641330
rect 41583 641325 41649 641328
rect 43407 641092 43473 641095
rect 41538 641090 43473 641092
rect 41538 641034 43412 641090
rect 43468 641034 43473 641090
rect 41538 641032 43473 641034
rect 41538 640988 41598 641032
rect 43407 641029 43473 641032
rect 649986 640796 650046 641194
rect 655503 640796 655569 640799
rect 649986 640794 655569 640796
rect 649986 640738 655508 640794
rect 655564 640738 655569 640794
rect 649986 640736 655569 640738
rect 655503 640733 655569 640736
rect 654159 640648 654225 640651
rect 649986 640646 654225 640648
rect 40770 640354 40830 640618
rect 649986 640590 654164 640646
rect 654220 640590 654225 640646
rect 649986 640588 654225 640590
rect 40762 640290 40768 640354
rect 40832 640290 40838 640354
rect 41538 639911 41598 640026
rect 649986 640012 650046 640588
rect 654159 640585 654225 640588
rect 675130 640290 675136 640354
rect 675200 640352 675206 640354
rect 675471 640352 675537 640355
rect 675200 640350 675537 640352
rect 675200 640294 675476 640350
rect 675532 640294 675537 640350
rect 675200 640292 675537 640294
rect 675200 640290 675206 640292
rect 675471 640289 675537 640292
rect 673978 640142 673984 640206
rect 674048 640204 674054 640206
rect 675183 640204 675249 640207
rect 674048 640202 675249 640204
rect 674048 640146 675188 640202
rect 675244 640146 675249 640202
rect 674048 640144 675249 640146
rect 674048 640142 674054 640144
rect 675183 640141 675249 640144
rect 41538 639906 41649 639911
rect 41538 639850 41588 639906
rect 41644 639850 41649 639906
rect 41538 639848 41649 639850
rect 41583 639845 41649 639848
rect 40578 639318 40638 639434
rect 40570 639254 40576 639318
rect 40640 639254 40646 639318
rect 41346 638726 41406 639138
rect 41338 638662 41344 638726
rect 41408 638662 41414 638726
rect 42682 638576 42688 638578
rect 41568 638516 42688 638576
rect 42682 638514 42688 638516
rect 42752 638514 42758 638578
rect 649986 638280 650046 638830
rect 674746 638366 674752 638430
rect 674816 638428 674822 638430
rect 675471 638428 675537 638431
rect 674816 638426 675537 638428
rect 674816 638370 675476 638426
rect 675532 638370 675537 638426
rect 674816 638368 675537 638370
rect 674816 638366 674822 638368
rect 675471 638365 675537 638368
rect 655791 638280 655857 638283
rect 649986 638278 655857 638280
rect 649986 638222 655796 638278
rect 655852 638222 655857 638278
rect 649986 638220 655857 638222
rect 655791 638217 655857 638220
rect 41871 637984 41937 637987
rect 41568 637982 41937 637984
rect 41568 637926 41876 637982
rect 41932 637926 41937 637982
rect 41568 637924 41937 637926
rect 41871 637921 41937 637924
rect 41538 637244 41598 637584
rect 42298 637244 42304 637246
rect 41538 637184 42304 637244
rect 42298 637182 42304 637184
rect 42368 637182 42374 637246
rect 43066 637096 43072 637098
rect 41568 637036 43072 637096
rect 43066 637034 43072 637036
rect 43136 637034 43142 637098
rect 649986 637096 650046 637648
rect 655887 637096 655953 637099
rect 649986 637094 655953 637096
rect 649986 637038 655892 637094
rect 655948 637038 655953 637094
rect 649986 637036 655953 637038
rect 655887 637033 655953 637036
rect 42106 636504 42112 636506
rect 41568 636444 42112 636504
rect 42106 636442 42112 636444
rect 42176 636442 42182 636506
rect 41775 636134 41841 636137
rect 41568 636132 41841 636134
rect 41568 636076 41780 636132
rect 41836 636076 41841 636132
rect 41568 636074 41841 636076
rect 41775 636071 41841 636074
rect 41722 635616 41728 635618
rect 41568 635556 41728 635616
rect 41722 635554 41728 635556
rect 41792 635554 41798 635618
rect 41914 635024 41920 635026
rect 41568 634964 41920 635024
rect 41914 634962 41920 634964
rect 41984 634962 41990 635026
rect 41538 634286 41598 634550
rect 41530 634222 41536 634286
rect 41600 634222 41606 634286
rect 41775 634136 41841 634139
rect 675375 634138 675441 634139
rect 675322 634136 675328 634138
rect 41568 634134 41841 634136
rect 41568 634078 41780 634134
rect 41836 634078 41841 634134
rect 41568 634076 41841 634078
rect 675284 634076 675328 634136
rect 675392 634134 675441 634138
rect 675436 634078 675441 634134
rect 41775 634073 41841 634076
rect 675322 634074 675328 634076
rect 675392 634074 675441 634078
rect 675375 634073 675441 634074
rect 41775 633544 41841 633547
rect 41568 633542 41841 633544
rect 41568 633486 41780 633542
rect 41836 633486 41841 633542
rect 41568 633484 41841 633486
rect 41775 633481 41841 633484
rect 28866 632807 28926 633070
rect 28815 632802 28926 632807
rect 28815 632746 28820 632802
rect 28876 632746 28926 632802
rect 28815 632744 28926 632746
rect 675759 632804 675825 632807
rect 676858 632804 676864 632806
rect 675759 632802 676864 632804
rect 675759 632746 675764 632802
rect 675820 632746 676864 632802
rect 675759 632744 676864 632746
rect 28815 632741 28881 632744
rect 675759 632741 675825 632744
rect 676858 632742 676864 632744
rect 676928 632742 676934 632806
rect 41775 632582 41841 632585
rect 41568 632580 41841 632582
rect 41568 632524 41780 632580
rect 41836 632524 41841 632580
rect 41568 632522 41841 632524
rect 41775 632519 41841 632522
rect 28815 632360 28881 632363
rect 28815 632358 28926 632360
rect 28815 632302 28820 632358
rect 28876 632302 28926 632358
rect 28815 632297 28926 632302
rect 28866 632034 28926 632297
rect 675759 629104 675825 629107
rect 676282 629104 676288 629106
rect 675759 629102 676288 629104
rect 675759 629046 675764 629102
rect 675820 629046 676288 629102
rect 675759 629044 676288 629046
rect 675759 629041 675825 629044
rect 676282 629042 676288 629044
rect 676352 629042 676358 629106
rect 675759 627328 675825 627331
rect 676474 627328 676480 627330
rect 675759 627326 676480 627328
rect 675759 627270 675764 627326
rect 675820 627270 676480 627326
rect 675759 627268 676480 627270
rect 675759 627265 675825 627268
rect 676474 627266 676480 627268
rect 676544 627266 676550 627330
rect 41530 625934 41536 625998
rect 41600 625996 41606 625998
rect 42927 625996 42993 625999
rect 41600 625994 42993 625996
rect 41600 625938 42932 625994
rect 42988 625938 42993 625994
rect 41600 625936 42993 625938
rect 41600 625934 41606 625936
rect 42927 625933 42993 625936
rect 41722 625046 41728 625110
rect 41792 625108 41798 625110
rect 42831 625108 42897 625111
rect 41792 625106 42897 625108
rect 41792 625050 42836 625106
rect 42892 625050 42897 625106
rect 41792 625048 42897 625050
rect 41792 625046 41798 625048
rect 42831 625045 42897 625048
rect 42106 623862 42112 623926
rect 42176 623924 42182 623926
rect 43023 623924 43089 623927
rect 42176 623922 43089 623924
rect 42176 623866 43028 623922
rect 43084 623866 43089 623922
rect 42176 623864 43089 623866
rect 42176 623862 42182 623864
rect 43023 623861 43089 623864
rect 41914 622086 41920 622150
rect 41984 622148 41990 622150
rect 42831 622148 42897 622151
rect 41984 622146 42897 622148
rect 41984 622090 42836 622146
rect 42892 622090 42897 622146
rect 41984 622088 42897 622090
rect 41984 622086 41990 622088
rect 42831 622085 42897 622088
rect 42298 621938 42304 622002
rect 42368 622000 42374 622002
rect 43119 622000 43185 622003
rect 42368 621998 43185 622000
rect 42368 621942 43124 621998
rect 43180 621942 43185 621998
rect 42368 621940 43185 621942
rect 42368 621938 42374 621940
rect 43119 621937 43185 621940
rect 40762 621346 40768 621410
rect 40832 621408 40838 621410
rect 42927 621408 42993 621411
rect 40832 621406 42993 621408
rect 40832 621350 42932 621406
rect 42988 621350 42993 621406
rect 40832 621348 42993 621350
rect 40832 621346 40838 621348
rect 42927 621345 42993 621348
rect 42159 620816 42225 620819
rect 42682 620816 42688 620818
rect 42159 620814 42688 620816
rect 42159 620758 42164 620814
rect 42220 620758 42688 620814
rect 42159 620756 42688 620758
rect 42159 620753 42225 620756
rect 42682 620754 42688 620756
rect 42752 620754 42758 620818
rect 58959 618004 59025 618007
rect 58959 618002 64638 618004
rect 58959 617946 58964 618002
rect 59020 617946 64638 618002
rect 58959 617944 64638 617946
rect 58959 617941 59025 617944
rect 40570 617646 40576 617710
rect 40640 617708 40646 617710
rect 43023 617708 43089 617711
rect 40640 617706 43089 617708
rect 40640 617650 43028 617706
rect 43084 617650 43089 617706
rect 40640 617648 43089 617650
rect 40640 617646 40646 617648
rect 43023 617645 43089 617648
rect 64578 617416 64638 617944
rect 42159 617264 42225 617267
rect 43066 617264 43072 617266
rect 42159 617262 43072 617264
rect 42159 617206 42164 617262
rect 42220 617206 43072 617262
rect 42159 617204 43072 617206
rect 42159 617201 42225 617204
rect 43066 617202 43072 617204
rect 43136 617202 43142 617266
rect 41338 616610 41344 616674
rect 41408 616672 41414 616674
rect 41775 616672 41841 616675
rect 41408 616670 41841 616672
rect 41408 616614 41780 616670
rect 41836 616614 41841 616670
rect 41408 616612 41841 616614
rect 41408 616610 41414 616612
rect 41775 616609 41841 616612
rect 59631 616228 59697 616231
rect 64578 616228 64638 616234
rect 59631 616226 64638 616228
rect 59631 616170 59636 616226
rect 59692 616170 64638 616226
rect 59631 616168 64638 616170
rect 59631 616165 59697 616168
rect 58191 615636 58257 615639
rect 58191 615634 64638 615636
rect 58191 615578 58196 615634
rect 58252 615578 64638 615634
rect 58191 615576 64638 615578
rect 58191 615573 58257 615576
rect 64578 615052 64638 615576
rect 58959 614452 59025 614455
rect 676143 614452 676209 614455
rect 676290 614452 676350 614718
rect 58959 614450 64638 614452
rect 58959 614394 58964 614450
rect 59020 614394 64638 614450
rect 58959 614392 64638 614394
rect 58959 614389 59025 614392
rect 64578 613870 64638 614392
rect 676143 614450 676350 614452
rect 676143 614394 676148 614450
rect 676204 614394 676350 614450
rect 676143 614392 676350 614394
rect 676143 614389 676209 614392
rect 676047 614156 676113 614159
rect 676047 614154 676320 614156
rect 676047 614098 676052 614154
rect 676108 614098 676320 614154
rect 676047 614096 676320 614098
rect 676047 614093 676113 614096
rect 676239 613860 676305 613863
rect 676239 613858 676350 613860
rect 676239 613802 676244 613858
rect 676300 613802 676350 613858
rect 676239 613797 676350 613802
rect 676290 613534 676350 613797
rect 59631 613268 59697 613271
rect 59631 613266 64638 613268
rect 59631 613210 59636 613266
rect 59692 613210 64638 613266
rect 59631 613208 64638 613210
rect 59631 613205 59697 613208
rect 64578 612688 64638 613208
rect 676047 613194 676113 613197
rect 676047 613192 676320 613194
rect 676047 613136 676052 613192
rect 676108 613136 676320 613192
rect 676047 613134 676320 613136
rect 676047 613131 676113 613134
rect 676047 612676 676113 612679
rect 676047 612674 676320 612676
rect 676047 612618 676052 612674
rect 676108 612618 676320 612674
rect 676047 612616 676320 612618
rect 676047 612613 676113 612616
rect 59535 612084 59601 612087
rect 59535 612082 64638 612084
rect 59535 612026 59540 612082
rect 59596 612026 64638 612082
rect 59535 612024 64638 612026
rect 59535 612021 59601 612024
rect 64578 611506 64638 612024
rect 676290 611939 676350 612054
rect 676239 611934 676350 611939
rect 676239 611878 676244 611934
rect 676300 611878 676350 611934
rect 676239 611876 676350 611878
rect 676239 611873 676305 611876
rect 676047 611714 676113 611717
rect 676047 611712 676320 611714
rect 676047 611656 676052 611712
rect 676108 611656 676320 611712
rect 676047 611654 676320 611656
rect 676047 611651 676113 611654
rect 676047 611196 676113 611199
rect 676047 611194 676320 611196
rect 676047 611138 676052 611194
rect 676108 611138 676320 611194
rect 676047 611136 676320 611138
rect 676047 611133 676113 611136
rect 676047 610604 676113 610607
rect 676047 610602 676320 610604
rect 676047 610546 676052 610602
rect 676108 610546 676320 610602
rect 676047 610544 676320 610546
rect 676047 610541 676113 610544
rect 675898 610098 675904 610162
rect 675968 610160 675974 610162
rect 675968 610100 676320 610160
rect 675968 610098 675974 610100
rect 674362 609654 674368 609718
rect 674432 609716 674438 609718
rect 674432 609656 676320 609716
rect 674432 609654 674438 609656
rect 674170 609062 674176 609126
rect 674240 609124 674246 609126
rect 674240 609064 676320 609124
rect 674240 609062 674246 609064
rect 675514 608618 675520 608682
rect 675584 608680 675590 608682
rect 675584 608620 676320 608680
rect 675584 608618 675590 608620
rect 676090 608470 676096 608534
rect 676160 608532 676166 608534
rect 676160 608472 676350 608532
rect 676160 608470 676166 608472
rect 676290 608132 676350 608472
rect 674554 607582 674560 607646
rect 674624 607644 674630 607646
rect 674624 607584 676320 607644
rect 674624 607582 674630 607584
rect 676047 607200 676113 607203
rect 676047 607198 676320 607200
rect 676047 607142 676052 607198
rect 676108 607142 676320 607198
rect 676047 607140 676320 607142
rect 676047 607137 676113 607140
rect 676047 606682 676113 606685
rect 676047 606680 676320 606682
rect 676047 606624 676052 606680
rect 676108 606624 676320 606680
rect 676047 606622 676320 606624
rect 676047 606619 676113 606622
rect 676239 606312 676305 606315
rect 676239 606310 676350 606312
rect 676239 606254 676244 606310
rect 676300 606254 676350 606310
rect 676239 606249 676350 606254
rect 676290 606134 676350 606249
rect 676047 605720 676113 605723
rect 676047 605718 676320 605720
rect 676047 605662 676052 605718
rect 676108 605662 676320 605718
rect 676047 605660 676320 605662
rect 676047 605657 676113 605660
rect 676047 605128 676113 605131
rect 676047 605126 676320 605128
rect 676047 605070 676052 605126
rect 676108 605070 676320 605126
rect 676047 605068 676320 605070
rect 676047 605065 676113 605068
rect 676047 604684 676113 604687
rect 676047 604682 676320 604684
rect 676047 604626 676052 604682
rect 676108 604626 676320 604682
rect 676047 604624 676320 604626
rect 676047 604621 676113 604624
rect 676239 604388 676305 604391
rect 676239 604386 676350 604388
rect 676239 604330 676244 604386
rect 676300 604330 676350 604386
rect 676239 604325 676350 604330
rect 676290 604210 676350 604325
rect 676047 603648 676113 603651
rect 676047 603646 676320 603648
rect 676047 603590 676052 603646
rect 676108 603590 676320 603646
rect 676047 603588 676320 603590
rect 676047 603585 676113 603588
rect 679938 602911 679998 603100
rect 679938 602906 680049 602911
rect 679938 602850 679988 602906
rect 680044 602850 680049 602906
rect 679938 602848 680049 602850
rect 679983 602845 680049 602848
rect 679746 602467 679806 602730
rect 679746 602462 679857 602467
rect 679983 602464 680049 602467
rect 679746 602406 679796 602462
rect 679852 602406 679857 602462
rect 679746 602404 679857 602406
rect 679791 602401 679857 602404
rect 679938 602462 680049 602464
rect 679938 602406 679988 602462
rect 680044 602406 680049 602462
rect 679938 602401 680049 602406
rect 679938 602138 679998 602401
rect 679791 602020 679857 602023
rect 679746 602018 679857 602020
rect 679746 601962 679796 602018
rect 679852 601962 679857 602018
rect 679746 601957 679857 601962
rect 40335 601726 40401 601727
rect 40335 601724 40384 601726
rect 40292 601722 40384 601724
rect 40292 601666 40340 601722
rect 40292 601664 40384 601666
rect 40335 601662 40384 601664
rect 40448 601662 40454 601726
rect 40335 601661 40401 601662
rect 41538 601579 41598 601842
rect 679746 601620 679806 601957
rect 41538 601574 41649 601579
rect 41538 601518 41588 601574
rect 41644 601518 41649 601574
rect 41538 601516 41649 601518
rect 41583 601513 41649 601516
rect 41775 601428 41841 601431
rect 41568 601426 41841 601428
rect 41568 601370 41780 601426
rect 41836 601370 41841 601426
rect 41568 601368 41841 601370
rect 41775 601365 41841 601368
rect 41775 600836 41841 600839
rect 41568 600834 41841 600836
rect 41568 600778 41780 600834
rect 41836 600778 41841 600834
rect 41568 600776 41841 600778
rect 41775 600773 41841 600776
rect 41775 600392 41841 600395
rect 41568 600390 41841 600392
rect 41568 600334 41780 600390
rect 41836 600334 41841 600390
rect 41568 600332 41841 600334
rect 41775 600329 41841 600332
rect 41775 599874 41841 599877
rect 41568 599872 41841 599874
rect 41568 599816 41780 599872
rect 41836 599816 41841 599872
rect 41568 599814 41841 599816
rect 41775 599811 41841 599814
rect 41775 599356 41841 599359
rect 41568 599354 41841 599356
rect 41568 599298 41780 599354
rect 41836 599298 41841 599354
rect 41568 599296 41841 599298
rect 41775 599293 41841 599296
rect 40386 598767 40446 598882
rect 40335 598762 40446 598767
rect 40335 598706 40340 598762
rect 40396 598706 40446 598762
rect 40335 598704 40446 598706
rect 40335 598701 40401 598704
rect 41775 598394 41841 598397
rect 41568 598392 41841 598394
rect 41568 598336 41780 598392
rect 41836 598336 41841 598392
rect 41568 598334 41841 598336
rect 41775 598331 41841 598334
rect 39759 598024 39825 598027
rect 39759 598022 39870 598024
rect 39759 597966 39764 598022
rect 39820 597966 39870 598022
rect 39759 597961 39870 597966
rect 39810 597846 39870 597961
rect 649986 597876 650046 598336
rect 655215 597876 655281 597879
rect 649986 597874 655281 597876
rect 649986 597818 655220 597874
rect 655276 597818 655281 597874
rect 649986 597816 655281 597818
rect 655215 597813 655281 597816
rect 40578 597138 40638 597402
rect 40570 597074 40576 597138
rect 40640 597074 40646 597138
rect 41538 596695 41598 596810
rect 41538 596690 41649 596695
rect 41538 596634 41588 596690
rect 41644 596634 41649 596690
rect 41538 596632 41649 596634
rect 649986 596692 650046 597154
rect 674170 597074 674176 597138
rect 674240 597136 674246 597138
rect 675375 597136 675441 597139
rect 674240 597134 675441 597136
rect 674240 597078 675380 597134
rect 675436 597078 675441 597134
rect 674240 597076 675441 597078
rect 674240 597074 674246 597076
rect 675375 597073 675441 597076
rect 655407 596692 655473 596695
rect 649986 596690 655473 596692
rect 649986 596634 655412 596690
rect 655468 596634 655473 596690
rect 649986 596632 655473 596634
rect 41583 596629 41649 596632
rect 655407 596629 655473 596632
rect 40386 596102 40446 596366
rect 40378 596038 40384 596102
rect 40448 596038 40454 596102
rect 674554 596038 674560 596102
rect 674624 596100 674630 596102
rect 675471 596100 675537 596103
rect 674624 596098 675537 596100
rect 674624 596042 675476 596098
rect 675532 596042 675537 596098
rect 674624 596040 675537 596042
rect 674624 596038 674630 596040
rect 675471 596037 675537 596040
rect 40770 595658 40830 595922
rect 40762 595594 40768 595658
rect 40832 595594 40838 595658
rect 649986 595508 650046 595972
rect 655599 595508 655665 595511
rect 649986 595506 655665 595508
rect 649986 595450 655604 595506
rect 655660 595450 655665 595506
rect 649986 595448 655665 595450
rect 655599 595445 655665 595448
rect 42874 595360 42880 595362
rect 41568 595300 42880 595360
rect 42874 595298 42880 595300
rect 42944 595298 42950 595362
rect 654543 595360 654609 595363
rect 649986 595358 654609 595360
rect 649986 595302 654548 595358
rect 654604 595302 654609 595358
rect 649986 595300 654609 595302
rect 41871 594842 41937 594845
rect 41568 594840 41937 594842
rect 41568 594784 41876 594840
rect 41932 594784 41937 594840
rect 649986 594790 650046 595300
rect 654543 595297 654609 595300
rect 41568 594782 41937 594784
rect 41871 594779 41937 594782
rect 40962 594178 41022 594442
rect 40954 594114 40960 594178
rect 41024 594114 41030 594178
rect 674938 593966 674944 594030
rect 675008 594028 675014 594030
rect 675471 594028 675537 594031
rect 675008 594026 675537 594028
rect 675008 593970 675476 594026
rect 675532 593970 675537 594026
rect 675008 593968 675537 593970
rect 675008 593966 675014 593968
rect 675471 593965 675537 593968
rect 42106 593880 42112 593882
rect 41568 593820 42112 593880
rect 42106 593818 42112 593820
rect 42176 593818 42182 593882
rect 42298 593436 42304 593438
rect 41538 593376 42304 593436
rect 41538 593332 41598 593376
rect 42298 593374 42304 593376
rect 42368 593374 42374 593438
rect 649986 593436 650046 593608
rect 654159 593436 654225 593439
rect 649986 593434 654225 593436
rect 649986 593378 654164 593434
rect 654220 593378 654225 593434
rect 649986 593376 654225 593378
rect 654159 593373 654225 593376
rect 41775 592992 41841 592995
rect 41568 592990 41841 592992
rect 41568 592934 41780 592990
rect 41836 592934 41841 592990
rect 41568 592932 41841 592934
rect 41775 592929 41841 592932
rect 41538 592106 41598 592370
rect 41530 592042 41536 592106
rect 41600 592042 41606 592106
rect 649986 591956 650046 592426
rect 654351 591956 654417 591959
rect 649986 591954 654417 591956
rect 649986 591898 654356 591954
rect 654412 591898 654417 591954
rect 649986 591896 654417 591898
rect 654351 591893 654417 591896
rect 41722 591808 41728 591810
rect 41568 591748 41728 591808
rect 41722 591746 41728 591748
rect 41792 591746 41798 591810
rect 41914 591438 41920 591440
rect 41568 591378 41920 591438
rect 41914 591376 41920 591378
rect 41984 591376 41990 591440
rect 41775 590920 41841 590923
rect 41568 590918 41841 590920
rect 41568 590862 41780 590918
rect 41836 590862 41841 590918
rect 41568 590860 41841 590862
rect 41775 590857 41841 590860
rect 41538 590180 41598 590298
rect 41538 590120 41790 590180
rect 28866 589591 28926 589928
rect 41730 589736 41790 590120
rect 28815 589586 28926 589591
rect 28815 589530 28820 589586
rect 28876 589530 28926 589586
rect 28815 589528 28926 589530
rect 41538 589676 41790 589736
rect 675471 589738 675537 589739
rect 675471 589734 675520 589738
rect 675584 589736 675590 589738
rect 675471 589678 675476 589734
rect 28815 589525 28881 589528
rect 41538 589147 41598 589676
rect 675471 589674 675520 589678
rect 675584 589676 675628 589736
rect 675584 589674 675590 589676
rect 675471 589673 675537 589674
rect 28815 589144 28881 589147
rect 28815 589142 28926 589144
rect 28815 589086 28820 589142
rect 28876 589086 28926 589142
rect 28815 589081 28926 589086
rect 41538 589142 41649 589147
rect 41538 589086 41588 589142
rect 41644 589086 41649 589142
rect 41538 589084 41649 589086
rect 41583 589081 41649 589084
rect 28866 588818 28926 589081
rect 675759 584704 675825 584707
rect 675898 584704 675904 584706
rect 675759 584702 675904 584704
rect 675759 584646 675764 584702
rect 675820 584646 675904 584702
rect 675759 584644 675904 584646
rect 675759 584641 675825 584644
rect 675898 584642 675904 584644
rect 675968 584642 675974 584706
rect 41530 583014 41536 583078
rect 41600 583076 41606 583078
rect 42447 583076 42513 583079
rect 41600 583074 42513 583076
rect 41600 583018 42452 583074
rect 42508 583018 42513 583074
rect 41600 583016 42513 583018
rect 41600 583014 41606 583016
rect 42447 583013 42513 583016
rect 675663 582930 675729 582931
rect 675663 582926 675712 582930
rect 675776 582928 675782 582930
rect 675663 582870 675668 582926
rect 675663 582866 675712 582870
rect 675776 582868 675820 582928
rect 675776 582866 675782 582868
rect 675663 582865 675729 582866
rect 41914 582570 41920 582634
rect 41984 582632 41990 582634
rect 43119 582632 43185 582635
rect 41984 582630 43185 582632
rect 41984 582574 43124 582630
rect 43180 582574 43185 582630
rect 41984 582572 43185 582574
rect 41984 582570 41990 582572
rect 43119 582569 43185 582572
rect 42106 581682 42112 581746
rect 42176 581744 42182 581746
rect 42831 581744 42897 581747
rect 42176 581742 42897 581744
rect 42176 581686 42836 581742
rect 42892 581686 42897 581742
rect 42176 581684 42897 581686
rect 42176 581682 42182 581684
rect 42831 581681 42897 581684
rect 42298 580498 42304 580562
rect 42368 580560 42374 580562
rect 43119 580560 43185 580563
rect 42368 580558 43185 580560
rect 42368 580502 43124 580558
rect 43180 580502 43185 580558
rect 42368 580500 43185 580502
rect 42368 580498 42374 580500
rect 43119 580497 43185 580500
rect 42927 579526 42993 579527
rect 42874 579524 42880 579526
rect 42836 579464 42880 579524
rect 42944 579522 42993 579526
rect 42988 579466 42993 579522
rect 42874 579462 42880 579464
rect 42944 579462 42993 579466
rect 42927 579461 42993 579462
rect 41722 578870 41728 578934
rect 41792 578932 41798 578934
rect 42447 578932 42513 578935
rect 41792 578930 42513 578932
rect 41792 578874 42452 578930
rect 42508 578874 42513 578930
rect 41792 578872 42513 578874
rect 41792 578870 41798 578872
rect 42447 578869 42513 578872
rect 40570 576354 40576 576418
rect 40640 576416 40646 576418
rect 43023 576416 43089 576419
rect 40640 576414 43089 576416
rect 40640 576358 43028 576414
rect 43084 576358 43089 576414
rect 40640 576356 43089 576358
rect 40640 576354 40646 576356
rect 43023 576353 43089 576356
rect 40954 576206 40960 576270
rect 41024 576268 41030 576270
rect 42927 576268 42993 576271
rect 41024 576266 42993 576268
rect 41024 576210 42932 576266
rect 42988 576210 42993 576266
rect 41024 576208 42993 576210
rect 41024 576206 41030 576208
rect 42927 576205 42993 576208
rect 40762 576058 40768 576122
rect 40832 576120 40838 576122
rect 42351 576120 42417 576123
rect 40832 576118 42417 576120
rect 40832 576062 42356 576118
rect 42412 576062 42417 576118
rect 40832 576060 42417 576062
rect 40832 576058 40838 576060
rect 42351 576057 42417 576060
rect 58959 574788 59025 574791
rect 58959 574786 64638 574788
rect 58959 574730 58964 574786
rect 59020 574730 64638 574786
rect 58959 574728 64638 574730
rect 58959 574725 59025 574728
rect 64578 574194 64638 574728
rect 40378 573838 40384 573902
rect 40448 573900 40454 573902
rect 42831 573900 42897 573903
rect 40448 573898 42897 573900
rect 40448 573842 42836 573898
rect 42892 573842 42897 573898
rect 40448 573840 42897 573842
rect 40448 573838 40454 573840
rect 42831 573837 42897 573840
rect 59631 573012 59697 573015
rect 59631 573010 64638 573012
rect 59631 572954 59636 573010
rect 59692 572954 64638 573010
rect 59631 572952 64638 572954
rect 59631 572949 59697 572952
rect 45039 572420 45105 572423
rect 45039 572418 64638 572420
rect 45039 572362 45044 572418
rect 45100 572362 64638 572418
rect 45039 572360 64638 572362
rect 45039 572357 45105 572360
rect 64578 571830 64638 572360
rect 58959 571236 59025 571239
rect 58959 571234 64638 571236
rect 58959 571178 58964 571234
rect 59020 571178 64638 571234
rect 58959 571176 64638 571178
rect 58959 571173 59025 571176
rect 64578 570648 64638 571176
rect 60399 570052 60465 570055
rect 60399 570050 64638 570052
rect 60399 569994 60404 570050
rect 60460 569994 64638 570050
rect 60399 569992 64638 569994
rect 60399 569989 60465 569992
rect 64578 569466 64638 569992
rect 676290 569315 676350 569430
rect 676239 569310 676350 569315
rect 676239 569254 676244 569310
rect 676300 569254 676350 569310
rect 676239 569252 676350 569254
rect 676239 569249 676305 569252
rect 59151 568868 59217 568871
rect 59151 568866 64638 568868
rect 59151 568810 59156 568866
rect 59212 568810 64638 568866
rect 59151 568808 64638 568810
rect 59151 568805 59217 568808
rect 64578 568284 64638 568808
rect 676143 568572 676209 568575
rect 676290 568572 676350 568912
rect 676143 568570 676350 568572
rect 676143 568514 676148 568570
rect 676204 568514 676350 568570
rect 676143 568512 676350 568514
rect 676143 568509 676209 568512
rect 676047 568424 676113 568427
rect 676047 568422 676320 568424
rect 676047 568366 676052 568422
rect 676108 568366 676320 568422
rect 676047 568364 676320 568366
rect 676047 568361 676113 568364
rect 679746 567835 679806 567950
rect 679695 567830 679806 567835
rect 679695 567774 679700 567830
rect 679756 567774 679806 567830
rect 679695 567772 679806 567774
rect 679695 567769 679761 567772
rect 676047 567462 676113 567465
rect 676047 567460 676320 567462
rect 676047 567404 676052 567460
rect 676108 567404 676320 567460
rect 676047 567402 676320 567404
rect 676047 567399 676113 567402
rect 674895 567240 674961 567243
rect 676090 567240 676096 567242
rect 674895 567238 676096 567240
rect 674895 567182 674900 567238
rect 674956 567182 676096 567238
rect 674895 567180 676096 567182
rect 674895 567177 674961 567180
rect 676090 567178 676096 567180
rect 676160 567178 676166 567242
rect 676239 567092 676305 567095
rect 676239 567090 676350 567092
rect 676239 567034 676244 567090
rect 676300 567034 676350 567090
rect 676239 567029 676350 567034
rect 676290 566914 676350 567029
rect 676290 566355 676350 566470
rect 676239 566350 676350 566355
rect 676239 566294 676244 566350
rect 676300 566294 676350 566350
rect 676239 566292 676350 566294
rect 676239 566289 676305 566292
rect 676047 565908 676113 565911
rect 676047 565906 676320 565908
rect 676047 565850 676052 565906
rect 676108 565850 676320 565906
rect 676047 565848 676320 565850
rect 676047 565845 676113 565848
rect 676047 565464 676113 565467
rect 676047 565462 676320 565464
rect 676047 565406 676052 565462
rect 676108 565406 676320 565462
rect 676047 565404 676320 565406
rect 676047 565401 676113 565404
rect 675130 564958 675136 565022
rect 675200 565020 675206 565022
rect 675200 564960 676320 565020
rect 675200 564958 675206 564960
rect 676282 564662 676288 564726
rect 676352 564662 676358 564726
rect 676290 564398 676350 564662
rect 676666 564218 676672 564282
rect 676736 564218 676742 564282
rect 676674 563880 676734 564218
rect 674746 563478 674752 563542
rect 674816 563540 674822 563542
rect 674816 563480 676320 563540
rect 674816 563478 674822 563480
rect 675322 562886 675328 562950
rect 675392 562948 675398 562950
rect 675392 562888 676320 562948
rect 675392 562886 675398 562888
rect 676474 562738 676480 562802
rect 676544 562738 676550 562802
rect 676482 562400 676542 562738
rect 673978 561998 673984 562062
rect 674048 562060 674054 562062
rect 674048 562000 676320 562060
rect 674048 561998 674054 562000
rect 676047 561468 676113 561471
rect 676047 561466 676320 561468
rect 676047 561410 676052 561466
rect 676108 561410 676320 561466
rect 676047 561408 676320 561410
rect 676047 561405 676113 561408
rect 676047 560876 676113 560879
rect 676047 560874 676320 560876
rect 676047 560818 676052 560874
rect 676108 560818 676320 560874
rect 676047 560816 676320 560818
rect 676047 560813 676113 560816
rect 676239 560728 676305 560731
rect 676239 560726 676350 560728
rect 676239 560670 676244 560726
rect 676300 560670 676350 560726
rect 676239 560665 676350 560670
rect 676290 560550 676350 560665
rect 676858 560222 676864 560286
rect 676928 560222 676934 560286
rect 676866 559958 676926 560222
rect 676047 559396 676113 559399
rect 676047 559394 676320 559396
rect 676047 559338 676052 559394
rect 676108 559338 676320 559394
rect 676047 559336 676320 559338
rect 676047 559333 676113 559336
rect 676047 559026 676113 559029
rect 676047 559024 676320 559026
rect 676047 558968 676052 559024
rect 676108 558968 676320 559024
rect 676047 558966 676320 558968
rect 676047 558963 676113 558966
rect 676239 558656 676305 558659
rect 676239 558654 676350 558656
rect 676239 558598 676244 558654
rect 676300 558598 676350 558654
rect 676239 558593 676350 558598
rect 676290 558478 676350 558593
rect 679746 557771 679806 557886
rect 679746 557766 679857 557771
rect 679746 557710 679796 557766
rect 679852 557710 679857 557766
rect 679746 557708 679857 557710
rect 679791 557705 679857 557708
rect 685506 557179 685566 557442
rect 679791 557176 679857 557179
rect 679746 557174 679857 557176
rect 679746 557118 679796 557174
rect 679852 557118 679857 557174
rect 679746 557113 679857 557118
rect 685455 557174 685566 557179
rect 685455 557118 685460 557174
rect 685516 557118 685566 557174
rect 685455 557116 685566 557118
rect 685455 557113 685521 557116
rect 679746 556998 679806 557113
rect 685455 556732 685521 556735
rect 685455 556730 685566 556732
rect 685455 556674 685460 556730
rect 685516 556674 685566 556730
rect 685455 556669 685566 556674
rect 685506 556406 685566 556669
rect 649986 553328 650046 553914
rect 655119 553328 655185 553331
rect 649986 553326 655185 553328
rect 649986 553270 655124 553326
rect 655180 553270 655185 553326
rect 649986 553268 655185 553270
rect 655119 553265 655185 553268
rect 674362 552970 674368 553034
rect 674432 553032 674438 553034
rect 675471 553032 675537 553035
rect 674432 553030 675537 553032
rect 674432 552974 675476 553030
rect 675532 552974 675537 553030
rect 674432 552972 675537 552974
rect 674432 552970 674438 552972
rect 675471 552969 675537 552972
rect 649986 552144 650046 552732
rect 673978 552230 673984 552294
rect 674048 552292 674054 552294
rect 675375 552292 675441 552295
rect 674048 552290 675441 552292
rect 674048 552234 675380 552290
rect 675436 552234 675441 552290
rect 674048 552232 675441 552234
rect 674048 552230 674054 552232
rect 675375 552229 675441 552232
rect 655311 552144 655377 552147
rect 649986 552142 655377 552144
rect 649986 552086 655316 552142
rect 655372 552086 655377 552142
rect 649986 552084 655377 552086
rect 655311 552081 655377 552084
rect 675183 551702 675249 551703
rect 675130 551700 675136 551702
rect 675092 551640 675136 551700
rect 675200 551698 675249 551702
rect 675244 551642 675249 551698
rect 675130 551638 675136 551640
rect 675200 551638 675249 551642
rect 675183 551637 675249 551638
rect 649986 551108 650046 551550
rect 655503 551108 655569 551111
rect 649986 551106 655569 551108
rect 649986 551050 655508 551106
rect 655564 551050 655569 551106
rect 649986 551048 655569 551050
rect 655503 551045 655569 551048
rect 653775 550960 653841 550963
rect 649986 550958 653841 550960
rect 649986 550902 653780 550958
rect 653836 550902 653841 550958
rect 649986 550900 653841 550902
rect 649986 550368 650046 550900
rect 653775 550897 653841 550900
rect 674746 550158 674752 550222
rect 674816 550220 674822 550222
rect 675279 550220 675345 550223
rect 674816 550218 675345 550220
rect 674816 550162 675284 550218
rect 675340 550162 675345 550218
rect 674816 550160 675345 550162
rect 674816 550158 674822 550160
rect 675279 550157 675345 550160
rect 649986 548592 650046 549186
rect 656271 548592 656337 548595
rect 649986 548590 656337 548592
rect 649986 548534 656276 548590
rect 656332 548534 656337 548590
rect 649986 548532 656337 548534
rect 656271 548529 656337 548532
rect 649986 547556 650046 548004
rect 654159 547556 654225 547559
rect 649986 547554 654225 547556
rect 649986 547498 654164 547554
rect 654220 547498 654225 547554
rect 649986 547496 654225 547498
rect 654159 547493 654225 547496
rect 675375 545486 675441 545487
rect 675322 545484 675328 545486
rect 675284 545424 675328 545484
rect 675392 545482 675441 545486
rect 675436 545426 675441 545482
rect 675322 545422 675328 545424
rect 675392 545422 675441 545426
rect 675375 545421 675441 545422
rect 675375 544300 675441 544303
rect 676858 544300 676864 544302
rect 675375 544298 676864 544300
rect 675375 544242 675380 544298
rect 675436 544242 676864 544298
rect 675375 544240 676864 544242
rect 675375 544237 675441 544240
rect 676858 544238 676864 544240
rect 676928 544238 676934 544302
rect 675759 540600 675825 540603
rect 676282 540600 676288 540602
rect 675759 540598 676288 540600
rect 675759 540542 675764 540598
rect 675820 540542 676288 540598
rect 675759 540540 676288 540542
rect 675759 540537 675825 540540
rect 676282 540538 676288 540540
rect 676352 540538 676358 540602
rect 40378 540390 40384 540454
rect 40448 540452 40454 540454
rect 41775 540452 41841 540455
rect 40448 540450 41841 540452
rect 40448 540394 41780 540450
rect 41836 540394 41841 540450
rect 40448 540392 41841 540394
rect 40448 540390 40454 540392
rect 41775 540389 41841 540392
rect 40570 538762 40576 538826
rect 40640 538824 40646 538826
rect 41775 538824 41841 538827
rect 40640 538822 41841 538824
rect 40640 538766 41780 538822
rect 41836 538766 41841 538822
rect 40640 538764 41841 538766
rect 40640 538762 40646 538764
rect 41775 538761 41841 538764
rect 675183 538676 675249 538679
rect 677050 538676 677056 538678
rect 675183 538674 677056 538676
rect 675183 538618 675188 538674
rect 675244 538618 677056 538674
rect 675183 538616 677056 538618
rect 675183 538613 675249 538616
rect 677050 538614 677056 538616
rect 677120 538614 677126 538678
rect 40954 536838 40960 536902
rect 41024 536900 41030 536902
rect 41775 536900 41841 536903
rect 41024 536898 41841 536900
rect 41024 536842 41780 536898
rect 41836 536842 41841 536898
rect 41024 536840 41841 536842
rect 41024 536838 41030 536840
rect 41775 536837 41841 536840
rect 41338 534766 41344 534830
rect 41408 534828 41414 534830
rect 41775 534828 41841 534831
rect 41408 534826 41841 534828
rect 41408 534770 41780 534826
rect 41836 534770 41841 534826
rect 41408 534768 41841 534770
rect 41408 534766 41414 534768
rect 41775 534765 41841 534768
rect 40762 534470 40768 534534
rect 40832 534532 40838 534534
rect 41775 534532 41841 534535
rect 40832 534530 41841 534532
rect 40832 534474 41780 534530
rect 41836 534474 41841 534530
rect 40832 534472 41841 534474
rect 40832 534470 40838 534472
rect 41775 534469 41841 534472
rect 41871 533646 41937 533647
rect 41871 533642 41920 533646
rect 41984 533644 41990 533646
rect 41871 533586 41876 533642
rect 41871 533582 41920 533586
rect 41984 533584 42028 533644
rect 41984 533582 41990 533584
rect 41871 533581 41937 533582
rect 57711 531720 57777 531723
rect 57711 531718 64638 531720
rect 57711 531662 57716 531718
rect 57772 531662 64638 531718
rect 57711 531660 64638 531662
rect 57711 531657 57777 531660
rect 41146 531362 41152 531426
rect 41216 531424 41222 531426
rect 41775 531424 41841 531427
rect 41216 531422 41841 531424
rect 41216 531366 41780 531422
rect 41836 531366 41841 531422
rect 41216 531364 41841 531366
rect 41216 531362 41222 531364
rect 41775 531361 41841 531364
rect 64578 531172 64638 531660
rect 41530 530622 41536 530686
rect 41600 530684 41606 530686
rect 41775 530684 41841 530687
rect 41600 530682 41841 530684
rect 41600 530626 41780 530682
rect 41836 530626 41841 530682
rect 41600 530624 41841 530626
rect 41600 530622 41606 530624
rect 41775 530621 41841 530624
rect 57615 530536 57681 530539
rect 57615 530534 64638 530536
rect 57615 530478 57620 530534
rect 57676 530478 64638 530534
rect 57615 530476 64638 530478
rect 57615 530473 57681 530476
rect 41775 530094 41841 530095
rect 41722 530092 41728 530094
rect 41684 530032 41728 530092
rect 41792 530090 41841 530094
rect 41836 530034 41841 530090
rect 41722 530030 41728 530032
rect 41792 530030 41841 530034
rect 41775 530029 41841 530030
rect 64578 529990 64638 530476
rect 42159 529352 42225 529355
rect 42298 529352 42304 529354
rect 42159 529350 42304 529352
rect 42159 529294 42164 529350
rect 42220 529294 42304 529350
rect 42159 529292 42304 529294
rect 42159 529289 42225 529292
rect 42298 529290 42304 529292
rect 42368 529290 42374 529354
rect 45039 529352 45105 529355
rect 45039 529350 64638 529352
rect 45039 529294 45044 529350
rect 45100 529294 64638 529350
rect 45039 529292 64638 529294
rect 45039 529289 45105 529292
rect 64578 528808 64638 529292
rect 42159 527724 42225 527727
rect 42490 527724 42496 527726
rect 42159 527722 42496 527724
rect 42159 527666 42164 527722
rect 42220 527666 42496 527722
rect 42159 527664 42496 527666
rect 42159 527661 42225 527664
rect 42490 527662 42496 527664
rect 42560 527662 42566 527726
rect 42063 527134 42129 527135
rect 42063 527130 42112 527134
rect 42176 527132 42182 527134
rect 58959 527132 59025 527135
rect 64578 527132 64638 527626
rect 42063 527074 42068 527130
rect 42063 527070 42112 527074
rect 42176 527072 42220 527132
rect 58959 527130 64638 527132
rect 58959 527074 58964 527130
rect 59020 527074 64638 527130
rect 58959 527072 64638 527074
rect 42176 527070 42182 527072
rect 42063 527069 42129 527070
rect 58959 527069 59025 527072
rect 42063 526540 42129 526543
rect 42682 526540 42688 526542
rect 42063 526538 42688 526540
rect 42063 526482 42068 526538
rect 42124 526482 42688 526538
rect 42063 526480 42688 526482
rect 42063 526477 42129 526480
rect 42682 526478 42688 526480
rect 42752 526478 42758 526542
rect 58575 525948 58641 525951
rect 64578 525948 64638 526444
rect 58575 525946 64638 525948
rect 58575 525890 58580 525946
rect 58636 525890 64638 525946
rect 58575 525888 64638 525890
rect 58575 525885 58641 525888
rect 59343 524764 59409 524767
rect 64578 524764 64638 525262
rect 676290 525211 676350 525474
rect 676290 525206 676401 525211
rect 676290 525150 676340 525206
rect 676396 525150 676401 525206
rect 676290 525148 676401 525150
rect 676335 525145 676401 525148
rect 59343 524762 64638 524764
rect 59343 524706 59348 524762
rect 59404 524706 64638 524762
rect 59343 524704 64638 524706
rect 676143 524764 676209 524767
rect 676290 524764 676350 524882
rect 676143 524762 676350 524764
rect 676143 524706 676148 524762
rect 676204 524706 676350 524762
rect 676143 524704 676350 524706
rect 59343 524701 59409 524704
rect 676143 524701 676209 524704
rect 676239 524616 676305 524619
rect 676239 524614 676350 524616
rect 676239 524558 676244 524614
rect 676300 524558 676350 524614
rect 676239 524553 676350 524558
rect 676290 524438 676350 524553
rect 676047 524024 676113 524027
rect 676047 524022 676320 524024
rect 676047 523966 676052 524022
rect 676108 523966 676320 524022
rect 676047 523964 676320 523966
rect 676047 523961 676113 523964
rect 676482 523287 676542 523402
rect 676482 523282 676593 523287
rect 676482 523226 676532 523282
rect 676588 523226 676593 523282
rect 676482 523224 676593 523226
rect 676527 523221 676593 523224
rect 676047 522914 676113 522917
rect 676047 522912 676320 522914
rect 676047 522856 676052 522912
rect 676108 522856 676320 522912
rect 676047 522854 676320 522856
rect 676047 522851 676113 522854
rect 676674 522251 676734 522514
rect 676623 522246 676734 522251
rect 676623 522190 676628 522246
rect 676684 522190 676734 522246
rect 676623 522188 676734 522190
rect 676623 522185 676689 522188
rect 676290 521807 676350 521922
rect 676239 521802 676350 521807
rect 676239 521746 676244 521802
rect 676300 521746 676350 521802
rect 676239 521744 676350 521746
rect 676239 521741 676305 521744
rect 676674 521215 676734 521330
rect 676674 521210 676785 521215
rect 676674 521154 676724 521210
rect 676780 521154 676785 521210
rect 676674 521152 676785 521154
rect 676719 521149 676785 521152
rect 674554 521002 674560 521066
rect 674624 521064 674630 521066
rect 674624 521004 676320 521064
rect 674624 521002 674630 521004
rect 675898 520410 675904 520474
rect 675968 520472 675974 520474
rect 675968 520412 676320 520472
rect 675968 520410 675974 520412
rect 674170 519818 674176 519882
rect 674240 519880 674246 519882
rect 674240 519820 676320 519880
rect 674240 519818 674246 519820
rect 674938 519670 674944 519734
rect 675008 519732 675014 519734
rect 675008 519672 676350 519732
rect 675008 519670 675014 519672
rect 676290 519480 676350 519672
rect 675514 518930 675520 518994
rect 675584 518992 675590 518994
rect 675584 518932 676320 518992
rect 675584 518930 675590 518932
rect 675706 518338 675712 518402
rect 675776 518400 675782 518402
rect 675776 518340 676320 518400
rect 675776 518338 675782 518340
rect 676090 518190 676096 518254
rect 676160 518252 676166 518254
rect 676160 518192 676350 518252
rect 676160 518190 676166 518192
rect 676290 518000 676350 518192
rect 676239 517660 676305 517663
rect 676239 517658 676350 517660
rect 676239 517602 676244 517658
rect 676300 517602 676350 517658
rect 676239 517597 676350 517602
rect 676290 517482 676350 517597
rect 676047 516920 676113 516923
rect 676047 516918 676320 516920
rect 676047 516862 676052 516918
rect 676108 516862 676320 516918
rect 676047 516860 676320 516862
rect 676047 516857 676113 516860
rect 676047 516476 676113 516479
rect 676047 516474 676320 516476
rect 676047 516418 676052 516474
rect 676108 516418 676320 516474
rect 676047 516416 676320 516418
rect 676047 516413 676113 516416
rect 676239 516180 676305 516183
rect 676239 516178 676350 516180
rect 676239 516122 676244 516178
rect 676300 516122 676350 516178
rect 676239 516117 676350 516122
rect 676290 516002 676350 516117
rect 676047 515440 676113 515443
rect 676047 515438 676320 515440
rect 676047 515382 676052 515438
rect 676108 515382 676320 515438
rect 676047 515380 676320 515382
rect 676047 515377 676113 515380
rect 676047 514996 676113 514999
rect 676047 514994 676320 514996
rect 676047 514938 676052 514994
rect 676108 514938 676320 514994
rect 676047 514936 676320 514938
rect 676047 514933 676113 514936
rect 676047 514478 676113 514481
rect 676047 514476 676320 514478
rect 676047 514420 676052 514476
rect 676108 514420 676320 514476
rect 676047 514418 676320 514420
rect 676047 514415 676113 514418
rect 679983 514108 680049 514111
rect 679938 514106 680049 514108
rect 679938 514050 679988 514106
rect 680044 514050 680049 514106
rect 679938 514045 680049 514050
rect 679938 513930 679998 514045
rect 679746 513223 679806 513486
rect 679746 513218 679857 513223
rect 679983 513220 680049 513223
rect 679746 513162 679796 513218
rect 679852 513162 679857 513218
rect 679746 513160 679857 513162
rect 679791 513157 679857 513160
rect 679938 513218 680049 513220
rect 679938 513162 679988 513218
rect 680044 513162 680049 513218
rect 679938 513157 680049 513162
rect 679938 512968 679998 513157
rect 679791 512776 679857 512779
rect 679746 512774 679857 512776
rect 679746 512718 679796 512774
rect 679852 512718 679857 512774
rect 679746 512713 679857 512718
rect 679746 512450 679806 512713
rect 676290 482439 676350 482702
rect 676290 482434 676401 482439
rect 676290 482378 676340 482434
rect 676396 482378 676401 482434
rect 676290 482376 676401 482378
rect 676335 482373 676401 482376
rect 676143 481844 676209 481847
rect 676290 481844 676350 482110
rect 676143 481842 676350 481844
rect 676143 481786 676148 481842
rect 676204 481786 676350 481842
rect 676143 481784 676350 481786
rect 676143 481781 676209 481784
rect 676290 481403 676350 481592
rect 676239 481398 676350 481403
rect 676527 481400 676593 481403
rect 676239 481342 676244 481398
rect 676300 481342 676350 481398
rect 676239 481340 676350 481342
rect 676482 481398 676593 481400
rect 676482 481342 676532 481398
rect 676588 481342 676593 481398
rect 676239 481337 676305 481340
rect 676482 481337 676593 481342
rect 676482 481222 676542 481337
rect 676674 480367 676734 480630
rect 676431 480364 676497 480367
rect 676431 480362 676542 480364
rect 676431 480306 676436 480362
rect 676492 480306 676542 480362
rect 676431 480301 676542 480306
rect 676674 480362 676785 480367
rect 676674 480306 676724 480362
rect 676780 480306 676785 480362
rect 676674 480304 676785 480306
rect 676719 480301 676785 480304
rect 676482 480038 676542 480301
rect 676047 479698 676113 479701
rect 676047 479696 676320 479698
rect 676047 479640 676052 479696
rect 676108 479640 676320 479696
rect 676047 479638 676320 479640
rect 676047 479635 676113 479638
rect 676623 479328 676689 479331
rect 676623 479326 676734 479328
rect 676623 479270 676628 479326
rect 676684 479270 676734 479326
rect 676623 479265 676734 479270
rect 676674 479150 676734 479265
rect 676290 478443 676350 478558
rect 676239 478438 676350 478443
rect 676239 478382 676244 478438
rect 676300 478382 676350 478438
rect 676239 478380 676350 478382
rect 676239 478377 676305 478380
rect 675130 478230 675136 478294
rect 675200 478292 675206 478294
rect 675200 478232 676350 478292
rect 675200 478230 675206 478232
rect 676290 478188 676350 478232
rect 676282 477786 676288 477850
rect 676352 477786 676358 477850
rect 676290 477670 676350 477786
rect 674362 477046 674368 477110
rect 674432 477108 674438 477110
rect 674432 477048 676320 477108
rect 674432 477046 674438 477048
rect 674746 476602 674752 476666
rect 674816 476664 674822 476666
rect 674816 476604 676320 476664
rect 674816 476602 674822 476604
rect 675322 476158 675328 476222
rect 675392 476220 675398 476222
rect 675392 476160 676320 476220
rect 675392 476158 675398 476160
rect 41775 476072 41841 476075
rect 41568 476070 41841 476072
rect 41568 476014 41780 476070
rect 41836 476014 41841 476070
rect 41568 476012 41841 476014
rect 41775 476009 41841 476012
rect 676047 475628 676113 475631
rect 676047 475626 676320 475628
rect 676047 475570 676052 475626
rect 676108 475570 676320 475626
rect 676047 475568 676320 475570
rect 676047 475565 676113 475568
rect 41775 475554 41841 475557
rect 41568 475552 41841 475554
rect 41568 475496 41780 475552
rect 41836 475496 41841 475552
rect 41568 475494 41841 475496
rect 41775 475491 41841 475494
rect 673978 475122 673984 475186
rect 674048 475184 674054 475186
rect 674048 475124 676320 475184
rect 674048 475122 674054 475124
rect 41775 475036 41841 475039
rect 41568 475034 41841 475036
rect 41568 474978 41780 475034
rect 41836 474978 41841 475034
rect 41568 474976 41841 474978
rect 41775 474973 41841 474976
rect 676047 474666 676113 474669
rect 676047 474664 676320 474666
rect 676047 474608 676052 474664
rect 676108 474608 676320 474664
rect 676047 474606 676320 474608
rect 676047 474603 676113 474606
rect 41871 474592 41937 474595
rect 41568 474590 41937 474592
rect 41568 474534 41876 474590
rect 41932 474534 41937 474590
rect 41568 474532 41937 474534
rect 41871 474529 41937 474532
rect 676239 474296 676305 474299
rect 676239 474294 676350 474296
rect 676239 474238 676244 474294
rect 676300 474238 676350 474294
rect 676239 474233 676350 474238
rect 676290 474118 676350 474233
rect 40386 473855 40446 473970
rect 40335 473850 40446 473855
rect 40335 473794 40340 473850
rect 40396 473794 40446 473850
rect 40335 473792 40446 473794
rect 40335 473789 40401 473792
rect 677058 473558 677118 473674
rect 41538 473260 41598 473526
rect 676858 473494 676864 473558
rect 676928 473494 676934 473558
rect 677050 473494 677056 473558
rect 677120 473494 677126 473558
rect 41679 473260 41745 473263
rect 41538 473258 41745 473260
rect 41538 473202 41684 473258
rect 41740 473202 41745 473258
rect 41538 473200 41745 473202
rect 41679 473197 41745 473200
rect 676866 473156 676926 473494
rect 43311 473112 43377 473115
rect 45039 473112 45105 473115
rect 41568 473110 45105 473112
rect 41568 473054 43316 473110
rect 43372 473054 45044 473110
rect 45100 473054 45105 473110
rect 41568 473052 45105 473054
rect 43311 473049 43377 473052
rect 45039 473049 45105 473052
rect 676239 472816 676305 472819
rect 676239 472814 676350 472816
rect 676239 472758 676244 472814
rect 676300 472758 676350 472814
rect 676239 472753 676350 472758
rect 676290 472638 676350 472753
rect 39618 472375 39678 472490
rect 39618 472370 39729 472375
rect 39618 472314 39668 472370
rect 39724 472314 39729 472370
rect 39618 472312 39729 472314
rect 39663 472309 39729 472312
rect 676047 472224 676113 472227
rect 676047 472222 676320 472224
rect 676047 472166 676052 472222
rect 676108 472166 676320 472222
rect 676047 472164 676320 472166
rect 676047 472161 676113 472164
rect 41775 472076 41841 472079
rect 41568 472074 41841 472076
rect 41568 472018 41780 472074
rect 41836 472018 41841 472074
rect 41568 472016 41841 472018
rect 41775 472013 41841 472016
rect 42490 471632 42496 471634
rect 41568 471572 42496 471632
rect 42490 471570 42496 471572
rect 42560 471570 42566 471634
rect 676047 471632 676113 471635
rect 676047 471630 676320 471632
rect 676047 471574 676052 471630
rect 676108 471574 676320 471630
rect 676047 471572 676320 471574
rect 676047 471569 676113 471572
rect 40570 471274 40576 471338
rect 40640 471274 40646 471338
rect 40578 471010 40638 471274
rect 679746 470895 679806 471158
rect 42682 470892 42688 470894
rect 41538 470832 42688 470892
rect 41538 470492 41598 470832
rect 42682 470830 42688 470832
rect 42752 470830 42758 470894
rect 679746 470890 679857 470895
rect 679746 470834 679796 470890
rect 679852 470834 679857 470890
rect 679746 470832 679857 470834
rect 679791 470829 679857 470832
rect 685506 470451 685566 470714
rect 679791 470448 679857 470451
rect 679746 470446 679857 470448
rect 679746 470390 679796 470446
rect 679852 470390 679857 470446
rect 679746 470385 679857 470390
rect 685455 470446 685566 470451
rect 685455 470390 685460 470446
rect 685516 470390 685566 470446
rect 685455 470388 685566 470390
rect 685455 470385 685521 470388
rect 42298 470152 42304 470154
rect 41568 470092 42304 470152
rect 42298 470090 42304 470092
rect 42368 470090 42374 470154
rect 679746 470122 679806 470385
rect 685455 470004 685521 470007
rect 685455 470002 685566 470004
rect 685455 469946 685460 470002
rect 685516 469946 685566 470002
rect 685455 469941 685566 469946
rect 685506 469604 685566 469941
rect 41914 469560 41920 469562
rect 41568 469500 41920 469560
rect 41914 469498 41920 469500
rect 41984 469498 41990 469562
rect 40378 469350 40384 469414
rect 40448 469350 40454 469414
rect 40386 468938 40446 469350
rect 42106 468672 42112 468674
rect 41568 468612 42112 468672
rect 42106 468610 42112 468612
rect 42176 468610 42182 468674
rect 41722 468080 41728 468082
rect 41568 468020 41728 468080
rect 41722 468018 41728 468020
rect 41792 468018 41798 468082
rect 41530 467722 41536 467786
rect 41600 467722 41606 467786
rect 41538 467458 41598 467722
rect 40954 467278 40960 467342
rect 41024 467278 41030 467342
rect 40962 467088 41022 467278
rect 41338 466834 41344 466898
rect 41408 466834 41414 466898
rect 41346 466570 41406 466834
rect 41146 466242 41152 466306
rect 41216 466242 41222 466306
rect 41154 465978 41214 466242
rect 40762 465798 40768 465862
rect 40832 465798 40838 465862
rect 40770 465608 40830 465798
rect 41583 465268 41649 465271
rect 41538 465266 41649 465268
rect 41538 465210 41588 465266
rect 41644 465210 41649 465266
rect 41538 465205 41649 465210
rect 41538 465090 41598 465205
rect 34434 464383 34494 464498
rect 34434 464378 34545 464383
rect 34434 464322 34484 464378
rect 34540 464322 34545 464378
rect 34434 464320 34545 464322
rect 34479 464317 34545 464320
rect 23106 463791 23166 464054
rect 23055 463786 23166 463791
rect 23055 463730 23060 463786
rect 23116 463730 23166 463786
rect 23055 463728 23166 463730
rect 23055 463725 23121 463728
rect 41775 463640 41841 463643
rect 41568 463638 41841 463640
rect 41568 463582 41780 463638
rect 41836 463582 41841 463638
rect 41568 463580 41841 463582
rect 41775 463577 41841 463580
rect 23055 463344 23121 463347
rect 23055 463342 23166 463344
rect 23055 463286 23060 463342
rect 23116 463286 23166 463342
rect 23055 463281 23166 463286
rect 23106 463018 23166 463281
rect 41775 429304 41841 429307
rect 41568 429302 41841 429304
rect 41568 429246 41780 429302
rect 41836 429246 41841 429302
rect 41568 429244 41841 429246
rect 41775 429241 41841 429244
rect 41538 428567 41598 428682
rect 41538 428562 41649 428567
rect 41538 428506 41588 428562
rect 41644 428506 41649 428562
rect 41538 428504 41649 428506
rect 41583 428501 41649 428504
rect 41775 428268 41841 428271
rect 41568 428266 41841 428268
rect 41568 428210 41780 428266
rect 41836 428210 41841 428266
rect 41568 428208 41841 428210
rect 41775 428205 41841 428208
rect 40335 427972 40401 427975
rect 40335 427970 40446 427972
rect 40335 427914 40340 427970
rect 40396 427914 40446 427970
rect 40335 427909 40446 427914
rect 40386 427794 40446 427909
rect 41538 427087 41598 427202
rect 41538 427082 41649 427087
rect 41538 427026 41588 427082
rect 41644 427026 41649 427082
rect 41538 427024 41649 427026
rect 41583 427021 41649 427024
rect 41775 426714 41841 426717
rect 41568 426712 41841 426714
rect 41568 426656 41780 426712
rect 41836 426656 41841 426712
rect 41568 426654 41841 426656
rect 41775 426651 41841 426654
rect 41679 426492 41745 426495
rect 41538 426490 41745 426492
rect 41538 426434 41684 426490
rect 41740 426434 41745 426490
rect 41538 426432 41745 426434
rect 41538 426314 41598 426432
rect 41679 426429 41745 426432
rect 41538 425607 41598 425722
rect 41538 425602 41649 425607
rect 41538 425546 41588 425602
rect 41644 425546 41649 425602
rect 41538 425544 41649 425546
rect 41583 425541 41649 425544
rect 41538 425012 41598 425130
rect 41679 425012 41745 425015
rect 41538 425010 41745 425012
rect 41538 424954 41684 425010
rect 41740 424954 41745 425010
rect 41538 424952 41745 424954
rect 41679 424949 41745 424952
rect 41538 424422 41598 424834
rect 41530 424358 41536 424422
rect 41600 424358 41606 424422
rect 41914 424272 41920 424274
rect 41568 424212 41920 424272
rect 41914 424210 41920 424212
rect 41984 424210 41990 424274
rect 42106 423680 42112 423682
rect 41568 423620 42112 423680
rect 42106 423618 42112 423620
rect 42176 423618 42182 423682
rect 41154 422942 41214 423280
rect 41146 422878 41152 422942
rect 41216 422878 41222 422942
rect 42682 422792 42688 422794
rect 41568 422732 42688 422792
rect 42682 422730 42688 422732
rect 42752 422730 42758 422794
rect 41775 422200 41841 422203
rect 41568 422198 41841 422200
rect 41568 422142 41780 422198
rect 41836 422142 41841 422198
rect 41568 422140 41841 422142
rect 41775 422137 41841 422140
rect 40770 421462 40830 421800
rect 40762 421398 40768 421462
rect 40832 421398 40838 421462
rect 40962 421018 41022 421282
rect 40954 420954 40960 421018
rect 41024 420954 41030 421018
rect 41346 420574 41406 420690
rect 41338 420510 41344 420574
rect 41408 420510 41414 420574
rect 41538 420131 41598 420246
rect 41538 420126 41649 420131
rect 41538 420070 41588 420126
rect 41644 420070 41649 420126
rect 41538 420068 41649 420070
rect 41583 420065 41649 420068
rect 41722 419832 41728 419834
rect 41568 419772 41728 419832
rect 41722 419770 41728 419772
rect 41792 419770 41798 419834
rect 40378 419326 40384 419390
rect 40448 419326 40454 419390
rect 40386 419210 40446 419326
rect 42490 418796 42496 418798
rect 41568 418736 42496 418796
rect 42490 418734 42496 418736
rect 42560 418734 42566 418798
rect 40578 417910 40638 418248
rect 40570 417846 40576 417910
rect 40640 417846 40646 417910
rect 41568 417700 41790 417760
rect 28866 417023 28926 417286
rect 41730 417168 41790 417700
rect 41538 417108 41790 417168
rect 28866 417018 28977 417023
rect 28866 416962 28916 417018
rect 28972 416962 28977 417018
rect 28866 416960 28977 416962
rect 28911 416957 28977 416960
rect 41538 416579 41598 417108
rect 28911 416576 28977 416579
rect 28866 416574 28977 416576
rect 28866 416518 28916 416574
rect 28972 416518 28977 416574
rect 28866 416513 28977 416518
rect 41538 416574 41649 416579
rect 41538 416518 41588 416574
rect 41644 416518 41649 416574
rect 41538 416516 41649 416518
rect 41583 416513 41649 416516
rect 28866 416250 28926 416513
rect 41871 411694 41937 411695
rect 41871 411690 41920 411694
rect 41984 411692 41990 411694
rect 41871 411634 41876 411690
rect 41871 411630 41920 411634
rect 41984 411632 42028 411692
rect 41984 411630 41990 411632
rect 41871 411629 41937 411630
rect 41722 411482 41728 411546
rect 41792 411482 41798 411546
rect 41730 411102 41790 411482
rect 41722 411038 41728 411102
rect 41792 411038 41798 411102
rect 40570 408374 40576 408438
rect 40640 408436 40646 408438
rect 41775 408436 41841 408439
rect 40640 408434 41841 408436
rect 40640 408378 41780 408434
rect 41836 408378 41841 408434
rect 40640 408376 41841 408378
rect 40640 408374 40646 408376
rect 41775 408373 41841 408376
rect 41775 407994 41841 407995
rect 41722 407992 41728 407994
rect 41684 407932 41728 407992
rect 41792 407990 41841 407994
rect 41836 407934 41841 407990
rect 41722 407930 41728 407932
rect 41792 407930 41841 407934
rect 41775 407929 41841 407930
rect 42159 407400 42225 407403
rect 42490 407400 42496 407402
rect 42159 407398 42496 407400
rect 42159 407342 42164 407398
rect 42220 407342 42496 407398
rect 42159 407340 42496 407342
rect 42159 407337 42225 407340
rect 42490 407338 42496 407340
rect 42560 407338 42566 407402
rect 42063 406512 42129 406515
rect 42682 406512 42688 406514
rect 42063 406510 42688 406512
rect 42063 406454 42068 406510
rect 42124 406454 42688 406510
rect 42063 406452 42688 406454
rect 42063 406449 42129 406452
rect 42682 406450 42688 406452
rect 42752 406450 42758 406514
rect 40378 404230 40384 404294
rect 40448 404292 40454 404294
rect 41775 404292 41841 404295
rect 40448 404290 41841 404292
rect 40448 404234 41780 404290
rect 41836 404234 41841 404290
rect 40448 404232 41841 404234
rect 40448 404230 40454 404232
rect 41775 404229 41841 404232
rect 58479 404144 58545 404147
rect 58479 404142 64638 404144
rect 58479 404086 58484 404142
rect 58540 404086 64638 404142
rect 58479 404084 64638 404086
rect 58479 404081 58545 404084
rect 41338 403638 41344 403702
rect 41408 403700 41414 403702
rect 41775 403700 41841 403703
rect 41408 403698 41841 403700
rect 41408 403642 41780 403698
rect 41836 403642 41841 403698
rect 41408 403640 41841 403642
rect 41408 403638 41414 403640
rect 41775 403637 41841 403640
rect 64578 403550 64638 404084
rect 40954 402898 40960 402962
rect 41024 402960 41030 402962
rect 41775 402960 41841 402963
rect 41024 402958 41841 402960
rect 41024 402902 41780 402958
rect 41836 402902 41841 402958
rect 41024 402900 41841 402902
rect 41024 402898 41030 402900
rect 41775 402897 41841 402900
rect 59631 402812 59697 402815
rect 59631 402810 64638 402812
rect 59631 402754 59636 402810
rect 59692 402754 64638 402810
rect 59631 402752 64638 402754
rect 59631 402749 59697 402752
rect 41146 402306 41152 402370
rect 41216 402368 41222 402370
rect 41775 402368 41841 402371
rect 64578 402368 64638 402752
rect 41216 402366 41841 402368
rect 41216 402310 41780 402366
rect 41836 402310 41841 402366
rect 41216 402308 41841 402310
rect 41216 402306 41222 402308
rect 41775 402305 41841 402308
rect 57615 400592 57681 400595
rect 64578 400592 64638 401186
rect 57615 400590 64638 400592
rect 57615 400534 57620 400590
rect 57676 400534 64638 400590
rect 57615 400532 64638 400534
rect 57615 400529 57681 400532
rect 41871 400298 41937 400299
rect 41871 400294 41920 400298
rect 41984 400296 41990 400298
rect 41871 400238 41876 400294
rect 41871 400234 41920 400238
rect 41984 400236 42028 400296
rect 41984 400234 41990 400236
rect 41871 400233 41937 400234
rect 59631 400000 59697 400003
rect 64578 400000 64638 400004
rect 59631 399998 64638 400000
rect 59631 399942 59636 399998
rect 59692 399942 64638 399998
rect 59631 399940 64638 399942
rect 59631 399937 59697 399940
rect 40762 399790 40768 399854
rect 40832 399852 40838 399854
rect 41775 399852 41841 399855
rect 40832 399850 41841 399852
rect 40832 399794 41780 399850
rect 41836 399794 41841 399850
rect 40832 399792 41841 399794
rect 40832 399790 40838 399792
rect 41775 399789 41841 399792
rect 42159 399410 42225 399411
rect 42106 399408 42112 399410
rect 42068 399348 42112 399408
rect 42176 399406 42225 399410
rect 42220 399350 42225 399406
rect 42106 399346 42112 399348
rect 42176 399346 42225 399350
rect 42159 399345 42225 399346
rect 59727 399408 59793 399411
rect 59727 399406 64638 399408
rect 59727 399350 59732 399406
rect 59788 399350 64638 399406
rect 59727 399348 64638 399350
rect 59727 399345 59793 399348
rect 64578 398822 64638 399348
rect 59535 398224 59601 398227
rect 59535 398222 64638 398224
rect 59535 398166 59540 398222
rect 59596 398166 64638 398222
rect 59535 398164 64638 398166
rect 59535 398161 59601 398164
rect 64578 397640 64638 398164
rect 676143 396448 676209 396451
rect 676290 396448 676350 396714
rect 676143 396446 676350 396448
rect 676143 396390 676148 396446
rect 676204 396390 676350 396446
rect 676143 396388 676350 396390
rect 676143 396385 676209 396388
rect 676290 395859 676350 396122
rect 676290 395854 676401 395859
rect 676290 395798 676340 395854
rect 676396 395798 676401 395854
rect 676290 395796 676401 395798
rect 676335 395793 676401 395796
rect 676290 395415 676350 395530
rect 676239 395410 676350 395415
rect 676719 395412 676785 395415
rect 676239 395354 676244 395410
rect 676300 395354 676350 395410
rect 676239 395352 676350 395354
rect 676674 395410 676785 395412
rect 676674 395354 676724 395410
rect 676780 395354 676785 395410
rect 676239 395349 676305 395352
rect 676674 395349 676785 395354
rect 676674 395160 676734 395349
rect 673978 394610 673984 394674
rect 674048 394672 674054 394674
rect 674048 394612 676320 394672
rect 674048 394610 674054 394612
rect 676290 393935 676350 394050
rect 676239 393930 676350 393935
rect 676239 393874 676244 393930
rect 676300 393874 676350 393930
rect 676239 393872 676350 393874
rect 676239 393869 676305 393872
rect 674362 393278 674368 393342
rect 674432 393340 674438 393342
rect 676290 393340 676350 393680
rect 674432 393280 676350 393340
rect 674432 393278 674438 393280
rect 675855 393192 675921 393195
rect 675855 393190 676320 393192
rect 675855 393134 675860 393190
rect 675916 393134 676320 393190
rect 675855 393132 676320 393134
rect 675855 393129 675921 393132
rect 674170 392538 674176 392602
rect 674240 392600 674246 392602
rect 674240 392540 676320 392600
rect 674240 392538 674246 392540
rect 676290 392011 676350 392126
rect 676239 392006 676350 392011
rect 676239 391950 676244 392006
rect 676300 391950 676350 392006
rect 676239 391948 676350 391950
rect 676239 391945 676305 391948
rect 674554 391650 674560 391714
rect 674624 391712 674630 391714
rect 674624 391652 676320 391712
rect 674624 391650 674630 391652
rect 675567 391120 675633 391123
rect 675567 391118 676320 391120
rect 675567 391062 675572 391118
rect 675628 391062 676320 391118
rect 675567 391060 676320 391062
rect 675567 391057 675633 391060
rect 676290 390531 676350 390646
rect 676239 390526 676350 390531
rect 676239 390470 676244 390526
rect 676300 390470 676350 390526
rect 676239 390468 676350 390470
rect 676239 390465 676305 390468
rect 676047 390158 676113 390161
rect 676047 390156 676320 390158
rect 676047 390100 676052 390156
rect 676108 390100 676320 390156
rect 676047 390098 676320 390100
rect 676047 390095 676113 390098
rect 676047 389640 676113 389643
rect 676047 389638 676320 389640
rect 676047 389582 676052 389638
rect 676108 389582 676320 389638
rect 676047 389580 676320 389582
rect 676047 389577 676113 389580
rect 676290 389051 676350 389166
rect 676239 389046 676350 389051
rect 676239 388990 676244 389046
rect 676300 388990 676350 389046
rect 676239 388988 676350 388990
rect 676239 388985 676305 388988
rect 676047 388678 676113 388681
rect 676047 388676 676320 388678
rect 676047 388620 676052 388676
rect 676108 388620 676320 388676
rect 676047 388618 676320 388620
rect 676047 388615 676113 388618
rect 675951 388160 676017 388163
rect 675951 388158 676320 388160
rect 675951 388102 675956 388158
rect 676012 388102 676320 388158
rect 675951 388100 676320 388102
rect 675951 388097 676017 388100
rect 676290 387571 676350 387686
rect 676239 387566 676350 387571
rect 676239 387510 676244 387566
rect 676300 387510 676350 387566
rect 676239 387508 676350 387510
rect 676239 387505 676305 387508
rect 676290 386979 676350 387094
rect 676239 386974 676350 386979
rect 676239 386918 676244 386974
rect 676300 386918 676350 386974
rect 676239 386916 676350 386918
rect 676239 386913 676305 386916
rect 676047 386680 676113 386683
rect 676047 386678 676320 386680
rect 676047 386622 676052 386678
rect 676108 386622 676320 386678
rect 676047 386620 676320 386622
rect 676047 386617 676113 386620
rect 675951 386236 676017 386239
rect 675951 386234 676320 386236
rect 675951 386178 675956 386234
rect 676012 386178 676320 386234
rect 675951 386176 676320 386178
rect 675951 386173 676017 386176
rect 41775 386088 41841 386091
rect 41568 386086 41841 386088
rect 41568 386030 41780 386086
rect 41836 386030 41841 386086
rect 41568 386028 41841 386030
rect 41775 386025 41841 386028
rect 676290 385499 676350 385614
rect 676239 385494 676350 385499
rect 41538 385351 41598 385466
rect 676239 385438 676244 385494
rect 676300 385438 676350 385494
rect 676239 385436 676350 385438
rect 676239 385433 676305 385436
rect 41538 385346 41649 385351
rect 41538 385290 41588 385346
rect 41644 385290 41649 385346
rect 41538 385288 41649 385290
rect 41583 385285 41649 385288
rect 41775 385052 41841 385055
rect 41568 385050 41841 385052
rect 41568 384994 41780 385050
rect 41836 384994 41841 385050
rect 41568 384992 41841 384994
rect 41775 384989 41841 384992
rect 679746 384907 679806 385096
rect 679695 384902 679806 384907
rect 679695 384846 679700 384902
rect 679756 384846 679806 384902
rect 679695 384844 679806 384846
rect 679695 384841 679761 384844
rect 41583 384756 41649 384759
rect 41538 384754 41649 384756
rect 41538 384698 41588 384754
rect 41644 384698 41649 384754
rect 41538 384693 41649 384698
rect 41538 384578 41598 384693
rect 685506 384463 685566 384726
rect 679695 384460 679761 384463
rect 679695 384458 679806 384460
rect 679695 384402 679700 384458
rect 679756 384402 679806 384458
rect 679695 384397 679806 384402
rect 685455 384458 685566 384463
rect 685455 384402 685460 384458
rect 685516 384402 685566 384458
rect 685455 384400 685566 384402
rect 685455 384397 685521 384400
rect 679746 384134 679806 384397
rect 685455 384016 685521 384019
rect 685455 384014 685566 384016
rect 41538 383871 41598 383986
rect 685455 383958 685460 384014
rect 685516 383958 685566 384014
rect 685455 383953 685566 383958
rect 41538 383866 41649 383871
rect 41538 383810 41588 383866
rect 41644 383810 41649 383866
rect 41538 383808 41649 383810
rect 41583 383805 41649 383808
rect 685506 383616 685566 383953
rect 41775 383572 41841 383575
rect 41568 383570 41841 383572
rect 41568 383514 41780 383570
rect 41836 383514 41841 383570
rect 41568 383512 41841 383514
rect 41775 383509 41841 383512
rect 41583 383276 41649 383279
rect 41538 383274 41649 383276
rect 41538 383218 41588 383274
rect 41644 383218 41649 383274
rect 41538 383213 41649 383218
rect 41538 383098 41598 383213
rect 40002 382243 40062 382506
rect 39951 382238 40062 382243
rect 39951 382182 39956 382238
rect 40012 382182 40062 382238
rect 39951 382180 40062 382182
rect 39951 382177 40017 382180
rect 41775 382018 41841 382021
rect 41568 382016 41841 382018
rect 41568 381960 41780 382016
rect 41836 381960 41841 382016
rect 41568 381958 41841 381960
rect 41775 381955 41841 381958
rect 40386 381354 40446 381618
rect 40378 381290 40384 381354
rect 40448 381290 40454 381354
rect 42106 381056 42112 381058
rect 41568 380996 42112 381056
rect 42106 380994 42112 380996
rect 42176 380994 42182 381058
rect 42682 380464 42688 380466
rect 41568 380404 42688 380464
rect 42682 380402 42688 380404
rect 42752 380402 42758 380466
rect 40962 379726 41022 380138
rect 40954 379662 40960 379726
rect 41024 379662 41030 379726
rect 42298 379576 42304 379578
rect 41568 379516 42304 379576
rect 42298 379514 42304 379516
rect 42368 379514 42374 379578
rect 41775 378984 41841 378987
rect 41568 378982 41841 378984
rect 41568 378926 41780 378982
rect 41836 378926 41841 378982
rect 41568 378924 41841 378926
rect 41775 378921 41841 378924
rect 40770 378246 40830 378584
rect 40762 378182 40768 378246
rect 40832 378182 40838 378246
rect 41154 377802 41214 378066
rect 41146 377738 41152 377802
rect 41216 377738 41222 377802
rect 41346 377312 41406 377474
rect 41338 377248 41344 377312
rect 41408 377248 41414 377312
rect 41538 376915 41598 377104
rect 41538 376910 41649 376915
rect 41538 376854 41588 376910
rect 41644 376854 41649 376910
rect 41538 376852 41649 376854
rect 41583 376849 41649 376852
rect 40954 376702 40960 376766
rect 41024 376764 41030 376766
rect 42490 376764 42496 376766
rect 41024 376704 42496 376764
rect 41024 376702 41030 376704
rect 42490 376702 42496 376704
rect 42560 376702 42566 376766
rect 41914 376616 41920 376618
rect 41568 376556 41920 376616
rect 41914 376554 41920 376556
rect 41984 376554 41990 376618
rect 40578 375878 40638 375994
rect 40570 375814 40576 375878
rect 40640 375814 40646 375878
rect 41538 375286 41598 375550
rect 41530 375222 41536 375286
rect 41600 375222 41606 375286
rect 41722 375136 41728 375138
rect 41568 375076 41728 375136
rect 41722 375074 41728 375076
rect 41792 375074 41798 375138
rect 41568 374484 41790 374544
rect 28866 373807 28926 374070
rect 41730 373952 41790 374484
rect 655119 374396 655185 374399
rect 28815 373802 28926 373807
rect 28815 373746 28820 373802
rect 28876 373746 28926 373802
rect 28815 373744 28926 373746
rect 41538 373892 41790 373952
rect 649986 374394 655185 374396
rect 649986 374338 655124 374394
rect 655180 374338 655185 374394
rect 649986 374336 655185 374338
rect 649986 373892 650046 374336
rect 655119 374333 655185 374336
rect 28815 373741 28881 373744
rect 41538 373363 41598 373892
rect 28815 373360 28881 373363
rect 28815 373358 28926 373360
rect 28815 373302 28820 373358
rect 28876 373302 28926 373358
rect 28815 373297 28926 373302
rect 41538 373358 41649 373363
rect 655503 373360 655569 373363
rect 41538 373302 41588 373358
rect 41644 373302 41649 373358
rect 41538 373300 41649 373302
rect 41583 373297 41649 373300
rect 649986 373358 655569 373360
rect 649986 373302 655508 373358
rect 655564 373302 655569 373358
rect 649986 373300 655569 373302
rect 28866 373034 28926 373297
rect 649986 372710 650046 373300
rect 655503 373297 655569 373300
rect 655311 372176 655377 372179
rect 649986 372174 655377 372176
rect 649986 372118 655316 372174
rect 655372 372118 655377 372174
rect 649986 372116 655377 372118
rect 649986 371528 650046 372116
rect 655311 372113 655377 372116
rect 654159 370992 654225 370995
rect 649986 370990 654225 370992
rect 649986 370934 654164 370990
rect 654220 370934 654225 370990
rect 649986 370932 654225 370934
rect 649986 370346 650046 370932
rect 654159 370929 654225 370932
rect 42063 368478 42129 368479
rect 42063 368474 42112 368478
rect 42176 368476 42182 368478
rect 42063 368418 42068 368474
rect 42063 368414 42112 368418
rect 42176 368416 42220 368476
rect 42176 368414 42182 368416
rect 42063 368413 42129 368414
rect 674554 367230 674560 367294
rect 674624 367292 674630 367294
rect 675471 367292 675537 367295
rect 674624 367290 675537 367292
rect 674624 367234 675476 367290
rect 675532 367234 675537 367290
rect 674624 367232 675537 367234
rect 674624 367230 674630 367232
rect 675471 367229 675537 367232
rect 41775 365222 41841 365223
rect 41722 365220 41728 365222
rect 41684 365160 41728 365220
rect 41792 365218 41841 365222
rect 41836 365162 41841 365218
rect 41722 365158 41728 365160
rect 41792 365158 41841 365162
rect 41775 365157 41841 365158
rect 41967 364630 42033 364631
rect 41914 364628 41920 364630
rect 41876 364568 41920 364628
rect 41984 364626 42033 364630
rect 42028 364570 42033 364626
rect 41914 364566 41920 364568
rect 41984 364566 42033 364570
rect 41967 364565 42033 364566
rect 41530 364122 41536 364186
rect 41600 364184 41606 364186
rect 41775 364184 41841 364187
rect 41600 364182 41841 364184
rect 41600 364126 41780 364182
rect 41836 364126 41841 364182
rect 41600 364124 41841 364126
rect 41600 364122 41606 364124
rect 41775 364121 41841 364124
rect 42159 363592 42225 363595
rect 42298 363592 42304 363594
rect 42159 363590 42304 363592
rect 42159 363534 42164 363590
rect 42220 363534 42304 363590
rect 42159 363532 42304 363534
rect 42159 363529 42225 363532
rect 42298 363530 42304 363532
rect 42368 363530 42374 363594
rect 40570 361014 40576 361078
rect 40640 361076 40646 361078
rect 41775 361076 41841 361079
rect 40640 361074 41841 361076
rect 40640 361018 41780 361074
rect 41836 361018 41841 361074
rect 40640 361016 41841 361018
rect 40640 361014 40646 361016
rect 41775 361013 41841 361016
rect 58287 360928 58353 360931
rect 58287 360926 64638 360928
rect 58287 360870 58292 360926
rect 58348 360870 64638 360926
rect 58287 360868 64638 360870
rect 58287 360865 58353 360868
rect 41338 360422 41344 360486
rect 41408 360484 41414 360486
rect 41775 360484 41841 360487
rect 41408 360482 41841 360484
rect 41408 360426 41780 360482
rect 41836 360426 41841 360482
rect 41408 360424 41841 360426
rect 41408 360422 41414 360424
rect 41775 360421 41841 360424
rect 64578 360328 64638 360868
rect 40954 359682 40960 359746
rect 41024 359744 41030 359746
rect 41775 359744 41841 359747
rect 41024 359742 41841 359744
rect 41024 359686 41780 359742
rect 41836 359686 41841 359742
rect 41024 359684 41841 359686
rect 41024 359682 41030 359684
rect 41775 359681 41841 359684
rect 59151 359744 59217 359747
rect 59151 359742 64638 359744
rect 59151 359686 59156 359742
rect 59212 359686 64638 359742
rect 59151 359684 64638 359686
rect 59151 359681 59217 359684
rect 64578 359146 64638 359684
rect 42063 359004 42129 359007
rect 42490 359004 42496 359006
rect 42063 359002 42496 359004
rect 42063 358946 42068 359002
rect 42124 358946 42496 359002
rect 42063 358944 42496 358946
rect 42063 358941 42129 358944
rect 42490 358942 42496 358944
rect 42560 358942 42566 359006
rect 57615 357524 57681 357527
rect 64578 357524 64638 357964
rect 57615 357522 64638 357524
rect 57615 357466 57620 357522
rect 57676 357466 64638 357522
rect 57615 357464 64638 357466
rect 57615 357461 57681 357464
rect 40378 357166 40384 357230
rect 40448 357228 40454 357230
rect 41775 357228 41841 357231
rect 40448 357226 41841 357228
rect 40448 357170 41780 357226
rect 41836 357170 41841 357226
rect 40448 357168 41841 357170
rect 40448 357166 40454 357168
rect 41775 357165 41841 357168
rect 59631 356784 59697 356787
rect 59631 356782 64638 356784
rect 59631 356726 59636 356782
rect 59692 356726 64638 356782
rect 59631 356724 64638 356726
rect 59631 356721 59697 356724
rect 40762 356574 40768 356638
rect 40832 356636 40838 356638
rect 41775 356636 41841 356639
rect 40832 356634 41841 356636
rect 40832 356578 41780 356634
rect 41836 356578 41841 356634
rect 40832 356576 41841 356578
rect 40832 356574 40838 356576
rect 41775 356573 41841 356576
rect 42159 356192 42225 356195
rect 42682 356192 42688 356194
rect 42159 356190 42688 356192
rect 42159 356134 42164 356190
rect 42220 356134 42688 356190
rect 42159 356132 42688 356134
rect 42159 356129 42225 356132
rect 42682 356130 42688 356132
rect 42752 356130 42758 356194
rect 58191 356192 58257 356195
rect 58191 356190 64638 356192
rect 58191 356134 58196 356190
rect 58252 356134 64638 356190
rect 58191 356132 64638 356134
rect 58191 356129 58257 356132
rect 64578 355600 64638 356132
rect 58575 355008 58641 355011
rect 58575 355006 64638 355008
rect 58575 354950 58580 355006
rect 58636 354950 64638 355006
rect 58575 354948 64638 354950
rect 58575 354945 58641 354948
rect 64578 354418 64638 354948
rect 676290 351755 676350 352018
rect 676239 351750 676350 351755
rect 676239 351694 676244 351750
rect 676300 351694 676350 351750
rect 676239 351692 676350 351694
rect 676239 351689 676305 351692
rect 676047 351604 676113 351607
rect 676047 351602 676320 351604
rect 676047 351546 676052 351602
rect 676108 351546 676320 351602
rect 676047 351544 676320 351546
rect 676047 351541 676113 351544
rect 676047 351012 676113 351015
rect 676047 351010 676320 351012
rect 676047 350954 676052 351010
rect 676108 350954 676320 351010
rect 676047 350952 676320 350954
rect 676047 350949 676113 350952
rect 673978 350506 673984 350570
rect 674048 350568 674054 350570
rect 674048 350508 676320 350568
rect 674048 350506 674054 350508
rect 674554 349618 674560 349682
rect 674624 349680 674630 349682
rect 676290 349680 676350 350020
rect 674624 349620 676350 349680
rect 674624 349618 674630 349620
rect 674362 349470 674368 349534
rect 674432 349532 674438 349534
rect 675514 349532 675520 349534
rect 674432 349472 675520 349532
rect 674432 349470 674438 349472
rect 675514 349470 675520 349472
rect 675584 349532 675590 349534
rect 675584 349472 676320 349532
rect 675584 349470 675590 349472
rect 675322 349026 675328 349090
rect 675392 349088 675398 349090
rect 675392 349028 676320 349088
rect 675392 349026 675398 349028
rect 670479 348644 670545 348647
rect 674170 348644 674176 348646
rect 670479 348642 674176 348644
rect 670479 348586 670484 348642
rect 670540 348586 674176 348642
rect 670479 348584 674176 348586
rect 670479 348581 670545 348584
rect 674170 348582 674176 348584
rect 674240 348644 674246 348646
rect 674240 348584 676350 348644
rect 674240 348582 674246 348584
rect 676290 348540 676350 348584
rect 674362 347990 674368 348054
rect 674432 348052 674438 348054
rect 674432 347992 676320 348052
rect 674432 347990 674438 347992
rect 675130 347546 675136 347610
rect 675200 347608 675206 347610
rect 675200 347548 676320 347608
rect 675200 347546 675206 347548
rect 677058 346871 677118 346986
rect 677007 346866 677118 346871
rect 677007 346810 677012 346866
rect 677068 346810 677118 346866
rect 677007 346808 677118 346810
rect 677007 346805 677073 346808
rect 676047 346572 676113 346575
rect 676047 346570 676320 346572
rect 676047 346514 676052 346570
rect 676108 346514 676320 346570
rect 676047 346512 676320 346514
rect 676047 346509 676113 346512
rect 673978 346066 673984 346130
rect 674048 346128 674054 346130
rect 674048 346068 676320 346128
rect 674048 346066 674054 346068
rect 674746 345474 674752 345538
rect 674816 345536 674822 345538
rect 674816 345476 676320 345536
rect 674816 345474 674822 345476
rect 676866 344799 676926 344988
rect 676866 344794 676977 344799
rect 676866 344738 676916 344794
rect 676972 344738 676977 344794
rect 676866 344736 676977 344738
rect 676911 344733 676977 344736
rect 676047 344648 676113 344651
rect 676047 344646 676320 344648
rect 676047 344590 676052 344646
rect 676108 344590 676320 344646
rect 676047 344588 676320 344590
rect 676047 344585 676113 344588
rect 676290 343911 676350 344026
rect 676239 343906 676350 343911
rect 676239 343850 676244 343906
rect 676300 343850 676350 343906
rect 676239 343848 676350 343850
rect 676239 343845 676305 343848
rect 674938 343254 674944 343318
rect 675008 343316 675014 343318
rect 676290 343316 676350 343508
rect 675008 343256 676350 343316
rect 675008 343254 675014 343256
rect 676866 342875 676926 343138
rect 41775 342872 41841 342875
rect 41568 342870 41841 342872
rect 41568 342814 41780 342870
rect 41836 342814 41841 342870
rect 41568 342812 41841 342814
rect 41775 342809 41841 342812
rect 676815 342870 676926 342875
rect 676815 342814 676820 342870
rect 676876 342814 676926 342870
rect 676815 342812 676926 342814
rect 676815 342809 676881 342812
rect 676047 342576 676113 342579
rect 676047 342574 676320 342576
rect 676047 342518 676052 342574
rect 676108 342518 676320 342574
rect 676047 342516 676320 342518
rect 676047 342513 676113 342516
rect 41775 342354 41841 342357
rect 41568 342352 41841 342354
rect 41568 342296 41780 342352
rect 41836 342296 41841 342352
rect 41568 342294 41841 342296
rect 41775 342291 41841 342294
rect 676290 341839 676350 341954
rect 41775 341836 41841 341839
rect 41568 341834 41841 341836
rect 41568 341778 41780 341834
rect 41836 341778 41841 341834
rect 41568 341776 41841 341778
rect 41775 341773 41841 341776
rect 676239 341834 676350 341839
rect 676239 341778 676244 341834
rect 676300 341778 676350 341834
rect 676239 341776 676350 341778
rect 676239 341773 676305 341776
rect 675951 341614 676017 341617
rect 675951 341612 676320 341614
rect 675951 341556 675956 341612
rect 676012 341556 676320 341612
rect 675951 341554 676320 341556
rect 675951 341551 676017 341554
rect 41775 341392 41841 341395
rect 41568 341390 41841 341392
rect 41568 341334 41780 341390
rect 41836 341334 41841 341390
rect 41568 341332 41841 341334
rect 41775 341329 41841 341332
rect 676047 341096 676113 341099
rect 676047 341094 676320 341096
rect 676047 341038 676052 341094
rect 676108 341038 676320 341094
rect 676047 341036 676320 341038
rect 676047 341033 676113 341036
rect 41538 340655 41598 340770
rect 41538 340650 41649 340655
rect 41538 340594 41588 340650
rect 41644 340594 41649 340650
rect 41538 340592 41649 340594
rect 41583 340589 41649 340592
rect 679938 340359 679998 340474
rect 41775 340356 41841 340359
rect 41568 340354 41841 340356
rect 41568 340298 41780 340354
rect 41836 340298 41841 340354
rect 41568 340296 41841 340298
rect 679938 340354 680049 340359
rect 679938 340298 679988 340354
rect 680044 340298 680049 340354
rect 679938 340296 680049 340298
rect 41775 340293 41841 340296
rect 679983 340293 680049 340296
rect 41583 340060 41649 340063
rect 41538 340058 41649 340060
rect 41538 340002 41588 340058
rect 41644 340002 41649 340058
rect 41538 339997 41649 340002
rect 41538 339882 41598 339997
rect 679746 339767 679806 340104
rect 675706 339702 675712 339766
rect 675776 339764 675782 339766
rect 676815 339764 676881 339767
rect 675776 339762 676881 339764
rect 675776 339706 676820 339762
rect 676876 339706 676881 339762
rect 675776 339704 676881 339706
rect 679746 339762 679857 339767
rect 679983 339764 680049 339767
rect 679746 339706 679796 339762
rect 679852 339706 679857 339762
rect 679746 339704 679857 339706
rect 675776 339702 675782 339704
rect 676815 339701 676881 339704
rect 679791 339701 679857 339704
rect 679938 339762 680049 339764
rect 679938 339706 679988 339762
rect 680044 339706 680049 339762
rect 679938 339701 680049 339706
rect 679938 339586 679998 339701
rect 41538 339175 41598 339290
rect 676666 339258 676672 339322
rect 676736 339320 676742 339322
rect 676911 339320 676977 339323
rect 679791 339320 679857 339323
rect 676736 339318 676977 339320
rect 676736 339262 676916 339318
rect 676972 339262 676977 339318
rect 676736 339260 676977 339262
rect 676736 339258 676742 339260
rect 676911 339257 676977 339260
rect 679746 339318 679857 339320
rect 679746 339262 679796 339318
rect 679852 339262 679857 339318
rect 679746 339257 679857 339262
rect 41538 339170 41649 339175
rect 41538 339114 41588 339170
rect 41644 339114 41649 339170
rect 41538 339112 41649 339114
rect 41583 339109 41649 339112
rect 679746 338994 679806 339257
rect 41775 338876 41841 338879
rect 41568 338874 41841 338876
rect 41568 338818 41780 338874
rect 41836 338818 41841 338874
rect 41568 338816 41841 338818
rect 41775 338813 41841 338816
rect 676474 338814 676480 338878
rect 676544 338876 676550 338878
rect 677007 338876 677073 338879
rect 676544 338874 677073 338876
rect 676544 338818 677012 338874
rect 677068 338818 677073 338874
rect 676544 338816 677073 338818
rect 676544 338814 676550 338816
rect 677007 338813 677073 338816
rect 42874 338432 42880 338434
rect 41568 338372 42880 338432
rect 42874 338370 42880 338372
rect 42944 338370 42950 338434
rect 40386 337546 40446 337810
rect 40378 337482 40384 337546
rect 40448 337482 40454 337546
rect 40578 337102 40638 337292
rect 40570 337038 40576 337102
rect 40640 337038 40646 337102
rect 42298 336952 42304 336954
rect 41568 336892 42304 336952
rect 42298 336890 42304 336892
rect 42368 336890 42374 336954
rect 42490 336360 42496 336362
rect 41568 336300 42496 336360
rect 42490 336298 42496 336300
rect 42560 336298 42566 336362
rect 34434 335623 34494 335738
rect 34434 335618 34545 335623
rect 34434 335562 34484 335618
rect 34540 335562 34545 335618
rect 34434 335560 34545 335562
rect 34479 335557 34545 335560
rect 40770 335030 40830 335442
rect 40762 334966 40768 335030
rect 40832 334966 40838 335030
rect 41154 334586 41214 334850
rect 41146 334522 41152 334586
rect 41216 334522 41222 334586
rect 40962 334142 41022 334258
rect 40954 334078 40960 334142
rect 41024 334078 41030 334142
rect 675130 333930 675136 333994
rect 675200 333992 675206 333994
rect 675375 333992 675441 333995
rect 675200 333990 675441 333992
rect 675200 333934 675380 333990
rect 675436 333934 675441 333990
rect 675200 333932 675441 333934
rect 675200 333930 675206 333932
rect 675375 333929 675441 333932
rect 41538 333550 41598 333888
rect 41530 333486 41536 333550
rect 41600 333486 41606 333550
rect 42106 333400 42112 333402
rect 41568 333340 42112 333400
rect 42106 333338 42112 333340
rect 42176 333338 42182 333402
rect 41346 332662 41406 332778
rect 41338 332598 41344 332662
rect 41408 332598 41414 332662
rect 41914 332438 41920 332440
rect 41568 332378 41920 332438
rect 41914 332376 41920 332378
rect 41984 332376 41990 332440
rect 673978 332302 673984 332366
rect 674048 332364 674054 332366
rect 675471 332364 675537 332367
rect 674048 332362 675537 332364
rect 674048 332306 675476 332362
rect 675532 332306 675537 332362
rect 674048 332304 675537 332306
rect 674048 332302 674054 332304
rect 675471 332301 675537 332304
rect 41722 331920 41728 331922
rect 41568 331860 41728 331920
rect 41722 331858 41728 331860
rect 41792 331858 41798 331922
rect 41538 331180 41598 331298
rect 41538 331120 41790 331180
rect 28866 330591 28926 330854
rect 41730 330736 41790 331120
rect 674938 331118 674944 331182
rect 675008 331180 675014 331182
rect 675375 331180 675441 331183
rect 675008 331178 675441 331180
rect 675008 331122 675380 331178
rect 675436 331122 675441 331178
rect 675008 331120 675441 331122
rect 675008 331118 675014 331120
rect 675375 331117 675441 331120
rect 28815 330586 28926 330591
rect 28815 330530 28820 330586
rect 28876 330530 28926 330586
rect 28815 330528 28926 330530
rect 41538 330676 41790 330736
rect 28815 330525 28881 330528
rect 41538 330440 41598 330676
rect 41775 330440 41841 330443
rect 41538 330438 41841 330440
rect 41538 330410 41780 330438
rect 41568 330382 41780 330410
rect 41836 330382 41841 330438
rect 41568 330380 41841 330382
rect 41775 330377 41841 330380
rect 28815 330144 28881 330147
rect 28815 330142 28926 330144
rect 28815 330086 28820 330142
rect 28876 330086 28926 330142
rect 28815 330081 28926 330086
rect 28866 329818 28926 330081
rect 655215 329848 655281 329851
rect 649986 329846 655281 329848
rect 649986 329790 655220 329846
rect 655276 329790 655281 329846
rect 649986 329788 655281 329790
rect 649986 329234 650046 329788
rect 655215 329785 655281 329788
rect 655119 328072 655185 328075
rect 649986 328070 655185 328072
rect 649986 328014 655124 328070
rect 655180 328014 655185 328070
rect 649986 328012 655185 328014
rect 655119 328009 655185 328012
rect 674746 327862 674752 327926
rect 674816 327924 674822 327926
rect 675375 327924 675441 327927
rect 674816 327922 675441 327924
rect 674816 327866 675380 327922
rect 675436 327866 675441 327922
rect 674816 327864 675441 327866
rect 674816 327862 674822 327864
rect 675375 327861 675441 327864
rect 655311 327480 655377 327483
rect 649986 327478 655377 327480
rect 649986 327422 655316 327478
rect 655372 327422 655377 327478
rect 649986 327420 655377 327422
rect 649986 326870 650046 327420
rect 655311 327417 655377 327420
rect 654159 326296 654225 326299
rect 649986 326294 654225 326296
rect 649986 326238 654164 326294
rect 654220 326238 654225 326294
rect 649986 326236 654225 326238
rect 649986 325688 650046 326236
rect 654159 326233 654225 326236
rect 40378 325050 40384 325114
rect 40448 325112 40454 325114
rect 41775 325112 41841 325115
rect 40448 325110 41841 325112
rect 40448 325054 41780 325110
rect 41836 325054 41841 325110
rect 40448 325052 41841 325054
rect 40448 325050 40454 325052
rect 41775 325049 41841 325052
rect 675663 324966 675729 324967
rect 675663 324962 675712 324966
rect 675776 324964 675782 324966
rect 675663 324906 675668 324962
rect 675663 324902 675712 324906
rect 675776 324904 675820 324964
rect 675776 324902 675782 324904
rect 675663 324901 675729 324902
rect 41530 323274 41536 323338
rect 41600 323336 41606 323338
rect 41775 323336 41841 323339
rect 41600 323334 41841 323336
rect 41600 323278 41780 323334
rect 41836 323278 41841 323334
rect 41600 323276 41841 323278
rect 41600 323274 41606 323276
rect 41775 323273 41841 323276
rect 675759 323040 675825 323043
rect 676474 323040 676480 323042
rect 675759 323038 676480 323040
rect 675759 322982 675764 323038
rect 675820 322982 676480 323038
rect 675759 322980 676480 322982
rect 675759 322977 675825 322980
rect 676474 322978 676480 322980
rect 676544 322978 676550 323042
rect 41775 321858 41841 321859
rect 41722 321856 41728 321858
rect 41684 321796 41728 321856
rect 41792 321854 41841 321858
rect 41836 321798 41841 321854
rect 41722 321794 41728 321796
rect 41792 321794 41841 321798
rect 41775 321793 41841 321794
rect 42063 321266 42129 321267
rect 42063 321262 42112 321266
rect 42176 321264 42182 321266
rect 675759 321264 675825 321267
rect 676666 321264 676672 321266
rect 42063 321206 42068 321262
rect 42063 321202 42112 321206
rect 42176 321204 42220 321264
rect 675759 321262 676672 321264
rect 675759 321206 675764 321262
rect 675820 321206 676672 321262
rect 675759 321204 676672 321206
rect 42176 321202 42182 321204
rect 42063 321201 42129 321202
rect 675759 321201 675825 321204
rect 676666 321202 676672 321204
rect 676736 321202 676742 321266
rect 41871 320822 41937 320823
rect 41871 320818 41920 320822
rect 41984 320820 41990 320822
rect 41871 320762 41876 320818
rect 41871 320758 41920 320762
rect 41984 320760 42028 320820
rect 41984 320758 41990 320760
rect 41871 320757 41937 320758
rect 42063 319932 42129 319935
rect 42490 319932 42496 319934
rect 42063 319930 42496 319932
rect 42063 319874 42068 319930
rect 42124 319874 42496 319930
rect 42063 319872 42496 319874
rect 42063 319869 42129 319872
rect 42490 319870 42496 319872
rect 42560 319870 42566 319934
rect 41338 317650 41344 317714
rect 41408 317712 41414 317714
rect 41871 317712 41937 317715
rect 41408 317710 41937 317712
rect 41408 317654 41876 317710
rect 41932 317654 41937 317710
rect 41408 317652 41937 317654
rect 41408 317650 41414 317652
rect 41871 317649 41937 317652
rect 58479 317712 58545 317715
rect 58479 317710 64638 317712
rect 58479 317654 58484 317710
rect 58540 317654 64638 317710
rect 58479 317652 64638 317654
rect 58479 317649 58545 317652
rect 64578 317106 64638 317652
rect 40954 316762 40960 316826
rect 41024 316824 41030 316826
rect 41775 316824 41841 316827
rect 41024 316822 41841 316824
rect 41024 316766 41780 316822
rect 41836 316766 41841 316822
rect 41024 316764 41841 316766
rect 41024 316762 41030 316764
rect 41775 316761 41841 316764
rect 59151 316528 59217 316531
rect 59151 316526 64638 316528
rect 59151 316470 59156 316526
rect 59212 316470 64638 316526
rect 59151 316468 64638 316470
rect 59151 316465 59217 316468
rect 41146 316170 41152 316234
rect 41216 316232 41222 316234
rect 41775 316232 41841 316235
rect 41216 316230 41841 316232
rect 41216 316174 41780 316230
rect 41836 316174 41841 316230
rect 41216 316172 41841 316174
rect 41216 316170 41222 316172
rect 41775 316169 41841 316172
rect 64578 315924 64638 316468
rect 41338 315578 41344 315642
rect 41408 315640 41414 315642
rect 41775 315640 41841 315643
rect 41408 315638 41841 315640
rect 41408 315582 41780 315638
rect 41836 315582 41841 315638
rect 41408 315580 41841 315582
rect 41408 315578 41414 315580
rect 41775 315577 41841 315580
rect 59055 314160 59121 314163
rect 64578 314160 64638 314742
rect 59055 314158 64638 314160
rect 59055 314102 59060 314158
rect 59116 314102 64638 314158
rect 59055 314100 64638 314102
rect 59055 314097 59121 314100
rect 674554 313950 674560 314014
rect 674624 314012 674630 314014
rect 679887 314012 679953 314015
rect 674624 314010 679953 314012
rect 674624 313954 679892 314010
rect 679948 313954 679953 314010
rect 674624 313952 679953 313954
rect 674624 313950 674630 313952
rect 679887 313949 679953 313952
rect 42159 313864 42225 313867
rect 42874 313864 42880 313866
rect 42159 313862 42880 313864
rect 42159 313806 42164 313862
rect 42220 313806 42880 313862
rect 42159 313804 42880 313806
rect 42159 313801 42225 313804
rect 42874 313802 42880 313804
rect 42944 313802 42950 313866
rect 59631 313568 59697 313571
rect 59631 313566 64638 313568
rect 59631 313510 59636 313566
rect 59692 313510 64638 313566
rect 59631 313508 64638 313510
rect 59631 313505 59697 313508
rect 40762 313210 40768 313274
rect 40832 313272 40838 313274
rect 41775 313272 41841 313275
rect 40832 313270 41841 313272
rect 40832 313214 41780 313270
rect 41836 313214 41841 313270
rect 40832 313212 41841 313214
rect 40832 313210 40838 313212
rect 41775 313209 41841 313212
rect 59727 312976 59793 312979
rect 59727 312974 64638 312976
rect 59727 312918 59732 312974
rect 59788 312918 64638 312974
rect 59727 312916 64638 312918
rect 59727 312913 59793 312916
rect 40570 312618 40576 312682
rect 40640 312680 40646 312682
rect 41775 312680 41841 312683
rect 40640 312678 41841 312680
rect 40640 312622 41780 312678
rect 41836 312622 41841 312678
rect 40640 312620 41841 312622
rect 40640 312618 40646 312620
rect 41775 312617 41841 312620
rect 64578 312378 64638 312916
rect 59535 311792 59601 311795
rect 59535 311790 64638 311792
rect 59535 311734 59540 311790
rect 59596 311734 64638 311790
rect 59535 311732 64638 311734
rect 59535 311729 59601 311732
rect 64578 311196 64638 311732
rect 676290 305727 676350 306064
rect 676239 305722 676350 305727
rect 676239 305666 676244 305722
rect 676300 305666 676350 305722
rect 676239 305664 676350 305666
rect 676239 305661 676305 305664
rect 676290 305283 676350 305546
rect 676239 305278 676350 305283
rect 676239 305222 676244 305278
rect 676300 305222 676350 305278
rect 676239 305220 676350 305222
rect 676239 305217 676305 305220
rect 676290 304839 676350 304954
rect 676239 304834 676350 304839
rect 676239 304778 676244 304834
rect 676300 304778 676350 304834
rect 676239 304776 676350 304778
rect 679887 304836 679953 304839
rect 679887 304834 679998 304836
rect 679887 304778 679892 304834
rect 679948 304778 679998 304834
rect 676239 304773 676305 304776
rect 679887 304773 679998 304778
rect 679938 304584 679998 304773
rect 676047 304096 676113 304099
rect 676047 304094 676320 304096
rect 676047 304038 676052 304094
rect 676108 304038 676320 304094
rect 676047 304036 676320 304038
rect 676047 304033 676113 304036
rect 672687 303504 672753 303507
rect 675322 303504 675328 303506
rect 672687 303502 675328 303504
rect 672687 303446 672692 303502
rect 672748 303446 675328 303502
rect 672687 303444 675328 303446
rect 672687 303441 672753 303444
rect 675322 303442 675328 303444
rect 675392 303504 675398 303506
rect 675392 303444 676320 303504
rect 675392 303442 675398 303444
rect 653775 303356 653841 303359
rect 649986 303354 653841 303356
rect 649986 303298 653780 303354
rect 653836 303298 653841 303354
rect 649986 303296 653841 303298
rect 649986 302776 650046 303296
rect 653775 303293 653841 303296
rect 676047 303060 676113 303063
rect 676047 303058 676320 303060
rect 676047 303002 676052 303058
rect 676108 303002 676320 303058
rect 676047 303000 676320 303002
rect 676047 302997 676113 303000
rect 672879 302616 672945 302619
rect 674362 302616 674368 302618
rect 672879 302614 674368 302616
rect 672879 302558 672884 302614
rect 672940 302558 674368 302614
rect 672879 302556 674368 302558
rect 672879 302553 672945 302556
rect 674362 302554 674368 302556
rect 674432 302616 674438 302618
rect 674432 302556 676320 302616
rect 674432 302554 674438 302556
rect 654063 302172 654129 302175
rect 649986 302170 654129 302172
rect 649986 302114 654068 302170
rect 654124 302114 654129 302170
rect 649986 302112 654129 302114
rect 649986 301594 650046 302112
rect 654063 302109 654129 302112
rect 676047 302024 676113 302027
rect 676047 302022 676320 302024
rect 676047 301966 676052 302022
rect 676108 301966 676320 302022
rect 676047 301964 676320 301966
rect 676047 301961 676113 301964
rect 675706 301518 675712 301582
rect 675776 301580 675782 301582
rect 675776 301520 676320 301580
rect 675776 301518 675782 301520
rect 654159 300988 654225 300991
rect 649986 300986 654225 300988
rect 649986 300930 654164 300986
rect 654220 300930 654225 300986
rect 649986 300928 654225 300930
rect 649986 300412 650046 300928
rect 654159 300925 654225 300928
rect 674170 300630 674176 300694
rect 674240 300692 674246 300694
rect 676290 300692 676350 301032
rect 674240 300632 676350 300692
rect 674240 300630 674246 300632
rect 675898 300482 675904 300546
rect 675968 300544 675974 300546
rect 675968 300484 676320 300544
rect 675968 300482 675974 300484
rect 676482 299806 676542 300070
rect 676474 299742 676480 299806
rect 676544 299742 676550 299806
rect 41775 299656 41841 299659
rect 41568 299654 41841 299656
rect 41568 299598 41780 299654
rect 41836 299598 41841 299654
rect 41568 299596 41841 299598
rect 41775 299593 41841 299596
rect 675130 299594 675136 299658
rect 675200 299656 675206 299658
rect 675200 299596 676350 299656
rect 675200 299594 675206 299596
rect 676290 299552 676350 299596
rect 41538 298771 41598 299182
rect 41538 298766 41649 298771
rect 41538 298710 41588 298766
rect 41644 298710 41649 298766
rect 41538 298708 41649 298710
rect 649986 298768 650046 299230
rect 674362 299002 674368 299066
rect 674432 299064 674438 299066
rect 674432 299004 676320 299064
rect 674432 299002 674438 299004
rect 656559 298768 656625 298771
rect 649986 298766 656625 298768
rect 649986 298710 656564 298766
rect 656620 298710 656625 298766
rect 649986 298708 656625 298710
rect 41583 298705 41649 298708
rect 656559 298705 656625 298708
rect 41775 298620 41841 298623
rect 41568 298618 41841 298620
rect 41568 298562 41780 298618
rect 41836 298562 41841 298618
rect 41568 298560 41841 298562
rect 41775 298557 41841 298560
rect 676047 298620 676113 298623
rect 676047 298618 676320 298620
rect 676047 298562 676052 298618
rect 676108 298562 676320 298618
rect 676047 298560 676320 298562
rect 676047 298557 676113 298560
rect 41775 298176 41841 298179
rect 41568 298174 41841 298176
rect 41568 298118 41780 298174
rect 41836 298118 41841 298174
rect 41568 298116 41841 298118
rect 41775 298113 41841 298116
rect 41775 297658 41841 297661
rect 41568 297656 41841 297658
rect 41568 297600 41780 297656
rect 41836 297600 41841 297656
rect 41568 297598 41841 297600
rect 41775 297595 41841 297598
rect 649986 297584 650046 298048
rect 676290 297734 676350 297998
rect 676282 297670 676288 297734
rect 676352 297670 676358 297734
rect 656367 297584 656433 297587
rect 649986 297582 656433 297584
rect 649986 297526 656372 297582
rect 656428 297526 656433 297582
rect 649986 297524 656433 297526
rect 656367 297521 656433 297524
rect 675322 297522 675328 297586
rect 675392 297584 675398 297586
rect 675392 297524 676320 297584
rect 675392 297522 675398 297524
rect 41775 297140 41841 297143
rect 41568 297138 41841 297140
rect 41568 297082 41780 297138
rect 41836 297082 41841 297138
rect 41568 297080 41841 297082
rect 41775 297077 41841 297080
rect 674746 297078 674752 297142
rect 674816 297140 674822 297142
rect 674816 297080 676320 297140
rect 674816 297078 674822 297080
rect 649986 296844 650046 296866
rect 656175 296844 656241 296847
rect 649986 296842 656241 296844
rect 649986 296786 656180 296842
rect 656236 296786 656241 296842
rect 649986 296784 656241 296786
rect 656175 296781 656241 296784
rect 39618 296551 39678 296670
rect 39618 296546 39729 296551
rect 39618 296490 39668 296546
rect 39724 296490 39729 296546
rect 39618 296488 39729 296490
rect 39663 296485 39729 296488
rect 676090 296190 676096 296254
rect 676160 296252 676166 296254
rect 676290 296252 676350 296518
rect 676160 296192 676350 296252
rect 676160 296190 676166 296192
rect 41538 295959 41598 296074
rect 676047 296030 676113 296033
rect 676047 296028 676320 296030
rect 676047 295972 676052 296028
rect 676108 295972 676320 296028
rect 676047 295970 676320 295972
rect 676047 295967 676113 295970
rect 39855 295956 39921 295959
rect 39810 295954 39921 295956
rect 39810 295898 39860 295954
rect 39916 295898 39921 295954
rect 39810 295893 39921 295898
rect 41538 295954 41649 295959
rect 41538 295898 41588 295954
rect 41644 295898 41649 295954
rect 41538 295896 41649 295898
rect 41583 295893 41649 295896
rect 39810 295630 39870 295893
rect 59631 295216 59697 295219
rect 64578 295216 64638 295684
rect 59631 295214 64638 295216
rect 40578 294922 40638 295186
rect 59631 295158 59636 295214
rect 59692 295158 64638 295214
rect 59631 295156 64638 295158
rect 649986 295216 650046 295684
rect 675514 295598 675520 295662
rect 675584 295660 675590 295662
rect 675584 295600 676320 295660
rect 675584 295598 675590 295600
rect 656079 295216 656145 295219
rect 649986 295214 656145 295216
rect 649986 295158 656084 295214
rect 656140 295158 656145 295214
rect 649986 295156 656145 295158
rect 59631 295153 59697 295156
rect 656079 295153 656145 295156
rect 40570 294858 40576 294922
rect 40640 294858 40646 294922
rect 676866 294774 676926 295038
rect 676858 294710 676864 294774
rect 676928 294710 676934 294774
rect 42298 294624 42304 294626
rect 41568 294564 42304 294624
rect 42298 294562 42304 294564
rect 42368 294562 42374 294626
rect 42682 294180 42688 294182
rect 41568 294120 42688 294180
rect 42682 294118 42688 294120
rect 42752 294118 42758 294182
rect 58191 294032 58257 294035
rect 64578 294032 64638 294502
rect 58191 294030 64638 294032
rect 58191 293974 58196 294030
rect 58252 293974 64638 294030
rect 58191 293972 64638 293974
rect 649986 294032 650046 294502
rect 679938 294331 679998 294520
rect 679887 294326 679998 294331
rect 679887 294270 679892 294326
rect 679948 294270 679998 294326
rect 679887 294268 679998 294270
rect 679887 294265 679953 294268
rect 655887 294032 655953 294035
rect 649986 294030 655953 294032
rect 649986 293974 655892 294030
rect 655948 293974 655953 294030
rect 649986 293972 655953 293974
rect 58191 293969 58257 293972
rect 655887 293969 655953 293972
rect 679746 293887 679806 294150
rect 679695 293882 679806 293887
rect 679695 293826 679700 293882
rect 679756 293826 679806 293882
rect 679695 293824 679806 293826
rect 679887 293884 679953 293887
rect 679887 293882 679998 293884
rect 679887 293826 679892 293882
rect 679948 293826 679998 293882
rect 679695 293821 679761 293824
rect 679887 293821 679998 293826
rect 40962 293442 41022 293706
rect 679938 293558 679998 293821
rect 40954 293378 40960 293442
rect 41024 293378 41030 293442
rect 42490 293144 42496 293146
rect 41568 293084 42496 293144
rect 42490 293082 42496 293084
rect 42560 293082 42566 293146
rect 59055 292848 59121 292851
rect 64578 292848 64638 293320
rect 59055 292846 64638 292848
rect 59055 292790 59060 292846
rect 59116 292790 64638 292846
rect 59055 292788 64638 292790
rect 649986 292848 650046 293320
rect 679695 293292 679761 293295
rect 679695 293290 679806 293292
rect 679695 293234 679700 293290
rect 679756 293234 679806 293290
rect 679695 293229 679806 293234
rect 679746 292966 679806 293229
rect 655791 292848 655857 292851
rect 649986 292846 655857 292848
rect 649986 292790 655796 292846
rect 655852 292790 655857 292846
rect 649986 292788 655857 292790
rect 59055 292785 59121 292788
rect 655791 292785 655857 292788
rect 34434 292407 34494 292596
rect 34434 292402 34545 292407
rect 34434 292346 34484 292402
rect 34540 292346 34545 292402
rect 34434 292344 34545 292346
rect 34479 292341 34545 292344
rect 40770 291962 40830 292226
rect 40762 291898 40768 291962
rect 40832 291898 40838 291962
rect 59631 291664 59697 291667
rect 64578 291664 64638 292138
rect 59631 291662 64638 291664
rect 41346 291370 41406 291634
rect 59631 291606 59636 291662
rect 59692 291606 64638 291662
rect 59631 291604 64638 291606
rect 649986 291664 650046 292138
rect 655983 291664 656049 291667
rect 649986 291662 656049 291664
rect 649986 291606 655988 291662
rect 656044 291606 656049 291662
rect 649986 291604 656049 291606
rect 59631 291601 59697 291604
rect 655983 291601 656049 291604
rect 60207 291516 60273 291519
rect 60207 291514 64638 291516
rect 60207 291458 60212 291514
rect 60268 291458 64638 291514
rect 60207 291456 64638 291458
rect 60207 291453 60273 291456
rect 41338 291306 41344 291370
rect 41408 291306 41414 291370
rect 41154 290926 41214 291042
rect 64578 290956 64638 291456
rect 41146 290862 41152 290926
rect 41216 290862 41222 290926
rect 649986 290924 650046 290956
rect 655599 290924 655665 290927
rect 649986 290922 655665 290924
rect 649986 290866 655604 290922
rect 655660 290866 655665 290922
rect 649986 290864 655665 290866
rect 655599 290861 655665 290864
rect 41538 290334 41598 290746
rect 675759 290628 675825 290631
rect 675898 290628 675904 290630
rect 675759 290626 675904 290628
rect 675759 290570 675764 290626
rect 675820 290570 675904 290626
rect 675759 290568 675904 290570
rect 675759 290565 675825 290568
rect 675898 290566 675904 290568
rect 675968 290566 675974 290630
rect 41530 290270 41536 290334
rect 41600 290270 41606 290334
rect 57519 290332 57585 290335
rect 57519 290330 64638 290332
rect 57519 290274 57524 290330
rect 57580 290274 64638 290330
rect 57519 290272 64638 290274
rect 57519 290269 57585 290272
rect 42106 290184 42112 290186
rect 41568 290124 42112 290184
rect 42106 290122 42112 290124
rect 42176 290122 42182 290186
rect 64578 289774 64638 290272
rect 40386 289446 40446 289562
rect 40378 289382 40384 289446
rect 40448 289382 40454 289446
rect 649986 289296 650046 289774
rect 675759 289742 675825 289743
rect 675706 289678 675712 289742
rect 675776 289740 675825 289742
rect 675776 289738 675868 289740
rect 675820 289682 675868 289738
rect 675776 289680 675868 289682
rect 675776 289678 675825 289680
rect 675759 289677 675825 289678
rect 654159 289296 654225 289299
rect 649986 289294 654225 289296
rect 649986 289238 654164 289294
rect 654220 289238 654225 289294
rect 649986 289236 654225 289238
rect 654159 289233 654225 289236
rect 41914 289222 41920 289224
rect 41568 289162 41920 289222
rect 41914 289160 41920 289162
rect 41984 289160 41990 289224
rect 41722 288704 41728 288706
rect 41568 288644 41728 288704
rect 41722 288642 41728 288644
rect 41792 288642 41798 288706
rect 59631 288112 59697 288115
rect 64578 288112 64638 288592
rect 59631 288110 64638 288112
rect 41538 287964 41598 288082
rect 59631 288054 59636 288110
rect 59692 288054 64638 288110
rect 59631 288052 64638 288054
rect 649986 288112 650046 288592
rect 655407 288112 655473 288115
rect 649986 288110 655473 288112
rect 649986 288054 655412 288110
rect 655468 288054 655473 288110
rect 649986 288052 655473 288054
rect 59631 288049 59697 288052
rect 655407 288049 655473 288052
rect 675759 287964 675825 287967
rect 676474 287964 676480 287966
rect 41538 287904 41790 287964
rect 28866 287375 28926 287712
rect 41730 287520 41790 287904
rect 675759 287962 676480 287964
rect 675759 287906 675764 287962
rect 675820 287906 676480 287962
rect 675759 287904 676480 287906
rect 675759 287901 675825 287904
rect 676474 287902 676480 287904
rect 676544 287902 676550 287966
rect 28815 287370 28926 287375
rect 28815 287314 28820 287370
rect 28876 287314 28926 287370
rect 28815 287312 28926 287314
rect 41538 287460 41790 287520
rect 675759 287520 675825 287523
rect 676282 287520 676288 287522
rect 675759 287518 676288 287520
rect 675759 287462 675764 287518
rect 675820 287462 676288 287518
rect 675759 287460 676288 287462
rect 28815 287309 28881 287312
rect 41538 287224 41598 287460
rect 675759 287457 675825 287460
rect 676282 287458 676288 287460
rect 676352 287458 676358 287522
rect 41775 287224 41841 287227
rect 41538 287222 41841 287224
rect 41538 287194 41780 287222
rect 41568 287166 41780 287194
rect 41836 287166 41841 287222
rect 41568 287164 41841 287166
rect 41775 287161 41841 287164
rect 28815 286928 28881 286931
rect 58095 286928 58161 286931
rect 64578 286928 64638 287410
rect 28815 286926 28926 286928
rect 28815 286870 28820 286926
rect 28876 286870 28926 286926
rect 28815 286865 28926 286870
rect 58095 286926 64638 286928
rect 58095 286870 58100 286926
rect 58156 286870 64638 286926
rect 58095 286868 64638 286870
rect 649986 286928 650046 287410
rect 655503 286928 655569 286931
rect 675375 286930 675441 286931
rect 675322 286928 675328 286930
rect 649986 286926 655569 286928
rect 649986 286870 655508 286926
rect 655564 286870 655569 286926
rect 649986 286868 655569 286870
rect 675284 286868 675328 286928
rect 675392 286926 675441 286930
rect 675436 286870 675441 286926
rect 58095 286865 58161 286868
rect 655503 286865 655569 286868
rect 675322 286866 675328 286868
rect 675392 286866 675441 286870
rect 675375 286865 675441 286866
rect 28866 286602 28926 286865
rect 59535 285744 59601 285747
rect 64578 285744 64638 286228
rect 59535 285742 64638 285744
rect 59535 285686 59540 285742
rect 59596 285686 64638 285742
rect 59535 285684 64638 285686
rect 649986 285744 650046 286228
rect 655695 285744 655761 285747
rect 649986 285742 655761 285744
rect 649986 285686 655700 285742
rect 655756 285686 655761 285742
rect 649986 285684 655761 285686
rect 59535 285681 59601 285684
rect 655695 285681 655761 285684
rect 57615 284560 57681 284563
rect 64578 284560 64638 285046
rect 57615 284558 64638 284560
rect 57615 284502 57620 284558
rect 57676 284502 64638 284558
rect 57615 284500 64638 284502
rect 649986 284560 650046 285046
rect 653775 284560 653841 284563
rect 649986 284558 653841 284560
rect 649986 284502 653780 284558
rect 653836 284502 653841 284558
rect 649986 284500 653841 284502
rect 57615 284497 57681 284500
rect 653775 284497 653841 284500
rect 59631 283376 59697 283379
rect 64578 283376 64638 283864
rect 59631 283374 64638 283376
rect 59631 283318 59636 283374
rect 59692 283318 64638 283374
rect 59631 283316 64638 283318
rect 649986 283376 650046 283864
rect 675130 283758 675136 283822
rect 675200 283820 675206 283822
rect 675375 283820 675441 283823
rect 675200 283818 675441 283820
rect 675200 283762 675380 283818
rect 675436 283762 675441 283818
rect 675200 283760 675441 283762
rect 675200 283758 675206 283760
rect 675375 283757 675441 283760
rect 655119 283376 655185 283379
rect 649986 283374 655185 283376
rect 649986 283318 655124 283374
rect 655180 283318 655185 283374
rect 649986 283316 655185 283318
rect 59631 283313 59697 283316
rect 655119 283313 655185 283316
rect 675567 282934 675633 282935
rect 675514 282870 675520 282934
rect 675584 282932 675633 282934
rect 675584 282930 675676 282932
rect 675628 282874 675676 282930
rect 675584 282872 675676 282874
rect 675584 282870 675633 282872
rect 675567 282869 675633 282870
rect 58959 282488 59025 282491
rect 64578 282488 64638 282682
rect 58959 282486 64638 282488
rect 58959 282430 58964 282486
rect 59020 282430 64638 282486
rect 58959 282428 64638 282430
rect 58959 282425 59025 282428
rect 649986 282340 650046 282682
rect 655311 282340 655377 282343
rect 676858 282340 676864 282342
rect 649986 282338 655377 282340
rect 649986 282282 655316 282338
rect 655372 282282 655377 282338
rect 649986 282280 655377 282282
rect 655311 282277 655377 282280
rect 675522 282280 676864 282340
rect 42063 281896 42129 281899
rect 42298 281896 42304 281898
rect 42063 281894 42304 281896
rect 42063 281838 42068 281894
rect 42124 281838 42304 281894
rect 42063 281836 42304 281838
rect 42063 281833 42129 281836
rect 42298 281834 42304 281836
rect 42368 281834 42374 281898
rect 675522 281751 675582 282280
rect 676858 282278 676864 282280
rect 676928 282278 676934 282342
rect 675663 281896 675729 281899
rect 676090 281896 676096 281898
rect 675663 281894 676096 281896
rect 675663 281838 675668 281894
rect 675724 281838 676096 281894
rect 675663 281836 676096 281838
rect 675663 281833 675729 281836
rect 676090 281834 676096 281836
rect 676160 281834 676166 281898
rect 675522 281746 675633 281751
rect 675522 281690 675572 281746
rect 675628 281690 675633 281746
rect 675522 281688 675633 281690
rect 675567 281685 675633 281688
rect 58191 281008 58257 281011
rect 64578 281008 64638 281500
rect 58191 281006 64638 281008
rect 58191 280950 58196 281006
rect 58252 280950 64638 281006
rect 58191 280948 64638 280950
rect 649986 281008 650046 281500
rect 655215 281008 655281 281011
rect 649986 281006 655281 281008
rect 649986 280950 655220 281006
rect 655276 280950 655281 281006
rect 649986 280948 655281 280950
rect 58191 280945 58257 280948
rect 655215 280945 655281 280948
rect 674746 280650 674752 280714
rect 674816 280712 674822 280714
rect 675375 280712 675441 280715
rect 674816 280710 675441 280712
rect 674816 280654 675380 280710
rect 675436 280654 675441 280710
rect 674816 280652 675441 280654
rect 674816 280650 674822 280652
rect 675375 280649 675441 280652
rect 41530 280058 41536 280122
rect 41600 280120 41606 280122
rect 41775 280120 41841 280123
rect 41600 280118 41841 280120
rect 41600 280062 41780 280118
rect 41836 280062 41841 280118
rect 41600 280060 41841 280062
rect 41600 280058 41606 280060
rect 41775 280057 41841 280060
rect 59631 279824 59697 279827
rect 64578 279824 64638 280318
rect 59631 279822 64638 279824
rect 59631 279766 59636 279822
rect 59692 279766 64638 279822
rect 59631 279764 64638 279766
rect 649986 279824 650046 280318
rect 654735 279824 654801 279827
rect 649986 279822 654801 279824
rect 649986 279766 654740 279822
rect 654796 279766 654801 279822
rect 649986 279764 654801 279766
rect 59631 279761 59697 279764
rect 654735 279761 654801 279764
rect 674170 278874 674176 278938
rect 674240 278936 674246 278938
rect 675375 278936 675441 278939
rect 674240 278934 675441 278936
rect 674240 278878 675380 278934
rect 675436 278878 675441 278934
rect 674240 278876 675441 278878
rect 674240 278874 674246 278876
rect 675375 278873 675441 278876
rect 41775 278790 41841 278791
rect 41722 278788 41728 278790
rect 41684 278728 41728 278788
rect 41792 278786 41841 278790
rect 41836 278730 41841 278786
rect 41722 278726 41728 278728
rect 41792 278726 41841 278730
rect 41775 278725 41841 278726
rect 45039 278640 45105 278643
rect 674938 278640 674944 278642
rect 45039 278638 674944 278640
rect 45039 278582 45044 278638
rect 45100 278582 674944 278638
rect 45039 278580 674944 278582
rect 45039 278577 45105 278580
rect 674938 278578 674944 278580
rect 675008 278578 675014 278642
rect 44463 278492 44529 278495
rect 672495 278492 672561 278495
rect 44463 278490 672561 278492
rect 44463 278434 44468 278490
rect 44524 278434 672500 278490
rect 672556 278434 672561 278490
rect 44463 278432 672561 278434
rect 44463 278429 44529 278432
rect 672495 278429 672561 278432
rect 45423 278344 45489 278347
rect 670287 278344 670353 278347
rect 45423 278342 670353 278344
rect 45423 278286 45428 278342
rect 45484 278286 670292 278342
rect 670348 278286 670353 278342
rect 45423 278284 670353 278286
rect 45423 278281 45489 278284
rect 670287 278281 670353 278284
rect 45999 278196 46065 278199
rect 670479 278196 670545 278199
rect 45999 278194 670545 278196
rect 45999 278138 46004 278194
rect 46060 278138 670484 278194
rect 670540 278138 670545 278194
rect 45999 278136 670545 278138
rect 45999 278133 46065 278136
rect 670479 278133 670545 278136
rect 42063 278050 42129 278051
rect 42063 278046 42112 278050
rect 42176 278048 42182 278050
rect 62127 278048 62193 278051
rect 672687 278048 672753 278051
rect 42063 277990 42068 278046
rect 42063 277986 42112 277990
rect 42176 277988 42220 278048
rect 62127 278046 672753 278048
rect 62127 277990 62132 278046
rect 62188 277990 672692 278046
rect 672748 277990 672753 278046
rect 62127 277988 672753 277990
rect 42176 277986 42182 277988
rect 42063 277985 42129 277986
rect 62127 277985 62193 277988
rect 672687 277985 672753 277988
rect 44847 277900 44913 277903
rect 668175 277900 668241 277903
rect 44847 277898 668241 277900
rect 44847 277842 44852 277898
rect 44908 277842 668180 277898
rect 668236 277842 668241 277898
rect 44847 277840 668241 277842
rect 44847 277837 44913 277840
rect 668175 277837 668241 277840
rect 62319 277752 62385 277755
rect 672879 277752 672945 277755
rect 62319 277750 672945 277752
rect 62319 277694 62324 277750
rect 62380 277694 672884 277750
rect 672940 277694 672945 277750
rect 62319 277692 672945 277694
rect 62319 277689 62385 277692
rect 672879 277689 672945 277692
rect 41871 277606 41937 277607
rect 41871 277602 41920 277606
rect 41984 277604 41990 277606
rect 62703 277604 62769 277607
rect 670095 277604 670161 277607
rect 41871 277546 41876 277602
rect 41871 277542 41920 277546
rect 41984 277544 42028 277604
rect 62703 277602 670161 277604
rect 62703 277546 62708 277602
rect 62764 277546 670100 277602
rect 670156 277546 670161 277602
rect 62703 277544 670161 277546
rect 41984 277542 41990 277544
rect 41871 277541 41937 277542
rect 62703 277541 62769 277544
rect 670095 277541 670161 277544
rect 40570 277394 40576 277458
rect 40640 277456 40646 277458
rect 41914 277456 41920 277458
rect 40640 277396 41920 277456
rect 40640 277394 40646 277396
rect 41914 277394 41920 277396
rect 41984 277394 41990 277458
rect 62799 277456 62865 277459
rect 669903 277456 669969 277459
rect 62799 277454 669969 277456
rect 62799 277398 62804 277454
rect 62860 277398 669908 277454
rect 669964 277398 669969 277454
rect 62799 277396 669969 277398
rect 62799 277393 62865 277396
rect 669903 277393 669969 277396
rect 44655 277308 44721 277311
rect 646575 277308 646641 277311
rect 44655 277306 646641 277308
rect 44655 277250 44660 277306
rect 44716 277250 646580 277306
rect 646636 277250 646641 277306
rect 44655 277248 646641 277250
rect 44655 277245 44721 277248
rect 646575 277245 646641 277248
rect 674362 276950 674368 277014
rect 674432 277012 674438 277014
rect 675375 277012 675441 277015
rect 674432 277010 675441 277012
rect 674432 276954 675380 277010
rect 675436 276954 675441 277010
rect 674432 276952 675441 276954
rect 674432 276950 674438 276952
rect 675375 276949 675441 276952
rect 42063 276716 42129 276719
rect 42490 276716 42496 276718
rect 42063 276714 42496 276716
rect 42063 276658 42068 276714
rect 42124 276658 42496 276714
rect 42063 276656 42496 276658
rect 42063 276653 42129 276656
rect 42490 276654 42496 276656
rect 42560 276654 42566 276718
rect 402543 276716 402609 276719
rect 529839 276716 529905 276719
rect 402543 276714 529905 276716
rect 402543 276658 402548 276714
rect 402604 276658 529844 276714
rect 529900 276658 529905 276714
rect 402543 276656 529905 276658
rect 402543 276653 402609 276656
rect 529839 276653 529905 276656
rect 396687 276568 396753 276571
rect 610767 276568 610833 276571
rect 396687 276566 610833 276568
rect 396687 276510 396692 276566
rect 396748 276510 610772 276566
rect 610828 276510 610833 276566
rect 396687 276508 610833 276510
rect 396687 276505 396753 276508
rect 610767 276505 610833 276508
rect 45135 276420 45201 276423
rect 673263 276420 673329 276423
rect 45135 276418 673329 276420
rect 45135 276362 45140 276418
rect 45196 276362 673268 276418
rect 673324 276362 673329 276418
rect 45135 276360 673329 276362
rect 45135 276357 45201 276360
rect 673263 276357 673329 276360
rect 44367 276272 44433 276275
rect 672399 276272 672465 276275
rect 44367 276270 672465 276272
rect 44367 276214 44372 276270
rect 44428 276214 672404 276270
rect 672460 276214 672465 276270
rect 44367 276212 672465 276214
rect 44367 276209 44433 276212
rect 672399 276209 672465 276212
rect 61935 276124 62001 276127
rect 673167 276124 673233 276127
rect 61935 276122 673233 276124
rect 61935 276066 61940 276122
rect 61996 276066 673172 276122
rect 673228 276066 673233 276122
rect 61935 276064 673233 276066
rect 61935 276061 62001 276064
rect 673167 276061 673233 276064
rect 381807 275976 381873 275979
rect 574095 275976 574161 275979
rect 381807 275974 574161 275976
rect 381807 275918 381812 275974
rect 381868 275918 574100 275974
rect 574156 275918 574161 275974
rect 381807 275916 574161 275918
rect 381807 275913 381873 275916
rect 574095 275913 574161 275916
rect 390351 275828 390417 275831
rect 595407 275828 595473 275831
rect 390351 275826 595473 275828
rect 390351 275770 390356 275826
rect 390412 275770 595412 275826
rect 595468 275770 595473 275826
rect 390351 275768 595473 275770
rect 390351 275765 390417 275768
rect 595407 275765 595473 275768
rect 408975 275680 409041 275683
rect 650415 275680 650481 275683
rect 408975 275678 650481 275680
rect 408975 275622 408980 275678
rect 409036 275622 650420 275678
rect 650476 275622 650481 275678
rect 408975 275620 650481 275622
rect 408975 275617 409041 275620
rect 650415 275617 650481 275620
rect 44559 275532 44625 275535
rect 646479 275532 646545 275535
rect 44559 275530 646545 275532
rect 44559 275474 44564 275530
rect 44620 275474 646484 275530
rect 646540 275474 646545 275530
rect 44559 275472 646545 275474
rect 44559 275469 44625 275472
rect 646479 275469 646545 275472
rect 50511 275384 50577 275387
rect 669519 275384 669585 275387
rect 50511 275382 669585 275384
rect 50511 275326 50516 275382
rect 50572 275326 669524 275382
rect 669580 275326 669585 275382
rect 50511 275324 669585 275326
rect 50511 275321 50577 275324
rect 669519 275321 669585 275324
rect 50319 275236 50385 275239
rect 669711 275236 669777 275239
rect 50319 275234 669777 275236
rect 50319 275178 50324 275234
rect 50380 275178 669716 275234
rect 669772 275178 669777 275234
rect 50319 275176 669777 275178
rect 50319 275173 50385 275176
rect 669711 275173 669777 275176
rect 44943 275088 45009 275091
rect 679887 275088 679953 275091
rect 44943 275086 679953 275088
rect 44943 275030 44948 275086
rect 45004 275030 679892 275086
rect 679948 275030 679953 275086
rect 44943 275028 679953 275030
rect 44943 275025 45009 275028
rect 679887 275025 679953 275028
rect 379119 274940 379185 274943
rect 566991 274940 567057 274943
rect 379119 274938 567057 274940
rect 379119 274882 379124 274938
rect 379180 274882 566996 274938
rect 567052 274882 567057 274938
rect 379119 274880 567057 274882
rect 379119 274877 379185 274880
rect 566991 274877 567057 274880
rect 376239 274792 376305 274795
rect 559887 274792 559953 274795
rect 376239 274790 559953 274792
rect 376239 274734 376244 274790
rect 376300 274734 559892 274790
rect 559948 274734 559953 274790
rect 376239 274732 559953 274734
rect 376239 274729 376305 274732
rect 559887 274729 559953 274732
rect 373455 274644 373521 274647
rect 552783 274644 552849 274647
rect 373455 274642 552849 274644
rect 373455 274586 373460 274642
rect 373516 274586 552788 274642
rect 552844 274586 552849 274642
rect 373455 274584 552849 274586
rect 373455 274581 373521 274584
rect 552783 274581 552849 274584
rect 40378 274434 40384 274498
rect 40448 274496 40454 274498
rect 41775 274496 41841 274499
rect 40448 274494 41841 274496
rect 40448 274438 41780 274494
rect 41836 274438 41841 274494
rect 40448 274436 41841 274438
rect 40448 274434 40454 274436
rect 41775 274433 41841 274436
rect 353391 274496 353457 274499
rect 503151 274496 503217 274499
rect 353391 274494 503217 274496
rect 353391 274438 353396 274494
rect 353452 274438 503156 274494
rect 503212 274438 503217 274494
rect 353391 274436 503217 274438
rect 353391 274433 353457 274436
rect 503151 274433 503217 274436
rect 347631 274348 347697 274351
rect 489039 274348 489105 274351
rect 347631 274346 489105 274348
rect 347631 274290 347636 274346
rect 347692 274290 489044 274346
rect 489100 274290 489105 274346
rect 347631 274288 489105 274290
rect 347631 274285 347697 274288
rect 489039 274285 489105 274288
rect 41146 273546 41152 273610
rect 41216 273608 41222 273610
rect 41775 273608 41841 273611
rect 41216 273606 41841 273608
rect 41216 273550 41780 273606
rect 41836 273550 41841 273606
rect 41216 273548 41841 273550
rect 41216 273546 41222 273548
rect 41775 273545 41841 273548
rect 381231 273608 381297 273611
rect 408975 273608 409041 273611
rect 381231 273606 409041 273608
rect 381231 273550 381236 273606
rect 381292 273550 408980 273606
rect 409036 273550 409041 273606
rect 381231 273548 409041 273550
rect 381231 273545 381297 273548
rect 408975 273545 409041 273548
rect 378639 273460 378705 273463
rect 565839 273460 565905 273463
rect 378639 273458 565905 273460
rect 378639 273402 378644 273458
rect 378700 273402 565844 273458
rect 565900 273402 565905 273458
rect 378639 273400 565905 273402
rect 378639 273397 378705 273400
rect 565839 273397 565905 273400
rect 41338 273250 41344 273314
rect 41408 273312 41414 273314
rect 41775 273312 41841 273315
rect 41408 273310 41841 273312
rect 41408 273254 41780 273310
rect 41836 273254 41841 273310
rect 41408 273252 41841 273254
rect 41408 273250 41414 273252
rect 41775 273249 41841 273252
rect 382959 273312 383025 273315
rect 576495 273312 576561 273315
rect 382959 273310 576561 273312
rect 382959 273254 382964 273310
rect 383020 273254 576500 273310
rect 576556 273254 576561 273310
rect 382959 273252 576561 273254
rect 382959 273249 383025 273252
rect 576495 273249 576561 273252
rect 387279 273164 387345 273167
rect 587151 273164 587217 273167
rect 387279 273162 587217 273164
rect 387279 273106 387284 273162
rect 387340 273106 587156 273162
rect 587212 273106 587217 273162
rect 387279 273104 587217 273106
rect 387279 273101 387345 273104
rect 587151 273101 587217 273104
rect 390159 273016 390225 273019
rect 594159 273016 594225 273019
rect 390159 273014 594225 273016
rect 390159 272958 390164 273014
rect 390220 272958 594164 273014
rect 594220 272958 594225 273014
rect 390159 272956 594225 272958
rect 390159 272953 390225 272956
rect 594159 272953 594225 272956
rect 392751 272868 392817 272871
rect 601263 272868 601329 272871
rect 392751 272866 601329 272868
rect 392751 272810 392756 272866
rect 392812 272810 601268 272866
rect 601324 272810 601329 272866
rect 392751 272808 601329 272810
rect 392751 272805 392817 272808
rect 601263 272805 601329 272808
rect 91887 272720 91953 272723
rect 200463 272720 200529 272723
rect 91887 272718 200529 272720
rect 91887 272662 91892 272718
rect 91948 272662 200468 272718
rect 200524 272662 200529 272718
rect 91887 272660 200529 272662
rect 91887 272657 91953 272660
rect 200463 272657 200529 272660
rect 398703 272720 398769 272723
rect 615471 272720 615537 272723
rect 398703 272718 615537 272720
rect 398703 272662 398708 272718
rect 398764 272662 615476 272718
rect 615532 272662 615537 272718
rect 398703 272660 615537 272662
rect 398703 272657 398769 272660
rect 615471 272657 615537 272660
rect 88335 272572 88401 272575
rect 199215 272572 199281 272575
rect 88335 272570 199281 272572
rect 88335 272514 88340 272570
rect 88396 272514 199220 272570
rect 199276 272514 199281 272570
rect 88335 272512 199281 272514
rect 88335 272509 88401 272512
rect 199215 272509 199281 272512
rect 401295 272572 401361 272575
rect 622575 272572 622641 272575
rect 401295 272570 622641 272572
rect 401295 272514 401300 272570
rect 401356 272514 622580 272570
rect 622636 272514 622641 272570
rect 401295 272512 622641 272514
rect 401295 272509 401361 272512
rect 622575 272509 622641 272512
rect 40954 272362 40960 272426
rect 41024 272424 41030 272426
rect 41775 272424 41841 272427
rect 41024 272422 41841 272424
rect 41024 272366 41780 272422
rect 41836 272366 41841 272422
rect 41024 272364 41841 272366
rect 41024 272362 41030 272364
rect 41775 272361 41841 272364
rect 78831 272424 78897 272427
rect 196623 272424 196689 272427
rect 78831 272422 196689 272424
rect 78831 272366 78836 272422
rect 78892 272366 196628 272422
rect 196684 272366 196689 272422
rect 78831 272364 196689 272366
rect 78831 272361 78897 272364
rect 196623 272361 196689 272364
rect 404175 272424 404241 272427
rect 629679 272424 629745 272427
rect 404175 272422 629745 272424
rect 404175 272366 404180 272422
rect 404236 272366 629684 272422
rect 629740 272366 629745 272422
rect 404175 272364 629745 272366
rect 404175 272361 404241 272364
rect 629679 272361 629745 272364
rect 72975 272276 73041 272279
rect 194415 272276 194481 272279
rect 72975 272274 194481 272276
rect 72975 272218 72980 272274
rect 73036 272218 194420 272274
rect 194476 272218 194481 272274
rect 72975 272216 194481 272218
rect 72975 272213 73041 272216
rect 194415 272213 194481 272216
rect 410895 272276 410961 272279
rect 646191 272276 646257 272279
rect 410895 272274 646257 272276
rect 410895 272218 410900 272274
rect 410956 272218 646196 272274
rect 646252 272218 646257 272274
rect 410895 272216 646257 272218
rect 410895 272213 410961 272216
rect 646191 272213 646257 272216
rect 70575 272128 70641 272131
rect 193743 272128 193809 272131
rect 70575 272126 193809 272128
rect 70575 272070 70580 272126
rect 70636 272070 193748 272126
rect 193804 272070 193809 272126
rect 70575 272068 193809 272070
rect 70575 272065 70641 272068
rect 193743 272065 193809 272068
rect 411759 272128 411825 272131
rect 648591 272128 648657 272131
rect 411759 272126 648657 272128
rect 411759 272070 411764 272126
rect 411820 272070 648596 272126
rect 648652 272070 648657 272126
rect 411759 272068 648657 272070
rect 411759 272065 411825 272068
rect 648591 272065 648657 272068
rect 375567 271980 375633 271983
rect 558735 271980 558801 271983
rect 375567 271978 558801 271980
rect 375567 271922 375572 271978
rect 375628 271922 558740 271978
rect 558796 271922 558801 271978
rect 375567 271920 558801 271922
rect 375567 271917 375633 271920
rect 558735 271917 558801 271920
rect 370095 271832 370161 271835
rect 544527 271832 544593 271835
rect 370095 271830 544593 271832
rect 370095 271774 370100 271830
rect 370156 271774 544532 271830
rect 544588 271774 544593 271830
rect 370095 271772 544593 271774
rect 370095 271769 370161 271772
rect 544527 271769 544593 271772
rect 369615 271684 369681 271687
rect 543375 271684 543441 271687
rect 369615 271682 543441 271684
rect 369615 271626 369620 271682
rect 369676 271626 543380 271682
rect 543436 271626 543441 271682
rect 369615 271624 543441 271626
rect 369615 271621 369681 271624
rect 543375 271621 543441 271624
rect 62511 271536 62577 271539
rect 672591 271536 672657 271539
rect 62511 271534 672657 271536
rect 62511 271478 62516 271534
rect 62572 271478 672596 271534
rect 672652 271478 672657 271534
rect 62511 271476 672657 271478
rect 62511 271473 62577 271476
rect 672591 271473 672657 271476
rect 41871 270650 41937 270651
rect 41871 270646 41920 270650
rect 41984 270648 41990 270650
rect 45231 270648 45297 270651
rect 669999 270648 670065 270651
rect 41871 270590 41876 270646
rect 41871 270586 41920 270590
rect 41984 270588 42028 270648
rect 45231 270646 670065 270648
rect 45231 270590 45236 270646
rect 45292 270590 670004 270646
rect 670060 270590 670065 270646
rect 45231 270588 670065 270590
rect 41984 270586 41990 270588
rect 41871 270585 41937 270586
rect 45231 270585 45297 270588
rect 669999 270585 670065 270588
rect 377007 270500 377073 270503
rect 562287 270500 562353 270503
rect 377007 270498 562353 270500
rect 377007 270442 377012 270498
rect 377068 270442 562292 270498
rect 562348 270442 562353 270498
rect 377007 270440 562353 270442
rect 377007 270437 377073 270440
rect 562287 270437 562353 270440
rect 385551 270352 385617 270355
rect 583599 270352 583665 270355
rect 385551 270350 583665 270352
rect 385551 270294 385556 270350
rect 385612 270294 583604 270350
rect 583660 270294 583665 270350
rect 385551 270292 583665 270294
rect 385551 270289 385617 270292
rect 583599 270289 583665 270292
rect 388431 270204 388497 270207
rect 590607 270204 590673 270207
rect 388431 270202 590673 270204
rect 388431 270146 388436 270202
rect 388492 270146 590612 270202
rect 590668 270146 590673 270202
rect 388431 270144 590673 270146
rect 388431 270141 388497 270144
rect 590607 270141 590673 270144
rect 40762 269994 40768 270058
rect 40832 270056 40838 270058
rect 41775 270056 41841 270059
rect 40832 270054 41841 270056
rect 40832 269998 41780 270054
rect 41836 269998 41841 270054
rect 40832 269996 41841 269998
rect 40832 269994 40838 269996
rect 41775 269993 41841 269996
rect 391503 270056 391569 270059
rect 597711 270056 597777 270059
rect 391503 270054 597777 270056
rect 391503 269998 391508 270054
rect 391564 269998 597716 270054
rect 597772 269998 597777 270054
rect 391503 269996 597777 269998
rect 391503 269993 391569 269996
rect 597711 269993 597777 269996
rect 139119 269908 139185 269911
rect 213327 269908 213393 269911
rect 139119 269906 213393 269908
rect 139119 269850 139124 269906
rect 139180 269850 213332 269906
rect 213388 269850 213393 269906
rect 139119 269848 213393 269850
rect 139119 269845 139185 269848
rect 213327 269845 213393 269848
rect 397071 269908 397137 269911
rect 611919 269908 611985 269911
rect 397071 269906 611985 269908
rect 397071 269850 397076 269906
rect 397132 269850 611924 269906
rect 611980 269850 611985 269906
rect 397071 269848 611985 269850
rect 397071 269845 397137 269848
rect 611919 269845 611985 269848
rect 77583 269760 77649 269763
rect 196143 269760 196209 269763
rect 77583 269758 196209 269760
rect 77583 269702 77588 269758
rect 77644 269702 196148 269758
rect 196204 269702 196209 269758
rect 77583 269700 196209 269702
rect 77583 269697 77649 269700
rect 196143 269697 196209 269700
rect 403023 269760 403089 269763
rect 626127 269760 626193 269763
rect 403023 269758 626193 269760
rect 403023 269702 403028 269758
rect 403084 269702 626132 269758
rect 626188 269702 626193 269758
rect 403023 269700 626193 269702
rect 403023 269697 403089 269700
rect 626127 269697 626193 269700
rect 42159 269612 42225 269615
rect 42682 269612 42688 269614
rect 42159 269610 42688 269612
rect 42159 269554 42164 269610
rect 42220 269554 42688 269610
rect 42159 269552 42688 269554
rect 42159 269549 42225 269552
rect 42682 269550 42688 269552
rect 42752 269550 42758 269614
rect 69423 269612 69489 269615
rect 193071 269612 193137 269615
rect 69423 269610 193137 269612
rect 69423 269554 69428 269610
rect 69484 269554 193076 269610
rect 193132 269554 193137 269610
rect 69423 269552 193137 269554
rect 69423 269549 69489 269552
rect 193071 269549 193137 269552
rect 405615 269612 405681 269615
rect 633231 269612 633297 269615
rect 405615 269610 633297 269612
rect 405615 269554 405620 269610
rect 405676 269554 633236 269610
rect 633292 269554 633297 269610
rect 405615 269552 633297 269554
rect 405615 269549 405681 269552
rect 633231 269549 633297 269552
rect 71727 269464 71793 269467
rect 194223 269464 194289 269467
rect 71727 269462 194289 269464
rect 71727 269406 71732 269462
rect 71788 269406 194228 269462
rect 194284 269406 194289 269462
rect 71727 269404 194289 269406
rect 71727 269401 71793 269404
rect 194223 269401 194289 269404
rect 410415 269464 410481 269467
rect 645039 269464 645105 269467
rect 410415 269462 645105 269464
rect 410415 269406 410420 269462
rect 410476 269406 645044 269462
rect 645100 269406 645105 269462
rect 410415 269404 645105 269406
rect 410415 269401 410481 269404
rect 645039 269401 645105 269404
rect 65871 269316 65937 269319
rect 192399 269316 192465 269319
rect 65871 269314 192465 269316
rect 65871 269258 65876 269314
rect 65932 269258 192404 269314
rect 192460 269258 192465 269314
rect 65871 269256 192465 269258
rect 65871 269253 65937 269256
rect 192399 269253 192465 269256
rect 411567 269316 411633 269319
rect 647343 269316 647409 269319
rect 411567 269314 647409 269316
rect 411567 269258 411572 269314
rect 411628 269258 647348 269314
rect 647404 269258 647409 269314
rect 411567 269256 647409 269258
rect 411567 269253 411633 269256
rect 647343 269253 647409 269256
rect 374319 269168 374385 269171
rect 555183 269168 555249 269171
rect 374319 269166 555249 269168
rect 374319 269110 374324 269166
rect 374380 269110 555188 269166
rect 555244 269110 555249 269166
rect 374319 269108 555249 269110
rect 374319 269105 374385 269108
rect 555183 269105 555249 269108
rect 368367 269020 368433 269023
rect 540975 269020 541041 269023
rect 368367 269018 541041 269020
rect 368367 268962 368372 269018
rect 368428 268962 540980 269018
rect 541036 268962 541041 269018
rect 368367 268960 541041 268962
rect 368367 268957 368433 268960
rect 540975 268957 541041 268960
rect 367887 268872 367953 268875
rect 539823 268872 539889 268875
rect 367887 268870 539889 268872
rect 367887 268814 367892 268870
rect 367948 268814 539828 268870
rect 539884 268814 539889 268870
rect 367887 268812 539889 268814
rect 367887 268809 367953 268812
rect 539823 268809 539889 268812
rect 209583 268132 209649 268135
rect 214287 268132 214353 268135
rect 209583 268130 214353 268132
rect 209583 268074 209588 268130
rect 209644 268074 214292 268130
rect 214348 268074 214353 268130
rect 209583 268072 214353 268074
rect 209583 268069 209649 268072
rect 214287 268069 214353 268072
rect 381231 267984 381297 267987
rect 388623 267984 388689 267987
rect 381231 267982 388689 267984
rect 381231 267926 381236 267982
rect 381292 267926 388628 267982
rect 388684 267926 388689 267982
rect 381231 267924 388689 267926
rect 381231 267921 381297 267924
rect 388623 267921 388689 267924
rect 61839 266948 61905 266951
rect 672399 266948 672465 266951
rect 61839 266946 672465 266948
rect 61839 266890 61844 266946
rect 61900 266890 672404 266946
rect 672460 266890 672465 266946
rect 61839 266888 672465 266890
rect 61839 266885 61905 266888
rect 672399 266885 672465 266888
rect 62031 266800 62097 266803
rect 672591 266800 672657 266803
rect 62031 266798 672657 266800
rect 62031 266742 62036 266798
rect 62092 266742 672596 266798
rect 672652 266742 672657 266798
rect 62031 266740 672657 266742
rect 62031 266737 62097 266740
rect 672591 266737 672657 266740
rect 62223 266652 62289 266655
rect 674362 266652 674368 266654
rect 62223 266650 674368 266652
rect 62223 266594 62228 266650
rect 62284 266594 674368 266650
rect 62223 266592 674368 266594
rect 62223 266589 62289 266592
rect 674362 266590 674368 266592
rect 674432 266590 674438 266654
rect 62895 266504 62961 266507
rect 674170 266504 674176 266506
rect 62895 266502 674176 266504
rect 62895 266446 62900 266502
rect 62956 266446 674176 266502
rect 62895 266444 674176 266446
rect 62895 266441 62961 266444
rect 674170 266442 674176 266444
rect 674240 266442 674246 266506
rect 44751 266356 44817 266359
rect 676282 266356 676288 266358
rect 44751 266354 676288 266356
rect 44751 266298 44756 266354
rect 44812 266298 676288 266354
rect 44751 266296 676288 266298
rect 44751 266293 44817 266296
rect 676282 266294 676288 266296
rect 676352 266294 676358 266358
rect 46287 263544 46353 263547
rect 669615 263544 669681 263547
rect 46287 263542 669681 263544
rect 46287 263486 46292 263542
rect 46348 263486 669620 263542
rect 669676 263486 669681 263542
rect 46287 263484 669681 263486
rect 46287 263481 46353 263484
rect 669615 263481 669681 263484
rect 46191 263396 46257 263399
rect 649743 263396 649809 263399
rect 46191 263394 649809 263396
rect 46191 263338 46196 263394
rect 46252 263338 649748 263394
rect 649804 263338 649809 263394
rect 46191 263336 649809 263338
rect 46191 263333 46257 263336
rect 649743 263333 649809 263336
rect 676290 262807 676350 263070
rect 676239 262802 676350 262807
rect 676239 262746 676244 262802
rect 676300 262746 676350 262802
rect 676239 262744 676350 262746
rect 676239 262741 676305 262744
rect 676047 262508 676113 262511
rect 676047 262506 676320 262508
rect 676047 262450 676052 262506
rect 676108 262450 676320 262506
rect 676047 262448 676320 262450
rect 676047 262445 676113 262448
rect 420399 262212 420465 262215
rect 412512 262210 420465 262212
rect 412512 262154 420404 262210
rect 420460 262154 420465 262210
rect 412512 262152 420465 262154
rect 420399 262149 420465 262152
rect 676290 261771 676350 262034
rect 676239 261766 676350 261771
rect 676239 261710 676244 261766
rect 676300 261710 676350 261766
rect 676239 261708 676350 261710
rect 676239 261705 676305 261708
rect 676047 261620 676113 261623
rect 676047 261618 676320 261620
rect 676047 261562 676052 261618
rect 676108 261562 676320 261618
rect 676047 261560 676320 261562
rect 676047 261557 676113 261560
rect 674554 260966 674560 261030
rect 674624 261028 674630 261030
rect 674624 260968 676320 261028
rect 674624 260966 674630 260968
rect 679695 260880 679761 260883
rect 679695 260878 679806 260880
rect 679695 260822 679700 260878
rect 679756 260822 679806 260878
rect 679695 260817 679806 260822
rect 679746 260480 679806 260817
rect 676282 260226 676288 260290
rect 676352 260226 676358 260290
rect 673978 260078 673984 260142
rect 674048 260140 674054 260142
rect 676290 260140 676350 260226
rect 674048 260110 676350 260140
rect 674048 260080 676320 260110
rect 674048 260078 674054 260080
rect 420399 259844 420465 259847
rect 679791 259844 679857 259847
rect 412512 259842 420465 259844
rect 412512 259786 420404 259842
rect 420460 259786 420465 259842
rect 412512 259784 420465 259786
rect 420399 259781 420465 259784
rect 679746 259842 679857 259844
rect 679746 259786 679796 259842
rect 679852 259786 679857 259842
rect 679746 259781 679857 259786
rect 679746 259518 679806 259781
rect 191535 259400 191601 259403
rect 191535 259398 191904 259400
rect 191535 259342 191540 259398
rect 191596 259342 191904 259398
rect 191535 259340 191904 259342
rect 191535 259337 191601 259340
rect 679746 258811 679806 259000
rect 679695 258806 679806 258811
rect 679695 258750 679700 258806
rect 679756 258750 679806 258806
rect 679695 258748 679806 258750
rect 679695 258745 679761 258748
rect 676047 258660 676113 258663
rect 676047 258658 676320 258660
rect 676047 258602 676052 258658
rect 676108 258602 676320 258658
rect 676047 258600 676320 258602
rect 676047 258597 676113 258600
rect 674938 258006 674944 258070
rect 675008 258068 675014 258070
rect 675008 258008 676320 258068
rect 675008 258006 675014 258008
rect 412482 257032 412542 257520
rect 675759 257476 675825 257479
rect 675759 257474 676320 257476
rect 675759 257418 675764 257474
rect 675820 257418 676320 257474
rect 675759 257416 676320 257418
rect 675759 257413 675825 257416
rect 675706 257044 675712 257108
rect 675776 257106 675782 257108
rect 675776 257046 676320 257106
rect 675776 257044 675782 257046
rect 420399 257032 420465 257035
rect 412482 257030 420465 257032
rect 412482 256974 420404 257030
rect 420460 256974 420465 257030
rect 412482 256972 420465 256974
rect 420399 256969 420465 256972
rect 675130 256526 675136 256590
rect 675200 256588 675206 256590
rect 675200 256528 676320 256588
rect 675200 256526 675206 256528
rect 40194 256295 40254 256410
rect 40194 256290 40305 256295
rect 40194 256234 40244 256290
rect 40300 256234 40305 256290
rect 40194 256232 40305 256234
rect 40239 256229 40305 256232
rect 41538 255703 41598 255966
rect 676866 255851 676926 255966
rect 676866 255846 676977 255851
rect 676866 255790 676916 255846
rect 676972 255790 676977 255846
rect 676866 255788 676977 255790
rect 676911 255785 676977 255788
rect 41538 255698 41649 255703
rect 41538 255642 41588 255698
rect 41644 255642 41649 255698
rect 41538 255640 41649 255642
rect 41583 255637 41649 255640
rect 676047 255626 676113 255629
rect 676047 255624 676320 255626
rect 676047 255568 676052 255624
rect 676108 255568 676320 255624
rect 676047 255566 676320 255568
rect 676047 255563 676113 255566
rect 41775 255404 41841 255407
rect 41568 255402 41841 255404
rect 41568 255346 41780 255402
rect 41836 255346 41841 255402
rect 41568 255344 41841 255346
rect 41775 255341 41841 255344
rect 420399 255256 420465 255259
rect 412512 255254 420465 255256
rect 412512 255198 420404 255254
rect 420460 255198 420465 255254
rect 412512 255196 420465 255198
rect 420399 255193 420465 255196
rect 675951 255108 676017 255111
rect 675951 255106 676320 255108
rect 675951 255050 675956 255106
rect 676012 255050 676320 255106
rect 675951 255048 676320 255050
rect 675951 255045 676017 255048
rect 41775 254960 41841 254963
rect 41568 254958 41841 254960
rect 41568 254902 41780 254958
rect 41836 254902 41841 254958
rect 41568 254900 41841 254902
rect 41775 254897 41841 254900
rect 41775 254516 41841 254519
rect 41568 254514 41841 254516
rect 41568 254458 41780 254514
rect 41836 254458 41841 254514
rect 41568 254456 41841 254458
rect 41775 254453 41841 254456
rect 676290 254371 676350 254486
rect 676239 254366 676350 254371
rect 676239 254310 676244 254366
rect 676300 254310 676350 254366
rect 676239 254308 676350 254310
rect 676239 254305 676305 254308
rect 23151 254220 23217 254223
rect 23106 254218 23217 254220
rect 23106 254162 23156 254218
rect 23212 254162 23217 254218
rect 23106 254157 23217 254162
rect 23106 253894 23166 254157
rect 676866 253927 676926 254042
rect 676815 253922 676926 253927
rect 676815 253866 676820 253922
rect 676876 253866 676926 253922
rect 676815 253864 676926 253866
rect 676815 253861 676881 253864
rect 675898 253566 675904 253630
rect 675968 253628 675974 253630
rect 675968 253568 676320 253628
rect 675968 253566 675974 253568
rect 23298 253335 23358 253450
rect 23055 253332 23121 253335
rect 23055 253330 23166 253332
rect 23055 253274 23060 253330
rect 23116 253274 23166 253330
rect 23055 253269 23166 253274
rect 23298 253330 23409 253335
rect 23298 253274 23348 253330
rect 23404 253274 23409 253330
rect 23298 253272 23409 253274
rect 23343 253269 23409 253272
rect 23106 252932 23166 253269
rect 676047 253036 676113 253039
rect 676047 253034 676320 253036
rect 676047 252978 676052 253034
rect 676108 252978 676320 253034
rect 676047 252976 676320 252978
rect 676047 252973 676113 252976
rect 420399 252888 420465 252891
rect 412512 252886 420465 252888
rect 412512 252830 420404 252886
rect 420460 252830 420465 252886
rect 412512 252828 420465 252830
rect 420399 252825 420465 252828
rect 23247 252740 23313 252743
rect 23247 252738 23358 252740
rect 23247 252682 23252 252738
rect 23308 252682 23358 252738
rect 23247 252677 23358 252682
rect 23298 252414 23358 252677
rect 676290 252447 676350 252562
rect 676239 252442 676350 252447
rect 676239 252386 676244 252442
rect 676300 252386 676350 252442
rect 676239 252384 676350 252386
rect 676239 252381 676305 252384
rect 675951 252074 676017 252077
rect 675951 252072 676320 252074
rect 675951 252016 675956 252072
rect 676012 252016 676320 252072
rect 675951 252014 676320 252016
rect 675951 252011 676017 252014
rect 40578 251706 40638 251970
rect 40570 251642 40576 251706
rect 40640 251642 40646 251706
rect 190191 251704 190257 251707
rect 679983 251704 680049 251707
rect 190191 251702 191904 251704
rect 190191 251646 190196 251702
rect 190252 251646 191904 251702
rect 190191 251644 191904 251646
rect 679938 251702 680049 251704
rect 679938 251646 679988 251702
rect 680044 251646 680049 251702
rect 190191 251641 190257 251644
rect 679938 251641 680049 251646
rect 679938 251526 679998 251641
rect 42106 251408 42112 251410
rect 41568 251348 42112 251408
rect 42106 251346 42112 251348
rect 42176 251346 42182 251410
rect 42682 250964 42688 250966
rect 41568 250904 42688 250964
rect 42682 250902 42688 250904
rect 42752 250902 42758 250966
rect 679746 250819 679806 251082
rect 679746 250814 679857 250819
rect 679983 250816 680049 250819
rect 679746 250758 679796 250814
rect 679852 250758 679857 250814
rect 679746 250756 679857 250758
rect 679791 250753 679857 250756
rect 679938 250814 680049 250816
rect 679938 250758 679988 250814
rect 680044 250758 680049 250814
rect 679938 250753 680049 250758
rect 679938 250564 679998 250753
rect 420303 250520 420369 250523
rect 412512 250518 420369 250520
rect 41346 250226 41406 250490
rect 412512 250462 420308 250518
rect 420364 250462 420369 250518
rect 412512 250460 420369 250462
rect 420303 250457 420369 250460
rect 679791 250372 679857 250375
rect 679746 250370 679857 250372
rect 679746 250314 679796 250370
rect 679852 250314 679857 250370
rect 679746 250309 679857 250314
rect 41338 250162 41344 250226
rect 41408 250162 41414 250226
rect 679746 250046 679806 250309
rect 42874 249928 42880 249930
rect 41568 249868 42880 249928
rect 42874 249866 42880 249868
rect 42944 249866 42950 249930
rect 41538 249188 41598 249454
rect 674746 249274 674752 249338
rect 674816 249336 674822 249338
rect 679695 249336 679761 249339
rect 674816 249334 679761 249336
rect 674816 249278 679700 249334
rect 679756 249278 679761 249334
rect 674816 249276 679761 249278
rect 674816 249274 674822 249276
rect 679695 249273 679761 249276
rect 41679 249188 41745 249191
rect 41538 249186 41745 249188
rect 41538 249130 41684 249186
rect 41740 249130 41745 249186
rect 41538 249128 41745 249130
rect 41679 249125 41745 249128
rect 40770 248746 40830 249010
rect 40762 248682 40768 248746
rect 40832 248682 40838 248746
rect 41154 248154 41214 248418
rect 41146 248090 41152 248154
rect 41216 248090 41222 248154
rect 420399 248152 420465 248155
rect 412512 248150 420465 248152
rect 412512 248094 420404 248150
rect 420460 248094 420465 248150
rect 412512 248092 420465 248094
rect 420399 248089 420465 248092
rect 676666 247942 676672 248006
rect 676736 248004 676742 248006
rect 676911 248004 676977 248007
rect 676736 248002 676977 248004
rect 676736 247946 676916 248002
rect 676972 247946 676977 248002
rect 676736 247944 676977 247946
rect 676736 247942 676742 247944
rect 676911 247941 676977 247944
rect 40962 247710 41022 247900
rect 676474 247794 676480 247858
rect 676544 247856 676550 247858
rect 676815 247856 676881 247859
rect 676544 247854 676881 247856
rect 676544 247798 676820 247854
rect 676876 247798 676881 247854
rect 676544 247796 676881 247798
rect 676544 247794 676550 247796
rect 676815 247793 676881 247796
rect 40954 247646 40960 247710
rect 41024 247646 41030 247710
rect 41914 247560 41920 247562
rect 41568 247500 41920 247560
rect 41914 247498 41920 247500
rect 41984 247498 41990 247562
rect 42490 246968 42496 246970
rect 41568 246908 42496 246968
rect 42490 246906 42496 246908
rect 42560 246906 42566 246970
rect 41538 246230 41598 246346
rect 41530 246166 41536 246230
rect 41600 246166 41606 246230
rect 42298 246080 42304 246082
rect 41568 246020 42304 246080
rect 42298 246018 42304 246020
rect 42368 246018 42374 246082
rect 41722 245488 41728 245490
rect 41568 245428 41728 245488
rect 41722 245426 41728 245428
rect 41792 245426 41798 245490
rect 412482 245340 412542 245828
rect 420399 245340 420465 245343
rect 412482 245338 420465 245340
rect 412482 245282 420404 245338
rect 420460 245282 420465 245338
rect 412482 245280 420465 245282
rect 420399 245277 420465 245280
rect 41775 244896 41841 244899
rect 41568 244894 41841 244896
rect 41568 244838 41780 244894
rect 41836 244838 41841 244894
rect 41568 244836 41841 244838
rect 41775 244833 41841 244836
rect 41583 244748 41649 244751
rect 41538 244746 41649 244748
rect 41538 244690 41588 244746
rect 41644 244690 41649 244746
rect 41538 244685 41649 244690
rect 41538 244496 41598 244685
rect 148335 244600 148401 244603
rect 143904 244598 148401 244600
rect 143904 244542 148340 244598
rect 148396 244542 148401 244598
rect 143904 244540 148401 244542
rect 148335 244537 148401 244540
rect 41538 243715 41598 243978
rect 41538 243710 41649 243715
rect 41538 243654 41588 243710
rect 41644 243654 41649 243710
rect 41538 243652 41649 243654
rect 41583 243649 41649 243652
rect 148719 243416 148785 243419
rect 143904 243414 148785 243416
rect 143904 243358 148724 243414
rect 148780 243358 148785 243414
rect 143904 243356 148785 243358
rect 148719 243353 148785 243356
rect 187119 243416 187185 243419
rect 191874 243416 191934 243904
rect 675663 243714 675729 243715
rect 675663 243710 675712 243714
rect 675776 243712 675782 243714
rect 675663 243654 675668 243710
rect 675663 243650 675712 243654
rect 675776 243652 675820 243712
rect 675776 243650 675782 243652
rect 675663 243649 675729 243650
rect 420399 243564 420465 243567
rect 412512 243562 420465 243564
rect 412512 243506 420404 243562
rect 420460 243506 420465 243562
rect 412512 243504 420465 243506
rect 420399 243501 420465 243504
rect 187119 243414 191934 243416
rect 187119 243358 187124 243414
rect 187180 243358 191934 243414
rect 187119 243356 191934 243358
rect 187119 243353 187185 243356
rect 143874 242084 143934 242128
rect 148527 242084 148593 242087
rect 143874 242082 148593 242084
rect 143874 242026 148532 242082
rect 148588 242026 148593 242082
rect 143874 242024 148593 242026
rect 148527 242021 148593 242024
rect 420399 241196 420465 241199
rect 412512 241194 420465 241196
rect 412512 241138 420404 241194
rect 420460 241138 420465 241194
rect 412512 241136 420465 241138
rect 420399 241133 420465 241136
rect 148911 240900 148977 240903
rect 143904 240898 148977 240900
rect 143904 240842 148916 240898
rect 148972 240842 148977 240898
rect 143904 240840 148977 240842
rect 148911 240837 148977 240840
rect 412143 240160 412209 240163
rect 627183 240160 627249 240163
rect 412143 240158 627249 240160
rect 412143 240102 412148 240158
rect 412204 240102 627188 240158
rect 627244 240102 627249 240158
rect 412143 240100 627249 240102
rect 412143 240097 412209 240100
rect 627183 240097 627249 240100
rect 412047 240012 412113 240015
rect 567375 240012 567441 240015
rect 412047 240010 567441 240012
rect 412047 239954 412052 240010
rect 412108 239954 567380 240010
rect 567436 239954 567441 240010
rect 412047 239952 567441 239954
rect 412047 239949 412113 239952
rect 567375 239949 567441 239952
rect 148239 239716 148305 239719
rect 143904 239714 148305 239716
rect 143904 239658 148244 239714
rect 148300 239658 148305 239714
rect 143904 239656 148305 239658
rect 148239 239653 148305 239656
rect 675130 239062 675136 239126
rect 675200 239124 675206 239126
rect 675375 239124 675441 239127
rect 675200 239122 675441 239124
rect 675200 239066 675380 239122
rect 675436 239066 675441 239122
rect 675200 239064 675441 239066
rect 675200 239062 675206 239064
rect 675375 239061 675441 239064
rect 413391 238976 413457 238979
rect 555375 238976 555441 238979
rect 413391 238974 555441 238976
rect 413391 238918 413396 238974
rect 413452 238918 555380 238974
rect 555436 238918 555441 238974
rect 413391 238916 555441 238918
rect 413391 238913 413457 238916
rect 555375 238913 555441 238916
rect 414063 238828 414129 238831
rect 581775 238828 581841 238831
rect 414063 238826 581841 238828
rect 414063 238770 414068 238826
rect 414124 238770 581780 238826
rect 581836 238770 581841 238826
rect 414063 238768 581841 238770
rect 414063 238765 414129 238768
rect 581775 238765 581841 238768
rect 42063 238682 42129 238683
rect 42063 238678 42112 238682
rect 42176 238680 42182 238682
rect 413679 238680 413745 238683
rect 550191 238680 550257 238683
rect 42063 238622 42068 238678
rect 42063 238618 42112 238622
rect 42176 238620 42220 238680
rect 413679 238678 550257 238680
rect 413679 238622 413684 238678
rect 413740 238622 550196 238678
rect 550252 238622 550257 238678
rect 413679 238620 550257 238622
rect 42176 238618 42182 238620
rect 42063 238617 42129 238618
rect 413679 238617 413745 238620
rect 550191 238617 550257 238620
rect 42106 238470 42112 238534
rect 42176 238532 42182 238534
rect 42682 238532 42688 238534
rect 42176 238472 42688 238532
rect 42176 238470 42182 238472
rect 42682 238470 42688 238472
rect 42752 238470 42758 238534
rect 148431 238532 148497 238535
rect 143904 238530 148497 238532
rect 143904 238474 148436 238530
rect 148492 238474 148497 238530
rect 143904 238472 148497 238474
rect 148431 238469 148497 238472
rect 413967 238384 414033 238387
rect 544335 238384 544401 238387
rect 413967 238382 544401 238384
rect 413967 238326 413972 238382
rect 414028 238326 544340 238382
rect 544396 238326 544401 238382
rect 413967 238324 544401 238326
rect 413967 238321 414033 238324
rect 544335 238321 544401 238324
rect 415215 238236 415281 238239
rect 559887 238236 559953 238239
rect 415215 238234 559953 238236
rect 415215 238178 415220 238234
rect 415276 238178 559892 238234
rect 559948 238178 559953 238234
rect 415215 238176 559953 238178
rect 415215 238173 415281 238176
rect 559887 238173 559953 238176
rect 414447 238088 414513 238091
rect 537999 238088 538065 238091
rect 414447 238086 538065 238088
rect 414447 238030 414452 238086
rect 414508 238030 538004 238086
rect 538060 238030 538065 238086
rect 414447 238028 538065 238030
rect 414447 238025 414513 238028
rect 537999 238025 538065 238028
rect 675759 238088 675825 238091
rect 675898 238088 675904 238090
rect 675759 238086 675904 238088
rect 675759 238030 675764 238086
rect 675820 238030 675904 238086
rect 675759 238028 675904 238030
rect 675759 238025 675825 238028
rect 675898 238026 675904 238028
rect 675968 238026 675974 238090
rect 41871 236906 41937 236907
rect 41871 236902 41920 236906
rect 41984 236904 41990 236906
rect 41871 236846 41876 236902
rect 41871 236842 41920 236846
rect 41984 236844 42028 236904
rect 41984 236842 41990 236844
rect 41871 236841 41937 236842
rect 40570 236694 40576 236758
rect 40640 236756 40646 236758
rect 41914 236756 41920 236758
rect 40640 236696 41920 236756
rect 40640 236694 40646 236696
rect 41914 236694 41920 236696
rect 41984 236694 41990 236758
rect 143874 236756 143934 237244
rect 372207 237052 372273 237055
rect 396975 237052 397041 237055
rect 372207 237050 397041 237052
rect 372207 236994 372212 237050
rect 372268 236994 396980 237050
rect 397036 236994 397041 237050
rect 372207 236992 397041 236994
rect 372207 236989 372273 236992
rect 396975 236989 397041 236992
rect 397114 236990 397120 237054
rect 397184 237052 397190 237054
rect 397498 237052 397504 237054
rect 397184 236992 397504 237052
rect 397184 236990 397190 236992
rect 397498 236990 397504 236992
rect 397568 236990 397574 237054
rect 397647 237052 397713 237055
rect 573135 237052 573201 237055
rect 397647 237050 573201 237052
rect 397647 236994 397652 237050
rect 397708 236994 573140 237050
rect 573196 236994 573201 237050
rect 397647 236992 573201 236994
rect 397647 236989 397713 236992
rect 573135 236989 573201 236992
rect 373455 236904 373521 236907
rect 387375 236904 387441 236907
rect 373455 236902 387441 236904
rect 373455 236846 373460 236902
rect 373516 236846 387380 236902
rect 387436 236846 387441 236902
rect 373455 236844 387441 236846
rect 373455 236841 373521 236844
rect 387375 236841 387441 236844
rect 387567 236904 387633 236907
rect 397071 236904 397137 236907
rect 398031 236904 398097 236907
rect 387567 236902 397137 236904
rect 387567 236846 387572 236902
rect 387628 236846 397076 236902
rect 397132 236846 397137 236902
rect 387567 236844 397137 236846
rect 387567 236841 387633 236844
rect 397071 236841 397137 236844
rect 397410 236902 398097 236904
rect 397410 236846 398036 236902
rect 398092 236846 398097 236902
rect 397410 236844 398097 236846
rect 148623 236756 148689 236759
rect 143874 236754 148689 236756
rect 143874 236698 148628 236754
rect 148684 236698 148689 236754
rect 143874 236696 148689 236698
rect 148623 236693 148689 236696
rect 370383 236756 370449 236759
rect 397410 236756 397470 236844
rect 398031 236841 398097 236844
rect 398319 236904 398385 236907
rect 567471 236904 567537 236907
rect 398319 236902 567537 236904
rect 398319 236846 398324 236902
rect 398380 236846 567476 236902
rect 567532 236846 567537 236902
rect 398319 236844 567537 236846
rect 398319 236841 398385 236844
rect 567471 236841 567537 236844
rect 370383 236754 397470 236756
rect 370383 236698 370388 236754
rect 370444 236698 397470 236754
rect 370383 236696 397470 236698
rect 370383 236693 370449 236696
rect 397690 236694 397696 236758
rect 397760 236756 397766 236758
rect 407290 236756 407296 236758
rect 397760 236696 407296 236756
rect 397760 236694 397766 236696
rect 407290 236694 407296 236696
rect 407360 236694 407366 236758
rect 407439 236756 407505 236759
rect 565263 236756 565329 236759
rect 407439 236754 565329 236756
rect 407439 236698 407444 236754
rect 407500 236698 565268 236754
rect 565324 236698 565329 236754
rect 407439 236696 565329 236698
rect 407439 236693 407505 236696
rect 565263 236693 565329 236696
rect 377967 236608 378033 236611
rect 559215 236608 559281 236611
rect 377967 236606 559281 236608
rect 377967 236550 377972 236606
rect 378028 236550 559220 236606
rect 559276 236550 559281 236606
rect 377967 236548 559281 236550
rect 377967 236545 378033 236548
rect 559215 236545 559281 236548
rect 368943 236460 369009 236463
rect 387375 236460 387441 236463
rect 557679 236460 557745 236463
rect 368943 236458 387198 236460
rect 368943 236402 368948 236458
rect 369004 236402 387198 236458
rect 368943 236400 387198 236402
rect 368943 236397 369009 236400
rect 374895 236312 374961 236315
rect 377967 236312 378033 236315
rect 374895 236310 378033 236312
rect 374895 236254 374900 236310
rect 374956 236254 377972 236310
rect 378028 236254 378033 236310
rect 374895 236252 378033 236254
rect 374895 236249 374961 236252
rect 377967 236249 378033 236252
rect 378159 236312 378225 236315
rect 382383 236312 382449 236315
rect 378159 236310 382449 236312
rect 378159 236254 378164 236310
rect 378220 236254 382388 236310
rect 382444 236254 382449 236310
rect 378159 236252 382449 236254
rect 378159 236249 378225 236252
rect 382383 236249 382449 236252
rect 382575 236312 382641 236315
rect 386991 236312 387057 236315
rect 382575 236310 387057 236312
rect 382575 236254 382580 236310
rect 382636 236254 386996 236310
rect 387052 236254 387057 236310
rect 382575 236252 387057 236254
rect 387138 236312 387198 236400
rect 387375 236458 557745 236460
rect 387375 236402 387380 236458
rect 387436 236402 557684 236458
rect 557740 236402 557745 236458
rect 387375 236400 557745 236402
rect 387375 236397 387441 236400
rect 557679 236397 557745 236400
rect 397114 236312 397120 236314
rect 387138 236252 397120 236312
rect 382575 236249 382641 236252
rect 386991 236249 387057 236252
rect 397114 236250 397120 236252
rect 397184 236250 397190 236314
rect 397359 236312 397425 236315
rect 407439 236312 407505 236315
rect 397359 236310 407505 236312
rect 397359 236254 397364 236310
rect 397420 236254 407444 236310
rect 407500 236254 407505 236310
rect 397359 236252 407505 236254
rect 397359 236249 397425 236252
rect 407439 236249 407505 236252
rect 407674 236250 407680 236314
rect 407744 236312 407750 236314
rect 413679 236312 413745 236315
rect 415215 236312 415281 236315
rect 407744 236310 413745 236312
rect 407744 236254 413684 236310
rect 413740 236254 413745 236310
rect 407744 236252 413745 236254
rect 407744 236250 407750 236252
rect 413679 236249 413745 236252
rect 413826 236310 415281 236312
rect 413826 236254 415220 236310
rect 415276 236254 415281 236310
rect 413826 236252 415281 236254
rect 413826 236167 413886 236252
rect 415215 236249 415281 236252
rect 415407 236312 415473 236315
rect 621135 236312 621201 236315
rect 415407 236310 621201 236312
rect 415407 236254 415412 236310
rect 415468 236254 621140 236310
rect 621196 236254 621201 236310
rect 415407 236252 621201 236254
rect 415407 236249 415473 236252
rect 621135 236249 621201 236252
rect 356847 236164 356913 236167
rect 406479 236164 406545 236167
rect 356847 236162 406545 236164
rect 356847 236106 356852 236162
rect 356908 236106 406484 236162
rect 406540 236106 406545 236162
rect 356847 236104 406545 236106
rect 356847 236101 356913 236104
rect 406479 236101 406545 236104
rect 409935 236164 410001 236167
rect 413626 236164 413632 236166
rect 409935 236162 413632 236164
rect 409935 236106 409940 236162
rect 409996 236106 413632 236162
rect 409935 236104 413632 236106
rect 409935 236101 410001 236104
rect 413626 236102 413632 236104
rect 413696 236102 413702 236166
rect 413826 236162 413937 236167
rect 413826 236106 413876 236162
rect 413932 236106 413937 236162
rect 413826 236104 413937 236106
rect 413871 236101 413937 236104
rect 414010 236102 414016 236166
rect 414080 236164 414086 236166
rect 591471 236164 591537 236167
rect 414080 236162 591537 236164
rect 414080 236106 591476 236162
rect 591532 236106 591537 236162
rect 414080 236104 591537 236106
rect 414080 236102 414086 236104
rect 591471 236101 591537 236104
rect 146991 236016 147057 236019
rect 143904 236014 147057 236016
rect 143904 235958 146996 236014
rect 147052 235958 147057 236014
rect 143904 235956 147057 235958
rect 146991 235953 147057 235956
rect 385839 236016 385905 236019
rect 580335 236016 580401 236019
rect 385839 236014 580401 236016
rect 385839 235958 385844 236014
rect 385900 235958 580340 236014
rect 580396 235958 580401 236014
rect 385839 235956 580401 235958
rect 385839 235953 385905 235956
rect 580335 235953 580401 235956
rect 675759 236016 675825 236019
rect 676474 236016 676480 236018
rect 675759 236014 676480 236016
rect 675759 235958 675764 236014
rect 675820 235958 676480 236014
rect 675759 235956 676480 235958
rect 675759 235953 675825 235956
rect 676474 235954 676480 235956
rect 676544 235954 676550 236018
rect 389871 235868 389937 235871
rect 587919 235868 587985 235871
rect 389871 235866 587985 235868
rect 389871 235810 389876 235866
rect 389932 235810 587924 235866
rect 587980 235810 587985 235866
rect 389871 235808 587985 235810
rect 389871 235805 389937 235808
rect 587919 235805 587985 235808
rect 342543 235720 342609 235723
rect 390735 235720 390801 235723
rect 342543 235718 390801 235720
rect 342543 235662 342548 235718
rect 342604 235662 390740 235718
rect 390796 235662 390801 235718
rect 342543 235660 390801 235662
rect 342543 235657 342609 235660
rect 390735 235657 390801 235660
rect 393039 235720 393105 235723
rect 590703 235720 590769 235723
rect 393039 235718 590769 235720
rect 393039 235662 393044 235718
rect 393100 235662 590708 235718
rect 590764 235662 590769 235718
rect 393039 235660 590769 235662
rect 393039 235657 393105 235660
rect 590703 235657 590769 235660
rect 41775 235574 41841 235575
rect 41722 235572 41728 235574
rect 41684 235512 41728 235572
rect 41792 235570 41841 235574
rect 41836 235514 41841 235570
rect 41722 235510 41728 235512
rect 41792 235510 41841 235514
rect 41775 235509 41841 235510
rect 367215 235572 367281 235575
rect 397743 235572 397809 235575
rect 367215 235570 397809 235572
rect 367215 235514 367220 235570
rect 367276 235514 397748 235570
rect 397804 235514 397809 235570
rect 367215 235512 397809 235514
rect 367215 235509 367281 235512
rect 397743 235509 397809 235512
rect 399855 235572 399921 235575
rect 608271 235572 608337 235575
rect 399855 235570 608337 235572
rect 399855 235514 399860 235570
rect 399916 235514 608276 235570
rect 608332 235514 608337 235570
rect 399855 235512 608337 235514
rect 399855 235509 399921 235512
rect 608271 235509 608337 235512
rect 401391 235424 401457 235427
rect 611247 235424 611313 235427
rect 401391 235422 611313 235424
rect 401391 235366 401396 235422
rect 401452 235366 611252 235422
rect 611308 235366 611313 235422
rect 401391 235364 611313 235366
rect 401391 235361 401457 235364
rect 611247 235361 611313 235364
rect 402639 235276 402705 235279
rect 614319 235276 614385 235279
rect 402639 235274 614385 235276
rect 402639 235218 402644 235274
rect 402700 235218 614324 235274
rect 614380 235218 614385 235274
rect 402639 235216 614385 235218
rect 402639 235213 402705 235216
rect 614319 235213 614385 235216
rect 405423 235128 405489 235131
rect 618831 235128 618897 235131
rect 405423 235126 618897 235128
rect 405423 235070 405428 235126
rect 405484 235070 618836 235126
rect 618892 235070 618897 235126
rect 405423 235068 618897 235070
rect 405423 235065 405489 235068
rect 618831 235065 618897 235068
rect 299439 234980 299505 234983
rect 354639 234980 354705 234983
rect 299439 234978 354705 234980
rect 299439 234922 299444 234978
rect 299500 234922 354644 234978
rect 354700 234922 354705 234978
rect 299439 234920 354705 234922
rect 299439 234917 299505 234920
rect 354639 234917 354705 234920
rect 356751 234980 356817 234983
rect 403119 234980 403185 234983
rect 356751 234978 403185 234980
rect 356751 234922 356756 234978
rect 356812 234922 403124 234978
rect 403180 234922 403185 234978
rect 356751 234920 403185 234922
rect 356751 234917 356817 234920
rect 403119 234917 403185 234920
rect 403983 234980 404049 234983
rect 616623 234980 616689 234983
rect 403983 234978 616689 234980
rect 403983 234922 403988 234978
rect 404044 234922 616628 234978
rect 616684 234922 616689 234978
rect 403983 234920 616689 234922
rect 403983 234917 404049 234920
rect 616623 234917 616689 234920
rect 42159 234832 42225 234835
rect 42490 234832 42496 234834
rect 42159 234830 42496 234832
rect 42159 234774 42164 234830
rect 42220 234774 42496 234830
rect 42159 234772 42496 234774
rect 42159 234769 42225 234772
rect 42490 234770 42496 234772
rect 42560 234770 42566 234834
rect 148815 234832 148881 234835
rect 143904 234830 148881 234832
rect 143904 234774 148820 234830
rect 148876 234774 148881 234830
rect 143904 234772 148881 234774
rect 148815 234769 148881 234772
rect 347631 234832 347697 234835
rect 405327 234832 405393 234835
rect 347631 234830 405393 234832
rect 347631 234774 347636 234830
rect 347692 234774 405332 234830
rect 405388 234774 405393 234830
rect 347631 234772 405393 234774
rect 347631 234769 347697 234772
rect 405327 234769 405393 234772
rect 405519 234832 405585 234835
rect 619599 234832 619665 234835
rect 405519 234830 619665 234832
rect 405519 234774 405524 234830
rect 405580 234774 619604 234830
rect 619660 234774 619665 234830
rect 405519 234772 619665 234774
rect 405519 234769 405585 234772
rect 619599 234769 619665 234772
rect 299343 234684 299409 234687
rect 405999 234684 406065 234687
rect 299343 234682 406065 234684
rect 299343 234626 299348 234682
rect 299404 234626 406004 234682
rect 406060 234626 406065 234682
rect 299343 234624 406065 234626
rect 299343 234621 299409 234624
rect 405999 234621 406065 234624
rect 408495 234684 408561 234687
rect 625551 234684 625617 234687
rect 408495 234682 625617 234684
rect 408495 234626 408500 234682
rect 408556 234626 625556 234682
rect 625612 234626 625617 234682
rect 408495 234624 625617 234626
rect 408495 234621 408561 234624
rect 625551 234621 625617 234624
rect 379119 234536 379185 234539
rect 409839 234536 409905 234539
rect 379119 234534 409905 234536
rect 379119 234478 379124 234534
rect 379180 234478 409844 234534
rect 409900 234478 409905 234534
rect 379119 234476 409905 234478
rect 379119 234473 379185 234476
rect 409839 234473 409905 234476
rect 411375 234536 411441 234539
rect 590895 234536 590961 234539
rect 411375 234534 590961 234536
rect 411375 234478 411380 234534
rect 411436 234478 590900 234534
rect 590956 234478 590961 234534
rect 411375 234476 590961 234478
rect 411375 234473 411441 234476
rect 590895 234473 590961 234476
rect 674938 234474 674944 234538
rect 675008 234536 675014 234538
rect 675375 234536 675441 234539
rect 675008 234534 675441 234536
rect 675008 234478 675380 234534
rect 675436 234478 675441 234534
rect 675008 234476 675441 234478
rect 675008 234474 675014 234476
rect 675375 234473 675441 234476
rect 42159 234388 42225 234391
rect 42298 234388 42304 234390
rect 42159 234386 42304 234388
rect 42159 234330 42164 234386
rect 42220 234330 42304 234386
rect 42159 234328 42304 234330
rect 42159 234325 42225 234328
rect 42298 234326 42304 234328
rect 42368 234326 42374 234390
rect 382095 234388 382161 234391
rect 410031 234388 410097 234391
rect 382095 234386 410097 234388
rect 382095 234330 382100 234386
rect 382156 234330 410036 234386
rect 410092 234330 410097 234386
rect 382095 234328 410097 234330
rect 382095 234325 382161 234328
rect 410031 234325 410097 234328
rect 410799 234388 410865 234391
rect 587439 234388 587505 234391
rect 410799 234386 587505 234388
rect 410799 234330 410804 234386
rect 410860 234330 587444 234386
rect 587500 234330 587505 234386
rect 410799 234328 587505 234330
rect 410799 234325 410865 234328
rect 587439 234325 587505 234328
rect 341583 234240 341649 234243
rect 490479 234240 490545 234243
rect 341583 234238 490545 234240
rect 341583 234182 341588 234238
rect 341644 234182 490484 234238
rect 490540 234182 490545 234238
rect 341583 234180 490545 234182
rect 341583 234177 341649 234180
rect 490479 234177 490545 234180
rect 332559 234092 332625 234095
rect 472335 234092 472401 234095
rect 332559 234090 472401 234092
rect 332559 234034 332564 234090
rect 332620 234034 472340 234090
rect 472396 234034 472401 234090
rect 332559 234032 472401 234034
rect 332559 234029 332625 234032
rect 472335 234029 472401 234032
rect 400239 233944 400305 233947
rect 480879 233944 480945 233947
rect 400239 233942 480945 233944
rect 400239 233886 400244 233942
rect 400300 233886 480884 233942
rect 480940 233886 480945 233942
rect 400239 233884 480945 233886
rect 400239 233881 400305 233884
rect 480879 233881 480945 233884
rect 364047 233796 364113 233799
rect 405903 233796 405969 233799
rect 364047 233794 405969 233796
rect 364047 233738 364052 233794
rect 364108 233738 405908 233794
rect 405964 233738 405969 233794
rect 364047 233736 405969 233738
rect 364047 233733 364113 233736
rect 405903 233733 405969 233736
rect 42159 233648 42225 233651
rect 42874 233648 42880 233650
rect 42159 233646 42880 233648
rect 42159 233590 42164 233646
rect 42220 233590 42880 233646
rect 42159 233588 42880 233590
rect 42159 233585 42225 233588
rect 42874 233586 42880 233588
rect 42944 233586 42950 233650
rect 149007 233648 149073 233651
rect 143904 233646 149073 233648
rect 143904 233590 149012 233646
rect 149068 233590 149073 233646
rect 143904 233588 149073 233590
rect 149007 233585 149073 233588
rect 365679 233352 365745 233355
rect 380079 233352 380145 233355
rect 365679 233350 380145 233352
rect 365679 233294 365684 233350
rect 365740 233294 380084 233350
rect 380140 233294 380145 233350
rect 365679 233292 380145 233294
rect 365679 233289 365745 233292
rect 380079 233289 380145 233292
rect 343983 233204 344049 233207
rect 495087 233204 495153 233207
rect 343983 233202 495153 233204
rect 343983 233146 343988 233202
rect 344044 233146 495092 233202
rect 495148 233146 495153 233202
rect 343983 233144 495153 233146
rect 343983 233141 344049 233144
rect 495087 233141 495153 233144
rect 371151 233056 371217 233059
rect 549423 233056 549489 233059
rect 371151 233054 549489 233056
rect 371151 232998 371156 233054
rect 371212 232998 549428 233054
rect 549484 232998 549489 233054
rect 371151 232996 549489 232998
rect 371151 232993 371217 232996
rect 549423 232993 549489 232996
rect 370767 232908 370833 232911
rect 551631 232908 551697 232911
rect 370767 232906 551697 232908
rect 370767 232850 370772 232906
rect 370828 232850 551636 232906
rect 551692 232850 551697 232906
rect 370767 232848 551697 232850
rect 370767 232845 370833 232848
rect 551631 232845 551697 232848
rect 374031 232760 374097 232763
rect 557583 232760 557649 232763
rect 374031 232758 557649 232760
rect 374031 232702 374036 232758
rect 374092 232702 557588 232758
rect 557644 232702 557649 232758
rect 374031 232700 557649 232702
rect 374031 232697 374097 232700
rect 557583 232697 557649 232700
rect 375375 232612 375441 232615
rect 560751 232612 560817 232615
rect 375375 232610 560817 232612
rect 375375 232554 375380 232610
rect 375436 232554 560756 232610
rect 560812 232554 560817 232610
rect 375375 232552 560817 232554
rect 375375 232549 375441 232552
rect 560751 232549 560817 232552
rect 675759 232612 675825 232615
rect 676666 232612 676672 232614
rect 675759 232610 676672 232612
rect 675759 232554 675764 232610
rect 675820 232554 676672 232610
rect 675759 232552 676672 232554
rect 675759 232549 675825 232552
rect 676666 232550 676672 232552
rect 676736 232550 676742 232614
rect 381711 232464 381777 232467
rect 570447 232464 570513 232467
rect 381711 232462 570513 232464
rect 381711 232406 381716 232462
rect 381772 232406 570452 232462
rect 570508 232406 570513 232462
rect 381711 232404 570513 232406
rect 381711 232401 381777 232404
rect 570447 232401 570513 232404
rect 149103 232316 149169 232319
rect 143904 232314 149169 232316
rect 143904 232258 149108 232314
rect 149164 232258 149169 232314
rect 143904 232256 149169 232258
rect 149103 232253 149169 232256
rect 384975 232316 385041 232319
rect 576591 232316 576657 232319
rect 384975 232314 576657 232316
rect 384975 232258 384980 232314
rect 385036 232258 576596 232314
rect 576652 232258 576657 232314
rect 384975 232256 576657 232258
rect 384975 232253 385041 232256
rect 576591 232253 576657 232256
rect 385263 232168 385329 232171
rect 578031 232168 578097 232171
rect 385263 232166 578097 232168
rect 385263 232110 385268 232166
rect 385324 232110 578036 232166
rect 578092 232110 578097 232166
rect 385263 232108 578097 232110
rect 385263 232105 385329 232108
rect 578031 232105 578097 232108
rect 382671 232020 382737 232023
rect 575823 232020 575889 232023
rect 382671 232018 575889 232020
rect 382671 231962 382676 232018
rect 382732 231962 575828 232018
rect 575884 231962 575889 232018
rect 382671 231960 575889 231962
rect 382671 231957 382737 231960
rect 575823 231957 575889 231960
rect 333807 231872 333873 231875
rect 368655 231872 368721 231875
rect 333807 231870 368721 231872
rect 333807 231814 333812 231870
rect 333868 231814 368660 231870
rect 368716 231814 368721 231870
rect 333807 231812 368721 231814
rect 333807 231809 333873 231812
rect 368655 231809 368721 231812
rect 405807 231872 405873 231875
rect 604527 231872 604593 231875
rect 405807 231870 604593 231872
rect 405807 231814 405812 231870
rect 405868 231814 604532 231870
rect 604588 231814 604593 231870
rect 405807 231812 604593 231814
rect 405807 231809 405873 231812
rect 604527 231809 604593 231812
rect 330255 231724 330321 231727
rect 470127 231724 470193 231727
rect 330255 231722 470193 231724
rect 330255 231666 330260 231722
rect 330316 231666 470132 231722
rect 470188 231666 470193 231722
rect 330255 231664 470193 231666
rect 330255 231661 330321 231664
rect 470127 231661 470193 231664
rect 322479 231576 322545 231579
rect 455247 231576 455313 231579
rect 322479 231574 455313 231576
rect 322479 231518 322484 231574
rect 322540 231518 455252 231574
rect 455308 231518 455313 231574
rect 322479 231516 455313 231518
rect 322479 231513 322545 231516
rect 455247 231513 455313 231516
rect 319503 231428 319569 231431
rect 448911 231428 448977 231431
rect 319503 231426 448977 231428
rect 319503 231370 319508 231426
rect 319564 231370 448916 231426
rect 448972 231370 448977 231426
rect 319503 231368 448977 231370
rect 319503 231365 319569 231368
rect 448911 231365 448977 231368
rect 41530 231218 41536 231282
rect 41600 231280 41606 231282
rect 41775 231280 41841 231283
rect 41600 231278 41841 231280
rect 41600 231222 41780 231278
rect 41836 231222 41841 231278
rect 41600 231220 41841 231222
rect 41600 231218 41606 231220
rect 41775 231217 41841 231220
rect 316719 231280 316785 231283
rect 442863 231280 442929 231283
rect 316719 231278 442929 231280
rect 316719 231222 316724 231278
rect 316780 231222 442868 231278
rect 442924 231222 442929 231278
rect 316719 231220 442929 231222
rect 316719 231217 316785 231220
rect 442863 231217 442929 231220
rect 147471 231132 147537 231135
rect 143904 231130 147537 231132
rect 143904 231074 147476 231130
rect 147532 231074 147537 231130
rect 143904 231072 147537 231074
rect 147471 231069 147537 231072
rect 307599 231132 307665 231135
rect 424719 231132 424785 231135
rect 307599 231130 424785 231132
rect 307599 231074 307604 231130
rect 307660 231074 424724 231130
rect 424780 231074 424785 231130
rect 307599 231072 424785 231074
rect 307599 231069 307665 231072
rect 424719 231069 424785 231072
rect 40954 230330 40960 230394
rect 41024 230392 41030 230394
rect 41775 230392 41841 230395
rect 41024 230390 41841 230392
rect 41024 230334 41780 230390
rect 41836 230334 41841 230390
rect 41024 230332 41841 230334
rect 41024 230330 41030 230332
rect 41775 230329 41841 230332
rect 408111 230392 408177 230395
rect 575055 230392 575121 230395
rect 408111 230390 575121 230392
rect 408111 230334 408116 230390
rect 408172 230334 575060 230390
rect 575116 230334 575121 230390
rect 408111 230332 575121 230334
rect 408111 230329 408177 230332
rect 575055 230329 575121 230332
rect 363567 230244 363633 230247
rect 534255 230244 534321 230247
rect 363567 230242 534321 230244
rect 363567 230186 363572 230242
rect 363628 230186 534260 230242
rect 534316 230186 534321 230242
rect 363567 230184 534321 230186
rect 363567 230181 363633 230184
rect 534255 230181 534321 230184
rect 41146 230034 41152 230098
rect 41216 230096 41222 230098
rect 41775 230096 41841 230099
rect 41216 230094 41841 230096
rect 41216 230038 41780 230094
rect 41836 230038 41841 230094
rect 41216 230036 41841 230038
rect 41216 230034 41222 230036
rect 41775 230033 41841 230036
rect 358959 230096 359025 230099
rect 527535 230096 527601 230099
rect 358959 230094 527601 230096
rect 358959 230038 358964 230094
rect 359020 230038 527540 230094
rect 527596 230038 527601 230094
rect 358959 230036 527601 230038
rect 358959 230033 359025 230036
rect 527535 230033 527601 230036
rect 147087 229948 147153 229951
rect 143904 229946 147153 229948
rect 143904 229890 147092 229946
rect 147148 229890 147153 229946
rect 143904 229888 147153 229890
rect 147087 229885 147153 229888
rect 366639 229948 366705 229951
rect 540303 229948 540369 229951
rect 366639 229946 540369 229948
rect 366639 229890 366644 229946
rect 366700 229890 540308 229946
rect 540364 229890 540369 229946
rect 366639 229888 540369 229890
rect 366639 229885 366705 229888
rect 540303 229885 540369 229888
rect 373071 229800 373137 229803
rect 553935 229800 554001 229803
rect 373071 229798 554001 229800
rect 373071 229742 373076 229798
rect 373132 229742 553940 229798
rect 553996 229742 554001 229798
rect 373071 229740 554001 229742
rect 373071 229737 373137 229740
rect 553935 229737 554001 229740
rect 379887 229652 379953 229655
rect 569775 229652 569841 229655
rect 379887 229650 569841 229652
rect 379887 229594 379892 229650
rect 379948 229594 569780 229650
rect 569836 229594 569841 229650
rect 379887 229592 569841 229594
rect 379887 229589 379953 229592
rect 569775 229589 569841 229592
rect 381327 229504 381393 229507
rect 572751 229504 572817 229507
rect 381327 229502 572817 229504
rect 381327 229446 381332 229502
rect 381388 229446 572756 229502
rect 572812 229446 572817 229502
rect 381327 229444 572817 229446
rect 381327 229441 381393 229444
rect 572751 229441 572817 229444
rect 41338 229294 41344 229358
rect 41408 229356 41414 229358
rect 41775 229356 41841 229359
rect 41408 229354 41841 229356
rect 41408 229298 41780 229354
rect 41836 229298 41841 229354
rect 41408 229296 41841 229298
rect 41408 229294 41414 229296
rect 41775 229293 41841 229296
rect 383535 229356 383601 229359
rect 573519 229356 573585 229359
rect 383535 229354 573585 229356
rect 383535 229298 383540 229354
rect 383596 229298 573524 229354
rect 573580 229298 573585 229354
rect 383535 229296 573585 229298
rect 383535 229293 383601 229296
rect 573519 229293 573585 229296
rect 296559 229208 296625 229211
rect 362799 229208 362865 229211
rect 296559 229206 362865 229208
rect 296559 229150 296564 229206
rect 296620 229150 362804 229206
rect 362860 229150 362865 229206
rect 296559 229148 362865 229150
rect 296559 229145 296625 229148
rect 362799 229145 362865 229148
rect 384399 229208 384465 229211
rect 578895 229208 578961 229211
rect 384399 229206 578961 229208
rect 384399 229150 384404 229206
rect 384460 229150 578900 229206
rect 578956 229150 578961 229206
rect 384399 229148 578961 229150
rect 384399 229145 384465 229148
rect 578895 229145 578961 229148
rect 292143 229060 292209 229063
rect 359823 229060 359889 229063
rect 292143 229058 359889 229060
rect 292143 229002 292148 229058
rect 292204 229002 359828 229058
rect 359884 229002 359889 229058
rect 292143 229000 359889 229002
rect 292143 228997 292209 229000
rect 359823 228997 359889 229000
rect 400239 229060 400305 229063
rect 599919 229060 599985 229063
rect 400239 229058 599985 229060
rect 400239 229002 400244 229058
rect 400300 229002 599924 229058
rect 599980 229002 599985 229058
rect 400239 229000 599985 229002
rect 400239 228997 400305 229000
rect 599919 228997 599985 229000
rect 293103 228912 293169 228915
rect 365679 228912 365745 228915
rect 293103 228910 365745 228912
rect 293103 228854 293108 228910
rect 293164 228854 365684 228910
rect 365740 228854 365745 228910
rect 293103 228852 365745 228854
rect 293103 228849 293169 228852
rect 365679 228849 365745 228852
rect 399471 228912 399537 228915
rect 607503 228912 607569 228915
rect 399471 228910 607569 228912
rect 399471 228854 399476 228910
rect 399532 228854 607508 228910
rect 607564 228854 607569 228910
rect 399471 228852 607569 228854
rect 399471 228849 399537 228852
rect 607503 228849 607569 228852
rect 360879 228764 360945 228767
rect 528303 228764 528369 228767
rect 360879 228762 528369 228764
rect 360879 228706 360884 228762
rect 360940 228706 528308 228762
rect 528364 228706 528369 228762
rect 360879 228704 528369 228706
rect 360879 228701 360945 228704
rect 528303 228701 528369 228704
rect 143874 228172 143934 228660
rect 342159 228616 342225 228619
rect 494223 228616 494289 228619
rect 342159 228614 494289 228616
rect 342159 228558 342164 228614
rect 342220 228558 494228 228614
rect 494284 228558 494289 228614
rect 342159 228556 494289 228558
rect 342159 228553 342225 228556
rect 494223 228553 494289 228556
rect 345423 228468 345489 228471
rect 497967 228468 498033 228471
rect 345423 228466 498033 228468
rect 345423 228410 345428 228466
rect 345484 228410 497972 228466
rect 498028 228410 498033 228466
rect 345423 228408 498033 228410
rect 345423 228405 345489 228408
rect 497967 228405 498033 228408
rect 339375 228320 339441 228323
rect 488271 228320 488337 228323
rect 339375 228318 488337 228320
rect 339375 228262 339380 228318
rect 339436 228262 488276 228318
rect 488332 228262 488337 228318
rect 339375 228260 488337 228262
rect 339375 228257 339441 228260
rect 488271 228257 488337 228260
rect 149391 228172 149457 228175
rect 143874 228170 149457 228172
rect 143874 228114 149396 228170
rect 149452 228114 149457 228170
rect 143874 228112 149457 228114
rect 149391 228109 149457 228112
rect 333039 228172 333105 228175
rect 476175 228172 476241 228175
rect 333039 228170 476241 228172
rect 333039 228114 333044 228170
rect 333100 228114 476180 228170
rect 476236 228114 476241 228170
rect 333039 228112 476241 228114
rect 333039 228109 333105 228112
rect 476175 228109 476241 228112
rect 41871 227434 41937 227435
rect 41871 227430 41920 227434
rect 41984 227432 41990 227434
rect 149487 227432 149553 227435
rect 41871 227374 41876 227430
rect 41871 227370 41920 227374
rect 41984 227372 42028 227432
rect 143904 227430 149553 227432
rect 143904 227374 149492 227430
rect 149548 227374 149553 227430
rect 143904 227372 149553 227374
rect 41984 227370 41990 227372
rect 41871 227369 41937 227370
rect 149487 227369 149553 227372
rect 336879 227432 336945 227435
rect 481455 227432 481521 227435
rect 336879 227430 481521 227432
rect 336879 227374 336884 227430
rect 336940 227374 481460 227430
rect 481516 227374 481521 227430
rect 336879 227372 481521 227374
rect 336879 227369 336945 227372
rect 481455 227369 481521 227372
rect 343119 227284 343185 227287
rect 493455 227284 493521 227287
rect 343119 227282 493521 227284
rect 343119 227226 343124 227282
rect 343180 227226 493460 227282
rect 493516 227226 493521 227282
rect 343119 227224 493521 227226
rect 343119 227221 343185 227224
rect 493455 227221 493521 227224
rect 344751 227136 344817 227139
rect 498831 227136 498897 227139
rect 344751 227134 498897 227136
rect 344751 227078 344756 227134
rect 344812 227078 498836 227134
rect 498892 227078 498897 227134
rect 344751 227076 498897 227078
rect 344751 227073 344817 227076
rect 498831 227073 498897 227076
rect 391599 226988 391665 226991
rect 591663 226988 591729 226991
rect 391599 226986 591729 226988
rect 391599 226930 391604 226986
rect 391660 226930 591668 226986
rect 591724 226930 591729 226986
rect 391599 226928 591729 226930
rect 391599 226925 391665 226928
rect 591663 226925 591729 226928
rect 40762 226778 40768 226842
rect 40832 226840 40838 226842
rect 41775 226840 41841 226843
rect 40832 226838 41841 226840
rect 40832 226782 41780 226838
rect 41836 226782 41841 226838
rect 40832 226780 41841 226782
rect 40832 226778 40838 226780
rect 41775 226777 41841 226780
rect 391215 226840 391281 226843
rect 590895 226840 590961 226843
rect 391215 226838 590961 226840
rect 391215 226782 391220 226838
rect 391276 226782 590900 226838
rect 590956 226782 590961 226838
rect 391215 226780 590961 226782
rect 391215 226777 391281 226780
rect 590895 226777 590961 226780
rect 394095 226692 394161 226695
rect 596175 226692 596241 226695
rect 394095 226690 596241 226692
rect 394095 226634 394100 226690
rect 394156 226634 596180 226690
rect 596236 226634 596241 226690
rect 394095 226632 596241 226634
rect 394095 226629 394161 226632
rect 596175 226629 596241 226632
rect 394479 226544 394545 226547
rect 596943 226544 597009 226547
rect 394479 226542 597009 226544
rect 394479 226486 394484 226542
rect 394540 226486 596948 226542
rect 597004 226486 597009 226542
rect 394479 226484 597009 226486
rect 394479 226481 394545 226484
rect 596943 226481 597009 226484
rect 42159 226398 42225 226399
rect 42106 226396 42112 226398
rect 42068 226336 42112 226396
rect 42176 226394 42225 226398
rect 147087 226396 147153 226399
rect 42220 226338 42225 226394
rect 42106 226334 42112 226336
rect 42176 226334 42225 226338
rect 143904 226394 147153 226396
rect 143904 226338 147092 226394
rect 147148 226338 147153 226394
rect 143904 226336 147153 226338
rect 42159 226333 42225 226334
rect 147087 226333 147153 226336
rect 404367 226396 404433 226399
rect 617295 226396 617361 226399
rect 404367 226394 617361 226396
rect 404367 226338 404372 226394
rect 404428 226338 617300 226394
rect 617356 226338 617361 226394
rect 404367 226336 617361 226338
rect 404367 226333 404433 226336
rect 617295 226333 617361 226336
rect 405711 226248 405777 226251
rect 620367 226248 620433 226251
rect 405711 226246 620433 226248
rect 405711 226190 405716 226246
rect 405772 226190 620372 226246
rect 620428 226190 620433 226246
rect 405711 226188 620433 226190
rect 405711 226185 405777 226188
rect 620367 226185 620433 226188
rect 407631 226100 407697 226103
rect 623343 226100 623409 226103
rect 407631 226098 623409 226100
rect 407631 226042 407636 226098
rect 407692 226042 623348 226098
rect 623404 226042 623409 226098
rect 407631 226040 623409 226042
rect 407631 226037 407697 226040
rect 623343 226037 623409 226040
rect 340143 225952 340209 225955
rect 487503 225952 487569 225955
rect 340143 225950 487569 225952
rect 340143 225894 340148 225950
rect 340204 225894 487508 225950
rect 487564 225894 487569 225950
rect 340143 225892 487569 225894
rect 340143 225889 340209 225892
rect 487503 225889 487569 225892
rect 330831 225804 330897 225807
rect 469359 225804 469425 225807
rect 330831 225802 469425 225804
rect 330831 225746 330836 225802
rect 330892 225746 469364 225802
rect 469420 225746 469425 225802
rect 330831 225744 469425 225746
rect 330831 225741 330897 225744
rect 469359 225741 469425 225744
rect 328047 225656 328113 225659
rect 463311 225656 463377 225659
rect 328047 225654 463377 225656
rect 328047 225598 328052 225654
rect 328108 225598 463316 225654
rect 463372 225598 463377 225654
rect 328047 225596 463377 225598
rect 328047 225593 328113 225596
rect 463311 225593 463377 225596
rect 327759 225508 327825 225511
rect 457263 225508 457329 225511
rect 327759 225506 457329 225508
rect 327759 225450 327764 225506
rect 327820 225450 457268 225506
rect 457324 225450 457329 225506
rect 327759 225448 457329 225450
rect 327759 225445 327825 225448
rect 457263 225445 457329 225448
rect 318927 225360 318993 225363
rect 445167 225360 445233 225363
rect 318927 225358 445233 225360
rect 318927 225302 318932 225358
rect 318988 225302 445172 225358
rect 445228 225302 445233 225358
rect 318927 225300 445233 225302
rect 318927 225297 318993 225300
rect 445167 225297 445233 225300
rect 149391 225212 149457 225215
rect 143904 225210 149457 225212
rect 143904 225154 149396 225210
rect 149452 225154 149457 225210
rect 143904 225152 149457 225154
rect 149391 225149 149457 225152
rect 368655 225212 368721 225215
rect 475311 225212 475377 225215
rect 368655 225210 475377 225212
rect 368655 225154 368660 225210
rect 368716 225154 475316 225210
rect 475372 225154 475377 225210
rect 368655 225152 475377 225154
rect 368655 225149 368721 225152
rect 475311 225149 475377 225152
rect 358575 224620 358641 224623
rect 525999 224620 526065 224623
rect 358575 224618 526065 224620
rect 358575 224562 358580 224618
rect 358636 224562 526004 224618
rect 526060 224562 526065 224618
rect 358575 224560 526065 224562
rect 358575 224557 358641 224560
rect 525999 224557 526065 224560
rect 359439 224472 359505 224475
rect 526671 224472 526737 224475
rect 359439 224470 526737 224472
rect 359439 224414 359444 224470
rect 359500 224414 526676 224470
rect 526732 224414 526737 224470
rect 359439 224412 526737 224414
rect 359439 224409 359505 224412
rect 526671 224409 526737 224412
rect 359727 224324 359793 224327
rect 528975 224324 529041 224327
rect 359727 224322 529041 224324
rect 359727 224266 359732 224322
rect 359788 224266 528980 224322
rect 529036 224266 529041 224322
rect 359727 224264 529041 224266
rect 359727 224261 359793 224264
rect 528975 224261 529041 224264
rect 360303 224176 360369 224179
rect 530511 224176 530577 224179
rect 360303 224174 530577 224176
rect 360303 224118 360308 224174
rect 360364 224118 530516 224174
rect 530572 224118 530577 224174
rect 360303 224116 530577 224118
rect 360303 224113 360369 224116
rect 530511 224113 530577 224116
rect 361455 224028 361521 224031
rect 532047 224028 532113 224031
rect 361455 224026 532113 224028
rect 361455 223970 361460 224026
rect 361516 223970 532052 224026
rect 532108 223970 532113 224026
rect 361455 223968 532113 223970
rect 361455 223965 361521 223968
rect 532047 223965 532113 223968
rect 149487 223880 149553 223883
rect 143904 223878 149553 223880
rect 143904 223822 149492 223878
rect 149548 223822 149553 223878
rect 143904 223820 149553 223822
rect 149487 223817 149553 223820
rect 364143 223880 364209 223883
rect 536559 223880 536625 223883
rect 364143 223878 536625 223880
rect 364143 223822 364148 223878
rect 364204 223822 536564 223878
rect 536620 223822 536625 223878
rect 364143 223820 536625 223822
rect 364143 223817 364209 223820
rect 536559 223817 536625 223820
rect 367599 223732 367665 223735
rect 544047 223732 544113 223735
rect 367599 223730 544113 223732
rect 367599 223674 367604 223730
rect 367660 223674 544052 223730
rect 544108 223674 544113 223730
rect 367599 223672 544113 223674
rect 367599 223669 367665 223672
rect 544047 223669 544113 223672
rect 377583 223584 377649 223587
rect 562959 223584 563025 223587
rect 377583 223582 563025 223584
rect 377583 223526 377588 223582
rect 377644 223526 562964 223582
rect 563020 223526 563025 223582
rect 377583 223524 563025 223526
rect 377583 223521 377649 223524
rect 562959 223521 563025 223524
rect 376719 223436 376785 223439
rect 562191 223436 562257 223439
rect 376719 223434 562257 223436
rect 376719 223378 376724 223434
rect 376780 223378 562196 223434
rect 562252 223378 562257 223434
rect 376719 223376 562257 223378
rect 376719 223373 376785 223376
rect 562191 223373 562257 223376
rect 381231 223288 381297 223291
rect 571311 223288 571377 223291
rect 381231 223286 571377 223288
rect 381231 223230 381236 223286
rect 381292 223230 571316 223286
rect 571372 223230 571377 223286
rect 381231 223228 571377 223230
rect 381231 223225 381297 223228
rect 571311 223225 571377 223228
rect 384303 223140 384369 223143
rect 577263 223140 577329 223143
rect 384303 223138 577329 223140
rect 384303 223082 384308 223138
rect 384364 223082 577268 223138
rect 577324 223082 577329 223138
rect 384303 223080 577329 223082
rect 384303 223077 384369 223080
rect 577263 223077 577329 223080
rect 354159 222992 354225 222995
rect 518415 222992 518481 222995
rect 354159 222990 518481 222992
rect 354159 222934 354164 222990
rect 354220 222934 518420 222990
rect 518476 222934 518481 222990
rect 354159 222932 518481 222934
rect 354159 222929 354225 222932
rect 518415 222929 518481 222932
rect 357231 222844 357297 222847
rect 524463 222844 524529 222847
rect 357231 222842 524529 222844
rect 357231 222786 357236 222842
rect 357292 222786 524468 222842
rect 524524 222786 524529 222842
rect 357231 222784 524529 222786
rect 357231 222781 357297 222784
rect 524463 222781 524529 222784
rect 149391 222696 149457 222699
rect 143904 222694 149457 222696
rect 143904 222638 149396 222694
rect 149452 222638 149457 222694
rect 143904 222636 149457 222638
rect 149391 222633 149457 222636
rect 355599 222696 355665 222699
rect 519855 222696 519921 222699
rect 355599 222694 519921 222696
rect 355599 222638 355604 222694
rect 355660 222638 519860 222694
rect 519916 222638 519921 222694
rect 355599 222636 519921 222638
rect 355599 222633 355665 222636
rect 519855 222633 519921 222636
rect 406479 222548 406545 222551
rect 522927 222548 522993 222551
rect 406479 222546 522993 222548
rect 406479 222490 406484 222546
rect 406540 222490 522932 222546
rect 522988 222490 522993 222546
rect 406479 222488 522993 222490
rect 406479 222485 406545 222488
rect 522927 222485 522993 222488
rect 149487 221512 149553 221515
rect 143904 221510 149553 221512
rect 143904 221454 149492 221510
rect 149548 221454 149553 221510
rect 143904 221452 149553 221454
rect 149487 221449 149553 221452
rect 186927 221068 186993 221071
rect 186927 221066 190560 221068
rect 186927 221010 186932 221066
rect 186988 221010 190560 221066
rect 186927 221008 190560 221010
rect 186927 221005 186993 221008
rect 185583 220328 185649 220331
rect 185583 220326 190560 220328
rect 185583 220270 185588 220326
rect 185644 220270 190560 220326
rect 185583 220268 190560 220270
rect 185583 220265 185649 220268
rect 143874 219736 143934 220224
rect 149391 219736 149457 219739
rect 143874 219734 149457 219736
rect 143874 219678 149396 219734
rect 149452 219678 149457 219734
rect 143874 219676 149457 219678
rect 149391 219673 149457 219676
rect 184335 219588 184401 219591
rect 184335 219586 190560 219588
rect 184335 219530 184340 219586
rect 184396 219530 190560 219586
rect 184335 219528 190560 219530
rect 184335 219525 184401 219528
rect 149391 218996 149457 218999
rect 143904 218994 149457 218996
rect 143904 218938 149396 218994
rect 149452 218938 149457 218994
rect 143904 218936 149457 218938
rect 149391 218933 149457 218936
rect 184335 218848 184401 218851
rect 184335 218846 190560 218848
rect 184335 218790 184340 218846
rect 184396 218790 190560 218846
rect 184335 218788 190560 218790
rect 184335 218785 184401 218788
rect 639810 218670 639870 220594
rect 676290 219739 676350 220076
rect 676239 219734 676350 219739
rect 676239 219678 676244 219734
rect 676300 219678 676350 219734
rect 676239 219676 676350 219678
rect 676239 219673 676305 219676
rect 676290 219295 676350 219558
rect 676239 219290 676350 219295
rect 676239 219234 676244 219290
rect 676300 219234 676350 219290
rect 676239 219232 676350 219234
rect 676239 219229 676305 219232
rect 676047 218996 676113 218999
rect 676047 218994 676320 218996
rect 676047 218938 676052 218994
rect 676108 218938 676320 218994
rect 676047 218936 676320 218938
rect 676047 218933 676113 218936
rect 674554 218490 674560 218554
rect 674624 218552 674630 218554
rect 674624 218492 676320 218552
rect 674624 218490 674630 218492
rect 674170 218342 674176 218406
rect 674240 218404 674246 218406
rect 674554 218404 674560 218406
rect 674240 218344 674560 218404
rect 674240 218342 674246 218344
rect 674554 218342 674560 218344
rect 674624 218342 674630 218406
rect 187023 218108 187089 218111
rect 187023 218106 190560 218108
rect 187023 218050 187028 218106
rect 187084 218050 190560 218106
rect 187023 218048 190560 218050
rect 187023 218045 187089 218048
rect 147279 217812 147345 217815
rect 143904 217810 147345 217812
rect 143904 217754 147284 217810
rect 147340 217754 147345 217810
rect 143904 217752 147345 217754
rect 147279 217749 147345 217752
rect 190146 217294 190206 218048
rect 674170 218046 674176 218110
rect 674240 218108 674246 218110
rect 674240 218048 676320 218108
rect 674240 218046 674246 218048
rect 673978 217454 673984 217518
rect 674048 217516 674054 217518
rect 674048 217456 676320 217516
rect 674048 217454 674054 217456
rect 673978 217306 673984 217370
rect 674048 217368 674054 217370
rect 674554 217368 674560 217370
rect 674048 217308 674560 217368
rect 674048 217306 674054 217308
rect 674554 217306 674560 217308
rect 674624 217306 674630 217370
rect 190146 217234 190560 217294
rect 674362 217010 674368 217074
rect 674432 217072 674438 217074
rect 674432 217012 676320 217072
rect 674432 217010 674438 217012
rect 674746 216862 674752 216926
rect 674816 216924 674822 216926
rect 674816 216864 676350 216924
rect 674816 216862 674822 216864
rect 149391 216628 149457 216631
rect 143904 216626 149457 216628
rect 143904 216570 149396 216626
rect 149452 216570 149457 216626
rect 143904 216568 149457 216570
rect 149391 216565 149457 216568
rect 186831 216480 186897 216483
rect 186831 216478 190560 216480
rect 186831 216422 186836 216478
rect 186892 216422 190560 216478
rect 186831 216420 190560 216422
rect 186831 216417 186897 216420
rect 190146 215814 190206 216420
rect 190146 215754 190560 215814
rect 143874 214852 143934 215340
rect 186543 215000 186609 215003
rect 186543 214998 190560 215000
rect 186543 214942 186548 214998
rect 186604 214942 190560 214998
rect 186543 214940 190560 214942
rect 186543 214937 186609 214940
rect 149487 214852 149553 214855
rect 143874 214850 149553 214852
rect 143874 214794 149492 214850
rect 149548 214794 149553 214850
rect 143874 214792 149553 214794
rect 149487 214789 149553 214792
rect 190146 214334 190206 214940
rect 640386 214822 640446 216746
rect 676290 216524 676350 216864
rect 673978 215974 673984 216038
rect 674048 216036 674054 216038
rect 674048 215976 676320 216036
rect 674048 215974 674054 215976
rect 676290 215447 676350 215562
rect 676239 215442 676350 215447
rect 676239 215386 676244 215442
rect 676300 215386 676350 215442
rect 676239 215384 676350 215386
rect 676239 215381 676305 215384
rect 674554 214642 674560 214706
rect 674624 214704 674630 214706
rect 676290 214704 676350 215044
rect 674624 214644 676350 214704
rect 674624 214642 674630 214644
rect 675567 214556 675633 214559
rect 675567 214554 676320 214556
rect 675567 214498 675572 214554
rect 675628 214498 676320 214554
rect 675567 214496 676320 214498
rect 675567 214493 675633 214496
rect 190146 214274 190560 214334
rect 149391 214112 149457 214115
rect 143904 214110 149457 214112
rect 143904 214054 149396 214110
rect 149452 214054 149457 214110
rect 143904 214052 149457 214054
rect 149391 214049 149457 214052
rect 676047 214112 676113 214115
rect 676047 214110 676320 214112
rect 676047 214054 676052 214110
rect 676108 214054 676320 214110
rect 676047 214052 676320 214054
rect 676047 214049 676113 214052
rect 186351 213520 186417 213523
rect 186351 213518 190560 213520
rect 186351 213462 186356 213518
rect 186412 213462 190560 213518
rect 186351 213460 190560 213462
rect 186351 213457 186417 213460
rect 41775 213298 41841 213301
rect 41568 213296 41841 213298
rect 41568 213240 41780 213296
rect 41836 213240 41841 213296
rect 41568 213238 41841 213240
rect 41775 213235 41841 213238
rect 41583 212928 41649 212931
rect 146895 212928 146961 212931
rect 41538 212926 41649 212928
rect 41538 212870 41588 212926
rect 41644 212870 41649 212926
rect 41538 212865 41649 212870
rect 143904 212926 146961 212928
rect 143904 212870 146900 212926
rect 146956 212870 146961 212926
rect 143904 212868 146961 212870
rect 146895 212865 146961 212868
rect 41538 212750 41598 212865
rect 190146 212706 190206 213460
rect 674746 213458 674752 213522
rect 674816 213520 674822 213522
rect 674816 213460 676320 213520
rect 674816 213458 674822 213460
rect 190146 212646 190560 212706
rect 640194 212339 640254 212898
rect 676866 212783 676926 213046
rect 676866 212778 676977 212783
rect 676866 212722 676916 212778
rect 676972 212722 676977 212778
rect 676866 212720 676977 212722
rect 676911 212717 676977 212720
rect 675279 212632 675345 212635
rect 675279 212630 676320 212632
rect 675279 212574 675284 212630
rect 675340 212574 676320 212630
rect 675279 212572 676320 212574
rect 675279 212569 675345 212572
rect 640143 212334 640254 212339
rect 640143 212278 640148 212334
rect 640204 212278 640254 212334
rect 640143 212276 640254 212278
rect 640143 212273 640209 212276
rect 41775 212188 41841 212191
rect 41568 212186 41841 212188
rect 41568 212130 41780 212186
rect 41836 212130 41841 212186
rect 41568 212128 41841 212130
rect 41775 212125 41841 212128
rect 186735 212040 186801 212043
rect 186735 212038 190560 212040
rect 186735 211982 186740 212038
rect 186796 211982 190560 212038
rect 186735 211980 190560 211982
rect 186735 211977 186801 211980
rect 41775 211744 41841 211747
rect 147087 211744 147153 211747
rect 41568 211742 41841 211744
rect 41568 211686 41780 211742
rect 41836 211686 41841 211742
rect 41568 211684 41841 211686
rect 143904 211742 147153 211744
rect 143904 211686 147092 211742
rect 147148 211686 147153 211742
rect 143904 211684 147153 211686
rect 41775 211681 41841 211684
rect 147087 211681 147153 211684
rect 41583 211448 41649 211451
rect 41538 211446 41649 211448
rect 41538 211390 41588 211446
rect 41644 211390 41649 211446
rect 41538 211385 41649 211390
rect 41538 211270 41598 211385
rect 190146 211152 190206 211980
rect 676290 211895 676350 212010
rect 676239 211890 676350 211895
rect 676239 211834 676244 211890
rect 676300 211834 676350 211890
rect 676239 211832 676350 211834
rect 676239 211829 676305 211832
rect 640143 211596 640209 211599
rect 640143 211594 640254 211596
rect 640143 211538 640148 211594
rect 640204 211538 640254 211594
rect 640143 211533 640254 211538
rect 190146 211092 190560 211152
rect 640194 210974 640254 211533
rect 676047 211522 676113 211525
rect 676047 211520 676320 211522
rect 676047 211464 676052 211520
rect 676108 211464 676320 211520
rect 676047 211462 676320 211464
rect 676047 211459 676113 211462
rect 676866 210859 676926 211122
rect 676815 210854 676926 210859
rect 676815 210798 676820 210854
rect 676876 210798 676926 210854
rect 676815 210796 676926 210798
rect 676815 210793 676881 210796
rect 41775 210708 41841 210711
rect 41568 210706 41841 210708
rect 41568 210650 41780 210706
rect 41836 210650 41841 210706
rect 41568 210648 41841 210650
rect 41775 210645 41841 210648
rect 186447 210560 186513 210563
rect 186447 210558 190206 210560
rect 186447 210502 186452 210558
rect 186508 210502 190206 210558
rect 186447 210500 190206 210502
rect 186447 210497 186513 210500
rect 190146 210486 190206 210500
rect 675130 210498 675136 210562
rect 675200 210560 675206 210562
rect 675200 210500 676320 210560
rect 675200 210498 675206 210500
rect 190146 210426 190560 210486
rect 147471 210412 147537 210415
rect 143904 210410 147537 210412
rect 143904 210354 147476 210410
rect 147532 210354 147537 210410
rect 143904 210352 147537 210354
rect 147471 210349 147537 210352
rect 41775 210264 41841 210267
rect 41568 210262 41841 210264
rect 41568 210206 41780 210262
rect 41836 210206 41841 210262
rect 41568 210204 41841 210206
rect 41775 210201 41841 210204
rect 41583 209968 41649 209971
rect 41538 209966 41649 209968
rect 41538 209910 41588 209966
rect 41644 209910 41649 209966
rect 41538 209905 41649 209910
rect 41538 209790 41598 209905
rect 190146 209672 190206 210426
rect 676047 210042 676113 210045
rect 676047 210040 676320 210042
rect 676047 209984 676052 210040
rect 676108 209984 676320 210040
rect 676047 209982 676320 209984
rect 676047 209979 676113 209982
rect 675951 209672 676017 209675
rect 190146 209612 190560 209672
rect 675951 209670 676320 209672
rect 675951 209614 675956 209670
rect 676012 209614 676320 209670
rect 675951 209612 676320 209614
rect 675951 209609 676017 209612
rect 41583 209376 41649 209379
rect 41538 209374 41649 209376
rect 41538 209318 41588 209374
rect 41644 209318 41649 209374
rect 41538 209313 41649 209318
rect 41538 209198 41598 209313
rect 146895 209228 146961 209231
rect 143904 209226 146961 209228
rect 143904 209170 146900 209226
rect 146956 209170 146961 209226
rect 143904 209168 146961 209170
rect 146895 209165 146961 209168
rect 186639 209080 186705 209083
rect 186639 209078 190206 209080
rect 186639 209022 186644 209078
rect 186700 209022 190206 209078
rect 186639 209020 190206 209022
rect 186639 209017 186705 209020
rect 190146 209006 190206 209020
rect 190146 208946 190560 209006
rect 42106 208784 42112 208786
rect 41568 208724 42112 208784
rect 42106 208722 42112 208724
rect 42176 208722 42182 208786
rect 41538 207898 41598 208236
rect 190146 208192 190206 208946
rect 190146 208132 190560 208192
rect 147183 208044 147249 208047
rect 143904 208042 147249 208044
rect 143904 207986 147188 208042
rect 147244 207986 147249 208042
rect 143904 207984 147249 207986
rect 147183 207981 147249 207984
rect 41530 207834 41536 207898
rect 41600 207834 41606 207898
rect 41914 207748 41920 207750
rect 41568 207688 41920 207748
rect 41914 207686 41920 207688
rect 41984 207686 41990 207750
rect 190146 207318 190560 207378
rect 186255 207304 186321 207307
rect 190146 207304 190206 207318
rect 186255 207302 190206 207304
rect 40962 207010 41022 207274
rect 186255 207246 186260 207302
rect 186316 207246 190206 207302
rect 639810 207274 639870 209124
rect 674938 209018 674944 209082
rect 675008 209080 675014 209082
rect 675008 209020 676320 209080
rect 675008 209018 675014 209020
rect 679938 208343 679998 208458
rect 679887 208338 679998 208343
rect 679887 208282 679892 208338
rect 679948 208282 679998 208338
rect 679887 208280 679998 208282
rect 679887 208277 679953 208280
rect 679746 207751 679806 208088
rect 679887 207896 679953 207899
rect 679887 207894 679998 207896
rect 679887 207838 679892 207894
rect 679948 207838 679998 207894
rect 679887 207833 679998 207838
rect 679746 207746 679857 207751
rect 679746 207690 679796 207746
rect 679852 207690 679857 207746
rect 679746 207688 679857 207690
rect 679791 207685 679857 207688
rect 679938 207570 679998 207833
rect 679791 207304 679857 207307
rect 679746 207302 679857 207304
rect 186255 207244 190206 207246
rect 186255 207241 186321 207244
rect 40954 206946 40960 207010
rect 41024 206946 41030 207010
rect 40578 206418 40638 206682
rect 40570 206354 40576 206418
rect 40640 206354 40646 206418
rect 143874 206416 143934 206904
rect 190146 206712 190206 207244
rect 679746 207246 679796 207302
rect 679852 207246 679857 207302
rect 679746 207241 679857 207246
rect 679746 206978 679806 207241
rect 190146 206652 190560 206712
rect 146895 206416 146961 206419
rect 143874 206414 146961 206416
rect 143874 206358 146900 206414
rect 146956 206358 146961 206414
rect 143874 206356 146961 206358
rect 146895 206353 146961 206356
rect 41775 206268 41841 206271
rect 41568 206266 41841 206268
rect 41568 206210 41780 206266
rect 41836 206210 41841 206266
rect 41568 206208 41841 206210
rect 41775 206205 41841 206208
rect 186063 205972 186129 205975
rect 186063 205970 190206 205972
rect 186063 205914 186068 205970
rect 186124 205914 190206 205970
rect 186063 205912 190206 205914
rect 186063 205909 186129 205912
rect 190146 205898 190206 205912
rect 190146 205838 190560 205898
rect 40770 205530 40830 205794
rect 149487 205676 149553 205679
rect 143904 205674 149553 205676
rect 143904 205618 149492 205674
rect 149548 205618 149553 205674
rect 143904 205616 149553 205618
rect 149487 205613 149553 205616
rect 40762 205466 40768 205530
rect 40832 205466 40838 205530
rect 190146 205232 190206 205838
rect 41346 204938 41406 205202
rect 190146 205172 190560 205232
rect 41338 204874 41344 204938
rect 41408 204874 41414 204938
rect 41154 204494 41214 204758
rect 41146 204430 41152 204494
rect 41216 204430 41222 204494
rect 149391 204492 149457 204495
rect 143904 204490 149457 204492
rect 143904 204434 149396 204490
rect 149452 204434 149457 204490
rect 143904 204432 149457 204434
rect 149391 204429 149457 204432
rect 185967 204344 186033 204347
rect 185967 204342 190560 204344
rect 40386 204050 40446 204314
rect 185967 204286 185972 204342
rect 186028 204286 190560 204342
rect 185967 204284 190560 204286
rect 185967 204281 186033 204284
rect 40378 203986 40384 204050
rect 40448 203986 40454 204050
rect 42490 203752 42496 203754
rect 41568 203692 42496 203752
rect 42490 203690 42496 203692
rect 42560 203690 42566 203754
rect 190146 203604 190206 204284
rect 190146 203544 190560 203604
rect 639810 203426 639870 205350
rect 675706 204726 675712 204790
rect 675776 204788 675782 204790
rect 676911 204788 676977 204791
rect 675776 204786 676977 204788
rect 675776 204730 676916 204786
rect 676972 204730 676977 204786
rect 675776 204728 676977 204730
rect 675776 204726 675782 204728
rect 676911 204725 676977 204728
rect 675898 204578 675904 204642
rect 675968 204640 675974 204642
rect 676815 204640 676881 204643
rect 675968 204638 676881 204640
rect 675968 204582 676820 204638
rect 676876 204582 676881 204638
rect 675968 204580 676881 204582
rect 675968 204578 675974 204580
rect 676815 204577 676881 204580
rect 147855 203308 147921 203311
rect 143904 203306 147921 203308
rect 143904 203250 147860 203306
rect 147916 203250 147921 203306
rect 143904 203248 147921 203250
rect 147855 203245 147921 203248
rect 41538 203012 41598 203204
rect 42682 203012 42688 203014
rect 41538 202952 42688 203012
rect 42682 202950 42688 202952
rect 42752 202950 42758 203014
rect 41722 202864 41728 202866
rect 41568 202804 41728 202864
rect 41722 202802 41728 202804
rect 41792 202802 41798 202866
rect 186159 202864 186225 202867
rect 186159 202862 190560 202864
rect 186159 202806 186164 202862
rect 186220 202806 190560 202862
rect 186159 202804 190560 202806
rect 186159 202801 186225 202804
rect 42298 202272 42304 202274
rect 41568 202212 42304 202272
rect 42298 202210 42304 202212
rect 42368 202210 42374 202274
rect 190146 202124 190206 202804
rect 190146 202064 190560 202124
rect 41871 201680 41937 201683
rect 41568 201678 41937 201680
rect 41568 201622 41876 201678
rect 41932 201622 41937 201678
rect 41568 201620 41937 201622
rect 143874 201680 143934 202020
rect 149391 201680 149457 201683
rect 143874 201678 149457 201680
rect 143874 201622 149396 201678
rect 149452 201622 149457 201678
rect 143874 201620 149457 201622
rect 41871 201617 41937 201620
rect 149391 201617 149457 201620
rect 41583 201532 41649 201535
rect 41538 201530 41649 201532
rect 41538 201474 41588 201530
rect 41644 201474 41649 201530
rect 41538 201469 41649 201474
rect 41538 201354 41598 201469
rect 190287 201384 190353 201387
rect 190287 201382 190560 201384
rect 190287 201326 190292 201382
rect 190348 201326 190560 201382
rect 190287 201324 190560 201326
rect 190287 201321 190353 201324
rect 640194 200943 640254 201502
rect 41583 200940 41649 200943
rect 41538 200938 41649 200940
rect 41538 200882 41588 200938
rect 41644 200882 41649 200938
rect 41538 200877 41649 200882
rect 640143 200938 640254 200943
rect 640143 200882 640148 200938
rect 640204 200882 640254 200938
rect 640143 200880 640254 200882
rect 640143 200877 640209 200880
rect 41538 200762 41598 200877
rect 149391 200792 149457 200795
rect 143904 200790 149457 200792
rect 143904 200734 149396 200790
rect 149452 200734 149457 200790
rect 143904 200732 149457 200734
rect 149391 200729 149457 200732
rect 190287 200570 190353 200573
rect 190287 200568 190560 200570
rect 190287 200512 190292 200568
rect 190348 200512 190560 200568
rect 190287 200510 190560 200512
rect 190287 200507 190353 200510
rect 640143 200200 640209 200203
rect 640143 200198 640254 200200
rect 640143 200142 640148 200198
rect 640204 200142 640254 200198
rect 640143 200137 640254 200142
rect 184335 199756 184401 199759
rect 184335 199754 190560 199756
rect 184335 199698 184340 199754
rect 184396 199698 190560 199754
rect 184335 199696 190560 199698
rect 184335 199693 184401 199696
rect 147567 199608 147633 199611
rect 143904 199606 147633 199608
rect 143904 199550 147572 199606
rect 147628 199550 147633 199606
rect 640194 199578 640254 200137
rect 143904 199548 147633 199550
rect 147567 199545 147633 199548
rect 187215 199164 187281 199167
rect 187215 199162 190014 199164
rect 187215 199106 187220 199162
rect 187276 199106 190014 199162
rect 187215 199104 190014 199106
rect 187215 199101 187281 199104
rect 189954 199090 190014 199104
rect 189954 199030 190560 199090
rect 149295 198424 149361 198427
rect 143904 198422 149361 198424
rect 143904 198366 149300 198422
rect 149356 198366 149361 198422
rect 143904 198364 149361 198366
rect 149295 198361 149361 198364
rect 185487 198276 185553 198279
rect 185487 198274 190560 198276
rect 185487 198218 185492 198274
rect 185548 198218 190560 198274
rect 185487 198216 190560 198218
rect 185487 198213 185553 198216
rect 184239 197684 184305 197687
rect 674170 197684 674176 197686
rect 184239 197682 190014 197684
rect 184239 197626 184244 197682
rect 184300 197626 190014 197682
rect 184239 197624 190014 197626
rect 184239 197621 184305 197624
rect 189954 197610 190014 197624
rect 189954 197550 190560 197610
rect 149391 197092 149457 197095
rect 143904 197090 149457 197092
rect 143904 197034 149396 197090
rect 149452 197034 149457 197090
rect 143904 197032 149457 197034
rect 149391 197029 149457 197032
rect 184335 196796 184401 196799
rect 184335 196794 190560 196796
rect 184335 196738 184340 196794
rect 184396 196738 190560 196794
rect 184335 196736 190560 196738
rect 184335 196733 184401 196736
rect 184431 196056 184497 196059
rect 184431 196054 190560 196056
rect 184431 195998 184436 196054
rect 184492 195998 190560 196054
rect 184431 195996 190560 195998
rect 184431 195993 184497 195996
rect 147279 195908 147345 195911
rect 143904 195906 147345 195908
rect 143904 195850 147284 195906
rect 147340 195850 147345 195906
rect 143904 195848 147345 195850
rect 147279 195845 147345 195848
rect 639810 195730 639870 197654
rect 673986 197624 674176 197684
rect 673986 197242 674046 197624
rect 674170 197622 674176 197624
rect 674240 197622 674246 197686
rect 673978 197178 673984 197242
rect 674048 197178 674054 197242
rect 41530 195402 41536 195466
rect 41600 195464 41606 195466
rect 41871 195464 41937 195467
rect 41600 195462 41937 195464
rect 41600 195406 41876 195462
rect 41932 195406 41937 195462
rect 41600 195404 41937 195406
rect 41600 195402 41606 195404
rect 41871 195401 41937 195404
rect 184335 195316 184401 195319
rect 184335 195314 190560 195316
rect 184335 195258 184340 195314
rect 184396 195258 190560 195314
rect 184335 195256 190560 195258
rect 184335 195253 184401 195256
rect 674746 195106 674752 195170
rect 674816 195168 674822 195170
rect 675471 195168 675537 195171
rect 674816 195166 675537 195168
rect 674816 195110 675476 195166
rect 675532 195110 675537 195166
rect 674816 195108 675537 195110
rect 674816 195106 674822 195108
rect 675471 195105 675537 195108
rect 149487 194724 149553 194727
rect 143904 194722 149553 194724
rect 143904 194666 149492 194722
rect 149548 194666 149553 194722
rect 143904 194664 149553 194666
rect 149487 194661 149553 194664
rect 184431 194428 184497 194431
rect 184431 194426 190560 194428
rect 184431 194370 184436 194426
rect 184492 194370 190560 194426
rect 184431 194368 190560 194370
rect 184431 194365 184497 194368
rect 675130 193922 675136 193986
rect 675200 193984 675206 193986
rect 675375 193984 675441 193987
rect 675200 193982 675441 193984
rect 675200 193926 675380 193982
rect 675436 193926 675441 193982
rect 675200 193924 675441 193926
rect 675200 193922 675206 193924
rect 675375 193921 675441 193924
rect 184527 193836 184593 193839
rect 184527 193834 190014 193836
rect 184527 193778 184532 193834
rect 184588 193778 190014 193834
rect 184527 193776 190014 193778
rect 184527 193773 184593 193776
rect 189954 193762 190014 193776
rect 189954 193702 190560 193762
rect 40378 193626 40384 193690
rect 40448 193688 40454 193690
rect 41775 193688 41841 193691
rect 40448 193686 41841 193688
rect 40448 193630 41780 193686
rect 41836 193630 41841 193686
rect 40448 193628 41841 193630
rect 40448 193626 40454 193628
rect 41775 193625 41841 193628
rect 143874 193244 143934 193436
rect 149391 193244 149457 193247
rect 143874 193242 149457 193244
rect 143874 193186 149396 193242
rect 149452 193186 149457 193242
rect 143874 193184 149457 193186
rect 149391 193181 149457 193184
rect 184431 192948 184497 192951
rect 184431 192946 190560 192948
rect 184431 192890 184436 192946
rect 184492 192890 190560 192946
rect 184431 192888 190560 192890
rect 184431 192885 184497 192888
rect 42159 192356 42225 192359
rect 42298 192356 42304 192358
rect 42159 192354 42304 192356
rect 42159 192298 42164 192354
rect 42220 192298 42304 192354
rect 42159 192296 42304 192298
rect 42159 192293 42225 192296
rect 42298 192294 42304 192296
rect 42368 192294 42374 192358
rect 184335 192356 184401 192359
rect 184335 192354 190014 192356
rect 184335 192298 184340 192354
rect 184396 192298 190014 192354
rect 184335 192296 190014 192298
rect 184335 192293 184401 192296
rect 189954 192282 190014 192296
rect 189954 192222 190560 192282
rect 149487 192208 149553 192211
rect 143904 192206 149553 192208
rect 143904 192150 149492 192206
rect 149548 192150 149553 192206
rect 143904 192148 149553 192150
rect 149487 192145 149553 192148
rect 639810 192030 639870 193880
rect 674938 193034 674944 193098
rect 675008 193096 675014 193098
rect 675471 193096 675537 193099
rect 675008 193094 675537 193096
rect 675008 193038 675476 193094
rect 675532 193038 675537 193094
rect 675008 193036 675537 193038
rect 675008 193034 675014 193036
rect 675471 193033 675537 193036
rect 675759 192208 675825 192211
rect 675898 192208 675904 192210
rect 675759 192206 675904 192208
rect 675759 192150 675764 192206
rect 675820 192150 675904 192206
rect 675759 192148 675904 192150
rect 675759 192145 675825 192148
rect 675898 192146 675904 192148
rect 675968 192146 675974 192210
rect 42159 191764 42225 191767
rect 42490 191764 42496 191766
rect 42159 191762 42496 191764
rect 42159 191706 42164 191762
rect 42220 191706 42496 191762
rect 42159 191704 42496 191706
rect 42159 191701 42225 191704
rect 42490 191702 42496 191704
rect 42560 191702 42566 191766
rect 184527 191468 184593 191471
rect 184527 191466 190560 191468
rect 184527 191410 184532 191466
rect 184588 191410 190560 191466
rect 184527 191408 190560 191410
rect 184527 191405 184593 191408
rect 41775 191174 41841 191175
rect 41722 191172 41728 191174
rect 41684 191112 41728 191172
rect 41792 191170 41841 191174
rect 41836 191114 41841 191170
rect 41722 191110 41728 191112
rect 41792 191110 41841 191114
rect 41775 191109 41841 191110
rect 149391 191024 149457 191027
rect 143904 191022 149457 191024
rect 143904 190966 149396 191022
rect 149452 190966 149457 191022
rect 143904 190964 149457 190966
rect 149391 190961 149457 190964
rect 184623 190728 184689 190731
rect 184623 190726 190014 190728
rect 184623 190670 184628 190726
rect 184684 190670 190014 190726
rect 184623 190668 190014 190670
rect 184623 190665 184689 190668
rect 189954 190654 190014 190668
rect 189954 190594 190560 190654
rect 40570 190370 40576 190434
rect 40640 190432 40646 190434
rect 41775 190432 41841 190435
rect 40640 190430 41841 190432
rect 40640 190374 41780 190430
rect 41836 190374 41841 190430
rect 40640 190372 41841 190374
rect 40640 190370 40646 190372
rect 41775 190369 41841 190372
rect 184335 189988 184401 189991
rect 184335 189986 190560 189988
rect 184335 189930 184340 189986
rect 184396 189930 190560 189986
rect 184335 189928 190560 189930
rect 184335 189925 184401 189928
rect 147663 189840 147729 189843
rect 143904 189838 147729 189840
rect 143904 189782 147668 189838
rect 147724 189782 147729 189838
rect 143904 189780 147729 189782
rect 147663 189777 147729 189780
rect 184527 189248 184593 189251
rect 184527 189246 190014 189248
rect 184527 189190 184532 189246
rect 184588 189190 190014 189246
rect 184527 189188 190014 189190
rect 184527 189185 184593 189188
rect 189954 189174 190014 189188
rect 189954 189114 190560 189174
rect 42063 188064 42129 188067
rect 42682 188064 42688 188066
rect 42063 188062 42688 188064
rect 42063 188006 42068 188062
rect 42124 188006 42688 188062
rect 42063 188004 42688 188006
rect 42063 188001 42129 188004
rect 42682 188002 42688 188004
rect 42752 188002 42758 188066
rect 143874 188064 143934 188552
rect 184335 188508 184401 188511
rect 184335 188506 190560 188508
rect 184335 188450 184340 188506
rect 184396 188450 190560 188506
rect 184335 188448 190560 188450
rect 184335 188445 184401 188448
rect 639810 188182 639870 190106
rect 674554 189926 674560 189990
rect 674624 189988 674630 189990
rect 675471 189988 675537 189991
rect 674624 189986 675537 189988
rect 674624 189930 675476 189986
rect 675532 189930 675537 189986
rect 674624 189928 675537 189930
rect 674624 189926 674630 189928
rect 675471 189925 675537 189928
rect 675759 188510 675825 188511
rect 675706 188446 675712 188510
rect 675776 188508 675825 188510
rect 675776 188506 675868 188508
rect 675820 188450 675868 188506
rect 675776 188448 675868 188450
rect 675776 188446 675825 188448
rect 675759 188445 675825 188446
rect 149295 188064 149361 188067
rect 143874 188062 149361 188064
rect 143874 188006 149300 188062
rect 149356 188006 149361 188062
rect 143874 188004 149361 188006
rect 149295 188001 149361 188004
rect 184431 187620 184497 187623
rect 184431 187618 190560 187620
rect 184431 187562 184436 187618
rect 184492 187562 190560 187618
rect 184431 187560 190560 187562
rect 184431 187557 184497 187560
rect 149391 187472 149457 187475
rect 143904 187470 149457 187472
rect 143904 187414 149396 187470
rect 149452 187414 149457 187470
rect 143904 187412 149457 187414
rect 149391 187409 149457 187412
rect 41146 187114 41152 187178
rect 41216 187176 41222 187178
rect 41775 187176 41841 187179
rect 41216 187174 41841 187176
rect 41216 187118 41780 187174
rect 41836 187118 41841 187174
rect 41216 187116 41841 187118
rect 41216 187114 41222 187116
rect 41775 187113 41841 187116
rect 41338 186818 41344 186882
rect 41408 186880 41414 186882
rect 41775 186880 41841 186883
rect 41408 186878 41841 186880
rect 41408 186822 41780 186878
rect 41836 186822 41841 186878
rect 41408 186820 41841 186822
rect 41408 186818 41414 186820
rect 41775 186817 41841 186820
rect 184335 186880 184401 186883
rect 184335 186878 190560 186880
rect 184335 186822 184340 186878
rect 184396 186822 190560 186878
rect 184335 186820 190560 186822
rect 184335 186817 184401 186820
rect 149583 186288 149649 186291
rect 143904 186286 149649 186288
rect 143904 186230 149588 186286
rect 149644 186230 149649 186286
rect 143904 186228 149649 186230
rect 149583 186225 149649 186228
rect 185391 186140 185457 186143
rect 185391 186138 190560 186140
rect 185391 186082 185396 186138
rect 185452 186082 190560 186138
rect 185391 186080 190560 186082
rect 185391 186077 185457 186080
rect 40954 185930 40960 185994
rect 41024 185992 41030 185994
rect 41775 185992 41841 185995
rect 41024 185990 41841 185992
rect 41024 185934 41780 185990
rect 41836 185934 41841 185990
rect 41024 185932 41841 185934
rect 41024 185930 41030 185932
rect 41775 185929 41841 185932
rect 640194 185699 640254 186258
rect 640194 185694 640305 185699
rect 640194 185638 640244 185694
rect 640300 185638 640305 185694
rect 640194 185636 640305 185638
rect 640239 185633 640305 185636
rect 184431 185400 184497 185403
rect 184431 185398 190014 185400
rect 184431 185342 184436 185398
rect 184492 185342 190014 185398
rect 184431 185340 190014 185342
rect 184431 185337 184497 185340
rect 189954 185326 190014 185340
rect 189954 185266 190560 185326
rect 143874 184512 143934 185000
rect 640239 184956 640305 184959
rect 640194 184954 640305 184956
rect 640194 184898 640244 184954
rect 640300 184898 640305 184954
rect 640194 184893 640305 184898
rect 184527 184660 184593 184663
rect 184527 184658 190560 184660
rect 184527 184602 184532 184658
rect 184588 184602 190560 184658
rect 184527 184600 190560 184602
rect 184527 184597 184593 184600
rect 149199 184512 149265 184515
rect 143874 184510 149265 184512
rect 143874 184454 149204 184510
rect 149260 184454 149265 184510
rect 143874 184452 149265 184454
rect 149199 184449 149265 184452
rect 640194 184334 640254 184893
rect 42159 184218 42225 184219
rect 42106 184216 42112 184218
rect 42068 184156 42112 184216
rect 42176 184214 42225 184218
rect 42220 184158 42225 184214
rect 42106 184154 42112 184156
rect 42176 184154 42225 184158
rect 42159 184153 42225 184154
rect 184335 183920 184401 183923
rect 184335 183918 190014 183920
rect 184335 183862 184340 183918
rect 184396 183862 190014 183918
rect 184335 183860 190014 183862
rect 184335 183857 184401 183860
rect 189954 183846 190014 183860
rect 189954 183786 190560 183846
rect 149487 183772 149553 183775
rect 143904 183770 149553 183772
rect 143904 183714 149492 183770
rect 149548 183714 149553 183770
rect 143904 183712 149553 183714
rect 149487 183709 149553 183712
rect 40762 183562 40768 183626
rect 40832 183624 40838 183626
rect 41775 183624 41841 183627
rect 40832 183622 41841 183624
rect 40832 183566 41780 183622
rect 41836 183566 41841 183622
rect 40832 183564 41841 183566
rect 40832 183562 40838 183564
rect 41775 183561 41841 183564
rect 41871 183182 41937 183183
rect 41871 183178 41920 183182
rect 41984 183180 41990 183182
rect 184431 183180 184497 183183
rect 41871 183122 41876 183178
rect 41871 183118 41920 183122
rect 41984 183120 42028 183180
rect 184431 183178 190560 183180
rect 184431 183122 184436 183178
rect 184492 183122 190560 183178
rect 184431 183120 190560 183122
rect 41984 183118 41990 183120
rect 41871 183117 41937 183118
rect 184431 183117 184497 183120
rect 645135 183032 645201 183035
rect 640386 183030 645201 183032
rect 640386 182974 645140 183030
rect 645196 182974 645201 183030
rect 640386 182972 645201 182974
rect 149391 182588 149457 182591
rect 143904 182586 149457 182588
rect 143904 182530 149396 182586
rect 149452 182530 149457 182586
rect 143904 182528 149457 182530
rect 149391 182525 149457 182528
rect 186255 182440 186321 182443
rect 640386 182440 640446 182972
rect 645135 182969 645201 182972
rect 186255 182438 190014 182440
rect 186255 182382 186260 182438
rect 186316 182382 190014 182438
rect 640224 182410 640446 182440
rect 186255 182380 190014 182382
rect 186255 182377 186321 182380
rect 189954 182366 190014 182380
rect 640194 182380 640416 182410
rect 189954 182306 190560 182366
rect 184527 181552 184593 181555
rect 184527 181550 190560 181552
rect 184527 181494 184532 181550
rect 184588 181494 190560 181550
rect 184527 181492 190560 181494
rect 184527 181489 184593 181492
rect 149487 181404 149553 181407
rect 143904 181402 149553 181404
rect 143904 181346 149492 181402
rect 149548 181346 149553 181402
rect 143904 181344 149553 181346
rect 149487 181341 149553 181344
rect 184335 180812 184401 180815
rect 184335 180810 190560 180812
rect 184335 180754 184340 180810
rect 184396 180754 190560 180810
rect 184335 180752 190560 180754
rect 184335 180749 184401 180752
rect 640194 180560 640254 182380
rect 143874 179628 143934 180116
rect 184431 180072 184497 180075
rect 184431 180070 190560 180072
rect 184431 180014 184436 180070
rect 184492 180014 190560 180070
rect 184431 180012 190560 180014
rect 184431 180009 184497 180012
rect 149295 179628 149361 179631
rect 143874 179626 149361 179628
rect 143874 179570 149300 179626
rect 149356 179570 149361 179626
rect 143874 179568 149361 179570
rect 149295 179565 149361 179568
rect 184527 179332 184593 179335
rect 645135 179332 645201 179335
rect 184527 179330 190560 179332
rect 184527 179274 184532 179330
rect 184588 179274 190560 179330
rect 184527 179272 190560 179274
rect 640194 179330 645201 179332
rect 640194 179274 645140 179330
rect 645196 179274 645201 179330
rect 640194 179272 645201 179274
rect 184527 179269 184593 179272
rect 149391 178888 149457 178891
rect 143904 178886 149457 178888
rect 143904 178830 149396 178886
rect 149452 178830 149457 178886
rect 143904 178828 149457 178830
rect 149391 178825 149457 178828
rect 184623 178592 184689 178595
rect 184623 178590 190560 178592
rect 184623 178534 184628 178590
rect 184684 178534 190560 178590
rect 184623 178532 190560 178534
rect 184623 178529 184689 178532
rect 149487 177704 149553 177707
rect 143904 177702 149553 177704
rect 143904 177646 149492 177702
rect 149548 177646 149553 177702
rect 143904 177644 149553 177646
rect 149487 177641 149553 177644
rect 184335 177704 184401 177707
rect 184335 177702 190560 177704
rect 184335 177646 184340 177702
rect 184396 177646 190560 177702
rect 184335 177644 190560 177646
rect 184335 177641 184401 177644
rect 184431 177112 184497 177115
rect 184431 177110 190014 177112
rect 184431 177054 184436 177110
rect 184492 177054 190014 177110
rect 184431 177052 190014 177054
rect 184431 177049 184497 177052
rect 189954 177038 190014 177052
rect 189954 176978 190560 177038
rect 640194 176786 640254 179272
rect 645135 179269 645201 179272
rect 149391 176520 149457 176523
rect 143904 176518 149457 176520
rect 143904 176462 149396 176518
rect 149452 176462 149457 176518
rect 143904 176460 149457 176462
rect 149391 176457 149457 176460
rect 184527 176224 184593 176227
rect 184527 176222 190560 176224
rect 184527 176166 184532 176222
rect 184588 176166 190560 176222
rect 184527 176164 190560 176166
rect 184527 176161 184593 176164
rect 184335 175632 184401 175635
rect 184335 175630 190014 175632
rect 184335 175574 184340 175630
rect 184396 175574 190014 175630
rect 184335 175572 190014 175574
rect 184335 175569 184401 175572
rect 189954 175558 190014 175572
rect 189954 175498 190560 175558
rect 147759 175188 147825 175191
rect 143904 175186 147825 175188
rect 143904 175130 147764 175186
rect 147820 175130 147825 175186
rect 143904 175128 147825 175130
rect 147759 175125 147825 175128
rect 645135 174892 645201 174895
rect 640416 174890 645201 174892
rect 640416 174862 645140 174890
rect 640386 174834 645140 174862
rect 645196 174834 645201 174890
rect 640386 174832 645201 174834
rect 185871 174744 185937 174747
rect 185871 174742 190560 174744
rect 185871 174686 185876 174742
rect 185932 174686 190560 174742
rect 185871 174684 190560 174686
rect 185871 174681 185937 174684
rect 149103 174004 149169 174007
rect 143904 174002 149169 174004
rect 143904 173946 149108 174002
rect 149164 173946 149169 174002
rect 143904 173944 149169 173946
rect 149103 173941 149169 173944
rect 184431 174004 184497 174007
rect 184431 174002 190014 174004
rect 184431 173946 184436 174002
rect 184492 173946 190014 174002
rect 184431 173944 190014 173946
rect 184431 173941 184497 173944
rect 189954 173930 190014 173944
rect 189954 173870 190560 173930
rect 185679 173264 185745 173267
rect 185679 173262 190560 173264
rect 185679 173206 185684 173262
rect 185740 173206 190560 173262
rect 185679 173204 190560 173206
rect 185679 173201 185745 173204
rect 640386 172938 640446 174832
rect 645135 174829 645201 174832
rect 676143 173856 676209 173859
rect 676290 173856 676350 174122
rect 676143 173854 676350 173856
rect 676143 173798 676148 173854
rect 676204 173798 676350 173854
rect 676143 173796 676350 173798
rect 676143 173793 676209 173796
rect 676047 173560 676113 173563
rect 676047 173558 676320 173560
rect 676047 173502 676052 173558
rect 676108 173502 676320 173558
rect 676047 173500 676320 173502
rect 676047 173497 676113 173500
rect 676239 173264 676305 173267
rect 676239 173262 676350 173264
rect 676239 173206 676244 173262
rect 676300 173206 676350 173262
rect 676239 173201 676350 173206
rect 676290 172938 676350 173201
rect 149583 172820 149649 172823
rect 143904 172818 149649 172820
rect 143904 172762 149588 172818
rect 149644 172762 149649 172818
rect 143904 172760 149649 172762
rect 149583 172757 149649 172760
rect 673978 172758 673984 172822
rect 674048 172820 674054 172822
rect 674048 172760 676350 172820
rect 674048 172758 674054 172760
rect 676290 172568 676350 172760
rect 184335 172524 184401 172527
rect 184335 172522 190014 172524
rect 184335 172466 184340 172522
rect 184396 172466 190014 172522
rect 184335 172464 190014 172466
rect 184335 172461 184401 172464
rect 189954 172450 190014 172464
rect 189954 172390 190560 172450
rect 673978 172018 673984 172082
rect 674048 172080 674054 172082
rect 674048 172020 676320 172080
rect 674048 172018 674054 172020
rect 184527 171784 184593 171787
rect 184527 171782 190560 171784
rect 184527 171726 184532 171782
rect 184588 171726 190560 171782
rect 184527 171724 190560 171726
rect 184527 171721 184593 171724
rect 143874 171044 143934 171532
rect 674362 171426 674368 171490
rect 674432 171488 674438 171490
rect 674432 171428 676320 171488
rect 674432 171426 674438 171428
rect 149295 171044 149361 171047
rect 645135 171044 645201 171047
rect 143874 171042 149361 171044
rect 143874 170986 149300 171042
rect 149356 170986 149361 171042
rect 640416 171042 645201 171044
rect 640416 171014 645140 171042
rect 143874 170984 149361 170986
rect 149295 170981 149361 170984
rect 640386 170986 645140 171014
rect 645196 170986 645201 171042
rect 640386 170984 645201 170986
rect 184431 170896 184497 170899
rect 184431 170894 190560 170896
rect 184431 170838 184436 170894
rect 184492 170838 190560 170894
rect 184431 170836 190560 170838
rect 184431 170833 184497 170836
rect 149199 170304 149265 170307
rect 143904 170302 149265 170304
rect 143904 170246 149204 170302
rect 149260 170246 149265 170302
rect 143904 170244 149265 170246
rect 149199 170241 149265 170244
rect 184623 170304 184689 170307
rect 184623 170302 190014 170304
rect 184623 170246 184628 170302
rect 184684 170246 190014 170302
rect 184623 170244 190014 170246
rect 184623 170241 184689 170244
rect 189954 170230 190014 170244
rect 189954 170170 190560 170230
rect 184335 169416 184401 169419
rect 184335 169414 190560 169416
rect 184335 169358 184340 169414
rect 184396 169358 190560 169414
rect 184335 169356 190560 169358
rect 184335 169353 184401 169356
rect 148719 169120 148785 169123
rect 143904 169118 148785 169120
rect 143904 169062 148724 169118
rect 148780 169062 148785 169118
rect 640386 169090 640446 170984
rect 645135 170981 645201 170984
rect 672399 171044 672465 171047
rect 674362 171044 674368 171046
rect 672399 171042 674368 171044
rect 672399 170986 672404 171042
rect 672460 170986 674368 171042
rect 672399 170984 674368 170986
rect 672399 170981 672465 170984
rect 674362 170982 674368 170984
rect 674432 171044 674438 171046
rect 676290 171044 676350 171088
rect 674432 170984 676350 171044
rect 674432 170982 674438 170984
rect 674170 170538 674176 170602
rect 674240 170600 674246 170602
rect 674240 170540 676320 170600
rect 674240 170538 674246 170540
rect 676047 170008 676113 170011
rect 676047 170006 676320 170008
rect 676047 169950 676052 170006
rect 676108 169950 676320 170006
rect 676047 169948 676320 169950
rect 676047 169945 676113 169948
rect 676290 169270 676350 169534
rect 676282 169206 676288 169270
rect 676352 169206 676358 169270
rect 676047 169120 676113 169123
rect 676047 169118 676320 169120
rect 143904 169060 148785 169062
rect 148719 169057 148785 169060
rect 676047 169062 676052 169118
rect 676108 169062 676320 169118
rect 676047 169060 676320 169062
rect 676047 169057 676113 169060
rect 184527 168676 184593 168679
rect 184527 168674 190014 168676
rect 184527 168618 184532 168674
rect 184588 168618 190014 168674
rect 184527 168616 190014 168618
rect 184527 168613 184593 168616
rect 189954 168602 190014 168616
rect 676090 168614 676096 168678
rect 676160 168676 676166 168678
rect 676160 168616 676350 168676
rect 676160 168614 676166 168616
rect 189954 168542 190560 168602
rect 676290 168498 676350 168616
rect 148527 168084 148593 168087
rect 143904 168082 148593 168084
rect 143904 168026 148532 168082
rect 148588 168026 148593 168082
rect 143904 168024 148593 168026
rect 148527 168021 148593 168024
rect 675514 168022 675520 168086
rect 675584 168084 675590 168086
rect 675584 168024 676320 168084
rect 675584 168022 675590 168024
rect 184623 167936 184689 167939
rect 184623 167934 190560 167936
rect 184623 167878 184628 167934
rect 184684 167878 190560 167934
rect 184623 167876 190560 167878
rect 184623 167873 184689 167876
rect 645135 167788 645201 167791
rect 640386 167786 645201 167788
rect 640386 167730 645140 167786
rect 645196 167730 645201 167786
rect 640386 167728 645201 167730
rect 184431 167196 184497 167199
rect 184431 167194 190014 167196
rect 184431 167138 184436 167194
rect 184492 167138 190014 167194
rect 184431 167136 190014 167138
rect 184431 167133 184497 167136
rect 189954 167122 190014 167136
rect 189954 167062 190560 167122
rect 143874 166308 143934 166796
rect 184335 166456 184401 166459
rect 184335 166454 190560 166456
rect 184335 166398 184340 166454
rect 184396 166398 190560 166454
rect 184335 166396 190560 166398
rect 184335 166393 184401 166396
rect 148623 166308 148689 166311
rect 143874 166306 148689 166308
rect 143874 166250 148628 166306
rect 148684 166250 148689 166306
rect 143874 166248 148689 166250
rect 148623 166245 148689 166248
rect 640386 166012 640446 167728
rect 645135 167725 645201 167728
rect 674554 167282 674560 167346
rect 674624 167344 674630 167346
rect 676290 167344 676350 167536
rect 674624 167284 676350 167344
rect 674624 167282 674630 167284
rect 674362 166986 674368 167050
rect 674432 167048 674438 167050
rect 674432 166988 676320 167048
rect 674432 166986 674438 166988
rect 675706 166542 675712 166606
rect 675776 166604 675782 166606
rect 675776 166544 676320 166604
rect 675776 166542 675782 166544
rect 640194 165952 640446 166012
rect 184527 165716 184593 165719
rect 184527 165714 190014 165716
rect 184527 165658 184532 165714
rect 184588 165658 190014 165714
rect 184527 165656 190014 165658
rect 184527 165653 184593 165656
rect 189954 165642 190014 165656
rect 189954 165582 190560 165642
rect 148431 165568 148497 165571
rect 143904 165566 148497 165568
rect 143904 165510 148436 165566
rect 148492 165510 148497 165566
rect 143904 165508 148497 165510
rect 148431 165505 148497 165508
rect 640194 165242 640254 165952
rect 675322 165654 675328 165718
rect 675392 165716 675398 165718
rect 676290 165716 676350 166056
rect 675392 165656 676350 165716
rect 675392 165654 675398 165656
rect 675898 165506 675904 165570
rect 675968 165568 675974 165570
rect 675968 165508 676320 165568
rect 675968 165506 675974 165508
rect 674938 165062 674944 165126
rect 675008 165124 675014 165126
rect 675008 165064 676320 165124
rect 675008 165062 675014 165064
rect 184431 164828 184497 164831
rect 184431 164826 190560 164828
rect 184431 164770 184436 164826
rect 184492 164770 190560 164826
rect 184431 164768 190560 164770
rect 184431 164765 184497 164768
rect 674746 164470 674752 164534
rect 674816 164532 674822 164534
rect 674816 164472 676320 164532
rect 674816 164470 674822 164472
rect 148239 164384 148305 164387
rect 143904 164382 148305 164384
rect 143904 164326 148244 164382
rect 148300 164326 148305 164382
rect 143904 164324 148305 164326
rect 148239 164321 148305 164324
rect 184335 164088 184401 164091
rect 676047 164088 676113 164091
rect 184335 164086 190560 164088
rect 184335 164030 184340 164086
rect 184396 164030 190560 164086
rect 184335 164028 190560 164030
rect 676047 164086 676320 164088
rect 676047 164030 676052 164086
rect 676108 164030 676320 164086
rect 676047 164028 676320 164030
rect 184335 164025 184401 164028
rect 676047 164025 676113 164028
rect 675130 163582 675136 163646
rect 675200 163644 675206 163646
rect 675200 163584 676320 163644
rect 675200 163582 675206 163584
rect 184527 163348 184593 163351
rect 645135 163348 645201 163351
rect 184527 163346 190560 163348
rect 184527 163290 184532 163346
rect 184588 163290 190560 163346
rect 640416 163346 645201 163348
rect 640416 163318 645140 163346
rect 184527 163288 190560 163290
rect 640386 163290 645140 163318
rect 645196 163290 645201 163346
rect 640386 163288 645201 163290
rect 184527 163285 184593 163288
rect 148911 163200 148977 163203
rect 143904 163198 148977 163200
rect 143904 163142 148916 163198
rect 148972 163142 148977 163198
rect 143904 163140 148977 163142
rect 148911 163137 148977 163140
rect 184335 162608 184401 162611
rect 184335 162606 190560 162608
rect 184335 162550 184340 162606
rect 184396 162550 190560 162606
rect 184335 162548 190560 162550
rect 184335 162545 184401 162548
rect 148335 161868 148401 161871
rect 143904 161866 148401 161868
rect 143904 161810 148340 161866
rect 148396 161810 148401 161866
rect 143904 161808 148401 161810
rect 148335 161805 148401 161808
rect 184431 161868 184497 161871
rect 184431 161866 190560 161868
rect 184431 161810 184436 161866
rect 184492 161810 190560 161866
rect 184431 161808 190560 161810
rect 184431 161805 184497 161808
rect 640386 161394 640446 163288
rect 645135 163285 645201 163288
rect 676866 162758 676926 163022
rect 676858 162694 676864 162758
rect 676928 162694 676934 162758
rect 676290 162315 676350 162504
rect 676239 162310 676350 162315
rect 676239 162254 676244 162310
rect 676300 162254 676350 162310
rect 676239 162252 676350 162254
rect 676239 162249 676305 162252
rect 676143 161868 676209 161871
rect 676290 161868 676350 162134
rect 676143 161866 676350 161868
rect 676143 161810 676148 161866
rect 676204 161810 676350 161866
rect 676143 161808 676350 161810
rect 676143 161805 676209 161808
rect 676290 161427 676350 161542
rect 676239 161422 676350 161427
rect 676239 161366 676244 161422
rect 676300 161366 676350 161422
rect 676239 161364 676350 161366
rect 676239 161361 676305 161364
rect 184335 160980 184401 160983
rect 184335 160978 190560 160980
rect 184335 160922 184340 160978
rect 184396 160922 190560 160978
rect 184335 160920 190560 160922
rect 184335 160917 184401 160920
rect 148815 160684 148881 160687
rect 143904 160682 148881 160684
rect 143904 160626 148820 160682
rect 148876 160626 148881 160682
rect 143904 160624 148881 160626
rect 148815 160621 148881 160624
rect 184431 160388 184497 160391
rect 184431 160386 190014 160388
rect 184431 160330 184436 160386
rect 184492 160330 190014 160386
rect 184431 160328 190014 160330
rect 184431 160325 184497 160328
rect 189954 160314 190014 160328
rect 189954 160254 190560 160314
rect 147087 159500 147153 159503
rect 143904 159498 147153 159500
rect 143904 159442 147092 159498
rect 147148 159442 147153 159498
rect 143904 159440 147153 159442
rect 147087 159437 147153 159440
rect 184623 159500 184689 159503
rect 645135 159500 645201 159503
rect 184623 159498 190560 159500
rect 184623 159442 184628 159498
rect 184684 159442 190560 159498
rect 640416 159498 645201 159500
rect 640416 159470 645140 159498
rect 184623 159440 190560 159442
rect 640386 159442 645140 159470
rect 645196 159442 645201 159498
rect 640386 159440 645201 159442
rect 184623 159437 184689 159440
rect 184527 158908 184593 158911
rect 184527 158906 190014 158908
rect 184527 158850 184532 158906
rect 184588 158850 190014 158906
rect 184527 158848 190014 158850
rect 184527 158845 184593 158848
rect 189954 158834 190014 158848
rect 189954 158774 190560 158834
rect 143874 158020 143934 158212
rect 149391 158020 149457 158023
rect 143874 158018 149457 158020
rect 143874 157962 149396 158018
rect 149452 157962 149457 158018
rect 143874 157960 149457 157962
rect 149391 157957 149457 157960
rect 184335 158020 184401 158023
rect 184335 158018 190560 158020
rect 184335 157962 184340 158018
rect 184396 157962 190560 158018
rect 184335 157960 190560 157962
rect 184335 157957 184401 157960
rect 640386 157546 640446 159440
rect 645135 159437 645201 159440
rect 675759 158168 675825 158171
rect 676090 158168 676096 158170
rect 675759 158166 676096 158168
rect 675759 158110 675764 158166
rect 675820 158110 676096 158166
rect 675759 158108 676096 158110
rect 675759 158105 675825 158108
rect 676090 158106 676096 158108
rect 676160 158106 676166 158170
rect 675759 157726 675825 157727
rect 675706 157662 675712 157726
rect 675776 157724 675825 157726
rect 675776 157722 675868 157724
rect 675820 157666 675868 157722
rect 675776 157664 675868 157666
rect 675776 157662 675825 157664
rect 675759 157661 675825 157662
rect 184431 157428 184497 157431
rect 184431 157426 190014 157428
rect 184431 157370 184436 157426
rect 184492 157370 190014 157426
rect 184431 157368 190014 157370
rect 184431 157365 184497 157368
rect 189954 157354 190014 157368
rect 189954 157294 190560 157354
rect 147087 156984 147153 156987
rect 143904 156982 147153 156984
rect 143904 156926 147092 156982
rect 147148 156926 147153 156982
rect 143904 156924 147153 156926
rect 147087 156921 147153 156924
rect 675759 156984 675825 156987
rect 676282 156984 676288 156986
rect 675759 156982 676288 156984
rect 675759 156926 675764 156982
rect 675820 156926 676288 156982
rect 675759 156924 676288 156926
rect 675759 156921 675825 156924
rect 676282 156922 676288 156924
rect 676352 156922 676358 156986
rect 184623 156540 184689 156543
rect 184623 156538 190560 156540
rect 184623 156482 184628 156538
rect 184684 156482 190560 156538
rect 184623 156480 190560 156482
rect 184623 156477 184689 156480
rect 149391 155800 149457 155803
rect 143904 155798 149457 155800
rect 143904 155742 149396 155798
rect 149452 155742 149457 155798
rect 143904 155740 149457 155742
rect 149391 155737 149457 155740
rect 184527 155652 184593 155655
rect 184527 155650 190560 155652
rect 184527 155594 184532 155650
rect 184588 155594 190560 155650
rect 184527 155592 190560 155594
rect 184527 155589 184593 155592
rect 640194 155504 640254 155622
rect 645135 155504 645201 155507
rect 640194 155502 645201 155504
rect 640194 155446 645140 155502
rect 645196 155446 645201 155502
rect 640194 155444 645201 155446
rect 184527 155060 184593 155063
rect 184527 155058 190560 155060
rect 184527 155002 184532 155058
rect 184588 155002 190560 155058
rect 184527 155000 190560 155002
rect 184527 154997 184593 155000
rect 149487 154616 149553 154619
rect 143904 154614 149553 154616
rect 143904 154558 149492 154614
rect 149548 154558 149553 154614
rect 143904 154556 149553 154558
rect 149487 154553 149553 154556
rect 184335 154172 184401 154175
rect 184335 154170 190560 154172
rect 184335 154114 184340 154170
rect 184396 154114 190560 154170
rect 184335 154112 190560 154114
rect 184335 154109 184401 154112
rect 640386 153772 640446 155444
rect 645135 155441 645201 155444
rect 675471 155210 675537 155211
rect 675471 155206 675520 155210
rect 675584 155208 675590 155210
rect 675471 155150 675476 155206
rect 675471 155146 675520 155150
rect 675584 155148 675628 155208
rect 675584 155146 675590 155148
rect 675471 155145 675537 155146
rect 675375 154470 675441 154471
rect 675322 154468 675328 154470
rect 675284 154408 675328 154468
rect 675392 154466 675441 154470
rect 675436 154410 675441 154466
rect 675322 154406 675328 154408
rect 675392 154406 675441 154410
rect 675375 154405 675441 154406
rect 675759 153876 675825 153879
rect 675898 153876 675904 153878
rect 675759 153874 675904 153876
rect 675759 153818 675764 153874
rect 675820 153818 675904 153874
rect 675759 153816 675904 153818
rect 675759 153813 675825 153816
rect 675898 153814 675904 153816
rect 675968 153814 675974 153878
rect 184431 153580 184497 153583
rect 184431 153578 190014 153580
rect 184431 153522 184436 153578
rect 184492 153522 190014 153578
rect 184431 153520 190014 153522
rect 184431 153517 184497 153520
rect 189954 153506 190014 153520
rect 189954 153446 190560 153506
rect 143874 152988 143934 153328
rect 149391 152988 149457 152991
rect 143874 152986 149457 152988
rect 143874 152930 149396 152986
rect 149452 152930 149457 152986
rect 143874 152928 149457 152930
rect 149391 152925 149457 152928
rect 184623 152692 184689 152695
rect 675183 152692 675249 152695
rect 676858 152692 676864 152694
rect 184623 152690 190560 152692
rect 184623 152634 184628 152690
rect 184684 152634 190560 152690
rect 184623 152632 190560 152634
rect 675183 152690 676864 152692
rect 675183 152634 675188 152690
rect 675244 152634 676864 152690
rect 675183 152632 676864 152634
rect 184623 152629 184689 152632
rect 675183 152629 675249 152632
rect 676858 152630 676864 152632
rect 676928 152630 676934 152694
rect 645135 152544 645201 152547
rect 640194 152542 645201 152544
rect 640194 152486 645140 152542
rect 645196 152486 645201 152542
rect 640194 152484 645201 152486
rect 149679 152100 149745 152103
rect 143904 152098 149745 152100
rect 143904 152042 149684 152098
rect 149740 152042 149745 152098
rect 143904 152040 149745 152042
rect 149679 152037 149745 152040
rect 184335 151952 184401 151955
rect 184335 151950 190014 151952
rect 184335 151894 184340 151950
rect 184396 151894 190014 151950
rect 184335 151892 190014 151894
rect 184335 151889 184401 151892
rect 189954 151878 190014 151892
rect 189954 151818 190560 151878
rect 184431 151212 184497 151215
rect 184431 151210 190560 151212
rect 184431 151154 184436 151210
rect 184492 151154 190560 151210
rect 184431 151152 190560 151154
rect 184431 151149 184497 151152
rect 149487 150916 149553 150919
rect 143904 150914 149553 150916
rect 143904 150858 149492 150914
rect 149548 150858 149553 150914
rect 143904 150856 149553 150858
rect 149487 150853 149553 150856
rect 184527 150472 184593 150475
rect 184527 150470 190014 150472
rect 184527 150414 184532 150470
rect 184588 150414 190014 150470
rect 184527 150412 190014 150414
rect 184527 150409 184593 150412
rect 189954 150398 190014 150412
rect 189954 150338 190560 150398
rect 640194 149998 640254 152484
rect 645135 152481 645201 152484
rect 674554 150854 674560 150918
rect 674624 150916 674630 150918
rect 675375 150916 675441 150919
rect 674624 150914 675441 150916
rect 674624 150858 675380 150914
rect 675436 150858 675441 150914
rect 674624 150856 675441 150858
rect 674624 150854 674630 150856
rect 675375 150853 675441 150856
rect 675130 150262 675136 150326
rect 675200 150324 675206 150326
rect 675471 150324 675537 150327
rect 675200 150322 675537 150324
rect 675200 150266 675476 150322
rect 675532 150266 675537 150322
rect 675200 150264 675537 150266
rect 675200 150262 675206 150264
rect 675471 150261 675537 150264
rect 149391 149880 149457 149883
rect 143874 149878 149457 149880
rect 143874 149822 149396 149878
rect 149452 149822 149457 149878
rect 143874 149820 149457 149822
rect 143874 149776 143934 149820
rect 149391 149817 149457 149820
rect 184335 149732 184401 149735
rect 184335 149730 190560 149732
rect 184335 149674 184340 149730
rect 184396 149674 190560 149730
rect 184335 149672 190560 149674
rect 184335 149669 184401 149672
rect 674746 149522 674752 149586
rect 674816 149584 674822 149586
rect 675375 149584 675441 149587
rect 674816 149582 675441 149584
rect 674816 149526 675380 149582
rect 675436 149526 675441 149582
rect 674816 149524 675441 149526
rect 674816 149522 674822 149524
rect 675375 149521 675441 149524
rect 184431 148992 184497 148995
rect 184431 148990 190014 148992
rect 184431 148934 184436 148990
rect 184492 148934 190014 148990
rect 184431 148932 190014 148934
rect 184431 148929 184497 148932
rect 189954 148918 190014 148932
rect 189954 148858 190560 148918
rect 149487 148548 149553 148551
rect 143904 148546 149553 148548
rect 143904 148490 149492 148546
rect 149548 148490 149553 148546
rect 143904 148488 149553 148490
rect 149487 148485 149553 148488
rect 184335 148104 184401 148107
rect 645135 148104 645201 148107
rect 184335 148102 190560 148104
rect 184335 148046 184340 148102
rect 184396 148046 190560 148102
rect 640416 148102 645201 148104
rect 640416 148074 645140 148102
rect 184335 148044 190560 148046
rect 640386 148046 645140 148074
rect 645196 148046 645201 148102
rect 640386 148044 645201 148046
rect 184335 148041 184401 148044
rect 149391 147364 149457 147367
rect 143904 147362 149457 147364
rect 143904 147306 149396 147362
rect 149452 147306 149457 147362
rect 143904 147304 149457 147306
rect 149391 147301 149457 147304
rect 184527 147364 184593 147367
rect 184527 147362 190560 147364
rect 184527 147306 184532 147362
rect 184588 147306 190560 147362
rect 184527 147304 190560 147306
rect 184527 147301 184593 147304
rect 184335 146624 184401 146627
rect 184335 146622 190560 146624
rect 184335 146566 184340 146622
rect 184396 146566 190560 146622
rect 184335 146564 190560 146566
rect 184335 146561 184401 146564
rect 149487 146180 149553 146183
rect 143904 146178 149553 146180
rect 143904 146122 149492 146178
rect 149548 146122 149553 146178
rect 640386 146150 640446 148044
rect 645135 148041 645201 148044
rect 674938 147894 674944 147958
rect 675008 147956 675014 147958
rect 675375 147956 675441 147959
rect 675008 147954 675441 147956
rect 675008 147898 675380 147954
rect 675436 147898 675441 147954
rect 675008 147896 675441 147898
rect 675008 147894 675014 147896
rect 675375 147893 675441 147896
rect 143904 146120 149553 146122
rect 149487 146117 149553 146120
rect 186735 145884 186801 145887
rect 186735 145882 190560 145884
rect 186735 145826 186740 145882
rect 186796 145826 190560 145882
rect 186735 145824 190560 145826
rect 186735 145821 186801 145824
rect 184431 145144 184497 145147
rect 184431 145142 190014 145144
rect 184431 145086 184436 145142
rect 184492 145086 190014 145142
rect 184431 145084 190014 145086
rect 184431 145081 184497 145084
rect 189954 145070 190014 145084
rect 189954 145010 190560 145070
rect 143874 144552 143934 144892
rect 149391 144552 149457 144555
rect 143874 144550 149457 144552
rect 143874 144494 149396 144550
rect 149452 144494 149457 144550
rect 143874 144492 149457 144494
rect 149391 144489 149457 144492
rect 184527 144404 184593 144407
rect 184527 144402 190560 144404
rect 184527 144346 184532 144402
rect 184588 144346 190560 144402
rect 184527 144344 190560 144346
rect 184527 144341 184593 144344
rect 646671 144256 646737 144259
rect 640416 144254 646737 144256
rect 640416 144226 646676 144254
rect 640386 144198 646676 144226
rect 646732 144198 646737 144254
rect 640386 144196 646737 144198
rect 149487 143664 149553 143667
rect 143904 143662 149553 143664
rect 143904 143606 149492 143662
rect 149548 143606 149553 143662
rect 143904 143604 149553 143606
rect 149487 143601 149553 143604
rect 185391 143664 185457 143667
rect 185391 143662 190014 143664
rect 185391 143606 185396 143662
rect 185452 143606 190014 143662
rect 185391 143604 190014 143606
rect 185391 143601 185457 143604
rect 189954 143590 190014 143604
rect 189954 143530 190560 143590
rect 184335 142776 184401 142779
rect 184335 142774 190560 142776
rect 184335 142718 184340 142774
rect 184396 142718 190560 142774
rect 184335 142716 190560 142718
rect 184335 142713 184401 142716
rect 149391 142480 149457 142483
rect 143904 142478 149457 142480
rect 143904 142422 149396 142478
rect 149452 142422 149457 142478
rect 143904 142420 149457 142422
rect 149391 142417 149457 142420
rect 640386 142302 640446 144196
rect 646671 144193 646737 144196
rect 674362 143898 674368 143962
rect 674432 143960 674438 143962
rect 675471 143960 675537 143963
rect 674432 143958 675537 143960
rect 674432 143902 675476 143958
rect 675532 143902 675537 143958
rect 674432 143900 675537 143902
rect 674432 143898 674438 143900
rect 675471 143897 675537 143900
rect 184431 142184 184497 142187
rect 184431 142182 190014 142184
rect 184431 142126 184436 142182
rect 184492 142126 190014 142182
rect 184431 142124 190014 142126
rect 184431 142121 184497 142124
rect 189954 142110 190014 142124
rect 189954 142050 190560 142110
rect 147087 141296 147153 141299
rect 143904 141294 147153 141296
rect 143904 141238 147092 141294
rect 147148 141238 147153 141294
rect 143904 141236 147153 141238
rect 147087 141233 147153 141236
rect 184527 141296 184593 141299
rect 184527 141294 190560 141296
rect 184527 141238 184532 141294
rect 184588 141238 190560 141294
rect 184527 141236 190560 141238
rect 184527 141233 184593 141236
rect 646767 141000 646833 141003
rect 640386 140998 646833 141000
rect 640386 140942 646772 140998
rect 646828 140942 646833 140998
rect 640386 140940 646833 140942
rect 184335 140556 184401 140559
rect 184335 140554 190560 140556
rect 184335 140498 184340 140554
rect 184396 140498 190560 140554
rect 184335 140496 190560 140498
rect 184335 140493 184401 140496
rect 640386 140408 640446 140940
rect 646767 140937 646833 140940
rect 640224 140378 640446 140408
rect 640194 140348 640416 140378
rect 146895 139964 146961 139967
rect 143904 139962 146961 139964
rect 143904 139906 146900 139962
rect 146956 139906 146961 139962
rect 143904 139904 146961 139906
rect 146895 139901 146961 139904
rect 184431 139816 184497 139819
rect 184431 139814 190560 139816
rect 184431 139758 184436 139814
rect 184492 139758 190560 139814
rect 184431 139756 190560 139758
rect 184431 139753 184497 139756
rect 184527 138928 184593 138931
rect 184527 138926 190560 138928
rect 184527 138870 184532 138926
rect 184588 138870 190560 138926
rect 184527 138868 190560 138870
rect 184527 138865 184593 138868
rect 149391 138780 149457 138783
rect 143904 138778 149457 138780
rect 143904 138722 149396 138778
rect 149452 138722 149457 138778
rect 143904 138720 149457 138722
rect 149391 138717 149457 138720
rect 640194 138528 640254 140348
rect 184623 138336 184689 138339
rect 184623 138334 190560 138336
rect 184623 138278 184628 138334
rect 184684 138278 190560 138334
rect 184623 138276 190560 138278
rect 184623 138273 184689 138276
rect 149679 137596 149745 137599
rect 143904 137594 149745 137596
rect 143904 137538 149684 137594
rect 149740 137538 149745 137594
rect 143904 137536 149745 137538
rect 149679 137533 149745 137536
rect 186159 137448 186225 137451
rect 186159 137446 190560 137448
rect 186159 137390 186164 137446
rect 186220 137390 190560 137446
rect 186159 137388 190560 137390
rect 186159 137385 186225 137388
rect 185967 136856 186033 136859
rect 185967 136854 190014 136856
rect 185967 136798 185972 136854
rect 186028 136798 190014 136854
rect 185967 136796 190014 136798
rect 185967 136793 186033 136796
rect 189954 136782 190014 136796
rect 189954 136722 190560 136782
rect 143874 135968 143934 136308
rect 149391 135968 149457 135971
rect 143874 135966 149457 135968
rect 143874 135910 149396 135966
rect 149452 135910 149457 135966
rect 143874 135908 149457 135910
rect 149391 135905 149457 135908
rect 185775 135968 185841 135971
rect 185775 135966 190560 135968
rect 185775 135910 185780 135966
rect 185836 135910 190560 135966
rect 185775 135908 190560 135910
rect 185775 135905 185841 135908
rect 186255 135228 186321 135231
rect 186255 135226 190014 135228
rect 186255 135170 186260 135226
rect 186316 135170 190014 135226
rect 186255 135168 190014 135170
rect 186255 135165 186321 135168
rect 189954 135154 190014 135168
rect 189954 135094 190560 135154
rect 149391 135080 149457 135083
rect 143904 135078 149457 135080
rect 143904 135022 149396 135078
rect 149452 135022 149457 135078
rect 143904 135020 149457 135022
rect 149391 135017 149457 135020
rect 647055 134784 647121 134787
rect 640416 134782 647121 134784
rect 640416 134726 647060 134782
rect 647116 134726 647121 134782
rect 640416 134724 647121 134726
rect 647055 134721 647121 134724
rect 184431 134488 184497 134491
rect 184431 134486 190560 134488
rect 184431 134430 184436 134486
rect 184492 134430 190560 134486
rect 184431 134428 190560 134430
rect 184431 134425 184497 134428
rect 148815 133896 148881 133899
rect 143904 133894 148881 133896
rect 143904 133838 148820 133894
rect 148876 133838 148881 133894
rect 143904 133836 148881 133838
rect 148815 133833 148881 133836
rect 184527 133748 184593 133751
rect 184527 133746 190014 133748
rect 184527 133690 184532 133746
rect 184588 133690 190014 133746
rect 184527 133688 190014 133690
rect 184527 133685 184593 133688
rect 189954 133674 190014 133688
rect 189954 133614 190560 133674
rect 184335 133008 184401 133011
rect 184335 133006 190560 133008
rect 184335 132950 184340 133006
rect 184396 132950 190560 133006
rect 184335 132948 190560 132950
rect 184335 132945 184401 132948
rect 149007 132712 149073 132715
rect 143904 132710 149073 132712
rect 143904 132654 149012 132710
rect 149068 132654 149073 132710
rect 143904 132652 149073 132654
rect 149007 132649 149073 132652
rect 184335 132268 184401 132271
rect 184335 132266 190014 132268
rect 184335 132210 184340 132266
rect 184396 132210 190014 132266
rect 184335 132208 190014 132210
rect 184335 132205 184401 132208
rect 189954 132194 190014 132208
rect 189954 132134 190560 132194
rect 184431 131528 184497 131531
rect 184431 131526 190560 131528
rect 184431 131470 184436 131526
rect 184492 131470 190560 131526
rect 184431 131468 190560 131470
rect 184431 131465 184497 131468
rect 143874 130936 143934 131424
rect 149295 130936 149361 130939
rect 647727 130936 647793 130939
rect 143874 130934 149361 130936
rect 143874 130878 149300 130934
rect 149356 130878 149361 130934
rect 143874 130876 149361 130878
rect 640416 130934 647793 130936
rect 640416 130878 647732 130934
rect 647788 130878 647793 130934
rect 640416 130876 647793 130878
rect 149295 130873 149361 130876
rect 647727 130873 647793 130876
rect 184527 130640 184593 130643
rect 184527 130638 190560 130640
rect 184527 130582 184532 130638
rect 184588 130582 190560 130638
rect 184527 130580 190560 130582
rect 184527 130577 184593 130580
rect 149391 130344 149457 130347
rect 143904 130342 149457 130344
rect 143904 130286 149396 130342
rect 149452 130286 149457 130342
rect 143904 130284 149457 130286
rect 149391 130281 149457 130284
rect 184623 129900 184689 129903
rect 184623 129898 190560 129900
rect 184623 129842 184628 129898
rect 184684 129842 190560 129898
rect 184623 129840 190560 129842
rect 184623 129837 184689 129840
rect 676290 129607 676350 129870
rect 676239 129602 676350 129607
rect 676239 129546 676244 129602
rect 676300 129546 676350 129602
rect 676239 129544 676350 129546
rect 676239 129541 676305 129544
rect 676290 129163 676350 129278
rect 149103 129160 149169 129163
rect 143904 129158 149169 129160
rect 143904 129102 149108 129158
rect 149164 129102 149169 129158
rect 143904 129100 149169 129102
rect 149103 129097 149169 129100
rect 184335 129160 184401 129163
rect 184335 129158 190560 129160
rect 184335 129102 184340 129158
rect 184396 129102 190560 129158
rect 184335 129100 190560 129102
rect 676290 129158 676401 129163
rect 676290 129102 676340 129158
rect 676396 129102 676401 129158
rect 676290 129100 676401 129102
rect 184335 129097 184401 129100
rect 676335 129097 676401 129100
rect 647919 129012 647985 129015
rect 640416 129010 647985 129012
rect 640416 128954 647924 129010
rect 647980 128954 647985 129010
rect 640416 128952 647985 128954
rect 647919 128949 647985 128952
rect 676290 128571 676350 128834
rect 676239 128566 676350 128571
rect 676239 128510 676244 128566
rect 676300 128510 676350 128566
rect 676239 128508 676350 128510
rect 676239 128505 676305 128508
rect 184431 128420 184497 128423
rect 184431 128418 190014 128420
rect 184431 128362 184436 128418
rect 184492 128362 190014 128418
rect 184431 128360 190014 128362
rect 184431 128357 184497 128360
rect 189954 128346 190014 128360
rect 673978 128358 673984 128422
rect 674048 128420 674054 128422
rect 674048 128360 676320 128420
rect 674048 128358 674054 128360
rect 189954 128286 190560 128346
rect 149391 127976 149457 127979
rect 143904 127974 149457 127976
rect 143904 127918 149396 127974
rect 149452 127918 149457 127974
rect 143904 127916 149457 127918
rect 149391 127913 149457 127916
rect 184527 127680 184593 127683
rect 646959 127680 647025 127683
rect 184527 127678 190560 127680
rect 184527 127622 184532 127678
rect 184588 127622 190560 127678
rect 184527 127620 190560 127622
rect 640386 127678 647025 127680
rect 640386 127622 646964 127678
rect 647020 127622 647025 127678
rect 640386 127620 647025 127622
rect 184527 127617 184593 127620
rect 640386 127058 640446 127620
rect 646959 127617 647025 127620
rect 676143 127532 676209 127535
rect 676290 127532 676350 127798
rect 676143 127530 676350 127532
rect 676143 127474 676148 127530
rect 676204 127474 676350 127530
rect 676143 127472 676350 127474
rect 676143 127469 676209 127472
rect 674170 127322 674176 127386
rect 674240 127384 674246 127386
rect 674240 127324 676350 127384
rect 674240 127322 674246 127324
rect 676290 127280 676350 127324
rect 184623 126940 184689 126943
rect 676047 126940 676113 126943
rect 184623 126938 190014 126940
rect 184623 126882 184628 126938
rect 184684 126882 190014 126938
rect 184623 126880 190014 126882
rect 184623 126877 184689 126880
rect 189954 126866 190014 126880
rect 676047 126938 676320 126940
rect 676047 126882 676052 126938
rect 676108 126882 676320 126938
rect 676047 126880 676320 126882
rect 676047 126877 676113 126880
rect 189954 126806 190560 126866
rect 149295 126644 149361 126647
rect 143904 126642 149361 126644
rect 143904 126586 149300 126642
rect 149356 126586 149361 126642
rect 143904 126584 149361 126586
rect 149295 126581 149361 126584
rect 676047 126348 676113 126351
rect 676047 126346 676320 126348
rect 676047 126290 676052 126346
rect 676108 126290 676320 126346
rect 676047 126288 676320 126290
rect 676047 126285 676113 126288
rect 184335 126052 184401 126055
rect 184335 126050 190560 126052
rect 184335 125994 184340 126050
rect 184396 125994 190560 126050
rect 184335 125992 190560 125994
rect 184335 125989 184401 125992
rect 646863 125756 646929 125759
rect 640386 125754 646929 125756
rect 640386 125698 646868 125754
rect 646924 125698 646929 125754
rect 640386 125696 646929 125698
rect 149583 125460 149649 125463
rect 143904 125458 149649 125460
rect 143904 125402 149588 125458
rect 149644 125402 149649 125458
rect 143904 125400 149649 125402
rect 149583 125397 149649 125400
rect 184431 125460 184497 125463
rect 184431 125458 190014 125460
rect 184431 125402 184436 125458
rect 184492 125402 190014 125458
rect 184431 125400 190014 125402
rect 184431 125397 184497 125400
rect 189954 125386 190014 125400
rect 189954 125326 190560 125386
rect 640386 125208 640446 125696
rect 646863 125693 646929 125696
rect 676290 125611 676350 125800
rect 676239 125606 676350 125611
rect 676239 125550 676244 125606
rect 676300 125550 676350 125606
rect 676239 125548 676350 125550
rect 676239 125545 676305 125548
rect 675514 125398 675520 125462
rect 675584 125460 675590 125462
rect 675584 125400 676320 125460
rect 675584 125398 675590 125400
rect 676866 124575 676926 124838
rect 184527 124572 184593 124575
rect 184527 124570 190560 124572
rect 184527 124514 184532 124570
rect 184588 124514 190560 124570
rect 184527 124512 190560 124514
rect 676815 124570 676926 124575
rect 676815 124514 676820 124570
rect 676876 124514 676926 124570
rect 676815 124512 676926 124514
rect 184527 124509 184593 124512
rect 676815 124509 676881 124512
rect 148431 124276 148497 124279
rect 143904 124274 148497 124276
rect 143904 124218 148436 124274
rect 148492 124218 148497 124274
rect 143904 124216 148497 124218
rect 148431 124213 148497 124216
rect 676047 124276 676113 124279
rect 676047 124274 676320 124276
rect 676047 124218 676052 124274
rect 676108 124218 676320 124274
rect 676047 124216 676320 124218
rect 676047 124213 676113 124216
rect 675898 123844 675904 123908
rect 675968 123906 675974 123908
rect 675968 123846 676320 123906
rect 675968 123844 675974 123846
rect 184335 123832 184401 123835
rect 646575 123832 646641 123835
rect 184335 123830 190560 123832
rect 184335 123774 184340 123830
rect 184396 123774 190560 123830
rect 184335 123772 190560 123774
rect 640194 123830 646641 123832
rect 640194 123774 646580 123830
rect 646636 123774 646641 123830
rect 640194 123772 646641 123774
rect 184335 123769 184401 123772
rect 640194 123358 640254 123772
rect 646575 123769 646641 123772
rect 674170 123326 674176 123390
rect 674240 123388 674246 123390
rect 674240 123328 676320 123388
rect 674240 123326 674246 123328
rect 184431 123092 184497 123095
rect 184431 123090 190560 123092
rect 184431 123034 184436 123090
rect 184492 123034 190560 123090
rect 184431 123032 190560 123034
rect 184431 123029 184497 123032
rect 143874 122500 143934 122988
rect 679746 122651 679806 122766
rect 679695 122646 679806 122651
rect 679695 122590 679700 122646
rect 679756 122590 679806 122646
rect 679695 122588 679806 122590
rect 679695 122585 679761 122588
rect 148527 122500 148593 122503
rect 143874 122498 148593 122500
rect 143874 122442 148532 122498
rect 148588 122442 148593 122498
rect 143874 122440 148593 122442
rect 148527 122437 148593 122440
rect 676047 122426 676113 122429
rect 676047 122424 676320 122426
rect 676047 122368 676052 122424
rect 676108 122368 676320 122424
rect 676047 122366 676320 122368
rect 676047 122363 676113 122366
rect 184623 122204 184689 122207
rect 184623 122202 190560 122204
rect 184623 122146 184628 122202
rect 184684 122146 190560 122202
rect 184623 122144 190560 122146
rect 184623 122141 184689 122144
rect 646479 122056 646545 122059
rect 640194 122054 646545 122056
rect 640194 121998 646484 122054
rect 646540 121998 646545 122054
rect 640194 121996 646545 121998
rect 148719 121760 148785 121763
rect 143904 121758 148785 121760
rect 143904 121702 148724 121758
rect 148780 121702 148785 121758
rect 143904 121700 148785 121702
rect 148719 121697 148785 121700
rect 184527 121612 184593 121615
rect 184527 121610 190560 121612
rect 184527 121554 184532 121610
rect 184588 121554 190560 121610
rect 184527 121552 190560 121554
rect 184527 121549 184593 121552
rect 640194 121434 640254 121996
rect 646479 121993 646545 121996
rect 675951 121908 676017 121911
rect 675951 121906 676320 121908
rect 675951 121850 675956 121906
rect 676012 121850 676320 121906
rect 675951 121848 676320 121850
rect 675951 121845 676017 121848
rect 676290 121171 676350 121286
rect 676239 121166 676350 121171
rect 676239 121110 676244 121166
rect 676300 121110 676350 121166
rect 676239 121108 676350 121110
rect 676239 121105 676305 121108
rect 675706 120810 675712 120874
rect 675776 120872 675782 120874
rect 675776 120812 676320 120872
rect 675776 120810 675782 120812
rect 184431 120724 184497 120727
rect 184431 120722 190560 120724
rect 184431 120666 184436 120722
rect 184492 120666 190560 120722
rect 184431 120664 190560 120666
rect 184431 120661 184497 120664
rect 149391 120576 149457 120579
rect 143904 120574 149457 120576
rect 143904 120518 149396 120574
rect 149452 120518 149457 120574
rect 143904 120516 149457 120518
rect 149391 120513 149457 120516
rect 676047 120428 676113 120431
rect 676047 120426 676320 120428
rect 676047 120370 676052 120426
rect 676108 120370 676320 120426
rect 676047 120368 676320 120370
rect 676047 120365 676113 120368
rect 184527 120132 184593 120135
rect 184527 120130 190014 120132
rect 184527 120074 184532 120130
rect 184588 120074 190014 120130
rect 184527 120072 190014 120074
rect 184527 120069 184593 120072
rect 189954 120058 190014 120072
rect 189954 119998 190560 120058
rect 676047 119836 676113 119839
rect 676047 119834 676320 119836
rect 676047 119778 676052 119834
rect 676108 119778 676320 119834
rect 676047 119776 676320 119778
rect 676047 119773 676113 119776
rect 647823 119540 647889 119543
rect 640416 119538 647889 119540
rect 640416 119482 647828 119538
rect 647884 119482 647889 119538
rect 640416 119480 647889 119482
rect 647823 119477 647889 119480
rect 149487 119392 149553 119395
rect 143904 119390 149553 119392
rect 143904 119334 149492 119390
rect 149548 119334 149553 119390
rect 143904 119332 149553 119334
rect 149487 119329 149553 119332
rect 676290 119247 676350 119362
rect 184335 119244 184401 119247
rect 184335 119242 190560 119244
rect 184335 119186 184340 119242
rect 184396 119186 190560 119242
rect 184335 119184 190560 119186
rect 676239 119242 676350 119247
rect 676239 119186 676244 119242
rect 676300 119186 676350 119242
rect 676239 119184 676350 119186
rect 184335 119181 184401 119184
rect 676239 119181 676305 119184
rect 675951 118874 676017 118877
rect 675951 118872 676320 118874
rect 675951 118816 675956 118872
rect 676012 118816 676320 118872
rect 675951 118814 676320 118816
rect 675951 118811 676017 118814
rect 184623 118652 184689 118655
rect 184623 118650 190014 118652
rect 184623 118594 184628 118650
rect 184684 118594 190014 118650
rect 184623 118592 190014 118594
rect 184623 118589 184689 118592
rect 189954 118578 190014 118592
rect 189954 118518 190560 118578
rect 676239 118504 676305 118507
rect 676239 118502 676350 118504
rect 676239 118446 676244 118502
rect 676300 118446 676350 118502
rect 676239 118441 676350 118446
rect 676290 118326 676350 118441
rect 149391 118208 149457 118211
rect 143874 118206 149457 118208
rect 143874 118150 149396 118206
rect 149452 118150 149457 118206
rect 143874 118148 149457 118150
rect 143874 118104 143934 118148
rect 149391 118145 149457 118148
rect 184335 117764 184401 117767
rect 676143 117764 676209 117767
rect 676290 117764 676350 117882
rect 184335 117762 190560 117764
rect 184335 117706 184340 117762
rect 184396 117706 190560 117762
rect 184335 117704 190560 117706
rect 676143 117762 676350 117764
rect 676143 117706 676148 117762
rect 676204 117706 676350 117762
rect 676143 117704 676350 117706
rect 184335 117701 184401 117704
rect 676143 117701 676209 117704
rect 646191 117616 646257 117619
rect 640416 117614 646257 117616
rect 640416 117558 646196 117614
rect 646252 117558 646257 117614
rect 640416 117556 646257 117558
rect 646191 117553 646257 117556
rect 676290 117175 676350 117364
rect 676239 117170 676350 117175
rect 676239 117114 676244 117170
rect 676300 117114 676350 117170
rect 676239 117112 676350 117114
rect 676239 117109 676305 117112
rect 184431 117024 184497 117027
rect 184431 117022 190014 117024
rect 184431 116966 184436 117022
rect 184492 116966 190014 117022
rect 184431 116964 190014 116966
rect 184431 116961 184497 116964
rect 189954 116950 190014 116964
rect 189954 116890 190560 116950
rect 149487 116876 149553 116879
rect 143904 116874 149553 116876
rect 143904 116818 149492 116874
rect 149548 116818 149553 116874
rect 143904 116816 149553 116818
rect 149487 116813 149553 116816
rect 184527 116284 184593 116287
rect 184527 116282 190560 116284
rect 184527 116226 184532 116282
rect 184588 116226 190560 116282
rect 184527 116224 190560 116226
rect 184527 116221 184593 116224
rect 149391 115692 149457 115695
rect 647919 115692 647985 115695
rect 143904 115690 149457 115692
rect 143904 115634 149396 115690
rect 149452 115634 149457 115690
rect 143904 115632 149457 115634
rect 640416 115690 647985 115692
rect 640416 115634 647924 115690
rect 647980 115634 647985 115690
rect 640416 115632 647985 115634
rect 149391 115629 149457 115632
rect 647919 115629 647985 115632
rect 676474 115630 676480 115694
rect 676544 115692 676550 115694
rect 676815 115692 676881 115695
rect 676544 115690 676881 115692
rect 676544 115634 676820 115690
rect 676876 115634 676881 115690
rect 676544 115632 676881 115634
rect 676544 115630 676550 115632
rect 676815 115629 676881 115632
rect 184623 115396 184689 115399
rect 184623 115394 190560 115396
rect 184623 115338 184628 115394
rect 184684 115338 190560 115394
rect 184623 115336 190560 115338
rect 184623 115333 184689 115336
rect 148815 115248 148881 115251
rect 149391 115248 149457 115251
rect 148815 115246 149457 115248
rect 148815 115190 148820 115246
rect 148876 115190 149396 115246
rect 149452 115190 149457 115246
rect 148815 115188 149457 115190
rect 148815 115185 148881 115188
rect 149391 115185 149457 115188
rect 676666 115186 676672 115250
rect 676736 115248 676742 115250
rect 679695 115248 679761 115251
rect 676736 115246 679761 115248
rect 676736 115190 679700 115246
rect 679756 115190 679761 115246
rect 676736 115188 679761 115190
rect 676736 115186 676742 115188
rect 679695 115185 679761 115188
rect 184335 114804 184401 114807
rect 184335 114802 190560 114804
rect 184335 114746 184340 114802
rect 184396 114746 190560 114802
rect 184335 114744 190560 114746
rect 184335 114741 184401 114744
rect 149487 114508 149553 114511
rect 143904 114506 149553 114508
rect 143904 114450 149492 114506
rect 149548 114450 149553 114506
rect 143904 114448 149553 114450
rect 149487 114445 149553 114448
rect 184431 113916 184497 113919
rect 184431 113914 190560 113916
rect 184431 113858 184436 113914
rect 184492 113858 190560 113914
rect 184431 113856 190560 113858
rect 184431 113853 184497 113856
rect 149391 113176 149457 113179
rect 143904 113174 149457 113176
rect 143904 113118 149396 113174
rect 149452 113118 149457 113174
rect 143904 113116 149457 113118
rect 149391 113113 149457 113116
rect 184623 113176 184689 113179
rect 640194 113176 640254 113738
rect 646575 113176 646641 113179
rect 184623 113174 190560 113176
rect 184623 113118 184628 113174
rect 184684 113118 190560 113174
rect 184623 113116 190560 113118
rect 640194 113174 646641 113176
rect 640194 113118 646580 113174
rect 646636 113118 646641 113174
rect 640194 113116 646641 113118
rect 184623 113113 184689 113116
rect 646575 113113 646641 113116
rect 184527 112436 184593 112439
rect 184527 112434 190560 112436
rect 184527 112378 184532 112434
rect 184588 112378 190560 112434
rect 184527 112376 190560 112378
rect 184527 112373 184593 112376
rect 675567 112142 675633 112143
rect 675514 112078 675520 112142
rect 675584 112140 675633 112142
rect 675584 112138 675676 112140
rect 675628 112082 675676 112138
rect 675584 112080 675676 112082
rect 675584 112078 675633 112080
rect 675567 112077 675633 112078
rect 148719 111992 148785 111995
rect 143904 111990 148785 111992
rect 143904 111934 148724 111990
rect 148780 111934 148785 111990
rect 143904 111932 148785 111934
rect 148719 111929 148785 111932
rect 184335 111696 184401 111699
rect 184335 111694 190014 111696
rect 184335 111638 184340 111694
rect 184396 111638 190014 111694
rect 184335 111636 190014 111638
rect 184335 111633 184401 111636
rect 189954 111622 190014 111636
rect 189954 111562 190560 111622
rect 640386 111400 640446 111888
rect 647151 111400 647217 111403
rect 640386 111398 647217 111400
rect 640386 111342 647156 111398
rect 647212 111342 647217 111398
rect 640386 111340 647217 111342
rect 647151 111337 647217 111340
rect 148335 110956 148401 110959
rect 143904 110954 148401 110956
rect 143904 110898 148340 110954
rect 148396 110898 148401 110954
rect 143904 110896 148401 110898
rect 148335 110893 148401 110896
rect 184527 110956 184593 110959
rect 675759 110956 675825 110959
rect 675898 110956 675904 110958
rect 184527 110954 190560 110956
rect 184527 110898 184532 110954
rect 184588 110898 190560 110954
rect 184527 110896 190560 110898
rect 675759 110954 675904 110956
rect 675759 110898 675764 110954
rect 675820 110898 675904 110954
rect 675759 110896 675904 110898
rect 184527 110893 184593 110896
rect 675759 110893 675825 110896
rect 675898 110894 675904 110896
rect 675968 110894 675974 110958
rect 185679 110216 185745 110219
rect 185679 110214 190014 110216
rect 185679 110158 185684 110214
rect 185740 110158 190014 110214
rect 185679 110156 190014 110158
rect 185679 110153 185745 110156
rect 189954 110142 190014 110156
rect 189954 110082 190560 110142
rect 143874 109624 143934 109668
rect 149391 109624 149457 109627
rect 143874 109622 149457 109624
rect 143874 109566 149396 109622
rect 149452 109566 149457 109622
rect 143874 109564 149457 109566
rect 149391 109561 149457 109564
rect 640386 109476 640446 109890
rect 646671 109476 646737 109479
rect 640386 109474 646737 109476
rect 640386 109418 646676 109474
rect 646732 109418 646737 109474
rect 640386 109416 646737 109418
rect 646671 109413 646737 109416
rect 185295 109328 185361 109331
rect 185295 109326 190560 109328
rect 185295 109270 185300 109326
rect 185356 109270 190560 109326
rect 185295 109268 190560 109270
rect 185295 109265 185361 109268
rect 186255 108736 186321 108739
rect 186255 108734 190014 108736
rect 186255 108678 186260 108734
rect 186316 108678 190014 108734
rect 186255 108676 190014 108678
rect 186255 108673 186321 108676
rect 189954 108662 190014 108676
rect 189954 108602 190560 108662
rect 147855 108440 147921 108443
rect 143904 108438 147921 108440
rect 143904 108382 147860 108438
rect 147916 108382 147921 108438
rect 143904 108380 147921 108382
rect 147855 108377 147921 108380
rect 646767 107996 646833 107999
rect 640416 107994 646833 107996
rect 640416 107938 646772 107994
rect 646828 107938 646833 107994
rect 640416 107936 646833 107938
rect 646767 107933 646833 107936
rect 184431 107848 184497 107851
rect 184431 107846 190560 107848
rect 184431 107790 184436 107846
rect 184492 107790 190560 107846
rect 184431 107788 190560 107790
rect 184431 107785 184497 107788
rect 147183 107256 147249 107259
rect 143904 107254 147249 107256
rect 143904 107198 147188 107254
rect 147244 107198 147249 107254
rect 143904 107196 147249 107198
rect 147183 107193 147249 107196
rect 184335 107108 184401 107111
rect 184335 107106 190560 107108
rect 184335 107050 184340 107106
rect 184396 107050 190560 107106
rect 184335 107048 190560 107050
rect 184335 107045 184401 107048
rect 674170 106454 674176 106518
rect 674240 106516 674246 106518
rect 675375 106516 675441 106519
rect 674240 106514 675441 106516
rect 674240 106458 675380 106514
rect 675436 106458 675441 106514
rect 674240 106456 675441 106458
rect 674240 106454 674246 106456
rect 675375 106453 675441 106456
rect 186639 106368 186705 106371
rect 668175 106368 668241 106371
rect 186639 106366 190560 106368
rect 186639 106310 186644 106366
rect 186700 106310 190560 106366
rect 186639 106308 190560 106310
rect 665346 106366 668241 106368
rect 665346 106310 668180 106366
rect 668236 106310 668241 106366
rect 665346 106308 668241 106310
rect 186639 106305 186705 106308
rect 665346 106082 665406 106308
rect 668175 106305 668241 106308
rect 148815 106072 148881 106075
rect 645903 106072 645969 106075
rect 143904 106070 148881 106072
rect 143904 106014 148820 106070
rect 148876 106014 148881 106070
rect 143904 106012 148881 106014
rect 640416 106070 645969 106072
rect 640416 106014 645908 106070
rect 645964 106014 645969 106070
rect 640416 106012 645969 106014
rect 148815 106009 148881 106012
rect 645903 106009 645969 106012
rect 184335 105628 184401 105631
rect 184335 105626 190560 105628
rect 184335 105570 184340 105626
rect 184396 105570 190560 105626
rect 184335 105568 190560 105570
rect 184335 105565 184401 105568
rect 665346 105332 665406 105361
rect 665583 105332 665649 105335
rect 665346 105330 665649 105332
rect 665346 105274 665588 105330
rect 665644 105274 665649 105330
rect 665346 105272 665649 105274
rect 665583 105269 665649 105272
rect 665295 105184 665361 105187
rect 665295 105182 665406 105184
rect 665295 105126 665300 105182
rect 665356 105126 665406 105182
rect 665295 105121 665406 105126
rect 665346 104996 665406 105121
rect 184527 104888 184593 104891
rect 184527 104886 190014 104888
rect 184527 104830 184532 104886
rect 184588 104830 190014 104886
rect 184527 104828 190014 104830
rect 184527 104825 184593 104828
rect 189954 104814 190014 104828
rect 189954 104754 190560 104814
rect 148239 104740 148305 104743
rect 143904 104738 148305 104740
rect 143904 104682 148244 104738
rect 148300 104682 148305 104738
rect 143904 104680 148305 104682
rect 148239 104677 148305 104680
rect 647919 104148 647985 104151
rect 640416 104146 647985 104148
rect 640416 104090 647924 104146
rect 647980 104090 647985 104146
rect 640416 104088 647985 104090
rect 647919 104085 647985 104088
rect 184431 104000 184497 104003
rect 184431 103998 190560 104000
rect 184431 103942 184436 103998
rect 184492 103942 190560 103998
rect 184431 103940 190560 103942
rect 184431 103937 184497 103940
rect 148431 103556 148497 103559
rect 143904 103554 148497 103556
rect 143904 103498 148436 103554
rect 148492 103498 148497 103554
rect 143904 103496 148497 103498
rect 148431 103493 148497 103496
rect 675663 103558 675729 103559
rect 675663 103554 675712 103558
rect 675776 103556 675782 103558
rect 675663 103498 675668 103554
rect 675663 103494 675712 103498
rect 675776 103496 675820 103556
rect 675776 103494 675782 103496
rect 675663 103493 675729 103494
rect 184335 103408 184401 103411
rect 184335 103406 190014 103408
rect 184335 103350 184340 103406
rect 184396 103350 190014 103406
rect 184335 103348 190014 103350
rect 184335 103345 184401 103348
rect 189954 103334 190014 103348
rect 189954 103274 190560 103334
rect 184719 102520 184785 102523
rect 184719 102518 190560 102520
rect 184719 102462 184724 102518
rect 184780 102462 190560 102518
rect 184719 102460 190560 102462
rect 184719 102457 184785 102460
rect 148911 102372 148977 102375
rect 143904 102370 148977 102372
rect 143904 102314 148916 102370
rect 148972 102314 148977 102370
rect 143904 102312 148977 102314
rect 148911 102309 148977 102312
rect 645135 102224 645201 102227
rect 640416 102222 645201 102224
rect 640416 102166 645140 102222
rect 645196 102166 645201 102222
rect 640416 102164 645201 102166
rect 645135 102161 645201 102164
rect 184431 101928 184497 101931
rect 184431 101926 190014 101928
rect 184431 101870 184436 101926
rect 184492 101870 190014 101926
rect 184431 101868 190014 101870
rect 184431 101865 184497 101868
rect 189954 101854 190014 101868
rect 189954 101794 190560 101854
rect 675759 101632 675825 101635
rect 676474 101632 676480 101634
rect 675759 101630 676480 101632
rect 675759 101574 675764 101630
rect 675820 101574 676480 101630
rect 675759 101572 676480 101574
rect 675759 101569 675825 101572
rect 676474 101570 676480 101572
rect 676544 101570 676550 101634
rect 143874 100892 143934 101084
rect 184527 101040 184593 101043
rect 184527 101038 190560 101040
rect 184527 100982 184532 101038
rect 184588 100982 190560 101038
rect 184527 100980 190560 100982
rect 184527 100977 184593 100980
rect 149391 100892 149457 100895
rect 143874 100890 149457 100892
rect 143874 100834 149396 100890
rect 149452 100834 149457 100890
rect 143874 100832 149457 100834
rect 149391 100829 149457 100832
rect 184335 100300 184401 100303
rect 184335 100298 190014 100300
rect 184335 100242 184340 100298
rect 184396 100242 190014 100298
rect 184335 100240 190014 100242
rect 184335 100237 184401 100240
rect 189954 100226 190014 100240
rect 189954 100166 190560 100226
rect 149487 99856 149553 99859
rect 143904 99854 149553 99856
rect 143904 99798 149492 99854
rect 149548 99798 149553 99854
rect 143904 99796 149553 99798
rect 149487 99793 149553 99796
rect 640194 99708 640254 100270
rect 675759 99856 675825 99859
rect 676666 99856 676672 99858
rect 675759 99854 676672 99856
rect 675759 99798 675764 99854
rect 675820 99798 676672 99854
rect 675759 99796 676672 99798
rect 675759 99793 675825 99796
rect 676666 99794 676672 99796
rect 676736 99794 676742 99858
rect 647919 99708 647985 99711
rect 640194 99706 647985 99708
rect 640194 99650 647924 99706
rect 647980 99650 647985 99706
rect 640194 99648 647985 99650
rect 647919 99645 647985 99648
rect 184431 99560 184497 99563
rect 184431 99558 190560 99560
rect 184431 99502 184436 99558
rect 184492 99502 190560 99558
rect 184431 99500 190560 99502
rect 184431 99497 184497 99500
rect 149391 98672 149457 98675
rect 143904 98670 149457 98672
rect 143904 98614 149396 98670
rect 149452 98614 149457 98670
rect 143904 98612 149457 98614
rect 149391 98609 149457 98612
rect 184527 98672 184593 98675
rect 184527 98670 190560 98672
rect 184527 98614 184532 98670
rect 184588 98614 190560 98670
rect 184527 98612 190560 98614
rect 184527 98609 184593 98612
rect 184623 98080 184689 98083
rect 640386 98080 640446 98420
rect 646959 98080 647025 98083
rect 184623 98078 190560 98080
rect 184623 98022 184628 98078
rect 184684 98022 190560 98078
rect 184623 98020 190560 98022
rect 640386 98078 647025 98080
rect 640386 98022 646964 98078
rect 647020 98022 647025 98078
rect 640386 98020 647025 98022
rect 184623 98017 184689 98020
rect 646959 98017 647025 98020
rect 149487 97488 149553 97491
rect 143904 97486 149553 97488
rect 143904 97430 149492 97486
rect 149548 97430 149553 97486
rect 143904 97428 149553 97430
rect 149487 97425 149553 97428
rect 184335 97192 184401 97195
rect 184335 97190 190560 97192
rect 184335 97134 184340 97190
rect 184396 97134 190560 97190
rect 184335 97132 190560 97134
rect 184335 97129 184401 97132
rect 184431 96452 184497 96455
rect 184431 96450 190560 96452
rect 184431 96394 184436 96450
rect 184492 96394 190560 96450
rect 184431 96392 190560 96394
rect 184431 96389 184497 96392
rect 143874 95712 143934 96200
rect 640386 96008 640446 96570
rect 645423 96008 645489 96011
rect 640386 96006 645489 96008
rect 640386 95950 645428 96006
rect 645484 95950 645489 96006
rect 640386 95948 645489 95950
rect 645423 95945 645489 95948
rect 149391 95712 149457 95715
rect 143874 95710 149457 95712
rect 143874 95654 149396 95710
rect 149452 95654 149457 95710
rect 143874 95652 149457 95654
rect 149391 95649 149457 95652
rect 184527 95712 184593 95715
rect 184527 95710 190560 95712
rect 184527 95654 184532 95710
rect 184588 95654 190560 95710
rect 184527 95652 190560 95654
rect 184527 95649 184593 95652
rect 149583 94972 149649 94975
rect 143904 94970 149649 94972
rect 143904 94914 149588 94970
rect 149644 94914 149649 94970
rect 143904 94912 149649 94914
rect 149583 94909 149649 94912
rect 189954 94838 190560 94898
rect 184335 94824 184401 94827
rect 189954 94824 190014 94838
rect 184335 94822 190014 94824
rect 184335 94766 184340 94822
rect 184396 94766 190014 94822
rect 184335 94764 190014 94766
rect 184335 94761 184401 94764
rect 184623 94232 184689 94235
rect 184623 94230 190560 94232
rect 184623 94174 184628 94230
rect 184684 94174 190560 94230
rect 184623 94172 190560 94174
rect 184623 94169 184689 94172
rect 640386 94084 640446 94646
rect 647823 94084 647889 94087
rect 640386 94082 647889 94084
rect 640386 94026 647828 94082
rect 647884 94026 647889 94082
rect 640386 94024 647889 94026
rect 647823 94021 647889 94024
rect 149487 93788 149553 93791
rect 143904 93786 149553 93788
rect 143904 93730 149492 93786
rect 149548 93730 149553 93786
rect 143904 93728 149553 93730
rect 149487 93725 149553 93728
rect 184431 93492 184497 93495
rect 184431 93490 190014 93492
rect 184431 93434 184436 93490
rect 184492 93434 190014 93490
rect 184431 93432 190014 93434
rect 184431 93429 184497 93432
rect 189954 93418 190014 93432
rect 189954 93358 190560 93418
rect 184527 92752 184593 92755
rect 647727 92752 647793 92755
rect 184527 92750 190560 92752
rect 184527 92694 184532 92750
rect 184588 92694 190560 92750
rect 184527 92692 190560 92694
rect 640416 92750 647793 92752
rect 640416 92694 647732 92750
rect 647788 92694 647793 92750
rect 640416 92692 647793 92694
rect 184527 92689 184593 92692
rect 647727 92689 647793 92692
rect 149391 92604 149457 92607
rect 143904 92602 149457 92604
rect 143904 92546 149396 92602
rect 149452 92546 149457 92602
rect 143904 92544 149457 92546
rect 149391 92541 149457 92544
rect 184335 92012 184401 92015
rect 184335 92010 190014 92012
rect 184335 91954 184340 92010
rect 184396 91954 190014 92010
rect 184335 91952 190014 91954
rect 184335 91949 184401 91952
rect 189954 91938 190014 91952
rect 189954 91878 190560 91938
rect 149295 91420 149361 91423
rect 143904 91418 149361 91420
rect 143904 91362 149300 91418
rect 149356 91362 149361 91418
rect 143904 91360 149361 91362
rect 149295 91357 149361 91360
rect 184623 91124 184689 91127
rect 184623 91122 190560 91124
rect 184623 91066 184628 91122
rect 184684 91066 190560 91122
rect 184623 91064 190560 91066
rect 184623 91061 184689 91064
rect 659343 90828 659409 90831
rect 640416 90826 659409 90828
rect 640416 90770 659348 90826
rect 659404 90770 659409 90826
rect 640416 90768 659409 90770
rect 659343 90765 659409 90768
rect 184431 90384 184497 90387
rect 184431 90382 190560 90384
rect 184431 90326 184436 90382
rect 184492 90326 190560 90382
rect 184431 90324 190560 90326
rect 184431 90321 184497 90324
rect 149199 90236 149265 90239
rect 143904 90234 149265 90236
rect 143904 90178 149204 90234
rect 149260 90178 149265 90234
rect 143904 90176 149265 90178
rect 149199 90173 149265 90176
rect 184527 89644 184593 89647
rect 184527 89642 190560 89644
rect 184527 89586 184532 89642
rect 184588 89586 190560 89642
rect 184527 89584 190560 89586
rect 184527 89581 184593 89584
rect 149391 89052 149457 89055
rect 143904 89050 149457 89052
rect 143904 88994 149396 89050
rect 149452 88994 149457 89050
rect 143904 88992 149457 88994
rect 149391 88989 149457 88992
rect 184335 88904 184401 88907
rect 645903 88904 645969 88907
rect 184335 88902 190560 88904
rect 184335 88846 184340 88902
rect 184396 88846 190560 88902
rect 184335 88844 190560 88846
rect 640416 88902 645969 88904
rect 640416 88846 645908 88902
rect 645964 88846 645969 88902
rect 640416 88844 645969 88846
rect 184335 88841 184401 88844
rect 645903 88841 645969 88844
rect 184431 88164 184497 88167
rect 184431 88162 190014 88164
rect 184431 88106 184436 88162
rect 184492 88106 190014 88162
rect 184431 88104 190014 88106
rect 184431 88101 184497 88104
rect 189954 88090 190014 88104
rect 189954 88030 190560 88090
rect 143874 87276 143934 87764
rect 149487 87276 149553 87279
rect 143874 87274 149553 87276
rect 143874 87218 149492 87274
rect 149548 87218 149553 87274
rect 143874 87216 149553 87218
rect 149487 87213 149553 87216
rect 184527 87276 184593 87279
rect 184527 87274 190560 87276
rect 184527 87218 184532 87274
rect 184588 87218 190560 87274
rect 184527 87216 190560 87218
rect 184527 87213 184593 87216
rect 647919 87128 647985 87131
rect 640386 87126 647985 87128
rect 640386 87070 647924 87126
rect 647980 87070 647985 87126
rect 640386 87068 647985 87070
rect 640386 86950 640446 87068
rect 647919 87065 647985 87068
rect 653679 86980 653745 86983
rect 653679 86978 656736 86980
rect 653679 86922 653684 86978
rect 653740 86922 656736 86978
rect 653679 86920 656736 86922
rect 653679 86917 653745 86920
rect 184623 86684 184689 86687
rect 184623 86682 190014 86684
rect 184623 86626 184628 86682
rect 184684 86626 190014 86682
rect 184623 86624 190014 86626
rect 184623 86621 184689 86624
rect 189954 86610 190014 86624
rect 189954 86550 190560 86610
rect 148719 86536 148785 86539
rect 143904 86534 148785 86536
rect 143904 86478 148724 86534
rect 148780 86478 148785 86534
rect 143904 86476 148785 86478
rect 148719 86473 148785 86476
rect 663279 86388 663345 86391
rect 663234 86386 663345 86388
rect 663234 86330 663284 86386
rect 663340 86330 663345 86386
rect 663234 86325 663345 86330
rect 650895 86240 650961 86243
rect 650895 86238 656736 86240
rect 650895 86182 650900 86238
rect 650956 86182 656736 86238
rect 663234 86210 663294 86325
rect 650895 86180 656736 86182
rect 650895 86177 650961 86180
rect 184335 85796 184401 85799
rect 184335 85794 190560 85796
rect 184335 85738 184340 85794
rect 184396 85738 190560 85794
rect 184335 85736 190560 85738
rect 184335 85733 184401 85736
rect 148623 85352 148689 85355
rect 143904 85350 148689 85352
rect 143904 85294 148628 85350
rect 148684 85294 148689 85350
rect 143904 85292 148689 85294
rect 148623 85289 148689 85292
rect 652335 85352 652401 85355
rect 652335 85350 656736 85352
rect 652335 85294 652340 85350
rect 652396 85294 656736 85350
rect 652335 85292 656736 85294
rect 652335 85289 652401 85292
rect 184527 85204 184593 85207
rect 184527 85202 190014 85204
rect 184527 85146 184532 85202
rect 184588 85146 190014 85202
rect 184527 85144 190014 85146
rect 184527 85141 184593 85144
rect 189954 85130 190014 85144
rect 189954 85070 190560 85130
rect 640194 84464 640254 85026
rect 663234 84763 663294 85322
rect 663234 84758 663345 84763
rect 663234 84702 663284 84758
rect 663340 84702 663345 84758
rect 663234 84700 663345 84702
rect 663279 84697 663345 84700
rect 645903 84464 645969 84467
rect 640194 84462 645969 84464
rect 640194 84406 645908 84462
rect 645964 84406 645969 84462
rect 640194 84404 645969 84406
rect 645903 84401 645969 84404
rect 184431 84316 184497 84319
rect 651759 84316 651825 84319
rect 184431 84314 190560 84316
rect 184431 84258 184436 84314
rect 184492 84258 190560 84314
rect 184431 84256 190560 84258
rect 651759 84314 656736 84316
rect 651759 84258 651764 84314
rect 651820 84258 656736 84314
rect 651759 84256 656736 84258
rect 184431 84253 184497 84256
rect 651759 84253 651825 84256
rect 146991 84168 147057 84171
rect 143904 84166 147057 84168
rect 143904 84110 146996 84166
rect 147052 84110 147057 84166
rect 143904 84108 147057 84110
rect 146991 84105 147057 84108
rect 663426 84023 663486 84582
rect 663375 84018 663486 84023
rect 663375 83962 663380 84018
rect 663436 83962 663486 84018
rect 663375 83960 663486 83962
rect 663375 83957 663441 83960
rect 189954 83442 190560 83502
rect 184335 83428 184401 83431
rect 189954 83428 190014 83442
rect 184335 83426 190014 83428
rect 184335 83370 184340 83426
rect 184396 83370 190014 83426
rect 184335 83368 190014 83370
rect 652239 83428 652305 83431
rect 652239 83426 656736 83428
rect 652239 83370 652244 83426
rect 652300 83370 656736 83426
rect 652239 83368 656736 83370
rect 184335 83365 184401 83368
rect 652239 83365 652305 83368
rect 143874 82392 143934 82880
rect 186159 82836 186225 82839
rect 186159 82834 190560 82836
rect 186159 82778 186164 82834
rect 186220 82778 190560 82834
rect 186159 82776 190560 82778
rect 186159 82773 186225 82776
rect 640386 82688 640446 83176
rect 663426 82839 663486 83398
rect 663426 82834 663537 82839
rect 663426 82778 663476 82834
rect 663532 82778 663537 82834
rect 663426 82776 663537 82778
rect 663471 82773 663537 82776
rect 647919 82688 647985 82691
rect 640386 82686 647985 82688
rect 640386 82630 647924 82686
rect 647980 82630 647985 82686
rect 640386 82628 647985 82630
rect 647919 82625 647985 82628
rect 652431 82688 652497 82691
rect 652431 82686 656736 82688
rect 652431 82630 652436 82686
rect 652492 82630 656736 82686
rect 652431 82628 656736 82630
rect 652431 82625 652497 82628
rect 148911 82392 148977 82395
rect 143874 82390 148977 82392
rect 143874 82334 148916 82390
rect 148972 82334 148977 82390
rect 143874 82332 148977 82334
rect 148911 82329 148977 82332
rect 663234 82099 663294 82658
rect 663234 82094 663345 82099
rect 663234 82038 663284 82094
rect 663340 82038 663345 82094
rect 663234 82036 663345 82038
rect 663279 82033 663345 82036
rect 184239 81948 184305 81951
rect 184239 81946 190560 81948
rect 184239 81890 184244 81946
rect 184300 81890 190560 81946
rect 184239 81888 190560 81890
rect 184239 81885 184305 81888
rect 148239 81652 148305 81655
rect 143904 81650 148305 81652
rect 143904 81594 148244 81650
rect 148300 81594 148305 81650
rect 143904 81592 148305 81594
rect 148239 81589 148305 81592
rect 662415 81652 662481 81655
rect 663042 81652 663102 81770
rect 662415 81650 663102 81652
rect 662415 81594 662420 81650
rect 662476 81594 663102 81650
rect 662415 81592 663102 81594
rect 662415 81589 662481 81592
rect 184431 81356 184497 81359
rect 184431 81354 190560 81356
rect 184431 81298 184436 81354
rect 184492 81298 190560 81354
rect 184431 81296 190560 81298
rect 184431 81293 184497 81296
rect 640386 81060 640446 81326
rect 647919 81060 647985 81063
rect 640386 81058 647985 81060
rect 640386 81002 647924 81058
rect 647980 81002 647985 81058
rect 640386 81000 647985 81002
rect 647919 80997 647985 81000
rect 149583 80468 149649 80471
rect 143904 80466 149649 80468
rect 143904 80410 149588 80466
rect 149644 80410 149649 80466
rect 143904 80408 149649 80410
rect 149583 80405 149649 80408
rect 184623 80468 184689 80471
rect 184623 80466 190560 80468
rect 184623 80410 184628 80466
rect 184684 80410 190560 80466
rect 184623 80408 190560 80410
rect 184623 80405 184689 80408
rect 184431 79876 184497 79879
rect 184431 79874 190014 79876
rect 184431 79818 184436 79874
rect 184492 79818 190014 79874
rect 184431 79816 190014 79818
rect 184431 79813 184497 79816
rect 189954 79802 190014 79816
rect 189954 79742 190560 79802
rect 645519 79432 645585 79435
rect 640416 79430 645585 79432
rect 640416 79374 645524 79430
rect 645580 79374 645585 79430
rect 640416 79372 645585 79374
rect 645519 79369 645585 79372
rect 149679 79284 149745 79287
rect 143904 79282 149745 79284
rect 143904 79226 149684 79282
rect 149740 79226 149745 79282
rect 143904 79224 149745 79226
rect 149679 79221 149745 79224
rect 184335 78988 184401 78991
rect 184335 78986 190560 78988
rect 184335 78930 184340 78986
rect 184396 78930 190560 78986
rect 184335 78928 190560 78930
rect 184335 78925 184401 78928
rect 184527 78248 184593 78251
rect 184527 78246 190014 78248
rect 184527 78190 184532 78246
rect 184588 78190 190014 78246
rect 184527 78188 190014 78190
rect 184527 78185 184593 78188
rect 189954 78174 190014 78188
rect 189954 78114 190560 78174
rect 148815 77952 148881 77955
rect 143904 77950 148881 77952
rect 143904 77894 148820 77950
rect 148876 77894 148881 77950
rect 143904 77892 148881 77894
rect 148815 77889 148881 77892
rect 184431 77508 184497 77511
rect 647919 77508 647985 77511
rect 184431 77506 190560 77508
rect 184431 77450 184436 77506
rect 184492 77450 190560 77506
rect 184431 77448 190560 77450
rect 640416 77506 647985 77508
rect 640416 77450 647924 77506
rect 647980 77450 647985 77506
rect 640416 77448 647985 77450
rect 184431 77445 184497 77448
rect 647919 77445 647985 77448
rect 149391 76768 149457 76771
rect 143904 76766 149457 76768
rect 143904 76710 149396 76766
rect 149452 76710 149457 76766
rect 143904 76708 149457 76710
rect 149391 76705 149457 76708
rect 184335 76768 184401 76771
rect 184335 76766 190014 76768
rect 184335 76710 184340 76766
rect 184396 76710 190014 76766
rect 184335 76708 190014 76710
rect 184335 76705 184401 76708
rect 189954 76694 190014 76708
rect 189954 76634 190560 76694
rect 184623 76028 184689 76031
rect 184623 76026 190560 76028
rect 184623 75970 184628 76026
rect 184684 75970 190560 76026
rect 184623 75968 190560 75970
rect 184623 75965 184689 75968
rect 149199 75584 149265 75587
rect 645999 75584 646065 75587
rect 143904 75582 149265 75584
rect 143904 75526 149204 75582
rect 149260 75526 149265 75582
rect 143904 75524 149265 75526
rect 640416 75582 646065 75584
rect 640416 75526 646004 75582
rect 646060 75526 646065 75582
rect 640416 75524 646065 75526
rect 149199 75521 149265 75524
rect 645999 75521 646065 75524
rect 184527 75140 184593 75143
rect 184527 75138 190560 75140
rect 184527 75082 184532 75138
rect 184588 75082 190560 75138
rect 184527 75080 190560 75082
rect 184527 75077 184593 75080
rect 184335 74400 184401 74403
rect 184335 74398 190560 74400
rect 184335 74342 184340 74398
rect 184396 74342 190560 74398
rect 184335 74340 190560 74342
rect 184335 74337 184401 74340
rect 143874 73808 143934 74296
rect 149295 73808 149361 73811
rect 143874 73806 149361 73808
rect 143874 73750 149300 73806
rect 149356 73750 149361 73806
rect 143874 73748 149361 73750
rect 149295 73745 149361 73748
rect 184527 73660 184593 73663
rect 647919 73660 647985 73663
rect 184527 73658 190560 73660
rect 184527 73602 184532 73658
rect 184588 73602 190560 73658
rect 184527 73600 190560 73602
rect 640416 73658 647985 73660
rect 640416 73602 647924 73658
rect 647980 73602 647985 73658
rect 640416 73600 647985 73602
rect 184527 73597 184593 73600
rect 647919 73597 647985 73600
rect 149007 73068 149073 73071
rect 143904 73066 149073 73068
rect 143904 73010 149012 73066
rect 149068 73010 149073 73066
rect 143904 73008 149073 73010
rect 149007 73005 149073 73008
rect 184431 72920 184497 72923
rect 184431 72918 190560 72920
rect 184431 72862 184436 72918
rect 184492 72862 190560 72918
rect 184431 72860 190560 72862
rect 184431 72857 184497 72860
rect 184623 72180 184689 72183
rect 184623 72178 190560 72180
rect 184623 72122 184628 72178
rect 184684 72122 190560 72178
rect 184623 72120 190560 72122
rect 184623 72117 184689 72120
rect 149103 72032 149169 72035
rect 143904 72030 149169 72032
rect 143904 71974 149108 72030
rect 149164 71974 149169 72030
rect 143904 71972 149169 71974
rect 149103 71969 149169 71972
rect 647055 71884 647121 71887
rect 640386 71882 647121 71884
rect 640386 71826 647060 71882
rect 647116 71826 647121 71882
rect 640386 71824 647121 71826
rect 640386 71706 640446 71824
rect 647055 71821 647121 71824
rect 184335 71440 184401 71443
rect 184335 71438 190014 71440
rect 184335 71382 184340 71438
rect 184396 71382 190014 71438
rect 184335 71380 190014 71382
rect 184335 71377 184401 71380
rect 189954 71366 190014 71380
rect 189954 71306 190560 71366
rect 149487 70848 149553 70851
rect 143904 70846 149553 70848
rect 143904 70790 149492 70846
rect 149548 70790 149553 70846
rect 143904 70788 149553 70790
rect 149487 70785 149553 70788
rect 184431 70552 184497 70555
rect 184431 70550 190560 70552
rect 184431 70494 184436 70550
rect 184492 70494 190560 70550
rect 184431 70492 190560 70494
rect 184431 70489 184497 70492
rect 184527 69960 184593 69963
rect 184527 69958 190014 69960
rect 184527 69902 184532 69958
rect 184588 69902 190014 69958
rect 184527 69900 190014 69902
rect 184527 69897 184593 69900
rect 189954 69886 190014 69900
rect 189954 69826 190560 69886
rect 640386 69664 640446 69856
rect 647919 69664 647985 69667
rect 640386 69662 647985 69664
rect 640386 69606 647924 69662
rect 647980 69606 647985 69662
rect 640386 69604 647985 69606
rect 647919 69601 647985 69604
rect 149391 69516 149457 69519
rect 143904 69514 149457 69516
rect 143904 69458 149396 69514
rect 149452 69458 149457 69514
rect 143904 69456 149457 69458
rect 149391 69453 149457 69456
rect 184335 69072 184401 69075
rect 184335 69070 190560 69072
rect 184335 69014 184340 69070
rect 184396 69014 190560 69070
rect 184335 69012 190560 69014
rect 184335 69009 184401 69012
rect 646863 68628 646929 68631
rect 640194 68626 646929 68628
rect 640194 68570 646868 68626
rect 646924 68570 646929 68626
rect 640194 68568 646929 68570
rect 184431 68480 184497 68483
rect 184431 68478 190014 68480
rect 184431 68422 184436 68478
rect 184492 68422 190014 68478
rect 184431 68420 190014 68422
rect 184431 68417 184497 68420
rect 189954 68406 190014 68420
rect 189954 68346 190560 68406
rect 149199 68332 149265 68335
rect 143904 68330 149265 68332
rect 143904 68274 149204 68330
rect 149260 68274 149265 68330
rect 143904 68272 149265 68274
rect 149199 68269 149265 68272
rect 640194 68006 640254 68568
rect 646863 68565 646929 68568
rect 184335 67592 184401 67595
rect 184335 67590 190560 67592
rect 184335 67534 184340 67590
rect 184396 67534 190560 67590
rect 184335 67532 190560 67534
rect 184335 67529 184401 67532
rect 149583 67148 149649 67151
rect 143904 67146 149649 67148
rect 143904 67090 149588 67146
rect 149644 67090 149649 67146
rect 143904 67088 149649 67090
rect 149583 67085 149649 67088
rect 184527 66852 184593 66855
rect 184527 66850 190560 66852
rect 184527 66794 184532 66850
rect 184588 66794 190560 66850
rect 184527 66792 190560 66794
rect 184527 66789 184593 66792
rect 645999 66260 646065 66263
rect 640194 66258 646065 66260
rect 640194 66202 646004 66258
rect 646060 66202 646065 66258
rect 640194 66200 646065 66202
rect 184335 66112 184401 66115
rect 184335 66110 190560 66112
rect 184335 66054 184340 66110
rect 184396 66054 190560 66110
rect 640194 66082 640254 66200
rect 645999 66197 646065 66200
rect 184335 66052 190560 66054
rect 184335 66049 184401 66052
rect 143874 65372 143934 65860
rect 149487 65372 149553 65375
rect 143874 65370 149553 65372
rect 143874 65314 149492 65370
rect 149548 65314 149553 65370
rect 143874 65312 149553 65314
rect 149487 65309 149553 65312
rect 184527 65224 184593 65227
rect 184527 65222 190560 65224
rect 184527 65166 184532 65222
rect 184588 65166 190560 65222
rect 184527 65164 190560 65166
rect 184527 65161 184593 65164
rect 149391 64632 149457 64635
rect 143904 64630 149457 64632
rect 143904 64574 149396 64630
rect 149452 64574 149457 64630
rect 143904 64572 149457 64574
rect 149391 64569 149457 64572
rect 184623 64632 184689 64635
rect 184623 64630 190014 64632
rect 184623 64574 184628 64630
rect 184684 64574 190014 64630
rect 184623 64572 190014 64574
rect 184623 64569 184689 64572
rect 189954 64558 190014 64572
rect 189954 64498 190560 64558
rect 647919 64188 647985 64191
rect 640416 64186 647985 64188
rect 640416 64130 647924 64186
rect 647980 64130 647985 64186
rect 640416 64128 647985 64130
rect 647919 64125 647985 64128
rect 184431 63744 184497 63747
rect 184431 63742 190560 63744
rect 184431 63686 184436 63742
rect 184492 63686 190560 63742
rect 184431 63684 190560 63686
rect 184431 63681 184497 63684
rect 149295 63448 149361 63451
rect 143904 63446 149361 63448
rect 143904 63390 149300 63446
rect 149356 63390 149361 63446
rect 143904 63388 149361 63390
rect 149295 63385 149361 63388
rect 184335 63152 184401 63155
rect 184335 63150 190014 63152
rect 184335 63094 184340 63150
rect 184396 63094 190014 63150
rect 184335 63092 190014 63094
rect 184335 63089 184401 63092
rect 189954 63078 190014 63092
rect 189954 63018 190560 63078
rect 149487 62264 149553 62267
rect 143904 62262 149553 62264
rect 143904 62206 149492 62262
rect 149548 62206 149553 62262
rect 143904 62204 149553 62206
rect 149487 62201 149553 62204
rect 184431 62264 184497 62267
rect 647919 62264 647985 62267
rect 184431 62262 190560 62264
rect 184431 62206 184436 62262
rect 184492 62206 190560 62262
rect 184431 62204 190560 62206
rect 640416 62262 647985 62264
rect 640416 62206 647924 62262
rect 647980 62206 647985 62262
rect 640416 62204 647985 62206
rect 184431 62201 184497 62204
rect 647919 62201 647985 62204
rect 184527 61524 184593 61527
rect 184527 61522 190014 61524
rect 184527 61466 184532 61522
rect 184588 61466 190014 61522
rect 184527 61464 190014 61466
rect 184527 61461 184593 61464
rect 189954 61450 190014 61464
rect 189954 61390 190560 61450
rect 143874 60636 143934 60976
rect 184623 60784 184689 60787
rect 184623 60782 190560 60784
rect 184623 60726 184628 60782
rect 184684 60726 190560 60782
rect 184623 60724 190560 60726
rect 184623 60721 184689 60724
rect 149391 60636 149457 60639
rect 143874 60634 149457 60636
rect 143874 60578 149396 60634
rect 149452 60578 149457 60634
rect 143874 60576 149457 60578
rect 149391 60573 149457 60576
rect 647151 60340 647217 60343
rect 640416 60338 647217 60340
rect 640416 60282 647156 60338
rect 647212 60282 647217 60338
rect 640416 60280 647217 60282
rect 647151 60277 647217 60280
rect 184335 60044 184401 60047
rect 184335 60042 190014 60044
rect 184335 59986 184340 60042
rect 184396 59986 190014 60042
rect 184335 59984 190014 59986
rect 184335 59981 184401 59984
rect 189954 59970 190014 59984
rect 189954 59910 190560 59970
rect 149391 59748 149457 59751
rect 143904 59746 149457 59748
rect 143904 59690 149396 59746
rect 149452 59690 149457 59746
rect 143904 59688 149457 59690
rect 149391 59685 149457 59688
rect 184431 59304 184497 59307
rect 184431 59302 190560 59304
rect 184431 59246 184436 59302
rect 184492 59246 190560 59302
rect 184431 59244 190560 59246
rect 184431 59241 184497 59244
rect 645999 59008 646065 59011
rect 640386 59006 646065 59008
rect 640386 58950 646004 59006
rect 646060 58950 646065 59006
rect 640386 58948 646065 58950
rect 149391 58564 149457 58567
rect 143904 58562 149457 58564
rect 143904 58506 149396 58562
rect 149452 58506 149457 58562
rect 143904 58504 149457 58506
rect 149391 58501 149457 58504
rect 184527 58416 184593 58419
rect 184527 58414 190560 58416
rect 184527 58358 184532 58414
rect 184588 58358 190560 58414
rect 640386 58386 640446 58948
rect 645999 58945 646065 58948
rect 184527 58356 190560 58358
rect 184527 58353 184593 58356
rect 184335 57676 184401 57679
rect 184335 57674 190560 57676
rect 184335 57618 184340 57674
rect 184396 57618 190560 57674
rect 184335 57616 190560 57618
rect 184335 57613 184401 57616
rect 149487 57380 149553 57383
rect 143904 57378 149553 57380
rect 143904 57322 149492 57378
rect 149548 57322 149553 57378
rect 143904 57320 149553 57322
rect 149487 57317 149553 57320
rect 646767 57084 646833 57087
rect 640386 57082 646833 57084
rect 640386 57026 646772 57082
rect 646828 57026 646833 57082
rect 640386 57024 646833 57026
rect 184335 56936 184401 56939
rect 184335 56934 190560 56936
rect 184335 56878 184340 56934
rect 184396 56878 190560 56934
rect 184335 56876 190560 56878
rect 184335 56873 184401 56876
rect 640386 56536 640446 57024
rect 646767 57021 646833 57024
rect 149391 56196 149457 56199
rect 143874 56194 149457 56196
rect 143874 56138 149396 56194
rect 149452 56138 149457 56194
rect 143874 56136 149457 56138
rect 143874 56092 143934 56136
rect 149391 56133 149457 56136
rect 184335 56196 184401 56199
rect 184335 56194 190560 56196
rect 184335 56138 184340 56194
rect 184396 56138 190560 56194
rect 184335 56136 190560 56138
rect 184335 56133 184401 56136
rect 184431 55456 184497 55459
rect 184431 55454 190560 55456
rect 184431 55398 184436 55454
rect 184492 55398 190560 55454
rect 184431 55396 190560 55398
rect 184431 55393 184497 55396
rect 149679 54864 149745 54867
rect 143904 54862 149745 54864
rect 143904 54806 149684 54862
rect 149740 54806 149745 54862
rect 143904 54804 149745 54806
rect 149679 54801 149745 54804
rect 184335 54716 184401 54719
rect 646479 54716 646545 54719
rect 184335 54714 190014 54716
rect 184335 54658 184340 54714
rect 184396 54658 190014 54714
rect 184335 54656 190014 54658
rect 184335 54653 184401 54656
rect 189954 54642 190014 54656
rect 640386 54714 646545 54716
rect 640386 54658 646484 54714
rect 646540 54658 646545 54714
rect 640386 54656 646545 54658
rect 189954 54582 190560 54642
rect 640386 54612 640446 54656
rect 646479 54653 646545 54656
rect 184335 53976 184401 53979
rect 184335 53974 190560 53976
rect 184335 53918 184340 53974
rect 184396 53918 190560 53974
rect 184335 53916 190560 53918
rect 184335 53913 184401 53916
rect 149391 53828 149457 53831
rect 143904 53826 149457 53828
rect 143904 53770 149396 53826
rect 149452 53770 149457 53826
rect 143904 53768 149457 53770
rect 149391 53765 149457 53768
rect 426159 44948 426225 44951
rect 472239 44948 472305 44951
rect 419394 44946 426225 44948
rect 419394 44890 426164 44946
rect 426220 44890 426225 44946
rect 419394 44888 426225 44890
rect 419394 44404 419454 44888
rect 426159 44885 426225 44888
rect 472194 44946 472305 44948
rect 472194 44890 472244 44946
rect 472300 44890 472305 44946
rect 472194 44885 472305 44890
rect 472194 44404 472254 44885
rect 415215 41988 415281 41991
rect 415215 41986 417630 41988
rect 415215 41930 415220 41986
rect 415276 41930 417630 41986
rect 415215 41928 417630 41930
rect 415215 41925 415281 41928
rect 416847 41840 416913 41843
rect 416847 41838 416958 41840
rect 416847 41782 416852 41838
rect 416908 41782 416958 41838
rect 416847 41777 416958 41782
rect 416898 40508 416958 41777
rect 417570 40656 417630 41928
rect 464847 41840 464913 41843
rect 457890 41838 464913 41840
rect 457890 41782 464852 41838
rect 464908 41782 464913 41838
rect 457890 41780 464913 41782
rect 457890 40656 457950 41780
rect 464847 41777 464913 41780
rect 470319 41840 470385 41843
rect 512175 41840 512241 41843
rect 525903 41840 525969 41843
rect 470319 41838 478110 41840
rect 470319 41782 470324 41838
rect 470380 41782 478110 41838
rect 470319 41780 478110 41782
rect 470319 41777 470385 41780
rect 417570 40596 457950 40656
rect 417466 40508 417472 40510
rect 416898 40448 417472 40508
rect 417466 40446 417472 40448
rect 417536 40446 417542 40510
rect 417658 40446 417664 40510
rect 417728 40508 417734 40510
rect 420783 40508 420849 40511
rect 417728 40506 420849 40508
rect 417728 40450 420788 40506
rect 420844 40450 420849 40506
rect 417728 40448 420849 40450
rect 478050 40508 478110 41780
rect 512175 41838 525969 41840
rect 512175 41782 512180 41838
rect 512236 41782 525908 41838
rect 525964 41782 525969 41838
rect 512175 41780 525969 41782
rect 512175 41777 512241 41780
rect 525903 41777 525969 41780
rect 539727 40508 539793 40511
rect 478050 40506 539793 40508
rect 478050 40450 539732 40506
rect 539788 40450 539793 40506
rect 478050 40448 539793 40450
rect 417728 40446 417734 40448
rect 420783 40445 420849 40448
rect 539727 40445 539793 40448
rect 142095 40212 142161 40215
rect 141762 40210 142161 40212
rect 141762 40154 142100 40210
rect 142156 40154 142161 40210
rect 141762 40152 142161 40154
rect 141762 39886 141822 40152
rect 142095 40149 142161 40152
rect 311055 37252 311121 37255
rect 328335 37252 328401 37255
rect 311055 37250 328401 37252
rect 311055 37194 311060 37250
rect 311116 37194 328340 37250
rect 328396 37194 328401 37250
rect 311055 37192 328401 37194
rect 311055 37189 311121 37192
rect 328335 37189 328401 37192
<< via3 >>
rect 673984 873390 674048 873454
rect 673984 852522 674048 852586
rect 40384 815078 40448 815142
rect 40576 814042 40640 814106
rect 40768 813006 40832 813070
rect 41536 805014 41600 805078
rect 41920 801078 41984 801082
rect 41920 801022 41932 801078
rect 41932 801022 41984 801078
rect 41920 801018 41984 801022
rect 42496 800722 42560 800786
rect 42304 800574 42368 800638
rect 42496 800426 42560 800490
rect 41920 798798 41984 798862
rect 40768 793914 40832 793978
rect 42304 790214 42368 790278
rect 41536 786366 41600 786430
rect 674752 774526 674816 774590
rect 674560 773638 674624 773702
rect 676096 773046 676160 773110
rect 40576 772306 40640 772370
rect 40192 771862 40256 771926
rect 40384 771862 40448 771926
rect 40576 770826 40640 770890
rect 675904 770678 675968 770742
rect 675520 769998 675584 770002
rect 675520 769942 675532 769998
rect 675532 769942 675584 769998
rect 675520 769938 675584 769942
rect 40768 769790 40832 769854
rect 674368 769346 674432 769410
rect 41344 768902 41408 768966
rect 41152 760170 41216 760234
rect 42112 757950 42176 758014
rect 42304 757802 42368 757866
rect 42304 752474 42368 752538
rect 42112 751142 42176 751206
rect 40768 748774 40832 748838
rect 41344 747294 41408 747358
rect 41152 746998 41216 747062
rect 677056 731606 677120 731670
rect 674944 729830 675008 729894
rect 40576 729238 40640 729302
rect 676288 729386 676352 729450
rect 40384 728706 40448 728710
rect 40384 728650 40436 728706
rect 40436 728650 40448 728706
rect 40384 728646 40448 728650
rect 675712 728706 675776 728710
rect 675712 728650 675724 728706
rect 675724 728650 675776 728706
rect 675712 728646 675776 728650
rect 40576 727610 40640 727674
rect 675328 726782 675392 726786
rect 675328 726726 675380 726782
rect 675380 726726 675392 726782
rect 675328 726722 675392 726726
rect 676480 726130 676544 726194
rect 673984 725834 674048 725898
rect 41152 725686 41216 725750
rect 40960 723762 41024 723826
rect 676864 721838 676928 721902
rect 42304 718582 42368 718646
rect 40384 717694 40448 717758
rect 40768 716954 40832 717018
rect 40576 716806 40640 716870
rect 40576 708814 40640 708878
rect 42304 708666 42368 708730
rect 40768 708518 40832 708582
rect 40960 705854 41024 705918
rect 41152 705410 41216 705474
rect 40384 701266 40448 701330
rect 676096 698898 676160 698962
rect 674752 697714 674816 697778
rect 674560 695790 674624 695854
rect 675904 695198 675968 695262
rect 675520 695050 675584 695114
rect 674368 693126 674432 693190
rect 677056 692534 677120 692598
rect 674176 685578 674240 685642
rect 40384 685430 40448 685494
rect 675904 684394 675968 684458
rect 40768 683358 40832 683422
rect 675520 682678 675584 682682
rect 675520 682622 675572 682678
rect 675572 682622 675584 682678
rect 675520 682618 675584 682622
rect 40576 682470 40640 682534
rect 41152 681878 41216 681942
rect 41920 681730 41984 681794
rect 40960 680398 41024 680462
rect 42304 680250 42368 680314
rect 42112 679658 42176 679722
rect 41728 678770 41792 678834
rect 676096 678326 676160 678390
rect 42304 678178 42368 678242
rect 41536 677438 41600 677502
rect 677056 676846 677120 676910
rect 674368 673294 674432 673358
rect 674560 671370 674624 671434
rect 41536 668558 41600 668622
rect 41920 668410 41984 668474
rect 41728 668262 41792 668326
rect 42304 666190 42368 666254
rect 42496 665450 42560 665514
rect 42112 665302 42176 665366
rect 40768 664266 40832 664330
rect 40960 663970 41024 664034
rect 41152 662490 41216 662554
rect 40576 661454 40640 661518
rect 675712 654498 675776 654562
rect 674944 653462 675008 653526
rect 675328 653018 675392 653082
rect 676288 651390 676352 651454
rect 676480 651390 676544 651454
rect 673984 650502 674048 650566
rect 677056 649762 677120 649826
rect 676864 648726 676928 648790
rect 40384 642214 40448 642278
rect 40576 642214 40640 642278
rect 676672 641622 676736 641686
rect 40768 640290 40832 640354
rect 675136 640290 675200 640354
rect 673984 640142 674048 640206
rect 40576 639254 40640 639318
rect 41344 638662 41408 638726
rect 42688 638514 42752 638578
rect 674752 638366 674816 638430
rect 42304 637182 42368 637246
rect 43072 637034 43136 637098
rect 42112 636442 42176 636506
rect 41728 635554 41792 635618
rect 41920 634962 41984 635026
rect 41536 634222 41600 634286
rect 675328 634134 675392 634138
rect 675328 634078 675380 634134
rect 675380 634078 675392 634134
rect 675328 634074 675392 634078
rect 676864 632742 676928 632806
rect 676288 629042 676352 629106
rect 676480 627266 676544 627330
rect 41536 625934 41600 625998
rect 41728 625046 41792 625110
rect 42112 623862 42176 623926
rect 41920 622086 41984 622150
rect 42304 621938 42368 622002
rect 40768 621346 40832 621410
rect 42688 620754 42752 620818
rect 40576 617646 40640 617710
rect 43072 617202 43136 617266
rect 41344 616610 41408 616674
rect 675904 610098 675968 610162
rect 674368 609654 674432 609718
rect 674176 609062 674240 609126
rect 675520 608618 675584 608682
rect 676096 608470 676160 608534
rect 674560 607582 674624 607646
rect 40384 601722 40448 601726
rect 40384 601666 40396 601722
rect 40396 601666 40448 601722
rect 40384 601662 40448 601666
rect 40576 597074 40640 597138
rect 674176 597074 674240 597138
rect 40384 596038 40448 596102
rect 674560 596038 674624 596102
rect 40768 595594 40832 595658
rect 42880 595298 42944 595362
rect 40960 594114 41024 594178
rect 674944 593966 675008 594030
rect 42112 593818 42176 593882
rect 42304 593374 42368 593438
rect 41536 592042 41600 592106
rect 41728 591746 41792 591810
rect 41920 591376 41984 591440
rect 675520 589734 675584 589738
rect 675520 589678 675532 589734
rect 675532 589678 675584 589734
rect 675520 589674 675584 589678
rect 675904 584642 675968 584706
rect 41536 583014 41600 583078
rect 675712 582926 675776 582930
rect 675712 582870 675724 582926
rect 675724 582870 675776 582926
rect 675712 582866 675776 582870
rect 41920 582570 41984 582634
rect 42112 581682 42176 581746
rect 42304 580498 42368 580562
rect 42880 579522 42944 579526
rect 42880 579466 42932 579522
rect 42932 579466 42944 579522
rect 42880 579462 42944 579466
rect 41728 578870 41792 578934
rect 40576 576354 40640 576418
rect 40960 576206 41024 576270
rect 40768 576058 40832 576122
rect 40384 573838 40448 573902
rect 676096 567178 676160 567242
rect 675136 564958 675200 565022
rect 676288 564662 676352 564726
rect 676672 564218 676736 564282
rect 674752 563478 674816 563542
rect 675328 562886 675392 562950
rect 676480 562738 676544 562802
rect 673984 561998 674048 562062
rect 676864 560222 676928 560286
rect 674368 552970 674432 553034
rect 673984 552230 674048 552294
rect 675136 551698 675200 551702
rect 675136 551642 675188 551698
rect 675188 551642 675200 551698
rect 675136 551638 675200 551642
rect 674752 550158 674816 550222
rect 675328 545482 675392 545486
rect 675328 545426 675380 545482
rect 675380 545426 675392 545482
rect 675328 545422 675392 545426
rect 676864 544238 676928 544302
rect 676288 540538 676352 540602
rect 40384 540390 40448 540454
rect 40576 538762 40640 538826
rect 677056 538614 677120 538678
rect 40960 536838 41024 536902
rect 41344 534766 41408 534830
rect 40768 534470 40832 534534
rect 41920 533642 41984 533646
rect 41920 533586 41932 533642
rect 41932 533586 41984 533642
rect 41920 533582 41984 533586
rect 41152 531362 41216 531426
rect 41536 530622 41600 530686
rect 41728 530090 41792 530094
rect 41728 530034 41780 530090
rect 41780 530034 41792 530090
rect 41728 530030 41792 530034
rect 42304 529290 42368 529354
rect 42496 527662 42560 527726
rect 42112 527130 42176 527134
rect 42112 527074 42124 527130
rect 42124 527074 42176 527130
rect 42112 527070 42176 527074
rect 42688 526478 42752 526542
rect 674560 521002 674624 521066
rect 675904 520410 675968 520474
rect 674176 519818 674240 519882
rect 674944 519670 675008 519734
rect 675520 518930 675584 518994
rect 675712 518338 675776 518402
rect 676096 518190 676160 518254
rect 675136 478230 675200 478294
rect 676288 477786 676352 477850
rect 674368 477046 674432 477110
rect 674752 476602 674816 476666
rect 675328 476158 675392 476222
rect 673984 475122 674048 475186
rect 676864 473494 676928 473558
rect 677056 473494 677120 473558
rect 42496 471570 42560 471634
rect 40576 471274 40640 471338
rect 42688 470830 42752 470894
rect 42304 470090 42368 470154
rect 41920 469498 41984 469562
rect 40384 469350 40448 469414
rect 42112 468610 42176 468674
rect 41728 468018 41792 468082
rect 41536 467722 41600 467786
rect 40960 467278 41024 467342
rect 41344 466834 41408 466898
rect 41152 466242 41216 466306
rect 40768 465798 40832 465862
rect 41536 424358 41600 424422
rect 41920 424210 41984 424274
rect 42112 423618 42176 423682
rect 41152 422878 41216 422942
rect 42688 422730 42752 422794
rect 40768 421398 40832 421462
rect 40960 420954 41024 421018
rect 41344 420510 41408 420574
rect 41728 419770 41792 419834
rect 40384 419326 40448 419390
rect 42496 418734 42560 418798
rect 40576 417846 40640 417910
rect 41920 411690 41984 411694
rect 41920 411634 41932 411690
rect 41932 411634 41984 411690
rect 41920 411630 41984 411634
rect 41728 411482 41792 411546
rect 41728 411038 41792 411102
rect 40576 408374 40640 408438
rect 41728 407990 41792 407994
rect 41728 407934 41780 407990
rect 41780 407934 41792 407990
rect 41728 407930 41792 407934
rect 42496 407338 42560 407402
rect 42688 406450 42752 406514
rect 40384 404230 40448 404294
rect 41344 403638 41408 403702
rect 40960 402898 41024 402962
rect 41152 402306 41216 402370
rect 41920 400294 41984 400298
rect 41920 400238 41932 400294
rect 41932 400238 41984 400294
rect 41920 400234 41984 400238
rect 40768 399790 40832 399854
rect 42112 399406 42176 399410
rect 42112 399350 42164 399406
rect 42164 399350 42176 399406
rect 42112 399346 42176 399350
rect 673984 394610 674048 394674
rect 674368 393278 674432 393342
rect 674176 392538 674240 392602
rect 674560 391650 674624 391714
rect 40384 381290 40448 381354
rect 42112 380994 42176 381058
rect 42688 380402 42752 380466
rect 40960 379662 41024 379726
rect 42304 379514 42368 379578
rect 40768 378182 40832 378246
rect 41152 377738 41216 377802
rect 41344 377248 41408 377312
rect 40960 376702 41024 376766
rect 42496 376702 42560 376766
rect 41920 376554 41984 376618
rect 40576 375814 40640 375878
rect 41536 375222 41600 375286
rect 41728 375074 41792 375138
rect 42112 368474 42176 368478
rect 42112 368418 42124 368474
rect 42124 368418 42176 368474
rect 42112 368414 42176 368418
rect 674560 367230 674624 367294
rect 41728 365218 41792 365222
rect 41728 365162 41780 365218
rect 41780 365162 41792 365218
rect 41728 365158 41792 365162
rect 41920 364626 41984 364630
rect 41920 364570 41972 364626
rect 41972 364570 41984 364626
rect 41920 364566 41984 364570
rect 41536 364122 41600 364186
rect 42304 363530 42368 363594
rect 40576 361014 40640 361078
rect 41344 360422 41408 360486
rect 40960 359682 41024 359746
rect 42496 358942 42560 359006
rect 40384 357166 40448 357230
rect 40768 356574 40832 356638
rect 42688 356130 42752 356194
rect 673984 350506 674048 350570
rect 674560 349618 674624 349682
rect 674368 349470 674432 349534
rect 675520 349470 675584 349534
rect 675328 349026 675392 349090
rect 674176 348582 674240 348646
rect 674368 347990 674432 348054
rect 675136 347546 675200 347610
rect 673984 346066 674048 346130
rect 674752 345474 674816 345538
rect 674944 343254 675008 343318
rect 675712 339702 675776 339766
rect 676672 339258 676736 339322
rect 676480 338814 676544 338878
rect 42880 338370 42944 338434
rect 40384 337482 40448 337546
rect 40576 337038 40640 337102
rect 42304 336890 42368 336954
rect 42496 336298 42560 336362
rect 40768 334966 40832 335030
rect 41152 334522 41216 334586
rect 40960 334078 41024 334142
rect 675136 333930 675200 333994
rect 41536 333486 41600 333550
rect 42112 333338 42176 333402
rect 41344 332598 41408 332662
rect 41920 332376 41984 332440
rect 673984 332302 674048 332366
rect 41728 331858 41792 331922
rect 674944 331118 675008 331182
rect 674752 327862 674816 327926
rect 40384 325050 40448 325114
rect 675712 324962 675776 324966
rect 675712 324906 675724 324962
rect 675724 324906 675776 324962
rect 675712 324902 675776 324906
rect 41536 323274 41600 323338
rect 676480 322978 676544 323042
rect 41728 321854 41792 321858
rect 41728 321798 41780 321854
rect 41780 321798 41792 321854
rect 41728 321794 41792 321798
rect 42112 321262 42176 321266
rect 42112 321206 42124 321262
rect 42124 321206 42176 321262
rect 42112 321202 42176 321206
rect 676672 321202 676736 321266
rect 41920 320818 41984 320822
rect 41920 320762 41932 320818
rect 41932 320762 41984 320818
rect 41920 320758 41984 320762
rect 42496 319870 42560 319934
rect 41344 317650 41408 317714
rect 40960 316762 41024 316826
rect 41152 316170 41216 316234
rect 41344 315578 41408 315642
rect 674560 313950 674624 314014
rect 42880 313802 42944 313866
rect 40768 313210 40832 313274
rect 40576 312618 40640 312682
rect 675328 303442 675392 303506
rect 674368 302554 674432 302618
rect 675712 301518 675776 301582
rect 674176 300630 674240 300694
rect 675904 300482 675968 300546
rect 676480 299742 676544 299806
rect 675136 299594 675200 299658
rect 674368 299002 674432 299066
rect 676288 297670 676352 297734
rect 675328 297522 675392 297586
rect 674752 297078 674816 297142
rect 676096 296190 676160 296254
rect 675520 295598 675584 295662
rect 40576 294858 40640 294922
rect 676864 294710 676928 294774
rect 42304 294562 42368 294626
rect 42688 294118 42752 294182
rect 40960 293378 41024 293442
rect 42496 293082 42560 293146
rect 40768 291898 40832 291962
rect 41344 291306 41408 291370
rect 41152 290862 41216 290926
rect 675904 290566 675968 290630
rect 41536 290270 41600 290334
rect 42112 290122 42176 290186
rect 40384 289382 40448 289446
rect 675712 289738 675776 289742
rect 675712 289682 675764 289738
rect 675764 289682 675776 289738
rect 675712 289678 675776 289682
rect 41920 289160 41984 289224
rect 41728 288642 41792 288706
rect 676480 287902 676544 287966
rect 676288 287458 676352 287522
rect 675328 286926 675392 286930
rect 675328 286870 675380 286926
rect 675380 286870 675392 286926
rect 675328 286866 675392 286870
rect 675136 283758 675200 283822
rect 675520 282930 675584 282934
rect 675520 282874 675572 282930
rect 675572 282874 675584 282930
rect 675520 282870 675584 282874
rect 42304 281834 42368 281898
rect 676864 282278 676928 282342
rect 676096 281834 676160 281898
rect 674752 280650 674816 280714
rect 41536 280058 41600 280122
rect 674176 278874 674240 278938
rect 41728 278786 41792 278790
rect 41728 278730 41780 278786
rect 41780 278730 41792 278786
rect 41728 278726 41792 278730
rect 674944 278578 675008 278642
rect 42112 278046 42176 278050
rect 42112 277990 42124 278046
rect 42124 277990 42176 278046
rect 42112 277986 42176 277990
rect 41920 277602 41984 277606
rect 41920 277546 41932 277602
rect 41932 277546 41984 277602
rect 41920 277542 41984 277546
rect 40576 277394 40640 277458
rect 41920 277394 41984 277458
rect 674368 276950 674432 277014
rect 42496 276654 42560 276718
rect 40384 274434 40448 274498
rect 41152 273546 41216 273610
rect 41344 273250 41408 273314
rect 40960 272362 41024 272426
rect 41920 270646 41984 270650
rect 41920 270590 41932 270646
rect 41932 270590 41984 270646
rect 41920 270586 41984 270590
rect 40768 269994 40832 270058
rect 42688 269550 42752 269614
rect 674368 266590 674432 266654
rect 674176 266442 674240 266506
rect 676288 266294 676352 266358
rect 674560 260966 674624 261030
rect 676288 260226 676352 260290
rect 673984 260078 674048 260142
rect 674944 258006 675008 258070
rect 675712 257044 675776 257108
rect 675136 256526 675200 256590
rect 675904 253566 675968 253630
rect 40576 251642 40640 251706
rect 42112 251346 42176 251410
rect 42688 250902 42752 250966
rect 41344 250162 41408 250226
rect 42880 249866 42944 249930
rect 674752 249274 674816 249338
rect 40768 248682 40832 248746
rect 41152 248090 41216 248154
rect 676672 247942 676736 248006
rect 676480 247794 676544 247858
rect 40960 247646 41024 247710
rect 41920 247498 41984 247562
rect 42496 246906 42560 246970
rect 41536 246166 41600 246230
rect 42304 246018 42368 246082
rect 41728 245426 41792 245490
rect 675712 243710 675776 243714
rect 675712 243654 675724 243710
rect 675724 243654 675776 243710
rect 675712 243650 675776 243654
rect 675136 239062 675200 239126
rect 42112 238678 42176 238682
rect 42112 238622 42124 238678
rect 42124 238622 42176 238678
rect 42112 238618 42176 238622
rect 42112 238470 42176 238534
rect 42688 238470 42752 238534
rect 675904 238026 675968 238090
rect 41920 236902 41984 236906
rect 41920 236846 41932 236902
rect 41932 236846 41984 236902
rect 41920 236842 41984 236846
rect 40576 236694 40640 236758
rect 41920 236694 41984 236758
rect 397120 236990 397184 237054
rect 397504 236990 397568 237054
rect 397696 236694 397760 236758
rect 407296 236694 407360 236758
rect 397120 236250 397184 236314
rect 407680 236250 407744 236314
rect 413632 236102 413696 236166
rect 414016 236102 414080 236166
rect 676480 235954 676544 236018
rect 41728 235570 41792 235574
rect 41728 235514 41780 235570
rect 41780 235514 41792 235570
rect 41728 235510 41792 235514
rect 42496 234770 42560 234834
rect 674944 234474 675008 234538
rect 42304 234326 42368 234390
rect 42880 233586 42944 233650
rect 676672 232550 676736 232614
rect 41536 231218 41600 231282
rect 40960 230330 41024 230394
rect 41152 230034 41216 230098
rect 41344 229294 41408 229358
rect 41920 227430 41984 227434
rect 41920 227374 41932 227430
rect 41932 227374 41984 227430
rect 41920 227370 41984 227374
rect 40768 226778 40832 226842
rect 42112 226394 42176 226398
rect 42112 226338 42164 226394
rect 42164 226338 42176 226394
rect 42112 226334 42176 226338
rect 674560 218490 674624 218554
rect 674176 218342 674240 218406
rect 674560 218342 674624 218406
rect 674176 218046 674240 218110
rect 673984 217454 674048 217518
rect 673984 217306 674048 217370
rect 674560 217306 674624 217370
rect 674368 217010 674432 217074
rect 674752 216862 674816 216926
rect 673984 215974 674048 216038
rect 674560 214642 674624 214706
rect 674752 213458 674816 213522
rect 675136 210498 675200 210562
rect 42112 208722 42176 208786
rect 41536 207834 41600 207898
rect 41920 207686 41984 207750
rect 674944 209018 675008 209082
rect 40960 206946 41024 207010
rect 40576 206354 40640 206418
rect 40768 205466 40832 205530
rect 41344 204874 41408 204938
rect 41152 204430 41216 204494
rect 40384 203986 40448 204050
rect 42496 203690 42560 203754
rect 675712 204726 675776 204790
rect 675904 204578 675968 204642
rect 42688 202950 42752 203014
rect 41728 202802 41792 202866
rect 42304 202210 42368 202274
rect 674176 197622 674240 197686
rect 673984 197178 674048 197242
rect 41536 195402 41600 195466
rect 674752 195106 674816 195170
rect 675136 193922 675200 193986
rect 40384 193626 40448 193690
rect 42304 192294 42368 192358
rect 674944 193034 675008 193098
rect 675904 192146 675968 192210
rect 42496 191702 42560 191766
rect 41728 191170 41792 191174
rect 41728 191114 41780 191170
rect 41780 191114 41792 191170
rect 41728 191110 41792 191114
rect 40576 190370 40640 190434
rect 42688 188002 42752 188066
rect 674560 189926 674624 189990
rect 675712 188506 675776 188510
rect 675712 188450 675764 188506
rect 675764 188450 675776 188506
rect 675712 188446 675776 188450
rect 41152 187114 41216 187178
rect 41344 186818 41408 186882
rect 40960 185930 41024 185994
rect 42112 184214 42176 184218
rect 42112 184158 42164 184214
rect 42164 184158 42176 184214
rect 42112 184154 42176 184158
rect 40768 183562 40832 183626
rect 41920 183178 41984 183182
rect 41920 183122 41932 183178
rect 41932 183122 41984 183178
rect 41920 183118 41984 183122
rect 673984 172758 674048 172822
rect 673984 172018 674048 172082
rect 674368 171426 674432 171490
rect 674368 170982 674432 171046
rect 674176 170538 674240 170602
rect 676288 169206 676352 169270
rect 676096 168614 676160 168678
rect 675520 168022 675584 168086
rect 674560 167282 674624 167346
rect 674368 166986 674432 167050
rect 675712 166542 675776 166606
rect 675328 165654 675392 165718
rect 675904 165506 675968 165570
rect 674944 165062 675008 165126
rect 674752 164470 674816 164534
rect 675136 163582 675200 163646
rect 676864 162694 676928 162758
rect 676096 158106 676160 158170
rect 675712 157722 675776 157726
rect 675712 157666 675764 157722
rect 675764 157666 675776 157722
rect 675712 157662 675776 157666
rect 676288 156922 676352 156986
rect 675520 155206 675584 155210
rect 675520 155150 675532 155206
rect 675532 155150 675584 155206
rect 675520 155146 675584 155150
rect 675328 154466 675392 154470
rect 675328 154410 675380 154466
rect 675380 154410 675392 154466
rect 675328 154406 675392 154410
rect 675904 153814 675968 153878
rect 676864 152630 676928 152694
rect 674560 150854 674624 150918
rect 675136 150262 675200 150326
rect 674752 149522 674816 149586
rect 674944 147894 675008 147958
rect 674368 143898 674432 143962
rect 673984 128358 674048 128422
rect 674176 127322 674240 127386
rect 675520 125398 675584 125462
rect 675904 123844 675968 123908
rect 674176 123326 674240 123390
rect 675712 120810 675776 120874
rect 676480 115630 676544 115694
rect 676672 115186 676736 115250
rect 675520 112138 675584 112142
rect 675520 112082 675572 112138
rect 675572 112082 675584 112138
rect 675520 112078 675584 112082
rect 675904 110894 675968 110958
rect 674176 106454 674240 106518
rect 675712 103554 675776 103558
rect 675712 103498 675724 103554
rect 675724 103498 675776 103554
rect 675712 103494 675776 103498
rect 676480 101570 676544 101634
rect 676672 99794 676736 99858
rect 417472 40446 417536 40510
rect 417664 40446 417728 40510
<< metal4 >>
rect 673983 873454 674049 873455
rect 673983 873390 673984 873454
rect 674048 873390 674049 873454
rect 673983 873389 674049 873390
rect 673986 852587 674046 873389
rect 673983 852586 674049 852587
rect 673983 852522 673984 852586
rect 674048 852522 674049 852586
rect 673983 852521 674049 852522
rect 40383 815142 40449 815143
rect 40383 815078 40384 815142
rect 40448 815078 40449 815142
rect 40383 815077 40449 815078
rect 40386 771927 40446 815077
rect 40575 814106 40641 814107
rect 40575 814042 40576 814106
rect 40640 814042 40641 814106
rect 40575 814041 40641 814042
rect 40578 772371 40638 814041
rect 40767 813070 40833 813071
rect 40767 813006 40768 813070
rect 40832 813006 40833 813070
rect 40767 813005 40833 813006
rect 40770 793979 40830 813005
rect 41535 805078 41601 805079
rect 41535 805014 41536 805078
rect 41600 805014 41601 805078
rect 41535 805013 41601 805014
rect 40767 793978 40833 793979
rect 40767 793914 40768 793978
rect 40832 793914 40833 793978
rect 40767 793913 40833 793914
rect 41538 786431 41598 805013
rect 41919 801082 41985 801083
rect 41919 801018 41920 801082
rect 41984 801018 41985 801082
rect 41919 801017 41985 801018
rect 41922 798863 41982 801017
rect 42495 800786 42561 800787
rect 42495 800722 42496 800786
rect 42560 800722 42561 800786
rect 42495 800721 42561 800722
rect 42303 800638 42369 800639
rect 42303 800574 42304 800638
rect 42368 800574 42369 800638
rect 42303 800573 42369 800574
rect 41919 798862 41985 798863
rect 41919 798798 41920 798862
rect 41984 798798 41985 798862
rect 41919 798797 41985 798798
rect 42306 790279 42366 800573
rect 42498 800491 42558 800721
rect 42495 800490 42561 800491
rect 42495 800426 42496 800490
rect 42560 800426 42561 800490
rect 42495 800425 42561 800426
rect 42303 790278 42369 790279
rect 42303 790214 42304 790278
rect 42368 790214 42369 790278
rect 42303 790213 42369 790214
rect 41535 786430 41601 786431
rect 41535 786366 41536 786430
rect 41600 786366 41601 786430
rect 41535 786365 41601 786366
rect 674751 774590 674817 774591
rect 674751 774526 674752 774590
rect 674816 774526 674817 774590
rect 674751 774525 674817 774526
rect 674559 773702 674625 773703
rect 674559 773638 674560 773702
rect 674624 773638 674625 773702
rect 674559 773637 674625 773638
rect 40575 772370 40641 772371
rect 40575 772306 40576 772370
rect 40640 772306 40641 772370
rect 40575 772305 40641 772306
rect 40191 771926 40257 771927
rect 40191 771862 40192 771926
rect 40256 771862 40257 771926
rect 40191 771861 40257 771862
rect 40383 771926 40449 771927
rect 40383 771862 40384 771926
rect 40448 771862 40449 771926
rect 40383 771861 40449 771862
rect 40194 771591 40254 771861
rect 40194 771531 40446 771591
rect 40386 728711 40446 771531
rect 40575 770890 40641 770891
rect 40575 770826 40576 770890
rect 40640 770826 40641 770890
rect 40575 770825 40641 770826
rect 40578 729303 40638 770825
rect 40767 769854 40833 769855
rect 40767 769790 40768 769854
rect 40832 769790 40833 769854
rect 40767 769789 40833 769790
rect 40770 748839 40830 769789
rect 674367 769410 674433 769411
rect 674367 769346 674368 769410
rect 674432 769346 674433 769410
rect 674367 769345 674433 769346
rect 41343 768966 41409 768967
rect 41343 768902 41344 768966
rect 41408 768902 41409 768966
rect 41343 768901 41409 768902
rect 41151 760234 41217 760235
rect 41151 760170 41152 760234
rect 41216 760170 41217 760234
rect 41151 760169 41217 760170
rect 40767 748838 40833 748839
rect 40767 748774 40768 748838
rect 40832 748774 40833 748838
rect 40767 748773 40833 748774
rect 41154 747063 41214 760169
rect 41346 747359 41406 768901
rect 42111 758014 42177 758015
rect 42111 757950 42112 758014
rect 42176 757950 42177 758014
rect 42111 757949 42177 757950
rect 42114 751207 42174 757949
rect 42303 757866 42369 757867
rect 42303 757802 42304 757866
rect 42368 757802 42369 757866
rect 42303 757801 42369 757802
rect 42306 752539 42366 757801
rect 42303 752538 42369 752539
rect 42303 752474 42304 752538
rect 42368 752474 42369 752538
rect 42303 752473 42369 752474
rect 42111 751206 42177 751207
rect 42111 751142 42112 751206
rect 42176 751142 42177 751206
rect 42111 751141 42177 751142
rect 41343 747358 41409 747359
rect 41343 747294 41344 747358
rect 41408 747294 41409 747358
rect 41343 747293 41409 747294
rect 41151 747062 41217 747063
rect 41151 746998 41152 747062
rect 41216 746998 41217 747062
rect 41151 746997 41217 746998
rect 40575 729302 40641 729303
rect 40575 729238 40576 729302
rect 40640 729238 40641 729302
rect 40575 729237 40641 729238
rect 40383 728710 40449 728711
rect 40383 728646 40384 728710
rect 40448 728646 40449 728710
rect 40383 728645 40449 728646
rect 40578 727675 40638 729237
rect 40575 727674 40641 727675
rect 40575 727610 40576 727674
rect 40640 727610 40641 727674
rect 40575 727609 40641 727610
rect 673983 725898 674049 725899
rect 673983 725834 673984 725898
rect 674048 725834 674049 725898
rect 673983 725833 674049 725834
rect 41151 725750 41217 725751
rect 41151 725686 41152 725750
rect 41216 725686 41217 725750
rect 41151 725685 41217 725686
rect 40959 723826 41025 723827
rect 40959 723762 40960 723826
rect 41024 723762 41025 723826
rect 40959 723761 41025 723762
rect 40383 717758 40449 717759
rect 40383 717694 40384 717758
rect 40448 717694 40449 717758
rect 40383 717693 40449 717694
rect 40386 701331 40446 717693
rect 40767 717018 40833 717019
rect 40767 716954 40768 717018
rect 40832 716954 40833 717018
rect 40767 716953 40833 716954
rect 40575 716870 40641 716871
rect 40575 716806 40576 716870
rect 40640 716806 40641 716870
rect 40575 716805 40641 716806
rect 40578 708879 40638 716805
rect 40575 708878 40641 708879
rect 40575 708814 40576 708878
rect 40640 708814 40641 708878
rect 40575 708813 40641 708814
rect 40770 708583 40830 716953
rect 40767 708582 40833 708583
rect 40767 708518 40768 708582
rect 40832 708518 40833 708582
rect 40767 708517 40833 708518
rect 40962 705919 41022 723761
rect 40959 705918 41025 705919
rect 40959 705854 40960 705918
rect 41024 705854 41025 705918
rect 40959 705853 41025 705854
rect 41154 705475 41214 725685
rect 42303 718646 42369 718647
rect 42303 718582 42304 718646
rect 42368 718582 42369 718646
rect 42303 718581 42369 718582
rect 42306 708731 42366 718581
rect 42303 708730 42369 708731
rect 42303 708666 42304 708730
rect 42368 708666 42369 708730
rect 42303 708665 42369 708666
rect 41151 705474 41217 705475
rect 41151 705410 41152 705474
rect 41216 705410 41217 705474
rect 41151 705409 41217 705410
rect 40383 701330 40449 701331
rect 40383 701266 40384 701330
rect 40448 701266 40449 701330
rect 40383 701265 40449 701266
rect 40383 685494 40449 685495
rect 40383 685430 40384 685494
rect 40448 685430 40449 685494
rect 40383 685429 40449 685430
rect 40386 650910 40446 685429
rect 40767 683422 40833 683423
rect 40767 683358 40768 683422
rect 40832 683358 40833 683422
rect 40767 683357 40833 683358
rect 40575 682534 40641 682535
rect 40575 682470 40576 682534
rect 40640 682470 40641 682534
rect 40575 682469 40641 682470
rect 40578 661519 40638 682469
rect 40770 664331 40830 683357
rect 41151 681942 41217 681943
rect 41151 681878 41152 681942
rect 41216 681878 41217 681942
rect 41151 681877 41217 681878
rect 40959 680462 41025 680463
rect 40959 680398 40960 680462
rect 41024 680398 41025 680462
rect 40959 680397 41025 680398
rect 40767 664330 40833 664331
rect 40767 664266 40768 664330
rect 40832 664266 40833 664330
rect 40767 664265 40833 664266
rect 40962 664035 41022 680397
rect 40959 664034 41025 664035
rect 40959 663970 40960 664034
rect 41024 663970 41025 664034
rect 40959 663969 41025 663970
rect 41154 662555 41214 681877
rect 41919 681794 41985 681795
rect 41919 681730 41920 681794
rect 41984 681730 41985 681794
rect 41919 681729 41985 681730
rect 41727 678834 41793 678835
rect 41727 678770 41728 678834
rect 41792 678770 41793 678834
rect 41727 678769 41793 678770
rect 41535 677502 41601 677503
rect 41535 677438 41536 677502
rect 41600 677438 41601 677502
rect 41535 677437 41601 677438
rect 41538 668623 41598 677437
rect 41535 668622 41601 668623
rect 41535 668558 41536 668622
rect 41600 668558 41601 668622
rect 41535 668557 41601 668558
rect 41730 668327 41790 678769
rect 41922 668475 41982 681729
rect 42303 680314 42369 680315
rect 42303 680250 42304 680314
rect 42368 680250 42369 680314
rect 42303 680249 42369 680250
rect 42111 679722 42177 679723
rect 42111 679658 42112 679722
rect 42176 679658 42177 679722
rect 42111 679657 42177 679658
rect 42306 679710 42366 680249
rect 41919 668474 41985 668475
rect 41919 668410 41920 668474
rect 41984 668410 41985 668474
rect 41919 668409 41985 668410
rect 41727 668326 41793 668327
rect 41727 668262 41728 668326
rect 41792 668262 41793 668326
rect 41727 668261 41793 668262
rect 42114 665367 42174 679657
rect 42306 679650 42558 679710
rect 42303 678242 42369 678243
rect 42303 678178 42304 678242
rect 42368 678178 42369 678242
rect 42303 678177 42369 678178
rect 42306 666255 42366 678177
rect 42303 666254 42369 666255
rect 42303 666190 42304 666254
rect 42368 666190 42369 666254
rect 42303 666189 42369 666190
rect 42498 665515 42558 679650
rect 42495 665514 42561 665515
rect 42495 665450 42496 665514
rect 42560 665450 42561 665514
rect 42495 665449 42561 665450
rect 42111 665366 42177 665367
rect 42111 665302 42112 665366
rect 42176 665302 42177 665366
rect 42111 665301 42177 665302
rect 41151 662554 41217 662555
rect 41151 662490 41152 662554
rect 41216 662490 41217 662554
rect 41151 662489 41217 662490
rect 40575 661518 40641 661519
rect 40575 661454 40576 661518
rect 40640 661454 40641 661518
rect 40575 661453 40641 661454
rect 40386 650850 40638 650910
rect 40578 642279 40638 650850
rect 673986 650567 674046 725833
rect 674370 693191 674430 769345
rect 674562 695855 674622 773637
rect 674754 697779 674814 774525
rect 676095 773110 676161 773111
rect 676095 773046 676096 773110
rect 676160 773046 676161 773110
rect 676095 773045 676161 773046
rect 675903 770742 675969 770743
rect 675903 770678 675904 770742
rect 675968 770678 675969 770742
rect 675903 770677 675969 770678
rect 675519 770002 675585 770003
rect 675519 769938 675520 770002
rect 675584 769938 675585 770002
rect 675519 769937 675585 769938
rect 674943 729894 675009 729895
rect 674943 729830 674944 729894
rect 675008 729830 675009 729894
rect 674943 729829 675009 729830
rect 674751 697778 674817 697779
rect 674751 697714 674752 697778
rect 674816 697714 674817 697778
rect 674751 697713 674817 697714
rect 674559 695854 674625 695855
rect 674559 695790 674560 695854
rect 674624 695790 674625 695854
rect 674559 695789 674625 695790
rect 674367 693190 674433 693191
rect 674367 693126 674368 693190
rect 674432 693126 674433 693190
rect 674367 693125 674433 693126
rect 674175 685642 674241 685643
rect 674175 685578 674176 685642
rect 674240 685578 674241 685642
rect 674175 685577 674241 685578
rect 673983 650566 674049 650567
rect 673983 650502 673984 650566
rect 674048 650502 674049 650566
rect 673983 650501 674049 650502
rect 40383 642278 40449 642279
rect 40383 642214 40384 642278
rect 40448 642214 40449 642278
rect 40383 642213 40449 642214
rect 40575 642278 40641 642279
rect 40575 642214 40576 642278
rect 40640 642214 40641 642278
rect 40575 642213 40641 642214
rect 40386 601727 40446 642213
rect 40767 640354 40833 640355
rect 40767 640290 40768 640354
rect 40832 640290 40833 640354
rect 40767 640289 40833 640290
rect 40575 639318 40641 639319
rect 40575 639254 40576 639318
rect 40640 639254 40641 639318
rect 40575 639253 40641 639254
rect 40578 617711 40638 639253
rect 40770 621411 40830 640289
rect 673983 640206 674049 640207
rect 673983 640142 673984 640206
rect 674048 640142 674049 640206
rect 673983 640141 674049 640142
rect 41343 638726 41409 638727
rect 41343 638662 41344 638726
rect 41408 638662 41409 638726
rect 41343 638661 41409 638662
rect 40767 621410 40833 621411
rect 40767 621346 40768 621410
rect 40832 621346 40833 621410
rect 40767 621345 40833 621346
rect 40575 617710 40641 617711
rect 40575 617646 40576 617710
rect 40640 617646 40641 617710
rect 40575 617645 40641 617646
rect 41346 616675 41406 638661
rect 42687 638578 42753 638579
rect 42687 638514 42688 638578
rect 42752 638514 42753 638578
rect 42687 638513 42753 638514
rect 42303 637246 42369 637247
rect 42303 637182 42304 637246
rect 42368 637182 42369 637246
rect 42303 637181 42369 637182
rect 42111 636506 42177 636507
rect 42111 636442 42112 636506
rect 42176 636442 42177 636506
rect 42111 636441 42177 636442
rect 41727 635618 41793 635619
rect 41727 635554 41728 635618
rect 41792 635554 41793 635618
rect 41727 635553 41793 635554
rect 41535 634286 41601 634287
rect 41535 634222 41536 634286
rect 41600 634222 41601 634286
rect 41535 634221 41601 634222
rect 41538 625999 41598 634221
rect 41535 625998 41601 625999
rect 41535 625934 41536 625998
rect 41600 625934 41601 625998
rect 41535 625933 41601 625934
rect 41730 625111 41790 635553
rect 41919 635026 41985 635027
rect 41919 634962 41920 635026
rect 41984 634962 41985 635026
rect 41919 634961 41985 634962
rect 41727 625110 41793 625111
rect 41727 625046 41728 625110
rect 41792 625046 41793 625110
rect 41727 625045 41793 625046
rect 41922 622151 41982 634961
rect 42114 623927 42174 636441
rect 42111 623926 42177 623927
rect 42111 623862 42112 623926
rect 42176 623862 42177 623926
rect 42111 623861 42177 623862
rect 41919 622150 41985 622151
rect 41919 622086 41920 622150
rect 41984 622086 41985 622150
rect 41919 622085 41985 622086
rect 42306 622003 42366 637181
rect 42303 622002 42369 622003
rect 42303 621938 42304 622002
rect 42368 621938 42369 622002
rect 42303 621937 42369 621938
rect 42690 620819 42750 638513
rect 43071 637098 43137 637099
rect 43071 637034 43072 637098
rect 43136 637034 43137 637098
rect 43071 637033 43137 637034
rect 42687 620818 42753 620819
rect 42687 620754 42688 620818
rect 42752 620754 42753 620818
rect 42687 620753 42753 620754
rect 43074 617267 43134 637033
rect 43071 617266 43137 617267
rect 43071 617202 43072 617266
rect 43136 617202 43137 617266
rect 43071 617201 43137 617202
rect 41343 616674 41409 616675
rect 41343 616610 41344 616674
rect 41408 616610 41409 616674
rect 41343 616609 41409 616610
rect 40383 601726 40449 601727
rect 40383 601662 40384 601726
rect 40448 601662 40449 601726
rect 40383 601661 40449 601662
rect 40575 597138 40641 597139
rect 40575 597074 40576 597138
rect 40640 597074 40641 597138
rect 40575 597073 40641 597074
rect 40383 596102 40449 596103
rect 40383 596038 40384 596102
rect 40448 596038 40449 596102
rect 40383 596037 40449 596038
rect 40386 573903 40446 596037
rect 40578 576419 40638 597073
rect 40767 595658 40833 595659
rect 40767 595594 40768 595658
rect 40832 595594 40833 595658
rect 40767 595593 40833 595594
rect 40575 576418 40641 576419
rect 40575 576354 40576 576418
rect 40640 576354 40641 576418
rect 40575 576353 40641 576354
rect 40770 576123 40830 595593
rect 42879 595362 42945 595363
rect 42879 595298 42880 595362
rect 42944 595298 42945 595362
rect 42879 595297 42945 595298
rect 40959 594178 41025 594179
rect 40959 594114 40960 594178
rect 41024 594114 41025 594178
rect 40959 594113 41025 594114
rect 40962 576271 41022 594113
rect 42111 593882 42177 593883
rect 42111 593818 42112 593882
rect 42176 593818 42177 593882
rect 42111 593817 42177 593818
rect 41535 592106 41601 592107
rect 41535 592042 41536 592106
rect 41600 592042 41601 592106
rect 41535 592041 41601 592042
rect 41538 583079 41598 592041
rect 41727 591810 41793 591811
rect 41727 591746 41728 591810
rect 41792 591746 41793 591810
rect 41727 591745 41793 591746
rect 41535 583078 41601 583079
rect 41535 583014 41536 583078
rect 41600 583014 41601 583078
rect 41535 583013 41601 583014
rect 41730 578935 41790 591745
rect 41919 591440 41985 591441
rect 41919 591376 41920 591440
rect 41984 591376 41985 591440
rect 41919 591375 41985 591376
rect 41922 582635 41982 591375
rect 41919 582634 41985 582635
rect 41919 582570 41920 582634
rect 41984 582570 41985 582634
rect 41919 582569 41985 582570
rect 42114 581747 42174 593817
rect 42303 593438 42369 593439
rect 42303 593374 42304 593438
rect 42368 593374 42369 593438
rect 42303 593373 42369 593374
rect 42111 581746 42177 581747
rect 42111 581682 42112 581746
rect 42176 581682 42177 581746
rect 42111 581681 42177 581682
rect 42306 580563 42366 593373
rect 42303 580562 42369 580563
rect 42303 580498 42304 580562
rect 42368 580498 42369 580562
rect 42303 580497 42369 580498
rect 42882 579527 42942 595297
rect 42879 579526 42945 579527
rect 42879 579462 42880 579526
rect 42944 579462 42945 579526
rect 42879 579461 42945 579462
rect 41727 578934 41793 578935
rect 41727 578870 41728 578934
rect 41792 578870 41793 578934
rect 41727 578869 41793 578870
rect 40959 576270 41025 576271
rect 40959 576206 40960 576270
rect 41024 576206 41025 576270
rect 40959 576205 41025 576206
rect 40767 576122 40833 576123
rect 40767 576058 40768 576122
rect 40832 576058 40833 576122
rect 40767 576057 40833 576058
rect 40383 573902 40449 573903
rect 40383 573838 40384 573902
rect 40448 573838 40449 573902
rect 40383 573837 40449 573838
rect 673986 562063 674046 640141
rect 674178 609127 674238 685577
rect 674367 673358 674433 673359
rect 674367 673294 674368 673358
rect 674432 673294 674433 673358
rect 674367 673293 674433 673294
rect 674370 609719 674430 673293
rect 674559 671434 674625 671435
rect 674559 671370 674560 671434
rect 674624 671370 674625 671434
rect 674559 671369 674625 671370
rect 674367 609718 674433 609719
rect 674367 609654 674368 609718
rect 674432 609654 674433 609718
rect 674367 609653 674433 609654
rect 674175 609126 674241 609127
rect 674175 609062 674176 609126
rect 674240 609062 674241 609126
rect 674175 609061 674241 609062
rect 674562 607647 674622 671369
rect 674946 653527 675006 729829
rect 675327 726786 675393 726787
rect 675327 726722 675328 726786
rect 675392 726722 675393 726786
rect 675327 726721 675393 726722
rect 674943 653526 675009 653527
rect 674943 653462 674944 653526
rect 675008 653462 675009 653526
rect 674943 653461 675009 653462
rect 675330 653083 675390 726721
rect 675522 695115 675582 769937
rect 675711 728710 675777 728711
rect 675711 728646 675712 728710
rect 675776 728646 675777 728710
rect 675711 728645 675777 728646
rect 675519 695114 675585 695115
rect 675519 695050 675520 695114
rect 675584 695050 675585 695114
rect 675519 695049 675585 695050
rect 675519 682682 675585 682683
rect 675519 682618 675520 682682
rect 675584 682618 675585 682682
rect 675519 682617 675585 682618
rect 675327 653082 675393 653083
rect 675327 653018 675328 653082
rect 675392 653018 675393 653082
rect 675327 653017 675393 653018
rect 675135 640354 675201 640355
rect 675135 640290 675136 640354
rect 675200 640290 675201 640354
rect 675135 640289 675201 640290
rect 674751 638430 674817 638431
rect 674751 638366 674752 638430
rect 674816 638366 674817 638430
rect 674751 638365 674817 638366
rect 674559 607646 674625 607647
rect 674559 607582 674560 607646
rect 674624 607582 674625 607646
rect 674559 607581 674625 607582
rect 674175 597138 674241 597139
rect 674175 597074 674176 597138
rect 674240 597074 674241 597138
rect 674175 597073 674241 597074
rect 673983 562062 674049 562063
rect 673983 561998 673984 562062
rect 674048 561998 674049 562062
rect 673983 561997 674049 561998
rect 673983 552294 674049 552295
rect 673983 552230 673984 552294
rect 674048 552230 674049 552294
rect 673983 552229 674049 552230
rect 40383 540454 40449 540455
rect 40383 540390 40384 540454
rect 40448 540390 40449 540454
rect 40383 540389 40449 540390
rect 40386 469415 40446 540389
rect 40575 538826 40641 538827
rect 40575 538762 40576 538826
rect 40640 538762 40641 538826
rect 40575 538761 40641 538762
rect 40578 471339 40638 538761
rect 40959 536902 41025 536903
rect 40959 536838 40960 536902
rect 41024 536838 41025 536902
rect 40959 536837 41025 536838
rect 40767 534534 40833 534535
rect 40767 534470 40768 534534
rect 40832 534470 40833 534534
rect 40767 534469 40833 534470
rect 40575 471338 40641 471339
rect 40575 471274 40576 471338
rect 40640 471274 40641 471338
rect 40575 471273 40641 471274
rect 40383 469414 40449 469415
rect 40383 469350 40384 469414
rect 40448 469350 40449 469414
rect 40383 469349 40449 469350
rect 40770 465863 40830 534469
rect 40962 467343 41022 536837
rect 41343 534830 41409 534831
rect 41343 534766 41344 534830
rect 41408 534766 41409 534830
rect 41343 534765 41409 534766
rect 41151 531426 41217 531427
rect 41151 531362 41152 531426
rect 41216 531362 41217 531426
rect 41151 531361 41217 531362
rect 40959 467342 41025 467343
rect 40959 467278 40960 467342
rect 41024 467278 41025 467342
rect 40959 467277 41025 467278
rect 41154 466307 41214 531361
rect 41346 466899 41406 534765
rect 41919 533646 41985 533647
rect 41919 533582 41920 533646
rect 41984 533582 41985 533646
rect 41919 533581 41985 533582
rect 41535 530686 41601 530687
rect 41535 530622 41536 530686
rect 41600 530622 41601 530686
rect 41535 530621 41601 530622
rect 41538 467787 41598 530621
rect 41727 530094 41793 530095
rect 41727 530030 41728 530094
rect 41792 530030 41793 530094
rect 41727 530029 41793 530030
rect 41730 468083 41790 530029
rect 41922 469563 41982 533581
rect 42303 529354 42369 529355
rect 42303 529290 42304 529354
rect 42368 529290 42369 529354
rect 42303 529289 42369 529290
rect 42111 527134 42177 527135
rect 42111 527070 42112 527134
rect 42176 527070 42177 527134
rect 42111 527069 42177 527070
rect 41919 469562 41985 469563
rect 41919 469498 41920 469562
rect 41984 469498 41985 469562
rect 41919 469497 41985 469498
rect 42114 468675 42174 527069
rect 42306 470155 42366 529289
rect 42495 527726 42561 527727
rect 42495 527662 42496 527726
rect 42560 527662 42561 527726
rect 42495 527661 42561 527662
rect 42498 471635 42558 527661
rect 42687 526542 42753 526543
rect 42687 526478 42688 526542
rect 42752 526478 42753 526542
rect 42687 526477 42753 526478
rect 42495 471634 42561 471635
rect 42495 471570 42496 471634
rect 42560 471570 42561 471634
rect 42495 471569 42561 471570
rect 42690 470895 42750 526477
rect 673986 475187 674046 552229
rect 674178 519883 674238 597073
rect 674559 596102 674625 596103
rect 674559 596038 674560 596102
rect 674624 596038 674625 596102
rect 674559 596037 674625 596038
rect 674367 553034 674433 553035
rect 674367 552970 674368 553034
rect 674432 552970 674433 553034
rect 674367 552969 674433 552970
rect 674175 519882 674241 519883
rect 674175 519818 674176 519882
rect 674240 519818 674241 519882
rect 674175 519817 674241 519818
rect 674370 477111 674430 552969
rect 674562 521067 674622 596037
rect 674754 563543 674814 638365
rect 674943 594030 675009 594031
rect 674943 593966 674944 594030
rect 675008 593966 675009 594030
rect 674943 593965 675009 593966
rect 674751 563542 674817 563543
rect 674751 563478 674752 563542
rect 674816 563478 674817 563542
rect 674751 563477 674817 563478
rect 674751 550222 674817 550223
rect 674751 550158 674752 550222
rect 674816 550158 674817 550222
rect 674751 550157 674817 550158
rect 674559 521066 674625 521067
rect 674559 521002 674560 521066
rect 674624 521002 674625 521066
rect 674559 521001 674625 521002
rect 674367 477110 674433 477111
rect 674367 477046 674368 477110
rect 674432 477046 674433 477110
rect 674367 477045 674433 477046
rect 674754 476667 674814 550157
rect 674946 519735 675006 593965
rect 675138 565023 675198 640289
rect 675327 634138 675393 634139
rect 675327 634074 675328 634138
rect 675392 634074 675393 634138
rect 675327 634073 675393 634074
rect 675135 565022 675201 565023
rect 675135 564958 675136 565022
rect 675200 564958 675201 565022
rect 675135 564957 675201 564958
rect 675330 562951 675390 634073
rect 675522 608683 675582 682617
rect 675714 654563 675774 728645
rect 675906 695263 675966 770677
rect 676098 698963 676158 773045
rect 677055 731670 677121 731671
rect 677055 731606 677056 731670
rect 677120 731606 677121 731670
rect 677055 731605 677121 731606
rect 676287 729450 676353 729451
rect 676287 729386 676288 729450
rect 676352 729386 676353 729450
rect 676287 729385 676353 729386
rect 676095 698962 676161 698963
rect 676095 698898 676096 698962
rect 676160 698898 676161 698962
rect 676095 698897 676161 698898
rect 675903 695262 675969 695263
rect 675903 695198 675904 695262
rect 675968 695198 675969 695262
rect 675903 695197 675969 695198
rect 675903 684458 675969 684459
rect 675903 684394 675904 684458
rect 675968 684394 675969 684458
rect 675903 684393 675969 684394
rect 675711 654562 675777 654563
rect 675711 654498 675712 654562
rect 675776 654498 675777 654562
rect 675711 654497 675777 654498
rect 675906 610163 675966 684393
rect 676095 678390 676161 678391
rect 676095 678326 676096 678390
rect 676160 678326 676161 678390
rect 676095 678325 676161 678326
rect 675903 610162 675969 610163
rect 675903 610098 675904 610162
rect 675968 610098 675969 610162
rect 675903 610097 675969 610098
rect 675519 608682 675585 608683
rect 675519 608618 675520 608682
rect 675584 608618 675585 608682
rect 675519 608617 675585 608618
rect 676098 608535 676158 678325
rect 676290 651455 676350 729385
rect 676479 726194 676545 726195
rect 676479 726130 676480 726194
rect 676544 726130 676545 726194
rect 676479 726129 676545 726130
rect 676482 651455 676542 726129
rect 676863 721902 676929 721903
rect 676863 721838 676864 721902
rect 676928 721838 676929 721902
rect 676863 721837 676929 721838
rect 676287 651454 676353 651455
rect 676287 651390 676288 651454
rect 676352 651390 676353 651454
rect 676287 651389 676353 651390
rect 676479 651454 676545 651455
rect 676479 651390 676480 651454
rect 676544 651390 676545 651454
rect 676479 651389 676545 651390
rect 676866 648791 676926 721837
rect 677058 692599 677118 731605
rect 677055 692598 677121 692599
rect 677055 692534 677056 692598
rect 677120 692534 677121 692598
rect 677055 692533 677121 692534
rect 677055 676910 677121 676911
rect 677055 676846 677056 676910
rect 677120 676846 677121 676910
rect 677055 676845 677121 676846
rect 677058 649827 677118 676845
rect 677055 649826 677121 649827
rect 677055 649762 677056 649826
rect 677120 649762 677121 649826
rect 677055 649761 677121 649762
rect 676863 648790 676929 648791
rect 676863 648726 676864 648790
rect 676928 648726 676929 648790
rect 676863 648725 676929 648726
rect 676671 641686 676737 641687
rect 676671 641622 676672 641686
rect 676736 641622 676737 641686
rect 676671 641621 676737 641622
rect 676287 629106 676353 629107
rect 676287 629042 676288 629106
rect 676352 629042 676353 629106
rect 676287 629041 676353 629042
rect 676095 608534 676161 608535
rect 676095 608470 676096 608534
rect 676160 608470 676161 608534
rect 676095 608469 676161 608470
rect 675519 589738 675585 589739
rect 675519 589674 675520 589738
rect 675584 589674 675585 589738
rect 675519 589673 675585 589674
rect 675327 562950 675393 562951
rect 675327 562886 675328 562950
rect 675392 562886 675393 562950
rect 675327 562885 675393 562886
rect 675135 551702 675201 551703
rect 675135 551638 675136 551702
rect 675200 551638 675201 551702
rect 675135 551637 675201 551638
rect 674943 519734 675009 519735
rect 674943 519670 674944 519734
rect 675008 519670 675009 519734
rect 674943 519669 675009 519670
rect 675138 478295 675198 551637
rect 675327 545486 675393 545487
rect 675327 545422 675328 545486
rect 675392 545422 675393 545486
rect 675327 545421 675393 545422
rect 675135 478294 675201 478295
rect 675135 478230 675136 478294
rect 675200 478230 675201 478294
rect 675135 478229 675201 478230
rect 674751 476666 674817 476667
rect 674751 476602 674752 476666
rect 674816 476602 674817 476666
rect 674751 476601 674817 476602
rect 675330 476223 675390 545421
rect 675522 518995 675582 589673
rect 675903 584706 675969 584707
rect 675903 584642 675904 584706
rect 675968 584642 675969 584706
rect 675903 584641 675969 584642
rect 675711 582930 675777 582931
rect 675711 582866 675712 582930
rect 675776 582866 675777 582930
rect 675711 582865 675777 582866
rect 675519 518994 675585 518995
rect 675519 518930 675520 518994
rect 675584 518930 675585 518994
rect 675519 518929 675585 518930
rect 675714 518403 675774 582865
rect 675906 520475 675966 584641
rect 676095 567242 676161 567243
rect 676095 567178 676096 567242
rect 676160 567178 676161 567242
rect 676095 567177 676161 567178
rect 675903 520474 675969 520475
rect 675903 520410 675904 520474
rect 675968 520410 675969 520474
rect 675903 520409 675969 520410
rect 675711 518402 675777 518403
rect 675711 518338 675712 518402
rect 675776 518338 675777 518402
rect 675711 518337 675777 518338
rect 676098 518255 676158 567177
rect 676290 564727 676350 629041
rect 676479 627330 676545 627331
rect 676479 627266 676480 627330
rect 676544 627266 676545 627330
rect 676479 627265 676545 627266
rect 676287 564726 676353 564727
rect 676287 564662 676288 564726
rect 676352 564662 676353 564726
rect 676287 564661 676353 564662
rect 676482 562803 676542 627265
rect 676674 564283 676734 641621
rect 676863 632806 676929 632807
rect 676863 632742 676864 632806
rect 676928 632742 676929 632806
rect 676863 632741 676929 632742
rect 676671 564282 676737 564283
rect 676671 564218 676672 564282
rect 676736 564218 676737 564282
rect 676671 564217 676737 564218
rect 676479 562802 676545 562803
rect 676479 562738 676480 562802
rect 676544 562738 676545 562802
rect 676479 562737 676545 562738
rect 676866 560287 676926 632741
rect 676863 560286 676929 560287
rect 676863 560222 676864 560286
rect 676928 560222 676929 560286
rect 676863 560221 676929 560222
rect 676863 544302 676929 544303
rect 676863 544238 676864 544302
rect 676928 544238 676929 544302
rect 676863 544237 676929 544238
rect 676287 540602 676353 540603
rect 676287 540538 676288 540602
rect 676352 540538 676353 540602
rect 676287 540537 676353 540538
rect 676095 518254 676161 518255
rect 676095 518190 676096 518254
rect 676160 518190 676161 518254
rect 676095 518189 676161 518190
rect 676290 477851 676350 540537
rect 676287 477850 676353 477851
rect 676287 477786 676288 477850
rect 676352 477786 676353 477850
rect 676287 477785 676353 477786
rect 675327 476222 675393 476223
rect 675327 476158 675328 476222
rect 675392 476158 675393 476222
rect 675327 476157 675393 476158
rect 673983 475186 674049 475187
rect 673983 475122 673984 475186
rect 674048 475122 674049 475186
rect 673983 475121 674049 475122
rect 676866 473559 676926 544237
rect 677055 538678 677121 538679
rect 677055 538614 677056 538678
rect 677120 538614 677121 538678
rect 677055 538613 677121 538614
rect 677058 473559 677118 538613
rect 676863 473558 676929 473559
rect 676863 473494 676864 473558
rect 676928 473494 676929 473558
rect 676863 473493 676929 473494
rect 677055 473558 677121 473559
rect 677055 473494 677056 473558
rect 677120 473494 677121 473558
rect 677055 473493 677121 473494
rect 42687 470894 42753 470895
rect 42687 470830 42688 470894
rect 42752 470830 42753 470894
rect 42687 470829 42753 470830
rect 42303 470154 42369 470155
rect 42303 470090 42304 470154
rect 42368 470090 42369 470154
rect 42303 470089 42369 470090
rect 42111 468674 42177 468675
rect 42111 468610 42112 468674
rect 42176 468610 42177 468674
rect 42111 468609 42177 468610
rect 41727 468082 41793 468083
rect 41727 468018 41728 468082
rect 41792 468018 41793 468082
rect 41727 468017 41793 468018
rect 41535 467786 41601 467787
rect 41535 467722 41536 467786
rect 41600 467722 41601 467786
rect 41535 467721 41601 467722
rect 41343 466898 41409 466899
rect 41343 466834 41344 466898
rect 41408 466834 41409 466898
rect 41343 466833 41409 466834
rect 41151 466306 41217 466307
rect 41151 466242 41152 466306
rect 41216 466242 41217 466306
rect 41151 466241 41217 466242
rect 40767 465862 40833 465863
rect 40767 465798 40768 465862
rect 40832 465798 40833 465862
rect 40767 465797 40833 465798
rect 41535 424422 41601 424423
rect 41535 424358 41536 424422
rect 41600 424358 41601 424422
rect 41535 424357 41601 424358
rect 41151 422942 41217 422943
rect 41151 422878 41152 422942
rect 41216 422878 41217 422942
rect 41151 422877 41217 422878
rect 40767 421462 40833 421463
rect 40767 421398 40768 421462
rect 40832 421398 40833 421462
rect 40767 421397 40833 421398
rect 40383 419390 40449 419391
rect 40383 419326 40384 419390
rect 40448 419326 40449 419390
rect 40383 419325 40449 419326
rect 40386 404295 40446 419325
rect 40575 417910 40641 417911
rect 40575 417846 40576 417910
rect 40640 417846 40641 417910
rect 40575 417845 40641 417846
rect 40578 408439 40638 417845
rect 40575 408438 40641 408439
rect 40575 408374 40576 408438
rect 40640 408374 40641 408438
rect 40575 408373 40641 408374
rect 40383 404294 40449 404295
rect 40383 404230 40384 404294
rect 40448 404230 40449 404294
rect 40383 404229 40449 404230
rect 40770 399855 40830 421397
rect 40959 421018 41025 421019
rect 40959 420954 40960 421018
rect 41024 420954 41025 421018
rect 40959 420953 41025 420954
rect 40962 402963 41022 420953
rect 40959 402962 41025 402963
rect 40959 402898 40960 402962
rect 41024 402898 41025 402962
rect 40959 402897 41025 402898
rect 41154 402371 41214 422877
rect 41343 420574 41409 420575
rect 41343 420510 41344 420574
rect 41408 420510 41409 420574
rect 41343 420509 41409 420510
rect 41346 403703 41406 420509
rect 41538 411285 41598 424357
rect 41919 424274 41985 424275
rect 41919 424210 41920 424274
rect 41984 424210 41985 424274
rect 41919 424209 41985 424210
rect 41727 419834 41793 419835
rect 41727 419770 41728 419834
rect 41792 419770 41793 419834
rect 41727 419769 41793 419770
rect 41730 411547 41790 419769
rect 41922 411695 41982 424209
rect 42111 423682 42177 423683
rect 42111 423618 42112 423682
rect 42176 423618 42177 423682
rect 42111 423617 42177 423618
rect 41919 411694 41985 411695
rect 41919 411630 41920 411694
rect 41984 411630 41985 411694
rect 41919 411629 41985 411630
rect 41727 411546 41793 411547
rect 41727 411482 41728 411546
rect 41792 411482 41793 411546
rect 41727 411481 41793 411482
rect 41538 411225 41982 411285
rect 41727 411102 41793 411103
rect 41727 411038 41728 411102
rect 41792 411038 41793 411102
rect 41727 411037 41793 411038
rect 41730 407995 41790 411037
rect 41727 407994 41793 407995
rect 41727 407930 41728 407994
rect 41792 407930 41793 407994
rect 41727 407929 41793 407930
rect 41343 403702 41409 403703
rect 41343 403638 41344 403702
rect 41408 403638 41409 403702
rect 41343 403637 41409 403638
rect 41151 402370 41217 402371
rect 41151 402306 41152 402370
rect 41216 402306 41217 402370
rect 41151 402305 41217 402306
rect 41922 400299 41982 411225
rect 41919 400298 41985 400299
rect 41919 400234 41920 400298
rect 41984 400234 41985 400298
rect 41919 400233 41985 400234
rect 40767 399854 40833 399855
rect 40767 399790 40768 399854
rect 40832 399790 40833 399854
rect 40767 399789 40833 399790
rect 42114 399411 42174 423617
rect 42687 422794 42753 422795
rect 42687 422730 42688 422794
rect 42752 422730 42753 422794
rect 42687 422729 42753 422730
rect 42495 418798 42561 418799
rect 42495 418734 42496 418798
rect 42560 418734 42561 418798
rect 42495 418733 42561 418734
rect 42498 407403 42558 418733
rect 42495 407402 42561 407403
rect 42495 407338 42496 407402
rect 42560 407338 42561 407402
rect 42495 407337 42561 407338
rect 42690 406515 42750 422729
rect 42687 406514 42753 406515
rect 42687 406450 42688 406514
rect 42752 406450 42753 406514
rect 42687 406449 42753 406450
rect 42111 399410 42177 399411
rect 42111 399346 42112 399410
rect 42176 399346 42177 399410
rect 42111 399345 42177 399346
rect 673983 394674 674049 394675
rect 673983 394610 673984 394674
rect 674048 394610 674049 394674
rect 673983 394609 674049 394610
rect 40383 381354 40449 381355
rect 40383 381290 40384 381354
rect 40448 381290 40449 381354
rect 40383 381289 40449 381290
rect 40386 357231 40446 381289
rect 42111 381058 42177 381059
rect 42111 380994 42112 381058
rect 42176 380994 42177 381058
rect 42111 380993 42177 380994
rect 40959 379726 41025 379727
rect 40959 379662 40960 379726
rect 41024 379662 41025 379726
rect 40959 379661 41025 379662
rect 40767 378246 40833 378247
rect 40767 378182 40768 378246
rect 40832 378182 40833 378246
rect 40767 378181 40833 378182
rect 40575 375878 40641 375879
rect 40575 375814 40576 375878
rect 40640 375814 40641 375878
rect 40575 375813 40641 375814
rect 40578 361079 40638 375813
rect 40575 361078 40641 361079
rect 40575 361014 40576 361078
rect 40640 361014 40641 361078
rect 40575 361013 40641 361014
rect 40383 357230 40449 357231
rect 40383 357166 40384 357230
rect 40448 357166 40449 357230
rect 40383 357165 40449 357166
rect 40770 356639 40830 378181
rect 40962 376767 41022 379661
rect 41151 377802 41217 377803
rect 41151 377738 41152 377802
rect 41216 377738 41217 377802
rect 41151 377737 41217 377738
rect 40959 376766 41025 376767
rect 40959 376702 40960 376766
rect 41024 376702 41025 376766
rect 40959 376701 41025 376702
rect 41154 375987 41214 377737
rect 41343 377312 41409 377313
rect 41343 377248 41344 377312
rect 41408 377248 41409 377312
rect 41343 377247 41409 377248
rect 40962 375927 41214 375987
rect 40962 359747 41022 375927
rect 41346 360487 41406 377247
rect 41919 376618 41985 376619
rect 41919 376554 41920 376618
rect 41984 376554 41985 376618
rect 41919 376553 41985 376554
rect 41535 375286 41601 375287
rect 41535 375222 41536 375286
rect 41600 375222 41601 375286
rect 41535 375221 41601 375222
rect 41538 364187 41598 375221
rect 41727 375138 41793 375139
rect 41727 375074 41728 375138
rect 41792 375074 41793 375138
rect 41727 375073 41793 375074
rect 41730 365223 41790 375073
rect 41727 365222 41793 365223
rect 41727 365158 41728 365222
rect 41792 365158 41793 365222
rect 41727 365157 41793 365158
rect 41922 364631 41982 376553
rect 42114 368479 42174 380993
rect 42687 380466 42753 380467
rect 42687 380402 42688 380466
rect 42752 380402 42753 380466
rect 42687 380401 42753 380402
rect 42303 379578 42369 379579
rect 42303 379514 42304 379578
rect 42368 379514 42369 379578
rect 42303 379513 42369 379514
rect 42111 368478 42177 368479
rect 42111 368414 42112 368478
rect 42176 368414 42177 368478
rect 42111 368413 42177 368414
rect 41919 364630 41985 364631
rect 41919 364566 41920 364630
rect 41984 364566 41985 364630
rect 41919 364565 41985 364566
rect 41535 364186 41601 364187
rect 41535 364122 41536 364186
rect 41600 364122 41601 364186
rect 41535 364121 41601 364122
rect 42306 363595 42366 379513
rect 42495 376766 42561 376767
rect 42495 376702 42496 376766
rect 42560 376702 42561 376766
rect 42495 376701 42561 376702
rect 42303 363594 42369 363595
rect 42303 363530 42304 363594
rect 42368 363530 42369 363594
rect 42303 363529 42369 363530
rect 41343 360486 41409 360487
rect 41343 360422 41344 360486
rect 41408 360422 41409 360486
rect 41343 360421 41409 360422
rect 40959 359746 41025 359747
rect 40959 359682 40960 359746
rect 41024 359682 41025 359746
rect 40959 359681 41025 359682
rect 42498 359007 42558 376701
rect 42495 359006 42561 359007
rect 42495 358942 42496 359006
rect 42560 358942 42561 359006
rect 42495 358941 42561 358942
rect 40767 356638 40833 356639
rect 40767 356574 40768 356638
rect 40832 356574 40833 356638
rect 40767 356573 40833 356574
rect 42690 356195 42750 380401
rect 42687 356194 42753 356195
rect 42687 356130 42688 356194
rect 42752 356130 42753 356194
rect 42687 356129 42753 356130
rect 673986 350571 674046 394609
rect 674367 393342 674433 393343
rect 674367 393278 674368 393342
rect 674432 393278 674433 393342
rect 674367 393277 674433 393278
rect 674175 392602 674241 392603
rect 674175 392538 674176 392602
rect 674240 392538 674241 392602
rect 674175 392537 674241 392538
rect 673983 350570 674049 350571
rect 673983 350506 673984 350570
rect 674048 350506 674049 350570
rect 673983 350505 674049 350506
rect 674178 348647 674238 392537
rect 674370 349535 674430 393277
rect 674559 391714 674625 391715
rect 674559 391650 674560 391714
rect 674624 391650 674625 391714
rect 674559 391649 674625 391650
rect 674562 367295 674622 391649
rect 674559 367294 674625 367295
rect 674559 367230 674560 367294
rect 674624 367230 674625 367294
rect 674559 367229 674625 367230
rect 674559 349682 674625 349683
rect 674559 349618 674560 349682
rect 674624 349618 674625 349682
rect 674559 349617 674625 349618
rect 674367 349534 674433 349535
rect 674367 349470 674368 349534
rect 674432 349470 674433 349534
rect 674367 349469 674433 349470
rect 674175 348646 674241 348647
rect 674175 348582 674176 348646
rect 674240 348582 674241 348646
rect 674175 348581 674241 348582
rect 674367 348054 674433 348055
rect 674367 347990 674368 348054
rect 674432 347990 674433 348054
rect 674367 347989 674433 347990
rect 673983 346130 674049 346131
rect 673983 346066 673984 346130
rect 674048 346066 674049 346130
rect 673983 346065 674049 346066
rect 42879 338434 42945 338435
rect 42879 338370 42880 338434
rect 42944 338370 42945 338434
rect 42879 338369 42945 338370
rect 40383 337546 40449 337547
rect 40383 337482 40384 337546
rect 40448 337482 40449 337546
rect 40383 337481 40449 337482
rect 40386 325115 40446 337481
rect 40575 337102 40641 337103
rect 40575 337038 40576 337102
rect 40640 337038 40641 337102
rect 40575 337037 40641 337038
rect 40383 325114 40449 325115
rect 40383 325050 40384 325114
rect 40448 325050 40449 325114
rect 40383 325049 40449 325050
rect 40578 312683 40638 337037
rect 42303 336954 42369 336955
rect 42303 336890 42304 336954
rect 42368 336890 42369 336954
rect 42303 336889 42369 336890
rect 40767 335030 40833 335031
rect 40767 334966 40768 335030
rect 40832 334966 40833 335030
rect 40767 334965 40833 334966
rect 40770 313275 40830 334965
rect 41151 334586 41217 334587
rect 41151 334522 41152 334586
rect 41216 334522 41217 334586
rect 41151 334521 41217 334522
rect 40959 334142 41025 334143
rect 40959 334078 40960 334142
rect 41024 334078 41025 334142
rect 40959 334077 41025 334078
rect 40962 316827 41022 334077
rect 40959 316826 41025 316827
rect 40959 316762 40960 316826
rect 41024 316762 41025 316826
rect 40959 316761 41025 316762
rect 41154 316235 41214 334521
rect 41535 333550 41601 333551
rect 41535 333486 41536 333550
rect 41600 333486 41601 333550
rect 41535 333485 41601 333486
rect 41343 332662 41409 332663
rect 41343 332598 41344 332662
rect 41408 332598 41409 332662
rect 41343 332597 41409 332598
rect 41346 317715 41406 332597
rect 41538 323339 41598 333485
rect 42111 333402 42177 333403
rect 42111 333338 42112 333402
rect 42176 333338 42177 333402
rect 42111 333337 42177 333338
rect 41919 332440 41985 332441
rect 41919 332376 41920 332440
rect 41984 332376 41985 332440
rect 41919 332375 41985 332376
rect 41727 331922 41793 331923
rect 41727 331858 41728 331922
rect 41792 331858 41793 331922
rect 41727 331857 41793 331858
rect 41535 323338 41601 323339
rect 41535 323274 41536 323338
rect 41600 323274 41601 323338
rect 41535 323273 41601 323274
rect 41730 321859 41790 331857
rect 41727 321858 41793 321859
rect 41727 321794 41728 321858
rect 41792 321794 41793 321858
rect 41727 321793 41793 321794
rect 41922 320823 41982 332375
rect 42114 321267 42174 333337
rect 42111 321266 42177 321267
rect 42111 321202 42112 321266
rect 42176 321202 42177 321266
rect 42111 321201 42177 321202
rect 41919 320822 41985 320823
rect 41919 320758 41920 320822
rect 41984 320758 41985 320822
rect 41919 320757 41985 320758
rect 41343 317714 41409 317715
rect 41343 317650 41344 317714
rect 41408 317650 41409 317714
rect 41343 317649 41409 317650
rect 42306 317379 42366 336889
rect 42495 336362 42561 336363
rect 42495 336298 42496 336362
rect 42560 336298 42561 336362
rect 42495 336297 42561 336298
rect 42498 319935 42558 336297
rect 42495 319934 42561 319935
rect 42495 319870 42496 319934
rect 42560 319870 42561 319934
rect 42495 319869 42561 319870
rect 41346 317319 42366 317379
rect 41151 316234 41217 316235
rect 41151 316170 41152 316234
rect 41216 316170 41217 316234
rect 41151 316169 41217 316170
rect 41346 315643 41406 317319
rect 41343 315642 41409 315643
rect 41343 315578 41344 315642
rect 41408 315578 41409 315642
rect 41343 315577 41409 315578
rect 42882 313867 42942 338369
rect 673986 332367 674046 346065
rect 673983 332366 674049 332367
rect 673983 332302 673984 332366
rect 674048 332302 674049 332366
rect 673983 332301 674049 332302
rect 42879 313866 42945 313867
rect 42879 313802 42880 313866
rect 42944 313802 42945 313866
rect 42879 313801 42945 313802
rect 40767 313274 40833 313275
rect 40767 313210 40768 313274
rect 40832 313210 40833 313274
rect 40767 313209 40833 313210
rect 40575 312682 40641 312683
rect 40575 312618 40576 312682
rect 40640 312618 40641 312682
rect 40575 312617 40641 312618
rect 674370 302619 674430 347989
rect 674562 314015 674622 349617
rect 675519 349534 675585 349535
rect 675519 349470 675520 349534
rect 675584 349470 675585 349534
rect 675519 349469 675585 349470
rect 675327 349090 675393 349091
rect 675327 349026 675328 349090
rect 675392 349026 675393 349090
rect 675327 349025 675393 349026
rect 675135 347610 675201 347611
rect 675135 347546 675136 347610
rect 675200 347546 675201 347610
rect 675135 347545 675201 347546
rect 674751 345538 674817 345539
rect 674751 345474 674752 345538
rect 674816 345474 674817 345538
rect 674751 345473 674817 345474
rect 674754 327927 674814 345473
rect 674943 343318 675009 343319
rect 674943 343254 674944 343318
rect 675008 343254 675009 343318
rect 674943 343253 675009 343254
rect 674946 331183 675006 343253
rect 675138 333995 675198 347545
rect 675135 333994 675201 333995
rect 675135 333930 675136 333994
rect 675200 333930 675201 333994
rect 675135 333929 675201 333930
rect 674943 331182 675009 331183
rect 674943 331118 674944 331182
rect 675008 331118 675009 331182
rect 674943 331117 675009 331118
rect 674751 327926 674817 327927
rect 674751 327862 674752 327926
rect 674816 327862 674817 327926
rect 674751 327861 674817 327862
rect 674559 314014 674625 314015
rect 674559 313950 674560 314014
rect 674624 313950 674625 314014
rect 674559 313949 674625 313950
rect 675330 303507 675390 349025
rect 675327 303506 675393 303507
rect 675327 303442 675328 303506
rect 675392 303442 675393 303506
rect 675327 303441 675393 303442
rect 674367 302618 674433 302619
rect 674367 302554 674368 302618
rect 674432 302554 674433 302618
rect 674367 302553 674433 302554
rect 674175 300694 674241 300695
rect 674175 300630 674176 300694
rect 674240 300630 674241 300694
rect 674175 300629 674241 300630
rect 40575 294922 40641 294923
rect 40575 294858 40576 294922
rect 40640 294858 40641 294922
rect 40575 294857 40641 294858
rect 40383 289446 40449 289447
rect 40383 289382 40384 289446
rect 40448 289382 40449 289446
rect 40383 289381 40449 289382
rect 40386 274499 40446 289381
rect 40578 277459 40638 294857
rect 42303 294626 42369 294627
rect 42303 294562 42304 294626
rect 42368 294562 42369 294626
rect 42303 294561 42369 294562
rect 40959 293442 41025 293443
rect 40959 293378 40960 293442
rect 41024 293378 41025 293442
rect 40959 293377 41025 293378
rect 40767 291962 40833 291963
rect 40767 291898 40768 291962
rect 40832 291898 40833 291962
rect 40767 291897 40833 291898
rect 40575 277458 40641 277459
rect 40575 277394 40576 277458
rect 40640 277394 40641 277458
rect 40575 277393 40641 277394
rect 40383 274498 40449 274499
rect 40383 274434 40384 274498
rect 40448 274434 40449 274498
rect 40383 274433 40449 274434
rect 40770 270059 40830 291897
rect 40962 272427 41022 293377
rect 41343 291370 41409 291371
rect 41343 291306 41344 291370
rect 41408 291306 41409 291370
rect 41343 291305 41409 291306
rect 41151 290926 41217 290927
rect 41151 290862 41152 290926
rect 41216 290862 41217 290926
rect 41151 290861 41217 290862
rect 41154 273611 41214 290861
rect 41151 273610 41217 273611
rect 41151 273546 41152 273610
rect 41216 273546 41217 273610
rect 41151 273545 41217 273546
rect 41346 273315 41406 291305
rect 41535 290334 41601 290335
rect 41535 290270 41536 290334
rect 41600 290270 41601 290334
rect 41535 290269 41601 290270
rect 41538 280123 41598 290269
rect 42111 290186 42177 290187
rect 42111 290122 42112 290186
rect 42176 290122 42177 290186
rect 42111 290121 42177 290122
rect 41919 289224 41985 289225
rect 41919 289160 41920 289224
rect 41984 289160 41985 289224
rect 41919 289159 41985 289160
rect 41727 288706 41793 288707
rect 41727 288642 41728 288706
rect 41792 288642 41793 288706
rect 41727 288641 41793 288642
rect 41535 280122 41601 280123
rect 41535 280058 41536 280122
rect 41600 280058 41601 280122
rect 41535 280057 41601 280058
rect 41730 278791 41790 288641
rect 41727 278790 41793 278791
rect 41727 278726 41728 278790
rect 41792 278726 41793 278790
rect 41727 278725 41793 278726
rect 41922 277607 41982 289159
rect 42114 278051 42174 290121
rect 42306 281899 42366 294561
rect 42687 294182 42753 294183
rect 42687 294118 42688 294182
rect 42752 294118 42753 294182
rect 42687 294117 42753 294118
rect 42495 293146 42561 293147
rect 42495 293082 42496 293146
rect 42560 293082 42561 293146
rect 42495 293081 42561 293082
rect 42303 281898 42369 281899
rect 42303 281834 42304 281898
rect 42368 281834 42369 281898
rect 42303 281833 42369 281834
rect 42111 278050 42177 278051
rect 42111 277986 42112 278050
rect 42176 277986 42177 278050
rect 42111 277985 42177 277986
rect 41919 277606 41985 277607
rect 41919 277542 41920 277606
rect 41984 277542 41985 277606
rect 41919 277541 41985 277542
rect 41919 277458 41985 277459
rect 41919 277394 41920 277458
rect 41984 277394 41985 277458
rect 41919 277393 41985 277394
rect 41343 273314 41409 273315
rect 41343 273250 41344 273314
rect 41408 273250 41409 273314
rect 41343 273249 41409 273250
rect 40959 272426 41025 272427
rect 40959 272362 40960 272426
rect 41024 272362 41025 272426
rect 40959 272361 41025 272362
rect 41922 270651 41982 277393
rect 42498 276719 42558 293081
rect 42495 276718 42561 276719
rect 42495 276654 42496 276718
rect 42560 276654 42561 276718
rect 42495 276653 42561 276654
rect 41919 270650 41985 270651
rect 41919 270586 41920 270650
rect 41984 270586 41985 270650
rect 41919 270585 41985 270586
rect 40767 270058 40833 270059
rect 40767 269994 40768 270058
rect 40832 269994 40833 270058
rect 40767 269993 40833 269994
rect 42690 269615 42750 294117
rect 674178 278939 674238 300629
rect 675522 300063 675582 349469
rect 675711 339766 675777 339767
rect 675711 339702 675712 339766
rect 675776 339702 675777 339766
rect 675711 339701 675777 339702
rect 675714 324967 675774 339701
rect 676671 339322 676737 339323
rect 676671 339258 676672 339322
rect 676736 339258 676737 339322
rect 676671 339257 676737 339258
rect 676479 338878 676545 338879
rect 676479 338814 676480 338878
rect 676544 338814 676545 338878
rect 676479 338813 676545 338814
rect 675711 324966 675777 324967
rect 675711 324902 675712 324966
rect 675776 324902 675777 324966
rect 675711 324901 675777 324902
rect 676482 323043 676542 338813
rect 676479 323042 676545 323043
rect 676479 322978 676480 323042
rect 676544 322978 676545 323042
rect 676479 322977 676545 322978
rect 676674 321267 676734 339257
rect 676671 321266 676737 321267
rect 676671 321202 676672 321266
rect 676736 321202 676737 321266
rect 676671 321201 676737 321202
rect 675711 301582 675777 301583
rect 675711 301518 675712 301582
rect 675776 301518 675777 301582
rect 675711 301517 675777 301518
rect 674946 300003 675582 300063
rect 674367 299066 674433 299067
rect 674367 299002 674368 299066
rect 674432 299002 674433 299066
rect 674367 299001 674433 299002
rect 674175 278938 674241 278939
rect 674175 278874 674176 278938
rect 674240 278874 674241 278938
rect 674175 278873 674241 278874
rect 674370 277015 674430 299001
rect 674751 297142 674817 297143
rect 674751 297078 674752 297142
rect 674816 297078 674817 297142
rect 674751 297077 674817 297078
rect 674754 280715 674814 297077
rect 674751 280714 674817 280715
rect 674751 280650 674752 280714
rect 674816 280650 674817 280714
rect 674751 280649 674817 280650
rect 674946 278643 675006 300003
rect 675135 299658 675201 299659
rect 675135 299594 675136 299658
rect 675200 299594 675201 299658
rect 675135 299593 675201 299594
rect 675138 283823 675198 299593
rect 675327 297586 675393 297587
rect 675327 297522 675328 297586
rect 675392 297522 675393 297586
rect 675327 297521 675393 297522
rect 675330 286931 675390 297521
rect 675519 295662 675585 295663
rect 675519 295598 675520 295662
rect 675584 295598 675585 295662
rect 675519 295597 675585 295598
rect 675327 286930 675393 286931
rect 675327 286866 675328 286930
rect 675392 286866 675393 286930
rect 675327 286865 675393 286866
rect 675135 283822 675201 283823
rect 675135 283758 675136 283822
rect 675200 283758 675201 283822
rect 675135 283757 675201 283758
rect 675522 282935 675582 295597
rect 675714 289743 675774 301517
rect 675903 300546 675969 300547
rect 675903 300482 675904 300546
rect 675968 300482 675969 300546
rect 675903 300481 675969 300482
rect 675906 290631 675966 300481
rect 676479 299806 676545 299807
rect 676479 299742 676480 299806
rect 676544 299742 676545 299806
rect 676479 299741 676545 299742
rect 676287 297734 676353 297735
rect 676287 297670 676288 297734
rect 676352 297670 676353 297734
rect 676287 297669 676353 297670
rect 676095 296254 676161 296255
rect 676095 296190 676096 296254
rect 676160 296190 676161 296254
rect 676095 296189 676161 296190
rect 675903 290630 675969 290631
rect 675903 290566 675904 290630
rect 675968 290566 675969 290630
rect 675903 290565 675969 290566
rect 675711 289742 675777 289743
rect 675711 289678 675712 289742
rect 675776 289678 675777 289742
rect 675711 289677 675777 289678
rect 675519 282934 675585 282935
rect 675519 282870 675520 282934
rect 675584 282870 675585 282934
rect 675519 282869 675585 282870
rect 676098 281899 676158 296189
rect 676290 287523 676350 297669
rect 676482 287967 676542 299741
rect 676863 294774 676929 294775
rect 676863 294710 676864 294774
rect 676928 294710 676929 294774
rect 676863 294709 676929 294710
rect 676479 287966 676545 287967
rect 676479 287902 676480 287966
rect 676544 287902 676545 287966
rect 676479 287901 676545 287902
rect 676287 287522 676353 287523
rect 676287 287458 676288 287522
rect 676352 287458 676353 287522
rect 676287 287457 676353 287458
rect 676866 282343 676926 294709
rect 676863 282342 676929 282343
rect 676863 282278 676864 282342
rect 676928 282278 676929 282342
rect 676863 282277 676929 282278
rect 676095 281898 676161 281899
rect 676095 281834 676096 281898
rect 676160 281834 676161 281898
rect 676095 281833 676161 281834
rect 674943 278642 675009 278643
rect 674943 278578 674944 278642
rect 675008 278578 675009 278642
rect 674943 278577 675009 278578
rect 674367 277014 674433 277015
rect 674367 276950 674368 277014
rect 674432 276950 674433 277014
rect 674367 276949 674433 276950
rect 42687 269614 42753 269615
rect 42687 269550 42688 269614
rect 42752 269550 42753 269614
rect 42687 269549 42753 269550
rect 674367 266654 674433 266655
rect 674367 266590 674368 266654
rect 674432 266590 674433 266654
rect 674367 266589 674433 266590
rect 674175 266506 674241 266507
rect 674175 266442 674176 266506
rect 674240 266442 674241 266506
rect 674175 266441 674241 266442
rect 673983 260142 674049 260143
rect 673983 260078 673984 260142
rect 674048 260078 674049 260142
rect 673983 260077 674049 260078
rect 40575 251706 40641 251707
rect 40575 251642 40576 251706
rect 40640 251642 40641 251706
rect 40575 251641 40641 251642
rect 40578 236759 40638 251641
rect 42111 251410 42177 251411
rect 42111 251346 42112 251410
rect 42176 251346 42177 251410
rect 42111 251345 42177 251346
rect 41343 250226 41409 250227
rect 41343 250162 41344 250226
rect 41408 250162 41409 250226
rect 41343 250161 41409 250162
rect 40767 248746 40833 248747
rect 40767 248682 40768 248746
rect 40832 248682 40833 248746
rect 40767 248681 40833 248682
rect 40575 236758 40641 236759
rect 40575 236694 40576 236758
rect 40640 236694 40641 236758
rect 40575 236693 40641 236694
rect 40770 226843 40830 248681
rect 41151 248154 41217 248155
rect 41151 248090 41152 248154
rect 41216 248090 41217 248154
rect 41151 248089 41217 248090
rect 40959 247710 41025 247711
rect 40959 247646 40960 247710
rect 41024 247646 41025 247710
rect 40959 247645 41025 247646
rect 40962 230395 41022 247645
rect 40959 230394 41025 230395
rect 40959 230330 40960 230394
rect 41024 230330 41025 230394
rect 40959 230329 41025 230330
rect 41154 230099 41214 248089
rect 41151 230098 41217 230099
rect 41151 230034 41152 230098
rect 41216 230034 41217 230098
rect 41151 230033 41217 230034
rect 41346 229359 41406 250161
rect 41919 247562 41985 247563
rect 41919 247498 41920 247562
rect 41984 247498 41985 247562
rect 41919 247497 41985 247498
rect 41535 246230 41601 246231
rect 41535 246166 41536 246230
rect 41600 246166 41601 246230
rect 41535 246165 41601 246166
rect 41538 231283 41598 246165
rect 41727 245490 41793 245491
rect 41727 245426 41728 245490
rect 41792 245426 41793 245490
rect 41727 245425 41793 245426
rect 41730 235575 41790 245425
rect 41922 236907 41982 247497
rect 42114 238683 42174 251345
rect 42687 250966 42753 250967
rect 42687 250902 42688 250966
rect 42752 250902 42753 250966
rect 42687 250901 42753 250902
rect 42495 246970 42561 246971
rect 42495 246906 42496 246970
rect 42560 246906 42561 246970
rect 42495 246905 42561 246906
rect 42303 246082 42369 246083
rect 42303 246018 42304 246082
rect 42368 246018 42369 246082
rect 42303 246017 42369 246018
rect 42111 238682 42177 238683
rect 42111 238618 42112 238682
rect 42176 238618 42177 238682
rect 42111 238617 42177 238618
rect 42111 238534 42177 238535
rect 42111 238470 42112 238534
rect 42176 238470 42177 238534
rect 42111 238469 42177 238470
rect 41919 236906 41985 236907
rect 41919 236842 41920 236906
rect 41984 236842 41985 236906
rect 41919 236841 41985 236842
rect 41919 236758 41985 236759
rect 41919 236694 41920 236758
rect 41984 236694 41985 236758
rect 41919 236693 41985 236694
rect 41727 235574 41793 235575
rect 41727 235510 41728 235574
rect 41792 235510 41793 235574
rect 41727 235509 41793 235510
rect 41535 231282 41601 231283
rect 41535 231218 41536 231282
rect 41600 231218 41601 231282
rect 41535 231217 41601 231218
rect 41343 229358 41409 229359
rect 41343 229294 41344 229358
rect 41408 229294 41409 229358
rect 41343 229293 41409 229294
rect 41922 227435 41982 236693
rect 41919 227434 41985 227435
rect 41919 227370 41920 227434
rect 41984 227370 41985 227434
rect 41919 227369 41985 227370
rect 40767 226842 40833 226843
rect 40767 226778 40768 226842
rect 40832 226778 40833 226842
rect 40767 226777 40833 226778
rect 42114 226399 42174 238469
rect 42306 234391 42366 246017
rect 42498 234835 42558 246905
rect 42690 238535 42750 250901
rect 42879 249930 42945 249931
rect 42879 249866 42880 249930
rect 42944 249866 42945 249930
rect 42879 249865 42945 249866
rect 42687 238534 42753 238535
rect 42687 238470 42688 238534
rect 42752 238470 42753 238534
rect 42687 238469 42753 238470
rect 42495 234834 42561 234835
rect 42495 234770 42496 234834
rect 42560 234770 42561 234834
rect 42495 234769 42561 234770
rect 42303 234390 42369 234391
rect 42303 234326 42304 234390
rect 42368 234326 42369 234390
rect 42303 234325 42369 234326
rect 42882 233651 42942 249865
rect 397119 237054 397185 237055
rect 397119 236990 397120 237054
rect 397184 236990 397185 237054
rect 397119 236989 397185 236990
rect 397503 237054 397569 237055
rect 397503 236990 397504 237054
rect 397568 236990 397569 237054
rect 397503 236989 397569 236990
rect 397122 236315 397182 236989
rect 397506 236793 397566 236989
rect 397506 236759 397758 236793
rect 407298 236759 407742 236793
rect 397506 236758 397761 236759
rect 397506 236733 397696 236758
rect 397695 236694 397696 236733
rect 397760 236694 397761 236758
rect 397695 236693 397761 236694
rect 407295 236758 407742 236759
rect 407295 236694 407296 236758
rect 407360 236733 407742 236758
rect 407360 236694 407361 236733
rect 407295 236693 407361 236694
rect 407682 236315 407742 236733
rect 397119 236314 397185 236315
rect 397119 236250 397120 236314
rect 397184 236250 397185 236314
rect 397119 236249 397185 236250
rect 407679 236314 407745 236315
rect 407679 236250 407680 236314
rect 407744 236250 407745 236314
rect 407679 236249 407745 236250
rect 413631 236166 413697 236167
rect 413631 236102 413632 236166
rect 413696 236127 413697 236166
rect 414015 236166 414081 236167
rect 414015 236127 414016 236166
rect 413696 236102 414016 236127
rect 414080 236102 414081 236166
rect 413631 236101 414081 236102
rect 413634 236067 414078 236101
rect 42879 233650 42945 233651
rect 42879 233586 42880 233650
rect 42944 233586 42945 233650
rect 42879 233585 42945 233586
rect 42111 226398 42177 226399
rect 42111 226334 42112 226398
rect 42176 226334 42177 226398
rect 42111 226333 42177 226334
rect 673986 217519 674046 260077
rect 674178 218407 674238 266441
rect 674175 218406 674241 218407
rect 674175 218342 674176 218406
rect 674240 218342 674241 218406
rect 674175 218341 674241 218342
rect 674175 218110 674241 218111
rect 674175 218046 674176 218110
rect 674240 218046 674241 218110
rect 674175 218045 674241 218046
rect 673983 217518 674049 217519
rect 673983 217454 673984 217518
rect 674048 217454 674049 217518
rect 673983 217453 674049 217454
rect 673983 217370 674049 217371
rect 673983 217306 673984 217370
rect 674048 217306 674049 217370
rect 673983 217305 674049 217306
rect 673986 216039 674046 217305
rect 673983 216038 674049 216039
rect 673983 215974 673984 216038
rect 674048 215974 674049 216038
rect 673983 215973 674049 215974
rect 42111 208786 42177 208787
rect 42111 208722 42112 208786
rect 42176 208722 42177 208786
rect 42111 208721 42177 208722
rect 41535 207898 41601 207899
rect 41535 207834 41536 207898
rect 41600 207834 41601 207898
rect 41535 207833 41601 207834
rect 40959 207010 41025 207011
rect 40959 206946 40960 207010
rect 41024 206946 41025 207010
rect 40959 206945 41025 206946
rect 40575 206418 40641 206419
rect 40575 206354 40576 206418
rect 40640 206354 40641 206418
rect 40575 206353 40641 206354
rect 40383 204050 40449 204051
rect 40383 203986 40384 204050
rect 40448 203986 40449 204050
rect 40383 203985 40449 203986
rect 40386 193691 40446 203985
rect 40383 193690 40449 193691
rect 40383 193626 40384 193690
rect 40448 193626 40449 193690
rect 40383 193625 40449 193626
rect 40578 190435 40638 206353
rect 40767 205530 40833 205531
rect 40767 205466 40768 205530
rect 40832 205466 40833 205530
rect 40767 205465 40833 205466
rect 40575 190434 40641 190435
rect 40575 190370 40576 190434
rect 40640 190370 40641 190434
rect 40575 190369 40641 190370
rect 40770 183627 40830 205465
rect 40962 185995 41022 206945
rect 41343 204938 41409 204939
rect 41343 204874 41344 204938
rect 41408 204874 41409 204938
rect 41343 204873 41409 204874
rect 41151 204494 41217 204495
rect 41151 204430 41152 204494
rect 41216 204430 41217 204494
rect 41151 204429 41217 204430
rect 41154 187179 41214 204429
rect 41151 187178 41217 187179
rect 41151 187114 41152 187178
rect 41216 187114 41217 187178
rect 41151 187113 41217 187114
rect 41346 186883 41406 204873
rect 41538 195467 41598 207833
rect 41919 207750 41985 207751
rect 41919 207686 41920 207750
rect 41984 207686 41985 207750
rect 41919 207685 41985 207686
rect 41727 202866 41793 202867
rect 41727 202802 41728 202866
rect 41792 202802 41793 202866
rect 41727 202801 41793 202802
rect 41535 195466 41601 195467
rect 41535 195402 41536 195466
rect 41600 195402 41601 195466
rect 41535 195401 41601 195402
rect 41730 191175 41790 202801
rect 41727 191174 41793 191175
rect 41727 191110 41728 191174
rect 41792 191110 41793 191174
rect 41727 191109 41793 191110
rect 41343 186882 41409 186883
rect 41343 186818 41344 186882
rect 41408 186818 41409 186882
rect 41343 186817 41409 186818
rect 40959 185994 41025 185995
rect 40959 185930 40960 185994
rect 41024 185930 41025 185994
rect 40959 185929 41025 185930
rect 40767 183626 40833 183627
rect 40767 183562 40768 183626
rect 40832 183562 40833 183626
rect 40767 183561 40833 183562
rect 41922 183183 41982 207685
rect 42114 184219 42174 208721
rect 42495 203754 42561 203755
rect 42495 203690 42496 203754
rect 42560 203690 42561 203754
rect 42495 203689 42561 203690
rect 42303 202274 42369 202275
rect 42303 202210 42304 202274
rect 42368 202210 42369 202274
rect 42303 202209 42369 202210
rect 42306 192359 42366 202209
rect 42303 192358 42369 192359
rect 42303 192294 42304 192358
rect 42368 192294 42369 192358
rect 42303 192293 42369 192294
rect 42498 191767 42558 203689
rect 42687 203014 42753 203015
rect 42687 202950 42688 203014
rect 42752 202950 42753 203014
rect 42687 202949 42753 202950
rect 42495 191766 42561 191767
rect 42495 191702 42496 191766
rect 42560 191702 42561 191766
rect 42495 191701 42561 191702
rect 42690 188067 42750 202949
rect 673986 197499 674046 215973
rect 674178 197687 674238 218045
rect 674370 217075 674430 266589
rect 676287 266358 676353 266359
rect 676287 266294 676288 266358
rect 676352 266294 676353 266358
rect 676287 266293 676353 266294
rect 674559 261030 674625 261031
rect 674559 260966 674560 261030
rect 674624 260966 674625 261030
rect 674559 260965 674625 260966
rect 674562 218555 674622 260965
rect 676290 260291 676350 266293
rect 676287 260290 676353 260291
rect 676287 260226 676288 260290
rect 676352 260226 676353 260290
rect 676287 260225 676353 260226
rect 674943 258070 675009 258071
rect 674943 258006 674944 258070
rect 675008 258006 675009 258070
rect 674943 258005 675009 258006
rect 674751 249338 674817 249339
rect 674751 249274 674752 249338
rect 674816 249274 674817 249338
rect 674751 249273 674817 249274
rect 674559 218554 674625 218555
rect 674559 218490 674560 218554
rect 674624 218490 674625 218554
rect 674559 218489 674625 218490
rect 674559 218406 674625 218407
rect 674559 218342 674560 218406
rect 674624 218342 674625 218406
rect 674559 218341 674625 218342
rect 674562 217371 674622 218341
rect 674559 217370 674625 217371
rect 674559 217306 674560 217370
rect 674624 217306 674625 217370
rect 674559 217305 674625 217306
rect 674367 217074 674433 217075
rect 674367 217010 674368 217074
rect 674432 217010 674433 217074
rect 674367 217009 674433 217010
rect 674175 197686 674241 197687
rect 674175 197622 674176 197686
rect 674240 197622 674241 197686
rect 674175 197621 674241 197622
rect 673986 197439 674238 197499
rect 673983 197242 674049 197243
rect 673983 197178 673984 197242
rect 674048 197178 674049 197242
rect 673983 197177 674049 197178
rect 42687 188066 42753 188067
rect 42687 188002 42688 188066
rect 42752 188002 42753 188066
rect 42687 188001 42753 188002
rect 42111 184218 42177 184219
rect 42111 184154 42112 184218
rect 42176 184154 42177 184218
rect 42111 184153 42177 184154
rect 41919 183182 41985 183183
rect 41919 183118 41920 183182
rect 41984 183118 41985 183182
rect 41919 183117 41985 183118
rect 673986 172823 674046 197177
rect 673983 172822 674049 172823
rect 673983 172758 673984 172822
rect 674048 172758 674049 172822
rect 673983 172757 674049 172758
rect 673983 172082 674049 172083
rect 673983 172018 673984 172082
rect 674048 172018 674049 172082
rect 673983 172017 674049 172018
rect 673986 128423 674046 172017
rect 674178 170603 674238 197439
rect 674370 171491 674430 217009
rect 674754 216927 674814 249273
rect 674946 234539 675006 258005
rect 675711 257108 675777 257109
rect 675711 257044 675712 257108
rect 675776 257044 675777 257108
rect 675711 257043 675777 257044
rect 675135 256590 675201 256591
rect 675135 256526 675136 256590
rect 675200 256526 675201 256590
rect 675135 256525 675201 256526
rect 675138 239127 675198 256525
rect 675714 243715 675774 257043
rect 675903 253630 675969 253631
rect 675903 253566 675904 253630
rect 675968 253566 675969 253630
rect 675903 253565 675969 253566
rect 675711 243714 675777 243715
rect 675711 243650 675712 243714
rect 675776 243650 675777 243714
rect 675711 243649 675777 243650
rect 675135 239126 675201 239127
rect 675135 239062 675136 239126
rect 675200 239062 675201 239126
rect 675135 239061 675201 239062
rect 675906 238091 675966 253565
rect 676671 248006 676737 248007
rect 676671 247942 676672 248006
rect 676736 247942 676737 248006
rect 676671 247941 676737 247942
rect 676479 247858 676545 247859
rect 676479 247794 676480 247858
rect 676544 247794 676545 247858
rect 676479 247793 676545 247794
rect 675903 238090 675969 238091
rect 675903 238026 675904 238090
rect 675968 238026 675969 238090
rect 675903 238025 675969 238026
rect 676482 236019 676542 247793
rect 676479 236018 676545 236019
rect 676479 235954 676480 236018
rect 676544 235954 676545 236018
rect 676479 235953 676545 235954
rect 674943 234538 675009 234539
rect 674943 234474 674944 234538
rect 675008 234474 675009 234538
rect 674943 234473 675009 234474
rect 676674 232615 676734 247941
rect 676671 232614 676737 232615
rect 676671 232550 676672 232614
rect 676736 232550 676737 232614
rect 676671 232549 676737 232550
rect 674751 216926 674817 216927
rect 674751 216862 674752 216926
rect 674816 216862 674817 216926
rect 674751 216861 674817 216862
rect 674559 214706 674625 214707
rect 674559 214642 674560 214706
rect 674624 214642 674625 214706
rect 674559 214641 674625 214642
rect 674562 189991 674622 214641
rect 674751 213522 674817 213523
rect 674751 213458 674752 213522
rect 674816 213458 674817 213522
rect 674751 213457 674817 213458
rect 674754 195171 674814 213457
rect 675135 210562 675201 210563
rect 675135 210498 675136 210562
rect 675200 210498 675201 210562
rect 675135 210497 675201 210498
rect 674943 209082 675009 209083
rect 674943 209018 674944 209082
rect 675008 209018 675009 209082
rect 674943 209017 675009 209018
rect 674751 195170 674817 195171
rect 674751 195106 674752 195170
rect 674816 195106 674817 195170
rect 674751 195105 674817 195106
rect 674946 193099 675006 209017
rect 675138 193987 675198 210497
rect 675711 204790 675777 204791
rect 675711 204726 675712 204790
rect 675776 204726 675777 204790
rect 675711 204725 675777 204726
rect 675135 193986 675201 193987
rect 675135 193922 675136 193986
rect 675200 193922 675201 193986
rect 675135 193921 675201 193922
rect 674943 193098 675009 193099
rect 674943 193034 674944 193098
rect 675008 193034 675009 193098
rect 674943 193033 675009 193034
rect 674559 189990 674625 189991
rect 674559 189926 674560 189990
rect 674624 189926 674625 189990
rect 674559 189925 674625 189926
rect 675714 188511 675774 204725
rect 675903 204642 675969 204643
rect 675903 204578 675904 204642
rect 675968 204578 675969 204642
rect 675903 204577 675969 204578
rect 675906 192211 675966 204577
rect 675903 192210 675969 192211
rect 675903 192146 675904 192210
rect 675968 192146 675969 192210
rect 675903 192145 675969 192146
rect 675711 188510 675777 188511
rect 675711 188446 675712 188510
rect 675776 188446 675777 188510
rect 675711 188445 675777 188446
rect 674367 171490 674433 171491
rect 674367 171426 674368 171490
rect 674432 171426 674433 171490
rect 674367 171425 674433 171426
rect 674367 171046 674433 171047
rect 674367 170982 674368 171046
rect 674432 170982 674433 171046
rect 674367 170981 674433 170982
rect 674175 170602 674241 170603
rect 674175 170538 674176 170602
rect 674240 170538 674241 170602
rect 674175 170537 674241 170538
rect 674370 170193 674430 170981
rect 674178 170133 674430 170193
rect 673983 128422 674049 128423
rect 673983 128358 673984 128422
rect 674048 128358 674049 128422
rect 673983 128357 674049 128358
rect 674178 127387 674238 170133
rect 676287 169270 676353 169271
rect 676287 169206 676288 169270
rect 676352 169206 676353 169270
rect 676287 169205 676353 169206
rect 676095 168678 676161 168679
rect 676095 168614 676096 168678
rect 676160 168614 676161 168678
rect 676095 168613 676161 168614
rect 675519 168086 675585 168087
rect 675519 168022 675520 168086
rect 675584 168022 675585 168086
rect 675519 168021 675585 168022
rect 674559 167346 674625 167347
rect 674559 167282 674560 167346
rect 674624 167282 674625 167346
rect 674559 167281 674625 167282
rect 674367 167050 674433 167051
rect 674367 166986 674368 167050
rect 674432 166986 674433 167050
rect 674367 166985 674433 166986
rect 674370 143963 674430 166985
rect 674562 150919 674622 167281
rect 675327 165718 675393 165719
rect 675327 165654 675328 165718
rect 675392 165654 675393 165718
rect 675327 165653 675393 165654
rect 674943 165126 675009 165127
rect 674943 165062 674944 165126
rect 675008 165062 675009 165126
rect 674943 165061 675009 165062
rect 674751 164534 674817 164535
rect 674751 164470 674752 164534
rect 674816 164470 674817 164534
rect 674751 164469 674817 164470
rect 674559 150918 674625 150919
rect 674559 150854 674560 150918
rect 674624 150854 674625 150918
rect 674559 150853 674625 150854
rect 674754 149587 674814 164469
rect 674751 149586 674817 149587
rect 674751 149522 674752 149586
rect 674816 149522 674817 149586
rect 674751 149521 674817 149522
rect 674946 147959 675006 165061
rect 675135 163646 675201 163647
rect 675135 163582 675136 163646
rect 675200 163582 675201 163646
rect 675135 163581 675201 163582
rect 675138 150327 675198 163581
rect 675330 154471 675390 165653
rect 675522 155211 675582 168021
rect 675711 166606 675777 166607
rect 675711 166542 675712 166606
rect 675776 166542 675777 166606
rect 675711 166541 675777 166542
rect 675714 157727 675774 166541
rect 675903 165570 675969 165571
rect 675903 165506 675904 165570
rect 675968 165506 675969 165570
rect 675903 165505 675969 165506
rect 675711 157726 675777 157727
rect 675711 157662 675712 157726
rect 675776 157662 675777 157726
rect 675711 157661 675777 157662
rect 675519 155210 675585 155211
rect 675519 155146 675520 155210
rect 675584 155146 675585 155210
rect 675519 155145 675585 155146
rect 675327 154470 675393 154471
rect 675327 154406 675328 154470
rect 675392 154406 675393 154470
rect 675327 154405 675393 154406
rect 675906 153879 675966 165505
rect 676098 158171 676158 168613
rect 676095 158170 676161 158171
rect 676095 158106 676096 158170
rect 676160 158106 676161 158170
rect 676095 158105 676161 158106
rect 676290 156987 676350 169205
rect 676863 162758 676929 162759
rect 676863 162694 676864 162758
rect 676928 162694 676929 162758
rect 676863 162693 676929 162694
rect 676287 156986 676353 156987
rect 676287 156922 676288 156986
rect 676352 156922 676353 156986
rect 676287 156921 676353 156922
rect 675903 153878 675969 153879
rect 675903 153814 675904 153878
rect 675968 153814 675969 153878
rect 675903 153813 675969 153814
rect 676866 152695 676926 162693
rect 676863 152694 676929 152695
rect 676863 152630 676864 152694
rect 676928 152630 676929 152694
rect 676863 152629 676929 152630
rect 675135 150326 675201 150327
rect 675135 150262 675136 150326
rect 675200 150262 675201 150326
rect 675135 150261 675201 150262
rect 674943 147958 675009 147959
rect 674943 147894 674944 147958
rect 675008 147894 675009 147958
rect 674943 147893 675009 147894
rect 674367 143962 674433 143963
rect 674367 143898 674368 143962
rect 674432 143898 674433 143962
rect 674367 143897 674433 143898
rect 674175 127386 674241 127387
rect 674175 127322 674176 127386
rect 674240 127322 674241 127386
rect 674175 127321 674241 127322
rect 675519 125462 675585 125463
rect 675519 125398 675520 125462
rect 675584 125398 675585 125462
rect 675519 125397 675585 125398
rect 674175 123390 674241 123391
rect 674175 123326 674176 123390
rect 674240 123326 674241 123390
rect 674175 123325 674241 123326
rect 674178 106519 674238 123325
rect 675522 112143 675582 125397
rect 675903 123908 675969 123909
rect 675903 123844 675904 123908
rect 675968 123844 675969 123908
rect 675903 123843 675969 123844
rect 675711 120874 675777 120875
rect 675711 120810 675712 120874
rect 675776 120810 675777 120874
rect 675711 120809 675777 120810
rect 675519 112142 675585 112143
rect 675519 112078 675520 112142
rect 675584 112078 675585 112142
rect 675519 112077 675585 112078
rect 674175 106518 674241 106519
rect 674175 106454 674176 106518
rect 674240 106454 674241 106518
rect 674175 106453 674241 106454
rect 675714 103559 675774 120809
rect 675906 110959 675966 123843
rect 676479 115694 676545 115695
rect 676479 115630 676480 115694
rect 676544 115630 676545 115694
rect 676479 115629 676545 115630
rect 675903 110958 675969 110959
rect 675903 110894 675904 110958
rect 675968 110894 675969 110958
rect 675903 110893 675969 110894
rect 675711 103558 675777 103559
rect 675711 103494 675712 103558
rect 675776 103494 675777 103558
rect 675711 103493 675777 103494
rect 676482 101635 676542 115629
rect 676671 115250 676737 115251
rect 676671 115186 676672 115250
rect 676736 115186 676737 115250
rect 676671 115185 676737 115186
rect 676479 101634 676545 101635
rect 676479 101570 676480 101634
rect 676544 101570 676545 101634
rect 676479 101569 676545 101570
rect 676674 99859 676734 115185
rect 676671 99858 676737 99859
rect 676671 99794 676672 99858
rect 676736 99794 676737 99858
rect 676671 99793 676737 99794
rect 417471 40510 417537 40511
rect 417471 40446 417472 40510
rect 417536 40446 417537 40510
rect 417471 40445 417537 40446
rect 417663 40510 417729 40511
rect 417663 40446 417664 40510
rect 417728 40446 417729 40510
rect 417663 40445 417729 40446
rect 417474 40323 417534 40445
rect 417666 40323 417726 40445
rect 417474 40263 417726 40323
<< metal5 >>
rect 76810 1018624 88978 1030788
rect 124810 1018624 136978 1030788
rect 172810 1018624 184978 1030788
rect 231210 1018624 243378 1030788
rect 282610 1018624 294778 1030788
rect 341210 1018624 353378 1030788
rect 427610 1018624 439778 1030788
rect 477410 1018624 489578 1030788
rect 527210 1018624 539378 1030788
rect 577010 1018624 589178 1030788
rect 628410 1018624 640578 1030788
rect 6811 956610 18975 968778
rect 698624 945422 710788 957590
rect 6167 915054 19619 925934
rect 697980 893466 711432 904346
rect 6811 872210 18975 884378
rect 698512 848240 711002 860780
rect 6811 829810 18975 841978
rect 698624 805222 710788 817390
rect 6598 787420 19088 799960
rect 698512 760840 711002 773380
rect 6598 744220 19088 756760
rect 698512 716440 711002 728980
rect 6598 701020 19088 713560
rect 698512 672240 711002 684780
rect 6598 657620 19088 670160
rect 698512 628040 711002 640580
rect 6598 614420 19088 626960
rect 6598 571220 19088 583760
rect 698512 583640 711002 596180
rect 6598 528020 19088 540560
rect 698512 539440 711002 551980
rect 6811 484810 18975 496978
rect 698624 496422 710788 508590
rect 6167 443254 19619 454134
rect 697980 453666 711432 464546
rect 6598 400220 19088 412760
rect 698624 409822 710788 421990
rect 6598 357020 19088 369560
rect 698512 365240 711002 377780
rect 6598 313620 19088 326160
rect 698512 321040 711002 333580
rect 6598 270420 19088 282960
rect 698512 276840 711002 289380
rect 6598 227220 19088 239760
rect 698512 232440 711002 244980
rect 6598 184020 19088 196560
rect 698512 188240 711002 200780
rect 698512 144040 711002 156580
rect 6811 111610 18975 123778
rect 698512 99640 711002 112180
rect 6167 70054 19619 80934
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200180 19088
rect 243266 6167 254146 19619
rect 296240 6598 308780 19088
rect 351040 6598 363580 19088
rect 405840 6598 418380 19088
rect 460640 6598 473180 19088
rect 515440 6598 527980 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use user_id_programming  user_id_value
timestamp 1625003591
transform 1 0 656624 0 1 80926
box 0 0 7109 7077
use storage  storage
timestamp 1625003591
transform 1 0 52032 0 1 53156
box 1066 70 92000 191480
use mgmt_core  soc
timestamp 1625003591
transform 1 0 190434 0 1 53602
box 0 0 450000 168026
use sky130_fd_sc_hvl__lsbufhv2lv_1_wrapped  rstb_level
timestamp 1625003591
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use simple_por  por
timestamp 1625003591
transform 1 0 654146 0 -1 112882
box 25 11 11344 8291
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1625003591
transform -1 0 710203 0 1 160400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1625003591
transform -1 0 710203 0 1 116200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1625003591
transform 1 0 7631 0 1 242800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1625003591
transform 1 0 7631 0 1 199600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1625003591
transform 1 0 7631 0 1 286000
box -1620 -364 34000 13964
use mgmt_protect  mgmt_buffers
timestamp 1625003591
transform 1 0 192180 0 1 240036
box -2762 -2778 222734 26170
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1625003591
transform -1 0 710203 0 1 206400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1625003591
transform -1 0 710203 0 1 249400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1625003591
transform 1 0 7631 0 1 372400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1625003591
transform 1 0 7631 0 1 329200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1625003591
transform -1 0 710203 0 1 292400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1625003591
transform -1 0 710203 0 1 338400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1625003591
transform -1 0 710203 0 1 383000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1625003591
transform 1 0 7631 0 1 415600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1625003591
transform 1 0 7631 0 1 462400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1625003591
transform -1 0 710203 0 1 511800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1625003591
transform -1 0 710203 0 1 469000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1625003591
transform 1 0 7631 0 1 588224
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1625003591
transform 1 0 7631 0 1 631400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1625003591
transform 1 0 7631 0 1 674600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1625003591
transform -1 0 710203 0 1 645400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1625003591
transform -1 0 710203 0 1 601000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1625003591
transform -1 0 710203 0 1 555800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1625003591
transform -1 0 710203 0 1 689600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1625003591
transform 1 0 7631 0 1 717800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1625003591
transform 1 0 7631 0 1 761000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1625003591
transform 1 0 7631 0 1 804200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in_1\[11\]
timestamp 1625003591
transform -1 0 710203 0 1 866800
box -1620 -364 34000 13964
use user_analog_project_wrapper  mprj
timestamp 1625003591
transform 1 0 65308 0 1 278718
box -800 -800 584800 704000
use chip_io_alt  padframe
timestamp 1625003591
transform 1 0 0 0 1 0
box 0 0 717600 1037600
<< labels >>
rlabel metal5 s 187640 6598 200180 19088 6 clock
port 0 nsew signal input
rlabel metal5 s 351040 6598 363580 19088 6 flash_clk
port 1 nsew signal tristate
rlabel metal5 s 296240 6598 308780 19088 6 flash_csb
port 2 nsew signal tristate
rlabel metal5 s 405840 6598 418380 19088 6 flash_io0
port 3 nsew signal tristate
rlabel metal5 s 460640 6598 473180 19088 6 flash_io1
port 4 nsew signal tristate
rlabel metal5 s 515440 6598 527980 19088 6 gpio
port 5 nsew signal bidirectional
rlabel metal5 s 698512 99640 711002 112180 6 mprj_io[0]
port 6 nsew signal bidirectional
rlabel metal5 s 698512 672240 711002 684780 6 mprj_io[10]
port 7 nsew signal bidirectional
rlabel metal5 s 698512 716440 711002 728980 6 mprj_io[11]
port 8 nsew signal bidirectional
rlabel metal5 s 698512 760840 711002 773380 6 mprj_io[12]
port 9 nsew signal bidirectional
rlabel metal5 s 698512 848240 711002 860780 6 mprj_io[13]
port 10 nsew signal bidirectional
rlabel metal5 s 698624 945422 710788 957590 6 mprj_io[14]
port 11 nsew signal bidirectional
rlabel metal5 s 628410 1018624 640578 1030788 6 mprj_io[15]
port 12 nsew signal bidirectional
rlabel metal5 s 527210 1018624 539378 1030788 6 mprj_io[16]
port 13 nsew signal bidirectional
rlabel metal5 s 477410 1018624 489578 1030788 6 mprj_io[17]
port 14 nsew signal bidirectional
rlabel metal5 s 427610 1018624 439778 1030788 6 mprj_io[18]
port 15 nsew signal bidirectional
rlabel metal5 s 282610 1018624 294778 1030788 6 mprj_io[19]
port 16 nsew signal bidirectional
rlabel metal5 s 698512 144040 711002 156580 6 mprj_io[1]
port 17 nsew signal bidirectional
rlabel metal5 s 231210 1018624 243378 1030788 6 mprj_io[20]
port 18 nsew signal bidirectional
rlabel metal5 s 172810 1018624 184978 1030788 6 mprj_io[21]
port 19 nsew signal bidirectional
rlabel metal5 s 124810 1018624 136978 1030788 6 mprj_io[22]
port 20 nsew signal bidirectional
rlabel metal5 s 76810 1018624 88978 1030788 6 mprj_io[23]
port 21 nsew signal bidirectional
rlabel metal5 s 6811 956610 18975 968778 6 mprj_io[24]
port 22 nsew signal bidirectional
rlabel metal5 s 6598 787420 19088 799960 6 mprj_io[25]
port 23 nsew signal bidirectional
rlabel metal5 s 6598 744220 19088 756760 6 mprj_io[26]
port 24 nsew signal bidirectional
rlabel metal5 s 6598 701020 19088 713560 6 mprj_io[27]
port 25 nsew signal bidirectional
rlabel metal5 s 6598 657620 19088 670160 6 mprj_io[28]
port 26 nsew signal bidirectional
rlabel metal5 s 6598 614420 19088 626960 6 mprj_io[29]
port 27 nsew signal bidirectional
rlabel metal5 s 698512 188240 711002 200780 6 mprj_io[2]
port 28 nsew signal bidirectional
rlabel metal5 s 6598 571220 19088 583760 6 mprj_io[30]
port 29 nsew signal bidirectional
rlabel metal5 s 6598 528020 19088 540560 6 mprj_io[31]
port 30 nsew signal bidirectional
rlabel metal5 s 6598 400220 19088 412760 6 mprj_io[32]
port 31 nsew signal bidirectional
rlabel metal5 s 6598 357020 19088 369560 6 mprj_io[33]
port 32 nsew signal bidirectional
rlabel metal5 s 6598 313620 19088 326160 6 mprj_io[34]
port 33 nsew signal bidirectional
rlabel metal5 s 6598 270420 19088 282960 6 mprj_io[35]
port 34 nsew signal bidirectional
rlabel metal5 s 6598 227220 19088 239760 6 mprj_io[36]
port 35 nsew signal bidirectional
rlabel metal5 s 6598 184020 19088 196560 6 mprj_io[37]
port 36 nsew signal bidirectional
rlabel metal5 s 698512 232440 711002 244980 6 mprj_io[3]
port 37 nsew signal bidirectional
rlabel metal5 s 698512 276840 711002 289380 6 mprj_io[4]
port 38 nsew signal bidirectional
rlabel metal5 s 698512 321040 711002 333580 6 mprj_io[5]
port 39 nsew signal bidirectional
rlabel metal5 s 698512 365240 711002 377780 6 mprj_io[6]
port 40 nsew signal bidirectional
rlabel metal5 s 698512 539440 711002 551980 6 mprj_io[7]
port 41 nsew signal bidirectional
rlabel metal5 s 698512 583640 711002 596180 6 mprj_io[8]
port 42 nsew signal bidirectional
rlabel metal5 s 698512 628040 711002 640580 6 mprj_io[9]
port 43 nsew signal bidirectional
rlabel metal5 s 136713 7143 144149 18309 6 resetb
port 44 nsew signal input
rlabel metal5 s 697980 893466 711432 904346 6 vccd1
port 45 nsew signal bidirectional
rlabel metal5 s 6167 915054 19619 925934 6 vccd2
port 46 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18975 6 vdda
port 47 nsew signal bidirectional
rlabel metal5 s 698624 805222 710788 817390 6 vdda1
port 48 nsew signal bidirectional
rlabel metal5 s 698624 496422 710788 508590 6 vdda1_2
port 49 nsew signal bidirectional
rlabel metal5 s 6811 484810 18975 496978 6 vdda2
port 50 nsew signal bidirectional
rlabel metal5 s 6811 872210 18975 884378 6 vddio_2
port 51 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030788 6 vssa1
port 52 nsew signal bidirectional
rlabel metal5 s 698624 409822 710788 421990 6 vssa1_2
port 53 nsew signal bidirectional
rlabel metal5 s 6811 829810 18975 841978 6 vssa2
port 54 nsew signal bidirectional
rlabel metal5 s 697980 453666 711432 464546 6 vssd1
port 55 nsew signal bidirectional
rlabel metal5 s 6167 443254 19619 454134 6 vssd2
port 56 nsew signal bidirectional
rlabel metal5 s 341210 1018624 353378 1030788 6 vssio_2
port 57 nsew signal bidirectional
rlabel metal5 s 6811 111610 18975 123778 6 vddio
port 58 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18975 6 vssio
port 59 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18975 6 vssa
port 60 nsew signal bidirectional
rlabel metal5 s 6167 70054 19619 80934 6 vccd
port 61 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19619 6 vssd
port 62 nsew signal bidirectional
rlabel metal2 s 579796 53602 579852 54402 6 pwr_ctrl_out[0]
port 63 nsew signal tristate
rlabel metal2 s 597092 53602 597148 54402 6 pwr_ctrl_out[1]
port 64 nsew signal tristate
rlabel metal2 s 614388 53602 614444 54402 6 pwr_ctrl_out[2]
port 65 nsew signal tristate
rlabel metal2 s 631684 53602 631740 54402 6 pwr_ctrl_out[3]
port 66 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
