magic
tech sky130A
timestamp 1602626256
<< metalrdl >>
tri -3800 11800 0 12400 se
tri 0 11800 3800 12400 sw
tri -7300 10100 -3800 11800 se
rect -3800 10100 3800 11800
tri 3800 10100 7300 11800 sw
tri -10100 7300 -7300 10100 se
rect -7300 7300 7300 10100
tri 7300 7300 10100 10100 sw
tri -11800 3800 -10100 7300 se
rect -10100 3800 10100 7300
tri 10100 3800 11800 7300 sw
tri -12400 0 -11800 3800 se
tri -12400 -3800 -11800 0 ne
rect -11800 -3800 11800 3800
tri 11800 0 12500 3800 sw
tri 11800 -3800 12500 0 nw
tri -11800 -7300 -10100 -3800 ne
rect -10100 -7300 10100 -3800
tri 10100 -7300 11800 -3800 nw
tri -10100 -10100 -7300 -7300 ne
rect -7300 -10100 7300 -7300
tri 7300 -10100 10100 -7300 nw
tri -7300 -11800 -3800 -10100 ne
rect -3800 -11800 3800 -10100
tri 3800 -11800 7300 -10100 nw
tri -3800 -12400 0 -11800 ne
tri 0 -12400 3800 -11800 nw
<< end >>
