magic
tech sky130A
magscale 12 1
timestamp 1598786680
<< metal5 >>
rect 15 60 30 75
rect 0 45 45 60
rect 15 30 30 45
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
