magic
tech sky130A
magscale 1 2
timestamp 1606422650
<< error_p >>
rect -265 1217 -207 1223
rect -147 1217 -89 1223
rect -29 1217 29 1223
rect 89 1217 147 1223
rect 207 1217 265 1223
rect -265 1183 -253 1217
rect -147 1183 -135 1217
rect -29 1183 -17 1217
rect 89 1183 101 1217
rect 207 1183 219 1217
rect -265 1177 -207 1183
rect -147 1177 -89 1183
rect -29 1177 29 1183
rect 89 1177 147 1183
rect 207 1177 265 1183
rect -265 489 -207 495
rect -147 489 -89 495
rect -29 489 29 495
rect 89 489 147 495
rect 207 489 265 495
rect -265 455 -253 489
rect -147 455 -135 489
rect -29 455 -17 489
rect 89 455 101 489
rect 207 455 219 489
rect -265 449 -207 455
rect -147 449 -89 455
rect -29 449 29 455
rect 89 449 147 455
rect 207 449 265 455
rect -265 381 -207 387
rect -147 381 -89 387
rect -29 381 29 387
rect 89 381 147 387
rect 207 381 265 387
rect -265 347 -253 381
rect -147 347 -135 381
rect -29 347 -17 381
rect 89 347 101 381
rect 207 347 219 381
rect -265 341 -207 347
rect -147 341 -89 347
rect -29 341 29 347
rect 89 341 147 347
rect 207 341 265 347
rect -265 -347 -207 -341
rect -147 -347 -89 -341
rect -29 -347 29 -341
rect 89 -347 147 -341
rect 207 -347 265 -341
rect -265 -381 -253 -347
rect -147 -381 -135 -347
rect -29 -381 -17 -347
rect 89 -381 101 -347
rect 207 -381 219 -347
rect -265 -387 -207 -381
rect -147 -387 -89 -381
rect -29 -387 29 -381
rect 89 -387 147 -381
rect 207 -387 265 -381
rect -265 -455 -207 -449
rect -147 -455 -89 -449
rect -29 -455 29 -449
rect 89 -455 147 -449
rect 207 -455 265 -449
rect -265 -489 -253 -455
rect -147 -489 -135 -455
rect -29 -489 -17 -455
rect 89 -489 101 -455
rect 207 -489 219 -455
rect -265 -495 -207 -489
rect -147 -495 -89 -489
rect -29 -495 29 -489
rect 89 -495 147 -489
rect 207 -495 265 -489
rect -265 -1183 -207 -1177
rect -147 -1183 -89 -1177
rect -29 -1183 29 -1177
rect 89 -1183 147 -1177
rect 207 -1183 265 -1177
rect -265 -1217 -253 -1183
rect -147 -1217 -135 -1183
rect -29 -1217 -17 -1183
rect 89 -1217 101 -1183
rect 207 -1217 219 -1183
rect -265 -1223 -207 -1217
rect -147 -1223 -89 -1217
rect -29 -1223 29 -1217
rect 89 -1223 147 -1217
rect 207 -1223 265 -1217
<< nwell >>
rect -462 -1355 462 1355
<< pmos >>
rect -266 536 -206 1136
rect -148 536 -88 1136
rect -30 536 30 1136
rect 88 536 148 1136
rect 206 536 266 1136
rect -266 -300 -206 300
rect -148 -300 -88 300
rect -30 -300 30 300
rect 88 -300 148 300
rect 206 -300 266 300
rect -266 -1136 -206 -536
rect -148 -1136 -88 -536
rect -30 -1136 30 -536
rect 88 -1136 148 -536
rect 206 -1136 266 -536
<< pdiff >>
rect -324 1124 -266 1136
rect -324 548 -312 1124
rect -278 548 -266 1124
rect -324 536 -266 548
rect -206 1124 -148 1136
rect -206 548 -194 1124
rect -160 548 -148 1124
rect -206 536 -148 548
rect -88 1124 -30 1136
rect -88 548 -76 1124
rect -42 548 -30 1124
rect -88 536 -30 548
rect 30 1124 88 1136
rect 30 548 42 1124
rect 76 548 88 1124
rect 30 536 88 548
rect 148 1124 206 1136
rect 148 548 160 1124
rect 194 548 206 1124
rect 148 536 206 548
rect 266 1124 324 1136
rect 266 548 278 1124
rect 312 548 324 1124
rect 266 536 324 548
rect -324 288 -266 300
rect -324 -288 -312 288
rect -278 -288 -266 288
rect -324 -300 -266 -288
rect -206 288 -148 300
rect -206 -288 -194 288
rect -160 -288 -148 288
rect -206 -300 -148 -288
rect -88 288 -30 300
rect -88 -288 -76 288
rect -42 -288 -30 288
rect -88 -300 -30 -288
rect 30 288 88 300
rect 30 -288 42 288
rect 76 -288 88 288
rect 30 -300 88 -288
rect 148 288 206 300
rect 148 -288 160 288
rect 194 -288 206 288
rect 148 -300 206 -288
rect 266 288 324 300
rect 266 -288 278 288
rect 312 -288 324 288
rect 266 -300 324 -288
rect -324 -548 -266 -536
rect -324 -1124 -312 -548
rect -278 -1124 -266 -548
rect -324 -1136 -266 -1124
rect -206 -548 -148 -536
rect -206 -1124 -194 -548
rect -160 -1124 -148 -548
rect -206 -1136 -148 -1124
rect -88 -548 -30 -536
rect -88 -1124 -76 -548
rect -42 -1124 -30 -548
rect -88 -1136 -30 -1124
rect 30 -548 88 -536
rect 30 -1124 42 -548
rect 76 -1124 88 -548
rect 30 -1136 88 -1124
rect 148 -548 206 -536
rect 148 -1124 160 -548
rect 194 -1124 206 -548
rect 148 -1136 206 -1124
rect 266 -548 324 -536
rect 266 -1124 278 -548
rect 312 -1124 324 -548
rect 266 -1136 324 -1124
<< pdiffc >>
rect -312 548 -278 1124
rect -194 548 -160 1124
rect -76 548 -42 1124
rect 42 548 76 1124
rect 160 548 194 1124
rect 278 548 312 1124
rect -312 -288 -278 288
rect -194 -288 -160 288
rect -76 -288 -42 288
rect 42 -288 76 288
rect 160 -288 194 288
rect 278 -288 312 288
rect -312 -1124 -278 -548
rect -194 -1124 -160 -548
rect -76 -1124 -42 -548
rect 42 -1124 76 -548
rect 160 -1124 194 -548
rect 278 -1124 312 -548
<< nsubdiff >>
rect -426 1285 -330 1319
rect 330 1285 426 1319
rect -426 1223 -392 1285
rect 392 1223 426 1285
rect -426 -1285 -392 -1223
rect 392 -1285 426 -1223
rect -426 -1319 -330 -1285
rect 330 -1319 426 -1285
<< nsubdiffcont >>
rect -330 1285 330 1319
rect -426 -1223 -392 1223
rect 392 -1223 426 1223
rect -330 -1319 330 -1285
<< poly >>
rect -269 1217 -203 1233
rect -269 1183 -253 1217
rect -219 1183 -203 1217
rect -269 1167 -203 1183
rect -151 1217 -85 1233
rect -151 1183 -135 1217
rect -101 1183 -85 1217
rect -151 1167 -85 1183
rect -33 1217 33 1233
rect -33 1183 -17 1217
rect 17 1183 33 1217
rect -33 1167 33 1183
rect 85 1217 151 1233
rect 85 1183 101 1217
rect 135 1183 151 1217
rect 85 1167 151 1183
rect 203 1217 269 1233
rect 203 1183 219 1217
rect 253 1183 269 1217
rect 203 1167 269 1183
rect -266 1136 -206 1167
rect -148 1136 -88 1167
rect -30 1136 30 1167
rect 88 1136 148 1167
rect 206 1136 266 1167
rect -266 505 -206 536
rect -148 505 -88 536
rect -30 505 30 536
rect 88 505 148 536
rect 206 505 266 536
rect -269 489 -203 505
rect -269 455 -253 489
rect -219 455 -203 489
rect -269 439 -203 455
rect -151 489 -85 505
rect -151 455 -135 489
rect -101 455 -85 489
rect -151 439 -85 455
rect -33 489 33 505
rect -33 455 -17 489
rect 17 455 33 489
rect -33 439 33 455
rect 85 489 151 505
rect 85 455 101 489
rect 135 455 151 489
rect 85 439 151 455
rect 203 489 269 505
rect 203 455 219 489
rect 253 455 269 489
rect 203 439 269 455
rect -269 381 -203 397
rect -269 347 -253 381
rect -219 347 -203 381
rect -269 331 -203 347
rect -151 381 -85 397
rect -151 347 -135 381
rect -101 347 -85 381
rect -151 331 -85 347
rect -33 381 33 397
rect -33 347 -17 381
rect 17 347 33 381
rect -33 331 33 347
rect 85 381 151 397
rect 85 347 101 381
rect 135 347 151 381
rect 85 331 151 347
rect 203 381 269 397
rect 203 347 219 381
rect 253 347 269 381
rect 203 331 269 347
rect -266 300 -206 331
rect -148 300 -88 331
rect -30 300 30 331
rect 88 300 148 331
rect 206 300 266 331
rect -266 -331 -206 -300
rect -148 -331 -88 -300
rect -30 -331 30 -300
rect 88 -331 148 -300
rect 206 -331 266 -300
rect -269 -347 -203 -331
rect -269 -381 -253 -347
rect -219 -381 -203 -347
rect -269 -397 -203 -381
rect -151 -347 -85 -331
rect -151 -381 -135 -347
rect -101 -381 -85 -347
rect -151 -397 -85 -381
rect -33 -347 33 -331
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect -33 -397 33 -381
rect 85 -347 151 -331
rect 85 -381 101 -347
rect 135 -381 151 -347
rect 85 -397 151 -381
rect 203 -347 269 -331
rect 203 -381 219 -347
rect 253 -381 269 -347
rect 203 -397 269 -381
rect -269 -455 -203 -439
rect -269 -489 -253 -455
rect -219 -489 -203 -455
rect -269 -505 -203 -489
rect -151 -455 -85 -439
rect -151 -489 -135 -455
rect -101 -489 -85 -455
rect -151 -505 -85 -489
rect -33 -455 33 -439
rect -33 -489 -17 -455
rect 17 -489 33 -455
rect -33 -505 33 -489
rect 85 -455 151 -439
rect 85 -489 101 -455
rect 135 -489 151 -455
rect 85 -505 151 -489
rect 203 -455 269 -439
rect 203 -489 219 -455
rect 253 -489 269 -455
rect 203 -505 269 -489
rect -266 -536 -206 -505
rect -148 -536 -88 -505
rect -30 -536 30 -505
rect 88 -536 148 -505
rect 206 -536 266 -505
rect -266 -1167 -206 -1136
rect -148 -1167 -88 -1136
rect -30 -1167 30 -1136
rect 88 -1167 148 -1136
rect 206 -1167 266 -1136
rect -269 -1183 -203 -1167
rect -269 -1217 -253 -1183
rect -219 -1217 -203 -1183
rect -269 -1233 -203 -1217
rect -151 -1183 -85 -1167
rect -151 -1217 -135 -1183
rect -101 -1217 -85 -1183
rect -151 -1233 -85 -1217
rect -33 -1183 33 -1167
rect -33 -1217 -17 -1183
rect 17 -1217 33 -1183
rect -33 -1233 33 -1217
rect 85 -1183 151 -1167
rect 85 -1217 101 -1183
rect 135 -1217 151 -1183
rect 85 -1233 151 -1217
rect 203 -1183 269 -1167
rect 203 -1217 219 -1183
rect 253 -1217 269 -1183
rect 203 -1233 269 -1217
<< polycont >>
rect -253 1183 -219 1217
rect -135 1183 -101 1217
rect -17 1183 17 1217
rect 101 1183 135 1217
rect 219 1183 253 1217
rect -253 455 -219 489
rect -135 455 -101 489
rect -17 455 17 489
rect 101 455 135 489
rect 219 455 253 489
rect -253 347 -219 381
rect -135 347 -101 381
rect -17 347 17 381
rect 101 347 135 381
rect 219 347 253 381
rect -253 -381 -219 -347
rect -135 -381 -101 -347
rect -17 -381 17 -347
rect 101 -381 135 -347
rect 219 -381 253 -347
rect -253 -489 -219 -455
rect -135 -489 -101 -455
rect -17 -489 17 -455
rect 101 -489 135 -455
rect 219 -489 253 -455
rect -253 -1217 -219 -1183
rect -135 -1217 -101 -1183
rect -17 -1217 17 -1183
rect 101 -1217 135 -1183
rect 219 -1217 253 -1183
<< locali >>
rect -426 1285 -330 1319
rect 330 1285 426 1319
rect -426 1223 -392 1285
rect 392 1223 426 1285
rect -269 1183 -253 1217
rect -219 1183 -203 1217
rect -151 1183 -135 1217
rect -101 1183 -85 1217
rect -33 1183 -17 1217
rect 17 1183 33 1217
rect 85 1183 101 1217
rect 135 1183 151 1217
rect 203 1183 219 1217
rect 253 1183 269 1217
rect -312 1124 -278 1140
rect -312 532 -278 548
rect -194 1124 -160 1140
rect -194 532 -160 548
rect -76 1124 -42 1140
rect -76 532 -42 548
rect 42 1124 76 1140
rect 42 532 76 548
rect 160 1124 194 1140
rect 160 532 194 548
rect 278 1124 312 1140
rect 278 532 312 548
rect -269 455 -253 489
rect -219 455 -203 489
rect -151 455 -135 489
rect -101 455 -85 489
rect -33 455 -17 489
rect 17 455 33 489
rect 85 455 101 489
rect 135 455 151 489
rect 203 455 219 489
rect 253 455 269 489
rect -269 347 -253 381
rect -219 347 -203 381
rect -151 347 -135 381
rect -101 347 -85 381
rect -33 347 -17 381
rect 17 347 33 381
rect 85 347 101 381
rect 135 347 151 381
rect 203 347 219 381
rect 253 347 269 381
rect -312 288 -278 304
rect -312 -304 -278 -288
rect -194 288 -160 304
rect -194 -304 -160 -288
rect -76 288 -42 304
rect -76 -304 -42 -288
rect 42 288 76 304
rect 42 -304 76 -288
rect 160 288 194 304
rect 160 -304 194 -288
rect 278 288 312 304
rect 278 -304 312 -288
rect -269 -381 -253 -347
rect -219 -381 -203 -347
rect -151 -381 -135 -347
rect -101 -381 -85 -347
rect -33 -381 -17 -347
rect 17 -381 33 -347
rect 85 -381 101 -347
rect 135 -381 151 -347
rect 203 -381 219 -347
rect 253 -381 269 -347
rect -269 -489 -253 -455
rect -219 -489 -203 -455
rect -151 -489 -135 -455
rect -101 -489 -85 -455
rect -33 -489 -17 -455
rect 17 -489 33 -455
rect 85 -489 101 -455
rect 135 -489 151 -455
rect 203 -489 219 -455
rect 253 -489 269 -455
rect -312 -548 -278 -532
rect -312 -1140 -278 -1124
rect -194 -548 -160 -532
rect -194 -1140 -160 -1124
rect -76 -548 -42 -532
rect -76 -1140 -42 -1124
rect 42 -548 76 -532
rect 42 -1140 76 -1124
rect 160 -548 194 -532
rect 160 -1140 194 -1124
rect 278 -548 312 -532
rect 278 -1140 312 -1124
rect -269 -1217 -253 -1183
rect -219 -1217 -203 -1183
rect -151 -1217 -135 -1183
rect -101 -1217 -85 -1183
rect -33 -1217 -17 -1183
rect 17 -1217 33 -1183
rect 85 -1217 101 -1183
rect 135 -1217 151 -1183
rect 203 -1217 219 -1183
rect 253 -1217 269 -1183
rect -426 -1285 -392 -1223
rect 392 -1285 426 -1223
rect -426 -1319 -330 -1285
rect 330 -1319 426 -1285
<< viali >>
rect -253 1183 -219 1217
rect -135 1183 -101 1217
rect -17 1183 17 1217
rect 101 1183 135 1217
rect 219 1183 253 1217
rect -312 548 -278 1124
rect -194 548 -160 1124
rect -76 548 -42 1124
rect 42 548 76 1124
rect 160 548 194 1124
rect 278 548 312 1124
rect -253 455 -219 489
rect -135 455 -101 489
rect -17 455 17 489
rect 101 455 135 489
rect 219 455 253 489
rect -253 347 -219 381
rect -135 347 -101 381
rect -17 347 17 381
rect 101 347 135 381
rect 219 347 253 381
rect -312 -288 -278 288
rect -194 -288 -160 288
rect -76 -288 -42 288
rect 42 -288 76 288
rect 160 -288 194 288
rect 278 -288 312 288
rect -253 -381 -219 -347
rect -135 -381 -101 -347
rect -17 -381 17 -347
rect 101 -381 135 -347
rect 219 -381 253 -347
rect -253 -489 -219 -455
rect -135 -489 -101 -455
rect -17 -489 17 -455
rect 101 -489 135 -455
rect 219 -489 253 -455
rect -312 -1124 -278 -548
rect -194 -1124 -160 -548
rect -76 -1124 -42 -548
rect 42 -1124 76 -548
rect 160 -1124 194 -548
rect 278 -1124 312 -548
rect -253 -1217 -219 -1183
rect -135 -1217 -101 -1183
rect -17 -1217 17 -1183
rect 101 -1217 135 -1183
rect 219 -1217 253 -1183
<< metal1 >>
rect -265 1217 -207 1223
rect -265 1183 -253 1217
rect -219 1183 -207 1217
rect -265 1177 -207 1183
rect -147 1217 -89 1223
rect -147 1183 -135 1217
rect -101 1183 -89 1217
rect -147 1177 -89 1183
rect -29 1217 29 1223
rect -29 1183 -17 1217
rect 17 1183 29 1217
rect -29 1177 29 1183
rect 89 1217 147 1223
rect 89 1183 101 1217
rect 135 1183 147 1217
rect 89 1177 147 1183
rect 207 1217 265 1223
rect 207 1183 219 1217
rect 253 1183 265 1217
rect 207 1177 265 1183
rect -318 1124 -272 1136
rect -318 548 -312 1124
rect -278 548 -272 1124
rect -318 536 -272 548
rect -200 1124 -154 1136
rect -200 548 -194 1124
rect -160 548 -154 1124
rect -200 536 -154 548
rect -82 1124 -36 1136
rect -82 548 -76 1124
rect -42 548 -36 1124
rect -82 536 -36 548
rect 36 1124 82 1136
rect 36 548 42 1124
rect 76 548 82 1124
rect 36 536 82 548
rect 154 1124 200 1136
rect 154 548 160 1124
rect 194 548 200 1124
rect 154 536 200 548
rect 272 1124 318 1136
rect 272 548 278 1124
rect 312 548 318 1124
rect 272 536 318 548
rect -265 489 -207 495
rect -265 455 -253 489
rect -219 455 -207 489
rect -265 449 -207 455
rect -147 489 -89 495
rect -147 455 -135 489
rect -101 455 -89 489
rect -147 449 -89 455
rect -29 489 29 495
rect -29 455 -17 489
rect 17 455 29 489
rect -29 449 29 455
rect 89 489 147 495
rect 89 455 101 489
rect 135 455 147 489
rect 89 449 147 455
rect 207 489 265 495
rect 207 455 219 489
rect 253 455 265 489
rect 207 449 265 455
rect -265 381 -207 387
rect -265 347 -253 381
rect -219 347 -207 381
rect -265 341 -207 347
rect -147 381 -89 387
rect -147 347 -135 381
rect -101 347 -89 381
rect -147 341 -89 347
rect -29 381 29 387
rect -29 347 -17 381
rect 17 347 29 381
rect -29 341 29 347
rect 89 381 147 387
rect 89 347 101 381
rect 135 347 147 381
rect 89 341 147 347
rect 207 381 265 387
rect 207 347 219 381
rect 253 347 265 381
rect 207 341 265 347
rect -318 288 -272 300
rect -318 -288 -312 288
rect -278 -288 -272 288
rect -318 -300 -272 -288
rect -200 288 -154 300
rect -200 -288 -194 288
rect -160 -288 -154 288
rect -200 -300 -154 -288
rect -82 288 -36 300
rect -82 -288 -76 288
rect -42 -288 -36 288
rect -82 -300 -36 -288
rect 36 288 82 300
rect 36 -288 42 288
rect 76 -288 82 288
rect 36 -300 82 -288
rect 154 288 200 300
rect 154 -288 160 288
rect 194 -288 200 288
rect 154 -300 200 -288
rect 272 288 318 300
rect 272 -288 278 288
rect 312 -288 318 288
rect 272 -300 318 -288
rect -265 -347 -207 -341
rect -265 -381 -253 -347
rect -219 -381 -207 -347
rect -265 -387 -207 -381
rect -147 -347 -89 -341
rect -147 -381 -135 -347
rect -101 -381 -89 -347
rect -147 -387 -89 -381
rect -29 -347 29 -341
rect -29 -381 -17 -347
rect 17 -381 29 -347
rect -29 -387 29 -381
rect 89 -347 147 -341
rect 89 -381 101 -347
rect 135 -381 147 -347
rect 89 -387 147 -381
rect 207 -347 265 -341
rect 207 -381 219 -347
rect 253 -381 265 -347
rect 207 -387 265 -381
rect -265 -455 -207 -449
rect -265 -489 -253 -455
rect -219 -489 -207 -455
rect -265 -495 -207 -489
rect -147 -455 -89 -449
rect -147 -489 -135 -455
rect -101 -489 -89 -455
rect -147 -495 -89 -489
rect -29 -455 29 -449
rect -29 -489 -17 -455
rect 17 -489 29 -455
rect -29 -495 29 -489
rect 89 -455 147 -449
rect 89 -489 101 -455
rect 135 -489 147 -455
rect 89 -495 147 -489
rect 207 -455 265 -449
rect 207 -489 219 -455
rect 253 -489 265 -455
rect 207 -495 265 -489
rect -318 -548 -272 -536
rect -318 -1124 -312 -548
rect -278 -1124 -272 -548
rect -318 -1136 -272 -1124
rect -200 -548 -154 -536
rect -200 -1124 -194 -548
rect -160 -1124 -154 -548
rect -200 -1136 -154 -1124
rect -82 -548 -36 -536
rect -82 -1124 -76 -548
rect -42 -1124 -36 -548
rect -82 -1136 -36 -1124
rect 36 -548 82 -536
rect 36 -1124 42 -548
rect 76 -1124 82 -548
rect 36 -1136 82 -1124
rect 154 -548 200 -536
rect 154 -1124 160 -548
rect 194 -1124 200 -548
rect 154 -1136 200 -1124
rect 272 -548 318 -536
rect 272 -1124 278 -548
rect 312 -1124 318 -548
rect 272 -1136 318 -1124
rect -265 -1183 -207 -1177
rect -265 -1217 -253 -1183
rect -219 -1217 -207 -1183
rect -265 -1223 -207 -1217
rect -147 -1183 -89 -1177
rect -147 -1217 -135 -1183
rect -101 -1217 -89 -1183
rect -147 -1223 -89 -1217
rect -29 -1183 29 -1177
rect -29 -1217 -17 -1183
rect 17 -1217 29 -1183
rect -29 -1223 29 -1217
rect 89 -1183 147 -1177
rect 89 -1217 101 -1183
rect 135 -1217 147 -1183
rect 89 -1223 147 -1217
rect 207 -1183 265 -1177
rect 207 -1217 219 -1183
rect 253 -1217 265 -1183
rect 207 -1223 265 -1217
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string FIXED_BBOX -409 -1302 409 1302
string parameters w 3 l 0.3 m 3 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viagl 0 viagr 0 viagt 0 viagb 0 viagate 100 viadrn 100 viasrc 100
string library sky130
<< end >>
