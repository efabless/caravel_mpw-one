magic
tech sky130A
magscale 12 1
timestamp 1598769811
<< metal5 >>
rect 0 70 15 105
rect 30 70 45 105
rect 0 60 45 70
rect 5 50 40 60
rect 10 40 35 50
rect 15 0 30 40
<< properties >>
string FIXED_BBOX 0 -30 60 105
<< end >>
