magic
tech sky130A
timestamp 1624145270
<< checkpaint >>
rect -4918 -4383 296880 356351
<< metal2 >>
rect 4043 351760 4099 352480
rect 12139 351760 12195 352480
rect 20235 351760 20291 352480
rect 28377 351760 28433 352480
rect 36473 351760 36529 352480
rect 44569 351760 44625 352480
rect 52711 351760 52767 352480
rect 60807 351760 60863 352480
rect 68903 351760 68959 352480
rect 77045 351760 77101 352480
rect 85141 351760 85197 352480
rect 93237 351760 93293 352480
rect 101379 351760 101435 352480
rect 109475 351760 109531 352480
rect 117571 351760 117627 352480
rect 125713 351760 125769 352480
rect 133809 351760 133865 352480
rect 141905 351760 141961 352480
rect 150047 351760 150103 352480
rect 158143 351760 158199 352480
rect 166239 351760 166295 352480
rect 174381 351760 174437 352480
rect 182477 351760 182533 352480
rect 190573 351760 190629 352480
rect 198715 351760 198771 352480
rect 206811 351760 206867 352480
rect 214907 351760 214963 352480
rect 223049 351760 223105 352480
rect 231145 351760 231201 352480
rect 239241 351760 239297 352480
rect 247383 351760 247439 352480
rect 255479 351760 255535 352480
rect 263575 351760 263631 352480
rect 271717 351760 271773 352480
rect 279813 351760 279869 352480
rect 287909 351760 287965 352480
rect 271 -480 327 240
rect 823 -480 879 240
rect 1421 -480 1477 240
rect 2019 -480 2075 240
rect 2617 -480 2673 240
rect 3215 -480 3271 240
rect 3813 -480 3869 240
rect 4411 -480 4467 240
rect 5009 -480 5065 240
rect 5607 -480 5663 240
rect 6205 -480 6261 240
rect 6803 -480 6859 240
rect 7401 -480 7457 240
rect 7999 -480 8055 240
rect 8597 -480 8653 240
rect 9149 -480 9205 240
rect 9747 -480 9803 240
rect 10345 -480 10401 240
rect 10943 -480 10999 240
rect 11541 -480 11597 240
rect 12139 -480 12195 240
rect 12737 -480 12793 240
rect 13335 -480 13391 240
rect 13933 -480 13989 240
rect 14531 -480 14587 240
rect 15129 -480 15185 240
rect 15727 -480 15783 240
rect 16325 -480 16381 240
rect 16923 -480 16979 240
rect 17475 -480 17531 240
rect 18073 -480 18129 240
rect 18671 -480 18727 240
rect 19269 -480 19325 240
rect 19867 -480 19923 240
rect 20465 -480 20521 240
rect 21063 -480 21119 240
rect 21661 -480 21717 240
rect 22259 -480 22315 240
rect 22857 -480 22913 240
rect 23455 -480 23511 240
rect 24053 -480 24109 240
rect 24651 -480 24707 240
rect 25249 -480 25305 240
rect 25801 -480 25857 240
rect 26399 -480 26455 240
rect 26997 -480 27053 240
rect 27595 -480 27651 240
rect 28193 -480 28249 240
rect 28791 -480 28847 240
rect 29389 -480 29445 240
rect 29987 -480 30043 240
rect 30585 -480 30641 240
rect 31183 -480 31239 240
rect 31781 -480 31837 240
rect 32379 -480 32435 240
rect 32977 -480 33033 240
rect 33575 -480 33631 240
rect 34127 -480 34183 240
rect 34725 -480 34781 240
rect 35323 -480 35379 240
rect 35921 -480 35977 240
rect 36519 -480 36575 240
rect 37117 -480 37173 240
rect 37715 -480 37771 240
rect 38313 -480 38369 240
rect 38911 -480 38967 240
rect 39509 -480 39565 240
rect 40107 -480 40163 240
rect 40705 -480 40761 240
rect 41303 -480 41359 240
rect 41901 -480 41957 240
rect 42453 -480 42509 240
rect 43051 -480 43107 240
rect 43649 -480 43705 240
rect 44247 -480 44303 240
rect 44845 -480 44901 240
rect 45443 -480 45499 240
rect 46041 -480 46097 240
rect 46639 -480 46695 240
rect 47237 -480 47293 240
rect 47835 -480 47891 240
rect 48433 -480 48489 240
rect 49031 -480 49087 240
rect 49629 -480 49685 240
rect 50227 -480 50283 240
rect 50779 -480 50835 240
rect 51377 -480 51433 240
rect 51975 -480 52031 240
rect 52573 -480 52629 240
rect 53171 -480 53227 240
rect 53769 -480 53825 240
rect 54367 -480 54423 240
rect 54965 -480 55021 240
rect 55563 -480 55619 240
rect 56161 -480 56217 240
rect 56759 -480 56815 240
rect 57357 -480 57413 240
rect 57955 -480 58011 240
rect 58553 -480 58609 240
rect 59105 -480 59161 240
rect 59703 -480 59759 240
rect 60301 -480 60357 240
rect 60899 -480 60955 240
rect 61497 -480 61553 240
rect 62095 -480 62151 240
rect 62693 -480 62749 240
rect 63291 -480 63347 240
rect 63889 -480 63945 240
rect 64487 -480 64543 240
rect 65085 -480 65141 240
rect 65683 -480 65739 240
rect 66281 -480 66337 240
rect 66879 -480 66935 240
rect 67431 -480 67487 240
rect 68029 -480 68085 240
rect 68627 -480 68683 240
rect 69225 -480 69281 240
rect 69823 -480 69879 240
rect 70421 -480 70477 240
rect 71019 -480 71075 240
rect 71617 -480 71673 240
rect 72215 -480 72271 240
rect 72813 -480 72869 240
rect 73411 -480 73467 240
rect 74009 -480 74065 240
rect 74607 -480 74663 240
rect 75205 -480 75261 240
rect 75757 -480 75813 240
rect 76355 -480 76411 240
rect 76953 -480 77009 240
rect 77551 -480 77607 240
rect 78149 -480 78205 240
rect 78747 -480 78803 240
rect 79345 -480 79401 240
rect 79943 -480 79999 240
rect 80541 -480 80597 240
rect 81139 -480 81195 240
rect 81737 -480 81793 240
rect 82335 -480 82391 240
rect 82933 -480 82989 240
rect 83531 -480 83587 240
rect 84083 -480 84139 240
rect 84681 -480 84737 240
rect 85279 -480 85335 240
rect 85877 -480 85933 240
rect 86475 -480 86531 240
rect 87073 -480 87129 240
rect 87671 -480 87727 240
rect 88269 -480 88325 240
rect 88867 -480 88923 240
rect 89465 -480 89521 240
rect 90063 -480 90119 240
rect 90661 -480 90717 240
rect 91259 -480 91315 240
rect 91857 -480 91913 240
rect 92409 -480 92465 240
rect 93007 -480 93063 240
rect 93605 -480 93661 240
rect 94203 -480 94259 240
rect 94801 -480 94857 240
rect 95399 -480 95455 240
rect 95997 -480 96053 240
rect 96595 -480 96651 240
rect 97193 -480 97249 240
rect 97791 -480 97847 240
rect 98389 -480 98445 240
rect 98987 -480 99043 240
rect 99585 -480 99641 240
rect 100183 -480 100239 240
rect 100735 -480 100791 240
rect 101333 -480 101389 240
rect 101931 -480 101987 240
rect 102529 -480 102585 240
rect 103127 -480 103183 240
rect 103725 -480 103781 240
rect 104323 -480 104379 240
rect 104921 -480 104977 240
rect 105519 -480 105575 240
rect 106117 -480 106173 240
rect 106715 -480 106771 240
rect 107313 -480 107369 240
rect 107911 -480 107967 240
rect 108509 -480 108565 240
rect 109061 -480 109117 240
rect 109659 -480 109715 240
rect 110257 -480 110313 240
rect 110855 -480 110911 240
rect 111453 -480 111509 240
rect 112051 -480 112107 240
rect 112649 -480 112705 240
rect 113247 -480 113303 240
rect 113845 -480 113901 240
rect 114443 -480 114499 240
rect 115041 -480 115097 240
rect 115639 -480 115695 240
rect 116237 -480 116293 240
rect 116835 -480 116891 240
rect 117387 -480 117443 240
rect 117985 -480 118041 240
rect 118583 -480 118639 240
rect 119181 -480 119237 240
rect 119779 -480 119835 240
rect 120377 -480 120433 240
rect 120975 -480 121031 240
rect 121573 -480 121629 240
rect 122171 -480 122227 240
rect 122769 -480 122825 240
rect 123367 -480 123423 240
rect 123965 -480 124021 240
rect 124563 -480 124619 240
rect 125161 -480 125217 240
rect 125713 -480 125769 240
rect 126311 -480 126367 240
rect 126909 -480 126965 240
rect 127507 -480 127563 240
rect 128105 -480 128161 240
rect 128703 -480 128759 240
rect 129301 -480 129357 240
rect 129899 -480 129955 240
rect 130497 -480 130553 240
rect 131095 -480 131151 240
rect 131693 -480 131749 240
rect 132291 -480 132347 240
rect 132889 -480 132945 240
rect 133487 -480 133543 240
rect 134039 -480 134095 240
rect 134637 -480 134693 240
rect 135235 -480 135291 240
rect 135833 -480 135889 240
rect 136431 -480 136487 240
rect 137029 -480 137085 240
rect 137627 -480 137683 240
rect 138225 -480 138281 240
rect 138823 -480 138879 240
rect 139421 -480 139477 240
rect 140019 -480 140075 240
rect 140617 -480 140673 240
rect 141215 -480 141271 240
rect 141813 -480 141869 240
rect 142365 -480 142421 240
rect 142963 -480 143019 240
rect 143561 -480 143617 240
rect 144159 -480 144215 240
rect 144757 -480 144813 240
rect 145355 -480 145411 240
rect 145953 -480 146009 240
rect 146551 -480 146607 240
rect 147149 -480 147205 240
rect 147747 -480 147803 240
rect 148345 -480 148401 240
rect 148943 -480 148999 240
rect 149541 -480 149597 240
rect 150139 -480 150195 240
rect 150691 -480 150747 240
rect 151289 -480 151345 240
rect 151887 -480 151943 240
rect 152485 -480 152541 240
rect 153083 -480 153139 240
rect 153681 -480 153737 240
rect 154279 -480 154335 240
rect 154877 -480 154933 240
rect 155475 -480 155531 240
rect 156073 -480 156129 240
rect 156671 -480 156727 240
rect 157269 -480 157325 240
rect 157867 -480 157923 240
rect 158465 -480 158521 240
rect 159017 -480 159073 240
rect 159615 -480 159671 240
rect 160213 -480 160269 240
rect 160811 -480 160867 240
rect 161409 -480 161465 240
rect 162007 -480 162063 240
rect 162605 -480 162661 240
rect 163203 -480 163259 240
rect 163801 -480 163857 240
rect 164399 -480 164455 240
rect 164997 -480 165053 240
rect 165595 -480 165651 240
rect 166193 -480 166249 240
rect 166791 -480 166847 240
rect 167343 -480 167399 240
rect 167941 -480 167997 240
rect 168539 -480 168595 240
rect 169137 -480 169193 240
rect 169735 -480 169791 240
rect 170333 -480 170389 240
rect 170931 -480 170987 240
rect 171529 -480 171585 240
rect 172127 -480 172183 240
rect 172725 -480 172781 240
rect 173323 -480 173379 240
rect 173921 -480 173977 240
rect 174519 -480 174575 240
rect 175117 -480 175173 240
rect 175669 -480 175725 240
rect 176267 -480 176323 240
rect 176865 -480 176921 240
rect 177463 -480 177519 240
rect 178061 -480 178117 240
rect 178659 -480 178715 240
rect 179257 -480 179313 240
rect 179855 -480 179911 240
rect 180453 -480 180509 240
rect 181051 -480 181107 240
rect 181649 -480 181705 240
rect 182247 -480 182303 240
rect 182845 -480 182901 240
rect 183443 -480 183499 240
rect 183995 -480 184051 240
rect 184593 -480 184649 240
rect 185191 -480 185247 240
rect 185789 -480 185845 240
rect 186387 -480 186443 240
rect 186985 -480 187041 240
rect 187583 -480 187639 240
rect 188181 -480 188237 240
rect 188779 -480 188835 240
rect 189377 -480 189433 240
rect 189975 -480 190031 240
rect 190573 -480 190629 240
rect 191171 -480 191227 240
rect 191769 -480 191825 240
rect 192321 -480 192377 240
rect 192919 -480 192975 240
rect 193517 -480 193573 240
rect 194115 -480 194171 240
rect 194713 -480 194769 240
rect 195311 -480 195367 240
rect 195909 -480 195965 240
rect 196507 -480 196563 240
rect 197105 -480 197161 240
rect 197703 -480 197759 240
rect 198301 -480 198357 240
rect 198899 -480 198955 240
rect 199497 -480 199553 240
rect 200095 -480 200151 240
rect 200647 -480 200703 240
rect 201245 -480 201301 240
rect 201843 -480 201899 240
rect 202441 -480 202497 240
rect 203039 -480 203095 240
rect 203637 -480 203693 240
rect 204235 -480 204291 240
rect 204833 -480 204889 240
rect 205431 -480 205487 240
rect 206029 -480 206085 240
rect 206627 -480 206683 240
rect 207225 -480 207281 240
rect 207823 -480 207879 240
rect 208421 -480 208477 240
rect 208973 -480 209029 240
rect 209571 -480 209627 240
rect 210169 -480 210225 240
rect 210767 -480 210823 240
rect 211365 -480 211421 240
rect 211963 -480 212019 240
rect 212561 -480 212617 240
rect 213159 -480 213215 240
rect 213757 -480 213813 240
rect 214355 -480 214411 240
rect 214953 -480 215009 240
rect 215551 -480 215607 240
rect 216149 -480 216205 240
rect 216747 -480 216803 240
rect 217299 -480 217355 240
rect 217897 -480 217953 240
rect 218495 -480 218551 240
rect 219093 -480 219149 240
rect 219691 -480 219747 240
rect 220289 -480 220345 240
rect 220887 -480 220943 240
rect 221485 -480 221541 240
rect 222083 -480 222139 240
rect 222681 -480 222737 240
rect 223279 -480 223335 240
rect 223877 -480 223933 240
rect 224475 -480 224531 240
rect 225073 -480 225129 240
rect 225625 -480 225681 240
rect 226223 -480 226279 240
rect 226821 -480 226877 240
rect 227419 -480 227475 240
rect 228017 -480 228073 240
rect 228615 -480 228671 240
rect 229213 -480 229269 240
rect 229811 -480 229867 240
rect 230409 -480 230465 240
rect 231007 -480 231063 240
rect 231605 -480 231661 240
rect 232203 -480 232259 240
rect 232801 -480 232857 240
rect 233399 -480 233455 240
rect 233951 -480 234007 240
rect 234549 -480 234605 240
rect 235147 -480 235203 240
rect 235745 -480 235801 240
rect 236343 -480 236399 240
rect 236941 -480 236997 240
rect 237539 -480 237595 240
rect 238137 -480 238193 240
rect 238735 -480 238791 240
rect 239333 -480 239389 240
rect 239931 -480 239987 240
rect 240529 -480 240585 240
rect 241127 -480 241183 240
rect 241725 -480 241781 240
rect 242277 -480 242333 240
rect 242875 -480 242931 240
rect 243473 -480 243529 240
rect 244071 -480 244127 240
rect 244669 -480 244725 240
rect 245267 -480 245323 240
rect 245865 -480 245921 240
rect 246463 -480 246519 240
rect 247061 -480 247117 240
rect 247659 -480 247715 240
rect 248257 -480 248313 240
rect 248855 -480 248911 240
rect 249453 -480 249509 240
rect 250051 -480 250107 240
rect 250603 -480 250659 240
rect 251201 -480 251257 240
rect 251799 -480 251855 240
rect 252397 -480 252453 240
rect 252995 -480 253051 240
rect 253593 -480 253649 240
rect 254191 -480 254247 240
rect 254789 -480 254845 240
rect 255387 -480 255443 240
rect 255985 -480 256041 240
rect 256583 -480 256639 240
rect 257181 -480 257237 240
rect 257779 -480 257835 240
rect 258377 -480 258433 240
rect 258929 -480 258985 240
rect 259527 -480 259583 240
rect 260125 -480 260181 240
rect 260723 -480 260779 240
rect 261321 -480 261377 240
rect 261919 -480 261975 240
rect 262517 -480 262573 240
rect 263115 -480 263171 240
rect 263713 -480 263769 240
rect 264311 -480 264367 240
rect 264909 -480 264965 240
rect 265507 -480 265563 240
rect 266105 -480 266161 240
rect 266703 -480 266759 240
rect 267255 -480 267311 240
rect 267853 -480 267909 240
rect 268451 -480 268507 240
rect 269049 -480 269105 240
rect 269647 -480 269703 240
rect 270245 -480 270301 240
rect 270843 -480 270899 240
rect 271441 -480 271497 240
rect 272039 -480 272095 240
rect 272637 -480 272693 240
rect 273235 -480 273291 240
rect 273833 -480 273889 240
rect 274431 -480 274487 240
rect 275029 -480 275085 240
rect 275581 -480 275637 240
rect 276179 -480 276235 240
rect 276777 -480 276833 240
rect 277375 -480 277431 240
rect 277973 -480 278029 240
rect 278571 -480 278627 240
rect 279169 -480 279225 240
rect 279767 -480 279823 240
rect 280365 -480 280421 240
rect 280963 -480 281019 240
rect 281561 -480 281617 240
rect 282159 -480 282215 240
rect 282757 -480 282813 240
rect 283355 -480 283411 240
rect 283907 -480 283963 240
rect 284505 -480 284561 240
rect 285103 -480 285159 240
rect 285701 -480 285757 240
rect 286299 -480 286355 240
rect 286897 -480 286953 240
rect 287495 -480 287551 240
rect 288093 -480 288149 240
rect 288691 -480 288747 240
rect 289289 -480 289345 240
rect 289887 -480 289943 240
rect 290485 -480 290541 240
rect 291083 -480 291139 240
rect 291681 -480 291737 240
<< metal3 >>
rect 291760 348950 292480 349070
rect -480 348270 240 348390
rect 291760 343102 292480 343222
rect -480 341062 240 341182
rect 291760 337254 292480 337374
rect -480 333922 240 334042
rect 291760 331338 292480 331458
rect -480 326714 240 326834
rect 291760 325490 292480 325610
rect 291760 319642 292480 319762
rect -480 319506 240 319626
rect 291760 313794 292480 313914
rect -480 312366 240 312486
rect 291760 307878 292480 307998
rect -480 305158 240 305278
rect 291760 302030 292480 302150
rect -480 297950 240 298070
rect 291760 296182 292480 296302
rect -480 290810 240 290930
rect 291760 290334 292480 290454
rect 291760 284418 292480 284538
rect -480 283602 240 283722
rect 291760 278570 292480 278690
rect -480 276462 240 276582
rect 291760 272722 292480 272842
rect -480 269254 240 269374
rect 291760 266874 292480 266994
rect -480 262046 240 262166
rect 291760 260958 292480 261078
rect 291760 255110 292480 255230
rect -480 254906 240 255026
rect 291760 249262 292480 249382
rect -480 247698 240 247818
rect 291760 243346 292480 243466
rect -480 240490 240 240610
rect 291760 237498 292480 237618
rect -480 233350 240 233470
rect 291760 231650 292480 231770
rect -480 226142 240 226262
rect 291760 225802 292480 225922
rect 291760 219886 292480 220006
rect -480 218934 240 219054
rect 291760 214038 292480 214158
rect -480 211794 240 211914
rect 291760 208190 292480 208310
rect -480 204586 240 204706
rect 291760 202342 292480 202462
rect -480 197446 240 197566
rect 291760 196426 292480 196546
rect 291760 190578 292480 190698
rect -480 190238 240 190358
rect 291760 184730 292480 184850
rect -480 183030 240 183150
rect 291760 178882 292480 179002
rect -480 175890 240 176010
rect 291760 172966 292480 173086
rect -480 168682 240 168802
rect 291760 167118 292480 167238
rect -480 161474 240 161594
rect 291760 161270 292480 161390
rect 291760 155354 292480 155474
rect -480 154334 240 154454
rect 291760 149506 292480 149626
rect -480 147126 240 147246
rect 291760 143658 292480 143778
rect -480 139986 240 140106
rect 291760 137810 292480 137930
rect -480 132778 240 132898
rect 291760 131894 292480 132014
rect 291760 126046 292480 126166
rect -480 125570 240 125690
rect 291760 120198 292480 120318
rect -480 118430 240 118550
rect 291760 114350 292480 114470
rect -480 111222 240 111342
rect 291760 108434 292480 108554
rect -480 104014 240 104134
rect 291760 102586 292480 102706
rect -480 96874 240 96994
rect 291760 96738 292480 96858
rect 291760 90890 292480 91010
rect -480 89666 240 89786
rect 291760 84974 292480 85094
rect -480 82458 240 82578
rect 291760 79126 292480 79246
rect -480 75318 240 75438
rect 291760 73278 292480 73398
rect -480 68110 240 68230
rect 291760 67362 292480 67482
rect 291760 61514 292480 61634
rect -480 60970 240 61090
rect 291760 55666 292480 55786
rect -480 53762 240 53882
rect 291760 49818 292480 49938
rect -480 46554 240 46674
rect 291760 43902 292480 44022
rect -480 39414 240 39534
rect 291760 38054 292480 38174
rect -480 32206 240 32326
rect 291760 32206 292480 32326
rect 291760 26358 292480 26478
rect -480 24998 240 25118
rect 291760 20442 292480 20562
rect -480 17858 240 17978
rect 291760 14594 292480 14714
rect -480 10650 240 10770
rect 291760 8746 292480 8866
rect -480 3510 240 3630
rect 291760 2898 292480 3018
<< metal4 >>
rect -4288 -3752 -3988 355720
rect -3818 -3282 -3518 355250
rect -3348 -2812 -3048 354780
rect -2878 -2342 -2578 354310
rect -2408 -1872 -2108 353840
rect -1938 -1402 -1638 353370
rect -1468 -932 -1168 352900
rect -998 -462 -698 352430
rect 402 351760 702 352900
rect 2202 351760 2502 353840
rect 4002 351760 4302 354780
rect 5802 351760 6102 355720
rect 9402 351760 9702 352900
rect 11202 351760 11502 353840
rect 13002 351760 13302 354780
rect 14802 351760 15102 355720
rect 18402 351760 18702 352900
rect 20202 351760 20502 353840
rect 22002 351760 22302 354780
rect 23802 351760 24102 355720
rect 27402 351760 27702 352900
rect 29202 351760 29502 353840
rect 31002 351760 31302 354780
rect 32802 351760 33102 355720
rect 36402 351760 36702 352900
rect 38202 351760 38502 353840
rect 40002 351760 40302 354780
rect 41802 351760 42102 355720
rect 45402 351760 45702 352900
rect 47202 351760 47502 353840
rect 49002 351760 49302 354780
rect 50802 351760 51102 355720
rect 54402 351760 54702 352900
rect 56202 351760 56502 353840
rect 58002 351760 58302 354780
rect 59802 351760 60102 355720
rect 63402 351760 63702 352900
rect 65202 351760 65502 353840
rect 67002 351760 67302 354780
rect 68802 351760 69102 355720
rect 72402 351760 72702 352900
rect 74202 351760 74502 353840
rect 76002 351760 76302 354780
rect 77802 351760 78102 355720
rect 81402 351760 81702 352900
rect 83202 351760 83502 353840
rect 85002 351760 85302 354780
rect 86802 351760 87102 355720
rect 90402 351760 90702 352900
rect 92202 351760 92502 353840
rect 94002 351760 94302 354780
rect 95802 351760 96102 355720
rect 99402 351760 99702 352900
rect 101202 351760 101502 353840
rect 103002 351760 103302 354780
rect 104802 351760 105102 355720
rect 108402 351760 108702 352900
rect 110202 351760 110502 353840
rect 112002 351760 112302 354780
rect 113802 351760 114102 355720
rect 117402 351760 117702 352900
rect 119202 351760 119502 353840
rect 121002 351760 121302 354780
rect 122802 351760 123102 355720
rect 126402 351760 126702 352900
rect 128202 351760 128502 353840
rect 130002 351760 130302 354780
rect 131802 351760 132102 355720
rect 135402 351760 135702 352900
rect 137202 351760 137502 353840
rect 139002 351760 139302 354780
rect 140802 351760 141102 355720
rect 144402 351760 144702 352900
rect 146202 351760 146502 353840
rect 148002 351760 148302 354780
rect 149802 351760 150102 355720
rect 153402 351760 153702 352900
rect 155202 351760 155502 353840
rect 157002 351760 157302 354780
rect 158802 351760 159102 355720
rect 162402 351760 162702 352900
rect 164202 351760 164502 353840
rect 166002 351760 166302 354780
rect 167802 351760 168102 355720
rect 171402 351760 171702 352900
rect 173202 351760 173502 353840
rect 175002 351760 175302 354780
rect 176802 351760 177102 355720
rect 180402 351760 180702 352900
rect 182202 351760 182502 353840
rect 184002 351760 184302 354780
rect 185802 351760 186102 355720
rect 189402 351760 189702 352900
rect 191202 351760 191502 353840
rect 193002 351760 193302 354780
rect 194802 351760 195102 355720
rect 198402 351760 198702 352900
rect 200202 351760 200502 353840
rect 202002 351760 202302 354780
rect 203802 351760 204102 355720
rect 207402 351760 207702 352900
rect 209202 351760 209502 353840
rect 211002 351760 211302 354780
rect 212802 351760 213102 355720
rect 216402 351760 216702 352900
rect 218202 351760 218502 353840
rect 220002 351760 220302 354780
rect 221802 351760 222102 355720
rect 225402 351760 225702 352900
rect 227202 351760 227502 353840
rect 229002 351760 229302 354780
rect 230802 351760 231102 355720
rect 234402 351760 234702 352900
rect 236202 351760 236502 353840
rect 238002 351760 238302 354780
rect 239802 351760 240102 355720
rect 243402 351760 243702 352900
rect 245202 351760 245502 353840
rect 247002 351760 247302 354780
rect 248802 351760 249102 355720
rect 252402 351760 252702 352900
rect 254202 351760 254502 353840
rect 256002 351760 256302 354780
rect 257802 351760 258102 355720
rect 261402 351760 261702 352900
rect 263202 351760 263502 353840
rect 265002 351760 265302 354780
rect 266802 351760 267102 355720
rect 270402 351760 270702 352900
rect 272202 351760 272502 353840
rect 274002 351760 274302 354780
rect 275802 351760 276102 355720
rect 279402 351760 279702 352900
rect 281202 351760 281502 353840
rect 283002 351760 283302 354780
rect 284802 351760 285102 355720
rect 288402 351760 288702 352900
rect 290202 351760 290502 353840
rect 402 -932 702 240
rect 2202 -1872 2502 240
rect 4002 -2812 4302 240
rect 5802 -3752 6102 240
rect 9402 -932 9702 240
rect 11202 -1872 11502 240
rect 13002 -2812 13302 240
rect 14802 -3752 15102 240
rect 18402 -932 18702 240
rect 20202 -1872 20502 240
rect 22002 -2812 22302 240
rect 23802 -3752 24102 240
rect 27402 -932 27702 240
rect 29202 -1872 29502 240
rect 31002 -2812 31302 240
rect 32802 -3752 33102 240
rect 36402 -932 36702 240
rect 38202 -1872 38502 240
rect 40002 -2812 40302 240
rect 41802 -3752 42102 240
rect 45402 -932 45702 240
rect 47202 -1872 47502 240
rect 49002 -2812 49302 240
rect 50802 -3752 51102 240
rect 54402 -932 54702 240
rect 56202 -1872 56502 240
rect 58002 -2812 58302 240
rect 59802 -3752 60102 240
rect 63402 -932 63702 240
rect 65202 -1872 65502 240
rect 67002 -2812 67302 240
rect 68802 -3752 69102 240
rect 72402 -932 72702 240
rect 74202 -1872 74502 240
rect 76002 -2812 76302 240
rect 77802 -3752 78102 240
rect 81402 -932 81702 240
rect 83202 -1872 83502 240
rect 85002 -2812 85302 240
rect 86802 -3752 87102 240
rect 90402 -932 90702 240
rect 92202 -1872 92502 240
rect 94002 -2812 94302 240
rect 95802 -3752 96102 240
rect 99402 -932 99702 240
rect 101202 -1872 101502 240
rect 103002 -2812 103302 240
rect 104802 -3752 105102 240
rect 108402 -932 108702 240
rect 110202 -1872 110502 240
rect 112002 -2812 112302 240
rect 113802 -3752 114102 240
rect 117402 -932 117702 240
rect 119202 -1872 119502 240
rect 121002 -2812 121302 240
rect 122802 -3752 123102 240
rect 126402 -932 126702 240
rect 128202 -1872 128502 240
rect 130002 -2812 130302 240
rect 131802 -3752 132102 240
rect 135402 -932 135702 240
rect 137202 -1872 137502 240
rect 139002 -2812 139302 240
rect 140802 -3752 141102 240
rect 144402 -932 144702 240
rect 146202 -1872 146502 240
rect 148002 -2812 148302 240
rect 149802 -3752 150102 240
rect 153402 -932 153702 240
rect 155202 -1872 155502 240
rect 157002 -2812 157302 240
rect 158802 -3752 159102 240
rect 162402 -932 162702 240
rect 164202 -1872 164502 240
rect 166002 -2812 166302 240
rect 167802 -3752 168102 240
rect 171402 -932 171702 240
rect 173202 -1872 173502 240
rect 175002 -2812 175302 240
rect 176802 -3752 177102 240
rect 180402 -932 180702 240
rect 182202 -1872 182502 240
rect 184002 -2812 184302 240
rect 185802 -3752 186102 240
rect 189402 -932 189702 240
rect 191202 -1872 191502 240
rect 193002 -2812 193302 240
rect 194802 -3752 195102 240
rect 198402 -932 198702 240
rect 200202 -1872 200502 240
rect 202002 -2812 202302 240
rect 203802 -3752 204102 240
rect 207402 -932 207702 240
rect 209202 -1872 209502 240
rect 211002 -2812 211302 240
rect 212802 -3752 213102 240
rect 216402 -932 216702 240
rect 218202 -1872 218502 240
rect 220002 -2812 220302 240
rect 221802 -3752 222102 240
rect 225402 -932 225702 240
rect 227202 -1872 227502 240
rect 229002 -2812 229302 240
rect 230802 -3752 231102 240
rect 234402 -932 234702 240
rect 236202 -1872 236502 240
rect 238002 -2812 238302 240
rect 239802 -3752 240102 240
rect 243402 -932 243702 240
rect 245202 -1872 245502 240
rect 247002 -2812 247302 240
rect 248802 -3752 249102 240
rect 252402 -932 252702 240
rect 254202 -1872 254502 240
rect 256002 -2812 256302 240
rect 257802 -3752 258102 240
rect 261402 -932 261702 240
rect 263202 -1872 263502 240
rect 265002 -2812 265302 240
rect 266802 -3752 267102 240
rect 270402 -932 270702 240
rect 272202 -1872 272502 240
rect 274002 -2812 274302 240
rect 275802 -3752 276102 240
rect 279402 -932 279702 240
rect 281202 -1872 281502 240
rect 283002 -2812 283302 240
rect 284802 -3752 285102 240
rect 288402 -932 288702 240
rect 290202 -1872 290502 240
rect 292660 -462 292960 352430
rect 293130 -932 293430 352900
rect 293600 -1402 293900 353370
rect 294070 -1872 294370 353840
rect 294540 -2342 294840 354310
rect 295010 -2812 295310 354780
rect 295480 -3282 295780 355250
rect 295950 -3752 296250 355720
<< metal5 >>
rect -4288 355420 296250 355720
rect -3818 354950 295780 355250
rect -3348 354480 295310 354780
rect -2878 354010 294840 354310
rect -2408 353540 294370 353840
rect -1938 353070 293900 353370
rect -1468 352600 293430 352900
rect -998 352130 292960 352430
rect -4288 348338 240 348638
rect 291760 348338 296250 348638
rect -3348 346538 240 346838
rect 291760 346538 295310 346838
rect -2408 344738 240 345038
rect 291760 344738 294370 345038
rect -1468 342938 240 343238
rect 291760 342938 293430 343238
rect -4288 339338 240 339638
rect 291760 339338 296250 339638
rect -3348 337538 240 337838
rect 291760 337538 295310 337838
rect -2408 335738 240 336038
rect 291760 335738 294370 336038
rect -1468 333938 240 334238
rect 291760 333938 293430 334238
rect -4288 330338 240 330638
rect 291760 330338 296250 330638
rect -3348 328538 240 328838
rect 291760 328538 295310 328838
rect -2408 326738 240 327038
rect 291760 326738 294370 327038
rect -1468 324938 240 325238
rect 291760 324938 293430 325238
rect -4288 321338 240 321638
rect 291760 321338 296250 321638
rect -3348 319538 240 319838
rect 291760 319538 295310 319838
rect -2408 317738 240 318038
rect 291760 317738 294370 318038
rect -1468 315938 240 316238
rect 291760 315938 293430 316238
rect -4288 312338 240 312638
rect 291760 312338 296250 312638
rect -3348 310538 240 310838
rect 291760 310538 295310 310838
rect -2408 308738 240 309038
rect 291760 308738 294370 309038
rect -1468 306938 240 307238
rect 291760 306938 293430 307238
rect -4288 303338 240 303638
rect 291760 303338 296250 303638
rect -3348 301538 240 301838
rect 291760 301538 295310 301838
rect -2408 299738 240 300038
rect 291760 299738 294370 300038
rect -1468 297938 240 298238
rect 291760 297938 293430 298238
rect -4288 294338 240 294638
rect 291760 294338 296250 294638
rect -3348 292538 240 292838
rect 291760 292538 295310 292838
rect -2408 290738 240 291038
rect 291760 290738 294370 291038
rect -1468 288938 240 289238
rect 291760 288938 293430 289238
rect -4288 285338 240 285638
rect 291760 285338 296250 285638
rect -3348 283538 240 283838
rect 291760 283538 295310 283838
rect -2408 281738 240 282038
rect 291760 281738 294370 282038
rect -1468 279938 240 280238
rect 291760 279938 293430 280238
rect -4288 276338 240 276638
rect 291760 276338 296250 276638
rect -3348 274538 240 274838
rect 291760 274538 295310 274838
rect -2408 272738 240 273038
rect 291760 272738 294370 273038
rect -1468 270938 240 271238
rect 291760 270938 293430 271238
rect -4288 267338 240 267638
rect 291760 267338 296250 267638
rect -3348 265538 240 265838
rect 291760 265538 295310 265838
rect -2408 263738 240 264038
rect 291760 263738 294370 264038
rect -1468 261938 240 262238
rect 291760 261938 293430 262238
rect -4288 258338 240 258638
rect 291760 258338 296250 258638
rect -3348 256538 240 256838
rect 291760 256538 295310 256838
rect -2408 254738 240 255038
rect 291760 254738 294370 255038
rect -1468 252938 240 253238
rect 291760 252938 293430 253238
rect -4288 249338 240 249638
rect 291760 249338 296250 249638
rect -3348 247538 240 247838
rect 291760 247538 295310 247838
rect -2408 245738 240 246038
rect 291760 245738 294370 246038
rect -1468 243938 240 244238
rect 291760 243938 293430 244238
rect -4288 240338 240 240638
rect 291760 240338 296250 240638
rect -3348 238538 240 238838
rect 291760 238538 295310 238838
rect -2408 236738 240 237038
rect 291760 236738 294370 237038
rect -1468 234938 240 235238
rect 291760 234938 293430 235238
rect -4288 231338 240 231638
rect 291760 231338 296250 231638
rect -3348 229538 240 229838
rect 291760 229538 295310 229838
rect -2408 227738 240 228038
rect 291760 227738 294370 228038
rect -1468 225938 240 226238
rect 291760 225938 293430 226238
rect -4288 222338 240 222638
rect 291760 222338 296250 222638
rect -3348 220538 240 220838
rect 291760 220538 295310 220838
rect -2408 218738 240 219038
rect 291760 218738 294370 219038
rect -1468 216938 240 217238
rect 291760 216938 293430 217238
rect -4288 213338 240 213638
rect 291760 213338 296250 213638
rect -3348 211538 240 211838
rect 291760 211538 295310 211838
rect -2408 209738 240 210038
rect 291760 209738 294370 210038
rect -1468 207938 240 208238
rect 291760 207938 293430 208238
rect -4288 204338 240 204638
rect 291760 204338 296250 204638
rect -3348 202538 240 202838
rect 291760 202538 295310 202838
rect -2408 200738 240 201038
rect 291760 200738 294370 201038
rect -1468 198938 240 199238
rect 291760 198938 293430 199238
rect -4288 195338 240 195638
rect 291760 195338 296250 195638
rect -3348 193538 240 193838
rect 291760 193538 295310 193838
rect -2408 191738 240 192038
rect 291760 191738 294370 192038
rect -1468 189938 240 190238
rect 291760 189938 293430 190238
rect -4288 186338 240 186638
rect 291760 186338 296250 186638
rect -3348 184538 240 184838
rect 291760 184538 295310 184838
rect -2408 182738 240 183038
rect 291760 182738 294370 183038
rect -1468 180938 240 181238
rect 291760 180938 293430 181238
rect -4288 177338 240 177638
rect 291760 177338 296250 177638
rect -3348 175538 240 175838
rect 291760 175538 295310 175838
rect -2408 173738 240 174038
rect 291760 173738 294370 174038
rect -1468 171938 240 172238
rect 291760 171938 293430 172238
rect -4288 168338 240 168638
rect 291760 168338 296250 168638
rect -3348 166538 240 166838
rect 291760 166538 295310 166838
rect -2408 164738 240 165038
rect 291760 164738 294370 165038
rect -1468 162938 240 163238
rect 291760 162938 293430 163238
rect -4288 159338 240 159638
rect 291760 159338 296250 159638
rect -3348 157538 240 157838
rect 291760 157538 295310 157838
rect -2408 155738 240 156038
rect 291760 155738 294370 156038
rect -1468 153938 240 154238
rect 291760 153938 293430 154238
rect -4288 150338 240 150638
rect 291760 150338 296250 150638
rect -3348 148538 240 148838
rect 291760 148538 295310 148838
rect -2408 146738 240 147038
rect 291760 146738 294370 147038
rect -1468 144938 240 145238
rect 291760 144938 293430 145238
rect -4288 141338 240 141638
rect 291760 141338 296250 141638
rect -3348 139538 240 139838
rect 291760 139538 295310 139838
rect -2408 137738 240 138038
rect 291760 137738 294370 138038
rect -1468 135938 240 136238
rect 291760 135938 293430 136238
rect -4288 132338 240 132638
rect 291760 132338 296250 132638
rect -3348 130538 240 130838
rect 291760 130538 295310 130838
rect -2408 128738 240 129038
rect 291760 128738 294370 129038
rect -1468 126938 240 127238
rect 291760 126938 293430 127238
rect -4288 123338 240 123638
rect 291760 123338 296250 123638
rect -3348 121538 240 121838
rect 291760 121538 295310 121838
rect -2408 119738 240 120038
rect 291760 119738 294370 120038
rect -1468 117938 240 118238
rect 291760 117938 293430 118238
rect -4288 114338 240 114638
rect 291760 114338 296250 114638
rect -3348 112538 240 112838
rect 291760 112538 295310 112838
rect -2408 110738 240 111038
rect 291760 110738 294370 111038
rect -1468 108938 240 109238
rect 291760 108938 293430 109238
rect -4288 105338 240 105638
rect 291760 105338 296250 105638
rect -3348 103538 240 103838
rect 291760 103538 295310 103838
rect -2408 101738 240 102038
rect 291760 101738 294370 102038
rect -1468 99938 240 100238
rect 291760 99938 293430 100238
rect -4288 96338 240 96638
rect 291760 96338 296250 96638
rect -3348 94538 240 94838
rect 291760 94538 295310 94838
rect -2408 92738 240 93038
rect 291760 92738 294370 93038
rect -1468 90938 240 91238
rect 291760 90938 293430 91238
rect -4288 87338 240 87638
rect 291760 87338 296250 87638
rect -3348 85538 240 85838
rect 291760 85538 295310 85838
rect -2408 83738 240 84038
rect 291760 83738 294370 84038
rect -1468 81938 240 82238
rect 291760 81938 293430 82238
rect -4288 78338 240 78638
rect 291760 78338 296250 78638
rect -3348 76538 240 76838
rect 291760 76538 295310 76838
rect -2408 74738 240 75038
rect 291760 74738 294370 75038
rect -1468 72938 240 73238
rect 291760 72938 293430 73238
rect -4288 69338 240 69638
rect 291760 69338 296250 69638
rect -3348 67538 240 67838
rect 291760 67538 295310 67838
rect -2408 65738 240 66038
rect 291760 65738 294370 66038
rect -1468 63938 240 64238
rect 291760 63938 293430 64238
rect -4288 60338 240 60638
rect 291760 60338 296250 60638
rect -3348 58538 240 58838
rect 291760 58538 295310 58838
rect -2408 56738 240 57038
rect 291760 56738 294370 57038
rect -1468 54938 240 55238
rect 291760 54938 293430 55238
rect -4288 51338 240 51638
rect 291760 51338 296250 51638
rect -3348 49538 240 49838
rect 291760 49538 295310 49838
rect -2408 47738 240 48038
rect 291760 47738 294370 48038
rect -1468 45938 240 46238
rect 291760 45938 293430 46238
rect -4288 42338 240 42638
rect 291760 42338 296250 42638
rect -3348 40538 240 40838
rect 291760 40538 295310 40838
rect -2408 38738 240 39038
rect 291760 38738 294370 39038
rect -1468 36938 240 37238
rect 291760 36938 293430 37238
rect -4288 33338 240 33638
rect 291760 33338 296250 33638
rect -3348 31538 240 31838
rect 291760 31538 295310 31838
rect -2408 29738 240 30038
rect 291760 29738 294370 30038
rect -1468 27938 240 28238
rect 291760 27938 293430 28238
rect -4288 24338 240 24638
rect 291760 24338 296250 24638
rect -3348 22538 240 22838
rect 291760 22538 295310 22838
rect -2408 20738 240 21038
rect 291760 20738 294370 21038
rect -1468 18938 240 19238
rect 291760 18938 293430 19238
rect -4288 15338 240 15638
rect 291760 15338 296250 15638
rect -3348 13538 240 13838
rect 291760 13538 295310 13838
rect -2408 11738 240 12038
rect 291760 11738 294370 12038
rect -1468 9938 240 10238
rect 291760 9938 293430 10238
rect -4288 6338 240 6638
rect 291760 6338 296250 6638
rect -3348 4538 240 4838
rect 291760 4538 295310 4838
rect -2408 2738 240 3038
rect 291760 2738 294370 3038
rect -1468 938 240 1238
rect 291760 938 293430 1238
rect -998 -462 292960 -162
rect -1468 -932 293430 -632
rect -1938 -1402 293900 -1102
rect -2408 -1872 294370 -1572
rect -2878 -2342 294840 -2042
rect -3348 -2812 295310 -2512
rect -3818 -3282 295780 -2982
rect -4288 -3752 296250 -3452
<< obsm5 >>
rect -4288 355720 -3988 355721
rect 14802 355720 15102 355721
rect 32802 355720 33102 355721
rect 50802 355720 51102 355721
rect 68802 355720 69102 355721
rect 86802 355720 87102 355721
rect 104802 355720 105102 355721
rect 122802 355720 123102 355721
rect 140802 355720 141102 355721
rect 158802 355720 159102 355721
rect 176802 355720 177102 355721
rect 194802 355720 195102 355721
rect 212802 355720 213102 355721
rect 230802 355720 231102 355721
rect 248802 355720 249102 355721
rect 266802 355720 267102 355721
rect 284802 355720 285102 355721
rect 295950 355720 296250 355721
rect -4288 355419 -3988 355420
rect 14802 355419 15102 355420
rect 32802 355419 33102 355420
rect 50802 355419 51102 355420
rect 68802 355419 69102 355420
rect 86802 355419 87102 355420
rect 104802 355419 105102 355420
rect 122802 355419 123102 355420
rect 140802 355419 141102 355420
rect 158802 355419 159102 355420
rect 176802 355419 177102 355420
rect 194802 355419 195102 355420
rect 212802 355419 213102 355420
rect 230802 355419 231102 355420
rect 248802 355419 249102 355420
rect 266802 355419 267102 355420
rect 284802 355419 285102 355420
rect 295950 355419 296250 355420
rect -3818 355250 -3518 355251
rect 5802 355250 6102 355251
rect 23802 355250 24102 355251
rect 41802 355250 42102 355251
rect 59802 355250 60102 355251
rect 77802 355250 78102 355251
rect 95802 355250 96102 355251
rect 113802 355250 114102 355251
rect 131802 355250 132102 355251
rect 149802 355250 150102 355251
rect 167802 355250 168102 355251
rect 185802 355250 186102 355251
rect 203802 355250 204102 355251
rect 221802 355250 222102 355251
rect 239802 355250 240102 355251
rect 257802 355250 258102 355251
rect 275802 355250 276102 355251
rect 295480 355250 295780 355251
rect -3818 354949 -3518 354950
rect 5802 354949 6102 354950
rect 23802 354949 24102 354950
rect 41802 354949 42102 354950
rect 59802 354949 60102 354950
rect 77802 354949 78102 354950
rect 95802 354949 96102 354950
rect 113802 354949 114102 354950
rect 131802 354949 132102 354950
rect 149802 354949 150102 354950
rect 167802 354949 168102 354950
rect 185802 354949 186102 354950
rect 203802 354949 204102 354950
rect 221802 354949 222102 354950
rect 239802 354949 240102 354950
rect 257802 354949 258102 354950
rect 275802 354949 276102 354950
rect 295480 354949 295780 354950
rect -3348 354780 -3048 354781
rect 13002 354780 13302 354781
rect 31002 354780 31302 354781
rect 49002 354780 49302 354781
rect 67002 354780 67302 354781
rect 85002 354780 85302 354781
rect 103002 354780 103302 354781
rect 121002 354780 121302 354781
rect 139002 354780 139302 354781
rect 157002 354780 157302 354781
rect 175002 354780 175302 354781
rect 193002 354780 193302 354781
rect 211002 354780 211302 354781
rect 229002 354780 229302 354781
rect 247002 354780 247302 354781
rect 265002 354780 265302 354781
rect 283002 354780 283302 354781
rect 295010 354780 295310 354781
rect -3348 354479 -3048 354480
rect 13002 354479 13302 354480
rect 31002 354479 31302 354480
rect 49002 354479 49302 354480
rect 67002 354479 67302 354480
rect 85002 354479 85302 354480
rect 103002 354479 103302 354480
rect 121002 354479 121302 354480
rect 139002 354479 139302 354480
rect 157002 354479 157302 354480
rect 175002 354479 175302 354480
rect 193002 354479 193302 354480
rect 211002 354479 211302 354480
rect 229002 354479 229302 354480
rect 247002 354479 247302 354480
rect 265002 354479 265302 354480
rect 283002 354479 283302 354480
rect 295010 354479 295310 354480
rect -2878 354310 -2578 354311
rect 4002 354310 4302 354311
rect 22002 354310 22302 354311
rect 40002 354310 40302 354311
rect 58002 354310 58302 354311
rect 76002 354310 76302 354311
rect 94002 354310 94302 354311
rect 112002 354310 112302 354311
rect 130002 354310 130302 354311
rect 148002 354310 148302 354311
rect 166002 354310 166302 354311
rect 184002 354310 184302 354311
rect 202002 354310 202302 354311
rect 220002 354310 220302 354311
rect 238002 354310 238302 354311
rect 256002 354310 256302 354311
rect 274002 354310 274302 354311
rect 294540 354310 294840 354311
rect -2878 354009 -2578 354010
rect 4002 354009 4302 354010
rect 22002 354009 22302 354010
rect 40002 354009 40302 354010
rect 58002 354009 58302 354010
rect 76002 354009 76302 354010
rect 94002 354009 94302 354010
rect 112002 354009 112302 354010
rect 130002 354009 130302 354010
rect 148002 354009 148302 354010
rect 166002 354009 166302 354010
rect 184002 354009 184302 354010
rect 202002 354009 202302 354010
rect 220002 354009 220302 354010
rect 238002 354009 238302 354010
rect 256002 354009 256302 354010
rect 274002 354009 274302 354010
rect 294540 354009 294840 354010
rect -2408 353840 -2108 353841
rect 11202 353840 11502 353841
rect 29202 353840 29502 353841
rect 47202 353840 47502 353841
rect 65202 353840 65502 353841
rect 83202 353840 83502 353841
rect 101202 353840 101502 353841
rect 119202 353840 119502 353841
rect 137202 353840 137502 353841
rect 155202 353840 155502 353841
rect 173202 353840 173502 353841
rect 191202 353840 191502 353841
rect 209202 353840 209502 353841
rect 227202 353840 227502 353841
rect 245202 353840 245502 353841
rect 263202 353840 263502 353841
rect 281202 353840 281502 353841
rect 294070 353840 294370 353841
rect -2408 353539 -2108 353540
rect 11202 353539 11502 353540
rect 29202 353539 29502 353540
rect 47202 353539 47502 353540
rect 65202 353539 65502 353540
rect 83202 353539 83502 353540
rect 101202 353539 101502 353540
rect 119202 353539 119502 353540
rect 137202 353539 137502 353540
rect 155202 353539 155502 353540
rect 173202 353539 173502 353540
rect 191202 353539 191502 353540
rect 209202 353539 209502 353540
rect 227202 353539 227502 353540
rect 245202 353539 245502 353540
rect 263202 353539 263502 353540
rect 281202 353539 281502 353540
rect 294070 353539 294370 353540
rect -1938 353370 -1638 353371
rect 2202 353370 2502 353371
rect 20202 353370 20502 353371
rect 38202 353370 38502 353371
rect 56202 353370 56502 353371
rect 74202 353370 74502 353371
rect 92202 353370 92502 353371
rect 110202 353370 110502 353371
rect 128202 353370 128502 353371
rect 146202 353370 146502 353371
rect 164202 353370 164502 353371
rect 182202 353370 182502 353371
rect 200202 353370 200502 353371
rect 218202 353370 218502 353371
rect 236202 353370 236502 353371
rect 254202 353370 254502 353371
rect 272202 353370 272502 353371
rect 290202 353370 290502 353371
rect 293600 353370 293900 353371
rect -1938 353069 -1638 353070
rect 2202 353069 2502 353070
rect 20202 353069 20502 353070
rect 38202 353069 38502 353070
rect 56202 353069 56502 353070
rect 74202 353069 74502 353070
rect 92202 353069 92502 353070
rect 110202 353069 110502 353070
rect 128202 353069 128502 353070
rect 146202 353069 146502 353070
rect 164202 353069 164502 353070
rect 182202 353069 182502 353070
rect 200202 353069 200502 353070
rect 218202 353069 218502 353070
rect 236202 353069 236502 353070
rect 254202 353069 254502 353070
rect 272202 353069 272502 353070
rect 290202 353069 290502 353070
rect 293600 353069 293900 353070
rect -1468 352900 -1168 352901
rect 9402 352900 9702 352901
rect 27402 352900 27702 352901
rect 45402 352900 45702 352901
rect 63402 352900 63702 352901
rect 81402 352900 81702 352901
rect 99402 352900 99702 352901
rect 117402 352900 117702 352901
rect 135402 352900 135702 352901
rect 153402 352900 153702 352901
rect 171402 352900 171702 352901
rect 189402 352900 189702 352901
rect 207402 352900 207702 352901
rect 225402 352900 225702 352901
rect 243402 352900 243702 352901
rect 261402 352900 261702 352901
rect 279402 352900 279702 352901
rect 293130 352900 293430 352901
rect -1468 352599 -1168 352600
rect 9402 352599 9702 352600
rect 27402 352599 27702 352600
rect 45402 352599 45702 352600
rect 63402 352599 63702 352600
rect 81402 352599 81702 352600
rect 99402 352599 99702 352600
rect 117402 352599 117702 352600
rect 135402 352599 135702 352600
rect 153402 352599 153702 352600
rect 171402 352599 171702 352600
rect 189402 352599 189702 352600
rect 207402 352599 207702 352600
rect 225402 352599 225702 352600
rect 243402 352599 243702 352600
rect 261402 352599 261702 352600
rect 279402 352599 279702 352600
rect 293130 352599 293430 352600
rect -998 352430 -698 352431
rect 402 352430 702 352431
rect 18402 352430 18702 352431
rect 36402 352430 36702 352431
rect 54402 352430 54702 352431
rect 72402 352430 72702 352431
rect 90402 352430 90702 352431
rect 108402 352430 108702 352431
rect 126402 352430 126702 352431
rect 144402 352430 144702 352431
rect 162402 352430 162702 352431
rect 180402 352430 180702 352431
rect 198402 352430 198702 352431
rect 216402 352430 216702 352431
rect 234402 352430 234702 352431
rect 252402 352430 252702 352431
rect 270402 352430 270702 352431
rect 288402 352430 288702 352431
rect 292660 352430 292960 352431
rect -998 352129 -698 352130
rect 402 352129 702 352130
rect 18402 352129 18702 352130
rect 36402 352129 36702 352130
rect 54402 352129 54702 352130
rect 72402 352129 72702 352130
rect 90402 352129 90702 352130
rect 108402 352129 108702 352130
rect 126402 352129 126702 352130
rect 144402 352129 144702 352130
rect 162402 352129 162702 352130
rect 180402 352129 180702 352130
rect 198402 352129 198702 352130
rect 216402 352129 216702 352130
rect 234402 352129 234702 352130
rect 252402 352129 252702 352130
rect 270402 352129 270702 352130
rect 288402 352129 288702 352130
rect 292660 352129 292960 352130
rect 0 348798 292000 351970
rect -3818 348638 -3518 348639
rect -3818 348337 -3518 348338
rect 400 348178 291600 348798
rect 295480 348638 295780 348639
rect 295480 348337 295780 348338
rect 0 346998 292000 348178
rect -2878 346838 -2578 346839
rect -2878 346537 -2578 346538
rect 400 346378 291600 346998
rect 294540 346838 294840 346839
rect 294540 346537 294840 346538
rect 0 345198 292000 346378
rect -1938 345038 -1638 345039
rect -1938 344737 -1638 344738
rect 400 344578 291600 345198
rect 293600 345038 293900 345039
rect 293600 344737 293900 344738
rect 0 343398 292000 344578
rect -998 343238 -698 343239
rect -998 342937 -698 342938
rect 400 342778 291600 343398
rect 292660 343238 292960 343239
rect 292660 342937 292960 342938
rect 0 339798 292000 342778
rect -4288 339638 -3988 339639
rect -4288 339337 -3988 339338
rect 400 339178 291600 339798
rect 295950 339638 296250 339639
rect 295950 339337 296250 339338
rect 0 337998 292000 339178
rect -3348 337838 -3048 337839
rect -3348 337537 -3048 337538
rect 400 337378 291600 337998
rect 295010 337838 295310 337839
rect 295010 337537 295310 337538
rect 0 336198 292000 337378
rect -2408 336038 -2108 336039
rect -2408 335737 -2108 335738
rect 400 335578 291600 336198
rect 294070 336038 294370 336039
rect 294070 335737 294370 335738
rect 0 334398 292000 335578
rect -1468 334238 -1168 334239
rect -1468 333937 -1168 333938
rect 400 333778 291600 334398
rect 293130 334238 293430 334239
rect 293130 333937 293430 333938
rect 0 330798 292000 333778
rect -3818 330638 -3518 330639
rect -3818 330337 -3518 330338
rect 400 330178 291600 330798
rect 295480 330638 295780 330639
rect 295480 330337 295780 330338
rect 0 328998 292000 330178
rect -2878 328838 -2578 328839
rect -2878 328537 -2578 328538
rect 400 328378 291600 328998
rect 294540 328838 294840 328839
rect 294540 328537 294840 328538
rect 0 327198 292000 328378
rect -1938 327038 -1638 327039
rect -1938 326737 -1638 326738
rect 400 326578 291600 327198
rect 293600 327038 293900 327039
rect 293600 326737 293900 326738
rect 0 325398 292000 326578
rect -998 325238 -698 325239
rect -998 324937 -698 324938
rect 400 324778 291600 325398
rect 292660 325238 292960 325239
rect 292660 324937 292960 324938
rect 0 321798 292000 324778
rect -4288 321638 -3988 321639
rect -4288 321337 -3988 321338
rect 400 321178 291600 321798
rect 295950 321638 296250 321639
rect 295950 321337 296250 321338
rect 0 319998 292000 321178
rect -3348 319838 -3048 319839
rect -3348 319537 -3048 319538
rect 400 319378 291600 319998
rect 295010 319838 295310 319839
rect 295010 319537 295310 319538
rect 0 318198 292000 319378
rect -2408 318038 -2108 318039
rect -2408 317737 -2108 317738
rect 400 317578 291600 318198
rect 294070 318038 294370 318039
rect 294070 317737 294370 317738
rect 0 316398 292000 317578
rect -1468 316238 -1168 316239
rect -1468 315937 -1168 315938
rect 400 315778 291600 316398
rect 293130 316238 293430 316239
rect 293130 315937 293430 315938
rect 0 312798 292000 315778
rect -3818 312638 -3518 312639
rect -3818 312337 -3518 312338
rect 400 312178 291600 312798
rect 295480 312638 295780 312639
rect 295480 312337 295780 312338
rect 0 310998 292000 312178
rect -2878 310838 -2578 310839
rect -2878 310537 -2578 310538
rect 400 310378 291600 310998
rect 294540 310838 294840 310839
rect 294540 310537 294840 310538
rect 0 309198 292000 310378
rect -1938 309038 -1638 309039
rect -1938 308737 -1638 308738
rect 400 308578 291600 309198
rect 293600 309038 293900 309039
rect 293600 308737 293900 308738
rect 0 307398 292000 308578
rect -998 307238 -698 307239
rect -998 306937 -698 306938
rect 400 306778 291600 307398
rect 292660 307238 292960 307239
rect 292660 306937 292960 306938
rect 0 303798 292000 306778
rect -4288 303638 -3988 303639
rect -4288 303337 -3988 303338
rect 400 303178 291600 303798
rect 295950 303638 296250 303639
rect 295950 303337 296250 303338
rect 0 301998 292000 303178
rect -3348 301838 -3048 301839
rect -3348 301537 -3048 301538
rect 400 301378 291600 301998
rect 295010 301838 295310 301839
rect 295010 301537 295310 301538
rect 0 300198 292000 301378
rect -2408 300038 -2108 300039
rect -2408 299737 -2108 299738
rect 400 299578 291600 300198
rect 294070 300038 294370 300039
rect 294070 299737 294370 299738
rect 0 298398 292000 299578
rect -1468 298238 -1168 298239
rect -1468 297937 -1168 297938
rect 400 297778 291600 298398
rect 293130 298238 293430 298239
rect 293130 297937 293430 297938
rect 0 294798 292000 297778
rect -3818 294638 -3518 294639
rect -3818 294337 -3518 294338
rect 400 294178 291600 294798
rect 295480 294638 295780 294639
rect 295480 294337 295780 294338
rect 0 292998 292000 294178
rect -2878 292838 -2578 292839
rect -2878 292537 -2578 292538
rect 400 292378 291600 292998
rect 294540 292838 294840 292839
rect 294540 292537 294840 292538
rect 0 291198 292000 292378
rect -1938 291038 -1638 291039
rect -1938 290737 -1638 290738
rect 400 290578 291600 291198
rect 293600 291038 293900 291039
rect 293600 290737 293900 290738
rect 0 289398 292000 290578
rect -998 289238 -698 289239
rect -998 288937 -698 288938
rect 400 288778 291600 289398
rect 292660 289238 292960 289239
rect 292660 288937 292960 288938
rect 0 285798 292000 288778
rect -4288 285638 -3988 285639
rect -4288 285337 -3988 285338
rect 400 285178 291600 285798
rect 295950 285638 296250 285639
rect 295950 285337 296250 285338
rect 0 283998 292000 285178
rect -3348 283838 -3048 283839
rect -3348 283537 -3048 283538
rect 400 283378 291600 283998
rect 295010 283838 295310 283839
rect 295010 283537 295310 283538
rect 0 282198 292000 283378
rect -2408 282038 -2108 282039
rect -2408 281737 -2108 281738
rect 400 281578 291600 282198
rect 294070 282038 294370 282039
rect 294070 281737 294370 281738
rect 0 280398 292000 281578
rect -1468 280238 -1168 280239
rect -1468 279937 -1168 279938
rect 400 279778 291600 280398
rect 293130 280238 293430 280239
rect 293130 279937 293430 279938
rect 0 276798 292000 279778
rect -3818 276638 -3518 276639
rect -3818 276337 -3518 276338
rect 400 276178 291600 276798
rect 295480 276638 295780 276639
rect 295480 276337 295780 276338
rect 0 274998 292000 276178
rect -2878 274838 -2578 274839
rect -2878 274537 -2578 274538
rect 400 274378 291600 274998
rect 294540 274838 294840 274839
rect 294540 274537 294840 274538
rect 0 273198 292000 274378
rect -1938 273038 -1638 273039
rect -1938 272737 -1638 272738
rect 400 272578 291600 273198
rect 293600 273038 293900 273039
rect 293600 272737 293900 272738
rect 0 271398 292000 272578
rect -998 271238 -698 271239
rect -998 270937 -698 270938
rect 400 270778 291600 271398
rect 292660 271238 292960 271239
rect 292660 270937 292960 270938
rect 0 267798 292000 270778
rect -4288 267638 -3988 267639
rect -4288 267337 -3988 267338
rect 400 267178 291600 267798
rect 295950 267638 296250 267639
rect 295950 267337 296250 267338
rect 0 265998 292000 267178
rect -3348 265838 -3048 265839
rect -3348 265537 -3048 265538
rect 400 265378 291600 265998
rect 295010 265838 295310 265839
rect 295010 265537 295310 265538
rect 0 264198 292000 265378
rect -2408 264038 -2108 264039
rect -2408 263737 -2108 263738
rect 400 263578 291600 264198
rect 294070 264038 294370 264039
rect 294070 263737 294370 263738
rect 0 262398 292000 263578
rect -1468 262238 -1168 262239
rect -1468 261937 -1168 261938
rect 400 261778 291600 262398
rect 293130 262238 293430 262239
rect 293130 261937 293430 261938
rect 0 258798 292000 261778
rect -3818 258638 -3518 258639
rect -3818 258337 -3518 258338
rect 400 258178 291600 258798
rect 295480 258638 295780 258639
rect 295480 258337 295780 258338
rect 0 256998 292000 258178
rect -2878 256838 -2578 256839
rect -2878 256537 -2578 256538
rect 400 256378 291600 256998
rect 294540 256838 294840 256839
rect 294540 256537 294840 256538
rect 0 255198 292000 256378
rect -1938 255038 -1638 255039
rect -1938 254737 -1638 254738
rect 400 254578 291600 255198
rect 293600 255038 293900 255039
rect 293600 254737 293900 254738
rect 0 253398 292000 254578
rect -998 253238 -698 253239
rect -998 252937 -698 252938
rect 400 252778 291600 253398
rect 292660 253238 292960 253239
rect 292660 252937 292960 252938
rect 0 249798 292000 252778
rect -4288 249638 -3988 249639
rect -4288 249337 -3988 249338
rect 400 249178 291600 249798
rect 295950 249638 296250 249639
rect 295950 249337 296250 249338
rect 0 247998 292000 249178
rect -3348 247838 -3048 247839
rect -3348 247537 -3048 247538
rect 400 247378 291600 247998
rect 295010 247838 295310 247839
rect 295010 247537 295310 247538
rect 0 246198 292000 247378
rect -2408 246038 -2108 246039
rect -2408 245737 -2108 245738
rect 400 245578 291600 246198
rect 294070 246038 294370 246039
rect 294070 245737 294370 245738
rect 0 244398 292000 245578
rect -1468 244238 -1168 244239
rect -1468 243937 -1168 243938
rect 400 243778 291600 244398
rect 293130 244238 293430 244239
rect 293130 243937 293430 243938
rect 0 240798 292000 243778
rect -3818 240638 -3518 240639
rect -3818 240337 -3518 240338
rect 400 240178 291600 240798
rect 295480 240638 295780 240639
rect 295480 240337 295780 240338
rect 0 238998 292000 240178
rect -2878 238838 -2578 238839
rect -2878 238537 -2578 238538
rect 400 238378 291600 238998
rect 294540 238838 294840 238839
rect 294540 238537 294840 238538
rect 0 237198 292000 238378
rect -1938 237038 -1638 237039
rect -1938 236737 -1638 236738
rect 400 236578 291600 237198
rect 293600 237038 293900 237039
rect 293600 236737 293900 236738
rect 0 235398 292000 236578
rect -998 235238 -698 235239
rect -998 234937 -698 234938
rect 400 234778 291600 235398
rect 292660 235238 292960 235239
rect 292660 234937 292960 234938
rect 0 231798 292000 234778
rect -4288 231638 -3988 231639
rect -4288 231337 -3988 231338
rect 400 231178 291600 231798
rect 295950 231638 296250 231639
rect 295950 231337 296250 231338
rect 0 229998 292000 231178
rect -3348 229838 -3048 229839
rect -3348 229537 -3048 229538
rect 400 229378 291600 229998
rect 295010 229838 295310 229839
rect 295010 229537 295310 229538
rect 0 228198 292000 229378
rect -2408 228038 -2108 228039
rect -2408 227737 -2108 227738
rect 400 227578 291600 228198
rect 294070 228038 294370 228039
rect 294070 227737 294370 227738
rect 0 226398 292000 227578
rect -1468 226238 -1168 226239
rect -1468 225937 -1168 225938
rect 400 225778 291600 226398
rect 293130 226238 293430 226239
rect 293130 225937 293430 225938
rect 0 222798 292000 225778
rect -3818 222638 -3518 222639
rect -3818 222337 -3518 222338
rect 400 222178 291600 222798
rect 295480 222638 295780 222639
rect 295480 222337 295780 222338
rect 0 220998 292000 222178
rect -2878 220838 -2578 220839
rect -2878 220537 -2578 220538
rect 400 220378 291600 220998
rect 294540 220838 294840 220839
rect 294540 220537 294840 220538
rect 0 219198 292000 220378
rect -1938 219038 -1638 219039
rect -1938 218737 -1638 218738
rect 400 218578 291600 219198
rect 293600 219038 293900 219039
rect 293600 218737 293900 218738
rect 0 217398 292000 218578
rect -998 217238 -698 217239
rect -998 216937 -698 216938
rect 400 216778 291600 217398
rect 292660 217238 292960 217239
rect 292660 216937 292960 216938
rect 0 213798 292000 216778
rect -4288 213638 -3988 213639
rect -4288 213337 -3988 213338
rect 400 213178 291600 213798
rect 295950 213638 296250 213639
rect 295950 213337 296250 213338
rect 0 211998 292000 213178
rect -3348 211838 -3048 211839
rect -3348 211537 -3048 211538
rect 400 211378 291600 211998
rect 295010 211838 295310 211839
rect 295010 211537 295310 211538
rect 0 210198 292000 211378
rect -2408 210038 -2108 210039
rect -2408 209737 -2108 209738
rect 400 209578 291600 210198
rect 294070 210038 294370 210039
rect 294070 209737 294370 209738
rect 0 208398 292000 209578
rect -1468 208238 -1168 208239
rect -1468 207937 -1168 207938
rect 400 207778 291600 208398
rect 293130 208238 293430 208239
rect 293130 207937 293430 207938
rect 0 204798 292000 207778
rect -3818 204638 -3518 204639
rect -3818 204337 -3518 204338
rect 400 204178 291600 204798
rect 295480 204638 295780 204639
rect 295480 204337 295780 204338
rect 0 202998 292000 204178
rect -2878 202838 -2578 202839
rect -2878 202537 -2578 202538
rect 400 202378 291600 202998
rect 294540 202838 294840 202839
rect 294540 202537 294840 202538
rect 0 201198 292000 202378
rect -1938 201038 -1638 201039
rect -1938 200737 -1638 200738
rect 400 200578 291600 201198
rect 293600 201038 293900 201039
rect 293600 200737 293900 200738
rect 0 199398 292000 200578
rect -998 199238 -698 199239
rect -998 198937 -698 198938
rect 400 198778 291600 199398
rect 292660 199238 292960 199239
rect 292660 198937 292960 198938
rect 0 195798 292000 198778
rect -4288 195638 -3988 195639
rect -4288 195337 -3988 195338
rect 400 195178 291600 195798
rect 295950 195638 296250 195639
rect 295950 195337 296250 195338
rect 0 193998 292000 195178
rect -3348 193838 -3048 193839
rect -3348 193537 -3048 193538
rect 400 193378 291600 193998
rect 295010 193838 295310 193839
rect 295010 193537 295310 193538
rect 0 192198 292000 193378
rect -2408 192038 -2108 192039
rect -2408 191737 -2108 191738
rect 400 191578 291600 192198
rect 294070 192038 294370 192039
rect 294070 191737 294370 191738
rect 0 190398 292000 191578
rect -1468 190238 -1168 190239
rect -1468 189937 -1168 189938
rect 400 189778 291600 190398
rect 293130 190238 293430 190239
rect 293130 189937 293430 189938
rect 0 186798 292000 189778
rect -3818 186638 -3518 186639
rect -3818 186337 -3518 186338
rect 400 186178 291600 186798
rect 295480 186638 295780 186639
rect 295480 186337 295780 186338
rect 0 184998 292000 186178
rect -2878 184838 -2578 184839
rect -2878 184537 -2578 184538
rect 400 184378 291600 184998
rect 294540 184838 294840 184839
rect 294540 184537 294840 184538
rect 0 183198 292000 184378
rect -1938 183038 -1638 183039
rect -1938 182737 -1638 182738
rect 400 182578 291600 183198
rect 293600 183038 293900 183039
rect 293600 182737 293900 182738
rect 0 181398 292000 182578
rect -998 181238 -698 181239
rect -998 180937 -698 180938
rect 400 180778 291600 181398
rect 292660 181238 292960 181239
rect 292660 180937 292960 180938
rect 0 177798 292000 180778
rect -4288 177638 -3988 177639
rect -4288 177337 -3988 177338
rect 400 177178 291600 177798
rect 295950 177638 296250 177639
rect 295950 177337 296250 177338
rect 0 175998 292000 177178
rect -3348 175838 -3048 175839
rect -3348 175537 -3048 175538
rect 400 175378 291600 175998
rect 295010 175838 295310 175839
rect 295010 175537 295310 175538
rect 0 174198 292000 175378
rect -2408 174038 -2108 174039
rect -2408 173737 -2108 173738
rect 400 173578 291600 174198
rect 294070 174038 294370 174039
rect 294070 173737 294370 173738
rect 0 172398 292000 173578
rect -1468 172238 -1168 172239
rect -1468 171937 -1168 171938
rect 400 171778 291600 172398
rect 293130 172238 293430 172239
rect 293130 171937 293430 171938
rect 0 168798 292000 171778
rect -3818 168638 -3518 168639
rect -3818 168337 -3518 168338
rect 400 168178 291600 168798
rect 295480 168638 295780 168639
rect 295480 168337 295780 168338
rect 0 166998 292000 168178
rect -2878 166838 -2578 166839
rect -2878 166537 -2578 166538
rect 400 166378 291600 166998
rect 294540 166838 294840 166839
rect 294540 166537 294840 166538
rect 0 165198 292000 166378
rect -1938 165038 -1638 165039
rect -1938 164737 -1638 164738
rect 400 164578 291600 165198
rect 293600 165038 293900 165039
rect 293600 164737 293900 164738
rect 0 163398 292000 164578
rect -998 163238 -698 163239
rect -998 162937 -698 162938
rect 400 162778 291600 163398
rect 292660 163238 292960 163239
rect 292660 162937 292960 162938
rect 0 159798 292000 162778
rect -4288 159638 -3988 159639
rect -4288 159337 -3988 159338
rect 400 159178 291600 159798
rect 295950 159638 296250 159639
rect 295950 159337 296250 159338
rect 0 157998 292000 159178
rect -3348 157838 -3048 157839
rect -3348 157537 -3048 157538
rect 400 157378 291600 157998
rect 295010 157838 295310 157839
rect 295010 157537 295310 157538
rect 0 156198 292000 157378
rect -2408 156038 -2108 156039
rect -2408 155737 -2108 155738
rect 400 155578 291600 156198
rect 294070 156038 294370 156039
rect 294070 155737 294370 155738
rect 0 154398 292000 155578
rect -1468 154238 -1168 154239
rect -1468 153937 -1168 153938
rect 400 153778 291600 154398
rect 293130 154238 293430 154239
rect 293130 153937 293430 153938
rect 0 150798 292000 153778
rect -3818 150638 -3518 150639
rect -3818 150337 -3518 150338
rect 400 150178 291600 150798
rect 295480 150638 295780 150639
rect 295480 150337 295780 150338
rect 0 148998 292000 150178
rect -2878 148838 -2578 148839
rect -2878 148537 -2578 148538
rect 400 148378 291600 148998
rect 294540 148838 294840 148839
rect 294540 148537 294840 148538
rect 0 147198 292000 148378
rect -1938 147038 -1638 147039
rect -1938 146737 -1638 146738
rect 400 146578 291600 147198
rect 293600 147038 293900 147039
rect 293600 146737 293900 146738
rect 0 145398 292000 146578
rect -998 145238 -698 145239
rect -998 144937 -698 144938
rect 400 144778 291600 145398
rect 292660 145238 292960 145239
rect 292660 144937 292960 144938
rect 0 141798 292000 144778
rect -4288 141638 -3988 141639
rect -4288 141337 -3988 141338
rect 400 141178 291600 141798
rect 295950 141638 296250 141639
rect 295950 141337 296250 141338
rect 0 139998 292000 141178
rect -3348 139838 -3048 139839
rect -3348 139537 -3048 139538
rect 400 139378 291600 139998
rect 295010 139838 295310 139839
rect 295010 139537 295310 139538
rect 0 138198 292000 139378
rect -2408 138038 -2108 138039
rect -2408 137737 -2108 137738
rect 400 137578 291600 138198
rect 294070 138038 294370 138039
rect 294070 137737 294370 137738
rect 0 136398 292000 137578
rect -1468 136238 -1168 136239
rect -1468 135937 -1168 135938
rect 400 135778 291600 136398
rect 293130 136238 293430 136239
rect 293130 135937 293430 135938
rect 0 132798 292000 135778
rect -3818 132638 -3518 132639
rect -3818 132337 -3518 132338
rect 400 132178 291600 132798
rect 295480 132638 295780 132639
rect 295480 132337 295780 132338
rect 0 130998 292000 132178
rect -2878 130838 -2578 130839
rect -2878 130537 -2578 130538
rect 400 130378 291600 130998
rect 294540 130838 294840 130839
rect 294540 130537 294840 130538
rect 0 129198 292000 130378
rect -1938 129038 -1638 129039
rect -1938 128737 -1638 128738
rect 400 128578 291600 129198
rect 293600 129038 293900 129039
rect 293600 128737 293900 128738
rect 0 127398 292000 128578
rect -998 127238 -698 127239
rect -998 126937 -698 126938
rect 400 126778 291600 127398
rect 292660 127238 292960 127239
rect 292660 126937 292960 126938
rect 0 123798 292000 126778
rect -4288 123638 -3988 123639
rect -4288 123337 -3988 123338
rect 400 123178 291600 123798
rect 295950 123638 296250 123639
rect 295950 123337 296250 123338
rect 0 121998 292000 123178
rect -3348 121838 -3048 121839
rect -3348 121537 -3048 121538
rect 400 121378 291600 121998
rect 295010 121838 295310 121839
rect 295010 121537 295310 121538
rect 0 120198 292000 121378
rect -2408 120038 -2108 120039
rect -2408 119737 -2108 119738
rect 400 119578 291600 120198
rect 294070 120038 294370 120039
rect 294070 119737 294370 119738
rect 0 118398 292000 119578
rect -1468 118238 -1168 118239
rect -1468 117937 -1168 117938
rect 400 117778 291600 118398
rect 293130 118238 293430 118239
rect 293130 117937 293430 117938
rect 0 114798 292000 117778
rect -3818 114638 -3518 114639
rect -3818 114337 -3518 114338
rect 400 114178 291600 114798
rect 295480 114638 295780 114639
rect 295480 114337 295780 114338
rect 0 112998 292000 114178
rect -2878 112838 -2578 112839
rect -2878 112537 -2578 112538
rect 400 112378 291600 112998
rect 294540 112838 294840 112839
rect 294540 112537 294840 112538
rect 0 111198 292000 112378
rect -1938 111038 -1638 111039
rect -1938 110737 -1638 110738
rect 400 110578 291600 111198
rect 293600 111038 293900 111039
rect 293600 110737 293900 110738
rect 0 109398 292000 110578
rect -998 109238 -698 109239
rect -998 108937 -698 108938
rect 400 108778 291600 109398
rect 292660 109238 292960 109239
rect 292660 108937 292960 108938
rect 0 105798 292000 108778
rect -4288 105638 -3988 105639
rect -4288 105337 -3988 105338
rect 400 105178 291600 105798
rect 295950 105638 296250 105639
rect 295950 105337 296250 105338
rect 0 103998 292000 105178
rect -3348 103838 -3048 103839
rect -3348 103537 -3048 103538
rect 400 103378 291600 103998
rect 295010 103838 295310 103839
rect 295010 103537 295310 103538
rect 0 102198 292000 103378
rect -2408 102038 -2108 102039
rect -2408 101737 -2108 101738
rect 400 101578 291600 102198
rect 294070 102038 294370 102039
rect 294070 101737 294370 101738
rect 0 100398 292000 101578
rect -1468 100238 -1168 100239
rect -1468 99937 -1168 99938
rect 400 99778 291600 100398
rect 293130 100238 293430 100239
rect 293130 99937 293430 99938
rect 0 96798 292000 99778
rect -3818 96638 -3518 96639
rect -3818 96337 -3518 96338
rect 400 96178 291600 96798
rect 295480 96638 295780 96639
rect 295480 96337 295780 96338
rect 0 94998 292000 96178
rect -2878 94838 -2578 94839
rect -2878 94537 -2578 94538
rect 400 94378 291600 94998
rect 294540 94838 294840 94839
rect 294540 94537 294840 94538
rect 0 93198 292000 94378
rect -1938 93038 -1638 93039
rect -1938 92737 -1638 92738
rect 400 92578 291600 93198
rect 293600 93038 293900 93039
rect 293600 92737 293900 92738
rect 0 91398 292000 92578
rect -998 91238 -698 91239
rect -998 90937 -698 90938
rect 400 90778 291600 91398
rect 292660 91238 292960 91239
rect 292660 90937 292960 90938
rect 0 87798 292000 90778
rect -4288 87638 -3988 87639
rect -4288 87337 -3988 87338
rect 400 87178 291600 87798
rect 295950 87638 296250 87639
rect 295950 87337 296250 87338
rect 0 85998 292000 87178
rect -3348 85838 -3048 85839
rect -3348 85537 -3048 85538
rect 400 85378 291600 85998
rect 295010 85838 295310 85839
rect 295010 85537 295310 85538
rect 0 84198 292000 85378
rect -2408 84038 -2108 84039
rect -2408 83737 -2108 83738
rect 400 83578 291600 84198
rect 294070 84038 294370 84039
rect 294070 83737 294370 83738
rect 0 82398 292000 83578
rect -1468 82238 -1168 82239
rect -1468 81937 -1168 81938
rect 400 81778 291600 82398
rect 293130 82238 293430 82239
rect 293130 81937 293430 81938
rect 0 78798 292000 81778
rect -3818 78638 -3518 78639
rect -3818 78337 -3518 78338
rect 400 78178 291600 78798
rect 295480 78638 295780 78639
rect 295480 78337 295780 78338
rect 0 76998 292000 78178
rect -2878 76838 -2578 76839
rect -2878 76537 -2578 76538
rect 400 76378 291600 76998
rect 294540 76838 294840 76839
rect 294540 76537 294840 76538
rect 0 75198 292000 76378
rect -1938 75038 -1638 75039
rect -1938 74737 -1638 74738
rect 400 74578 291600 75198
rect 293600 75038 293900 75039
rect 293600 74737 293900 74738
rect 0 73398 292000 74578
rect -998 73238 -698 73239
rect -998 72937 -698 72938
rect 400 72778 291600 73398
rect 292660 73238 292960 73239
rect 292660 72937 292960 72938
rect 0 69798 292000 72778
rect -4288 69638 -3988 69639
rect -4288 69337 -3988 69338
rect 400 69178 291600 69798
rect 295950 69638 296250 69639
rect 295950 69337 296250 69338
rect 0 67998 292000 69178
rect -3348 67838 -3048 67839
rect -3348 67537 -3048 67538
rect 400 67378 291600 67998
rect 295010 67838 295310 67839
rect 295010 67537 295310 67538
rect 0 66198 292000 67378
rect -2408 66038 -2108 66039
rect -2408 65737 -2108 65738
rect 400 65578 291600 66198
rect 294070 66038 294370 66039
rect 294070 65737 294370 65738
rect 0 64398 292000 65578
rect -1468 64238 -1168 64239
rect -1468 63937 -1168 63938
rect 400 63778 291600 64398
rect 293130 64238 293430 64239
rect 293130 63937 293430 63938
rect 0 60798 292000 63778
rect -3818 60638 -3518 60639
rect -3818 60337 -3518 60338
rect 400 60178 291600 60798
rect 295480 60638 295780 60639
rect 295480 60337 295780 60338
rect 0 58998 292000 60178
rect -2878 58838 -2578 58839
rect -2878 58537 -2578 58538
rect 400 58378 291600 58998
rect 294540 58838 294840 58839
rect 294540 58537 294840 58538
rect 0 57198 292000 58378
rect -1938 57038 -1638 57039
rect -1938 56737 -1638 56738
rect 400 56578 291600 57198
rect 293600 57038 293900 57039
rect 293600 56737 293900 56738
rect 0 55398 292000 56578
rect -998 55238 -698 55239
rect -998 54937 -698 54938
rect 400 54778 291600 55398
rect 292660 55238 292960 55239
rect 292660 54937 292960 54938
rect 0 51798 292000 54778
rect -4288 51638 -3988 51639
rect -4288 51337 -3988 51338
rect 400 51178 291600 51798
rect 295950 51638 296250 51639
rect 295950 51337 296250 51338
rect 0 49998 292000 51178
rect -3348 49838 -3048 49839
rect -3348 49537 -3048 49538
rect 400 49378 291600 49998
rect 295010 49838 295310 49839
rect 295010 49537 295310 49538
rect 0 48198 292000 49378
rect -2408 48038 -2108 48039
rect -2408 47737 -2108 47738
rect 400 47578 291600 48198
rect 294070 48038 294370 48039
rect 294070 47737 294370 47738
rect 0 46398 292000 47578
rect -1468 46238 -1168 46239
rect -1468 45937 -1168 45938
rect 400 45778 291600 46398
rect 293130 46238 293430 46239
rect 293130 45937 293430 45938
rect 0 42798 292000 45778
rect -3818 42638 -3518 42639
rect -3818 42337 -3518 42338
rect 400 42178 291600 42798
rect 295480 42638 295780 42639
rect 295480 42337 295780 42338
rect 0 40998 292000 42178
rect -2878 40838 -2578 40839
rect -2878 40537 -2578 40538
rect 400 40378 291600 40998
rect 294540 40838 294840 40839
rect 294540 40537 294840 40538
rect 0 39198 292000 40378
rect -1938 39038 -1638 39039
rect -1938 38737 -1638 38738
rect 400 38578 291600 39198
rect 293600 39038 293900 39039
rect 293600 38737 293900 38738
rect 0 37398 292000 38578
rect -998 37238 -698 37239
rect -998 36937 -698 36938
rect 400 36778 291600 37398
rect 292660 37238 292960 37239
rect 292660 36937 292960 36938
rect 0 33798 292000 36778
rect -4288 33638 -3988 33639
rect -4288 33337 -3988 33338
rect 400 33178 291600 33798
rect 295950 33638 296250 33639
rect 295950 33337 296250 33338
rect 0 31998 292000 33178
rect -3348 31838 -3048 31839
rect -3348 31537 -3048 31538
rect 400 31378 291600 31998
rect 295010 31838 295310 31839
rect 295010 31537 295310 31538
rect 0 30198 292000 31378
rect -2408 30038 -2108 30039
rect -2408 29737 -2108 29738
rect 400 29578 291600 30198
rect 294070 30038 294370 30039
rect 294070 29737 294370 29738
rect 0 28398 292000 29578
rect -1468 28238 -1168 28239
rect -1468 27937 -1168 27938
rect 400 27778 291600 28398
rect 293130 28238 293430 28239
rect 293130 27937 293430 27938
rect 0 24798 292000 27778
rect -3818 24638 -3518 24639
rect -3818 24337 -3518 24338
rect 400 24178 291600 24798
rect 295480 24638 295780 24639
rect 295480 24337 295780 24338
rect 0 22998 292000 24178
rect -2878 22838 -2578 22839
rect -2878 22537 -2578 22538
rect 400 22378 291600 22998
rect 294540 22838 294840 22839
rect 294540 22537 294840 22538
rect 0 21198 292000 22378
rect -1938 21038 -1638 21039
rect -1938 20737 -1638 20738
rect 400 20578 291600 21198
rect 293600 21038 293900 21039
rect 293600 20737 293900 20738
rect 0 19398 292000 20578
rect -998 19238 -698 19239
rect -998 18937 -698 18938
rect 400 18778 291600 19398
rect 292660 19238 292960 19239
rect 292660 18937 292960 18938
rect 0 15798 292000 18778
rect -4288 15638 -3988 15639
rect -4288 15337 -3988 15338
rect 400 15178 291600 15798
rect 295950 15638 296250 15639
rect 295950 15337 296250 15338
rect 0 13998 292000 15178
rect -3348 13838 -3048 13839
rect -3348 13537 -3048 13538
rect 400 13378 291600 13998
rect 295010 13838 295310 13839
rect 295010 13537 295310 13538
rect 0 12198 292000 13378
rect -2408 12038 -2108 12039
rect -2408 11737 -2108 11738
rect 400 11578 291600 12198
rect 294070 12038 294370 12039
rect 294070 11737 294370 11738
rect 0 10398 292000 11578
rect -1468 10238 -1168 10239
rect -1468 9937 -1168 9938
rect 400 9778 291600 10398
rect 293130 10238 293430 10239
rect 293130 9937 293430 9938
rect 0 6798 292000 9778
rect -3818 6638 -3518 6639
rect -3818 6337 -3518 6338
rect 400 6178 291600 6798
rect 295480 6638 295780 6639
rect 295480 6337 295780 6338
rect 0 4998 292000 6178
rect -2878 4838 -2578 4839
rect -2878 4537 -2578 4538
rect 400 4378 291600 4998
rect 294540 4838 294840 4839
rect 294540 4537 294840 4538
rect 0 3198 292000 4378
rect -1938 3038 -1638 3039
rect -1938 2737 -1638 2738
rect 400 2578 291600 3198
rect 293600 3038 293900 3039
rect 293600 2737 293900 2738
rect 0 1398 292000 2578
rect -998 1238 -698 1239
rect -998 937 -698 938
rect 400 778 291600 1398
rect 292660 1238 292960 1239
rect 292660 937 292960 938
rect 0 0 292000 778
rect -998 -162 -698 -161
rect 402 -162 702 -161
rect 18402 -162 18702 -161
rect 36402 -162 36702 -161
rect 54402 -162 54702 -161
rect 72402 -162 72702 -161
rect 90402 -162 90702 -161
rect 108402 -162 108702 -161
rect 126402 -162 126702 -161
rect 144402 -162 144702 -161
rect 162402 -162 162702 -161
rect 180402 -162 180702 -161
rect 198402 -162 198702 -161
rect 216402 -162 216702 -161
rect 234402 -162 234702 -161
rect 252402 -162 252702 -161
rect 270402 -162 270702 -161
rect 288402 -162 288702 -161
rect 292660 -162 292960 -161
rect -998 -463 -698 -462
rect 402 -463 702 -462
rect 18402 -463 18702 -462
rect 36402 -463 36702 -462
rect 54402 -463 54702 -462
rect 72402 -463 72702 -462
rect 90402 -463 90702 -462
rect 108402 -463 108702 -462
rect 126402 -463 126702 -462
rect 144402 -463 144702 -462
rect 162402 -463 162702 -462
rect 180402 -463 180702 -462
rect 198402 -463 198702 -462
rect 216402 -463 216702 -462
rect 234402 -463 234702 -462
rect 252402 -463 252702 -462
rect 270402 -463 270702 -462
rect 288402 -463 288702 -462
rect 292660 -463 292960 -462
rect -1468 -632 -1168 -631
rect 9402 -632 9702 -631
rect 27402 -632 27702 -631
rect 45402 -632 45702 -631
rect 63402 -632 63702 -631
rect 81402 -632 81702 -631
rect 99402 -632 99702 -631
rect 117402 -632 117702 -631
rect 135402 -632 135702 -631
rect 153402 -632 153702 -631
rect 171402 -632 171702 -631
rect 189402 -632 189702 -631
rect 207402 -632 207702 -631
rect 225402 -632 225702 -631
rect 243402 -632 243702 -631
rect 261402 -632 261702 -631
rect 279402 -632 279702 -631
rect 293130 -632 293430 -631
rect -1468 -933 -1168 -932
rect 9402 -933 9702 -932
rect 27402 -933 27702 -932
rect 45402 -933 45702 -932
rect 63402 -933 63702 -932
rect 81402 -933 81702 -932
rect 99402 -933 99702 -932
rect 117402 -933 117702 -932
rect 135402 -933 135702 -932
rect 153402 -933 153702 -932
rect 171402 -933 171702 -932
rect 189402 -933 189702 -932
rect 207402 -933 207702 -932
rect 225402 -933 225702 -932
rect 243402 -933 243702 -932
rect 261402 -933 261702 -932
rect 279402 -933 279702 -932
rect 293130 -933 293430 -932
rect -1938 -1102 -1638 -1101
rect 2202 -1102 2502 -1101
rect 20202 -1102 20502 -1101
rect 38202 -1102 38502 -1101
rect 56202 -1102 56502 -1101
rect 74202 -1102 74502 -1101
rect 92202 -1102 92502 -1101
rect 110202 -1102 110502 -1101
rect 128202 -1102 128502 -1101
rect 146202 -1102 146502 -1101
rect 164202 -1102 164502 -1101
rect 182202 -1102 182502 -1101
rect 200202 -1102 200502 -1101
rect 218202 -1102 218502 -1101
rect 236202 -1102 236502 -1101
rect 254202 -1102 254502 -1101
rect 272202 -1102 272502 -1101
rect 290202 -1102 290502 -1101
rect 293600 -1102 293900 -1101
rect -1938 -1403 -1638 -1402
rect 2202 -1403 2502 -1402
rect 20202 -1403 20502 -1402
rect 38202 -1403 38502 -1402
rect 56202 -1403 56502 -1402
rect 74202 -1403 74502 -1402
rect 92202 -1403 92502 -1402
rect 110202 -1403 110502 -1402
rect 128202 -1403 128502 -1402
rect 146202 -1403 146502 -1402
rect 164202 -1403 164502 -1402
rect 182202 -1403 182502 -1402
rect 200202 -1403 200502 -1402
rect 218202 -1403 218502 -1402
rect 236202 -1403 236502 -1402
rect 254202 -1403 254502 -1402
rect 272202 -1403 272502 -1402
rect 290202 -1403 290502 -1402
rect 293600 -1403 293900 -1402
rect -2408 -1572 -2108 -1571
rect 11202 -1572 11502 -1571
rect 29202 -1572 29502 -1571
rect 47202 -1572 47502 -1571
rect 65202 -1572 65502 -1571
rect 83202 -1572 83502 -1571
rect 101202 -1572 101502 -1571
rect 119202 -1572 119502 -1571
rect 137202 -1572 137502 -1571
rect 155202 -1572 155502 -1571
rect 173202 -1572 173502 -1571
rect 191202 -1572 191502 -1571
rect 209202 -1572 209502 -1571
rect 227202 -1572 227502 -1571
rect 245202 -1572 245502 -1571
rect 263202 -1572 263502 -1571
rect 281202 -1572 281502 -1571
rect 294070 -1572 294370 -1571
rect -2408 -1873 -2108 -1872
rect 11202 -1873 11502 -1872
rect 29202 -1873 29502 -1872
rect 47202 -1873 47502 -1872
rect 65202 -1873 65502 -1872
rect 83202 -1873 83502 -1872
rect 101202 -1873 101502 -1872
rect 119202 -1873 119502 -1872
rect 137202 -1873 137502 -1872
rect 155202 -1873 155502 -1872
rect 173202 -1873 173502 -1872
rect 191202 -1873 191502 -1872
rect 209202 -1873 209502 -1872
rect 227202 -1873 227502 -1872
rect 245202 -1873 245502 -1872
rect 263202 -1873 263502 -1872
rect 281202 -1873 281502 -1872
rect 294070 -1873 294370 -1872
rect -2878 -2042 -2578 -2041
rect 4002 -2042 4302 -2041
rect 22002 -2042 22302 -2041
rect 40002 -2042 40302 -2041
rect 58002 -2042 58302 -2041
rect 76002 -2042 76302 -2041
rect 94002 -2042 94302 -2041
rect 112002 -2042 112302 -2041
rect 130002 -2042 130302 -2041
rect 148002 -2042 148302 -2041
rect 166002 -2042 166302 -2041
rect 184002 -2042 184302 -2041
rect 202002 -2042 202302 -2041
rect 220002 -2042 220302 -2041
rect 238002 -2042 238302 -2041
rect 256002 -2042 256302 -2041
rect 274002 -2042 274302 -2041
rect 294540 -2042 294840 -2041
rect -2878 -2343 -2578 -2342
rect 4002 -2343 4302 -2342
rect 22002 -2343 22302 -2342
rect 40002 -2343 40302 -2342
rect 58002 -2343 58302 -2342
rect 76002 -2343 76302 -2342
rect 94002 -2343 94302 -2342
rect 112002 -2343 112302 -2342
rect 130002 -2343 130302 -2342
rect 148002 -2343 148302 -2342
rect 166002 -2343 166302 -2342
rect 184002 -2343 184302 -2342
rect 202002 -2343 202302 -2342
rect 220002 -2343 220302 -2342
rect 238002 -2343 238302 -2342
rect 256002 -2343 256302 -2342
rect 274002 -2343 274302 -2342
rect 294540 -2343 294840 -2342
rect -3348 -2512 -3048 -2511
rect 13002 -2512 13302 -2511
rect 31002 -2512 31302 -2511
rect 49002 -2512 49302 -2511
rect 67002 -2512 67302 -2511
rect 85002 -2512 85302 -2511
rect 103002 -2512 103302 -2511
rect 121002 -2512 121302 -2511
rect 139002 -2512 139302 -2511
rect 157002 -2512 157302 -2511
rect 175002 -2512 175302 -2511
rect 193002 -2512 193302 -2511
rect 211002 -2512 211302 -2511
rect 229002 -2512 229302 -2511
rect 247002 -2512 247302 -2511
rect 265002 -2512 265302 -2511
rect 283002 -2512 283302 -2511
rect 295010 -2512 295310 -2511
rect -3348 -2813 -3048 -2812
rect 13002 -2813 13302 -2812
rect 31002 -2813 31302 -2812
rect 49002 -2813 49302 -2812
rect 67002 -2813 67302 -2812
rect 85002 -2813 85302 -2812
rect 103002 -2813 103302 -2812
rect 121002 -2813 121302 -2812
rect 139002 -2813 139302 -2812
rect 157002 -2813 157302 -2812
rect 175002 -2813 175302 -2812
rect 193002 -2813 193302 -2812
rect 211002 -2813 211302 -2812
rect 229002 -2813 229302 -2812
rect 247002 -2813 247302 -2812
rect 265002 -2813 265302 -2812
rect 283002 -2813 283302 -2812
rect 295010 -2813 295310 -2812
rect -3818 -2982 -3518 -2981
rect 5802 -2982 6102 -2981
rect 23802 -2982 24102 -2981
rect 41802 -2982 42102 -2981
rect 59802 -2982 60102 -2981
rect 77802 -2982 78102 -2981
rect 95802 -2982 96102 -2981
rect 113802 -2982 114102 -2981
rect 131802 -2982 132102 -2981
rect 149802 -2982 150102 -2981
rect 167802 -2982 168102 -2981
rect 185802 -2982 186102 -2981
rect 203802 -2982 204102 -2981
rect 221802 -2982 222102 -2981
rect 239802 -2982 240102 -2981
rect 257802 -2982 258102 -2981
rect 275802 -2982 276102 -2981
rect 295480 -2982 295780 -2981
rect -3818 -3283 -3518 -3282
rect 5802 -3283 6102 -3282
rect 23802 -3283 24102 -3282
rect 41802 -3283 42102 -3282
rect 59802 -3283 60102 -3282
rect 77802 -3283 78102 -3282
rect 95802 -3283 96102 -3282
rect 113802 -3283 114102 -3282
rect 131802 -3283 132102 -3282
rect 149802 -3283 150102 -3282
rect 167802 -3283 168102 -3282
rect 185802 -3283 186102 -3282
rect 203802 -3283 204102 -3282
rect 221802 -3283 222102 -3282
rect 239802 -3283 240102 -3282
rect 257802 -3283 258102 -3282
rect 275802 -3283 276102 -3282
rect 295480 -3283 295780 -3282
rect -4288 -3452 -3988 -3451
rect 14802 -3452 15102 -3451
rect 32802 -3452 33102 -3451
rect 50802 -3452 51102 -3451
rect 68802 -3452 69102 -3451
rect 86802 -3452 87102 -3451
rect 104802 -3452 105102 -3451
rect 122802 -3452 123102 -3451
rect 140802 -3452 141102 -3451
rect 158802 -3452 159102 -3451
rect 176802 -3452 177102 -3451
rect 194802 -3452 195102 -3451
rect 212802 -3452 213102 -3451
rect 230802 -3452 231102 -3451
rect 248802 -3452 249102 -3451
rect 266802 -3452 267102 -3451
rect 284802 -3452 285102 -3451
rect 295950 -3452 296250 -3451
rect -4288 -3753 -3988 -3752
rect 14802 -3753 15102 -3752
rect 32802 -3753 33102 -3752
rect 50802 -3753 51102 -3752
rect 68802 -3753 69102 -3752
rect 86802 -3753 87102 -3752
rect 104802 -3753 105102 -3752
rect 122802 -3753 123102 -3752
rect 140802 -3753 141102 -3752
rect 158802 -3753 159102 -3752
rect 176802 -3753 177102 -3752
rect 194802 -3753 195102 -3752
rect 212802 -3753 213102 -3752
rect 230802 -3753 231102 -3752
rect 248802 -3753 249102 -3752
rect 266802 -3753 267102 -3752
rect 284802 -3753 285102 -3752
rect 295950 -3753 296250 -3752
<< labels >>
rlabel metal3 s 291760 2898 292480 3018 6 analog_io[0]
port 1 nsew default bidirectional
rlabel metal3 s 291760 237498 292480 237618 6 analog_io[10]
port 2 nsew default bidirectional
rlabel metal3 s 291760 260958 292480 261078 6 analog_io[11]
port 3 nsew default bidirectional
rlabel metal3 s 291760 284418 292480 284538 6 analog_io[12]
port 4 nsew default bidirectional
rlabel metal3 s 291760 307878 292480 307998 6 analog_io[13]
port 5 nsew default bidirectional
rlabel metal3 s 291760 331338 292480 331458 6 analog_io[14]
port 6 nsew default bidirectional
rlabel metal2 s 287909 351760 287965 352480 6 analog_io[15]
port 7 nsew default bidirectional
rlabel metal2 s 255479 351760 255535 352480 6 analog_io[16]
port 8 nsew default bidirectional
rlabel metal2 s 223049 351760 223105 352480 6 analog_io[17]
port 9 nsew default bidirectional
rlabel metal2 s 190573 351760 190629 352480 6 analog_io[18]
port 10 nsew default bidirectional
rlabel metal2 s 158143 351760 158199 352480 6 analog_io[19]
port 11 nsew default bidirectional
rlabel metal3 s 291760 26358 292480 26478 6 analog_io[1]
port 12 nsew default bidirectional
rlabel metal2 s 125713 351760 125769 352480 6 analog_io[20]
port 13 nsew default bidirectional
rlabel metal2 s 93237 351760 93293 352480 6 analog_io[21]
port 14 nsew default bidirectional
rlabel metal2 s 60807 351760 60863 352480 6 analog_io[22]
port 15 nsew default bidirectional
rlabel metal2 s 28377 351760 28433 352480 6 analog_io[23]
port 16 nsew default bidirectional
rlabel metal3 s -480 348270 240 348390 4 analog_io[24]
port 17 nsew default bidirectional
rlabel metal3 s -480 319506 240 319626 4 analog_io[25]
port 18 nsew default bidirectional
rlabel metal3 s -480 290810 240 290930 4 analog_io[26]
port 19 nsew default bidirectional
rlabel metal3 s -480 262046 240 262166 4 analog_io[27]
port 20 nsew default bidirectional
rlabel metal3 s -480 233350 240 233470 4 analog_io[28]
port 21 nsew default bidirectional
rlabel metal3 s -480 204586 240 204706 4 analog_io[29]
port 22 nsew default bidirectional
rlabel metal3 s 291760 49818 292480 49938 6 analog_io[2]
port 23 nsew default bidirectional
rlabel metal3 s -480 175890 240 176010 4 analog_io[30]
port 24 nsew default bidirectional
rlabel metal3 s 291760 73278 292480 73398 6 analog_io[3]
port 25 nsew default bidirectional
rlabel metal3 s 291760 96738 292480 96858 6 analog_io[4]
port 26 nsew default bidirectional
rlabel metal3 s 291760 120198 292480 120318 6 analog_io[5]
port 27 nsew default bidirectional
rlabel metal3 s 291760 143658 292480 143778 6 analog_io[6]
port 28 nsew default bidirectional
rlabel metal3 s 291760 167118 292480 167238 6 analog_io[7]
port 29 nsew default bidirectional
rlabel metal3 s 291760 190578 292480 190698 6 analog_io[8]
port 30 nsew default bidirectional
rlabel metal3 s 291760 214038 292480 214158 6 analog_io[9]
port 31 nsew default bidirectional
rlabel metal3 s 291760 8746 292480 8866 6 io_in[0]
port 32 nsew default input
rlabel metal3 s 291760 243346 292480 243466 6 io_in[10]
port 33 nsew default input
rlabel metal3 s 291760 266874 292480 266994 6 io_in[11]
port 34 nsew default input
rlabel metal3 s 291760 290334 292480 290454 6 io_in[12]
port 35 nsew default input
rlabel metal3 s 291760 313794 292480 313914 6 io_in[13]
port 36 nsew default input
rlabel metal3 s 291760 337254 292480 337374 6 io_in[14]
port 37 nsew default input
rlabel metal2 s 279813 351760 279869 352480 6 io_in[15]
port 38 nsew default input
rlabel metal2 s 247383 351760 247439 352480 6 io_in[16]
port 39 nsew default input
rlabel metal2 s 214907 351760 214963 352480 6 io_in[17]
port 40 nsew default input
rlabel metal2 s 182477 351760 182533 352480 6 io_in[18]
port 41 nsew default input
rlabel metal2 s 150047 351760 150103 352480 6 io_in[19]
port 42 nsew default input
rlabel metal3 s 291760 32206 292480 32326 6 io_in[1]
port 43 nsew default input
rlabel metal2 s 117571 351760 117627 352480 6 io_in[20]
port 44 nsew default input
rlabel metal2 s 85141 351760 85197 352480 6 io_in[21]
port 45 nsew default input
rlabel metal2 s 52711 351760 52767 352480 6 io_in[22]
port 46 nsew default input
rlabel metal2 s 20235 351760 20291 352480 6 io_in[23]
port 47 nsew default input
rlabel metal3 s -480 341062 240 341182 4 io_in[24]
port 48 nsew default input
rlabel metal3 s -480 312366 240 312486 4 io_in[25]
port 49 nsew default input
rlabel metal3 s -480 283602 240 283722 4 io_in[26]
port 50 nsew default input
rlabel metal3 s -480 254906 240 255026 4 io_in[27]
port 51 nsew default input
rlabel metal3 s -480 226142 240 226262 4 io_in[28]
port 52 nsew default input
rlabel metal3 s -480 197446 240 197566 4 io_in[29]
port 53 nsew default input
rlabel metal3 s 291760 55666 292480 55786 6 io_in[2]
port 54 nsew default input
rlabel metal3 s -480 168682 240 168802 4 io_in[30]
port 55 nsew default input
rlabel metal3 s -480 147126 240 147246 4 io_in[31]
port 56 nsew default input
rlabel metal3 s -480 125570 240 125690 4 io_in[32]
port 57 nsew default input
rlabel metal3 s -480 104014 240 104134 4 io_in[33]
port 58 nsew default input
rlabel metal3 s -480 82458 240 82578 4 io_in[34]
port 59 nsew default input
rlabel metal3 s -480 60970 240 61090 4 io_in[35]
port 60 nsew default input
rlabel metal3 s -480 39414 240 39534 4 io_in[36]
port 61 nsew default input
rlabel metal3 s -480 17858 240 17978 4 io_in[37]
port 62 nsew default input
rlabel metal3 s 291760 79126 292480 79246 6 io_in[3]
port 63 nsew default input
rlabel metal3 s 291760 102586 292480 102706 6 io_in[4]
port 64 nsew default input
rlabel metal3 s 291760 126046 292480 126166 6 io_in[5]
port 65 nsew default input
rlabel metal3 s 291760 149506 292480 149626 6 io_in[6]
port 66 nsew default input
rlabel metal3 s 291760 172966 292480 173086 6 io_in[7]
port 67 nsew default input
rlabel metal3 s 291760 196426 292480 196546 6 io_in[8]
port 68 nsew default input
rlabel metal3 s 291760 219886 292480 220006 6 io_in[9]
port 69 nsew default input
rlabel metal3 s 291760 20442 292480 20562 6 io_oeb[0]
port 70 nsew default output
rlabel metal3 s 291760 255110 292480 255230 6 io_oeb[10]
port 71 nsew default output
rlabel metal3 s 291760 278570 292480 278690 6 io_oeb[11]
port 72 nsew default output
rlabel metal3 s 291760 302030 292480 302150 6 io_oeb[12]
port 73 nsew default output
rlabel metal3 s 291760 325490 292480 325610 6 io_oeb[13]
port 74 nsew default output
rlabel metal3 s 291760 348950 292480 349070 6 io_oeb[14]
port 75 nsew default output
rlabel metal2 s 263575 351760 263631 352480 6 io_oeb[15]
port 76 nsew default output
rlabel metal2 s 231145 351760 231201 352480 6 io_oeb[16]
port 77 nsew default output
rlabel metal2 s 198715 351760 198771 352480 6 io_oeb[17]
port 78 nsew default output
rlabel metal2 s 166239 351760 166295 352480 6 io_oeb[18]
port 79 nsew default output
rlabel metal2 s 133809 351760 133865 352480 6 io_oeb[19]
port 80 nsew default output
rlabel metal3 s 291760 43902 292480 44022 6 io_oeb[1]
port 81 nsew default output
rlabel metal2 s 101379 351760 101435 352480 6 io_oeb[20]
port 82 nsew default output
rlabel metal2 s 68903 351760 68959 352480 6 io_oeb[21]
port 83 nsew default output
rlabel metal2 s 36473 351760 36529 352480 6 io_oeb[22]
port 84 nsew default output
rlabel metal2 s 4043 351760 4099 352480 6 io_oeb[23]
port 85 nsew default output
rlabel metal3 s -480 326714 240 326834 4 io_oeb[24]
port 86 nsew default output
rlabel metal3 s -480 297950 240 298070 4 io_oeb[25]
port 87 nsew default output
rlabel metal3 s -480 269254 240 269374 4 io_oeb[26]
port 88 nsew default output
rlabel metal3 s -480 240490 240 240610 4 io_oeb[27]
port 89 nsew default output
rlabel metal3 s -480 211794 240 211914 4 io_oeb[28]
port 90 nsew default output
rlabel metal3 s -480 183030 240 183150 4 io_oeb[29]
port 91 nsew default output
rlabel metal3 s 291760 67362 292480 67482 6 io_oeb[2]
port 92 nsew default output
rlabel metal3 s -480 154334 240 154454 4 io_oeb[30]
port 93 nsew default output
rlabel metal3 s -480 132778 240 132898 4 io_oeb[31]
port 94 nsew default output
rlabel metal3 s -480 111222 240 111342 4 io_oeb[32]
port 95 nsew default output
rlabel metal3 s -480 89666 240 89786 4 io_oeb[33]
port 96 nsew default output
rlabel metal3 s -480 68110 240 68230 4 io_oeb[34]
port 97 nsew default output
rlabel metal3 s -480 46554 240 46674 4 io_oeb[35]
port 98 nsew default output
rlabel metal3 s -480 24998 240 25118 4 io_oeb[36]
port 99 nsew default output
rlabel metal3 s -480 3510 240 3630 4 io_oeb[37]
port 100 nsew default output
rlabel metal3 s 291760 90890 292480 91010 6 io_oeb[3]
port 101 nsew default output
rlabel metal3 s 291760 114350 292480 114470 6 io_oeb[4]
port 102 nsew default output
rlabel metal3 s 291760 137810 292480 137930 6 io_oeb[5]
port 103 nsew default output
rlabel metal3 s 291760 161270 292480 161390 6 io_oeb[6]
port 104 nsew default output
rlabel metal3 s 291760 184730 292480 184850 6 io_oeb[7]
port 105 nsew default output
rlabel metal3 s 291760 208190 292480 208310 6 io_oeb[8]
port 106 nsew default output
rlabel metal3 s 291760 231650 292480 231770 6 io_oeb[9]
port 107 nsew default output
rlabel metal3 s 291760 14594 292480 14714 6 io_out[0]
port 108 nsew default output
rlabel metal3 s 291760 249262 292480 249382 6 io_out[10]
port 109 nsew default output
rlabel metal3 s 291760 272722 292480 272842 6 io_out[11]
port 110 nsew default output
rlabel metal3 s 291760 296182 292480 296302 6 io_out[12]
port 111 nsew default output
rlabel metal3 s 291760 319642 292480 319762 6 io_out[13]
port 112 nsew default output
rlabel metal3 s 291760 343102 292480 343222 6 io_out[14]
port 113 nsew default output
rlabel metal2 s 271717 351760 271773 352480 6 io_out[15]
port 114 nsew default output
rlabel metal2 s 239241 351760 239297 352480 6 io_out[16]
port 115 nsew default output
rlabel metal2 s 206811 351760 206867 352480 6 io_out[17]
port 116 nsew default output
rlabel metal2 s 174381 351760 174437 352480 6 io_out[18]
port 117 nsew default output
rlabel metal2 s 141905 351760 141961 352480 6 io_out[19]
port 118 nsew default output
rlabel metal3 s 291760 38054 292480 38174 6 io_out[1]
port 119 nsew default output
rlabel metal2 s 109475 351760 109531 352480 6 io_out[20]
port 120 nsew default output
rlabel metal2 s 77045 351760 77101 352480 6 io_out[21]
port 121 nsew default output
rlabel metal2 s 44569 351760 44625 352480 6 io_out[22]
port 122 nsew default output
rlabel metal2 s 12139 351760 12195 352480 6 io_out[23]
port 123 nsew default output
rlabel metal3 s -480 333922 240 334042 4 io_out[24]
port 124 nsew default output
rlabel metal3 s -480 305158 240 305278 4 io_out[25]
port 125 nsew default output
rlabel metal3 s -480 276462 240 276582 4 io_out[26]
port 126 nsew default output
rlabel metal3 s -480 247698 240 247818 4 io_out[27]
port 127 nsew default output
rlabel metal3 s -480 218934 240 219054 4 io_out[28]
port 128 nsew default output
rlabel metal3 s -480 190238 240 190358 4 io_out[29]
port 129 nsew default output
rlabel metal3 s 291760 61514 292480 61634 6 io_out[2]
port 130 nsew default output
rlabel metal3 s -480 161474 240 161594 4 io_out[30]
port 131 nsew default output
rlabel metal3 s -480 139986 240 140106 4 io_out[31]
port 132 nsew default output
rlabel metal3 s -480 118430 240 118550 4 io_out[32]
port 133 nsew default output
rlabel metal3 s -480 96874 240 96994 4 io_out[33]
port 134 nsew default output
rlabel metal3 s -480 75318 240 75438 4 io_out[34]
port 135 nsew default output
rlabel metal3 s -480 53762 240 53882 4 io_out[35]
port 136 nsew default output
rlabel metal3 s -480 32206 240 32326 4 io_out[36]
port 137 nsew default output
rlabel metal3 s -480 10650 240 10770 4 io_out[37]
port 138 nsew default output
rlabel metal3 s 291760 84974 292480 85094 6 io_out[3]
port 139 nsew default output
rlabel metal3 s 291760 108434 292480 108554 6 io_out[4]
port 140 nsew default output
rlabel metal3 s 291760 131894 292480 132014 6 io_out[5]
port 141 nsew default output
rlabel metal3 s 291760 155354 292480 155474 6 io_out[6]
port 142 nsew default output
rlabel metal3 s 291760 178882 292480 179002 6 io_out[7]
port 143 nsew default output
rlabel metal3 s 291760 202342 292480 202462 6 io_out[8]
port 144 nsew default output
rlabel metal3 s 291760 225802 292480 225922 6 io_out[9]
port 145 nsew default output
rlabel metal2 s 63291 -480 63347 240 8 la_data_in[0]
port 146 nsew default input
rlabel metal2 s 241725 -480 241781 240 8 la_data_in[100]
port 147 nsew default input
rlabel metal2 s 243473 -480 243529 240 8 la_data_in[101]
port 148 nsew default input
rlabel metal2 s 245267 -480 245323 240 8 la_data_in[102]
port 149 nsew default input
rlabel metal2 s 247061 -480 247117 240 8 la_data_in[103]
port 150 nsew default input
rlabel metal2 s 248855 -480 248911 240 8 la_data_in[104]
port 151 nsew default input
rlabel metal2 s 250603 -480 250659 240 8 la_data_in[105]
port 152 nsew default input
rlabel metal2 s 252397 -480 252453 240 8 la_data_in[106]
port 153 nsew default input
rlabel metal2 s 254191 -480 254247 240 8 la_data_in[107]
port 154 nsew default input
rlabel metal2 s 255985 -480 256041 240 8 la_data_in[108]
port 155 nsew default input
rlabel metal2 s 257779 -480 257835 240 8 la_data_in[109]
port 156 nsew default input
rlabel metal2 s 81139 -480 81195 240 8 la_data_in[10]
port 157 nsew default input
rlabel metal2 s 259527 -480 259583 240 8 la_data_in[110]
port 158 nsew default input
rlabel metal2 s 261321 -480 261377 240 8 la_data_in[111]
port 159 nsew default input
rlabel metal2 s 263115 -480 263171 240 8 la_data_in[112]
port 160 nsew default input
rlabel metal2 s 264909 -480 264965 240 8 la_data_in[113]
port 161 nsew default input
rlabel metal2 s 266703 -480 266759 240 8 la_data_in[114]
port 162 nsew default input
rlabel metal2 s 268451 -480 268507 240 8 la_data_in[115]
port 163 nsew default input
rlabel metal2 s 270245 -480 270301 240 8 la_data_in[116]
port 164 nsew default input
rlabel metal2 s 272039 -480 272095 240 8 la_data_in[117]
port 165 nsew default input
rlabel metal2 s 273833 -480 273889 240 8 la_data_in[118]
port 166 nsew default input
rlabel metal2 s 275581 -480 275637 240 8 la_data_in[119]
port 167 nsew default input
rlabel metal2 s 82933 -480 82989 240 8 la_data_in[11]
port 168 nsew default input
rlabel metal2 s 277375 -480 277431 240 8 la_data_in[120]
port 169 nsew default input
rlabel metal2 s 279169 -480 279225 240 8 la_data_in[121]
port 170 nsew default input
rlabel metal2 s 280963 -480 281019 240 8 la_data_in[122]
port 171 nsew default input
rlabel metal2 s 282757 -480 282813 240 8 la_data_in[123]
port 172 nsew default input
rlabel metal2 s 284505 -480 284561 240 8 la_data_in[124]
port 173 nsew default input
rlabel metal2 s 286299 -480 286355 240 8 la_data_in[125]
port 174 nsew default input
rlabel metal2 s 288093 -480 288149 240 8 la_data_in[126]
port 175 nsew default input
rlabel metal2 s 289887 -480 289943 240 8 la_data_in[127]
port 176 nsew default input
rlabel metal2 s 84681 -480 84737 240 8 la_data_in[12]
port 177 nsew default input
rlabel metal2 s 86475 -480 86531 240 8 la_data_in[13]
port 178 nsew default input
rlabel metal2 s 88269 -480 88325 240 8 la_data_in[14]
port 179 nsew default input
rlabel metal2 s 90063 -480 90119 240 8 la_data_in[15]
port 180 nsew default input
rlabel metal2 s 91857 -480 91913 240 8 la_data_in[16]
port 181 nsew default input
rlabel metal2 s 93605 -480 93661 240 8 la_data_in[17]
port 182 nsew default input
rlabel metal2 s 95399 -480 95455 240 8 la_data_in[18]
port 183 nsew default input
rlabel metal2 s 97193 -480 97249 240 8 la_data_in[19]
port 184 nsew default input
rlabel metal2 s 65085 -480 65141 240 8 la_data_in[1]
port 185 nsew default input
rlabel metal2 s 98987 -480 99043 240 8 la_data_in[20]
port 186 nsew default input
rlabel metal2 s 100735 -480 100791 240 8 la_data_in[21]
port 187 nsew default input
rlabel metal2 s 102529 -480 102585 240 8 la_data_in[22]
port 188 nsew default input
rlabel metal2 s 104323 -480 104379 240 8 la_data_in[23]
port 189 nsew default input
rlabel metal2 s 106117 -480 106173 240 8 la_data_in[24]
port 190 nsew default input
rlabel metal2 s 107911 -480 107967 240 8 la_data_in[25]
port 191 nsew default input
rlabel metal2 s 109659 -480 109715 240 8 la_data_in[26]
port 192 nsew default input
rlabel metal2 s 111453 -480 111509 240 8 la_data_in[27]
port 193 nsew default input
rlabel metal2 s 113247 -480 113303 240 8 la_data_in[28]
port 194 nsew default input
rlabel metal2 s 115041 -480 115097 240 8 la_data_in[29]
port 195 nsew default input
rlabel metal2 s 66879 -480 66935 240 8 la_data_in[2]
port 196 nsew default input
rlabel metal2 s 116835 -480 116891 240 8 la_data_in[30]
port 197 nsew default input
rlabel metal2 s 118583 -480 118639 240 8 la_data_in[31]
port 198 nsew default input
rlabel metal2 s 120377 -480 120433 240 8 la_data_in[32]
port 199 nsew default input
rlabel metal2 s 122171 -480 122227 240 8 la_data_in[33]
port 200 nsew default input
rlabel metal2 s 123965 -480 124021 240 8 la_data_in[34]
port 201 nsew default input
rlabel metal2 s 125713 -480 125769 240 8 la_data_in[35]
port 202 nsew default input
rlabel metal2 s 127507 -480 127563 240 8 la_data_in[36]
port 203 nsew default input
rlabel metal2 s 129301 -480 129357 240 8 la_data_in[37]
port 204 nsew default input
rlabel metal2 s 131095 -480 131151 240 8 la_data_in[38]
port 205 nsew default input
rlabel metal2 s 132889 -480 132945 240 8 la_data_in[39]
port 206 nsew default input
rlabel metal2 s 68627 -480 68683 240 8 la_data_in[3]
port 207 nsew default input
rlabel metal2 s 134637 -480 134693 240 8 la_data_in[40]
port 208 nsew default input
rlabel metal2 s 136431 -480 136487 240 8 la_data_in[41]
port 209 nsew default input
rlabel metal2 s 138225 -480 138281 240 8 la_data_in[42]
port 210 nsew default input
rlabel metal2 s 140019 -480 140075 240 8 la_data_in[43]
port 211 nsew default input
rlabel metal2 s 141813 -480 141869 240 8 la_data_in[44]
port 212 nsew default input
rlabel metal2 s 143561 -480 143617 240 8 la_data_in[45]
port 213 nsew default input
rlabel metal2 s 145355 -480 145411 240 8 la_data_in[46]
port 214 nsew default input
rlabel metal2 s 147149 -480 147205 240 8 la_data_in[47]
port 215 nsew default input
rlabel metal2 s 148943 -480 148999 240 8 la_data_in[48]
port 216 nsew default input
rlabel metal2 s 150691 -480 150747 240 8 la_data_in[49]
port 217 nsew default input
rlabel metal2 s 70421 -480 70477 240 8 la_data_in[4]
port 218 nsew default input
rlabel metal2 s 152485 -480 152541 240 8 la_data_in[50]
port 219 nsew default input
rlabel metal2 s 154279 -480 154335 240 8 la_data_in[51]
port 220 nsew default input
rlabel metal2 s 156073 -480 156129 240 8 la_data_in[52]
port 221 nsew default input
rlabel metal2 s 157867 -480 157923 240 8 la_data_in[53]
port 222 nsew default input
rlabel metal2 s 159615 -480 159671 240 8 la_data_in[54]
port 223 nsew default input
rlabel metal2 s 161409 -480 161465 240 8 la_data_in[55]
port 224 nsew default input
rlabel metal2 s 163203 -480 163259 240 8 la_data_in[56]
port 225 nsew default input
rlabel metal2 s 164997 -480 165053 240 8 la_data_in[57]
port 226 nsew default input
rlabel metal2 s 166791 -480 166847 240 8 la_data_in[58]
port 227 nsew default input
rlabel metal2 s 168539 -480 168595 240 8 la_data_in[59]
port 228 nsew default input
rlabel metal2 s 72215 -480 72271 240 8 la_data_in[5]
port 229 nsew default input
rlabel metal2 s 170333 -480 170389 240 8 la_data_in[60]
port 230 nsew default input
rlabel metal2 s 172127 -480 172183 240 8 la_data_in[61]
port 231 nsew default input
rlabel metal2 s 173921 -480 173977 240 8 la_data_in[62]
port 232 nsew default input
rlabel metal2 s 175669 -480 175725 240 8 la_data_in[63]
port 233 nsew default input
rlabel metal2 s 177463 -480 177519 240 8 la_data_in[64]
port 234 nsew default input
rlabel metal2 s 179257 -480 179313 240 8 la_data_in[65]
port 235 nsew default input
rlabel metal2 s 181051 -480 181107 240 8 la_data_in[66]
port 236 nsew default input
rlabel metal2 s 182845 -480 182901 240 8 la_data_in[67]
port 237 nsew default input
rlabel metal2 s 184593 -480 184649 240 8 la_data_in[68]
port 238 nsew default input
rlabel metal2 s 186387 -480 186443 240 8 la_data_in[69]
port 239 nsew default input
rlabel metal2 s 74009 -480 74065 240 8 la_data_in[6]
port 240 nsew default input
rlabel metal2 s 188181 -480 188237 240 8 la_data_in[70]
port 241 nsew default input
rlabel metal2 s 189975 -480 190031 240 8 la_data_in[71]
port 242 nsew default input
rlabel metal2 s 191769 -480 191825 240 8 la_data_in[72]
port 243 nsew default input
rlabel metal2 s 193517 -480 193573 240 8 la_data_in[73]
port 244 nsew default input
rlabel metal2 s 195311 -480 195367 240 8 la_data_in[74]
port 245 nsew default input
rlabel metal2 s 197105 -480 197161 240 8 la_data_in[75]
port 246 nsew default input
rlabel metal2 s 198899 -480 198955 240 8 la_data_in[76]
port 247 nsew default input
rlabel metal2 s 200647 -480 200703 240 8 la_data_in[77]
port 248 nsew default input
rlabel metal2 s 202441 -480 202497 240 8 la_data_in[78]
port 249 nsew default input
rlabel metal2 s 204235 -480 204291 240 8 la_data_in[79]
port 250 nsew default input
rlabel metal2 s 75757 -480 75813 240 8 la_data_in[7]
port 251 nsew default input
rlabel metal2 s 206029 -480 206085 240 8 la_data_in[80]
port 252 nsew default input
rlabel metal2 s 207823 -480 207879 240 8 la_data_in[81]
port 253 nsew default input
rlabel metal2 s 209571 -480 209627 240 8 la_data_in[82]
port 254 nsew default input
rlabel metal2 s 211365 -480 211421 240 8 la_data_in[83]
port 255 nsew default input
rlabel metal2 s 213159 -480 213215 240 8 la_data_in[84]
port 256 nsew default input
rlabel metal2 s 214953 -480 215009 240 8 la_data_in[85]
port 257 nsew default input
rlabel metal2 s 216747 -480 216803 240 8 la_data_in[86]
port 258 nsew default input
rlabel metal2 s 218495 -480 218551 240 8 la_data_in[87]
port 259 nsew default input
rlabel metal2 s 220289 -480 220345 240 8 la_data_in[88]
port 260 nsew default input
rlabel metal2 s 222083 -480 222139 240 8 la_data_in[89]
port 261 nsew default input
rlabel metal2 s 77551 -480 77607 240 8 la_data_in[8]
port 262 nsew default input
rlabel metal2 s 223877 -480 223933 240 8 la_data_in[90]
port 263 nsew default input
rlabel metal2 s 225625 -480 225681 240 8 la_data_in[91]
port 264 nsew default input
rlabel metal2 s 227419 -480 227475 240 8 la_data_in[92]
port 265 nsew default input
rlabel metal2 s 229213 -480 229269 240 8 la_data_in[93]
port 266 nsew default input
rlabel metal2 s 231007 -480 231063 240 8 la_data_in[94]
port 267 nsew default input
rlabel metal2 s 232801 -480 232857 240 8 la_data_in[95]
port 268 nsew default input
rlabel metal2 s 234549 -480 234605 240 8 la_data_in[96]
port 269 nsew default input
rlabel metal2 s 236343 -480 236399 240 8 la_data_in[97]
port 270 nsew default input
rlabel metal2 s 238137 -480 238193 240 8 la_data_in[98]
port 271 nsew default input
rlabel metal2 s 239931 -480 239987 240 8 la_data_in[99]
port 272 nsew default input
rlabel metal2 s 79345 -480 79401 240 8 la_data_in[9]
port 273 nsew default input
rlabel metal2 s 63889 -480 63945 240 8 la_data_out[0]
port 274 nsew default output
rlabel metal2 s 242277 -480 242333 240 8 la_data_out[100]
port 275 nsew default output
rlabel metal2 s 244071 -480 244127 240 8 la_data_out[101]
port 276 nsew default output
rlabel metal2 s 245865 -480 245921 240 8 la_data_out[102]
port 277 nsew default output
rlabel metal2 s 247659 -480 247715 240 8 la_data_out[103]
port 278 nsew default output
rlabel metal2 s 249453 -480 249509 240 8 la_data_out[104]
port 279 nsew default output
rlabel metal2 s 251201 -480 251257 240 8 la_data_out[105]
port 280 nsew default output
rlabel metal2 s 252995 -480 253051 240 8 la_data_out[106]
port 281 nsew default output
rlabel metal2 s 254789 -480 254845 240 8 la_data_out[107]
port 282 nsew default output
rlabel metal2 s 256583 -480 256639 240 8 la_data_out[108]
port 283 nsew default output
rlabel metal2 s 258377 -480 258433 240 8 la_data_out[109]
port 284 nsew default output
rlabel metal2 s 81737 -480 81793 240 8 la_data_out[10]
port 285 nsew default output
rlabel metal2 s 260125 -480 260181 240 8 la_data_out[110]
port 286 nsew default output
rlabel metal2 s 261919 -480 261975 240 8 la_data_out[111]
port 287 nsew default output
rlabel metal2 s 263713 -480 263769 240 8 la_data_out[112]
port 288 nsew default output
rlabel metal2 s 265507 -480 265563 240 8 la_data_out[113]
port 289 nsew default output
rlabel metal2 s 267255 -480 267311 240 8 la_data_out[114]
port 290 nsew default output
rlabel metal2 s 269049 -480 269105 240 8 la_data_out[115]
port 291 nsew default output
rlabel metal2 s 270843 -480 270899 240 8 la_data_out[116]
port 292 nsew default output
rlabel metal2 s 272637 -480 272693 240 8 la_data_out[117]
port 293 nsew default output
rlabel metal2 s 274431 -480 274487 240 8 la_data_out[118]
port 294 nsew default output
rlabel metal2 s 276179 -480 276235 240 8 la_data_out[119]
port 295 nsew default output
rlabel metal2 s 83531 -480 83587 240 8 la_data_out[11]
port 296 nsew default output
rlabel metal2 s 277973 -480 278029 240 8 la_data_out[120]
port 297 nsew default output
rlabel metal2 s 279767 -480 279823 240 8 la_data_out[121]
port 298 nsew default output
rlabel metal2 s 281561 -480 281617 240 8 la_data_out[122]
port 299 nsew default output
rlabel metal2 s 283355 -480 283411 240 8 la_data_out[123]
port 300 nsew default output
rlabel metal2 s 285103 -480 285159 240 8 la_data_out[124]
port 301 nsew default output
rlabel metal2 s 286897 -480 286953 240 8 la_data_out[125]
port 302 nsew default output
rlabel metal2 s 288691 -480 288747 240 8 la_data_out[126]
port 303 nsew default output
rlabel metal2 s 290485 -480 290541 240 8 la_data_out[127]
port 304 nsew default output
rlabel metal2 s 85279 -480 85335 240 8 la_data_out[12]
port 305 nsew default output
rlabel metal2 s 87073 -480 87129 240 8 la_data_out[13]
port 306 nsew default output
rlabel metal2 s 88867 -480 88923 240 8 la_data_out[14]
port 307 nsew default output
rlabel metal2 s 90661 -480 90717 240 8 la_data_out[15]
port 308 nsew default output
rlabel metal2 s 92409 -480 92465 240 8 la_data_out[16]
port 309 nsew default output
rlabel metal2 s 94203 -480 94259 240 8 la_data_out[17]
port 310 nsew default output
rlabel metal2 s 95997 -480 96053 240 8 la_data_out[18]
port 311 nsew default output
rlabel metal2 s 97791 -480 97847 240 8 la_data_out[19]
port 312 nsew default output
rlabel metal2 s 65683 -480 65739 240 8 la_data_out[1]
port 313 nsew default output
rlabel metal2 s 99585 -480 99641 240 8 la_data_out[20]
port 314 nsew default output
rlabel metal2 s 101333 -480 101389 240 8 la_data_out[21]
port 315 nsew default output
rlabel metal2 s 103127 -480 103183 240 8 la_data_out[22]
port 316 nsew default output
rlabel metal2 s 104921 -480 104977 240 8 la_data_out[23]
port 317 nsew default output
rlabel metal2 s 106715 -480 106771 240 8 la_data_out[24]
port 318 nsew default output
rlabel metal2 s 108509 -480 108565 240 8 la_data_out[25]
port 319 nsew default output
rlabel metal2 s 110257 -480 110313 240 8 la_data_out[26]
port 320 nsew default output
rlabel metal2 s 112051 -480 112107 240 8 la_data_out[27]
port 321 nsew default output
rlabel metal2 s 113845 -480 113901 240 8 la_data_out[28]
port 322 nsew default output
rlabel metal2 s 115639 -480 115695 240 8 la_data_out[29]
port 323 nsew default output
rlabel metal2 s 67431 -480 67487 240 8 la_data_out[2]
port 324 nsew default output
rlabel metal2 s 117387 -480 117443 240 8 la_data_out[30]
port 325 nsew default output
rlabel metal2 s 119181 -480 119237 240 8 la_data_out[31]
port 326 nsew default output
rlabel metal2 s 120975 -480 121031 240 8 la_data_out[32]
port 327 nsew default output
rlabel metal2 s 122769 -480 122825 240 8 la_data_out[33]
port 328 nsew default output
rlabel metal2 s 124563 -480 124619 240 8 la_data_out[34]
port 329 nsew default output
rlabel metal2 s 126311 -480 126367 240 8 la_data_out[35]
port 330 nsew default output
rlabel metal2 s 128105 -480 128161 240 8 la_data_out[36]
port 331 nsew default output
rlabel metal2 s 129899 -480 129955 240 8 la_data_out[37]
port 332 nsew default output
rlabel metal2 s 131693 -480 131749 240 8 la_data_out[38]
port 333 nsew default output
rlabel metal2 s 133487 -480 133543 240 8 la_data_out[39]
port 334 nsew default output
rlabel metal2 s 69225 -480 69281 240 8 la_data_out[3]
port 335 nsew default output
rlabel metal2 s 135235 -480 135291 240 8 la_data_out[40]
port 336 nsew default output
rlabel metal2 s 137029 -480 137085 240 8 la_data_out[41]
port 337 nsew default output
rlabel metal2 s 138823 -480 138879 240 8 la_data_out[42]
port 338 nsew default output
rlabel metal2 s 140617 -480 140673 240 8 la_data_out[43]
port 339 nsew default output
rlabel metal2 s 142365 -480 142421 240 8 la_data_out[44]
port 340 nsew default output
rlabel metal2 s 144159 -480 144215 240 8 la_data_out[45]
port 341 nsew default output
rlabel metal2 s 145953 -480 146009 240 8 la_data_out[46]
port 342 nsew default output
rlabel metal2 s 147747 -480 147803 240 8 la_data_out[47]
port 343 nsew default output
rlabel metal2 s 149541 -480 149597 240 8 la_data_out[48]
port 344 nsew default output
rlabel metal2 s 151289 -480 151345 240 8 la_data_out[49]
port 345 nsew default output
rlabel metal2 s 71019 -480 71075 240 8 la_data_out[4]
port 346 nsew default output
rlabel metal2 s 153083 -480 153139 240 8 la_data_out[50]
port 347 nsew default output
rlabel metal2 s 154877 -480 154933 240 8 la_data_out[51]
port 348 nsew default output
rlabel metal2 s 156671 -480 156727 240 8 la_data_out[52]
port 349 nsew default output
rlabel metal2 s 158465 -480 158521 240 8 la_data_out[53]
port 350 nsew default output
rlabel metal2 s 160213 -480 160269 240 8 la_data_out[54]
port 351 nsew default output
rlabel metal2 s 162007 -480 162063 240 8 la_data_out[55]
port 352 nsew default output
rlabel metal2 s 163801 -480 163857 240 8 la_data_out[56]
port 353 nsew default output
rlabel metal2 s 165595 -480 165651 240 8 la_data_out[57]
port 354 nsew default output
rlabel metal2 s 167343 -480 167399 240 8 la_data_out[58]
port 355 nsew default output
rlabel metal2 s 169137 -480 169193 240 8 la_data_out[59]
port 356 nsew default output
rlabel metal2 s 72813 -480 72869 240 8 la_data_out[5]
port 357 nsew default output
rlabel metal2 s 170931 -480 170987 240 8 la_data_out[60]
port 358 nsew default output
rlabel metal2 s 172725 -480 172781 240 8 la_data_out[61]
port 359 nsew default output
rlabel metal2 s 174519 -480 174575 240 8 la_data_out[62]
port 360 nsew default output
rlabel metal2 s 176267 -480 176323 240 8 la_data_out[63]
port 361 nsew default output
rlabel metal2 s 178061 -480 178117 240 8 la_data_out[64]
port 362 nsew default output
rlabel metal2 s 179855 -480 179911 240 8 la_data_out[65]
port 363 nsew default output
rlabel metal2 s 181649 -480 181705 240 8 la_data_out[66]
port 364 nsew default output
rlabel metal2 s 183443 -480 183499 240 8 la_data_out[67]
port 365 nsew default output
rlabel metal2 s 185191 -480 185247 240 8 la_data_out[68]
port 366 nsew default output
rlabel metal2 s 186985 -480 187041 240 8 la_data_out[69]
port 367 nsew default output
rlabel metal2 s 74607 -480 74663 240 8 la_data_out[6]
port 368 nsew default output
rlabel metal2 s 188779 -480 188835 240 8 la_data_out[70]
port 369 nsew default output
rlabel metal2 s 190573 -480 190629 240 8 la_data_out[71]
port 370 nsew default output
rlabel metal2 s 192321 -480 192377 240 8 la_data_out[72]
port 371 nsew default output
rlabel metal2 s 194115 -480 194171 240 8 la_data_out[73]
port 372 nsew default output
rlabel metal2 s 195909 -480 195965 240 8 la_data_out[74]
port 373 nsew default output
rlabel metal2 s 197703 -480 197759 240 8 la_data_out[75]
port 374 nsew default output
rlabel metal2 s 199497 -480 199553 240 8 la_data_out[76]
port 375 nsew default output
rlabel metal2 s 201245 -480 201301 240 8 la_data_out[77]
port 376 nsew default output
rlabel metal2 s 203039 -480 203095 240 8 la_data_out[78]
port 377 nsew default output
rlabel metal2 s 204833 -480 204889 240 8 la_data_out[79]
port 378 nsew default output
rlabel metal2 s 76355 -480 76411 240 8 la_data_out[7]
port 379 nsew default output
rlabel metal2 s 206627 -480 206683 240 8 la_data_out[80]
port 380 nsew default output
rlabel metal2 s 208421 -480 208477 240 8 la_data_out[81]
port 381 nsew default output
rlabel metal2 s 210169 -480 210225 240 8 la_data_out[82]
port 382 nsew default output
rlabel metal2 s 211963 -480 212019 240 8 la_data_out[83]
port 383 nsew default output
rlabel metal2 s 213757 -480 213813 240 8 la_data_out[84]
port 384 nsew default output
rlabel metal2 s 215551 -480 215607 240 8 la_data_out[85]
port 385 nsew default output
rlabel metal2 s 217299 -480 217355 240 8 la_data_out[86]
port 386 nsew default output
rlabel metal2 s 219093 -480 219149 240 8 la_data_out[87]
port 387 nsew default output
rlabel metal2 s 220887 -480 220943 240 8 la_data_out[88]
port 388 nsew default output
rlabel metal2 s 222681 -480 222737 240 8 la_data_out[89]
port 389 nsew default output
rlabel metal2 s 78149 -480 78205 240 8 la_data_out[8]
port 390 nsew default output
rlabel metal2 s 224475 -480 224531 240 8 la_data_out[90]
port 391 nsew default output
rlabel metal2 s 226223 -480 226279 240 8 la_data_out[91]
port 392 nsew default output
rlabel metal2 s 228017 -480 228073 240 8 la_data_out[92]
port 393 nsew default output
rlabel metal2 s 229811 -480 229867 240 8 la_data_out[93]
port 394 nsew default output
rlabel metal2 s 231605 -480 231661 240 8 la_data_out[94]
port 395 nsew default output
rlabel metal2 s 233399 -480 233455 240 8 la_data_out[95]
port 396 nsew default output
rlabel metal2 s 235147 -480 235203 240 8 la_data_out[96]
port 397 nsew default output
rlabel metal2 s 236941 -480 236997 240 8 la_data_out[97]
port 398 nsew default output
rlabel metal2 s 238735 -480 238791 240 8 la_data_out[98]
port 399 nsew default output
rlabel metal2 s 240529 -480 240585 240 8 la_data_out[99]
port 400 nsew default output
rlabel metal2 s 79943 -480 79999 240 8 la_data_out[9]
port 401 nsew default output
rlabel metal2 s 64487 -480 64543 240 8 la_oen[0]
port 402 nsew default input
rlabel metal2 s 242875 -480 242931 240 8 la_oen[100]
port 403 nsew default input
rlabel metal2 s 244669 -480 244725 240 8 la_oen[101]
port 404 nsew default input
rlabel metal2 s 246463 -480 246519 240 8 la_oen[102]
port 405 nsew default input
rlabel metal2 s 248257 -480 248313 240 8 la_oen[103]
port 406 nsew default input
rlabel metal2 s 250051 -480 250107 240 8 la_oen[104]
port 407 nsew default input
rlabel metal2 s 251799 -480 251855 240 8 la_oen[105]
port 408 nsew default input
rlabel metal2 s 253593 -480 253649 240 8 la_oen[106]
port 409 nsew default input
rlabel metal2 s 255387 -480 255443 240 8 la_oen[107]
port 410 nsew default input
rlabel metal2 s 257181 -480 257237 240 8 la_oen[108]
port 411 nsew default input
rlabel metal2 s 258929 -480 258985 240 8 la_oen[109]
port 412 nsew default input
rlabel metal2 s 82335 -480 82391 240 8 la_oen[10]
port 413 nsew default input
rlabel metal2 s 260723 -480 260779 240 8 la_oen[110]
port 414 nsew default input
rlabel metal2 s 262517 -480 262573 240 8 la_oen[111]
port 415 nsew default input
rlabel metal2 s 264311 -480 264367 240 8 la_oen[112]
port 416 nsew default input
rlabel metal2 s 266105 -480 266161 240 8 la_oen[113]
port 417 nsew default input
rlabel metal2 s 267853 -480 267909 240 8 la_oen[114]
port 418 nsew default input
rlabel metal2 s 269647 -480 269703 240 8 la_oen[115]
port 419 nsew default input
rlabel metal2 s 271441 -480 271497 240 8 la_oen[116]
port 420 nsew default input
rlabel metal2 s 273235 -480 273291 240 8 la_oen[117]
port 421 nsew default input
rlabel metal2 s 275029 -480 275085 240 8 la_oen[118]
port 422 nsew default input
rlabel metal2 s 276777 -480 276833 240 8 la_oen[119]
port 423 nsew default input
rlabel metal2 s 84083 -480 84139 240 8 la_oen[11]
port 424 nsew default input
rlabel metal2 s 278571 -480 278627 240 8 la_oen[120]
port 425 nsew default input
rlabel metal2 s 280365 -480 280421 240 8 la_oen[121]
port 426 nsew default input
rlabel metal2 s 282159 -480 282215 240 8 la_oen[122]
port 427 nsew default input
rlabel metal2 s 283907 -480 283963 240 8 la_oen[123]
port 428 nsew default input
rlabel metal2 s 285701 -480 285757 240 8 la_oen[124]
port 429 nsew default input
rlabel metal2 s 287495 -480 287551 240 8 la_oen[125]
port 430 nsew default input
rlabel metal2 s 289289 -480 289345 240 8 la_oen[126]
port 431 nsew default input
rlabel metal2 s 291083 -480 291139 240 8 la_oen[127]
port 432 nsew default input
rlabel metal2 s 85877 -480 85933 240 8 la_oen[12]
port 433 nsew default input
rlabel metal2 s 87671 -480 87727 240 8 la_oen[13]
port 434 nsew default input
rlabel metal2 s 89465 -480 89521 240 8 la_oen[14]
port 435 nsew default input
rlabel metal2 s 91259 -480 91315 240 8 la_oen[15]
port 436 nsew default input
rlabel metal2 s 93007 -480 93063 240 8 la_oen[16]
port 437 nsew default input
rlabel metal2 s 94801 -480 94857 240 8 la_oen[17]
port 438 nsew default input
rlabel metal2 s 96595 -480 96651 240 8 la_oen[18]
port 439 nsew default input
rlabel metal2 s 98389 -480 98445 240 8 la_oen[19]
port 440 nsew default input
rlabel metal2 s 66281 -480 66337 240 8 la_oen[1]
port 441 nsew default input
rlabel metal2 s 100183 -480 100239 240 8 la_oen[20]
port 442 nsew default input
rlabel metal2 s 101931 -480 101987 240 8 la_oen[21]
port 443 nsew default input
rlabel metal2 s 103725 -480 103781 240 8 la_oen[22]
port 444 nsew default input
rlabel metal2 s 105519 -480 105575 240 8 la_oen[23]
port 445 nsew default input
rlabel metal2 s 107313 -480 107369 240 8 la_oen[24]
port 446 nsew default input
rlabel metal2 s 109061 -480 109117 240 8 la_oen[25]
port 447 nsew default input
rlabel metal2 s 110855 -480 110911 240 8 la_oen[26]
port 448 nsew default input
rlabel metal2 s 112649 -480 112705 240 8 la_oen[27]
port 449 nsew default input
rlabel metal2 s 114443 -480 114499 240 8 la_oen[28]
port 450 nsew default input
rlabel metal2 s 116237 -480 116293 240 8 la_oen[29]
port 451 nsew default input
rlabel metal2 s 68029 -480 68085 240 8 la_oen[2]
port 452 nsew default input
rlabel metal2 s 117985 -480 118041 240 8 la_oen[30]
port 453 nsew default input
rlabel metal2 s 119779 -480 119835 240 8 la_oen[31]
port 454 nsew default input
rlabel metal2 s 121573 -480 121629 240 8 la_oen[32]
port 455 nsew default input
rlabel metal2 s 123367 -480 123423 240 8 la_oen[33]
port 456 nsew default input
rlabel metal2 s 125161 -480 125217 240 8 la_oen[34]
port 457 nsew default input
rlabel metal2 s 126909 -480 126965 240 8 la_oen[35]
port 458 nsew default input
rlabel metal2 s 128703 -480 128759 240 8 la_oen[36]
port 459 nsew default input
rlabel metal2 s 130497 -480 130553 240 8 la_oen[37]
port 460 nsew default input
rlabel metal2 s 132291 -480 132347 240 8 la_oen[38]
port 461 nsew default input
rlabel metal2 s 134039 -480 134095 240 8 la_oen[39]
port 462 nsew default input
rlabel metal2 s 69823 -480 69879 240 8 la_oen[3]
port 463 nsew default input
rlabel metal2 s 135833 -480 135889 240 8 la_oen[40]
port 464 nsew default input
rlabel metal2 s 137627 -480 137683 240 8 la_oen[41]
port 465 nsew default input
rlabel metal2 s 139421 -480 139477 240 8 la_oen[42]
port 466 nsew default input
rlabel metal2 s 141215 -480 141271 240 8 la_oen[43]
port 467 nsew default input
rlabel metal2 s 142963 -480 143019 240 8 la_oen[44]
port 468 nsew default input
rlabel metal2 s 144757 -480 144813 240 8 la_oen[45]
port 469 nsew default input
rlabel metal2 s 146551 -480 146607 240 8 la_oen[46]
port 470 nsew default input
rlabel metal2 s 148345 -480 148401 240 8 la_oen[47]
port 471 nsew default input
rlabel metal2 s 150139 -480 150195 240 8 la_oen[48]
port 472 nsew default input
rlabel metal2 s 151887 -480 151943 240 8 la_oen[49]
port 473 nsew default input
rlabel metal2 s 71617 -480 71673 240 8 la_oen[4]
port 474 nsew default input
rlabel metal2 s 153681 -480 153737 240 8 la_oen[50]
port 475 nsew default input
rlabel metal2 s 155475 -480 155531 240 8 la_oen[51]
port 476 nsew default input
rlabel metal2 s 157269 -480 157325 240 8 la_oen[52]
port 477 nsew default input
rlabel metal2 s 159017 -480 159073 240 8 la_oen[53]
port 478 nsew default input
rlabel metal2 s 160811 -480 160867 240 8 la_oen[54]
port 479 nsew default input
rlabel metal2 s 162605 -480 162661 240 8 la_oen[55]
port 480 nsew default input
rlabel metal2 s 164399 -480 164455 240 8 la_oen[56]
port 481 nsew default input
rlabel metal2 s 166193 -480 166249 240 8 la_oen[57]
port 482 nsew default input
rlabel metal2 s 167941 -480 167997 240 8 la_oen[58]
port 483 nsew default input
rlabel metal2 s 169735 -480 169791 240 8 la_oen[59]
port 484 nsew default input
rlabel metal2 s 73411 -480 73467 240 8 la_oen[5]
port 485 nsew default input
rlabel metal2 s 171529 -480 171585 240 8 la_oen[60]
port 486 nsew default input
rlabel metal2 s 173323 -480 173379 240 8 la_oen[61]
port 487 nsew default input
rlabel metal2 s 175117 -480 175173 240 8 la_oen[62]
port 488 nsew default input
rlabel metal2 s 176865 -480 176921 240 8 la_oen[63]
port 489 nsew default input
rlabel metal2 s 178659 -480 178715 240 8 la_oen[64]
port 490 nsew default input
rlabel metal2 s 180453 -480 180509 240 8 la_oen[65]
port 491 nsew default input
rlabel metal2 s 182247 -480 182303 240 8 la_oen[66]
port 492 nsew default input
rlabel metal2 s 183995 -480 184051 240 8 la_oen[67]
port 493 nsew default input
rlabel metal2 s 185789 -480 185845 240 8 la_oen[68]
port 494 nsew default input
rlabel metal2 s 187583 -480 187639 240 8 la_oen[69]
port 495 nsew default input
rlabel metal2 s 75205 -480 75261 240 8 la_oen[6]
port 496 nsew default input
rlabel metal2 s 189377 -480 189433 240 8 la_oen[70]
port 497 nsew default input
rlabel metal2 s 191171 -480 191227 240 8 la_oen[71]
port 498 nsew default input
rlabel metal2 s 192919 -480 192975 240 8 la_oen[72]
port 499 nsew default input
rlabel metal2 s 194713 -480 194769 240 8 la_oen[73]
port 500 nsew default input
rlabel metal2 s 196507 -480 196563 240 8 la_oen[74]
port 501 nsew default input
rlabel metal2 s 198301 -480 198357 240 8 la_oen[75]
port 502 nsew default input
rlabel metal2 s 200095 -480 200151 240 8 la_oen[76]
port 503 nsew default input
rlabel metal2 s 201843 -480 201899 240 8 la_oen[77]
port 504 nsew default input
rlabel metal2 s 203637 -480 203693 240 8 la_oen[78]
port 505 nsew default input
rlabel metal2 s 205431 -480 205487 240 8 la_oen[79]
port 506 nsew default input
rlabel metal2 s 76953 -480 77009 240 8 la_oen[7]
port 507 nsew default input
rlabel metal2 s 207225 -480 207281 240 8 la_oen[80]
port 508 nsew default input
rlabel metal2 s 208973 -480 209029 240 8 la_oen[81]
port 509 nsew default input
rlabel metal2 s 210767 -480 210823 240 8 la_oen[82]
port 510 nsew default input
rlabel metal2 s 212561 -480 212617 240 8 la_oen[83]
port 511 nsew default input
rlabel metal2 s 214355 -480 214411 240 8 la_oen[84]
port 512 nsew default input
rlabel metal2 s 216149 -480 216205 240 8 la_oen[85]
port 513 nsew default input
rlabel metal2 s 217897 -480 217953 240 8 la_oen[86]
port 514 nsew default input
rlabel metal2 s 219691 -480 219747 240 8 la_oen[87]
port 515 nsew default input
rlabel metal2 s 221485 -480 221541 240 8 la_oen[88]
port 516 nsew default input
rlabel metal2 s 223279 -480 223335 240 8 la_oen[89]
port 517 nsew default input
rlabel metal2 s 78747 -480 78803 240 8 la_oen[8]
port 518 nsew default input
rlabel metal2 s 225073 -480 225129 240 8 la_oen[90]
port 519 nsew default input
rlabel metal2 s 226821 -480 226877 240 8 la_oen[91]
port 520 nsew default input
rlabel metal2 s 228615 -480 228671 240 8 la_oen[92]
port 521 nsew default input
rlabel metal2 s 230409 -480 230465 240 8 la_oen[93]
port 522 nsew default input
rlabel metal2 s 232203 -480 232259 240 8 la_oen[94]
port 523 nsew default input
rlabel metal2 s 233951 -480 234007 240 8 la_oen[95]
port 524 nsew default input
rlabel metal2 s 235745 -480 235801 240 8 la_oen[96]
port 525 nsew default input
rlabel metal2 s 237539 -480 237595 240 8 la_oen[97]
port 526 nsew default input
rlabel metal2 s 239333 -480 239389 240 8 la_oen[98]
port 527 nsew default input
rlabel metal2 s 241127 -480 241183 240 8 la_oen[99]
port 528 nsew default input
rlabel metal2 s 80541 -480 80597 240 8 la_oen[9]
port 529 nsew default input
rlabel metal2 s 291681 -480 291737 240 8 user_clock2
port 530 nsew default input
rlabel metal2 s 271 -480 327 240 8 wb_clk_i
port 531 nsew default input
rlabel metal2 s 823 -480 879 240 8 wb_rst_i
port 532 nsew default input
rlabel metal2 s 1421 -480 1477 240 8 wbs_ack_o
port 533 nsew default output
rlabel metal2 s 3813 -480 3869 240 8 wbs_adr_i[0]
port 534 nsew default input
rlabel metal2 s 24053 -480 24109 240 8 wbs_adr_i[10]
port 535 nsew default input
rlabel metal2 s 25801 -480 25857 240 8 wbs_adr_i[11]
port 536 nsew default input
rlabel metal2 s 27595 -480 27651 240 8 wbs_adr_i[12]
port 537 nsew default input
rlabel metal2 s 29389 -480 29445 240 8 wbs_adr_i[13]
port 538 nsew default input
rlabel metal2 s 31183 -480 31239 240 8 wbs_adr_i[14]
port 539 nsew default input
rlabel metal2 s 32977 -480 33033 240 8 wbs_adr_i[15]
port 540 nsew default input
rlabel metal2 s 34725 -480 34781 240 8 wbs_adr_i[16]
port 541 nsew default input
rlabel metal2 s 36519 -480 36575 240 8 wbs_adr_i[17]
port 542 nsew default input
rlabel metal2 s 38313 -480 38369 240 8 wbs_adr_i[18]
port 543 nsew default input
rlabel metal2 s 40107 -480 40163 240 8 wbs_adr_i[19]
port 544 nsew default input
rlabel metal2 s 6205 -480 6261 240 8 wbs_adr_i[1]
port 545 nsew default input
rlabel metal2 s 41901 -480 41957 240 8 wbs_adr_i[20]
port 546 nsew default input
rlabel metal2 s 43649 -480 43705 240 8 wbs_adr_i[21]
port 547 nsew default input
rlabel metal2 s 45443 -480 45499 240 8 wbs_adr_i[22]
port 548 nsew default input
rlabel metal2 s 47237 -480 47293 240 8 wbs_adr_i[23]
port 549 nsew default input
rlabel metal2 s 49031 -480 49087 240 8 wbs_adr_i[24]
port 550 nsew default input
rlabel metal2 s 50779 -480 50835 240 8 wbs_adr_i[25]
port 551 nsew default input
rlabel metal2 s 52573 -480 52629 240 8 wbs_adr_i[26]
port 552 nsew default input
rlabel metal2 s 54367 -480 54423 240 8 wbs_adr_i[27]
port 553 nsew default input
rlabel metal2 s 56161 -480 56217 240 8 wbs_adr_i[28]
port 554 nsew default input
rlabel metal2 s 57955 -480 58011 240 8 wbs_adr_i[29]
port 555 nsew default input
rlabel metal2 s 8597 -480 8653 240 8 wbs_adr_i[2]
port 556 nsew default input
rlabel metal2 s 59703 -480 59759 240 8 wbs_adr_i[30]
port 557 nsew default input
rlabel metal2 s 61497 -480 61553 240 8 wbs_adr_i[31]
port 558 nsew default input
rlabel metal2 s 10943 -480 10999 240 8 wbs_adr_i[3]
port 559 nsew default input
rlabel metal2 s 13335 -480 13391 240 8 wbs_adr_i[4]
port 560 nsew default input
rlabel metal2 s 15129 -480 15185 240 8 wbs_adr_i[5]
port 561 nsew default input
rlabel metal2 s 16923 -480 16979 240 8 wbs_adr_i[6]
port 562 nsew default input
rlabel metal2 s 18671 -480 18727 240 8 wbs_adr_i[7]
port 563 nsew default input
rlabel metal2 s 20465 -480 20521 240 8 wbs_adr_i[8]
port 564 nsew default input
rlabel metal2 s 22259 -480 22315 240 8 wbs_adr_i[9]
port 565 nsew default input
rlabel metal2 s 2019 -480 2075 240 8 wbs_cyc_i
port 566 nsew default input
rlabel metal2 s 4411 -480 4467 240 8 wbs_dat_i[0]
port 567 nsew default input
rlabel metal2 s 24651 -480 24707 240 8 wbs_dat_i[10]
port 568 nsew default input
rlabel metal2 s 26399 -480 26455 240 8 wbs_dat_i[11]
port 569 nsew default input
rlabel metal2 s 28193 -480 28249 240 8 wbs_dat_i[12]
port 570 nsew default input
rlabel metal2 s 29987 -480 30043 240 8 wbs_dat_i[13]
port 571 nsew default input
rlabel metal2 s 31781 -480 31837 240 8 wbs_dat_i[14]
port 572 nsew default input
rlabel metal2 s 33575 -480 33631 240 8 wbs_dat_i[15]
port 573 nsew default input
rlabel metal2 s 35323 -480 35379 240 8 wbs_dat_i[16]
port 574 nsew default input
rlabel metal2 s 37117 -480 37173 240 8 wbs_dat_i[17]
port 575 nsew default input
rlabel metal2 s 38911 -480 38967 240 8 wbs_dat_i[18]
port 576 nsew default input
rlabel metal2 s 40705 -480 40761 240 8 wbs_dat_i[19]
port 577 nsew default input
rlabel metal2 s 6803 -480 6859 240 8 wbs_dat_i[1]
port 578 nsew default input
rlabel metal2 s 42453 -480 42509 240 8 wbs_dat_i[20]
port 579 nsew default input
rlabel metal2 s 44247 -480 44303 240 8 wbs_dat_i[21]
port 580 nsew default input
rlabel metal2 s 46041 -480 46097 240 8 wbs_dat_i[22]
port 581 nsew default input
rlabel metal2 s 47835 -480 47891 240 8 wbs_dat_i[23]
port 582 nsew default input
rlabel metal2 s 49629 -480 49685 240 8 wbs_dat_i[24]
port 583 nsew default input
rlabel metal2 s 51377 -480 51433 240 8 wbs_dat_i[25]
port 584 nsew default input
rlabel metal2 s 53171 -480 53227 240 8 wbs_dat_i[26]
port 585 nsew default input
rlabel metal2 s 54965 -480 55021 240 8 wbs_dat_i[27]
port 586 nsew default input
rlabel metal2 s 56759 -480 56815 240 8 wbs_dat_i[28]
port 587 nsew default input
rlabel metal2 s 58553 -480 58609 240 8 wbs_dat_i[29]
port 588 nsew default input
rlabel metal2 s 9149 -480 9205 240 8 wbs_dat_i[2]
port 589 nsew default input
rlabel metal2 s 60301 -480 60357 240 8 wbs_dat_i[30]
port 590 nsew default input
rlabel metal2 s 62095 -480 62151 240 8 wbs_dat_i[31]
port 591 nsew default input
rlabel metal2 s 11541 -480 11597 240 8 wbs_dat_i[3]
port 592 nsew default input
rlabel metal2 s 13933 -480 13989 240 8 wbs_dat_i[4]
port 593 nsew default input
rlabel metal2 s 15727 -480 15783 240 8 wbs_dat_i[5]
port 594 nsew default input
rlabel metal2 s 17475 -480 17531 240 8 wbs_dat_i[6]
port 595 nsew default input
rlabel metal2 s 19269 -480 19325 240 8 wbs_dat_i[7]
port 596 nsew default input
rlabel metal2 s 21063 -480 21119 240 8 wbs_dat_i[8]
port 597 nsew default input
rlabel metal2 s 22857 -480 22913 240 8 wbs_dat_i[9]
port 598 nsew default input
rlabel metal2 s 5009 -480 5065 240 8 wbs_dat_o[0]
port 599 nsew default output
rlabel metal2 s 25249 -480 25305 240 8 wbs_dat_o[10]
port 600 nsew default output
rlabel metal2 s 26997 -480 27053 240 8 wbs_dat_o[11]
port 601 nsew default output
rlabel metal2 s 28791 -480 28847 240 8 wbs_dat_o[12]
port 602 nsew default output
rlabel metal2 s 30585 -480 30641 240 8 wbs_dat_o[13]
port 603 nsew default output
rlabel metal2 s 32379 -480 32435 240 8 wbs_dat_o[14]
port 604 nsew default output
rlabel metal2 s 34127 -480 34183 240 8 wbs_dat_o[15]
port 605 nsew default output
rlabel metal2 s 35921 -480 35977 240 8 wbs_dat_o[16]
port 606 nsew default output
rlabel metal2 s 37715 -480 37771 240 8 wbs_dat_o[17]
port 607 nsew default output
rlabel metal2 s 39509 -480 39565 240 8 wbs_dat_o[18]
port 608 nsew default output
rlabel metal2 s 41303 -480 41359 240 8 wbs_dat_o[19]
port 609 nsew default output
rlabel metal2 s 7401 -480 7457 240 8 wbs_dat_o[1]
port 610 nsew default output
rlabel metal2 s 43051 -480 43107 240 8 wbs_dat_o[20]
port 611 nsew default output
rlabel metal2 s 44845 -480 44901 240 8 wbs_dat_o[21]
port 612 nsew default output
rlabel metal2 s 46639 -480 46695 240 8 wbs_dat_o[22]
port 613 nsew default output
rlabel metal2 s 48433 -480 48489 240 8 wbs_dat_o[23]
port 614 nsew default output
rlabel metal2 s 50227 -480 50283 240 8 wbs_dat_o[24]
port 615 nsew default output
rlabel metal2 s 51975 -480 52031 240 8 wbs_dat_o[25]
port 616 nsew default output
rlabel metal2 s 53769 -480 53825 240 8 wbs_dat_o[26]
port 617 nsew default output
rlabel metal2 s 55563 -480 55619 240 8 wbs_dat_o[27]
port 618 nsew default output
rlabel metal2 s 57357 -480 57413 240 8 wbs_dat_o[28]
port 619 nsew default output
rlabel metal2 s 59105 -480 59161 240 8 wbs_dat_o[29]
port 620 nsew default output
rlabel metal2 s 9747 -480 9803 240 8 wbs_dat_o[2]
port 621 nsew default output
rlabel metal2 s 60899 -480 60955 240 8 wbs_dat_o[30]
port 622 nsew default output
rlabel metal2 s 62693 -480 62749 240 8 wbs_dat_o[31]
port 623 nsew default output
rlabel metal2 s 12139 -480 12195 240 8 wbs_dat_o[3]
port 624 nsew default output
rlabel metal2 s 14531 -480 14587 240 8 wbs_dat_o[4]
port 625 nsew default output
rlabel metal2 s 16325 -480 16381 240 8 wbs_dat_o[5]
port 626 nsew default output
rlabel metal2 s 18073 -480 18129 240 8 wbs_dat_o[6]
port 627 nsew default output
rlabel metal2 s 19867 -480 19923 240 8 wbs_dat_o[7]
port 628 nsew default output
rlabel metal2 s 21661 -480 21717 240 8 wbs_dat_o[8]
port 629 nsew default output
rlabel metal2 s 23455 -480 23511 240 8 wbs_dat_o[9]
port 630 nsew default output
rlabel metal2 s 5607 -480 5663 240 8 wbs_sel_i[0]
port 631 nsew default input
rlabel metal2 s 7999 -480 8055 240 8 wbs_sel_i[1]
port 632 nsew default input
rlabel metal2 s 10345 -480 10401 240 8 wbs_sel_i[2]
port 633 nsew default input
rlabel metal2 s 12737 -480 12793 240 8 wbs_sel_i[3]
port 634 nsew default input
rlabel metal2 s 2617 -480 2673 240 8 wbs_stb_i
port 635 nsew default input
rlabel metal2 s 3215 -480 3271 240 8 wbs_we_i
port 636 nsew default input
rlabel metal4 s 288402 351760 288702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 270402 351760 270702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 252402 351760 252702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 234402 351760 234702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 216402 351760 216702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 198402 351760 198702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 180402 351760 180702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 162402 351760 162702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 144402 351760 144702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 126402 351760 126702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 108402 351760 108702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 90402 351760 90702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 72402 351760 72702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 54402 351760 54702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 36402 351760 36702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 18402 351760 18702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 402 351760 702 352900 6 vccd1
port 637 nsew default input
rlabel metal4 s 292660 -462 292960 352430 6 vccd1
port 637 nsew default input
rlabel metal4 s -998 -462 -698 352430 4 vccd1
port 637 nsew default input
rlabel metal4 s 288402 -932 288702 240 8 vccd1
port 637 nsew default input
rlabel metal4 s 270402 -932 270702 240 8 vccd1
port 637 nsew default input
rlabel metal4 s 252402 -932 252702 240 8 vccd1
port 637 nsew default input
rlabel metal4 s 234402 -932 234702 240 8 vccd1
port 637 nsew default input
rlabel metal4 s 216402 -932 216702 240 8 vccd1
port 637 nsew default input
rlabel metal4 s 198402 -932 198702 240 8 vccd1
port 637 nsew default input
rlabel metal4 s 180402 -932 180702 240 8 vccd1
port 637 nsew default input
rlabel metal4 s 162402 -932 162702 240 8 vccd1
port 637 nsew default input
rlabel metal4 s 144402 -932 144702 240 8 vccd1
port 637 nsew default input
rlabel metal4 s 126402 -932 126702 240 8 vccd1
port 637 nsew default input
rlabel metal4 s 108402 -932 108702 240 8 vccd1
port 637 nsew default input
rlabel metal4 s 90402 -932 90702 240 8 vccd1
port 637 nsew default input
rlabel metal4 s 72402 -932 72702 240 8 vccd1
port 637 nsew default input
rlabel metal4 s 54402 -932 54702 240 8 vccd1
port 637 nsew default input
rlabel metal4 s 36402 -932 36702 240 8 vccd1
port 637 nsew default input
rlabel metal4 s 18402 -932 18702 240 8 vccd1
port 637 nsew default input
rlabel metal4 s 402 -932 702 240 8 vccd1
port 637 nsew default input
rlabel metal5 s -998 352130 292960 352430 6 vccd1
port 637 nsew default input
rlabel metal5 s 291760 342938 293430 343238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 342938 240 343238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 324938 293430 325238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 324938 240 325238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 306938 293430 307238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 306938 240 307238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 288938 293430 289238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 288938 240 289238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 270938 293430 271238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 270938 240 271238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 252938 293430 253238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 252938 240 253238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 234938 293430 235238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 234938 240 235238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 216938 293430 217238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 216938 240 217238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 198938 293430 199238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 198938 240 199238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 180938 293430 181238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 180938 240 181238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 162938 293430 163238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 162938 240 163238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 144938 293430 145238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 144938 240 145238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 126938 293430 127238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 126938 240 127238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 108938 293430 109238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 108938 240 109238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 90938 293430 91238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 90938 240 91238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 72938 293430 73238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 72938 240 73238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 54938 293430 55238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 54938 240 55238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 36938 293430 37238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 36938 240 37238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 18938 293430 19238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 18938 240 19238 4 vccd1
port 637 nsew default input
rlabel metal5 s 291760 938 293430 1238 6 vccd1
port 637 nsew default input
rlabel metal5 s -1468 938 240 1238 4 vccd1
port 637 nsew default input
rlabel metal5 s -998 -462 292960 -162 8 vccd1
port 637 nsew default input
rlabel metal4 s 293130 -932 293430 352900 6 vssd1
port 638 nsew default input
rlabel metal4 s 279402 351760 279702 352900 6 vssd1
port 638 nsew default input
rlabel metal4 s 261402 351760 261702 352900 6 vssd1
port 638 nsew default input
rlabel metal4 s 243402 351760 243702 352900 6 vssd1
port 638 nsew default input
rlabel metal4 s 225402 351760 225702 352900 6 vssd1
port 638 nsew default input
rlabel metal4 s 207402 351760 207702 352900 6 vssd1
port 638 nsew default input
rlabel metal4 s 189402 351760 189702 352900 6 vssd1
port 638 nsew default input
rlabel metal4 s 171402 351760 171702 352900 6 vssd1
port 638 nsew default input
rlabel metal4 s 153402 351760 153702 352900 6 vssd1
port 638 nsew default input
rlabel metal4 s 135402 351760 135702 352900 6 vssd1
port 638 nsew default input
rlabel metal4 s 117402 351760 117702 352900 6 vssd1
port 638 nsew default input
rlabel metal4 s 99402 351760 99702 352900 6 vssd1
port 638 nsew default input
rlabel metal4 s 81402 351760 81702 352900 6 vssd1
port 638 nsew default input
rlabel metal4 s 63402 351760 63702 352900 6 vssd1
port 638 nsew default input
rlabel metal4 s 45402 351760 45702 352900 6 vssd1
port 638 nsew default input
rlabel metal4 s 27402 351760 27702 352900 6 vssd1
port 638 nsew default input
rlabel metal4 s 9402 351760 9702 352900 6 vssd1
port 638 nsew default input
rlabel metal4 s -1468 -932 -1168 352900 4 vssd1
port 638 nsew default input
rlabel metal4 s 279402 -932 279702 240 8 vssd1
port 638 nsew default input
rlabel metal4 s 261402 -932 261702 240 8 vssd1
port 638 nsew default input
rlabel metal4 s 243402 -932 243702 240 8 vssd1
port 638 nsew default input
rlabel metal4 s 225402 -932 225702 240 8 vssd1
port 638 nsew default input
rlabel metal4 s 207402 -932 207702 240 8 vssd1
port 638 nsew default input
rlabel metal4 s 189402 -932 189702 240 8 vssd1
port 638 nsew default input
rlabel metal4 s 171402 -932 171702 240 8 vssd1
port 638 nsew default input
rlabel metal4 s 153402 -932 153702 240 8 vssd1
port 638 nsew default input
rlabel metal4 s 135402 -932 135702 240 8 vssd1
port 638 nsew default input
rlabel metal4 s 117402 -932 117702 240 8 vssd1
port 638 nsew default input
rlabel metal4 s 99402 -932 99702 240 8 vssd1
port 638 nsew default input
rlabel metal4 s 81402 -932 81702 240 8 vssd1
port 638 nsew default input
rlabel metal4 s 63402 -932 63702 240 8 vssd1
port 638 nsew default input
rlabel metal4 s 45402 -932 45702 240 8 vssd1
port 638 nsew default input
rlabel metal4 s 27402 -932 27702 240 8 vssd1
port 638 nsew default input
rlabel metal4 s 9402 -932 9702 240 8 vssd1
port 638 nsew default input
rlabel metal5 s -1468 352600 293430 352900 6 vssd1
port 638 nsew default input
rlabel metal5 s 291760 333938 293430 334238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 333938 240 334238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 315938 293430 316238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 315938 240 316238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 297938 293430 298238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 297938 240 298238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 279938 293430 280238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 279938 240 280238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 261938 293430 262238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 261938 240 262238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 243938 293430 244238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 243938 240 244238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 225938 293430 226238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 225938 240 226238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 207938 293430 208238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 207938 240 208238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 189938 293430 190238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 189938 240 190238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 171938 293430 172238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 171938 240 172238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 153938 293430 154238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 153938 240 154238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 135938 293430 136238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 135938 240 136238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 117938 293430 118238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 117938 240 118238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 99938 293430 100238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 99938 240 100238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 81938 293430 82238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 81938 240 82238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 63938 293430 64238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 63938 240 64238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 45938 293430 46238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 45938 240 46238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 27938 293430 28238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 27938 240 28238 4 vssd1
port 638 nsew default input
rlabel metal5 s 291760 9938 293430 10238 6 vssd1
port 638 nsew default input
rlabel metal5 s -1468 9938 240 10238 4 vssd1
port 638 nsew default input
rlabel metal5 s -1468 -932 293430 -632 8 vssd1
port 638 nsew default input
rlabel metal4 s 290202 351760 290502 353840 6 vccd2
port 639 nsew default input
rlabel metal4 s 272202 351760 272502 353840 6 vccd2
port 639 nsew default input
rlabel metal4 s 254202 351760 254502 353840 6 vccd2
port 639 nsew default input
rlabel metal4 s 236202 351760 236502 353840 6 vccd2
port 639 nsew default input
rlabel metal4 s 218202 351760 218502 353840 6 vccd2
port 639 nsew default input
rlabel metal4 s 200202 351760 200502 353840 6 vccd2
port 639 nsew default input
rlabel metal4 s 182202 351760 182502 353840 6 vccd2
port 639 nsew default input
rlabel metal4 s 164202 351760 164502 353840 6 vccd2
port 639 nsew default input
rlabel metal4 s 146202 351760 146502 353840 6 vccd2
port 639 nsew default input
rlabel metal4 s 128202 351760 128502 353840 6 vccd2
port 639 nsew default input
rlabel metal4 s 110202 351760 110502 353840 6 vccd2
port 639 nsew default input
rlabel metal4 s 92202 351760 92502 353840 6 vccd2
port 639 nsew default input
rlabel metal4 s 74202 351760 74502 353840 6 vccd2
port 639 nsew default input
rlabel metal4 s 56202 351760 56502 353840 6 vccd2
port 639 nsew default input
rlabel metal4 s 38202 351760 38502 353840 6 vccd2
port 639 nsew default input
rlabel metal4 s 20202 351760 20502 353840 6 vccd2
port 639 nsew default input
rlabel metal4 s 2202 351760 2502 353840 6 vccd2
port 639 nsew default input
rlabel metal4 s 293600 -1402 293900 353370 6 vccd2
port 639 nsew default input
rlabel metal4 s -1938 -1402 -1638 353370 4 vccd2
port 639 nsew default input
rlabel metal4 s 290202 -1872 290502 240 8 vccd2
port 639 nsew default input
rlabel metal4 s 272202 -1872 272502 240 8 vccd2
port 639 nsew default input
rlabel metal4 s 254202 -1872 254502 240 8 vccd2
port 639 nsew default input
rlabel metal4 s 236202 -1872 236502 240 8 vccd2
port 639 nsew default input
rlabel metal4 s 218202 -1872 218502 240 8 vccd2
port 639 nsew default input
rlabel metal4 s 200202 -1872 200502 240 8 vccd2
port 639 nsew default input
rlabel metal4 s 182202 -1872 182502 240 8 vccd2
port 639 nsew default input
rlabel metal4 s 164202 -1872 164502 240 8 vccd2
port 639 nsew default input
rlabel metal4 s 146202 -1872 146502 240 8 vccd2
port 639 nsew default input
rlabel metal4 s 128202 -1872 128502 240 8 vccd2
port 639 nsew default input
rlabel metal4 s 110202 -1872 110502 240 8 vccd2
port 639 nsew default input
rlabel metal4 s 92202 -1872 92502 240 8 vccd2
port 639 nsew default input
rlabel metal4 s 74202 -1872 74502 240 8 vccd2
port 639 nsew default input
rlabel metal4 s 56202 -1872 56502 240 8 vccd2
port 639 nsew default input
rlabel metal4 s 38202 -1872 38502 240 8 vccd2
port 639 nsew default input
rlabel metal4 s 20202 -1872 20502 240 8 vccd2
port 639 nsew default input
rlabel metal4 s 2202 -1872 2502 240 8 vccd2
port 639 nsew default input
rlabel metal5 s -1938 353070 293900 353370 6 vccd2
port 639 nsew default input
rlabel metal5 s 291760 344738 294370 345038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 344738 240 345038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 326738 294370 327038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 326738 240 327038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 308738 294370 309038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 308738 240 309038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 290738 294370 291038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 290738 240 291038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 272738 294370 273038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 272738 240 273038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 254738 294370 255038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 254738 240 255038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 236738 294370 237038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 236738 240 237038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 218738 294370 219038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 218738 240 219038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 200738 294370 201038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 200738 240 201038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 182738 294370 183038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 182738 240 183038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 164738 294370 165038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 164738 240 165038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 146738 294370 147038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 146738 240 147038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 128738 294370 129038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 128738 240 129038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 110738 294370 111038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 110738 240 111038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 92738 294370 93038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 92738 240 93038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 74738 294370 75038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 74738 240 75038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 56738 294370 57038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 56738 240 57038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 38738 294370 39038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 38738 240 39038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 20738 294370 21038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 20738 240 21038 4 vccd2
port 639 nsew default input
rlabel metal5 s 291760 2738 294370 3038 6 vccd2
port 639 nsew default input
rlabel metal5 s -2408 2738 240 3038 4 vccd2
port 639 nsew default input
rlabel metal5 s -1938 -1402 293900 -1102 8 vccd2
port 639 nsew default input
rlabel metal4 s 294070 -1872 294370 353840 6 vssd2
port 640 nsew default input
rlabel metal4 s 281202 351760 281502 353840 6 vssd2
port 640 nsew default input
rlabel metal4 s 263202 351760 263502 353840 6 vssd2
port 640 nsew default input
rlabel metal4 s 245202 351760 245502 353840 6 vssd2
port 640 nsew default input
rlabel metal4 s 227202 351760 227502 353840 6 vssd2
port 640 nsew default input
rlabel metal4 s 209202 351760 209502 353840 6 vssd2
port 640 nsew default input
rlabel metal4 s 191202 351760 191502 353840 6 vssd2
port 640 nsew default input
rlabel metal4 s 173202 351760 173502 353840 6 vssd2
port 640 nsew default input
rlabel metal4 s 155202 351760 155502 353840 6 vssd2
port 640 nsew default input
rlabel metal4 s 137202 351760 137502 353840 6 vssd2
port 640 nsew default input
rlabel metal4 s 119202 351760 119502 353840 6 vssd2
port 640 nsew default input
rlabel metal4 s 101202 351760 101502 353840 6 vssd2
port 640 nsew default input
rlabel metal4 s 83202 351760 83502 353840 6 vssd2
port 640 nsew default input
rlabel metal4 s 65202 351760 65502 353840 6 vssd2
port 640 nsew default input
rlabel metal4 s 47202 351760 47502 353840 6 vssd2
port 640 nsew default input
rlabel metal4 s 29202 351760 29502 353840 6 vssd2
port 640 nsew default input
rlabel metal4 s 11202 351760 11502 353840 6 vssd2
port 640 nsew default input
rlabel metal4 s -2408 -1872 -2108 353840 4 vssd2
port 640 nsew default input
rlabel metal4 s 281202 -1872 281502 240 8 vssd2
port 640 nsew default input
rlabel metal4 s 263202 -1872 263502 240 8 vssd2
port 640 nsew default input
rlabel metal4 s 245202 -1872 245502 240 8 vssd2
port 640 nsew default input
rlabel metal4 s 227202 -1872 227502 240 8 vssd2
port 640 nsew default input
rlabel metal4 s 209202 -1872 209502 240 8 vssd2
port 640 nsew default input
rlabel metal4 s 191202 -1872 191502 240 8 vssd2
port 640 nsew default input
rlabel metal4 s 173202 -1872 173502 240 8 vssd2
port 640 nsew default input
rlabel metal4 s 155202 -1872 155502 240 8 vssd2
port 640 nsew default input
rlabel metal4 s 137202 -1872 137502 240 8 vssd2
port 640 nsew default input
rlabel metal4 s 119202 -1872 119502 240 8 vssd2
port 640 nsew default input
rlabel metal4 s 101202 -1872 101502 240 8 vssd2
port 640 nsew default input
rlabel metal4 s 83202 -1872 83502 240 8 vssd2
port 640 nsew default input
rlabel metal4 s 65202 -1872 65502 240 8 vssd2
port 640 nsew default input
rlabel metal4 s 47202 -1872 47502 240 8 vssd2
port 640 nsew default input
rlabel metal4 s 29202 -1872 29502 240 8 vssd2
port 640 nsew default input
rlabel metal4 s 11202 -1872 11502 240 8 vssd2
port 640 nsew default input
rlabel metal5 s -2408 353540 294370 353840 6 vssd2
port 640 nsew default input
rlabel metal5 s 291760 335738 294370 336038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 335738 240 336038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 317738 294370 318038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 317738 240 318038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 299738 294370 300038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 299738 240 300038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 281738 294370 282038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 281738 240 282038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 263738 294370 264038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 263738 240 264038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 245738 294370 246038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 245738 240 246038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 227738 294370 228038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 227738 240 228038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 209738 294370 210038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 209738 240 210038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 191738 294370 192038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 191738 240 192038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 173738 294370 174038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 173738 240 174038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 155738 294370 156038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 155738 240 156038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 137738 294370 138038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 137738 240 138038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 119738 294370 120038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 119738 240 120038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 101738 294370 102038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 101738 240 102038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 83738 294370 84038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 83738 240 84038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 65738 294370 66038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 65738 240 66038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 47738 294370 48038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 47738 240 48038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 29738 294370 30038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 29738 240 30038 4 vssd2
port 640 nsew default input
rlabel metal5 s 291760 11738 294370 12038 6 vssd2
port 640 nsew default input
rlabel metal5 s -2408 11738 240 12038 4 vssd2
port 640 nsew default input
rlabel metal5 s -2408 -1872 294370 -1572 8 vssd2
port 640 nsew default input
rlabel metal4 s 274002 351760 274302 354780 6 vdda1
port 641 nsew default input
rlabel metal4 s 256002 351760 256302 354780 6 vdda1
port 641 nsew default input
rlabel metal4 s 238002 351760 238302 354780 6 vdda1
port 641 nsew default input
rlabel metal4 s 220002 351760 220302 354780 6 vdda1
port 641 nsew default input
rlabel metal4 s 202002 351760 202302 354780 6 vdda1
port 641 nsew default input
rlabel metal4 s 184002 351760 184302 354780 6 vdda1
port 641 nsew default input
rlabel metal4 s 166002 351760 166302 354780 6 vdda1
port 641 nsew default input
rlabel metal4 s 148002 351760 148302 354780 6 vdda1
port 641 nsew default input
rlabel metal4 s 130002 351760 130302 354780 6 vdda1
port 641 nsew default input
rlabel metal4 s 112002 351760 112302 354780 6 vdda1
port 641 nsew default input
rlabel metal4 s 94002 351760 94302 354780 6 vdda1
port 641 nsew default input
rlabel metal4 s 76002 351760 76302 354780 6 vdda1
port 641 nsew default input
rlabel metal4 s 58002 351760 58302 354780 6 vdda1
port 641 nsew default input
rlabel metal4 s 40002 351760 40302 354780 6 vdda1
port 641 nsew default input
rlabel metal4 s 22002 351760 22302 354780 6 vdda1
port 641 nsew default input
rlabel metal4 s 4002 351760 4302 354780 6 vdda1
port 641 nsew default input
rlabel metal4 s 294540 -2342 294840 354310 6 vdda1
port 641 nsew default input
rlabel metal4 s -2878 -2342 -2578 354310 4 vdda1
port 641 nsew default input
rlabel metal4 s 274002 -2812 274302 240 8 vdda1
port 641 nsew default input
rlabel metal4 s 256002 -2812 256302 240 8 vdda1
port 641 nsew default input
rlabel metal4 s 238002 -2812 238302 240 8 vdda1
port 641 nsew default input
rlabel metal4 s 220002 -2812 220302 240 8 vdda1
port 641 nsew default input
rlabel metal4 s 202002 -2812 202302 240 8 vdda1
port 641 nsew default input
rlabel metal4 s 184002 -2812 184302 240 8 vdda1
port 641 nsew default input
rlabel metal4 s 166002 -2812 166302 240 8 vdda1
port 641 nsew default input
rlabel metal4 s 148002 -2812 148302 240 8 vdda1
port 641 nsew default input
rlabel metal4 s 130002 -2812 130302 240 8 vdda1
port 641 nsew default input
rlabel metal4 s 112002 -2812 112302 240 8 vdda1
port 641 nsew default input
rlabel metal4 s 94002 -2812 94302 240 8 vdda1
port 641 nsew default input
rlabel metal4 s 76002 -2812 76302 240 8 vdda1
port 641 nsew default input
rlabel metal4 s 58002 -2812 58302 240 8 vdda1
port 641 nsew default input
rlabel metal4 s 40002 -2812 40302 240 8 vdda1
port 641 nsew default input
rlabel metal4 s 22002 -2812 22302 240 8 vdda1
port 641 nsew default input
rlabel metal4 s 4002 -2812 4302 240 8 vdda1
port 641 nsew default input
rlabel metal5 s -2878 354010 294840 354310 6 vdda1
port 641 nsew default input
rlabel metal5 s 291760 346538 295310 346838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 346538 240 346838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 328538 295310 328838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 328538 240 328838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 310538 295310 310838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 310538 240 310838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 292538 295310 292838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 292538 240 292838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 274538 295310 274838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 274538 240 274838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 256538 295310 256838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 256538 240 256838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 238538 295310 238838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 238538 240 238838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 220538 295310 220838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 220538 240 220838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 202538 295310 202838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 202538 240 202838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 184538 295310 184838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 184538 240 184838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 166538 295310 166838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 166538 240 166838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 148538 295310 148838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 148538 240 148838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 130538 295310 130838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 130538 240 130838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 112538 295310 112838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 112538 240 112838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 94538 295310 94838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 94538 240 94838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 76538 295310 76838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 76538 240 76838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 58538 295310 58838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 58538 240 58838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 40538 295310 40838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 40538 240 40838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 22538 295310 22838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 22538 240 22838 4 vdda1
port 641 nsew default input
rlabel metal5 s 291760 4538 295310 4838 6 vdda1
port 641 nsew default input
rlabel metal5 s -3348 4538 240 4838 4 vdda1
port 641 nsew default input
rlabel metal5 s -2878 -2342 294840 -2042 8 vdda1
port 641 nsew default input
rlabel metal4 s 295010 -2812 295310 354780 6 vssa1
port 642 nsew default input
rlabel metal4 s 283002 351760 283302 354780 6 vssa1
port 642 nsew default input
rlabel metal4 s 265002 351760 265302 354780 6 vssa1
port 642 nsew default input
rlabel metal4 s 247002 351760 247302 354780 6 vssa1
port 642 nsew default input
rlabel metal4 s 229002 351760 229302 354780 6 vssa1
port 642 nsew default input
rlabel metal4 s 211002 351760 211302 354780 6 vssa1
port 642 nsew default input
rlabel metal4 s 193002 351760 193302 354780 6 vssa1
port 642 nsew default input
rlabel metal4 s 175002 351760 175302 354780 6 vssa1
port 642 nsew default input
rlabel metal4 s 157002 351760 157302 354780 6 vssa1
port 642 nsew default input
rlabel metal4 s 139002 351760 139302 354780 6 vssa1
port 642 nsew default input
rlabel metal4 s 121002 351760 121302 354780 6 vssa1
port 642 nsew default input
rlabel metal4 s 103002 351760 103302 354780 6 vssa1
port 642 nsew default input
rlabel metal4 s 85002 351760 85302 354780 6 vssa1
port 642 nsew default input
rlabel metal4 s 67002 351760 67302 354780 6 vssa1
port 642 nsew default input
rlabel metal4 s 49002 351760 49302 354780 6 vssa1
port 642 nsew default input
rlabel metal4 s 31002 351760 31302 354780 6 vssa1
port 642 nsew default input
rlabel metal4 s 13002 351760 13302 354780 6 vssa1
port 642 nsew default input
rlabel metal4 s -3348 -2812 -3048 354780 4 vssa1
port 642 nsew default input
rlabel metal4 s 283002 -2812 283302 240 8 vssa1
port 642 nsew default input
rlabel metal4 s 265002 -2812 265302 240 8 vssa1
port 642 nsew default input
rlabel metal4 s 247002 -2812 247302 240 8 vssa1
port 642 nsew default input
rlabel metal4 s 229002 -2812 229302 240 8 vssa1
port 642 nsew default input
rlabel metal4 s 211002 -2812 211302 240 8 vssa1
port 642 nsew default input
rlabel metal4 s 193002 -2812 193302 240 8 vssa1
port 642 nsew default input
rlabel metal4 s 175002 -2812 175302 240 8 vssa1
port 642 nsew default input
rlabel metal4 s 157002 -2812 157302 240 8 vssa1
port 642 nsew default input
rlabel metal4 s 139002 -2812 139302 240 8 vssa1
port 642 nsew default input
rlabel metal4 s 121002 -2812 121302 240 8 vssa1
port 642 nsew default input
rlabel metal4 s 103002 -2812 103302 240 8 vssa1
port 642 nsew default input
rlabel metal4 s 85002 -2812 85302 240 8 vssa1
port 642 nsew default input
rlabel metal4 s 67002 -2812 67302 240 8 vssa1
port 642 nsew default input
rlabel metal4 s 49002 -2812 49302 240 8 vssa1
port 642 nsew default input
rlabel metal4 s 31002 -2812 31302 240 8 vssa1
port 642 nsew default input
rlabel metal4 s 13002 -2812 13302 240 8 vssa1
port 642 nsew default input
rlabel metal5 s -3348 354480 295310 354780 6 vssa1
port 642 nsew default input
rlabel metal5 s 291760 337538 295310 337838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 337538 240 337838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 319538 295310 319838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 319538 240 319838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 301538 295310 301838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 301538 240 301838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 283538 295310 283838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 283538 240 283838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 265538 295310 265838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 265538 240 265838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 247538 295310 247838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 247538 240 247838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 229538 295310 229838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 229538 240 229838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 211538 295310 211838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 211538 240 211838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 193538 295310 193838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 193538 240 193838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 175538 295310 175838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 175538 240 175838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 157538 295310 157838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 157538 240 157838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 139538 295310 139838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 139538 240 139838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 121538 295310 121838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 121538 240 121838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 103538 295310 103838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 103538 240 103838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 85538 295310 85838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 85538 240 85838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 67538 295310 67838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 67538 240 67838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 49538 295310 49838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 49538 240 49838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 31538 295310 31838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 31538 240 31838 4 vssa1
port 642 nsew default input
rlabel metal5 s 291760 13538 295310 13838 6 vssa1
port 642 nsew default input
rlabel metal5 s -3348 13538 240 13838 4 vssa1
port 642 nsew default input
rlabel metal5 s -3348 -2812 295310 -2512 8 vssa1
port 642 nsew default input
rlabel metal4 s 275802 351760 276102 355720 6 vdda2
port 643 nsew default input
rlabel metal4 s 257802 351760 258102 355720 6 vdda2
port 643 nsew default input
rlabel metal4 s 239802 351760 240102 355720 6 vdda2
port 643 nsew default input
rlabel metal4 s 221802 351760 222102 355720 6 vdda2
port 643 nsew default input
rlabel metal4 s 203802 351760 204102 355720 6 vdda2
port 643 nsew default input
rlabel metal4 s 185802 351760 186102 355720 6 vdda2
port 643 nsew default input
rlabel metal4 s 167802 351760 168102 355720 6 vdda2
port 643 nsew default input
rlabel metal4 s 149802 351760 150102 355720 6 vdda2
port 643 nsew default input
rlabel metal4 s 131802 351760 132102 355720 6 vdda2
port 643 nsew default input
rlabel metal4 s 113802 351760 114102 355720 6 vdda2
port 643 nsew default input
rlabel metal4 s 95802 351760 96102 355720 6 vdda2
port 643 nsew default input
rlabel metal4 s 77802 351760 78102 355720 6 vdda2
port 643 nsew default input
rlabel metal4 s 59802 351760 60102 355720 6 vdda2
port 643 nsew default input
rlabel metal4 s 41802 351760 42102 355720 6 vdda2
port 643 nsew default input
rlabel metal4 s 23802 351760 24102 355720 6 vdda2
port 643 nsew default input
rlabel metal4 s 5802 351760 6102 355720 6 vdda2
port 643 nsew default input
rlabel metal4 s 295480 -3282 295780 355250 6 vdda2
port 643 nsew default input
rlabel metal4 s -3818 -3282 -3518 355250 4 vdda2
port 643 nsew default input
rlabel metal4 s 275802 -3752 276102 240 8 vdda2
port 643 nsew default input
rlabel metal4 s 257802 -3752 258102 240 8 vdda2
port 643 nsew default input
rlabel metal4 s 239802 -3752 240102 240 8 vdda2
port 643 nsew default input
rlabel metal4 s 221802 -3752 222102 240 8 vdda2
port 643 nsew default input
rlabel metal4 s 203802 -3752 204102 240 8 vdda2
port 643 nsew default input
rlabel metal4 s 185802 -3752 186102 240 8 vdda2
port 643 nsew default input
rlabel metal4 s 167802 -3752 168102 240 8 vdda2
port 643 nsew default input
rlabel metal4 s 149802 -3752 150102 240 8 vdda2
port 643 nsew default input
rlabel metal4 s 131802 -3752 132102 240 8 vdda2
port 643 nsew default input
rlabel metal4 s 113802 -3752 114102 240 8 vdda2
port 643 nsew default input
rlabel metal4 s 95802 -3752 96102 240 8 vdda2
port 643 nsew default input
rlabel metal4 s 77802 -3752 78102 240 8 vdda2
port 643 nsew default input
rlabel metal4 s 59802 -3752 60102 240 8 vdda2
port 643 nsew default input
rlabel metal4 s 41802 -3752 42102 240 8 vdda2
port 643 nsew default input
rlabel metal4 s 23802 -3752 24102 240 8 vdda2
port 643 nsew default input
rlabel metal4 s 5802 -3752 6102 240 8 vdda2
port 643 nsew default input
rlabel metal5 s -3818 354950 295780 355250 6 vdda2
port 643 nsew default input
rlabel metal5 s 291760 348338 296250 348638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 348338 240 348638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 330338 296250 330638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 330338 240 330638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 312338 296250 312638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 312338 240 312638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 294338 296250 294638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 294338 240 294638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 276338 296250 276638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 276338 240 276638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 258338 296250 258638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 258338 240 258638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 240338 296250 240638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 240338 240 240638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 222338 296250 222638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 222338 240 222638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 204338 296250 204638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 204338 240 204638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 186338 296250 186638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 186338 240 186638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 168338 296250 168638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 168338 240 168638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 150338 296250 150638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 150338 240 150638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 132338 296250 132638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 132338 240 132638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 114338 296250 114638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 114338 240 114638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 96338 296250 96638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 96338 240 96638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 78338 296250 78638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 78338 240 78638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 60338 296250 60638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 60338 240 60638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 42338 296250 42638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 42338 240 42638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 24338 296250 24638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 24338 240 24638 4 vdda2
port 643 nsew default input
rlabel metal5 s 291760 6338 296250 6638 6 vdda2
port 643 nsew default input
rlabel metal5 s -4288 6338 240 6638 4 vdda2
port 643 nsew default input
rlabel metal5 s -3818 -3282 295780 -2982 8 vdda2
port 643 nsew default input
rlabel metal4 s 295950 -3752 296250 355720 6 vssa2
port 644 nsew default input
rlabel metal4 s 284802 351760 285102 355720 6 vssa2
port 644 nsew default input
rlabel metal4 s 266802 351760 267102 355720 6 vssa2
port 644 nsew default input
rlabel metal4 s 248802 351760 249102 355720 6 vssa2
port 644 nsew default input
rlabel metal4 s 230802 351760 231102 355720 6 vssa2
port 644 nsew default input
rlabel metal4 s 212802 351760 213102 355720 6 vssa2
port 644 nsew default input
rlabel metal4 s 194802 351760 195102 355720 6 vssa2
port 644 nsew default input
rlabel metal4 s 176802 351760 177102 355720 6 vssa2
port 644 nsew default input
rlabel metal4 s 158802 351760 159102 355720 6 vssa2
port 644 nsew default input
rlabel metal4 s 140802 351760 141102 355720 6 vssa2
port 644 nsew default input
rlabel metal4 s 122802 351760 123102 355720 6 vssa2
port 644 nsew default input
rlabel metal4 s 104802 351760 105102 355720 6 vssa2
port 644 nsew default input
rlabel metal4 s 86802 351760 87102 355720 6 vssa2
port 644 nsew default input
rlabel metal4 s 68802 351760 69102 355720 6 vssa2
port 644 nsew default input
rlabel metal4 s 50802 351760 51102 355720 6 vssa2
port 644 nsew default input
rlabel metal4 s 32802 351760 33102 355720 6 vssa2
port 644 nsew default input
rlabel metal4 s 14802 351760 15102 355720 6 vssa2
port 644 nsew default input
rlabel metal4 s -4288 -3752 -3988 355720 4 vssa2
port 644 nsew default input
rlabel metal4 s 284802 -3752 285102 240 8 vssa2
port 644 nsew default input
rlabel metal4 s 266802 -3752 267102 240 8 vssa2
port 644 nsew default input
rlabel metal4 s 248802 -3752 249102 240 8 vssa2
port 644 nsew default input
rlabel metal4 s 230802 -3752 231102 240 8 vssa2
port 644 nsew default input
rlabel metal4 s 212802 -3752 213102 240 8 vssa2
port 644 nsew default input
rlabel metal4 s 194802 -3752 195102 240 8 vssa2
port 644 nsew default input
rlabel metal4 s 176802 -3752 177102 240 8 vssa2
port 644 nsew default input
rlabel metal4 s 158802 -3752 159102 240 8 vssa2
port 644 nsew default input
rlabel metal4 s 140802 -3752 141102 240 8 vssa2
port 644 nsew default input
rlabel metal4 s 122802 -3752 123102 240 8 vssa2
port 644 nsew default input
rlabel metal4 s 104802 -3752 105102 240 8 vssa2
port 644 nsew default input
rlabel metal4 s 86802 -3752 87102 240 8 vssa2
port 644 nsew default input
rlabel metal4 s 68802 -3752 69102 240 8 vssa2
port 644 nsew default input
rlabel metal4 s 50802 -3752 51102 240 8 vssa2
port 644 nsew default input
rlabel metal4 s 32802 -3752 33102 240 8 vssa2
port 644 nsew default input
rlabel metal4 s 14802 -3752 15102 240 8 vssa2
port 644 nsew default input
rlabel metal5 s -4288 355420 296250 355720 6 vssa2
port 644 nsew default input
rlabel metal5 s 291760 339338 296250 339638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 339338 240 339638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 321338 296250 321638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 321338 240 321638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 303338 296250 303638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 303338 240 303638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 285338 296250 285638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 285338 240 285638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 267338 296250 267638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 267338 240 267638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 249338 296250 249638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 249338 240 249638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 231338 296250 231638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 231338 240 231638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 213338 296250 213638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 213338 240 213638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 195338 296250 195638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 195338 240 195638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 177338 296250 177638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 177338 240 177638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 159338 296250 159638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 159338 240 159638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 141338 296250 141638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 141338 240 141638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 123338 296250 123638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 123338 240 123638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 105338 296250 105638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 105338 240 105638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 87338 296250 87638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 87338 240 87638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 69338 296250 69638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 69338 240 69638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 51338 296250 51638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 51338 240 51638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 33338 296250 33638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 33338 240 33638 4 vssa2
port 644 nsew default input
rlabel metal5 s 291760 15338 296250 15638 6 vssa2
port 644 nsew default input
rlabel metal5 s -4288 15338 240 15638 4 vssa2
port 644 nsew default input
rlabel metal5 s -4288 -3752 296250 -3452 8 vssa2
port 644 nsew default input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 292000 352000
string GDS_FILE ../gds/user_project_wrapper.gds
string GDS_END 370014
string GDS_START 130
string LEFview TRUE
<< end >>
