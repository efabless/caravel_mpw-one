VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO digital_pll
  CLASS BLOCK ;
  FOREIGN digital_pll ;
  ORIGIN 0.000 0.000 ;
  SIZE 205.680 BY 205.200 ;
  PIN clockp[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 138.810 157.880 139.090 161.880 ;
        RECT 138.880 151.200 139.020 157.880 ;
    END
  END clockp[0]
  PIN clockp[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.520 48.120 108.660 54.000 ;
        RECT 108.450 44.120 108.730 48.120 ;
    END
  END clockp[1]
  PIN dco
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.600 48.120 61.740 54.000 ;
        RECT 61.530 44.120 61.810 48.120 ;
    END
  END dco
  PIN div[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 52.310 58.980 52.630 59.040 ;
        RECT 52.310 58.840 54.000 58.980 ;
        RECT 52.310 58.780 52.630 58.840 ;
      LAYER via ;
        RECT 52.340 58.780 52.600 59.040 ;
      LAYER met2 ;
        RECT 52.340 58.750 52.600 59.070 ;
        RECT 52.400 48.120 52.540 58.750 ;
        RECT 52.330 44.120 52.610 48.120 ;
    END
  END div[0]
  PIN div[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 89.490 53.480 89.640 ;
        RECT 49.480 89.190 54.000 89.490 ;
        RECT 49.480 89.040 53.480 89.190 ;
    END
  END div[1]
  PIN div[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.040 48.120 137.180 54.000 ;
        RECT 136.970 44.120 137.250 48.120 ;
    END
  END div[2]
  PIN div[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.880 52.805 139.020 54.000 ;
        RECT 138.810 52.435 139.090 52.805 ;
      LAYER via2 ;
        RECT 138.810 52.480 139.090 52.760 ;
      LAYER met3 ;
        RECT 138.785 52.770 139.115 52.785 ;
        RECT 152.520 52.770 156.520 52.920 ;
        RECT 138.785 52.470 156.520 52.770 ;
        RECT 138.785 52.455 139.115 52.470 ;
        RECT 152.520 52.320 156.520 52.470 ;
    END
  END div[3]
  PIN div[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 62.290 53.480 62.440 ;
        RECT 49.480 61.990 54.000 62.290 ;
        RECT 49.480 61.840 53.480 61.990 ;
    END
  END div[4]
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.090 157.880 101.370 161.880 ;
        RECT 101.160 151.200 101.300 157.880 ;
    END
  END enable
  PIN ext_trim[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.570 157.880 72.850 161.880 ;
        RECT 72.640 151.200 72.780 157.880 ;
    END
  END ext_trim[0]
  PIN ext_trim[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.490 157.880 119.770 161.880 ;
        RECT 119.560 151.200 119.700 157.880 ;
    END
  END ext_trim[10]
  PIN ext_trim[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 118.050 53.480 118.200 ;
        RECT 49.480 117.750 54.000 118.050 ;
        RECT 49.480 117.600 53.480 117.750 ;
    END
  END ext_trim[11]
  PIN ext_trim[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 152.520 66.370 156.520 66.520 ;
        RECT 151.680 66.070 156.520 66.370 ;
        RECT 152.520 65.920 156.520 66.070 ;
    END
  END ext_trim[12]
  PIN ext_trim[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 147.620 48.610 147.760 54.000 ;
        RECT 147.160 48.470 147.760 48.610 ;
        RECT 147.160 48.120 147.300 48.470 ;
        RECT 147.090 44.120 147.370 48.120 ;
    END
  END ext_trim[13]
  PIN ext_trim[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 104.450 53.480 104.600 ;
        RECT 49.480 104.150 54.000 104.450 ;
        RECT 49.480 104.000 53.480 104.150 ;
    END
  END ext_trim[14]
  PIN ext_trim[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.800 53.910 72.780 54.000 ;
        RECT 70.800 48.120 70.940 53.910 ;
        RECT 70.730 44.120 71.010 48.120 ;
    END
  END ext_trim[15]
  PIN ext_trim[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 152.520 137.090 156.520 137.240 ;
        RECT 151.680 136.790 156.520 137.090 ;
        RECT 152.520 136.640 156.520 136.790 ;
    END
  END ext_trim[16]
  PIN ext_trim[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 131.650 53.480 131.800 ;
        RECT 49.480 131.350 54.000 131.650 ;
        RECT 49.480 131.200 53.480 131.350 ;
    END
  END ext_trim[17]
  PIN ext_trim[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 148.010 157.880 148.290 161.880 ;
        RECT 148.080 151.200 148.220 157.880 ;
    END
  END ext_trim[18]
  PIN ext_trim[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.970 157.880 91.250 161.880 ;
        RECT 91.040 151.200 91.180 157.880 ;
    END
  END ext_trim[19]
  PIN ext_trim[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 152.520 123.490 156.520 123.640 ;
        RECT 151.680 123.190 156.520 123.490 ;
        RECT 152.520 123.040 156.520 123.190 ;
    END
  END ext_trim[1]
  PIN ext_trim[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 128.760 50.650 128.900 54.000 ;
        RECT 127.840 50.510 128.900 50.650 ;
        RECT 127.840 48.120 127.980 50.510 ;
        RECT 127.770 44.120 128.050 48.120 ;
    END
  END ext_trim[20]
  PIN ext_trim[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 146.610 53.480 146.760 ;
        RECT 49.480 146.310 54.000 146.610 ;
        RECT 49.480 146.160 53.480 146.310 ;
    END
  END ext_trim[21]
  PIN ext_trim[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 152.520 108.530 156.520 108.680 ;
        RECT 151.680 108.230 156.520 108.530 ;
        RECT 152.520 108.080 156.520 108.230 ;
    END
  END ext_trim[22]
  PIN ext_trim[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 49.480 75.890 53.480 76.040 ;
        RECT 49.480 75.590 54.000 75.890 ;
        RECT 49.480 75.440 53.480 75.590 ;
    END
  END ext_trim[23]
  PIN ext_trim[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 99.320 48.120 99.460 54.000 ;
        RECT 99.250 44.120 99.530 48.120 ;
    END
  END ext_trim[24]
  PIN ext_trim[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 152.520 81.330 156.520 81.480 ;
        RECT 151.680 81.030 156.520 81.330 ;
        RECT 152.520 80.880 156.520 81.030 ;
    END
  END ext_trim[25]
  PIN ext_trim[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 152.520 94.930 156.520 95.080 ;
        RECT 151.680 94.630 156.520 94.930 ;
        RECT 152.520 94.480 156.520 94.630 ;
    END
  END ext_trim[2]
  PIN ext_trim[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.450 157.880 62.730 161.880 ;
        RECT 62.520 151.200 62.660 157.880 ;
    END
  END ext_trim[3]
  PIN ext_trim[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.610 157.880 129.890 161.880 ;
        RECT 129.680 151.200 129.820 157.880 ;
    END
  END ext_trim[4]
  PIN ext_trim[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 118.640 48.120 118.780 54.000 ;
        RECT 118.570 44.120 118.850 48.120 ;
    END
  END ext_trim[5]
  PIN ext_trim[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.290 157.880 110.570 161.880 ;
        RECT 110.360 151.200 110.500 157.880 ;
    END
  END ext_trim[6]
  PIN ext_trim[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 53.230 143.640 53.550 143.700 ;
        RECT 53.230 143.500 54.000 143.640 ;
        RECT 53.230 143.440 53.550 143.500 ;
      LAYER via ;
        RECT 53.260 143.440 53.520 143.700 ;
      LAYER met2 ;
        RECT 53.250 157.880 53.530 161.880 ;
        RECT 53.320 143.730 53.460 157.880 ;
        RECT 53.260 143.410 53.520 143.730 ;
    END
  END ext_trim[7]
  PIN ext_trim[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.770 157.880 82.050 161.880 ;
        RECT 81.840 151.200 81.980 157.880 ;
    END
  END ext_trim[8]
  PIN ext_trim[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 152.520 150.690 156.520 150.840 ;
        RECT 151.680 150.390 156.520 150.690 ;
        RECT 152.520 150.240 156.520 150.390 ;
    END
  END ext_trim[9]
  PIN osc
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.120 48.120 90.260 54.000 ;
        RECT 90.050 44.120 90.330 48.120 ;
    END
  END osc
  PIN resetb
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 80.000 48.120 80.140 54.000 ;
        RECT 79.930 44.120 80.210 48.120 ;
    END
  END resetb
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 25.000 160.200 180.680 180.200 ;
        RECT 25.000 25.000 180.680 45.000 ;
      LAYER via3 ;
        RECT 25.040 179.840 25.360 180.160 ;
        RECT 25.440 179.840 25.760 180.160 ;
        RECT 25.840 179.840 26.160 180.160 ;
        RECT 26.240 179.840 26.560 180.160 ;
        RECT 26.640 179.840 26.960 180.160 ;
        RECT 27.040 179.840 27.360 180.160 ;
        RECT 27.440 179.840 27.760 180.160 ;
        RECT 27.840 179.840 28.160 180.160 ;
        RECT 28.240 179.840 28.560 180.160 ;
        RECT 28.640 179.840 28.960 180.160 ;
        RECT 29.040 179.840 29.360 180.160 ;
        RECT 29.440 179.840 29.760 180.160 ;
        RECT 29.840 179.840 30.160 180.160 ;
        RECT 30.240 179.840 30.560 180.160 ;
        RECT 30.640 179.840 30.960 180.160 ;
        RECT 31.040 179.840 31.360 180.160 ;
        RECT 31.440 179.840 31.760 180.160 ;
        RECT 31.840 179.840 32.160 180.160 ;
        RECT 32.240 179.840 32.560 180.160 ;
        RECT 32.640 179.840 32.960 180.160 ;
        RECT 33.040 179.840 33.360 180.160 ;
        RECT 33.440 179.840 33.760 180.160 ;
        RECT 33.840 179.840 34.160 180.160 ;
        RECT 34.240 179.840 34.560 180.160 ;
        RECT 34.640 179.840 34.960 180.160 ;
        RECT 35.040 179.840 35.360 180.160 ;
        RECT 35.440 179.840 35.760 180.160 ;
        RECT 35.840 179.840 36.160 180.160 ;
        RECT 36.240 179.840 36.560 180.160 ;
        RECT 36.640 179.840 36.960 180.160 ;
        RECT 37.040 179.840 37.360 180.160 ;
        RECT 37.440 179.840 37.760 180.160 ;
        RECT 37.840 179.840 38.160 180.160 ;
        RECT 38.240 179.840 38.560 180.160 ;
        RECT 38.640 179.840 38.960 180.160 ;
        RECT 39.040 179.840 39.360 180.160 ;
        RECT 39.440 179.840 39.760 180.160 ;
        RECT 39.840 179.840 40.160 180.160 ;
        RECT 40.240 179.840 40.560 180.160 ;
        RECT 40.640 179.840 40.960 180.160 ;
        RECT 41.040 179.840 41.360 180.160 ;
        RECT 41.440 179.840 41.760 180.160 ;
        RECT 41.840 179.840 42.160 180.160 ;
        RECT 42.240 179.840 42.560 180.160 ;
        RECT 42.640 179.840 42.960 180.160 ;
        RECT 43.040 179.840 43.360 180.160 ;
        RECT 43.440 179.840 43.760 180.160 ;
        RECT 43.840 179.840 44.160 180.160 ;
        RECT 44.240 179.840 44.560 180.160 ;
        RECT 44.640 179.840 44.960 180.160 ;
        RECT 70.560 179.840 70.880 180.160 ;
        RECT 70.960 179.840 71.280 180.160 ;
        RECT 71.360 179.840 71.680 180.160 ;
        RECT 71.760 179.840 72.080 180.160 ;
        RECT 120.560 179.840 120.880 180.160 ;
        RECT 120.960 179.840 121.280 180.160 ;
        RECT 121.360 179.840 121.680 180.160 ;
        RECT 121.760 179.840 122.080 180.160 ;
        RECT 160.720 179.840 161.040 180.160 ;
        RECT 161.120 179.840 161.440 180.160 ;
        RECT 161.520 179.840 161.840 180.160 ;
        RECT 161.920 179.840 162.240 180.160 ;
        RECT 162.320 179.840 162.640 180.160 ;
        RECT 162.720 179.840 163.040 180.160 ;
        RECT 163.120 179.840 163.440 180.160 ;
        RECT 163.520 179.840 163.840 180.160 ;
        RECT 163.920 179.840 164.240 180.160 ;
        RECT 164.320 179.840 164.640 180.160 ;
        RECT 164.720 179.840 165.040 180.160 ;
        RECT 165.120 179.840 165.440 180.160 ;
        RECT 165.520 179.840 165.840 180.160 ;
        RECT 165.920 179.840 166.240 180.160 ;
        RECT 166.320 179.840 166.640 180.160 ;
        RECT 166.720 179.840 167.040 180.160 ;
        RECT 167.120 179.840 167.440 180.160 ;
        RECT 167.520 179.840 167.840 180.160 ;
        RECT 167.920 179.840 168.240 180.160 ;
        RECT 168.320 179.840 168.640 180.160 ;
        RECT 168.720 179.840 169.040 180.160 ;
        RECT 169.120 179.840 169.440 180.160 ;
        RECT 169.520 179.840 169.840 180.160 ;
        RECT 169.920 179.840 170.240 180.160 ;
        RECT 170.320 179.840 170.640 180.160 ;
        RECT 170.720 179.840 171.040 180.160 ;
        RECT 171.120 179.840 171.440 180.160 ;
        RECT 171.520 179.840 171.840 180.160 ;
        RECT 171.920 179.840 172.240 180.160 ;
        RECT 172.320 179.840 172.640 180.160 ;
        RECT 172.720 179.840 173.040 180.160 ;
        RECT 173.120 179.840 173.440 180.160 ;
        RECT 173.520 179.840 173.840 180.160 ;
        RECT 173.920 179.840 174.240 180.160 ;
        RECT 174.320 179.840 174.640 180.160 ;
        RECT 174.720 179.840 175.040 180.160 ;
        RECT 175.120 179.840 175.440 180.160 ;
        RECT 175.520 179.840 175.840 180.160 ;
        RECT 175.920 179.840 176.240 180.160 ;
        RECT 176.320 179.840 176.640 180.160 ;
        RECT 176.720 179.840 177.040 180.160 ;
        RECT 177.120 179.840 177.440 180.160 ;
        RECT 177.520 179.840 177.840 180.160 ;
        RECT 177.920 179.840 178.240 180.160 ;
        RECT 178.320 179.840 178.640 180.160 ;
        RECT 178.720 179.840 179.040 180.160 ;
        RECT 179.120 179.840 179.440 180.160 ;
        RECT 179.520 179.840 179.840 180.160 ;
        RECT 179.920 179.840 180.240 180.160 ;
        RECT 180.320 179.840 180.640 180.160 ;
        RECT 25.040 179.440 25.360 179.760 ;
        RECT 25.440 179.440 25.760 179.760 ;
        RECT 25.840 179.440 26.160 179.760 ;
        RECT 26.240 179.440 26.560 179.760 ;
        RECT 26.640 179.440 26.960 179.760 ;
        RECT 27.040 179.440 27.360 179.760 ;
        RECT 27.440 179.440 27.760 179.760 ;
        RECT 27.840 179.440 28.160 179.760 ;
        RECT 28.240 179.440 28.560 179.760 ;
        RECT 28.640 179.440 28.960 179.760 ;
        RECT 29.040 179.440 29.360 179.760 ;
        RECT 29.440 179.440 29.760 179.760 ;
        RECT 29.840 179.440 30.160 179.760 ;
        RECT 30.240 179.440 30.560 179.760 ;
        RECT 30.640 179.440 30.960 179.760 ;
        RECT 31.040 179.440 31.360 179.760 ;
        RECT 31.440 179.440 31.760 179.760 ;
        RECT 31.840 179.440 32.160 179.760 ;
        RECT 32.240 179.440 32.560 179.760 ;
        RECT 32.640 179.440 32.960 179.760 ;
        RECT 33.040 179.440 33.360 179.760 ;
        RECT 33.440 179.440 33.760 179.760 ;
        RECT 33.840 179.440 34.160 179.760 ;
        RECT 34.240 179.440 34.560 179.760 ;
        RECT 34.640 179.440 34.960 179.760 ;
        RECT 35.040 179.440 35.360 179.760 ;
        RECT 35.440 179.440 35.760 179.760 ;
        RECT 35.840 179.440 36.160 179.760 ;
        RECT 36.240 179.440 36.560 179.760 ;
        RECT 36.640 179.440 36.960 179.760 ;
        RECT 37.040 179.440 37.360 179.760 ;
        RECT 37.440 179.440 37.760 179.760 ;
        RECT 37.840 179.440 38.160 179.760 ;
        RECT 38.240 179.440 38.560 179.760 ;
        RECT 38.640 179.440 38.960 179.760 ;
        RECT 39.040 179.440 39.360 179.760 ;
        RECT 39.440 179.440 39.760 179.760 ;
        RECT 39.840 179.440 40.160 179.760 ;
        RECT 40.240 179.440 40.560 179.760 ;
        RECT 40.640 179.440 40.960 179.760 ;
        RECT 41.040 179.440 41.360 179.760 ;
        RECT 41.440 179.440 41.760 179.760 ;
        RECT 41.840 179.440 42.160 179.760 ;
        RECT 42.240 179.440 42.560 179.760 ;
        RECT 42.640 179.440 42.960 179.760 ;
        RECT 43.040 179.440 43.360 179.760 ;
        RECT 43.440 179.440 43.760 179.760 ;
        RECT 43.840 179.440 44.160 179.760 ;
        RECT 44.240 179.440 44.560 179.760 ;
        RECT 44.640 179.440 44.960 179.760 ;
        RECT 70.560 179.440 70.880 179.760 ;
        RECT 70.960 179.440 71.280 179.760 ;
        RECT 71.360 179.440 71.680 179.760 ;
        RECT 71.760 179.440 72.080 179.760 ;
        RECT 120.560 179.440 120.880 179.760 ;
        RECT 120.960 179.440 121.280 179.760 ;
        RECT 121.360 179.440 121.680 179.760 ;
        RECT 121.760 179.440 122.080 179.760 ;
        RECT 160.720 179.440 161.040 179.760 ;
        RECT 161.120 179.440 161.440 179.760 ;
        RECT 161.520 179.440 161.840 179.760 ;
        RECT 161.920 179.440 162.240 179.760 ;
        RECT 162.320 179.440 162.640 179.760 ;
        RECT 162.720 179.440 163.040 179.760 ;
        RECT 163.120 179.440 163.440 179.760 ;
        RECT 163.520 179.440 163.840 179.760 ;
        RECT 163.920 179.440 164.240 179.760 ;
        RECT 164.320 179.440 164.640 179.760 ;
        RECT 164.720 179.440 165.040 179.760 ;
        RECT 165.120 179.440 165.440 179.760 ;
        RECT 165.520 179.440 165.840 179.760 ;
        RECT 165.920 179.440 166.240 179.760 ;
        RECT 166.320 179.440 166.640 179.760 ;
        RECT 166.720 179.440 167.040 179.760 ;
        RECT 167.120 179.440 167.440 179.760 ;
        RECT 167.520 179.440 167.840 179.760 ;
        RECT 167.920 179.440 168.240 179.760 ;
        RECT 168.320 179.440 168.640 179.760 ;
        RECT 168.720 179.440 169.040 179.760 ;
        RECT 169.120 179.440 169.440 179.760 ;
        RECT 169.520 179.440 169.840 179.760 ;
        RECT 169.920 179.440 170.240 179.760 ;
        RECT 170.320 179.440 170.640 179.760 ;
        RECT 170.720 179.440 171.040 179.760 ;
        RECT 171.120 179.440 171.440 179.760 ;
        RECT 171.520 179.440 171.840 179.760 ;
        RECT 171.920 179.440 172.240 179.760 ;
        RECT 172.320 179.440 172.640 179.760 ;
        RECT 172.720 179.440 173.040 179.760 ;
        RECT 173.120 179.440 173.440 179.760 ;
        RECT 173.520 179.440 173.840 179.760 ;
        RECT 173.920 179.440 174.240 179.760 ;
        RECT 174.320 179.440 174.640 179.760 ;
        RECT 174.720 179.440 175.040 179.760 ;
        RECT 175.120 179.440 175.440 179.760 ;
        RECT 175.520 179.440 175.840 179.760 ;
        RECT 175.920 179.440 176.240 179.760 ;
        RECT 176.320 179.440 176.640 179.760 ;
        RECT 176.720 179.440 177.040 179.760 ;
        RECT 177.120 179.440 177.440 179.760 ;
        RECT 177.520 179.440 177.840 179.760 ;
        RECT 177.920 179.440 178.240 179.760 ;
        RECT 178.320 179.440 178.640 179.760 ;
        RECT 178.720 179.440 179.040 179.760 ;
        RECT 179.120 179.440 179.440 179.760 ;
        RECT 179.520 179.440 179.840 179.760 ;
        RECT 179.920 179.440 180.240 179.760 ;
        RECT 180.320 179.440 180.640 179.760 ;
        RECT 25.040 179.040 25.360 179.360 ;
        RECT 25.440 179.040 25.760 179.360 ;
        RECT 25.840 179.040 26.160 179.360 ;
        RECT 26.240 179.040 26.560 179.360 ;
        RECT 26.640 179.040 26.960 179.360 ;
        RECT 27.040 179.040 27.360 179.360 ;
        RECT 27.440 179.040 27.760 179.360 ;
        RECT 27.840 179.040 28.160 179.360 ;
        RECT 28.240 179.040 28.560 179.360 ;
        RECT 28.640 179.040 28.960 179.360 ;
        RECT 29.040 179.040 29.360 179.360 ;
        RECT 29.440 179.040 29.760 179.360 ;
        RECT 29.840 179.040 30.160 179.360 ;
        RECT 30.240 179.040 30.560 179.360 ;
        RECT 30.640 179.040 30.960 179.360 ;
        RECT 31.040 179.040 31.360 179.360 ;
        RECT 31.440 179.040 31.760 179.360 ;
        RECT 31.840 179.040 32.160 179.360 ;
        RECT 32.240 179.040 32.560 179.360 ;
        RECT 32.640 179.040 32.960 179.360 ;
        RECT 33.040 179.040 33.360 179.360 ;
        RECT 33.440 179.040 33.760 179.360 ;
        RECT 33.840 179.040 34.160 179.360 ;
        RECT 34.240 179.040 34.560 179.360 ;
        RECT 34.640 179.040 34.960 179.360 ;
        RECT 35.040 179.040 35.360 179.360 ;
        RECT 35.440 179.040 35.760 179.360 ;
        RECT 35.840 179.040 36.160 179.360 ;
        RECT 36.240 179.040 36.560 179.360 ;
        RECT 36.640 179.040 36.960 179.360 ;
        RECT 37.040 179.040 37.360 179.360 ;
        RECT 37.440 179.040 37.760 179.360 ;
        RECT 37.840 179.040 38.160 179.360 ;
        RECT 38.240 179.040 38.560 179.360 ;
        RECT 38.640 179.040 38.960 179.360 ;
        RECT 39.040 179.040 39.360 179.360 ;
        RECT 39.440 179.040 39.760 179.360 ;
        RECT 39.840 179.040 40.160 179.360 ;
        RECT 40.240 179.040 40.560 179.360 ;
        RECT 40.640 179.040 40.960 179.360 ;
        RECT 41.040 179.040 41.360 179.360 ;
        RECT 41.440 179.040 41.760 179.360 ;
        RECT 41.840 179.040 42.160 179.360 ;
        RECT 42.240 179.040 42.560 179.360 ;
        RECT 42.640 179.040 42.960 179.360 ;
        RECT 43.040 179.040 43.360 179.360 ;
        RECT 43.440 179.040 43.760 179.360 ;
        RECT 43.840 179.040 44.160 179.360 ;
        RECT 44.240 179.040 44.560 179.360 ;
        RECT 44.640 179.040 44.960 179.360 ;
        RECT 70.560 179.040 70.880 179.360 ;
        RECT 70.960 179.040 71.280 179.360 ;
        RECT 71.360 179.040 71.680 179.360 ;
        RECT 71.760 179.040 72.080 179.360 ;
        RECT 120.560 179.040 120.880 179.360 ;
        RECT 120.960 179.040 121.280 179.360 ;
        RECT 121.360 179.040 121.680 179.360 ;
        RECT 121.760 179.040 122.080 179.360 ;
        RECT 160.720 179.040 161.040 179.360 ;
        RECT 161.120 179.040 161.440 179.360 ;
        RECT 161.520 179.040 161.840 179.360 ;
        RECT 161.920 179.040 162.240 179.360 ;
        RECT 162.320 179.040 162.640 179.360 ;
        RECT 162.720 179.040 163.040 179.360 ;
        RECT 163.120 179.040 163.440 179.360 ;
        RECT 163.520 179.040 163.840 179.360 ;
        RECT 163.920 179.040 164.240 179.360 ;
        RECT 164.320 179.040 164.640 179.360 ;
        RECT 164.720 179.040 165.040 179.360 ;
        RECT 165.120 179.040 165.440 179.360 ;
        RECT 165.520 179.040 165.840 179.360 ;
        RECT 165.920 179.040 166.240 179.360 ;
        RECT 166.320 179.040 166.640 179.360 ;
        RECT 166.720 179.040 167.040 179.360 ;
        RECT 167.120 179.040 167.440 179.360 ;
        RECT 167.520 179.040 167.840 179.360 ;
        RECT 167.920 179.040 168.240 179.360 ;
        RECT 168.320 179.040 168.640 179.360 ;
        RECT 168.720 179.040 169.040 179.360 ;
        RECT 169.120 179.040 169.440 179.360 ;
        RECT 169.520 179.040 169.840 179.360 ;
        RECT 169.920 179.040 170.240 179.360 ;
        RECT 170.320 179.040 170.640 179.360 ;
        RECT 170.720 179.040 171.040 179.360 ;
        RECT 171.120 179.040 171.440 179.360 ;
        RECT 171.520 179.040 171.840 179.360 ;
        RECT 171.920 179.040 172.240 179.360 ;
        RECT 172.320 179.040 172.640 179.360 ;
        RECT 172.720 179.040 173.040 179.360 ;
        RECT 173.120 179.040 173.440 179.360 ;
        RECT 173.520 179.040 173.840 179.360 ;
        RECT 173.920 179.040 174.240 179.360 ;
        RECT 174.320 179.040 174.640 179.360 ;
        RECT 174.720 179.040 175.040 179.360 ;
        RECT 175.120 179.040 175.440 179.360 ;
        RECT 175.520 179.040 175.840 179.360 ;
        RECT 175.920 179.040 176.240 179.360 ;
        RECT 176.320 179.040 176.640 179.360 ;
        RECT 176.720 179.040 177.040 179.360 ;
        RECT 177.120 179.040 177.440 179.360 ;
        RECT 177.520 179.040 177.840 179.360 ;
        RECT 177.920 179.040 178.240 179.360 ;
        RECT 178.320 179.040 178.640 179.360 ;
        RECT 178.720 179.040 179.040 179.360 ;
        RECT 179.120 179.040 179.440 179.360 ;
        RECT 179.520 179.040 179.840 179.360 ;
        RECT 179.920 179.040 180.240 179.360 ;
        RECT 180.320 179.040 180.640 179.360 ;
        RECT 25.040 178.640 25.360 178.960 ;
        RECT 25.440 178.640 25.760 178.960 ;
        RECT 25.840 178.640 26.160 178.960 ;
        RECT 26.240 178.640 26.560 178.960 ;
        RECT 26.640 178.640 26.960 178.960 ;
        RECT 27.040 178.640 27.360 178.960 ;
        RECT 27.440 178.640 27.760 178.960 ;
        RECT 27.840 178.640 28.160 178.960 ;
        RECT 28.240 178.640 28.560 178.960 ;
        RECT 28.640 178.640 28.960 178.960 ;
        RECT 29.040 178.640 29.360 178.960 ;
        RECT 29.440 178.640 29.760 178.960 ;
        RECT 29.840 178.640 30.160 178.960 ;
        RECT 30.240 178.640 30.560 178.960 ;
        RECT 30.640 178.640 30.960 178.960 ;
        RECT 31.040 178.640 31.360 178.960 ;
        RECT 31.440 178.640 31.760 178.960 ;
        RECT 31.840 178.640 32.160 178.960 ;
        RECT 32.240 178.640 32.560 178.960 ;
        RECT 32.640 178.640 32.960 178.960 ;
        RECT 33.040 178.640 33.360 178.960 ;
        RECT 33.440 178.640 33.760 178.960 ;
        RECT 33.840 178.640 34.160 178.960 ;
        RECT 34.240 178.640 34.560 178.960 ;
        RECT 34.640 178.640 34.960 178.960 ;
        RECT 35.040 178.640 35.360 178.960 ;
        RECT 35.440 178.640 35.760 178.960 ;
        RECT 35.840 178.640 36.160 178.960 ;
        RECT 36.240 178.640 36.560 178.960 ;
        RECT 36.640 178.640 36.960 178.960 ;
        RECT 37.040 178.640 37.360 178.960 ;
        RECT 37.440 178.640 37.760 178.960 ;
        RECT 37.840 178.640 38.160 178.960 ;
        RECT 38.240 178.640 38.560 178.960 ;
        RECT 38.640 178.640 38.960 178.960 ;
        RECT 39.040 178.640 39.360 178.960 ;
        RECT 39.440 178.640 39.760 178.960 ;
        RECT 39.840 178.640 40.160 178.960 ;
        RECT 40.240 178.640 40.560 178.960 ;
        RECT 40.640 178.640 40.960 178.960 ;
        RECT 41.040 178.640 41.360 178.960 ;
        RECT 41.440 178.640 41.760 178.960 ;
        RECT 41.840 178.640 42.160 178.960 ;
        RECT 42.240 178.640 42.560 178.960 ;
        RECT 42.640 178.640 42.960 178.960 ;
        RECT 43.040 178.640 43.360 178.960 ;
        RECT 43.440 178.640 43.760 178.960 ;
        RECT 43.840 178.640 44.160 178.960 ;
        RECT 44.240 178.640 44.560 178.960 ;
        RECT 44.640 178.640 44.960 178.960 ;
        RECT 70.560 178.640 70.880 178.960 ;
        RECT 70.960 178.640 71.280 178.960 ;
        RECT 71.360 178.640 71.680 178.960 ;
        RECT 71.760 178.640 72.080 178.960 ;
        RECT 120.560 178.640 120.880 178.960 ;
        RECT 120.960 178.640 121.280 178.960 ;
        RECT 121.360 178.640 121.680 178.960 ;
        RECT 121.760 178.640 122.080 178.960 ;
        RECT 160.720 178.640 161.040 178.960 ;
        RECT 161.120 178.640 161.440 178.960 ;
        RECT 161.520 178.640 161.840 178.960 ;
        RECT 161.920 178.640 162.240 178.960 ;
        RECT 162.320 178.640 162.640 178.960 ;
        RECT 162.720 178.640 163.040 178.960 ;
        RECT 163.120 178.640 163.440 178.960 ;
        RECT 163.520 178.640 163.840 178.960 ;
        RECT 163.920 178.640 164.240 178.960 ;
        RECT 164.320 178.640 164.640 178.960 ;
        RECT 164.720 178.640 165.040 178.960 ;
        RECT 165.120 178.640 165.440 178.960 ;
        RECT 165.520 178.640 165.840 178.960 ;
        RECT 165.920 178.640 166.240 178.960 ;
        RECT 166.320 178.640 166.640 178.960 ;
        RECT 166.720 178.640 167.040 178.960 ;
        RECT 167.120 178.640 167.440 178.960 ;
        RECT 167.520 178.640 167.840 178.960 ;
        RECT 167.920 178.640 168.240 178.960 ;
        RECT 168.320 178.640 168.640 178.960 ;
        RECT 168.720 178.640 169.040 178.960 ;
        RECT 169.120 178.640 169.440 178.960 ;
        RECT 169.520 178.640 169.840 178.960 ;
        RECT 169.920 178.640 170.240 178.960 ;
        RECT 170.320 178.640 170.640 178.960 ;
        RECT 170.720 178.640 171.040 178.960 ;
        RECT 171.120 178.640 171.440 178.960 ;
        RECT 171.520 178.640 171.840 178.960 ;
        RECT 171.920 178.640 172.240 178.960 ;
        RECT 172.320 178.640 172.640 178.960 ;
        RECT 172.720 178.640 173.040 178.960 ;
        RECT 173.120 178.640 173.440 178.960 ;
        RECT 173.520 178.640 173.840 178.960 ;
        RECT 173.920 178.640 174.240 178.960 ;
        RECT 174.320 178.640 174.640 178.960 ;
        RECT 174.720 178.640 175.040 178.960 ;
        RECT 175.120 178.640 175.440 178.960 ;
        RECT 175.520 178.640 175.840 178.960 ;
        RECT 175.920 178.640 176.240 178.960 ;
        RECT 176.320 178.640 176.640 178.960 ;
        RECT 176.720 178.640 177.040 178.960 ;
        RECT 177.120 178.640 177.440 178.960 ;
        RECT 177.520 178.640 177.840 178.960 ;
        RECT 177.920 178.640 178.240 178.960 ;
        RECT 178.320 178.640 178.640 178.960 ;
        RECT 178.720 178.640 179.040 178.960 ;
        RECT 179.120 178.640 179.440 178.960 ;
        RECT 179.520 178.640 179.840 178.960 ;
        RECT 179.920 178.640 180.240 178.960 ;
        RECT 180.320 178.640 180.640 178.960 ;
        RECT 25.040 178.240 25.360 178.560 ;
        RECT 25.440 178.240 25.760 178.560 ;
        RECT 25.840 178.240 26.160 178.560 ;
        RECT 26.240 178.240 26.560 178.560 ;
        RECT 26.640 178.240 26.960 178.560 ;
        RECT 27.040 178.240 27.360 178.560 ;
        RECT 27.440 178.240 27.760 178.560 ;
        RECT 27.840 178.240 28.160 178.560 ;
        RECT 28.240 178.240 28.560 178.560 ;
        RECT 28.640 178.240 28.960 178.560 ;
        RECT 29.040 178.240 29.360 178.560 ;
        RECT 29.440 178.240 29.760 178.560 ;
        RECT 29.840 178.240 30.160 178.560 ;
        RECT 30.240 178.240 30.560 178.560 ;
        RECT 30.640 178.240 30.960 178.560 ;
        RECT 31.040 178.240 31.360 178.560 ;
        RECT 31.440 178.240 31.760 178.560 ;
        RECT 31.840 178.240 32.160 178.560 ;
        RECT 32.240 178.240 32.560 178.560 ;
        RECT 32.640 178.240 32.960 178.560 ;
        RECT 33.040 178.240 33.360 178.560 ;
        RECT 33.440 178.240 33.760 178.560 ;
        RECT 33.840 178.240 34.160 178.560 ;
        RECT 34.240 178.240 34.560 178.560 ;
        RECT 34.640 178.240 34.960 178.560 ;
        RECT 35.040 178.240 35.360 178.560 ;
        RECT 35.440 178.240 35.760 178.560 ;
        RECT 35.840 178.240 36.160 178.560 ;
        RECT 36.240 178.240 36.560 178.560 ;
        RECT 36.640 178.240 36.960 178.560 ;
        RECT 37.040 178.240 37.360 178.560 ;
        RECT 37.440 178.240 37.760 178.560 ;
        RECT 37.840 178.240 38.160 178.560 ;
        RECT 38.240 178.240 38.560 178.560 ;
        RECT 38.640 178.240 38.960 178.560 ;
        RECT 39.040 178.240 39.360 178.560 ;
        RECT 39.440 178.240 39.760 178.560 ;
        RECT 39.840 178.240 40.160 178.560 ;
        RECT 40.240 178.240 40.560 178.560 ;
        RECT 40.640 178.240 40.960 178.560 ;
        RECT 41.040 178.240 41.360 178.560 ;
        RECT 41.440 178.240 41.760 178.560 ;
        RECT 41.840 178.240 42.160 178.560 ;
        RECT 42.240 178.240 42.560 178.560 ;
        RECT 42.640 178.240 42.960 178.560 ;
        RECT 43.040 178.240 43.360 178.560 ;
        RECT 43.440 178.240 43.760 178.560 ;
        RECT 43.840 178.240 44.160 178.560 ;
        RECT 44.240 178.240 44.560 178.560 ;
        RECT 44.640 178.240 44.960 178.560 ;
        RECT 70.560 178.240 70.880 178.560 ;
        RECT 70.960 178.240 71.280 178.560 ;
        RECT 71.360 178.240 71.680 178.560 ;
        RECT 71.760 178.240 72.080 178.560 ;
        RECT 120.560 178.240 120.880 178.560 ;
        RECT 120.960 178.240 121.280 178.560 ;
        RECT 121.360 178.240 121.680 178.560 ;
        RECT 121.760 178.240 122.080 178.560 ;
        RECT 160.720 178.240 161.040 178.560 ;
        RECT 161.120 178.240 161.440 178.560 ;
        RECT 161.520 178.240 161.840 178.560 ;
        RECT 161.920 178.240 162.240 178.560 ;
        RECT 162.320 178.240 162.640 178.560 ;
        RECT 162.720 178.240 163.040 178.560 ;
        RECT 163.120 178.240 163.440 178.560 ;
        RECT 163.520 178.240 163.840 178.560 ;
        RECT 163.920 178.240 164.240 178.560 ;
        RECT 164.320 178.240 164.640 178.560 ;
        RECT 164.720 178.240 165.040 178.560 ;
        RECT 165.120 178.240 165.440 178.560 ;
        RECT 165.520 178.240 165.840 178.560 ;
        RECT 165.920 178.240 166.240 178.560 ;
        RECT 166.320 178.240 166.640 178.560 ;
        RECT 166.720 178.240 167.040 178.560 ;
        RECT 167.120 178.240 167.440 178.560 ;
        RECT 167.520 178.240 167.840 178.560 ;
        RECT 167.920 178.240 168.240 178.560 ;
        RECT 168.320 178.240 168.640 178.560 ;
        RECT 168.720 178.240 169.040 178.560 ;
        RECT 169.120 178.240 169.440 178.560 ;
        RECT 169.520 178.240 169.840 178.560 ;
        RECT 169.920 178.240 170.240 178.560 ;
        RECT 170.320 178.240 170.640 178.560 ;
        RECT 170.720 178.240 171.040 178.560 ;
        RECT 171.120 178.240 171.440 178.560 ;
        RECT 171.520 178.240 171.840 178.560 ;
        RECT 171.920 178.240 172.240 178.560 ;
        RECT 172.320 178.240 172.640 178.560 ;
        RECT 172.720 178.240 173.040 178.560 ;
        RECT 173.120 178.240 173.440 178.560 ;
        RECT 173.520 178.240 173.840 178.560 ;
        RECT 173.920 178.240 174.240 178.560 ;
        RECT 174.320 178.240 174.640 178.560 ;
        RECT 174.720 178.240 175.040 178.560 ;
        RECT 175.120 178.240 175.440 178.560 ;
        RECT 175.520 178.240 175.840 178.560 ;
        RECT 175.920 178.240 176.240 178.560 ;
        RECT 176.320 178.240 176.640 178.560 ;
        RECT 176.720 178.240 177.040 178.560 ;
        RECT 177.120 178.240 177.440 178.560 ;
        RECT 177.520 178.240 177.840 178.560 ;
        RECT 177.920 178.240 178.240 178.560 ;
        RECT 178.320 178.240 178.640 178.560 ;
        RECT 178.720 178.240 179.040 178.560 ;
        RECT 179.120 178.240 179.440 178.560 ;
        RECT 179.520 178.240 179.840 178.560 ;
        RECT 179.920 178.240 180.240 178.560 ;
        RECT 180.320 178.240 180.640 178.560 ;
        RECT 25.040 177.840 25.360 178.160 ;
        RECT 25.440 177.840 25.760 178.160 ;
        RECT 25.840 177.840 26.160 178.160 ;
        RECT 26.240 177.840 26.560 178.160 ;
        RECT 26.640 177.840 26.960 178.160 ;
        RECT 27.040 177.840 27.360 178.160 ;
        RECT 27.440 177.840 27.760 178.160 ;
        RECT 27.840 177.840 28.160 178.160 ;
        RECT 28.240 177.840 28.560 178.160 ;
        RECT 28.640 177.840 28.960 178.160 ;
        RECT 29.040 177.840 29.360 178.160 ;
        RECT 29.440 177.840 29.760 178.160 ;
        RECT 29.840 177.840 30.160 178.160 ;
        RECT 30.240 177.840 30.560 178.160 ;
        RECT 30.640 177.840 30.960 178.160 ;
        RECT 31.040 177.840 31.360 178.160 ;
        RECT 31.440 177.840 31.760 178.160 ;
        RECT 31.840 177.840 32.160 178.160 ;
        RECT 32.240 177.840 32.560 178.160 ;
        RECT 32.640 177.840 32.960 178.160 ;
        RECT 33.040 177.840 33.360 178.160 ;
        RECT 33.440 177.840 33.760 178.160 ;
        RECT 33.840 177.840 34.160 178.160 ;
        RECT 34.240 177.840 34.560 178.160 ;
        RECT 34.640 177.840 34.960 178.160 ;
        RECT 35.040 177.840 35.360 178.160 ;
        RECT 35.440 177.840 35.760 178.160 ;
        RECT 35.840 177.840 36.160 178.160 ;
        RECT 36.240 177.840 36.560 178.160 ;
        RECT 36.640 177.840 36.960 178.160 ;
        RECT 37.040 177.840 37.360 178.160 ;
        RECT 37.440 177.840 37.760 178.160 ;
        RECT 37.840 177.840 38.160 178.160 ;
        RECT 38.240 177.840 38.560 178.160 ;
        RECT 38.640 177.840 38.960 178.160 ;
        RECT 39.040 177.840 39.360 178.160 ;
        RECT 39.440 177.840 39.760 178.160 ;
        RECT 39.840 177.840 40.160 178.160 ;
        RECT 40.240 177.840 40.560 178.160 ;
        RECT 40.640 177.840 40.960 178.160 ;
        RECT 41.040 177.840 41.360 178.160 ;
        RECT 41.440 177.840 41.760 178.160 ;
        RECT 41.840 177.840 42.160 178.160 ;
        RECT 42.240 177.840 42.560 178.160 ;
        RECT 42.640 177.840 42.960 178.160 ;
        RECT 43.040 177.840 43.360 178.160 ;
        RECT 43.440 177.840 43.760 178.160 ;
        RECT 43.840 177.840 44.160 178.160 ;
        RECT 44.240 177.840 44.560 178.160 ;
        RECT 44.640 177.840 44.960 178.160 ;
        RECT 70.560 177.840 70.880 178.160 ;
        RECT 70.960 177.840 71.280 178.160 ;
        RECT 71.360 177.840 71.680 178.160 ;
        RECT 71.760 177.840 72.080 178.160 ;
        RECT 120.560 177.840 120.880 178.160 ;
        RECT 120.960 177.840 121.280 178.160 ;
        RECT 121.360 177.840 121.680 178.160 ;
        RECT 121.760 177.840 122.080 178.160 ;
        RECT 160.720 177.840 161.040 178.160 ;
        RECT 161.120 177.840 161.440 178.160 ;
        RECT 161.520 177.840 161.840 178.160 ;
        RECT 161.920 177.840 162.240 178.160 ;
        RECT 162.320 177.840 162.640 178.160 ;
        RECT 162.720 177.840 163.040 178.160 ;
        RECT 163.120 177.840 163.440 178.160 ;
        RECT 163.520 177.840 163.840 178.160 ;
        RECT 163.920 177.840 164.240 178.160 ;
        RECT 164.320 177.840 164.640 178.160 ;
        RECT 164.720 177.840 165.040 178.160 ;
        RECT 165.120 177.840 165.440 178.160 ;
        RECT 165.520 177.840 165.840 178.160 ;
        RECT 165.920 177.840 166.240 178.160 ;
        RECT 166.320 177.840 166.640 178.160 ;
        RECT 166.720 177.840 167.040 178.160 ;
        RECT 167.120 177.840 167.440 178.160 ;
        RECT 167.520 177.840 167.840 178.160 ;
        RECT 167.920 177.840 168.240 178.160 ;
        RECT 168.320 177.840 168.640 178.160 ;
        RECT 168.720 177.840 169.040 178.160 ;
        RECT 169.120 177.840 169.440 178.160 ;
        RECT 169.520 177.840 169.840 178.160 ;
        RECT 169.920 177.840 170.240 178.160 ;
        RECT 170.320 177.840 170.640 178.160 ;
        RECT 170.720 177.840 171.040 178.160 ;
        RECT 171.120 177.840 171.440 178.160 ;
        RECT 171.520 177.840 171.840 178.160 ;
        RECT 171.920 177.840 172.240 178.160 ;
        RECT 172.320 177.840 172.640 178.160 ;
        RECT 172.720 177.840 173.040 178.160 ;
        RECT 173.120 177.840 173.440 178.160 ;
        RECT 173.520 177.840 173.840 178.160 ;
        RECT 173.920 177.840 174.240 178.160 ;
        RECT 174.320 177.840 174.640 178.160 ;
        RECT 174.720 177.840 175.040 178.160 ;
        RECT 175.120 177.840 175.440 178.160 ;
        RECT 175.520 177.840 175.840 178.160 ;
        RECT 175.920 177.840 176.240 178.160 ;
        RECT 176.320 177.840 176.640 178.160 ;
        RECT 176.720 177.840 177.040 178.160 ;
        RECT 177.120 177.840 177.440 178.160 ;
        RECT 177.520 177.840 177.840 178.160 ;
        RECT 177.920 177.840 178.240 178.160 ;
        RECT 178.320 177.840 178.640 178.160 ;
        RECT 178.720 177.840 179.040 178.160 ;
        RECT 179.120 177.840 179.440 178.160 ;
        RECT 179.520 177.840 179.840 178.160 ;
        RECT 179.920 177.840 180.240 178.160 ;
        RECT 180.320 177.840 180.640 178.160 ;
        RECT 25.040 177.440 25.360 177.760 ;
        RECT 25.440 177.440 25.760 177.760 ;
        RECT 25.840 177.440 26.160 177.760 ;
        RECT 26.240 177.440 26.560 177.760 ;
        RECT 26.640 177.440 26.960 177.760 ;
        RECT 27.040 177.440 27.360 177.760 ;
        RECT 27.440 177.440 27.760 177.760 ;
        RECT 27.840 177.440 28.160 177.760 ;
        RECT 28.240 177.440 28.560 177.760 ;
        RECT 28.640 177.440 28.960 177.760 ;
        RECT 29.040 177.440 29.360 177.760 ;
        RECT 29.440 177.440 29.760 177.760 ;
        RECT 29.840 177.440 30.160 177.760 ;
        RECT 30.240 177.440 30.560 177.760 ;
        RECT 30.640 177.440 30.960 177.760 ;
        RECT 31.040 177.440 31.360 177.760 ;
        RECT 31.440 177.440 31.760 177.760 ;
        RECT 31.840 177.440 32.160 177.760 ;
        RECT 32.240 177.440 32.560 177.760 ;
        RECT 32.640 177.440 32.960 177.760 ;
        RECT 33.040 177.440 33.360 177.760 ;
        RECT 33.440 177.440 33.760 177.760 ;
        RECT 33.840 177.440 34.160 177.760 ;
        RECT 34.240 177.440 34.560 177.760 ;
        RECT 34.640 177.440 34.960 177.760 ;
        RECT 35.040 177.440 35.360 177.760 ;
        RECT 35.440 177.440 35.760 177.760 ;
        RECT 35.840 177.440 36.160 177.760 ;
        RECT 36.240 177.440 36.560 177.760 ;
        RECT 36.640 177.440 36.960 177.760 ;
        RECT 37.040 177.440 37.360 177.760 ;
        RECT 37.440 177.440 37.760 177.760 ;
        RECT 37.840 177.440 38.160 177.760 ;
        RECT 38.240 177.440 38.560 177.760 ;
        RECT 38.640 177.440 38.960 177.760 ;
        RECT 39.040 177.440 39.360 177.760 ;
        RECT 39.440 177.440 39.760 177.760 ;
        RECT 39.840 177.440 40.160 177.760 ;
        RECT 40.240 177.440 40.560 177.760 ;
        RECT 40.640 177.440 40.960 177.760 ;
        RECT 41.040 177.440 41.360 177.760 ;
        RECT 41.440 177.440 41.760 177.760 ;
        RECT 41.840 177.440 42.160 177.760 ;
        RECT 42.240 177.440 42.560 177.760 ;
        RECT 42.640 177.440 42.960 177.760 ;
        RECT 43.040 177.440 43.360 177.760 ;
        RECT 43.440 177.440 43.760 177.760 ;
        RECT 43.840 177.440 44.160 177.760 ;
        RECT 44.240 177.440 44.560 177.760 ;
        RECT 44.640 177.440 44.960 177.760 ;
        RECT 70.560 177.440 70.880 177.760 ;
        RECT 70.960 177.440 71.280 177.760 ;
        RECT 71.360 177.440 71.680 177.760 ;
        RECT 71.760 177.440 72.080 177.760 ;
        RECT 120.560 177.440 120.880 177.760 ;
        RECT 120.960 177.440 121.280 177.760 ;
        RECT 121.360 177.440 121.680 177.760 ;
        RECT 121.760 177.440 122.080 177.760 ;
        RECT 160.720 177.440 161.040 177.760 ;
        RECT 161.120 177.440 161.440 177.760 ;
        RECT 161.520 177.440 161.840 177.760 ;
        RECT 161.920 177.440 162.240 177.760 ;
        RECT 162.320 177.440 162.640 177.760 ;
        RECT 162.720 177.440 163.040 177.760 ;
        RECT 163.120 177.440 163.440 177.760 ;
        RECT 163.520 177.440 163.840 177.760 ;
        RECT 163.920 177.440 164.240 177.760 ;
        RECT 164.320 177.440 164.640 177.760 ;
        RECT 164.720 177.440 165.040 177.760 ;
        RECT 165.120 177.440 165.440 177.760 ;
        RECT 165.520 177.440 165.840 177.760 ;
        RECT 165.920 177.440 166.240 177.760 ;
        RECT 166.320 177.440 166.640 177.760 ;
        RECT 166.720 177.440 167.040 177.760 ;
        RECT 167.120 177.440 167.440 177.760 ;
        RECT 167.520 177.440 167.840 177.760 ;
        RECT 167.920 177.440 168.240 177.760 ;
        RECT 168.320 177.440 168.640 177.760 ;
        RECT 168.720 177.440 169.040 177.760 ;
        RECT 169.120 177.440 169.440 177.760 ;
        RECT 169.520 177.440 169.840 177.760 ;
        RECT 169.920 177.440 170.240 177.760 ;
        RECT 170.320 177.440 170.640 177.760 ;
        RECT 170.720 177.440 171.040 177.760 ;
        RECT 171.120 177.440 171.440 177.760 ;
        RECT 171.520 177.440 171.840 177.760 ;
        RECT 171.920 177.440 172.240 177.760 ;
        RECT 172.320 177.440 172.640 177.760 ;
        RECT 172.720 177.440 173.040 177.760 ;
        RECT 173.120 177.440 173.440 177.760 ;
        RECT 173.520 177.440 173.840 177.760 ;
        RECT 173.920 177.440 174.240 177.760 ;
        RECT 174.320 177.440 174.640 177.760 ;
        RECT 174.720 177.440 175.040 177.760 ;
        RECT 175.120 177.440 175.440 177.760 ;
        RECT 175.520 177.440 175.840 177.760 ;
        RECT 175.920 177.440 176.240 177.760 ;
        RECT 176.320 177.440 176.640 177.760 ;
        RECT 176.720 177.440 177.040 177.760 ;
        RECT 177.120 177.440 177.440 177.760 ;
        RECT 177.520 177.440 177.840 177.760 ;
        RECT 177.920 177.440 178.240 177.760 ;
        RECT 178.320 177.440 178.640 177.760 ;
        RECT 178.720 177.440 179.040 177.760 ;
        RECT 179.120 177.440 179.440 177.760 ;
        RECT 179.520 177.440 179.840 177.760 ;
        RECT 179.920 177.440 180.240 177.760 ;
        RECT 180.320 177.440 180.640 177.760 ;
        RECT 25.040 177.040 25.360 177.360 ;
        RECT 25.440 177.040 25.760 177.360 ;
        RECT 25.840 177.040 26.160 177.360 ;
        RECT 26.240 177.040 26.560 177.360 ;
        RECT 26.640 177.040 26.960 177.360 ;
        RECT 27.040 177.040 27.360 177.360 ;
        RECT 27.440 177.040 27.760 177.360 ;
        RECT 27.840 177.040 28.160 177.360 ;
        RECT 28.240 177.040 28.560 177.360 ;
        RECT 28.640 177.040 28.960 177.360 ;
        RECT 29.040 177.040 29.360 177.360 ;
        RECT 29.440 177.040 29.760 177.360 ;
        RECT 29.840 177.040 30.160 177.360 ;
        RECT 30.240 177.040 30.560 177.360 ;
        RECT 30.640 177.040 30.960 177.360 ;
        RECT 31.040 177.040 31.360 177.360 ;
        RECT 31.440 177.040 31.760 177.360 ;
        RECT 31.840 177.040 32.160 177.360 ;
        RECT 32.240 177.040 32.560 177.360 ;
        RECT 32.640 177.040 32.960 177.360 ;
        RECT 33.040 177.040 33.360 177.360 ;
        RECT 33.440 177.040 33.760 177.360 ;
        RECT 33.840 177.040 34.160 177.360 ;
        RECT 34.240 177.040 34.560 177.360 ;
        RECT 34.640 177.040 34.960 177.360 ;
        RECT 35.040 177.040 35.360 177.360 ;
        RECT 35.440 177.040 35.760 177.360 ;
        RECT 35.840 177.040 36.160 177.360 ;
        RECT 36.240 177.040 36.560 177.360 ;
        RECT 36.640 177.040 36.960 177.360 ;
        RECT 37.040 177.040 37.360 177.360 ;
        RECT 37.440 177.040 37.760 177.360 ;
        RECT 37.840 177.040 38.160 177.360 ;
        RECT 38.240 177.040 38.560 177.360 ;
        RECT 38.640 177.040 38.960 177.360 ;
        RECT 39.040 177.040 39.360 177.360 ;
        RECT 39.440 177.040 39.760 177.360 ;
        RECT 39.840 177.040 40.160 177.360 ;
        RECT 40.240 177.040 40.560 177.360 ;
        RECT 40.640 177.040 40.960 177.360 ;
        RECT 41.040 177.040 41.360 177.360 ;
        RECT 41.440 177.040 41.760 177.360 ;
        RECT 41.840 177.040 42.160 177.360 ;
        RECT 42.240 177.040 42.560 177.360 ;
        RECT 42.640 177.040 42.960 177.360 ;
        RECT 43.040 177.040 43.360 177.360 ;
        RECT 43.440 177.040 43.760 177.360 ;
        RECT 43.840 177.040 44.160 177.360 ;
        RECT 44.240 177.040 44.560 177.360 ;
        RECT 44.640 177.040 44.960 177.360 ;
        RECT 70.560 177.040 70.880 177.360 ;
        RECT 70.960 177.040 71.280 177.360 ;
        RECT 71.360 177.040 71.680 177.360 ;
        RECT 71.760 177.040 72.080 177.360 ;
        RECT 120.560 177.040 120.880 177.360 ;
        RECT 120.960 177.040 121.280 177.360 ;
        RECT 121.360 177.040 121.680 177.360 ;
        RECT 121.760 177.040 122.080 177.360 ;
        RECT 160.720 177.040 161.040 177.360 ;
        RECT 161.120 177.040 161.440 177.360 ;
        RECT 161.520 177.040 161.840 177.360 ;
        RECT 161.920 177.040 162.240 177.360 ;
        RECT 162.320 177.040 162.640 177.360 ;
        RECT 162.720 177.040 163.040 177.360 ;
        RECT 163.120 177.040 163.440 177.360 ;
        RECT 163.520 177.040 163.840 177.360 ;
        RECT 163.920 177.040 164.240 177.360 ;
        RECT 164.320 177.040 164.640 177.360 ;
        RECT 164.720 177.040 165.040 177.360 ;
        RECT 165.120 177.040 165.440 177.360 ;
        RECT 165.520 177.040 165.840 177.360 ;
        RECT 165.920 177.040 166.240 177.360 ;
        RECT 166.320 177.040 166.640 177.360 ;
        RECT 166.720 177.040 167.040 177.360 ;
        RECT 167.120 177.040 167.440 177.360 ;
        RECT 167.520 177.040 167.840 177.360 ;
        RECT 167.920 177.040 168.240 177.360 ;
        RECT 168.320 177.040 168.640 177.360 ;
        RECT 168.720 177.040 169.040 177.360 ;
        RECT 169.120 177.040 169.440 177.360 ;
        RECT 169.520 177.040 169.840 177.360 ;
        RECT 169.920 177.040 170.240 177.360 ;
        RECT 170.320 177.040 170.640 177.360 ;
        RECT 170.720 177.040 171.040 177.360 ;
        RECT 171.120 177.040 171.440 177.360 ;
        RECT 171.520 177.040 171.840 177.360 ;
        RECT 171.920 177.040 172.240 177.360 ;
        RECT 172.320 177.040 172.640 177.360 ;
        RECT 172.720 177.040 173.040 177.360 ;
        RECT 173.120 177.040 173.440 177.360 ;
        RECT 173.520 177.040 173.840 177.360 ;
        RECT 173.920 177.040 174.240 177.360 ;
        RECT 174.320 177.040 174.640 177.360 ;
        RECT 174.720 177.040 175.040 177.360 ;
        RECT 175.120 177.040 175.440 177.360 ;
        RECT 175.520 177.040 175.840 177.360 ;
        RECT 175.920 177.040 176.240 177.360 ;
        RECT 176.320 177.040 176.640 177.360 ;
        RECT 176.720 177.040 177.040 177.360 ;
        RECT 177.120 177.040 177.440 177.360 ;
        RECT 177.520 177.040 177.840 177.360 ;
        RECT 177.920 177.040 178.240 177.360 ;
        RECT 178.320 177.040 178.640 177.360 ;
        RECT 178.720 177.040 179.040 177.360 ;
        RECT 179.120 177.040 179.440 177.360 ;
        RECT 179.520 177.040 179.840 177.360 ;
        RECT 179.920 177.040 180.240 177.360 ;
        RECT 180.320 177.040 180.640 177.360 ;
        RECT 25.040 176.640 25.360 176.960 ;
        RECT 25.440 176.640 25.760 176.960 ;
        RECT 25.840 176.640 26.160 176.960 ;
        RECT 26.240 176.640 26.560 176.960 ;
        RECT 26.640 176.640 26.960 176.960 ;
        RECT 27.040 176.640 27.360 176.960 ;
        RECT 27.440 176.640 27.760 176.960 ;
        RECT 27.840 176.640 28.160 176.960 ;
        RECT 28.240 176.640 28.560 176.960 ;
        RECT 28.640 176.640 28.960 176.960 ;
        RECT 29.040 176.640 29.360 176.960 ;
        RECT 29.440 176.640 29.760 176.960 ;
        RECT 29.840 176.640 30.160 176.960 ;
        RECT 30.240 176.640 30.560 176.960 ;
        RECT 30.640 176.640 30.960 176.960 ;
        RECT 31.040 176.640 31.360 176.960 ;
        RECT 31.440 176.640 31.760 176.960 ;
        RECT 31.840 176.640 32.160 176.960 ;
        RECT 32.240 176.640 32.560 176.960 ;
        RECT 32.640 176.640 32.960 176.960 ;
        RECT 33.040 176.640 33.360 176.960 ;
        RECT 33.440 176.640 33.760 176.960 ;
        RECT 33.840 176.640 34.160 176.960 ;
        RECT 34.240 176.640 34.560 176.960 ;
        RECT 34.640 176.640 34.960 176.960 ;
        RECT 35.040 176.640 35.360 176.960 ;
        RECT 35.440 176.640 35.760 176.960 ;
        RECT 35.840 176.640 36.160 176.960 ;
        RECT 36.240 176.640 36.560 176.960 ;
        RECT 36.640 176.640 36.960 176.960 ;
        RECT 37.040 176.640 37.360 176.960 ;
        RECT 37.440 176.640 37.760 176.960 ;
        RECT 37.840 176.640 38.160 176.960 ;
        RECT 38.240 176.640 38.560 176.960 ;
        RECT 38.640 176.640 38.960 176.960 ;
        RECT 39.040 176.640 39.360 176.960 ;
        RECT 39.440 176.640 39.760 176.960 ;
        RECT 39.840 176.640 40.160 176.960 ;
        RECT 40.240 176.640 40.560 176.960 ;
        RECT 40.640 176.640 40.960 176.960 ;
        RECT 41.040 176.640 41.360 176.960 ;
        RECT 41.440 176.640 41.760 176.960 ;
        RECT 41.840 176.640 42.160 176.960 ;
        RECT 42.240 176.640 42.560 176.960 ;
        RECT 42.640 176.640 42.960 176.960 ;
        RECT 43.040 176.640 43.360 176.960 ;
        RECT 43.440 176.640 43.760 176.960 ;
        RECT 43.840 176.640 44.160 176.960 ;
        RECT 44.240 176.640 44.560 176.960 ;
        RECT 44.640 176.640 44.960 176.960 ;
        RECT 70.560 176.640 70.880 176.960 ;
        RECT 70.960 176.640 71.280 176.960 ;
        RECT 71.360 176.640 71.680 176.960 ;
        RECT 71.760 176.640 72.080 176.960 ;
        RECT 120.560 176.640 120.880 176.960 ;
        RECT 120.960 176.640 121.280 176.960 ;
        RECT 121.360 176.640 121.680 176.960 ;
        RECT 121.760 176.640 122.080 176.960 ;
        RECT 160.720 176.640 161.040 176.960 ;
        RECT 161.120 176.640 161.440 176.960 ;
        RECT 161.520 176.640 161.840 176.960 ;
        RECT 161.920 176.640 162.240 176.960 ;
        RECT 162.320 176.640 162.640 176.960 ;
        RECT 162.720 176.640 163.040 176.960 ;
        RECT 163.120 176.640 163.440 176.960 ;
        RECT 163.520 176.640 163.840 176.960 ;
        RECT 163.920 176.640 164.240 176.960 ;
        RECT 164.320 176.640 164.640 176.960 ;
        RECT 164.720 176.640 165.040 176.960 ;
        RECT 165.120 176.640 165.440 176.960 ;
        RECT 165.520 176.640 165.840 176.960 ;
        RECT 165.920 176.640 166.240 176.960 ;
        RECT 166.320 176.640 166.640 176.960 ;
        RECT 166.720 176.640 167.040 176.960 ;
        RECT 167.120 176.640 167.440 176.960 ;
        RECT 167.520 176.640 167.840 176.960 ;
        RECT 167.920 176.640 168.240 176.960 ;
        RECT 168.320 176.640 168.640 176.960 ;
        RECT 168.720 176.640 169.040 176.960 ;
        RECT 169.120 176.640 169.440 176.960 ;
        RECT 169.520 176.640 169.840 176.960 ;
        RECT 169.920 176.640 170.240 176.960 ;
        RECT 170.320 176.640 170.640 176.960 ;
        RECT 170.720 176.640 171.040 176.960 ;
        RECT 171.120 176.640 171.440 176.960 ;
        RECT 171.520 176.640 171.840 176.960 ;
        RECT 171.920 176.640 172.240 176.960 ;
        RECT 172.320 176.640 172.640 176.960 ;
        RECT 172.720 176.640 173.040 176.960 ;
        RECT 173.120 176.640 173.440 176.960 ;
        RECT 173.520 176.640 173.840 176.960 ;
        RECT 173.920 176.640 174.240 176.960 ;
        RECT 174.320 176.640 174.640 176.960 ;
        RECT 174.720 176.640 175.040 176.960 ;
        RECT 175.120 176.640 175.440 176.960 ;
        RECT 175.520 176.640 175.840 176.960 ;
        RECT 175.920 176.640 176.240 176.960 ;
        RECT 176.320 176.640 176.640 176.960 ;
        RECT 176.720 176.640 177.040 176.960 ;
        RECT 177.120 176.640 177.440 176.960 ;
        RECT 177.520 176.640 177.840 176.960 ;
        RECT 177.920 176.640 178.240 176.960 ;
        RECT 178.320 176.640 178.640 176.960 ;
        RECT 178.720 176.640 179.040 176.960 ;
        RECT 179.120 176.640 179.440 176.960 ;
        RECT 179.520 176.640 179.840 176.960 ;
        RECT 179.920 176.640 180.240 176.960 ;
        RECT 180.320 176.640 180.640 176.960 ;
        RECT 25.040 176.240 25.360 176.560 ;
        RECT 25.440 176.240 25.760 176.560 ;
        RECT 25.840 176.240 26.160 176.560 ;
        RECT 26.240 176.240 26.560 176.560 ;
        RECT 26.640 176.240 26.960 176.560 ;
        RECT 27.040 176.240 27.360 176.560 ;
        RECT 27.440 176.240 27.760 176.560 ;
        RECT 27.840 176.240 28.160 176.560 ;
        RECT 28.240 176.240 28.560 176.560 ;
        RECT 28.640 176.240 28.960 176.560 ;
        RECT 29.040 176.240 29.360 176.560 ;
        RECT 29.440 176.240 29.760 176.560 ;
        RECT 29.840 176.240 30.160 176.560 ;
        RECT 30.240 176.240 30.560 176.560 ;
        RECT 30.640 176.240 30.960 176.560 ;
        RECT 31.040 176.240 31.360 176.560 ;
        RECT 31.440 176.240 31.760 176.560 ;
        RECT 31.840 176.240 32.160 176.560 ;
        RECT 32.240 176.240 32.560 176.560 ;
        RECT 32.640 176.240 32.960 176.560 ;
        RECT 33.040 176.240 33.360 176.560 ;
        RECT 33.440 176.240 33.760 176.560 ;
        RECT 33.840 176.240 34.160 176.560 ;
        RECT 34.240 176.240 34.560 176.560 ;
        RECT 34.640 176.240 34.960 176.560 ;
        RECT 35.040 176.240 35.360 176.560 ;
        RECT 35.440 176.240 35.760 176.560 ;
        RECT 35.840 176.240 36.160 176.560 ;
        RECT 36.240 176.240 36.560 176.560 ;
        RECT 36.640 176.240 36.960 176.560 ;
        RECT 37.040 176.240 37.360 176.560 ;
        RECT 37.440 176.240 37.760 176.560 ;
        RECT 37.840 176.240 38.160 176.560 ;
        RECT 38.240 176.240 38.560 176.560 ;
        RECT 38.640 176.240 38.960 176.560 ;
        RECT 39.040 176.240 39.360 176.560 ;
        RECT 39.440 176.240 39.760 176.560 ;
        RECT 39.840 176.240 40.160 176.560 ;
        RECT 40.240 176.240 40.560 176.560 ;
        RECT 40.640 176.240 40.960 176.560 ;
        RECT 41.040 176.240 41.360 176.560 ;
        RECT 41.440 176.240 41.760 176.560 ;
        RECT 41.840 176.240 42.160 176.560 ;
        RECT 42.240 176.240 42.560 176.560 ;
        RECT 42.640 176.240 42.960 176.560 ;
        RECT 43.040 176.240 43.360 176.560 ;
        RECT 43.440 176.240 43.760 176.560 ;
        RECT 43.840 176.240 44.160 176.560 ;
        RECT 44.240 176.240 44.560 176.560 ;
        RECT 44.640 176.240 44.960 176.560 ;
        RECT 70.560 176.240 70.880 176.560 ;
        RECT 70.960 176.240 71.280 176.560 ;
        RECT 71.360 176.240 71.680 176.560 ;
        RECT 71.760 176.240 72.080 176.560 ;
        RECT 120.560 176.240 120.880 176.560 ;
        RECT 120.960 176.240 121.280 176.560 ;
        RECT 121.360 176.240 121.680 176.560 ;
        RECT 121.760 176.240 122.080 176.560 ;
        RECT 160.720 176.240 161.040 176.560 ;
        RECT 161.120 176.240 161.440 176.560 ;
        RECT 161.520 176.240 161.840 176.560 ;
        RECT 161.920 176.240 162.240 176.560 ;
        RECT 162.320 176.240 162.640 176.560 ;
        RECT 162.720 176.240 163.040 176.560 ;
        RECT 163.120 176.240 163.440 176.560 ;
        RECT 163.520 176.240 163.840 176.560 ;
        RECT 163.920 176.240 164.240 176.560 ;
        RECT 164.320 176.240 164.640 176.560 ;
        RECT 164.720 176.240 165.040 176.560 ;
        RECT 165.120 176.240 165.440 176.560 ;
        RECT 165.520 176.240 165.840 176.560 ;
        RECT 165.920 176.240 166.240 176.560 ;
        RECT 166.320 176.240 166.640 176.560 ;
        RECT 166.720 176.240 167.040 176.560 ;
        RECT 167.120 176.240 167.440 176.560 ;
        RECT 167.520 176.240 167.840 176.560 ;
        RECT 167.920 176.240 168.240 176.560 ;
        RECT 168.320 176.240 168.640 176.560 ;
        RECT 168.720 176.240 169.040 176.560 ;
        RECT 169.120 176.240 169.440 176.560 ;
        RECT 169.520 176.240 169.840 176.560 ;
        RECT 169.920 176.240 170.240 176.560 ;
        RECT 170.320 176.240 170.640 176.560 ;
        RECT 170.720 176.240 171.040 176.560 ;
        RECT 171.120 176.240 171.440 176.560 ;
        RECT 171.520 176.240 171.840 176.560 ;
        RECT 171.920 176.240 172.240 176.560 ;
        RECT 172.320 176.240 172.640 176.560 ;
        RECT 172.720 176.240 173.040 176.560 ;
        RECT 173.120 176.240 173.440 176.560 ;
        RECT 173.520 176.240 173.840 176.560 ;
        RECT 173.920 176.240 174.240 176.560 ;
        RECT 174.320 176.240 174.640 176.560 ;
        RECT 174.720 176.240 175.040 176.560 ;
        RECT 175.120 176.240 175.440 176.560 ;
        RECT 175.520 176.240 175.840 176.560 ;
        RECT 175.920 176.240 176.240 176.560 ;
        RECT 176.320 176.240 176.640 176.560 ;
        RECT 176.720 176.240 177.040 176.560 ;
        RECT 177.120 176.240 177.440 176.560 ;
        RECT 177.520 176.240 177.840 176.560 ;
        RECT 177.920 176.240 178.240 176.560 ;
        RECT 178.320 176.240 178.640 176.560 ;
        RECT 178.720 176.240 179.040 176.560 ;
        RECT 179.120 176.240 179.440 176.560 ;
        RECT 179.520 176.240 179.840 176.560 ;
        RECT 179.920 176.240 180.240 176.560 ;
        RECT 180.320 176.240 180.640 176.560 ;
        RECT 25.040 175.840 25.360 176.160 ;
        RECT 25.440 175.840 25.760 176.160 ;
        RECT 25.840 175.840 26.160 176.160 ;
        RECT 26.240 175.840 26.560 176.160 ;
        RECT 26.640 175.840 26.960 176.160 ;
        RECT 27.040 175.840 27.360 176.160 ;
        RECT 27.440 175.840 27.760 176.160 ;
        RECT 27.840 175.840 28.160 176.160 ;
        RECT 28.240 175.840 28.560 176.160 ;
        RECT 28.640 175.840 28.960 176.160 ;
        RECT 29.040 175.840 29.360 176.160 ;
        RECT 29.440 175.840 29.760 176.160 ;
        RECT 29.840 175.840 30.160 176.160 ;
        RECT 30.240 175.840 30.560 176.160 ;
        RECT 30.640 175.840 30.960 176.160 ;
        RECT 31.040 175.840 31.360 176.160 ;
        RECT 31.440 175.840 31.760 176.160 ;
        RECT 31.840 175.840 32.160 176.160 ;
        RECT 32.240 175.840 32.560 176.160 ;
        RECT 32.640 175.840 32.960 176.160 ;
        RECT 33.040 175.840 33.360 176.160 ;
        RECT 33.440 175.840 33.760 176.160 ;
        RECT 33.840 175.840 34.160 176.160 ;
        RECT 34.240 175.840 34.560 176.160 ;
        RECT 34.640 175.840 34.960 176.160 ;
        RECT 35.040 175.840 35.360 176.160 ;
        RECT 35.440 175.840 35.760 176.160 ;
        RECT 35.840 175.840 36.160 176.160 ;
        RECT 36.240 175.840 36.560 176.160 ;
        RECT 36.640 175.840 36.960 176.160 ;
        RECT 37.040 175.840 37.360 176.160 ;
        RECT 37.440 175.840 37.760 176.160 ;
        RECT 37.840 175.840 38.160 176.160 ;
        RECT 38.240 175.840 38.560 176.160 ;
        RECT 38.640 175.840 38.960 176.160 ;
        RECT 39.040 175.840 39.360 176.160 ;
        RECT 39.440 175.840 39.760 176.160 ;
        RECT 39.840 175.840 40.160 176.160 ;
        RECT 40.240 175.840 40.560 176.160 ;
        RECT 40.640 175.840 40.960 176.160 ;
        RECT 41.040 175.840 41.360 176.160 ;
        RECT 41.440 175.840 41.760 176.160 ;
        RECT 41.840 175.840 42.160 176.160 ;
        RECT 42.240 175.840 42.560 176.160 ;
        RECT 42.640 175.840 42.960 176.160 ;
        RECT 43.040 175.840 43.360 176.160 ;
        RECT 43.440 175.840 43.760 176.160 ;
        RECT 43.840 175.840 44.160 176.160 ;
        RECT 44.240 175.840 44.560 176.160 ;
        RECT 44.640 175.840 44.960 176.160 ;
        RECT 70.560 175.840 70.880 176.160 ;
        RECT 70.960 175.840 71.280 176.160 ;
        RECT 71.360 175.840 71.680 176.160 ;
        RECT 71.760 175.840 72.080 176.160 ;
        RECT 120.560 175.840 120.880 176.160 ;
        RECT 120.960 175.840 121.280 176.160 ;
        RECT 121.360 175.840 121.680 176.160 ;
        RECT 121.760 175.840 122.080 176.160 ;
        RECT 160.720 175.840 161.040 176.160 ;
        RECT 161.120 175.840 161.440 176.160 ;
        RECT 161.520 175.840 161.840 176.160 ;
        RECT 161.920 175.840 162.240 176.160 ;
        RECT 162.320 175.840 162.640 176.160 ;
        RECT 162.720 175.840 163.040 176.160 ;
        RECT 163.120 175.840 163.440 176.160 ;
        RECT 163.520 175.840 163.840 176.160 ;
        RECT 163.920 175.840 164.240 176.160 ;
        RECT 164.320 175.840 164.640 176.160 ;
        RECT 164.720 175.840 165.040 176.160 ;
        RECT 165.120 175.840 165.440 176.160 ;
        RECT 165.520 175.840 165.840 176.160 ;
        RECT 165.920 175.840 166.240 176.160 ;
        RECT 166.320 175.840 166.640 176.160 ;
        RECT 166.720 175.840 167.040 176.160 ;
        RECT 167.120 175.840 167.440 176.160 ;
        RECT 167.520 175.840 167.840 176.160 ;
        RECT 167.920 175.840 168.240 176.160 ;
        RECT 168.320 175.840 168.640 176.160 ;
        RECT 168.720 175.840 169.040 176.160 ;
        RECT 169.120 175.840 169.440 176.160 ;
        RECT 169.520 175.840 169.840 176.160 ;
        RECT 169.920 175.840 170.240 176.160 ;
        RECT 170.320 175.840 170.640 176.160 ;
        RECT 170.720 175.840 171.040 176.160 ;
        RECT 171.120 175.840 171.440 176.160 ;
        RECT 171.520 175.840 171.840 176.160 ;
        RECT 171.920 175.840 172.240 176.160 ;
        RECT 172.320 175.840 172.640 176.160 ;
        RECT 172.720 175.840 173.040 176.160 ;
        RECT 173.120 175.840 173.440 176.160 ;
        RECT 173.520 175.840 173.840 176.160 ;
        RECT 173.920 175.840 174.240 176.160 ;
        RECT 174.320 175.840 174.640 176.160 ;
        RECT 174.720 175.840 175.040 176.160 ;
        RECT 175.120 175.840 175.440 176.160 ;
        RECT 175.520 175.840 175.840 176.160 ;
        RECT 175.920 175.840 176.240 176.160 ;
        RECT 176.320 175.840 176.640 176.160 ;
        RECT 176.720 175.840 177.040 176.160 ;
        RECT 177.120 175.840 177.440 176.160 ;
        RECT 177.520 175.840 177.840 176.160 ;
        RECT 177.920 175.840 178.240 176.160 ;
        RECT 178.320 175.840 178.640 176.160 ;
        RECT 178.720 175.840 179.040 176.160 ;
        RECT 179.120 175.840 179.440 176.160 ;
        RECT 179.520 175.840 179.840 176.160 ;
        RECT 179.920 175.840 180.240 176.160 ;
        RECT 180.320 175.840 180.640 176.160 ;
        RECT 25.040 175.440 25.360 175.760 ;
        RECT 25.440 175.440 25.760 175.760 ;
        RECT 25.840 175.440 26.160 175.760 ;
        RECT 26.240 175.440 26.560 175.760 ;
        RECT 26.640 175.440 26.960 175.760 ;
        RECT 27.040 175.440 27.360 175.760 ;
        RECT 27.440 175.440 27.760 175.760 ;
        RECT 27.840 175.440 28.160 175.760 ;
        RECT 28.240 175.440 28.560 175.760 ;
        RECT 28.640 175.440 28.960 175.760 ;
        RECT 29.040 175.440 29.360 175.760 ;
        RECT 29.440 175.440 29.760 175.760 ;
        RECT 29.840 175.440 30.160 175.760 ;
        RECT 30.240 175.440 30.560 175.760 ;
        RECT 30.640 175.440 30.960 175.760 ;
        RECT 31.040 175.440 31.360 175.760 ;
        RECT 31.440 175.440 31.760 175.760 ;
        RECT 31.840 175.440 32.160 175.760 ;
        RECT 32.240 175.440 32.560 175.760 ;
        RECT 32.640 175.440 32.960 175.760 ;
        RECT 33.040 175.440 33.360 175.760 ;
        RECT 33.440 175.440 33.760 175.760 ;
        RECT 33.840 175.440 34.160 175.760 ;
        RECT 34.240 175.440 34.560 175.760 ;
        RECT 34.640 175.440 34.960 175.760 ;
        RECT 35.040 175.440 35.360 175.760 ;
        RECT 35.440 175.440 35.760 175.760 ;
        RECT 35.840 175.440 36.160 175.760 ;
        RECT 36.240 175.440 36.560 175.760 ;
        RECT 36.640 175.440 36.960 175.760 ;
        RECT 37.040 175.440 37.360 175.760 ;
        RECT 37.440 175.440 37.760 175.760 ;
        RECT 37.840 175.440 38.160 175.760 ;
        RECT 38.240 175.440 38.560 175.760 ;
        RECT 38.640 175.440 38.960 175.760 ;
        RECT 39.040 175.440 39.360 175.760 ;
        RECT 39.440 175.440 39.760 175.760 ;
        RECT 39.840 175.440 40.160 175.760 ;
        RECT 40.240 175.440 40.560 175.760 ;
        RECT 40.640 175.440 40.960 175.760 ;
        RECT 41.040 175.440 41.360 175.760 ;
        RECT 41.440 175.440 41.760 175.760 ;
        RECT 41.840 175.440 42.160 175.760 ;
        RECT 42.240 175.440 42.560 175.760 ;
        RECT 42.640 175.440 42.960 175.760 ;
        RECT 43.040 175.440 43.360 175.760 ;
        RECT 43.440 175.440 43.760 175.760 ;
        RECT 43.840 175.440 44.160 175.760 ;
        RECT 44.240 175.440 44.560 175.760 ;
        RECT 44.640 175.440 44.960 175.760 ;
        RECT 70.560 175.440 70.880 175.760 ;
        RECT 70.960 175.440 71.280 175.760 ;
        RECT 71.360 175.440 71.680 175.760 ;
        RECT 71.760 175.440 72.080 175.760 ;
        RECT 120.560 175.440 120.880 175.760 ;
        RECT 120.960 175.440 121.280 175.760 ;
        RECT 121.360 175.440 121.680 175.760 ;
        RECT 121.760 175.440 122.080 175.760 ;
        RECT 160.720 175.440 161.040 175.760 ;
        RECT 161.120 175.440 161.440 175.760 ;
        RECT 161.520 175.440 161.840 175.760 ;
        RECT 161.920 175.440 162.240 175.760 ;
        RECT 162.320 175.440 162.640 175.760 ;
        RECT 162.720 175.440 163.040 175.760 ;
        RECT 163.120 175.440 163.440 175.760 ;
        RECT 163.520 175.440 163.840 175.760 ;
        RECT 163.920 175.440 164.240 175.760 ;
        RECT 164.320 175.440 164.640 175.760 ;
        RECT 164.720 175.440 165.040 175.760 ;
        RECT 165.120 175.440 165.440 175.760 ;
        RECT 165.520 175.440 165.840 175.760 ;
        RECT 165.920 175.440 166.240 175.760 ;
        RECT 166.320 175.440 166.640 175.760 ;
        RECT 166.720 175.440 167.040 175.760 ;
        RECT 167.120 175.440 167.440 175.760 ;
        RECT 167.520 175.440 167.840 175.760 ;
        RECT 167.920 175.440 168.240 175.760 ;
        RECT 168.320 175.440 168.640 175.760 ;
        RECT 168.720 175.440 169.040 175.760 ;
        RECT 169.120 175.440 169.440 175.760 ;
        RECT 169.520 175.440 169.840 175.760 ;
        RECT 169.920 175.440 170.240 175.760 ;
        RECT 170.320 175.440 170.640 175.760 ;
        RECT 170.720 175.440 171.040 175.760 ;
        RECT 171.120 175.440 171.440 175.760 ;
        RECT 171.520 175.440 171.840 175.760 ;
        RECT 171.920 175.440 172.240 175.760 ;
        RECT 172.320 175.440 172.640 175.760 ;
        RECT 172.720 175.440 173.040 175.760 ;
        RECT 173.120 175.440 173.440 175.760 ;
        RECT 173.520 175.440 173.840 175.760 ;
        RECT 173.920 175.440 174.240 175.760 ;
        RECT 174.320 175.440 174.640 175.760 ;
        RECT 174.720 175.440 175.040 175.760 ;
        RECT 175.120 175.440 175.440 175.760 ;
        RECT 175.520 175.440 175.840 175.760 ;
        RECT 175.920 175.440 176.240 175.760 ;
        RECT 176.320 175.440 176.640 175.760 ;
        RECT 176.720 175.440 177.040 175.760 ;
        RECT 177.120 175.440 177.440 175.760 ;
        RECT 177.520 175.440 177.840 175.760 ;
        RECT 177.920 175.440 178.240 175.760 ;
        RECT 178.320 175.440 178.640 175.760 ;
        RECT 178.720 175.440 179.040 175.760 ;
        RECT 179.120 175.440 179.440 175.760 ;
        RECT 179.520 175.440 179.840 175.760 ;
        RECT 179.920 175.440 180.240 175.760 ;
        RECT 180.320 175.440 180.640 175.760 ;
        RECT 25.040 175.040 25.360 175.360 ;
        RECT 25.440 175.040 25.760 175.360 ;
        RECT 25.840 175.040 26.160 175.360 ;
        RECT 26.240 175.040 26.560 175.360 ;
        RECT 26.640 175.040 26.960 175.360 ;
        RECT 27.040 175.040 27.360 175.360 ;
        RECT 27.440 175.040 27.760 175.360 ;
        RECT 27.840 175.040 28.160 175.360 ;
        RECT 28.240 175.040 28.560 175.360 ;
        RECT 28.640 175.040 28.960 175.360 ;
        RECT 29.040 175.040 29.360 175.360 ;
        RECT 29.440 175.040 29.760 175.360 ;
        RECT 29.840 175.040 30.160 175.360 ;
        RECT 30.240 175.040 30.560 175.360 ;
        RECT 30.640 175.040 30.960 175.360 ;
        RECT 31.040 175.040 31.360 175.360 ;
        RECT 31.440 175.040 31.760 175.360 ;
        RECT 31.840 175.040 32.160 175.360 ;
        RECT 32.240 175.040 32.560 175.360 ;
        RECT 32.640 175.040 32.960 175.360 ;
        RECT 33.040 175.040 33.360 175.360 ;
        RECT 33.440 175.040 33.760 175.360 ;
        RECT 33.840 175.040 34.160 175.360 ;
        RECT 34.240 175.040 34.560 175.360 ;
        RECT 34.640 175.040 34.960 175.360 ;
        RECT 35.040 175.040 35.360 175.360 ;
        RECT 35.440 175.040 35.760 175.360 ;
        RECT 35.840 175.040 36.160 175.360 ;
        RECT 36.240 175.040 36.560 175.360 ;
        RECT 36.640 175.040 36.960 175.360 ;
        RECT 37.040 175.040 37.360 175.360 ;
        RECT 37.440 175.040 37.760 175.360 ;
        RECT 37.840 175.040 38.160 175.360 ;
        RECT 38.240 175.040 38.560 175.360 ;
        RECT 38.640 175.040 38.960 175.360 ;
        RECT 39.040 175.040 39.360 175.360 ;
        RECT 39.440 175.040 39.760 175.360 ;
        RECT 39.840 175.040 40.160 175.360 ;
        RECT 40.240 175.040 40.560 175.360 ;
        RECT 40.640 175.040 40.960 175.360 ;
        RECT 41.040 175.040 41.360 175.360 ;
        RECT 41.440 175.040 41.760 175.360 ;
        RECT 41.840 175.040 42.160 175.360 ;
        RECT 42.240 175.040 42.560 175.360 ;
        RECT 42.640 175.040 42.960 175.360 ;
        RECT 43.040 175.040 43.360 175.360 ;
        RECT 43.440 175.040 43.760 175.360 ;
        RECT 43.840 175.040 44.160 175.360 ;
        RECT 44.240 175.040 44.560 175.360 ;
        RECT 44.640 175.040 44.960 175.360 ;
        RECT 70.560 175.040 70.880 175.360 ;
        RECT 70.960 175.040 71.280 175.360 ;
        RECT 71.360 175.040 71.680 175.360 ;
        RECT 71.760 175.040 72.080 175.360 ;
        RECT 120.560 175.040 120.880 175.360 ;
        RECT 120.960 175.040 121.280 175.360 ;
        RECT 121.360 175.040 121.680 175.360 ;
        RECT 121.760 175.040 122.080 175.360 ;
        RECT 160.720 175.040 161.040 175.360 ;
        RECT 161.120 175.040 161.440 175.360 ;
        RECT 161.520 175.040 161.840 175.360 ;
        RECT 161.920 175.040 162.240 175.360 ;
        RECT 162.320 175.040 162.640 175.360 ;
        RECT 162.720 175.040 163.040 175.360 ;
        RECT 163.120 175.040 163.440 175.360 ;
        RECT 163.520 175.040 163.840 175.360 ;
        RECT 163.920 175.040 164.240 175.360 ;
        RECT 164.320 175.040 164.640 175.360 ;
        RECT 164.720 175.040 165.040 175.360 ;
        RECT 165.120 175.040 165.440 175.360 ;
        RECT 165.520 175.040 165.840 175.360 ;
        RECT 165.920 175.040 166.240 175.360 ;
        RECT 166.320 175.040 166.640 175.360 ;
        RECT 166.720 175.040 167.040 175.360 ;
        RECT 167.120 175.040 167.440 175.360 ;
        RECT 167.520 175.040 167.840 175.360 ;
        RECT 167.920 175.040 168.240 175.360 ;
        RECT 168.320 175.040 168.640 175.360 ;
        RECT 168.720 175.040 169.040 175.360 ;
        RECT 169.120 175.040 169.440 175.360 ;
        RECT 169.520 175.040 169.840 175.360 ;
        RECT 169.920 175.040 170.240 175.360 ;
        RECT 170.320 175.040 170.640 175.360 ;
        RECT 170.720 175.040 171.040 175.360 ;
        RECT 171.120 175.040 171.440 175.360 ;
        RECT 171.520 175.040 171.840 175.360 ;
        RECT 171.920 175.040 172.240 175.360 ;
        RECT 172.320 175.040 172.640 175.360 ;
        RECT 172.720 175.040 173.040 175.360 ;
        RECT 173.120 175.040 173.440 175.360 ;
        RECT 173.520 175.040 173.840 175.360 ;
        RECT 173.920 175.040 174.240 175.360 ;
        RECT 174.320 175.040 174.640 175.360 ;
        RECT 174.720 175.040 175.040 175.360 ;
        RECT 175.120 175.040 175.440 175.360 ;
        RECT 175.520 175.040 175.840 175.360 ;
        RECT 175.920 175.040 176.240 175.360 ;
        RECT 176.320 175.040 176.640 175.360 ;
        RECT 176.720 175.040 177.040 175.360 ;
        RECT 177.120 175.040 177.440 175.360 ;
        RECT 177.520 175.040 177.840 175.360 ;
        RECT 177.920 175.040 178.240 175.360 ;
        RECT 178.320 175.040 178.640 175.360 ;
        RECT 178.720 175.040 179.040 175.360 ;
        RECT 179.120 175.040 179.440 175.360 ;
        RECT 179.520 175.040 179.840 175.360 ;
        RECT 179.920 175.040 180.240 175.360 ;
        RECT 180.320 175.040 180.640 175.360 ;
        RECT 25.040 174.640 25.360 174.960 ;
        RECT 25.440 174.640 25.760 174.960 ;
        RECT 25.840 174.640 26.160 174.960 ;
        RECT 26.240 174.640 26.560 174.960 ;
        RECT 26.640 174.640 26.960 174.960 ;
        RECT 27.040 174.640 27.360 174.960 ;
        RECT 27.440 174.640 27.760 174.960 ;
        RECT 27.840 174.640 28.160 174.960 ;
        RECT 28.240 174.640 28.560 174.960 ;
        RECT 28.640 174.640 28.960 174.960 ;
        RECT 29.040 174.640 29.360 174.960 ;
        RECT 29.440 174.640 29.760 174.960 ;
        RECT 29.840 174.640 30.160 174.960 ;
        RECT 30.240 174.640 30.560 174.960 ;
        RECT 30.640 174.640 30.960 174.960 ;
        RECT 31.040 174.640 31.360 174.960 ;
        RECT 31.440 174.640 31.760 174.960 ;
        RECT 31.840 174.640 32.160 174.960 ;
        RECT 32.240 174.640 32.560 174.960 ;
        RECT 32.640 174.640 32.960 174.960 ;
        RECT 33.040 174.640 33.360 174.960 ;
        RECT 33.440 174.640 33.760 174.960 ;
        RECT 33.840 174.640 34.160 174.960 ;
        RECT 34.240 174.640 34.560 174.960 ;
        RECT 34.640 174.640 34.960 174.960 ;
        RECT 35.040 174.640 35.360 174.960 ;
        RECT 35.440 174.640 35.760 174.960 ;
        RECT 35.840 174.640 36.160 174.960 ;
        RECT 36.240 174.640 36.560 174.960 ;
        RECT 36.640 174.640 36.960 174.960 ;
        RECT 37.040 174.640 37.360 174.960 ;
        RECT 37.440 174.640 37.760 174.960 ;
        RECT 37.840 174.640 38.160 174.960 ;
        RECT 38.240 174.640 38.560 174.960 ;
        RECT 38.640 174.640 38.960 174.960 ;
        RECT 39.040 174.640 39.360 174.960 ;
        RECT 39.440 174.640 39.760 174.960 ;
        RECT 39.840 174.640 40.160 174.960 ;
        RECT 40.240 174.640 40.560 174.960 ;
        RECT 40.640 174.640 40.960 174.960 ;
        RECT 41.040 174.640 41.360 174.960 ;
        RECT 41.440 174.640 41.760 174.960 ;
        RECT 41.840 174.640 42.160 174.960 ;
        RECT 42.240 174.640 42.560 174.960 ;
        RECT 42.640 174.640 42.960 174.960 ;
        RECT 43.040 174.640 43.360 174.960 ;
        RECT 43.440 174.640 43.760 174.960 ;
        RECT 43.840 174.640 44.160 174.960 ;
        RECT 44.240 174.640 44.560 174.960 ;
        RECT 44.640 174.640 44.960 174.960 ;
        RECT 70.560 174.640 70.880 174.960 ;
        RECT 70.960 174.640 71.280 174.960 ;
        RECT 71.360 174.640 71.680 174.960 ;
        RECT 71.760 174.640 72.080 174.960 ;
        RECT 120.560 174.640 120.880 174.960 ;
        RECT 120.960 174.640 121.280 174.960 ;
        RECT 121.360 174.640 121.680 174.960 ;
        RECT 121.760 174.640 122.080 174.960 ;
        RECT 160.720 174.640 161.040 174.960 ;
        RECT 161.120 174.640 161.440 174.960 ;
        RECT 161.520 174.640 161.840 174.960 ;
        RECT 161.920 174.640 162.240 174.960 ;
        RECT 162.320 174.640 162.640 174.960 ;
        RECT 162.720 174.640 163.040 174.960 ;
        RECT 163.120 174.640 163.440 174.960 ;
        RECT 163.520 174.640 163.840 174.960 ;
        RECT 163.920 174.640 164.240 174.960 ;
        RECT 164.320 174.640 164.640 174.960 ;
        RECT 164.720 174.640 165.040 174.960 ;
        RECT 165.120 174.640 165.440 174.960 ;
        RECT 165.520 174.640 165.840 174.960 ;
        RECT 165.920 174.640 166.240 174.960 ;
        RECT 166.320 174.640 166.640 174.960 ;
        RECT 166.720 174.640 167.040 174.960 ;
        RECT 167.120 174.640 167.440 174.960 ;
        RECT 167.520 174.640 167.840 174.960 ;
        RECT 167.920 174.640 168.240 174.960 ;
        RECT 168.320 174.640 168.640 174.960 ;
        RECT 168.720 174.640 169.040 174.960 ;
        RECT 169.120 174.640 169.440 174.960 ;
        RECT 169.520 174.640 169.840 174.960 ;
        RECT 169.920 174.640 170.240 174.960 ;
        RECT 170.320 174.640 170.640 174.960 ;
        RECT 170.720 174.640 171.040 174.960 ;
        RECT 171.120 174.640 171.440 174.960 ;
        RECT 171.520 174.640 171.840 174.960 ;
        RECT 171.920 174.640 172.240 174.960 ;
        RECT 172.320 174.640 172.640 174.960 ;
        RECT 172.720 174.640 173.040 174.960 ;
        RECT 173.120 174.640 173.440 174.960 ;
        RECT 173.520 174.640 173.840 174.960 ;
        RECT 173.920 174.640 174.240 174.960 ;
        RECT 174.320 174.640 174.640 174.960 ;
        RECT 174.720 174.640 175.040 174.960 ;
        RECT 175.120 174.640 175.440 174.960 ;
        RECT 175.520 174.640 175.840 174.960 ;
        RECT 175.920 174.640 176.240 174.960 ;
        RECT 176.320 174.640 176.640 174.960 ;
        RECT 176.720 174.640 177.040 174.960 ;
        RECT 177.120 174.640 177.440 174.960 ;
        RECT 177.520 174.640 177.840 174.960 ;
        RECT 177.920 174.640 178.240 174.960 ;
        RECT 178.320 174.640 178.640 174.960 ;
        RECT 178.720 174.640 179.040 174.960 ;
        RECT 179.120 174.640 179.440 174.960 ;
        RECT 179.520 174.640 179.840 174.960 ;
        RECT 179.920 174.640 180.240 174.960 ;
        RECT 180.320 174.640 180.640 174.960 ;
        RECT 25.040 174.240 25.360 174.560 ;
        RECT 25.440 174.240 25.760 174.560 ;
        RECT 25.840 174.240 26.160 174.560 ;
        RECT 26.240 174.240 26.560 174.560 ;
        RECT 26.640 174.240 26.960 174.560 ;
        RECT 27.040 174.240 27.360 174.560 ;
        RECT 27.440 174.240 27.760 174.560 ;
        RECT 27.840 174.240 28.160 174.560 ;
        RECT 28.240 174.240 28.560 174.560 ;
        RECT 28.640 174.240 28.960 174.560 ;
        RECT 29.040 174.240 29.360 174.560 ;
        RECT 29.440 174.240 29.760 174.560 ;
        RECT 29.840 174.240 30.160 174.560 ;
        RECT 30.240 174.240 30.560 174.560 ;
        RECT 30.640 174.240 30.960 174.560 ;
        RECT 31.040 174.240 31.360 174.560 ;
        RECT 31.440 174.240 31.760 174.560 ;
        RECT 31.840 174.240 32.160 174.560 ;
        RECT 32.240 174.240 32.560 174.560 ;
        RECT 32.640 174.240 32.960 174.560 ;
        RECT 33.040 174.240 33.360 174.560 ;
        RECT 33.440 174.240 33.760 174.560 ;
        RECT 33.840 174.240 34.160 174.560 ;
        RECT 34.240 174.240 34.560 174.560 ;
        RECT 34.640 174.240 34.960 174.560 ;
        RECT 35.040 174.240 35.360 174.560 ;
        RECT 35.440 174.240 35.760 174.560 ;
        RECT 35.840 174.240 36.160 174.560 ;
        RECT 36.240 174.240 36.560 174.560 ;
        RECT 36.640 174.240 36.960 174.560 ;
        RECT 37.040 174.240 37.360 174.560 ;
        RECT 37.440 174.240 37.760 174.560 ;
        RECT 37.840 174.240 38.160 174.560 ;
        RECT 38.240 174.240 38.560 174.560 ;
        RECT 38.640 174.240 38.960 174.560 ;
        RECT 39.040 174.240 39.360 174.560 ;
        RECT 39.440 174.240 39.760 174.560 ;
        RECT 39.840 174.240 40.160 174.560 ;
        RECT 40.240 174.240 40.560 174.560 ;
        RECT 40.640 174.240 40.960 174.560 ;
        RECT 41.040 174.240 41.360 174.560 ;
        RECT 41.440 174.240 41.760 174.560 ;
        RECT 41.840 174.240 42.160 174.560 ;
        RECT 42.240 174.240 42.560 174.560 ;
        RECT 42.640 174.240 42.960 174.560 ;
        RECT 43.040 174.240 43.360 174.560 ;
        RECT 43.440 174.240 43.760 174.560 ;
        RECT 43.840 174.240 44.160 174.560 ;
        RECT 44.240 174.240 44.560 174.560 ;
        RECT 44.640 174.240 44.960 174.560 ;
        RECT 70.560 174.240 70.880 174.560 ;
        RECT 70.960 174.240 71.280 174.560 ;
        RECT 71.360 174.240 71.680 174.560 ;
        RECT 71.760 174.240 72.080 174.560 ;
        RECT 120.560 174.240 120.880 174.560 ;
        RECT 120.960 174.240 121.280 174.560 ;
        RECT 121.360 174.240 121.680 174.560 ;
        RECT 121.760 174.240 122.080 174.560 ;
        RECT 160.720 174.240 161.040 174.560 ;
        RECT 161.120 174.240 161.440 174.560 ;
        RECT 161.520 174.240 161.840 174.560 ;
        RECT 161.920 174.240 162.240 174.560 ;
        RECT 162.320 174.240 162.640 174.560 ;
        RECT 162.720 174.240 163.040 174.560 ;
        RECT 163.120 174.240 163.440 174.560 ;
        RECT 163.520 174.240 163.840 174.560 ;
        RECT 163.920 174.240 164.240 174.560 ;
        RECT 164.320 174.240 164.640 174.560 ;
        RECT 164.720 174.240 165.040 174.560 ;
        RECT 165.120 174.240 165.440 174.560 ;
        RECT 165.520 174.240 165.840 174.560 ;
        RECT 165.920 174.240 166.240 174.560 ;
        RECT 166.320 174.240 166.640 174.560 ;
        RECT 166.720 174.240 167.040 174.560 ;
        RECT 167.120 174.240 167.440 174.560 ;
        RECT 167.520 174.240 167.840 174.560 ;
        RECT 167.920 174.240 168.240 174.560 ;
        RECT 168.320 174.240 168.640 174.560 ;
        RECT 168.720 174.240 169.040 174.560 ;
        RECT 169.120 174.240 169.440 174.560 ;
        RECT 169.520 174.240 169.840 174.560 ;
        RECT 169.920 174.240 170.240 174.560 ;
        RECT 170.320 174.240 170.640 174.560 ;
        RECT 170.720 174.240 171.040 174.560 ;
        RECT 171.120 174.240 171.440 174.560 ;
        RECT 171.520 174.240 171.840 174.560 ;
        RECT 171.920 174.240 172.240 174.560 ;
        RECT 172.320 174.240 172.640 174.560 ;
        RECT 172.720 174.240 173.040 174.560 ;
        RECT 173.120 174.240 173.440 174.560 ;
        RECT 173.520 174.240 173.840 174.560 ;
        RECT 173.920 174.240 174.240 174.560 ;
        RECT 174.320 174.240 174.640 174.560 ;
        RECT 174.720 174.240 175.040 174.560 ;
        RECT 175.120 174.240 175.440 174.560 ;
        RECT 175.520 174.240 175.840 174.560 ;
        RECT 175.920 174.240 176.240 174.560 ;
        RECT 176.320 174.240 176.640 174.560 ;
        RECT 176.720 174.240 177.040 174.560 ;
        RECT 177.120 174.240 177.440 174.560 ;
        RECT 177.520 174.240 177.840 174.560 ;
        RECT 177.920 174.240 178.240 174.560 ;
        RECT 178.320 174.240 178.640 174.560 ;
        RECT 178.720 174.240 179.040 174.560 ;
        RECT 179.120 174.240 179.440 174.560 ;
        RECT 179.520 174.240 179.840 174.560 ;
        RECT 179.920 174.240 180.240 174.560 ;
        RECT 180.320 174.240 180.640 174.560 ;
        RECT 25.040 173.840 25.360 174.160 ;
        RECT 25.440 173.840 25.760 174.160 ;
        RECT 25.840 173.840 26.160 174.160 ;
        RECT 26.240 173.840 26.560 174.160 ;
        RECT 26.640 173.840 26.960 174.160 ;
        RECT 27.040 173.840 27.360 174.160 ;
        RECT 27.440 173.840 27.760 174.160 ;
        RECT 27.840 173.840 28.160 174.160 ;
        RECT 28.240 173.840 28.560 174.160 ;
        RECT 28.640 173.840 28.960 174.160 ;
        RECT 29.040 173.840 29.360 174.160 ;
        RECT 29.440 173.840 29.760 174.160 ;
        RECT 29.840 173.840 30.160 174.160 ;
        RECT 30.240 173.840 30.560 174.160 ;
        RECT 30.640 173.840 30.960 174.160 ;
        RECT 31.040 173.840 31.360 174.160 ;
        RECT 31.440 173.840 31.760 174.160 ;
        RECT 31.840 173.840 32.160 174.160 ;
        RECT 32.240 173.840 32.560 174.160 ;
        RECT 32.640 173.840 32.960 174.160 ;
        RECT 33.040 173.840 33.360 174.160 ;
        RECT 33.440 173.840 33.760 174.160 ;
        RECT 33.840 173.840 34.160 174.160 ;
        RECT 34.240 173.840 34.560 174.160 ;
        RECT 34.640 173.840 34.960 174.160 ;
        RECT 35.040 173.840 35.360 174.160 ;
        RECT 35.440 173.840 35.760 174.160 ;
        RECT 35.840 173.840 36.160 174.160 ;
        RECT 36.240 173.840 36.560 174.160 ;
        RECT 36.640 173.840 36.960 174.160 ;
        RECT 37.040 173.840 37.360 174.160 ;
        RECT 37.440 173.840 37.760 174.160 ;
        RECT 37.840 173.840 38.160 174.160 ;
        RECT 38.240 173.840 38.560 174.160 ;
        RECT 38.640 173.840 38.960 174.160 ;
        RECT 39.040 173.840 39.360 174.160 ;
        RECT 39.440 173.840 39.760 174.160 ;
        RECT 39.840 173.840 40.160 174.160 ;
        RECT 40.240 173.840 40.560 174.160 ;
        RECT 40.640 173.840 40.960 174.160 ;
        RECT 41.040 173.840 41.360 174.160 ;
        RECT 41.440 173.840 41.760 174.160 ;
        RECT 41.840 173.840 42.160 174.160 ;
        RECT 42.240 173.840 42.560 174.160 ;
        RECT 42.640 173.840 42.960 174.160 ;
        RECT 43.040 173.840 43.360 174.160 ;
        RECT 43.440 173.840 43.760 174.160 ;
        RECT 43.840 173.840 44.160 174.160 ;
        RECT 44.240 173.840 44.560 174.160 ;
        RECT 44.640 173.840 44.960 174.160 ;
        RECT 70.560 173.840 70.880 174.160 ;
        RECT 70.960 173.840 71.280 174.160 ;
        RECT 71.360 173.840 71.680 174.160 ;
        RECT 71.760 173.840 72.080 174.160 ;
        RECT 120.560 173.840 120.880 174.160 ;
        RECT 120.960 173.840 121.280 174.160 ;
        RECT 121.360 173.840 121.680 174.160 ;
        RECT 121.760 173.840 122.080 174.160 ;
        RECT 160.720 173.840 161.040 174.160 ;
        RECT 161.120 173.840 161.440 174.160 ;
        RECT 161.520 173.840 161.840 174.160 ;
        RECT 161.920 173.840 162.240 174.160 ;
        RECT 162.320 173.840 162.640 174.160 ;
        RECT 162.720 173.840 163.040 174.160 ;
        RECT 163.120 173.840 163.440 174.160 ;
        RECT 163.520 173.840 163.840 174.160 ;
        RECT 163.920 173.840 164.240 174.160 ;
        RECT 164.320 173.840 164.640 174.160 ;
        RECT 164.720 173.840 165.040 174.160 ;
        RECT 165.120 173.840 165.440 174.160 ;
        RECT 165.520 173.840 165.840 174.160 ;
        RECT 165.920 173.840 166.240 174.160 ;
        RECT 166.320 173.840 166.640 174.160 ;
        RECT 166.720 173.840 167.040 174.160 ;
        RECT 167.120 173.840 167.440 174.160 ;
        RECT 167.520 173.840 167.840 174.160 ;
        RECT 167.920 173.840 168.240 174.160 ;
        RECT 168.320 173.840 168.640 174.160 ;
        RECT 168.720 173.840 169.040 174.160 ;
        RECT 169.120 173.840 169.440 174.160 ;
        RECT 169.520 173.840 169.840 174.160 ;
        RECT 169.920 173.840 170.240 174.160 ;
        RECT 170.320 173.840 170.640 174.160 ;
        RECT 170.720 173.840 171.040 174.160 ;
        RECT 171.120 173.840 171.440 174.160 ;
        RECT 171.520 173.840 171.840 174.160 ;
        RECT 171.920 173.840 172.240 174.160 ;
        RECT 172.320 173.840 172.640 174.160 ;
        RECT 172.720 173.840 173.040 174.160 ;
        RECT 173.120 173.840 173.440 174.160 ;
        RECT 173.520 173.840 173.840 174.160 ;
        RECT 173.920 173.840 174.240 174.160 ;
        RECT 174.320 173.840 174.640 174.160 ;
        RECT 174.720 173.840 175.040 174.160 ;
        RECT 175.120 173.840 175.440 174.160 ;
        RECT 175.520 173.840 175.840 174.160 ;
        RECT 175.920 173.840 176.240 174.160 ;
        RECT 176.320 173.840 176.640 174.160 ;
        RECT 176.720 173.840 177.040 174.160 ;
        RECT 177.120 173.840 177.440 174.160 ;
        RECT 177.520 173.840 177.840 174.160 ;
        RECT 177.920 173.840 178.240 174.160 ;
        RECT 178.320 173.840 178.640 174.160 ;
        RECT 178.720 173.840 179.040 174.160 ;
        RECT 179.120 173.840 179.440 174.160 ;
        RECT 179.520 173.840 179.840 174.160 ;
        RECT 179.920 173.840 180.240 174.160 ;
        RECT 180.320 173.840 180.640 174.160 ;
        RECT 25.040 173.440 25.360 173.760 ;
        RECT 25.440 173.440 25.760 173.760 ;
        RECT 25.840 173.440 26.160 173.760 ;
        RECT 26.240 173.440 26.560 173.760 ;
        RECT 26.640 173.440 26.960 173.760 ;
        RECT 27.040 173.440 27.360 173.760 ;
        RECT 27.440 173.440 27.760 173.760 ;
        RECT 27.840 173.440 28.160 173.760 ;
        RECT 28.240 173.440 28.560 173.760 ;
        RECT 28.640 173.440 28.960 173.760 ;
        RECT 29.040 173.440 29.360 173.760 ;
        RECT 29.440 173.440 29.760 173.760 ;
        RECT 29.840 173.440 30.160 173.760 ;
        RECT 30.240 173.440 30.560 173.760 ;
        RECT 30.640 173.440 30.960 173.760 ;
        RECT 31.040 173.440 31.360 173.760 ;
        RECT 31.440 173.440 31.760 173.760 ;
        RECT 31.840 173.440 32.160 173.760 ;
        RECT 32.240 173.440 32.560 173.760 ;
        RECT 32.640 173.440 32.960 173.760 ;
        RECT 33.040 173.440 33.360 173.760 ;
        RECT 33.440 173.440 33.760 173.760 ;
        RECT 33.840 173.440 34.160 173.760 ;
        RECT 34.240 173.440 34.560 173.760 ;
        RECT 34.640 173.440 34.960 173.760 ;
        RECT 35.040 173.440 35.360 173.760 ;
        RECT 35.440 173.440 35.760 173.760 ;
        RECT 35.840 173.440 36.160 173.760 ;
        RECT 36.240 173.440 36.560 173.760 ;
        RECT 36.640 173.440 36.960 173.760 ;
        RECT 37.040 173.440 37.360 173.760 ;
        RECT 37.440 173.440 37.760 173.760 ;
        RECT 37.840 173.440 38.160 173.760 ;
        RECT 38.240 173.440 38.560 173.760 ;
        RECT 38.640 173.440 38.960 173.760 ;
        RECT 39.040 173.440 39.360 173.760 ;
        RECT 39.440 173.440 39.760 173.760 ;
        RECT 39.840 173.440 40.160 173.760 ;
        RECT 40.240 173.440 40.560 173.760 ;
        RECT 40.640 173.440 40.960 173.760 ;
        RECT 41.040 173.440 41.360 173.760 ;
        RECT 41.440 173.440 41.760 173.760 ;
        RECT 41.840 173.440 42.160 173.760 ;
        RECT 42.240 173.440 42.560 173.760 ;
        RECT 42.640 173.440 42.960 173.760 ;
        RECT 43.040 173.440 43.360 173.760 ;
        RECT 43.440 173.440 43.760 173.760 ;
        RECT 43.840 173.440 44.160 173.760 ;
        RECT 44.240 173.440 44.560 173.760 ;
        RECT 44.640 173.440 44.960 173.760 ;
        RECT 70.560 173.440 70.880 173.760 ;
        RECT 70.960 173.440 71.280 173.760 ;
        RECT 71.360 173.440 71.680 173.760 ;
        RECT 71.760 173.440 72.080 173.760 ;
        RECT 120.560 173.440 120.880 173.760 ;
        RECT 120.960 173.440 121.280 173.760 ;
        RECT 121.360 173.440 121.680 173.760 ;
        RECT 121.760 173.440 122.080 173.760 ;
        RECT 160.720 173.440 161.040 173.760 ;
        RECT 161.120 173.440 161.440 173.760 ;
        RECT 161.520 173.440 161.840 173.760 ;
        RECT 161.920 173.440 162.240 173.760 ;
        RECT 162.320 173.440 162.640 173.760 ;
        RECT 162.720 173.440 163.040 173.760 ;
        RECT 163.120 173.440 163.440 173.760 ;
        RECT 163.520 173.440 163.840 173.760 ;
        RECT 163.920 173.440 164.240 173.760 ;
        RECT 164.320 173.440 164.640 173.760 ;
        RECT 164.720 173.440 165.040 173.760 ;
        RECT 165.120 173.440 165.440 173.760 ;
        RECT 165.520 173.440 165.840 173.760 ;
        RECT 165.920 173.440 166.240 173.760 ;
        RECT 166.320 173.440 166.640 173.760 ;
        RECT 166.720 173.440 167.040 173.760 ;
        RECT 167.120 173.440 167.440 173.760 ;
        RECT 167.520 173.440 167.840 173.760 ;
        RECT 167.920 173.440 168.240 173.760 ;
        RECT 168.320 173.440 168.640 173.760 ;
        RECT 168.720 173.440 169.040 173.760 ;
        RECT 169.120 173.440 169.440 173.760 ;
        RECT 169.520 173.440 169.840 173.760 ;
        RECT 169.920 173.440 170.240 173.760 ;
        RECT 170.320 173.440 170.640 173.760 ;
        RECT 170.720 173.440 171.040 173.760 ;
        RECT 171.120 173.440 171.440 173.760 ;
        RECT 171.520 173.440 171.840 173.760 ;
        RECT 171.920 173.440 172.240 173.760 ;
        RECT 172.320 173.440 172.640 173.760 ;
        RECT 172.720 173.440 173.040 173.760 ;
        RECT 173.120 173.440 173.440 173.760 ;
        RECT 173.520 173.440 173.840 173.760 ;
        RECT 173.920 173.440 174.240 173.760 ;
        RECT 174.320 173.440 174.640 173.760 ;
        RECT 174.720 173.440 175.040 173.760 ;
        RECT 175.120 173.440 175.440 173.760 ;
        RECT 175.520 173.440 175.840 173.760 ;
        RECT 175.920 173.440 176.240 173.760 ;
        RECT 176.320 173.440 176.640 173.760 ;
        RECT 176.720 173.440 177.040 173.760 ;
        RECT 177.120 173.440 177.440 173.760 ;
        RECT 177.520 173.440 177.840 173.760 ;
        RECT 177.920 173.440 178.240 173.760 ;
        RECT 178.320 173.440 178.640 173.760 ;
        RECT 178.720 173.440 179.040 173.760 ;
        RECT 179.120 173.440 179.440 173.760 ;
        RECT 179.520 173.440 179.840 173.760 ;
        RECT 179.920 173.440 180.240 173.760 ;
        RECT 180.320 173.440 180.640 173.760 ;
        RECT 25.040 173.040 25.360 173.360 ;
        RECT 25.440 173.040 25.760 173.360 ;
        RECT 25.840 173.040 26.160 173.360 ;
        RECT 26.240 173.040 26.560 173.360 ;
        RECT 26.640 173.040 26.960 173.360 ;
        RECT 27.040 173.040 27.360 173.360 ;
        RECT 27.440 173.040 27.760 173.360 ;
        RECT 27.840 173.040 28.160 173.360 ;
        RECT 28.240 173.040 28.560 173.360 ;
        RECT 28.640 173.040 28.960 173.360 ;
        RECT 29.040 173.040 29.360 173.360 ;
        RECT 29.440 173.040 29.760 173.360 ;
        RECT 29.840 173.040 30.160 173.360 ;
        RECT 30.240 173.040 30.560 173.360 ;
        RECT 30.640 173.040 30.960 173.360 ;
        RECT 31.040 173.040 31.360 173.360 ;
        RECT 31.440 173.040 31.760 173.360 ;
        RECT 31.840 173.040 32.160 173.360 ;
        RECT 32.240 173.040 32.560 173.360 ;
        RECT 32.640 173.040 32.960 173.360 ;
        RECT 33.040 173.040 33.360 173.360 ;
        RECT 33.440 173.040 33.760 173.360 ;
        RECT 33.840 173.040 34.160 173.360 ;
        RECT 34.240 173.040 34.560 173.360 ;
        RECT 34.640 173.040 34.960 173.360 ;
        RECT 35.040 173.040 35.360 173.360 ;
        RECT 35.440 173.040 35.760 173.360 ;
        RECT 35.840 173.040 36.160 173.360 ;
        RECT 36.240 173.040 36.560 173.360 ;
        RECT 36.640 173.040 36.960 173.360 ;
        RECT 37.040 173.040 37.360 173.360 ;
        RECT 37.440 173.040 37.760 173.360 ;
        RECT 37.840 173.040 38.160 173.360 ;
        RECT 38.240 173.040 38.560 173.360 ;
        RECT 38.640 173.040 38.960 173.360 ;
        RECT 39.040 173.040 39.360 173.360 ;
        RECT 39.440 173.040 39.760 173.360 ;
        RECT 39.840 173.040 40.160 173.360 ;
        RECT 40.240 173.040 40.560 173.360 ;
        RECT 40.640 173.040 40.960 173.360 ;
        RECT 41.040 173.040 41.360 173.360 ;
        RECT 41.440 173.040 41.760 173.360 ;
        RECT 41.840 173.040 42.160 173.360 ;
        RECT 42.240 173.040 42.560 173.360 ;
        RECT 42.640 173.040 42.960 173.360 ;
        RECT 43.040 173.040 43.360 173.360 ;
        RECT 43.440 173.040 43.760 173.360 ;
        RECT 43.840 173.040 44.160 173.360 ;
        RECT 44.240 173.040 44.560 173.360 ;
        RECT 44.640 173.040 44.960 173.360 ;
        RECT 70.560 173.040 70.880 173.360 ;
        RECT 70.960 173.040 71.280 173.360 ;
        RECT 71.360 173.040 71.680 173.360 ;
        RECT 71.760 173.040 72.080 173.360 ;
        RECT 120.560 173.040 120.880 173.360 ;
        RECT 120.960 173.040 121.280 173.360 ;
        RECT 121.360 173.040 121.680 173.360 ;
        RECT 121.760 173.040 122.080 173.360 ;
        RECT 160.720 173.040 161.040 173.360 ;
        RECT 161.120 173.040 161.440 173.360 ;
        RECT 161.520 173.040 161.840 173.360 ;
        RECT 161.920 173.040 162.240 173.360 ;
        RECT 162.320 173.040 162.640 173.360 ;
        RECT 162.720 173.040 163.040 173.360 ;
        RECT 163.120 173.040 163.440 173.360 ;
        RECT 163.520 173.040 163.840 173.360 ;
        RECT 163.920 173.040 164.240 173.360 ;
        RECT 164.320 173.040 164.640 173.360 ;
        RECT 164.720 173.040 165.040 173.360 ;
        RECT 165.120 173.040 165.440 173.360 ;
        RECT 165.520 173.040 165.840 173.360 ;
        RECT 165.920 173.040 166.240 173.360 ;
        RECT 166.320 173.040 166.640 173.360 ;
        RECT 166.720 173.040 167.040 173.360 ;
        RECT 167.120 173.040 167.440 173.360 ;
        RECT 167.520 173.040 167.840 173.360 ;
        RECT 167.920 173.040 168.240 173.360 ;
        RECT 168.320 173.040 168.640 173.360 ;
        RECT 168.720 173.040 169.040 173.360 ;
        RECT 169.120 173.040 169.440 173.360 ;
        RECT 169.520 173.040 169.840 173.360 ;
        RECT 169.920 173.040 170.240 173.360 ;
        RECT 170.320 173.040 170.640 173.360 ;
        RECT 170.720 173.040 171.040 173.360 ;
        RECT 171.120 173.040 171.440 173.360 ;
        RECT 171.520 173.040 171.840 173.360 ;
        RECT 171.920 173.040 172.240 173.360 ;
        RECT 172.320 173.040 172.640 173.360 ;
        RECT 172.720 173.040 173.040 173.360 ;
        RECT 173.120 173.040 173.440 173.360 ;
        RECT 173.520 173.040 173.840 173.360 ;
        RECT 173.920 173.040 174.240 173.360 ;
        RECT 174.320 173.040 174.640 173.360 ;
        RECT 174.720 173.040 175.040 173.360 ;
        RECT 175.120 173.040 175.440 173.360 ;
        RECT 175.520 173.040 175.840 173.360 ;
        RECT 175.920 173.040 176.240 173.360 ;
        RECT 176.320 173.040 176.640 173.360 ;
        RECT 176.720 173.040 177.040 173.360 ;
        RECT 177.120 173.040 177.440 173.360 ;
        RECT 177.520 173.040 177.840 173.360 ;
        RECT 177.920 173.040 178.240 173.360 ;
        RECT 178.320 173.040 178.640 173.360 ;
        RECT 178.720 173.040 179.040 173.360 ;
        RECT 179.120 173.040 179.440 173.360 ;
        RECT 179.520 173.040 179.840 173.360 ;
        RECT 179.920 173.040 180.240 173.360 ;
        RECT 180.320 173.040 180.640 173.360 ;
        RECT 25.040 172.640 25.360 172.960 ;
        RECT 25.440 172.640 25.760 172.960 ;
        RECT 25.840 172.640 26.160 172.960 ;
        RECT 26.240 172.640 26.560 172.960 ;
        RECT 26.640 172.640 26.960 172.960 ;
        RECT 27.040 172.640 27.360 172.960 ;
        RECT 27.440 172.640 27.760 172.960 ;
        RECT 27.840 172.640 28.160 172.960 ;
        RECT 28.240 172.640 28.560 172.960 ;
        RECT 28.640 172.640 28.960 172.960 ;
        RECT 29.040 172.640 29.360 172.960 ;
        RECT 29.440 172.640 29.760 172.960 ;
        RECT 29.840 172.640 30.160 172.960 ;
        RECT 30.240 172.640 30.560 172.960 ;
        RECT 30.640 172.640 30.960 172.960 ;
        RECT 31.040 172.640 31.360 172.960 ;
        RECT 31.440 172.640 31.760 172.960 ;
        RECT 31.840 172.640 32.160 172.960 ;
        RECT 32.240 172.640 32.560 172.960 ;
        RECT 32.640 172.640 32.960 172.960 ;
        RECT 33.040 172.640 33.360 172.960 ;
        RECT 33.440 172.640 33.760 172.960 ;
        RECT 33.840 172.640 34.160 172.960 ;
        RECT 34.240 172.640 34.560 172.960 ;
        RECT 34.640 172.640 34.960 172.960 ;
        RECT 35.040 172.640 35.360 172.960 ;
        RECT 35.440 172.640 35.760 172.960 ;
        RECT 35.840 172.640 36.160 172.960 ;
        RECT 36.240 172.640 36.560 172.960 ;
        RECT 36.640 172.640 36.960 172.960 ;
        RECT 37.040 172.640 37.360 172.960 ;
        RECT 37.440 172.640 37.760 172.960 ;
        RECT 37.840 172.640 38.160 172.960 ;
        RECT 38.240 172.640 38.560 172.960 ;
        RECT 38.640 172.640 38.960 172.960 ;
        RECT 39.040 172.640 39.360 172.960 ;
        RECT 39.440 172.640 39.760 172.960 ;
        RECT 39.840 172.640 40.160 172.960 ;
        RECT 40.240 172.640 40.560 172.960 ;
        RECT 40.640 172.640 40.960 172.960 ;
        RECT 41.040 172.640 41.360 172.960 ;
        RECT 41.440 172.640 41.760 172.960 ;
        RECT 41.840 172.640 42.160 172.960 ;
        RECT 42.240 172.640 42.560 172.960 ;
        RECT 42.640 172.640 42.960 172.960 ;
        RECT 43.040 172.640 43.360 172.960 ;
        RECT 43.440 172.640 43.760 172.960 ;
        RECT 43.840 172.640 44.160 172.960 ;
        RECT 44.240 172.640 44.560 172.960 ;
        RECT 44.640 172.640 44.960 172.960 ;
        RECT 70.560 172.640 70.880 172.960 ;
        RECT 70.960 172.640 71.280 172.960 ;
        RECT 71.360 172.640 71.680 172.960 ;
        RECT 71.760 172.640 72.080 172.960 ;
        RECT 120.560 172.640 120.880 172.960 ;
        RECT 120.960 172.640 121.280 172.960 ;
        RECT 121.360 172.640 121.680 172.960 ;
        RECT 121.760 172.640 122.080 172.960 ;
        RECT 160.720 172.640 161.040 172.960 ;
        RECT 161.120 172.640 161.440 172.960 ;
        RECT 161.520 172.640 161.840 172.960 ;
        RECT 161.920 172.640 162.240 172.960 ;
        RECT 162.320 172.640 162.640 172.960 ;
        RECT 162.720 172.640 163.040 172.960 ;
        RECT 163.120 172.640 163.440 172.960 ;
        RECT 163.520 172.640 163.840 172.960 ;
        RECT 163.920 172.640 164.240 172.960 ;
        RECT 164.320 172.640 164.640 172.960 ;
        RECT 164.720 172.640 165.040 172.960 ;
        RECT 165.120 172.640 165.440 172.960 ;
        RECT 165.520 172.640 165.840 172.960 ;
        RECT 165.920 172.640 166.240 172.960 ;
        RECT 166.320 172.640 166.640 172.960 ;
        RECT 166.720 172.640 167.040 172.960 ;
        RECT 167.120 172.640 167.440 172.960 ;
        RECT 167.520 172.640 167.840 172.960 ;
        RECT 167.920 172.640 168.240 172.960 ;
        RECT 168.320 172.640 168.640 172.960 ;
        RECT 168.720 172.640 169.040 172.960 ;
        RECT 169.120 172.640 169.440 172.960 ;
        RECT 169.520 172.640 169.840 172.960 ;
        RECT 169.920 172.640 170.240 172.960 ;
        RECT 170.320 172.640 170.640 172.960 ;
        RECT 170.720 172.640 171.040 172.960 ;
        RECT 171.120 172.640 171.440 172.960 ;
        RECT 171.520 172.640 171.840 172.960 ;
        RECT 171.920 172.640 172.240 172.960 ;
        RECT 172.320 172.640 172.640 172.960 ;
        RECT 172.720 172.640 173.040 172.960 ;
        RECT 173.120 172.640 173.440 172.960 ;
        RECT 173.520 172.640 173.840 172.960 ;
        RECT 173.920 172.640 174.240 172.960 ;
        RECT 174.320 172.640 174.640 172.960 ;
        RECT 174.720 172.640 175.040 172.960 ;
        RECT 175.120 172.640 175.440 172.960 ;
        RECT 175.520 172.640 175.840 172.960 ;
        RECT 175.920 172.640 176.240 172.960 ;
        RECT 176.320 172.640 176.640 172.960 ;
        RECT 176.720 172.640 177.040 172.960 ;
        RECT 177.120 172.640 177.440 172.960 ;
        RECT 177.520 172.640 177.840 172.960 ;
        RECT 177.920 172.640 178.240 172.960 ;
        RECT 178.320 172.640 178.640 172.960 ;
        RECT 178.720 172.640 179.040 172.960 ;
        RECT 179.120 172.640 179.440 172.960 ;
        RECT 179.520 172.640 179.840 172.960 ;
        RECT 179.920 172.640 180.240 172.960 ;
        RECT 180.320 172.640 180.640 172.960 ;
        RECT 25.040 172.240 25.360 172.560 ;
        RECT 25.440 172.240 25.760 172.560 ;
        RECT 25.840 172.240 26.160 172.560 ;
        RECT 26.240 172.240 26.560 172.560 ;
        RECT 26.640 172.240 26.960 172.560 ;
        RECT 27.040 172.240 27.360 172.560 ;
        RECT 27.440 172.240 27.760 172.560 ;
        RECT 27.840 172.240 28.160 172.560 ;
        RECT 28.240 172.240 28.560 172.560 ;
        RECT 28.640 172.240 28.960 172.560 ;
        RECT 29.040 172.240 29.360 172.560 ;
        RECT 29.440 172.240 29.760 172.560 ;
        RECT 29.840 172.240 30.160 172.560 ;
        RECT 30.240 172.240 30.560 172.560 ;
        RECT 30.640 172.240 30.960 172.560 ;
        RECT 31.040 172.240 31.360 172.560 ;
        RECT 31.440 172.240 31.760 172.560 ;
        RECT 31.840 172.240 32.160 172.560 ;
        RECT 32.240 172.240 32.560 172.560 ;
        RECT 32.640 172.240 32.960 172.560 ;
        RECT 33.040 172.240 33.360 172.560 ;
        RECT 33.440 172.240 33.760 172.560 ;
        RECT 33.840 172.240 34.160 172.560 ;
        RECT 34.240 172.240 34.560 172.560 ;
        RECT 34.640 172.240 34.960 172.560 ;
        RECT 35.040 172.240 35.360 172.560 ;
        RECT 35.440 172.240 35.760 172.560 ;
        RECT 35.840 172.240 36.160 172.560 ;
        RECT 36.240 172.240 36.560 172.560 ;
        RECT 36.640 172.240 36.960 172.560 ;
        RECT 37.040 172.240 37.360 172.560 ;
        RECT 37.440 172.240 37.760 172.560 ;
        RECT 37.840 172.240 38.160 172.560 ;
        RECT 38.240 172.240 38.560 172.560 ;
        RECT 38.640 172.240 38.960 172.560 ;
        RECT 39.040 172.240 39.360 172.560 ;
        RECT 39.440 172.240 39.760 172.560 ;
        RECT 39.840 172.240 40.160 172.560 ;
        RECT 40.240 172.240 40.560 172.560 ;
        RECT 40.640 172.240 40.960 172.560 ;
        RECT 41.040 172.240 41.360 172.560 ;
        RECT 41.440 172.240 41.760 172.560 ;
        RECT 41.840 172.240 42.160 172.560 ;
        RECT 42.240 172.240 42.560 172.560 ;
        RECT 42.640 172.240 42.960 172.560 ;
        RECT 43.040 172.240 43.360 172.560 ;
        RECT 43.440 172.240 43.760 172.560 ;
        RECT 43.840 172.240 44.160 172.560 ;
        RECT 44.240 172.240 44.560 172.560 ;
        RECT 44.640 172.240 44.960 172.560 ;
        RECT 70.560 172.240 70.880 172.560 ;
        RECT 70.960 172.240 71.280 172.560 ;
        RECT 71.360 172.240 71.680 172.560 ;
        RECT 71.760 172.240 72.080 172.560 ;
        RECT 120.560 172.240 120.880 172.560 ;
        RECT 120.960 172.240 121.280 172.560 ;
        RECT 121.360 172.240 121.680 172.560 ;
        RECT 121.760 172.240 122.080 172.560 ;
        RECT 160.720 172.240 161.040 172.560 ;
        RECT 161.120 172.240 161.440 172.560 ;
        RECT 161.520 172.240 161.840 172.560 ;
        RECT 161.920 172.240 162.240 172.560 ;
        RECT 162.320 172.240 162.640 172.560 ;
        RECT 162.720 172.240 163.040 172.560 ;
        RECT 163.120 172.240 163.440 172.560 ;
        RECT 163.520 172.240 163.840 172.560 ;
        RECT 163.920 172.240 164.240 172.560 ;
        RECT 164.320 172.240 164.640 172.560 ;
        RECT 164.720 172.240 165.040 172.560 ;
        RECT 165.120 172.240 165.440 172.560 ;
        RECT 165.520 172.240 165.840 172.560 ;
        RECT 165.920 172.240 166.240 172.560 ;
        RECT 166.320 172.240 166.640 172.560 ;
        RECT 166.720 172.240 167.040 172.560 ;
        RECT 167.120 172.240 167.440 172.560 ;
        RECT 167.520 172.240 167.840 172.560 ;
        RECT 167.920 172.240 168.240 172.560 ;
        RECT 168.320 172.240 168.640 172.560 ;
        RECT 168.720 172.240 169.040 172.560 ;
        RECT 169.120 172.240 169.440 172.560 ;
        RECT 169.520 172.240 169.840 172.560 ;
        RECT 169.920 172.240 170.240 172.560 ;
        RECT 170.320 172.240 170.640 172.560 ;
        RECT 170.720 172.240 171.040 172.560 ;
        RECT 171.120 172.240 171.440 172.560 ;
        RECT 171.520 172.240 171.840 172.560 ;
        RECT 171.920 172.240 172.240 172.560 ;
        RECT 172.320 172.240 172.640 172.560 ;
        RECT 172.720 172.240 173.040 172.560 ;
        RECT 173.120 172.240 173.440 172.560 ;
        RECT 173.520 172.240 173.840 172.560 ;
        RECT 173.920 172.240 174.240 172.560 ;
        RECT 174.320 172.240 174.640 172.560 ;
        RECT 174.720 172.240 175.040 172.560 ;
        RECT 175.120 172.240 175.440 172.560 ;
        RECT 175.520 172.240 175.840 172.560 ;
        RECT 175.920 172.240 176.240 172.560 ;
        RECT 176.320 172.240 176.640 172.560 ;
        RECT 176.720 172.240 177.040 172.560 ;
        RECT 177.120 172.240 177.440 172.560 ;
        RECT 177.520 172.240 177.840 172.560 ;
        RECT 177.920 172.240 178.240 172.560 ;
        RECT 178.320 172.240 178.640 172.560 ;
        RECT 178.720 172.240 179.040 172.560 ;
        RECT 179.120 172.240 179.440 172.560 ;
        RECT 179.520 172.240 179.840 172.560 ;
        RECT 179.920 172.240 180.240 172.560 ;
        RECT 180.320 172.240 180.640 172.560 ;
        RECT 25.040 171.840 25.360 172.160 ;
        RECT 25.440 171.840 25.760 172.160 ;
        RECT 25.840 171.840 26.160 172.160 ;
        RECT 26.240 171.840 26.560 172.160 ;
        RECT 26.640 171.840 26.960 172.160 ;
        RECT 27.040 171.840 27.360 172.160 ;
        RECT 27.440 171.840 27.760 172.160 ;
        RECT 27.840 171.840 28.160 172.160 ;
        RECT 28.240 171.840 28.560 172.160 ;
        RECT 28.640 171.840 28.960 172.160 ;
        RECT 29.040 171.840 29.360 172.160 ;
        RECT 29.440 171.840 29.760 172.160 ;
        RECT 29.840 171.840 30.160 172.160 ;
        RECT 30.240 171.840 30.560 172.160 ;
        RECT 30.640 171.840 30.960 172.160 ;
        RECT 31.040 171.840 31.360 172.160 ;
        RECT 31.440 171.840 31.760 172.160 ;
        RECT 31.840 171.840 32.160 172.160 ;
        RECT 32.240 171.840 32.560 172.160 ;
        RECT 32.640 171.840 32.960 172.160 ;
        RECT 33.040 171.840 33.360 172.160 ;
        RECT 33.440 171.840 33.760 172.160 ;
        RECT 33.840 171.840 34.160 172.160 ;
        RECT 34.240 171.840 34.560 172.160 ;
        RECT 34.640 171.840 34.960 172.160 ;
        RECT 35.040 171.840 35.360 172.160 ;
        RECT 35.440 171.840 35.760 172.160 ;
        RECT 35.840 171.840 36.160 172.160 ;
        RECT 36.240 171.840 36.560 172.160 ;
        RECT 36.640 171.840 36.960 172.160 ;
        RECT 37.040 171.840 37.360 172.160 ;
        RECT 37.440 171.840 37.760 172.160 ;
        RECT 37.840 171.840 38.160 172.160 ;
        RECT 38.240 171.840 38.560 172.160 ;
        RECT 38.640 171.840 38.960 172.160 ;
        RECT 39.040 171.840 39.360 172.160 ;
        RECT 39.440 171.840 39.760 172.160 ;
        RECT 39.840 171.840 40.160 172.160 ;
        RECT 40.240 171.840 40.560 172.160 ;
        RECT 40.640 171.840 40.960 172.160 ;
        RECT 41.040 171.840 41.360 172.160 ;
        RECT 41.440 171.840 41.760 172.160 ;
        RECT 41.840 171.840 42.160 172.160 ;
        RECT 42.240 171.840 42.560 172.160 ;
        RECT 42.640 171.840 42.960 172.160 ;
        RECT 43.040 171.840 43.360 172.160 ;
        RECT 43.440 171.840 43.760 172.160 ;
        RECT 43.840 171.840 44.160 172.160 ;
        RECT 44.240 171.840 44.560 172.160 ;
        RECT 44.640 171.840 44.960 172.160 ;
        RECT 70.560 171.840 70.880 172.160 ;
        RECT 70.960 171.840 71.280 172.160 ;
        RECT 71.360 171.840 71.680 172.160 ;
        RECT 71.760 171.840 72.080 172.160 ;
        RECT 120.560 171.840 120.880 172.160 ;
        RECT 120.960 171.840 121.280 172.160 ;
        RECT 121.360 171.840 121.680 172.160 ;
        RECT 121.760 171.840 122.080 172.160 ;
        RECT 160.720 171.840 161.040 172.160 ;
        RECT 161.120 171.840 161.440 172.160 ;
        RECT 161.520 171.840 161.840 172.160 ;
        RECT 161.920 171.840 162.240 172.160 ;
        RECT 162.320 171.840 162.640 172.160 ;
        RECT 162.720 171.840 163.040 172.160 ;
        RECT 163.120 171.840 163.440 172.160 ;
        RECT 163.520 171.840 163.840 172.160 ;
        RECT 163.920 171.840 164.240 172.160 ;
        RECT 164.320 171.840 164.640 172.160 ;
        RECT 164.720 171.840 165.040 172.160 ;
        RECT 165.120 171.840 165.440 172.160 ;
        RECT 165.520 171.840 165.840 172.160 ;
        RECT 165.920 171.840 166.240 172.160 ;
        RECT 166.320 171.840 166.640 172.160 ;
        RECT 166.720 171.840 167.040 172.160 ;
        RECT 167.120 171.840 167.440 172.160 ;
        RECT 167.520 171.840 167.840 172.160 ;
        RECT 167.920 171.840 168.240 172.160 ;
        RECT 168.320 171.840 168.640 172.160 ;
        RECT 168.720 171.840 169.040 172.160 ;
        RECT 169.120 171.840 169.440 172.160 ;
        RECT 169.520 171.840 169.840 172.160 ;
        RECT 169.920 171.840 170.240 172.160 ;
        RECT 170.320 171.840 170.640 172.160 ;
        RECT 170.720 171.840 171.040 172.160 ;
        RECT 171.120 171.840 171.440 172.160 ;
        RECT 171.520 171.840 171.840 172.160 ;
        RECT 171.920 171.840 172.240 172.160 ;
        RECT 172.320 171.840 172.640 172.160 ;
        RECT 172.720 171.840 173.040 172.160 ;
        RECT 173.120 171.840 173.440 172.160 ;
        RECT 173.520 171.840 173.840 172.160 ;
        RECT 173.920 171.840 174.240 172.160 ;
        RECT 174.320 171.840 174.640 172.160 ;
        RECT 174.720 171.840 175.040 172.160 ;
        RECT 175.120 171.840 175.440 172.160 ;
        RECT 175.520 171.840 175.840 172.160 ;
        RECT 175.920 171.840 176.240 172.160 ;
        RECT 176.320 171.840 176.640 172.160 ;
        RECT 176.720 171.840 177.040 172.160 ;
        RECT 177.120 171.840 177.440 172.160 ;
        RECT 177.520 171.840 177.840 172.160 ;
        RECT 177.920 171.840 178.240 172.160 ;
        RECT 178.320 171.840 178.640 172.160 ;
        RECT 178.720 171.840 179.040 172.160 ;
        RECT 179.120 171.840 179.440 172.160 ;
        RECT 179.520 171.840 179.840 172.160 ;
        RECT 179.920 171.840 180.240 172.160 ;
        RECT 180.320 171.840 180.640 172.160 ;
        RECT 25.040 171.440 25.360 171.760 ;
        RECT 25.440 171.440 25.760 171.760 ;
        RECT 25.840 171.440 26.160 171.760 ;
        RECT 26.240 171.440 26.560 171.760 ;
        RECT 26.640 171.440 26.960 171.760 ;
        RECT 27.040 171.440 27.360 171.760 ;
        RECT 27.440 171.440 27.760 171.760 ;
        RECT 27.840 171.440 28.160 171.760 ;
        RECT 28.240 171.440 28.560 171.760 ;
        RECT 28.640 171.440 28.960 171.760 ;
        RECT 29.040 171.440 29.360 171.760 ;
        RECT 29.440 171.440 29.760 171.760 ;
        RECT 29.840 171.440 30.160 171.760 ;
        RECT 30.240 171.440 30.560 171.760 ;
        RECT 30.640 171.440 30.960 171.760 ;
        RECT 31.040 171.440 31.360 171.760 ;
        RECT 31.440 171.440 31.760 171.760 ;
        RECT 31.840 171.440 32.160 171.760 ;
        RECT 32.240 171.440 32.560 171.760 ;
        RECT 32.640 171.440 32.960 171.760 ;
        RECT 33.040 171.440 33.360 171.760 ;
        RECT 33.440 171.440 33.760 171.760 ;
        RECT 33.840 171.440 34.160 171.760 ;
        RECT 34.240 171.440 34.560 171.760 ;
        RECT 34.640 171.440 34.960 171.760 ;
        RECT 35.040 171.440 35.360 171.760 ;
        RECT 35.440 171.440 35.760 171.760 ;
        RECT 35.840 171.440 36.160 171.760 ;
        RECT 36.240 171.440 36.560 171.760 ;
        RECT 36.640 171.440 36.960 171.760 ;
        RECT 37.040 171.440 37.360 171.760 ;
        RECT 37.440 171.440 37.760 171.760 ;
        RECT 37.840 171.440 38.160 171.760 ;
        RECT 38.240 171.440 38.560 171.760 ;
        RECT 38.640 171.440 38.960 171.760 ;
        RECT 39.040 171.440 39.360 171.760 ;
        RECT 39.440 171.440 39.760 171.760 ;
        RECT 39.840 171.440 40.160 171.760 ;
        RECT 40.240 171.440 40.560 171.760 ;
        RECT 40.640 171.440 40.960 171.760 ;
        RECT 41.040 171.440 41.360 171.760 ;
        RECT 41.440 171.440 41.760 171.760 ;
        RECT 41.840 171.440 42.160 171.760 ;
        RECT 42.240 171.440 42.560 171.760 ;
        RECT 42.640 171.440 42.960 171.760 ;
        RECT 43.040 171.440 43.360 171.760 ;
        RECT 43.440 171.440 43.760 171.760 ;
        RECT 43.840 171.440 44.160 171.760 ;
        RECT 44.240 171.440 44.560 171.760 ;
        RECT 44.640 171.440 44.960 171.760 ;
        RECT 70.560 171.440 70.880 171.760 ;
        RECT 70.960 171.440 71.280 171.760 ;
        RECT 71.360 171.440 71.680 171.760 ;
        RECT 71.760 171.440 72.080 171.760 ;
        RECT 120.560 171.440 120.880 171.760 ;
        RECT 120.960 171.440 121.280 171.760 ;
        RECT 121.360 171.440 121.680 171.760 ;
        RECT 121.760 171.440 122.080 171.760 ;
        RECT 160.720 171.440 161.040 171.760 ;
        RECT 161.120 171.440 161.440 171.760 ;
        RECT 161.520 171.440 161.840 171.760 ;
        RECT 161.920 171.440 162.240 171.760 ;
        RECT 162.320 171.440 162.640 171.760 ;
        RECT 162.720 171.440 163.040 171.760 ;
        RECT 163.120 171.440 163.440 171.760 ;
        RECT 163.520 171.440 163.840 171.760 ;
        RECT 163.920 171.440 164.240 171.760 ;
        RECT 164.320 171.440 164.640 171.760 ;
        RECT 164.720 171.440 165.040 171.760 ;
        RECT 165.120 171.440 165.440 171.760 ;
        RECT 165.520 171.440 165.840 171.760 ;
        RECT 165.920 171.440 166.240 171.760 ;
        RECT 166.320 171.440 166.640 171.760 ;
        RECT 166.720 171.440 167.040 171.760 ;
        RECT 167.120 171.440 167.440 171.760 ;
        RECT 167.520 171.440 167.840 171.760 ;
        RECT 167.920 171.440 168.240 171.760 ;
        RECT 168.320 171.440 168.640 171.760 ;
        RECT 168.720 171.440 169.040 171.760 ;
        RECT 169.120 171.440 169.440 171.760 ;
        RECT 169.520 171.440 169.840 171.760 ;
        RECT 169.920 171.440 170.240 171.760 ;
        RECT 170.320 171.440 170.640 171.760 ;
        RECT 170.720 171.440 171.040 171.760 ;
        RECT 171.120 171.440 171.440 171.760 ;
        RECT 171.520 171.440 171.840 171.760 ;
        RECT 171.920 171.440 172.240 171.760 ;
        RECT 172.320 171.440 172.640 171.760 ;
        RECT 172.720 171.440 173.040 171.760 ;
        RECT 173.120 171.440 173.440 171.760 ;
        RECT 173.520 171.440 173.840 171.760 ;
        RECT 173.920 171.440 174.240 171.760 ;
        RECT 174.320 171.440 174.640 171.760 ;
        RECT 174.720 171.440 175.040 171.760 ;
        RECT 175.120 171.440 175.440 171.760 ;
        RECT 175.520 171.440 175.840 171.760 ;
        RECT 175.920 171.440 176.240 171.760 ;
        RECT 176.320 171.440 176.640 171.760 ;
        RECT 176.720 171.440 177.040 171.760 ;
        RECT 177.120 171.440 177.440 171.760 ;
        RECT 177.520 171.440 177.840 171.760 ;
        RECT 177.920 171.440 178.240 171.760 ;
        RECT 178.320 171.440 178.640 171.760 ;
        RECT 178.720 171.440 179.040 171.760 ;
        RECT 179.120 171.440 179.440 171.760 ;
        RECT 179.520 171.440 179.840 171.760 ;
        RECT 179.920 171.440 180.240 171.760 ;
        RECT 180.320 171.440 180.640 171.760 ;
        RECT 25.040 171.040 25.360 171.360 ;
        RECT 25.440 171.040 25.760 171.360 ;
        RECT 25.840 171.040 26.160 171.360 ;
        RECT 26.240 171.040 26.560 171.360 ;
        RECT 26.640 171.040 26.960 171.360 ;
        RECT 27.040 171.040 27.360 171.360 ;
        RECT 27.440 171.040 27.760 171.360 ;
        RECT 27.840 171.040 28.160 171.360 ;
        RECT 28.240 171.040 28.560 171.360 ;
        RECT 28.640 171.040 28.960 171.360 ;
        RECT 29.040 171.040 29.360 171.360 ;
        RECT 29.440 171.040 29.760 171.360 ;
        RECT 29.840 171.040 30.160 171.360 ;
        RECT 30.240 171.040 30.560 171.360 ;
        RECT 30.640 171.040 30.960 171.360 ;
        RECT 31.040 171.040 31.360 171.360 ;
        RECT 31.440 171.040 31.760 171.360 ;
        RECT 31.840 171.040 32.160 171.360 ;
        RECT 32.240 171.040 32.560 171.360 ;
        RECT 32.640 171.040 32.960 171.360 ;
        RECT 33.040 171.040 33.360 171.360 ;
        RECT 33.440 171.040 33.760 171.360 ;
        RECT 33.840 171.040 34.160 171.360 ;
        RECT 34.240 171.040 34.560 171.360 ;
        RECT 34.640 171.040 34.960 171.360 ;
        RECT 35.040 171.040 35.360 171.360 ;
        RECT 35.440 171.040 35.760 171.360 ;
        RECT 35.840 171.040 36.160 171.360 ;
        RECT 36.240 171.040 36.560 171.360 ;
        RECT 36.640 171.040 36.960 171.360 ;
        RECT 37.040 171.040 37.360 171.360 ;
        RECT 37.440 171.040 37.760 171.360 ;
        RECT 37.840 171.040 38.160 171.360 ;
        RECT 38.240 171.040 38.560 171.360 ;
        RECT 38.640 171.040 38.960 171.360 ;
        RECT 39.040 171.040 39.360 171.360 ;
        RECT 39.440 171.040 39.760 171.360 ;
        RECT 39.840 171.040 40.160 171.360 ;
        RECT 40.240 171.040 40.560 171.360 ;
        RECT 40.640 171.040 40.960 171.360 ;
        RECT 41.040 171.040 41.360 171.360 ;
        RECT 41.440 171.040 41.760 171.360 ;
        RECT 41.840 171.040 42.160 171.360 ;
        RECT 42.240 171.040 42.560 171.360 ;
        RECT 42.640 171.040 42.960 171.360 ;
        RECT 43.040 171.040 43.360 171.360 ;
        RECT 43.440 171.040 43.760 171.360 ;
        RECT 43.840 171.040 44.160 171.360 ;
        RECT 44.240 171.040 44.560 171.360 ;
        RECT 44.640 171.040 44.960 171.360 ;
        RECT 70.560 171.040 70.880 171.360 ;
        RECT 70.960 171.040 71.280 171.360 ;
        RECT 71.360 171.040 71.680 171.360 ;
        RECT 71.760 171.040 72.080 171.360 ;
        RECT 120.560 171.040 120.880 171.360 ;
        RECT 120.960 171.040 121.280 171.360 ;
        RECT 121.360 171.040 121.680 171.360 ;
        RECT 121.760 171.040 122.080 171.360 ;
        RECT 160.720 171.040 161.040 171.360 ;
        RECT 161.120 171.040 161.440 171.360 ;
        RECT 161.520 171.040 161.840 171.360 ;
        RECT 161.920 171.040 162.240 171.360 ;
        RECT 162.320 171.040 162.640 171.360 ;
        RECT 162.720 171.040 163.040 171.360 ;
        RECT 163.120 171.040 163.440 171.360 ;
        RECT 163.520 171.040 163.840 171.360 ;
        RECT 163.920 171.040 164.240 171.360 ;
        RECT 164.320 171.040 164.640 171.360 ;
        RECT 164.720 171.040 165.040 171.360 ;
        RECT 165.120 171.040 165.440 171.360 ;
        RECT 165.520 171.040 165.840 171.360 ;
        RECT 165.920 171.040 166.240 171.360 ;
        RECT 166.320 171.040 166.640 171.360 ;
        RECT 166.720 171.040 167.040 171.360 ;
        RECT 167.120 171.040 167.440 171.360 ;
        RECT 167.520 171.040 167.840 171.360 ;
        RECT 167.920 171.040 168.240 171.360 ;
        RECT 168.320 171.040 168.640 171.360 ;
        RECT 168.720 171.040 169.040 171.360 ;
        RECT 169.120 171.040 169.440 171.360 ;
        RECT 169.520 171.040 169.840 171.360 ;
        RECT 169.920 171.040 170.240 171.360 ;
        RECT 170.320 171.040 170.640 171.360 ;
        RECT 170.720 171.040 171.040 171.360 ;
        RECT 171.120 171.040 171.440 171.360 ;
        RECT 171.520 171.040 171.840 171.360 ;
        RECT 171.920 171.040 172.240 171.360 ;
        RECT 172.320 171.040 172.640 171.360 ;
        RECT 172.720 171.040 173.040 171.360 ;
        RECT 173.120 171.040 173.440 171.360 ;
        RECT 173.520 171.040 173.840 171.360 ;
        RECT 173.920 171.040 174.240 171.360 ;
        RECT 174.320 171.040 174.640 171.360 ;
        RECT 174.720 171.040 175.040 171.360 ;
        RECT 175.120 171.040 175.440 171.360 ;
        RECT 175.520 171.040 175.840 171.360 ;
        RECT 175.920 171.040 176.240 171.360 ;
        RECT 176.320 171.040 176.640 171.360 ;
        RECT 176.720 171.040 177.040 171.360 ;
        RECT 177.120 171.040 177.440 171.360 ;
        RECT 177.520 171.040 177.840 171.360 ;
        RECT 177.920 171.040 178.240 171.360 ;
        RECT 178.320 171.040 178.640 171.360 ;
        RECT 178.720 171.040 179.040 171.360 ;
        RECT 179.120 171.040 179.440 171.360 ;
        RECT 179.520 171.040 179.840 171.360 ;
        RECT 179.920 171.040 180.240 171.360 ;
        RECT 180.320 171.040 180.640 171.360 ;
        RECT 25.040 170.640 25.360 170.960 ;
        RECT 25.440 170.640 25.760 170.960 ;
        RECT 25.840 170.640 26.160 170.960 ;
        RECT 26.240 170.640 26.560 170.960 ;
        RECT 26.640 170.640 26.960 170.960 ;
        RECT 27.040 170.640 27.360 170.960 ;
        RECT 27.440 170.640 27.760 170.960 ;
        RECT 27.840 170.640 28.160 170.960 ;
        RECT 28.240 170.640 28.560 170.960 ;
        RECT 28.640 170.640 28.960 170.960 ;
        RECT 29.040 170.640 29.360 170.960 ;
        RECT 29.440 170.640 29.760 170.960 ;
        RECT 29.840 170.640 30.160 170.960 ;
        RECT 30.240 170.640 30.560 170.960 ;
        RECT 30.640 170.640 30.960 170.960 ;
        RECT 31.040 170.640 31.360 170.960 ;
        RECT 31.440 170.640 31.760 170.960 ;
        RECT 31.840 170.640 32.160 170.960 ;
        RECT 32.240 170.640 32.560 170.960 ;
        RECT 32.640 170.640 32.960 170.960 ;
        RECT 33.040 170.640 33.360 170.960 ;
        RECT 33.440 170.640 33.760 170.960 ;
        RECT 33.840 170.640 34.160 170.960 ;
        RECT 34.240 170.640 34.560 170.960 ;
        RECT 34.640 170.640 34.960 170.960 ;
        RECT 35.040 170.640 35.360 170.960 ;
        RECT 35.440 170.640 35.760 170.960 ;
        RECT 35.840 170.640 36.160 170.960 ;
        RECT 36.240 170.640 36.560 170.960 ;
        RECT 36.640 170.640 36.960 170.960 ;
        RECT 37.040 170.640 37.360 170.960 ;
        RECT 37.440 170.640 37.760 170.960 ;
        RECT 37.840 170.640 38.160 170.960 ;
        RECT 38.240 170.640 38.560 170.960 ;
        RECT 38.640 170.640 38.960 170.960 ;
        RECT 39.040 170.640 39.360 170.960 ;
        RECT 39.440 170.640 39.760 170.960 ;
        RECT 39.840 170.640 40.160 170.960 ;
        RECT 40.240 170.640 40.560 170.960 ;
        RECT 40.640 170.640 40.960 170.960 ;
        RECT 41.040 170.640 41.360 170.960 ;
        RECT 41.440 170.640 41.760 170.960 ;
        RECT 41.840 170.640 42.160 170.960 ;
        RECT 42.240 170.640 42.560 170.960 ;
        RECT 42.640 170.640 42.960 170.960 ;
        RECT 43.040 170.640 43.360 170.960 ;
        RECT 43.440 170.640 43.760 170.960 ;
        RECT 43.840 170.640 44.160 170.960 ;
        RECT 44.240 170.640 44.560 170.960 ;
        RECT 44.640 170.640 44.960 170.960 ;
        RECT 70.560 170.640 70.880 170.960 ;
        RECT 70.960 170.640 71.280 170.960 ;
        RECT 71.360 170.640 71.680 170.960 ;
        RECT 71.760 170.640 72.080 170.960 ;
        RECT 120.560 170.640 120.880 170.960 ;
        RECT 120.960 170.640 121.280 170.960 ;
        RECT 121.360 170.640 121.680 170.960 ;
        RECT 121.760 170.640 122.080 170.960 ;
        RECT 160.720 170.640 161.040 170.960 ;
        RECT 161.120 170.640 161.440 170.960 ;
        RECT 161.520 170.640 161.840 170.960 ;
        RECT 161.920 170.640 162.240 170.960 ;
        RECT 162.320 170.640 162.640 170.960 ;
        RECT 162.720 170.640 163.040 170.960 ;
        RECT 163.120 170.640 163.440 170.960 ;
        RECT 163.520 170.640 163.840 170.960 ;
        RECT 163.920 170.640 164.240 170.960 ;
        RECT 164.320 170.640 164.640 170.960 ;
        RECT 164.720 170.640 165.040 170.960 ;
        RECT 165.120 170.640 165.440 170.960 ;
        RECT 165.520 170.640 165.840 170.960 ;
        RECT 165.920 170.640 166.240 170.960 ;
        RECT 166.320 170.640 166.640 170.960 ;
        RECT 166.720 170.640 167.040 170.960 ;
        RECT 167.120 170.640 167.440 170.960 ;
        RECT 167.520 170.640 167.840 170.960 ;
        RECT 167.920 170.640 168.240 170.960 ;
        RECT 168.320 170.640 168.640 170.960 ;
        RECT 168.720 170.640 169.040 170.960 ;
        RECT 169.120 170.640 169.440 170.960 ;
        RECT 169.520 170.640 169.840 170.960 ;
        RECT 169.920 170.640 170.240 170.960 ;
        RECT 170.320 170.640 170.640 170.960 ;
        RECT 170.720 170.640 171.040 170.960 ;
        RECT 171.120 170.640 171.440 170.960 ;
        RECT 171.520 170.640 171.840 170.960 ;
        RECT 171.920 170.640 172.240 170.960 ;
        RECT 172.320 170.640 172.640 170.960 ;
        RECT 172.720 170.640 173.040 170.960 ;
        RECT 173.120 170.640 173.440 170.960 ;
        RECT 173.520 170.640 173.840 170.960 ;
        RECT 173.920 170.640 174.240 170.960 ;
        RECT 174.320 170.640 174.640 170.960 ;
        RECT 174.720 170.640 175.040 170.960 ;
        RECT 175.120 170.640 175.440 170.960 ;
        RECT 175.520 170.640 175.840 170.960 ;
        RECT 175.920 170.640 176.240 170.960 ;
        RECT 176.320 170.640 176.640 170.960 ;
        RECT 176.720 170.640 177.040 170.960 ;
        RECT 177.120 170.640 177.440 170.960 ;
        RECT 177.520 170.640 177.840 170.960 ;
        RECT 177.920 170.640 178.240 170.960 ;
        RECT 178.320 170.640 178.640 170.960 ;
        RECT 178.720 170.640 179.040 170.960 ;
        RECT 179.120 170.640 179.440 170.960 ;
        RECT 179.520 170.640 179.840 170.960 ;
        RECT 179.920 170.640 180.240 170.960 ;
        RECT 180.320 170.640 180.640 170.960 ;
        RECT 25.040 170.240 25.360 170.560 ;
        RECT 25.440 170.240 25.760 170.560 ;
        RECT 25.840 170.240 26.160 170.560 ;
        RECT 26.240 170.240 26.560 170.560 ;
        RECT 26.640 170.240 26.960 170.560 ;
        RECT 27.040 170.240 27.360 170.560 ;
        RECT 27.440 170.240 27.760 170.560 ;
        RECT 27.840 170.240 28.160 170.560 ;
        RECT 28.240 170.240 28.560 170.560 ;
        RECT 28.640 170.240 28.960 170.560 ;
        RECT 29.040 170.240 29.360 170.560 ;
        RECT 29.440 170.240 29.760 170.560 ;
        RECT 29.840 170.240 30.160 170.560 ;
        RECT 30.240 170.240 30.560 170.560 ;
        RECT 30.640 170.240 30.960 170.560 ;
        RECT 31.040 170.240 31.360 170.560 ;
        RECT 31.440 170.240 31.760 170.560 ;
        RECT 31.840 170.240 32.160 170.560 ;
        RECT 32.240 170.240 32.560 170.560 ;
        RECT 32.640 170.240 32.960 170.560 ;
        RECT 33.040 170.240 33.360 170.560 ;
        RECT 33.440 170.240 33.760 170.560 ;
        RECT 33.840 170.240 34.160 170.560 ;
        RECT 34.240 170.240 34.560 170.560 ;
        RECT 34.640 170.240 34.960 170.560 ;
        RECT 35.040 170.240 35.360 170.560 ;
        RECT 35.440 170.240 35.760 170.560 ;
        RECT 35.840 170.240 36.160 170.560 ;
        RECT 36.240 170.240 36.560 170.560 ;
        RECT 36.640 170.240 36.960 170.560 ;
        RECT 37.040 170.240 37.360 170.560 ;
        RECT 37.440 170.240 37.760 170.560 ;
        RECT 37.840 170.240 38.160 170.560 ;
        RECT 38.240 170.240 38.560 170.560 ;
        RECT 38.640 170.240 38.960 170.560 ;
        RECT 39.040 170.240 39.360 170.560 ;
        RECT 39.440 170.240 39.760 170.560 ;
        RECT 39.840 170.240 40.160 170.560 ;
        RECT 40.240 170.240 40.560 170.560 ;
        RECT 40.640 170.240 40.960 170.560 ;
        RECT 41.040 170.240 41.360 170.560 ;
        RECT 41.440 170.240 41.760 170.560 ;
        RECT 41.840 170.240 42.160 170.560 ;
        RECT 42.240 170.240 42.560 170.560 ;
        RECT 42.640 170.240 42.960 170.560 ;
        RECT 43.040 170.240 43.360 170.560 ;
        RECT 43.440 170.240 43.760 170.560 ;
        RECT 43.840 170.240 44.160 170.560 ;
        RECT 44.240 170.240 44.560 170.560 ;
        RECT 44.640 170.240 44.960 170.560 ;
        RECT 70.560 170.240 70.880 170.560 ;
        RECT 70.960 170.240 71.280 170.560 ;
        RECT 71.360 170.240 71.680 170.560 ;
        RECT 71.760 170.240 72.080 170.560 ;
        RECT 120.560 170.240 120.880 170.560 ;
        RECT 120.960 170.240 121.280 170.560 ;
        RECT 121.360 170.240 121.680 170.560 ;
        RECT 121.760 170.240 122.080 170.560 ;
        RECT 160.720 170.240 161.040 170.560 ;
        RECT 161.120 170.240 161.440 170.560 ;
        RECT 161.520 170.240 161.840 170.560 ;
        RECT 161.920 170.240 162.240 170.560 ;
        RECT 162.320 170.240 162.640 170.560 ;
        RECT 162.720 170.240 163.040 170.560 ;
        RECT 163.120 170.240 163.440 170.560 ;
        RECT 163.520 170.240 163.840 170.560 ;
        RECT 163.920 170.240 164.240 170.560 ;
        RECT 164.320 170.240 164.640 170.560 ;
        RECT 164.720 170.240 165.040 170.560 ;
        RECT 165.120 170.240 165.440 170.560 ;
        RECT 165.520 170.240 165.840 170.560 ;
        RECT 165.920 170.240 166.240 170.560 ;
        RECT 166.320 170.240 166.640 170.560 ;
        RECT 166.720 170.240 167.040 170.560 ;
        RECT 167.120 170.240 167.440 170.560 ;
        RECT 167.520 170.240 167.840 170.560 ;
        RECT 167.920 170.240 168.240 170.560 ;
        RECT 168.320 170.240 168.640 170.560 ;
        RECT 168.720 170.240 169.040 170.560 ;
        RECT 169.120 170.240 169.440 170.560 ;
        RECT 169.520 170.240 169.840 170.560 ;
        RECT 169.920 170.240 170.240 170.560 ;
        RECT 170.320 170.240 170.640 170.560 ;
        RECT 170.720 170.240 171.040 170.560 ;
        RECT 171.120 170.240 171.440 170.560 ;
        RECT 171.520 170.240 171.840 170.560 ;
        RECT 171.920 170.240 172.240 170.560 ;
        RECT 172.320 170.240 172.640 170.560 ;
        RECT 172.720 170.240 173.040 170.560 ;
        RECT 173.120 170.240 173.440 170.560 ;
        RECT 173.520 170.240 173.840 170.560 ;
        RECT 173.920 170.240 174.240 170.560 ;
        RECT 174.320 170.240 174.640 170.560 ;
        RECT 174.720 170.240 175.040 170.560 ;
        RECT 175.120 170.240 175.440 170.560 ;
        RECT 175.520 170.240 175.840 170.560 ;
        RECT 175.920 170.240 176.240 170.560 ;
        RECT 176.320 170.240 176.640 170.560 ;
        RECT 176.720 170.240 177.040 170.560 ;
        RECT 177.120 170.240 177.440 170.560 ;
        RECT 177.520 170.240 177.840 170.560 ;
        RECT 177.920 170.240 178.240 170.560 ;
        RECT 178.320 170.240 178.640 170.560 ;
        RECT 178.720 170.240 179.040 170.560 ;
        RECT 179.120 170.240 179.440 170.560 ;
        RECT 179.520 170.240 179.840 170.560 ;
        RECT 179.920 170.240 180.240 170.560 ;
        RECT 180.320 170.240 180.640 170.560 ;
        RECT 25.040 169.840 25.360 170.160 ;
        RECT 25.440 169.840 25.760 170.160 ;
        RECT 25.840 169.840 26.160 170.160 ;
        RECT 26.240 169.840 26.560 170.160 ;
        RECT 26.640 169.840 26.960 170.160 ;
        RECT 27.040 169.840 27.360 170.160 ;
        RECT 27.440 169.840 27.760 170.160 ;
        RECT 27.840 169.840 28.160 170.160 ;
        RECT 28.240 169.840 28.560 170.160 ;
        RECT 28.640 169.840 28.960 170.160 ;
        RECT 29.040 169.840 29.360 170.160 ;
        RECT 29.440 169.840 29.760 170.160 ;
        RECT 29.840 169.840 30.160 170.160 ;
        RECT 30.240 169.840 30.560 170.160 ;
        RECT 30.640 169.840 30.960 170.160 ;
        RECT 31.040 169.840 31.360 170.160 ;
        RECT 31.440 169.840 31.760 170.160 ;
        RECT 31.840 169.840 32.160 170.160 ;
        RECT 32.240 169.840 32.560 170.160 ;
        RECT 32.640 169.840 32.960 170.160 ;
        RECT 33.040 169.840 33.360 170.160 ;
        RECT 33.440 169.840 33.760 170.160 ;
        RECT 33.840 169.840 34.160 170.160 ;
        RECT 34.240 169.840 34.560 170.160 ;
        RECT 34.640 169.840 34.960 170.160 ;
        RECT 35.040 169.840 35.360 170.160 ;
        RECT 35.440 169.840 35.760 170.160 ;
        RECT 35.840 169.840 36.160 170.160 ;
        RECT 36.240 169.840 36.560 170.160 ;
        RECT 36.640 169.840 36.960 170.160 ;
        RECT 37.040 169.840 37.360 170.160 ;
        RECT 37.440 169.840 37.760 170.160 ;
        RECT 37.840 169.840 38.160 170.160 ;
        RECT 38.240 169.840 38.560 170.160 ;
        RECT 38.640 169.840 38.960 170.160 ;
        RECT 39.040 169.840 39.360 170.160 ;
        RECT 39.440 169.840 39.760 170.160 ;
        RECT 39.840 169.840 40.160 170.160 ;
        RECT 40.240 169.840 40.560 170.160 ;
        RECT 40.640 169.840 40.960 170.160 ;
        RECT 41.040 169.840 41.360 170.160 ;
        RECT 41.440 169.840 41.760 170.160 ;
        RECT 41.840 169.840 42.160 170.160 ;
        RECT 42.240 169.840 42.560 170.160 ;
        RECT 42.640 169.840 42.960 170.160 ;
        RECT 43.040 169.840 43.360 170.160 ;
        RECT 43.440 169.840 43.760 170.160 ;
        RECT 43.840 169.840 44.160 170.160 ;
        RECT 44.240 169.840 44.560 170.160 ;
        RECT 44.640 169.840 44.960 170.160 ;
        RECT 70.560 169.840 70.880 170.160 ;
        RECT 70.960 169.840 71.280 170.160 ;
        RECT 71.360 169.840 71.680 170.160 ;
        RECT 71.760 169.840 72.080 170.160 ;
        RECT 120.560 169.840 120.880 170.160 ;
        RECT 120.960 169.840 121.280 170.160 ;
        RECT 121.360 169.840 121.680 170.160 ;
        RECT 121.760 169.840 122.080 170.160 ;
        RECT 160.720 169.840 161.040 170.160 ;
        RECT 161.120 169.840 161.440 170.160 ;
        RECT 161.520 169.840 161.840 170.160 ;
        RECT 161.920 169.840 162.240 170.160 ;
        RECT 162.320 169.840 162.640 170.160 ;
        RECT 162.720 169.840 163.040 170.160 ;
        RECT 163.120 169.840 163.440 170.160 ;
        RECT 163.520 169.840 163.840 170.160 ;
        RECT 163.920 169.840 164.240 170.160 ;
        RECT 164.320 169.840 164.640 170.160 ;
        RECT 164.720 169.840 165.040 170.160 ;
        RECT 165.120 169.840 165.440 170.160 ;
        RECT 165.520 169.840 165.840 170.160 ;
        RECT 165.920 169.840 166.240 170.160 ;
        RECT 166.320 169.840 166.640 170.160 ;
        RECT 166.720 169.840 167.040 170.160 ;
        RECT 167.120 169.840 167.440 170.160 ;
        RECT 167.520 169.840 167.840 170.160 ;
        RECT 167.920 169.840 168.240 170.160 ;
        RECT 168.320 169.840 168.640 170.160 ;
        RECT 168.720 169.840 169.040 170.160 ;
        RECT 169.120 169.840 169.440 170.160 ;
        RECT 169.520 169.840 169.840 170.160 ;
        RECT 169.920 169.840 170.240 170.160 ;
        RECT 170.320 169.840 170.640 170.160 ;
        RECT 170.720 169.840 171.040 170.160 ;
        RECT 171.120 169.840 171.440 170.160 ;
        RECT 171.520 169.840 171.840 170.160 ;
        RECT 171.920 169.840 172.240 170.160 ;
        RECT 172.320 169.840 172.640 170.160 ;
        RECT 172.720 169.840 173.040 170.160 ;
        RECT 173.120 169.840 173.440 170.160 ;
        RECT 173.520 169.840 173.840 170.160 ;
        RECT 173.920 169.840 174.240 170.160 ;
        RECT 174.320 169.840 174.640 170.160 ;
        RECT 174.720 169.840 175.040 170.160 ;
        RECT 175.120 169.840 175.440 170.160 ;
        RECT 175.520 169.840 175.840 170.160 ;
        RECT 175.920 169.840 176.240 170.160 ;
        RECT 176.320 169.840 176.640 170.160 ;
        RECT 176.720 169.840 177.040 170.160 ;
        RECT 177.120 169.840 177.440 170.160 ;
        RECT 177.520 169.840 177.840 170.160 ;
        RECT 177.920 169.840 178.240 170.160 ;
        RECT 178.320 169.840 178.640 170.160 ;
        RECT 178.720 169.840 179.040 170.160 ;
        RECT 179.120 169.840 179.440 170.160 ;
        RECT 179.520 169.840 179.840 170.160 ;
        RECT 179.920 169.840 180.240 170.160 ;
        RECT 180.320 169.840 180.640 170.160 ;
        RECT 25.040 169.440 25.360 169.760 ;
        RECT 25.440 169.440 25.760 169.760 ;
        RECT 25.840 169.440 26.160 169.760 ;
        RECT 26.240 169.440 26.560 169.760 ;
        RECT 26.640 169.440 26.960 169.760 ;
        RECT 27.040 169.440 27.360 169.760 ;
        RECT 27.440 169.440 27.760 169.760 ;
        RECT 27.840 169.440 28.160 169.760 ;
        RECT 28.240 169.440 28.560 169.760 ;
        RECT 28.640 169.440 28.960 169.760 ;
        RECT 29.040 169.440 29.360 169.760 ;
        RECT 29.440 169.440 29.760 169.760 ;
        RECT 29.840 169.440 30.160 169.760 ;
        RECT 30.240 169.440 30.560 169.760 ;
        RECT 30.640 169.440 30.960 169.760 ;
        RECT 31.040 169.440 31.360 169.760 ;
        RECT 31.440 169.440 31.760 169.760 ;
        RECT 31.840 169.440 32.160 169.760 ;
        RECT 32.240 169.440 32.560 169.760 ;
        RECT 32.640 169.440 32.960 169.760 ;
        RECT 33.040 169.440 33.360 169.760 ;
        RECT 33.440 169.440 33.760 169.760 ;
        RECT 33.840 169.440 34.160 169.760 ;
        RECT 34.240 169.440 34.560 169.760 ;
        RECT 34.640 169.440 34.960 169.760 ;
        RECT 35.040 169.440 35.360 169.760 ;
        RECT 35.440 169.440 35.760 169.760 ;
        RECT 35.840 169.440 36.160 169.760 ;
        RECT 36.240 169.440 36.560 169.760 ;
        RECT 36.640 169.440 36.960 169.760 ;
        RECT 37.040 169.440 37.360 169.760 ;
        RECT 37.440 169.440 37.760 169.760 ;
        RECT 37.840 169.440 38.160 169.760 ;
        RECT 38.240 169.440 38.560 169.760 ;
        RECT 38.640 169.440 38.960 169.760 ;
        RECT 39.040 169.440 39.360 169.760 ;
        RECT 39.440 169.440 39.760 169.760 ;
        RECT 39.840 169.440 40.160 169.760 ;
        RECT 40.240 169.440 40.560 169.760 ;
        RECT 40.640 169.440 40.960 169.760 ;
        RECT 41.040 169.440 41.360 169.760 ;
        RECT 41.440 169.440 41.760 169.760 ;
        RECT 41.840 169.440 42.160 169.760 ;
        RECT 42.240 169.440 42.560 169.760 ;
        RECT 42.640 169.440 42.960 169.760 ;
        RECT 43.040 169.440 43.360 169.760 ;
        RECT 43.440 169.440 43.760 169.760 ;
        RECT 43.840 169.440 44.160 169.760 ;
        RECT 44.240 169.440 44.560 169.760 ;
        RECT 44.640 169.440 44.960 169.760 ;
        RECT 70.560 169.440 70.880 169.760 ;
        RECT 70.960 169.440 71.280 169.760 ;
        RECT 71.360 169.440 71.680 169.760 ;
        RECT 71.760 169.440 72.080 169.760 ;
        RECT 120.560 169.440 120.880 169.760 ;
        RECT 120.960 169.440 121.280 169.760 ;
        RECT 121.360 169.440 121.680 169.760 ;
        RECT 121.760 169.440 122.080 169.760 ;
        RECT 160.720 169.440 161.040 169.760 ;
        RECT 161.120 169.440 161.440 169.760 ;
        RECT 161.520 169.440 161.840 169.760 ;
        RECT 161.920 169.440 162.240 169.760 ;
        RECT 162.320 169.440 162.640 169.760 ;
        RECT 162.720 169.440 163.040 169.760 ;
        RECT 163.120 169.440 163.440 169.760 ;
        RECT 163.520 169.440 163.840 169.760 ;
        RECT 163.920 169.440 164.240 169.760 ;
        RECT 164.320 169.440 164.640 169.760 ;
        RECT 164.720 169.440 165.040 169.760 ;
        RECT 165.120 169.440 165.440 169.760 ;
        RECT 165.520 169.440 165.840 169.760 ;
        RECT 165.920 169.440 166.240 169.760 ;
        RECT 166.320 169.440 166.640 169.760 ;
        RECT 166.720 169.440 167.040 169.760 ;
        RECT 167.120 169.440 167.440 169.760 ;
        RECT 167.520 169.440 167.840 169.760 ;
        RECT 167.920 169.440 168.240 169.760 ;
        RECT 168.320 169.440 168.640 169.760 ;
        RECT 168.720 169.440 169.040 169.760 ;
        RECT 169.120 169.440 169.440 169.760 ;
        RECT 169.520 169.440 169.840 169.760 ;
        RECT 169.920 169.440 170.240 169.760 ;
        RECT 170.320 169.440 170.640 169.760 ;
        RECT 170.720 169.440 171.040 169.760 ;
        RECT 171.120 169.440 171.440 169.760 ;
        RECT 171.520 169.440 171.840 169.760 ;
        RECT 171.920 169.440 172.240 169.760 ;
        RECT 172.320 169.440 172.640 169.760 ;
        RECT 172.720 169.440 173.040 169.760 ;
        RECT 173.120 169.440 173.440 169.760 ;
        RECT 173.520 169.440 173.840 169.760 ;
        RECT 173.920 169.440 174.240 169.760 ;
        RECT 174.320 169.440 174.640 169.760 ;
        RECT 174.720 169.440 175.040 169.760 ;
        RECT 175.120 169.440 175.440 169.760 ;
        RECT 175.520 169.440 175.840 169.760 ;
        RECT 175.920 169.440 176.240 169.760 ;
        RECT 176.320 169.440 176.640 169.760 ;
        RECT 176.720 169.440 177.040 169.760 ;
        RECT 177.120 169.440 177.440 169.760 ;
        RECT 177.520 169.440 177.840 169.760 ;
        RECT 177.920 169.440 178.240 169.760 ;
        RECT 178.320 169.440 178.640 169.760 ;
        RECT 178.720 169.440 179.040 169.760 ;
        RECT 179.120 169.440 179.440 169.760 ;
        RECT 179.520 169.440 179.840 169.760 ;
        RECT 179.920 169.440 180.240 169.760 ;
        RECT 180.320 169.440 180.640 169.760 ;
        RECT 25.040 169.040 25.360 169.360 ;
        RECT 25.440 169.040 25.760 169.360 ;
        RECT 25.840 169.040 26.160 169.360 ;
        RECT 26.240 169.040 26.560 169.360 ;
        RECT 26.640 169.040 26.960 169.360 ;
        RECT 27.040 169.040 27.360 169.360 ;
        RECT 27.440 169.040 27.760 169.360 ;
        RECT 27.840 169.040 28.160 169.360 ;
        RECT 28.240 169.040 28.560 169.360 ;
        RECT 28.640 169.040 28.960 169.360 ;
        RECT 29.040 169.040 29.360 169.360 ;
        RECT 29.440 169.040 29.760 169.360 ;
        RECT 29.840 169.040 30.160 169.360 ;
        RECT 30.240 169.040 30.560 169.360 ;
        RECT 30.640 169.040 30.960 169.360 ;
        RECT 31.040 169.040 31.360 169.360 ;
        RECT 31.440 169.040 31.760 169.360 ;
        RECT 31.840 169.040 32.160 169.360 ;
        RECT 32.240 169.040 32.560 169.360 ;
        RECT 32.640 169.040 32.960 169.360 ;
        RECT 33.040 169.040 33.360 169.360 ;
        RECT 33.440 169.040 33.760 169.360 ;
        RECT 33.840 169.040 34.160 169.360 ;
        RECT 34.240 169.040 34.560 169.360 ;
        RECT 34.640 169.040 34.960 169.360 ;
        RECT 35.040 169.040 35.360 169.360 ;
        RECT 35.440 169.040 35.760 169.360 ;
        RECT 35.840 169.040 36.160 169.360 ;
        RECT 36.240 169.040 36.560 169.360 ;
        RECT 36.640 169.040 36.960 169.360 ;
        RECT 37.040 169.040 37.360 169.360 ;
        RECT 37.440 169.040 37.760 169.360 ;
        RECT 37.840 169.040 38.160 169.360 ;
        RECT 38.240 169.040 38.560 169.360 ;
        RECT 38.640 169.040 38.960 169.360 ;
        RECT 39.040 169.040 39.360 169.360 ;
        RECT 39.440 169.040 39.760 169.360 ;
        RECT 39.840 169.040 40.160 169.360 ;
        RECT 40.240 169.040 40.560 169.360 ;
        RECT 40.640 169.040 40.960 169.360 ;
        RECT 41.040 169.040 41.360 169.360 ;
        RECT 41.440 169.040 41.760 169.360 ;
        RECT 41.840 169.040 42.160 169.360 ;
        RECT 42.240 169.040 42.560 169.360 ;
        RECT 42.640 169.040 42.960 169.360 ;
        RECT 43.040 169.040 43.360 169.360 ;
        RECT 43.440 169.040 43.760 169.360 ;
        RECT 43.840 169.040 44.160 169.360 ;
        RECT 44.240 169.040 44.560 169.360 ;
        RECT 44.640 169.040 44.960 169.360 ;
        RECT 70.560 169.040 70.880 169.360 ;
        RECT 70.960 169.040 71.280 169.360 ;
        RECT 71.360 169.040 71.680 169.360 ;
        RECT 71.760 169.040 72.080 169.360 ;
        RECT 120.560 169.040 120.880 169.360 ;
        RECT 120.960 169.040 121.280 169.360 ;
        RECT 121.360 169.040 121.680 169.360 ;
        RECT 121.760 169.040 122.080 169.360 ;
        RECT 160.720 169.040 161.040 169.360 ;
        RECT 161.120 169.040 161.440 169.360 ;
        RECT 161.520 169.040 161.840 169.360 ;
        RECT 161.920 169.040 162.240 169.360 ;
        RECT 162.320 169.040 162.640 169.360 ;
        RECT 162.720 169.040 163.040 169.360 ;
        RECT 163.120 169.040 163.440 169.360 ;
        RECT 163.520 169.040 163.840 169.360 ;
        RECT 163.920 169.040 164.240 169.360 ;
        RECT 164.320 169.040 164.640 169.360 ;
        RECT 164.720 169.040 165.040 169.360 ;
        RECT 165.120 169.040 165.440 169.360 ;
        RECT 165.520 169.040 165.840 169.360 ;
        RECT 165.920 169.040 166.240 169.360 ;
        RECT 166.320 169.040 166.640 169.360 ;
        RECT 166.720 169.040 167.040 169.360 ;
        RECT 167.120 169.040 167.440 169.360 ;
        RECT 167.520 169.040 167.840 169.360 ;
        RECT 167.920 169.040 168.240 169.360 ;
        RECT 168.320 169.040 168.640 169.360 ;
        RECT 168.720 169.040 169.040 169.360 ;
        RECT 169.120 169.040 169.440 169.360 ;
        RECT 169.520 169.040 169.840 169.360 ;
        RECT 169.920 169.040 170.240 169.360 ;
        RECT 170.320 169.040 170.640 169.360 ;
        RECT 170.720 169.040 171.040 169.360 ;
        RECT 171.120 169.040 171.440 169.360 ;
        RECT 171.520 169.040 171.840 169.360 ;
        RECT 171.920 169.040 172.240 169.360 ;
        RECT 172.320 169.040 172.640 169.360 ;
        RECT 172.720 169.040 173.040 169.360 ;
        RECT 173.120 169.040 173.440 169.360 ;
        RECT 173.520 169.040 173.840 169.360 ;
        RECT 173.920 169.040 174.240 169.360 ;
        RECT 174.320 169.040 174.640 169.360 ;
        RECT 174.720 169.040 175.040 169.360 ;
        RECT 175.120 169.040 175.440 169.360 ;
        RECT 175.520 169.040 175.840 169.360 ;
        RECT 175.920 169.040 176.240 169.360 ;
        RECT 176.320 169.040 176.640 169.360 ;
        RECT 176.720 169.040 177.040 169.360 ;
        RECT 177.120 169.040 177.440 169.360 ;
        RECT 177.520 169.040 177.840 169.360 ;
        RECT 177.920 169.040 178.240 169.360 ;
        RECT 178.320 169.040 178.640 169.360 ;
        RECT 178.720 169.040 179.040 169.360 ;
        RECT 179.120 169.040 179.440 169.360 ;
        RECT 179.520 169.040 179.840 169.360 ;
        RECT 179.920 169.040 180.240 169.360 ;
        RECT 180.320 169.040 180.640 169.360 ;
        RECT 25.040 168.640 25.360 168.960 ;
        RECT 25.440 168.640 25.760 168.960 ;
        RECT 25.840 168.640 26.160 168.960 ;
        RECT 26.240 168.640 26.560 168.960 ;
        RECT 26.640 168.640 26.960 168.960 ;
        RECT 27.040 168.640 27.360 168.960 ;
        RECT 27.440 168.640 27.760 168.960 ;
        RECT 27.840 168.640 28.160 168.960 ;
        RECT 28.240 168.640 28.560 168.960 ;
        RECT 28.640 168.640 28.960 168.960 ;
        RECT 29.040 168.640 29.360 168.960 ;
        RECT 29.440 168.640 29.760 168.960 ;
        RECT 29.840 168.640 30.160 168.960 ;
        RECT 30.240 168.640 30.560 168.960 ;
        RECT 30.640 168.640 30.960 168.960 ;
        RECT 31.040 168.640 31.360 168.960 ;
        RECT 31.440 168.640 31.760 168.960 ;
        RECT 31.840 168.640 32.160 168.960 ;
        RECT 32.240 168.640 32.560 168.960 ;
        RECT 32.640 168.640 32.960 168.960 ;
        RECT 33.040 168.640 33.360 168.960 ;
        RECT 33.440 168.640 33.760 168.960 ;
        RECT 33.840 168.640 34.160 168.960 ;
        RECT 34.240 168.640 34.560 168.960 ;
        RECT 34.640 168.640 34.960 168.960 ;
        RECT 35.040 168.640 35.360 168.960 ;
        RECT 35.440 168.640 35.760 168.960 ;
        RECT 35.840 168.640 36.160 168.960 ;
        RECT 36.240 168.640 36.560 168.960 ;
        RECT 36.640 168.640 36.960 168.960 ;
        RECT 37.040 168.640 37.360 168.960 ;
        RECT 37.440 168.640 37.760 168.960 ;
        RECT 37.840 168.640 38.160 168.960 ;
        RECT 38.240 168.640 38.560 168.960 ;
        RECT 38.640 168.640 38.960 168.960 ;
        RECT 39.040 168.640 39.360 168.960 ;
        RECT 39.440 168.640 39.760 168.960 ;
        RECT 39.840 168.640 40.160 168.960 ;
        RECT 40.240 168.640 40.560 168.960 ;
        RECT 40.640 168.640 40.960 168.960 ;
        RECT 41.040 168.640 41.360 168.960 ;
        RECT 41.440 168.640 41.760 168.960 ;
        RECT 41.840 168.640 42.160 168.960 ;
        RECT 42.240 168.640 42.560 168.960 ;
        RECT 42.640 168.640 42.960 168.960 ;
        RECT 43.040 168.640 43.360 168.960 ;
        RECT 43.440 168.640 43.760 168.960 ;
        RECT 43.840 168.640 44.160 168.960 ;
        RECT 44.240 168.640 44.560 168.960 ;
        RECT 44.640 168.640 44.960 168.960 ;
        RECT 70.560 168.640 70.880 168.960 ;
        RECT 70.960 168.640 71.280 168.960 ;
        RECT 71.360 168.640 71.680 168.960 ;
        RECT 71.760 168.640 72.080 168.960 ;
        RECT 120.560 168.640 120.880 168.960 ;
        RECT 120.960 168.640 121.280 168.960 ;
        RECT 121.360 168.640 121.680 168.960 ;
        RECT 121.760 168.640 122.080 168.960 ;
        RECT 160.720 168.640 161.040 168.960 ;
        RECT 161.120 168.640 161.440 168.960 ;
        RECT 161.520 168.640 161.840 168.960 ;
        RECT 161.920 168.640 162.240 168.960 ;
        RECT 162.320 168.640 162.640 168.960 ;
        RECT 162.720 168.640 163.040 168.960 ;
        RECT 163.120 168.640 163.440 168.960 ;
        RECT 163.520 168.640 163.840 168.960 ;
        RECT 163.920 168.640 164.240 168.960 ;
        RECT 164.320 168.640 164.640 168.960 ;
        RECT 164.720 168.640 165.040 168.960 ;
        RECT 165.120 168.640 165.440 168.960 ;
        RECT 165.520 168.640 165.840 168.960 ;
        RECT 165.920 168.640 166.240 168.960 ;
        RECT 166.320 168.640 166.640 168.960 ;
        RECT 166.720 168.640 167.040 168.960 ;
        RECT 167.120 168.640 167.440 168.960 ;
        RECT 167.520 168.640 167.840 168.960 ;
        RECT 167.920 168.640 168.240 168.960 ;
        RECT 168.320 168.640 168.640 168.960 ;
        RECT 168.720 168.640 169.040 168.960 ;
        RECT 169.120 168.640 169.440 168.960 ;
        RECT 169.520 168.640 169.840 168.960 ;
        RECT 169.920 168.640 170.240 168.960 ;
        RECT 170.320 168.640 170.640 168.960 ;
        RECT 170.720 168.640 171.040 168.960 ;
        RECT 171.120 168.640 171.440 168.960 ;
        RECT 171.520 168.640 171.840 168.960 ;
        RECT 171.920 168.640 172.240 168.960 ;
        RECT 172.320 168.640 172.640 168.960 ;
        RECT 172.720 168.640 173.040 168.960 ;
        RECT 173.120 168.640 173.440 168.960 ;
        RECT 173.520 168.640 173.840 168.960 ;
        RECT 173.920 168.640 174.240 168.960 ;
        RECT 174.320 168.640 174.640 168.960 ;
        RECT 174.720 168.640 175.040 168.960 ;
        RECT 175.120 168.640 175.440 168.960 ;
        RECT 175.520 168.640 175.840 168.960 ;
        RECT 175.920 168.640 176.240 168.960 ;
        RECT 176.320 168.640 176.640 168.960 ;
        RECT 176.720 168.640 177.040 168.960 ;
        RECT 177.120 168.640 177.440 168.960 ;
        RECT 177.520 168.640 177.840 168.960 ;
        RECT 177.920 168.640 178.240 168.960 ;
        RECT 178.320 168.640 178.640 168.960 ;
        RECT 178.720 168.640 179.040 168.960 ;
        RECT 179.120 168.640 179.440 168.960 ;
        RECT 179.520 168.640 179.840 168.960 ;
        RECT 179.920 168.640 180.240 168.960 ;
        RECT 180.320 168.640 180.640 168.960 ;
        RECT 25.040 168.240 25.360 168.560 ;
        RECT 25.440 168.240 25.760 168.560 ;
        RECT 25.840 168.240 26.160 168.560 ;
        RECT 26.240 168.240 26.560 168.560 ;
        RECT 26.640 168.240 26.960 168.560 ;
        RECT 27.040 168.240 27.360 168.560 ;
        RECT 27.440 168.240 27.760 168.560 ;
        RECT 27.840 168.240 28.160 168.560 ;
        RECT 28.240 168.240 28.560 168.560 ;
        RECT 28.640 168.240 28.960 168.560 ;
        RECT 29.040 168.240 29.360 168.560 ;
        RECT 29.440 168.240 29.760 168.560 ;
        RECT 29.840 168.240 30.160 168.560 ;
        RECT 30.240 168.240 30.560 168.560 ;
        RECT 30.640 168.240 30.960 168.560 ;
        RECT 31.040 168.240 31.360 168.560 ;
        RECT 31.440 168.240 31.760 168.560 ;
        RECT 31.840 168.240 32.160 168.560 ;
        RECT 32.240 168.240 32.560 168.560 ;
        RECT 32.640 168.240 32.960 168.560 ;
        RECT 33.040 168.240 33.360 168.560 ;
        RECT 33.440 168.240 33.760 168.560 ;
        RECT 33.840 168.240 34.160 168.560 ;
        RECT 34.240 168.240 34.560 168.560 ;
        RECT 34.640 168.240 34.960 168.560 ;
        RECT 35.040 168.240 35.360 168.560 ;
        RECT 35.440 168.240 35.760 168.560 ;
        RECT 35.840 168.240 36.160 168.560 ;
        RECT 36.240 168.240 36.560 168.560 ;
        RECT 36.640 168.240 36.960 168.560 ;
        RECT 37.040 168.240 37.360 168.560 ;
        RECT 37.440 168.240 37.760 168.560 ;
        RECT 37.840 168.240 38.160 168.560 ;
        RECT 38.240 168.240 38.560 168.560 ;
        RECT 38.640 168.240 38.960 168.560 ;
        RECT 39.040 168.240 39.360 168.560 ;
        RECT 39.440 168.240 39.760 168.560 ;
        RECT 39.840 168.240 40.160 168.560 ;
        RECT 40.240 168.240 40.560 168.560 ;
        RECT 40.640 168.240 40.960 168.560 ;
        RECT 41.040 168.240 41.360 168.560 ;
        RECT 41.440 168.240 41.760 168.560 ;
        RECT 41.840 168.240 42.160 168.560 ;
        RECT 42.240 168.240 42.560 168.560 ;
        RECT 42.640 168.240 42.960 168.560 ;
        RECT 43.040 168.240 43.360 168.560 ;
        RECT 43.440 168.240 43.760 168.560 ;
        RECT 43.840 168.240 44.160 168.560 ;
        RECT 44.240 168.240 44.560 168.560 ;
        RECT 44.640 168.240 44.960 168.560 ;
        RECT 70.560 168.240 70.880 168.560 ;
        RECT 70.960 168.240 71.280 168.560 ;
        RECT 71.360 168.240 71.680 168.560 ;
        RECT 71.760 168.240 72.080 168.560 ;
        RECT 120.560 168.240 120.880 168.560 ;
        RECT 120.960 168.240 121.280 168.560 ;
        RECT 121.360 168.240 121.680 168.560 ;
        RECT 121.760 168.240 122.080 168.560 ;
        RECT 160.720 168.240 161.040 168.560 ;
        RECT 161.120 168.240 161.440 168.560 ;
        RECT 161.520 168.240 161.840 168.560 ;
        RECT 161.920 168.240 162.240 168.560 ;
        RECT 162.320 168.240 162.640 168.560 ;
        RECT 162.720 168.240 163.040 168.560 ;
        RECT 163.120 168.240 163.440 168.560 ;
        RECT 163.520 168.240 163.840 168.560 ;
        RECT 163.920 168.240 164.240 168.560 ;
        RECT 164.320 168.240 164.640 168.560 ;
        RECT 164.720 168.240 165.040 168.560 ;
        RECT 165.120 168.240 165.440 168.560 ;
        RECT 165.520 168.240 165.840 168.560 ;
        RECT 165.920 168.240 166.240 168.560 ;
        RECT 166.320 168.240 166.640 168.560 ;
        RECT 166.720 168.240 167.040 168.560 ;
        RECT 167.120 168.240 167.440 168.560 ;
        RECT 167.520 168.240 167.840 168.560 ;
        RECT 167.920 168.240 168.240 168.560 ;
        RECT 168.320 168.240 168.640 168.560 ;
        RECT 168.720 168.240 169.040 168.560 ;
        RECT 169.120 168.240 169.440 168.560 ;
        RECT 169.520 168.240 169.840 168.560 ;
        RECT 169.920 168.240 170.240 168.560 ;
        RECT 170.320 168.240 170.640 168.560 ;
        RECT 170.720 168.240 171.040 168.560 ;
        RECT 171.120 168.240 171.440 168.560 ;
        RECT 171.520 168.240 171.840 168.560 ;
        RECT 171.920 168.240 172.240 168.560 ;
        RECT 172.320 168.240 172.640 168.560 ;
        RECT 172.720 168.240 173.040 168.560 ;
        RECT 173.120 168.240 173.440 168.560 ;
        RECT 173.520 168.240 173.840 168.560 ;
        RECT 173.920 168.240 174.240 168.560 ;
        RECT 174.320 168.240 174.640 168.560 ;
        RECT 174.720 168.240 175.040 168.560 ;
        RECT 175.120 168.240 175.440 168.560 ;
        RECT 175.520 168.240 175.840 168.560 ;
        RECT 175.920 168.240 176.240 168.560 ;
        RECT 176.320 168.240 176.640 168.560 ;
        RECT 176.720 168.240 177.040 168.560 ;
        RECT 177.120 168.240 177.440 168.560 ;
        RECT 177.520 168.240 177.840 168.560 ;
        RECT 177.920 168.240 178.240 168.560 ;
        RECT 178.320 168.240 178.640 168.560 ;
        RECT 178.720 168.240 179.040 168.560 ;
        RECT 179.120 168.240 179.440 168.560 ;
        RECT 179.520 168.240 179.840 168.560 ;
        RECT 179.920 168.240 180.240 168.560 ;
        RECT 180.320 168.240 180.640 168.560 ;
        RECT 25.040 167.840 25.360 168.160 ;
        RECT 25.440 167.840 25.760 168.160 ;
        RECT 25.840 167.840 26.160 168.160 ;
        RECT 26.240 167.840 26.560 168.160 ;
        RECT 26.640 167.840 26.960 168.160 ;
        RECT 27.040 167.840 27.360 168.160 ;
        RECT 27.440 167.840 27.760 168.160 ;
        RECT 27.840 167.840 28.160 168.160 ;
        RECT 28.240 167.840 28.560 168.160 ;
        RECT 28.640 167.840 28.960 168.160 ;
        RECT 29.040 167.840 29.360 168.160 ;
        RECT 29.440 167.840 29.760 168.160 ;
        RECT 29.840 167.840 30.160 168.160 ;
        RECT 30.240 167.840 30.560 168.160 ;
        RECT 30.640 167.840 30.960 168.160 ;
        RECT 31.040 167.840 31.360 168.160 ;
        RECT 31.440 167.840 31.760 168.160 ;
        RECT 31.840 167.840 32.160 168.160 ;
        RECT 32.240 167.840 32.560 168.160 ;
        RECT 32.640 167.840 32.960 168.160 ;
        RECT 33.040 167.840 33.360 168.160 ;
        RECT 33.440 167.840 33.760 168.160 ;
        RECT 33.840 167.840 34.160 168.160 ;
        RECT 34.240 167.840 34.560 168.160 ;
        RECT 34.640 167.840 34.960 168.160 ;
        RECT 35.040 167.840 35.360 168.160 ;
        RECT 35.440 167.840 35.760 168.160 ;
        RECT 35.840 167.840 36.160 168.160 ;
        RECT 36.240 167.840 36.560 168.160 ;
        RECT 36.640 167.840 36.960 168.160 ;
        RECT 37.040 167.840 37.360 168.160 ;
        RECT 37.440 167.840 37.760 168.160 ;
        RECT 37.840 167.840 38.160 168.160 ;
        RECT 38.240 167.840 38.560 168.160 ;
        RECT 38.640 167.840 38.960 168.160 ;
        RECT 39.040 167.840 39.360 168.160 ;
        RECT 39.440 167.840 39.760 168.160 ;
        RECT 39.840 167.840 40.160 168.160 ;
        RECT 40.240 167.840 40.560 168.160 ;
        RECT 40.640 167.840 40.960 168.160 ;
        RECT 41.040 167.840 41.360 168.160 ;
        RECT 41.440 167.840 41.760 168.160 ;
        RECT 41.840 167.840 42.160 168.160 ;
        RECT 42.240 167.840 42.560 168.160 ;
        RECT 42.640 167.840 42.960 168.160 ;
        RECT 43.040 167.840 43.360 168.160 ;
        RECT 43.440 167.840 43.760 168.160 ;
        RECT 43.840 167.840 44.160 168.160 ;
        RECT 44.240 167.840 44.560 168.160 ;
        RECT 44.640 167.840 44.960 168.160 ;
        RECT 70.560 167.840 70.880 168.160 ;
        RECT 70.960 167.840 71.280 168.160 ;
        RECT 71.360 167.840 71.680 168.160 ;
        RECT 71.760 167.840 72.080 168.160 ;
        RECT 120.560 167.840 120.880 168.160 ;
        RECT 120.960 167.840 121.280 168.160 ;
        RECT 121.360 167.840 121.680 168.160 ;
        RECT 121.760 167.840 122.080 168.160 ;
        RECT 160.720 167.840 161.040 168.160 ;
        RECT 161.120 167.840 161.440 168.160 ;
        RECT 161.520 167.840 161.840 168.160 ;
        RECT 161.920 167.840 162.240 168.160 ;
        RECT 162.320 167.840 162.640 168.160 ;
        RECT 162.720 167.840 163.040 168.160 ;
        RECT 163.120 167.840 163.440 168.160 ;
        RECT 163.520 167.840 163.840 168.160 ;
        RECT 163.920 167.840 164.240 168.160 ;
        RECT 164.320 167.840 164.640 168.160 ;
        RECT 164.720 167.840 165.040 168.160 ;
        RECT 165.120 167.840 165.440 168.160 ;
        RECT 165.520 167.840 165.840 168.160 ;
        RECT 165.920 167.840 166.240 168.160 ;
        RECT 166.320 167.840 166.640 168.160 ;
        RECT 166.720 167.840 167.040 168.160 ;
        RECT 167.120 167.840 167.440 168.160 ;
        RECT 167.520 167.840 167.840 168.160 ;
        RECT 167.920 167.840 168.240 168.160 ;
        RECT 168.320 167.840 168.640 168.160 ;
        RECT 168.720 167.840 169.040 168.160 ;
        RECT 169.120 167.840 169.440 168.160 ;
        RECT 169.520 167.840 169.840 168.160 ;
        RECT 169.920 167.840 170.240 168.160 ;
        RECT 170.320 167.840 170.640 168.160 ;
        RECT 170.720 167.840 171.040 168.160 ;
        RECT 171.120 167.840 171.440 168.160 ;
        RECT 171.520 167.840 171.840 168.160 ;
        RECT 171.920 167.840 172.240 168.160 ;
        RECT 172.320 167.840 172.640 168.160 ;
        RECT 172.720 167.840 173.040 168.160 ;
        RECT 173.120 167.840 173.440 168.160 ;
        RECT 173.520 167.840 173.840 168.160 ;
        RECT 173.920 167.840 174.240 168.160 ;
        RECT 174.320 167.840 174.640 168.160 ;
        RECT 174.720 167.840 175.040 168.160 ;
        RECT 175.120 167.840 175.440 168.160 ;
        RECT 175.520 167.840 175.840 168.160 ;
        RECT 175.920 167.840 176.240 168.160 ;
        RECT 176.320 167.840 176.640 168.160 ;
        RECT 176.720 167.840 177.040 168.160 ;
        RECT 177.120 167.840 177.440 168.160 ;
        RECT 177.520 167.840 177.840 168.160 ;
        RECT 177.920 167.840 178.240 168.160 ;
        RECT 178.320 167.840 178.640 168.160 ;
        RECT 178.720 167.840 179.040 168.160 ;
        RECT 179.120 167.840 179.440 168.160 ;
        RECT 179.520 167.840 179.840 168.160 ;
        RECT 179.920 167.840 180.240 168.160 ;
        RECT 180.320 167.840 180.640 168.160 ;
        RECT 25.040 167.440 25.360 167.760 ;
        RECT 25.440 167.440 25.760 167.760 ;
        RECT 25.840 167.440 26.160 167.760 ;
        RECT 26.240 167.440 26.560 167.760 ;
        RECT 26.640 167.440 26.960 167.760 ;
        RECT 27.040 167.440 27.360 167.760 ;
        RECT 27.440 167.440 27.760 167.760 ;
        RECT 27.840 167.440 28.160 167.760 ;
        RECT 28.240 167.440 28.560 167.760 ;
        RECT 28.640 167.440 28.960 167.760 ;
        RECT 29.040 167.440 29.360 167.760 ;
        RECT 29.440 167.440 29.760 167.760 ;
        RECT 29.840 167.440 30.160 167.760 ;
        RECT 30.240 167.440 30.560 167.760 ;
        RECT 30.640 167.440 30.960 167.760 ;
        RECT 31.040 167.440 31.360 167.760 ;
        RECT 31.440 167.440 31.760 167.760 ;
        RECT 31.840 167.440 32.160 167.760 ;
        RECT 32.240 167.440 32.560 167.760 ;
        RECT 32.640 167.440 32.960 167.760 ;
        RECT 33.040 167.440 33.360 167.760 ;
        RECT 33.440 167.440 33.760 167.760 ;
        RECT 33.840 167.440 34.160 167.760 ;
        RECT 34.240 167.440 34.560 167.760 ;
        RECT 34.640 167.440 34.960 167.760 ;
        RECT 35.040 167.440 35.360 167.760 ;
        RECT 35.440 167.440 35.760 167.760 ;
        RECT 35.840 167.440 36.160 167.760 ;
        RECT 36.240 167.440 36.560 167.760 ;
        RECT 36.640 167.440 36.960 167.760 ;
        RECT 37.040 167.440 37.360 167.760 ;
        RECT 37.440 167.440 37.760 167.760 ;
        RECT 37.840 167.440 38.160 167.760 ;
        RECT 38.240 167.440 38.560 167.760 ;
        RECT 38.640 167.440 38.960 167.760 ;
        RECT 39.040 167.440 39.360 167.760 ;
        RECT 39.440 167.440 39.760 167.760 ;
        RECT 39.840 167.440 40.160 167.760 ;
        RECT 40.240 167.440 40.560 167.760 ;
        RECT 40.640 167.440 40.960 167.760 ;
        RECT 41.040 167.440 41.360 167.760 ;
        RECT 41.440 167.440 41.760 167.760 ;
        RECT 41.840 167.440 42.160 167.760 ;
        RECT 42.240 167.440 42.560 167.760 ;
        RECT 42.640 167.440 42.960 167.760 ;
        RECT 43.040 167.440 43.360 167.760 ;
        RECT 43.440 167.440 43.760 167.760 ;
        RECT 43.840 167.440 44.160 167.760 ;
        RECT 44.240 167.440 44.560 167.760 ;
        RECT 44.640 167.440 44.960 167.760 ;
        RECT 70.560 167.440 70.880 167.760 ;
        RECT 70.960 167.440 71.280 167.760 ;
        RECT 71.360 167.440 71.680 167.760 ;
        RECT 71.760 167.440 72.080 167.760 ;
        RECT 120.560 167.440 120.880 167.760 ;
        RECT 120.960 167.440 121.280 167.760 ;
        RECT 121.360 167.440 121.680 167.760 ;
        RECT 121.760 167.440 122.080 167.760 ;
        RECT 160.720 167.440 161.040 167.760 ;
        RECT 161.120 167.440 161.440 167.760 ;
        RECT 161.520 167.440 161.840 167.760 ;
        RECT 161.920 167.440 162.240 167.760 ;
        RECT 162.320 167.440 162.640 167.760 ;
        RECT 162.720 167.440 163.040 167.760 ;
        RECT 163.120 167.440 163.440 167.760 ;
        RECT 163.520 167.440 163.840 167.760 ;
        RECT 163.920 167.440 164.240 167.760 ;
        RECT 164.320 167.440 164.640 167.760 ;
        RECT 164.720 167.440 165.040 167.760 ;
        RECT 165.120 167.440 165.440 167.760 ;
        RECT 165.520 167.440 165.840 167.760 ;
        RECT 165.920 167.440 166.240 167.760 ;
        RECT 166.320 167.440 166.640 167.760 ;
        RECT 166.720 167.440 167.040 167.760 ;
        RECT 167.120 167.440 167.440 167.760 ;
        RECT 167.520 167.440 167.840 167.760 ;
        RECT 167.920 167.440 168.240 167.760 ;
        RECT 168.320 167.440 168.640 167.760 ;
        RECT 168.720 167.440 169.040 167.760 ;
        RECT 169.120 167.440 169.440 167.760 ;
        RECT 169.520 167.440 169.840 167.760 ;
        RECT 169.920 167.440 170.240 167.760 ;
        RECT 170.320 167.440 170.640 167.760 ;
        RECT 170.720 167.440 171.040 167.760 ;
        RECT 171.120 167.440 171.440 167.760 ;
        RECT 171.520 167.440 171.840 167.760 ;
        RECT 171.920 167.440 172.240 167.760 ;
        RECT 172.320 167.440 172.640 167.760 ;
        RECT 172.720 167.440 173.040 167.760 ;
        RECT 173.120 167.440 173.440 167.760 ;
        RECT 173.520 167.440 173.840 167.760 ;
        RECT 173.920 167.440 174.240 167.760 ;
        RECT 174.320 167.440 174.640 167.760 ;
        RECT 174.720 167.440 175.040 167.760 ;
        RECT 175.120 167.440 175.440 167.760 ;
        RECT 175.520 167.440 175.840 167.760 ;
        RECT 175.920 167.440 176.240 167.760 ;
        RECT 176.320 167.440 176.640 167.760 ;
        RECT 176.720 167.440 177.040 167.760 ;
        RECT 177.120 167.440 177.440 167.760 ;
        RECT 177.520 167.440 177.840 167.760 ;
        RECT 177.920 167.440 178.240 167.760 ;
        RECT 178.320 167.440 178.640 167.760 ;
        RECT 178.720 167.440 179.040 167.760 ;
        RECT 179.120 167.440 179.440 167.760 ;
        RECT 179.520 167.440 179.840 167.760 ;
        RECT 179.920 167.440 180.240 167.760 ;
        RECT 180.320 167.440 180.640 167.760 ;
        RECT 25.040 167.040 25.360 167.360 ;
        RECT 25.440 167.040 25.760 167.360 ;
        RECT 25.840 167.040 26.160 167.360 ;
        RECT 26.240 167.040 26.560 167.360 ;
        RECT 26.640 167.040 26.960 167.360 ;
        RECT 27.040 167.040 27.360 167.360 ;
        RECT 27.440 167.040 27.760 167.360 ;
        RECT 27.840 167.040 28.160 167.360 ;
        RECT 28.240 167.040 28.560 167.360 ;
        RECT 28.640 167.040 28.960 167.360 ;
        RECT 29.040 167.040 29.360 167.360 ;
        RECT 29.440 167.040 29.760 167.360 ;
        RECT 29.840 167.040 30.160 167.360 ;
        RECT 30.240 167.040 30.560 167.360 ;
        RECT 30.640 167.040 30.960 167.360 ;
        RECT 31.040 167.040 31.360 167.360 ;
        RECT 31.440 167.040 31.760 167.360 ;
        RECT 31.840 167.040 32.160 167.360 ;
        RECT 32.240 167.040 32.560 167.360 ;
        RECT 32.640 167.040 32.960 167.360 ;
        RECT 33.040 167.040 33.360 167.360 ;
        RECT 33.440 167.040 33.760 167.360 ;
        RECT 33.840 167.040 34.160 167.360 ;
        RECT 34.240 167.040 34.560 167.360 ;
        RECT 34.640 167.040 34.960 167.360 ;
        RECT 35.040 167.040 35.360 167.360 ;
        RECT 35.440 167.040 35.760 167.360 ;
        RECT 35.840 167.040 36.160 167.360 ;
        RECT 36.240 167.040 36.560 167.360 ;
        RECT 36.640 167.040 36.960 167.360 ;
        RECT 37.040 167.040 37.360 167.360 ;
        RECT 37.440 167.040 37.760 167.360 ;
        RECT 37.840 167.040 38.160 167.360 ;
        RECT 38.240 167.040 38.560 167.360 ;
        RECT 38.640 167.040 38.960 167.360 ;
        RECT 39.040 167.040 39.360 167.360 ;
        RECT 39.440 167.040 39.760 167.360 ;
        RECT 39.840 167.040 40.160 167.360 ;
        RECT 40.240 167.040 40.560 167.360 ;
        RECT 40.640 167.040 40.960 167.360 ;
        RECT 41.040 167.040 41.360 167.360 ;
        RECT 41.440 167.040 41.760 167.360 ;
        RECT 41.840 167.040 42.160 167.360 ;
        RECT 42.240 167.040 42.560 167.360 ;
        RECT 42.640 167.040 42.960 167.360 ;
        RECT 43.040 167.040 43.360 167.360 ;
        RECT 43.440 167.040 43.760 167.360 ;
        RECT 43.840 167.040 44.160 167.360 ;
        RECT 44.240 167.040 44.560 167.360 ;
        RECT 44.640 167.040 44.960 167.360 ;
        RECT 70.560 167.040 70.880 167.360 ;
        RECT 70.960 167.040 71.280 167.360 ;
        RECT 71.360 167.040 71.680 167.360 ;
        RECT 71.760 167.040 72.080 167.360 ;
        RECT 120.560 167.040 120.880 167.360 ;
        RECT 120.960 167.040 121.280 167.360 ;
        RECT 121.360 167.040 121.680 167.360 ;
        RECT 121.760 167.040 122.080 167.360 ;
        RECT 160.720 167.040 161.040 167.360 ;
        RECT 161.120 167.040 161.440 167.360 ;
        RECT 161.520 167.040 161.840 167.360 ;
        RECT 161.920 167.040 162.240 167.360 ;
        RECT 162.320 167.040 162.640 167.360 ;
        RECT 162.720 167.040 163.040 167.360 ;
        RECT 163.120 167.040 163.440 167.360 ;
        RECT 163.520 167.040 163.840 167.360 ;
        RECT 163.920 167.040 164.240 167.360 ;
        RECT 164.320 167.040 164.640 167.360 ;
        RECT 164.720 167.040 165.040 167.360 ;
        RECT 165.120 167.040 165.440 167.360 ;
        RECT 165.520 167.040 165.840 167.360 ;
        RECT 165.920 167.040 166.240 167.360 ;
        RECT 166.320 167.040 166.640 167.360 ;
        RECT 166.720 167.040 167.040 167.360 ;
        RECT 167.120 167.040 167.440 167.360 ;
        RECT 167.520 167.040 167.840 167.360 ;
        RECT 167.920 167.040 168.240 167.360 ;
        RECT 168.320 167.040 168.640 167.360 ;
        RECT 168.720 167.040 169.040 167.360 ;
        RECT 169.120 167.040 169.440 167.360 ;
        RECT 169.520 167.040 169.840 167.360 ;
        RECT 169.920 167.040 170.240 167.360 ;
        RECT 170.320 167.040 170.640 167.360 ;
        RECT 170.720 167.040 171.040 167.360 ;
        RECT 171.120 167.040 171.440 167.360 ;
        RECT 171.520 167.040 171.840 167.360 ;
        RECT 171.920 167.040 172.240 167.360 ;
        RECT 172.320 167.040 172.640 167.360 ;
        RECT 172.720 167.040 173.040 167.360 ;
        RECT 173.120 167.040 173.440 167.360 ;
        RECT 173.520 167.040 173.840 167.360 ;
        RECT 173.920 167.040 174.240 167.360 ;
        RECT 174.320 167.040 174.640 167.360 ;
        RECT 174.720 167.040 175.040 167.360 ;
        RECT 175.120 167.040 175.440 167.360 ;
        RECT 175.520 167.040 175.840 167.360 ;
        RECT 175.920 167.040 176.240 167.360 ;
        RECT 176.320 167.040 176.640 167.360 ;
        RECT 176.720 167.040 177.040 167.360 ;
        RECT 177.120 167.040 177.440 167.360 ;
        RECT 177.520 167.040 177.840 167.360 ;
        RECT 177.920 167.040 178.240 167.360 ;
        RECT 178.320 167.040 178.640 167.360 ;
        RECT 178.720 167.040 179.040 167.360 ;
        RECT 179.120 167.040 179.440 167.360 ;
        RECT 179.520 167.040 179.840 167.360 ;
        RECT 179.920 167.040 180.240 167.360 ;
        RECT 180.320 167.040 180.640 167.360 ;
        RECT 25.040 166.640 25.360 166.960 ;
        RECT 25.440 166.640 25.760 166.960 ;
        RECT 25.840 166.640 26.160 166.960 ;
        RECT 26.240 166.640 26.560 166.960 ;
        RECT 26.640 166.640 26.960 166.960 ;
        RECT 27.040 166.640 27.360 166.960 ;
        RECT 27.440 166.640 27.760 166.960 ;
        RECT 27.840 166.640 28.160 166.960 ;
        RECT 28.240 166.640 28.560 166.960 ;
        RECT 28.640 166.640 28.960 166.960 ;
        RECT 29.040 166.640 29.360 166.960 ;
        RECT 29.440 166.640 29.760 166.960 ;
        RECT 29.840 166.640 30.160 166.960 ;
        RECT 30.240 166.640 30.560 166.960 ;
        RECT 30.640 166.640 30.960 166.960 ;
        RECT 31.040 166.640 31.360 166.960 ;
        RECT 31.440 166.640 31.760 166.960 ;
        RECT 31.840 166.640 32.160 166.960 ;
        RECT 32.240 166.640 32.560 166.960 ;
        RECT 32.640 166.640 32.960 166.960 ;
        RECT 33.040 166.640 33.360 166.960 ;
        RECT 33.440 166.640 33.760 166.960 ;
        RECT 33.840 166.640 34.160 166.960 ;
        RECT 34.240 166.640 34.560 166.960 ;
        RECT 34.640 166.640 34.960 166.960 ;
        RECT 35.040 166.640 35.360 166.960 ;
        RECT 35.440 166.640 35.760 166.960 ;
        RECT 35.840 166.640 36.160 166.960 ;
        RECT 36.240 166.640 36.560 166.960 ;
        RECT 36.640 166.640 36.960 166.960 ;
        RECT 37.040 166.640 37.360 166.960 ;
        RECT 37.440 166.640 37.760 166.960 ;
        RECT 37.840 166.640 38.160 166.960 ;
        RECT 38.240 166.640 38.560 166.960 ;
        RECT 38.640 166.640 38.960 166.960 ;
        RECT 39.040 166.640 39.360 166.960 ;
        RECT 39.440 166.640 39.760 166.960 ;
        RECT 39.840 166.640 40.160 166.960 ;
        RECT 40.240 166.640 40.560 166.960 ;
        RECT 40.640 166.640 40.960 166.960 ;
        RECT 41.040 166.640 41.360 166.960 ;
        RECT 41.440 166.640 41.760 166.960 ;
        RECT 41.840 166.640 42.160 166.960 ;
        RECT 42.240 166.640 42.560 166.960 ;
        RECT 42.640 166.640 42.960 166.960 ;
        RECT 43.040 166.640 43.360 166.960 ;
        RECT 43.440 166.640 43.760 166.960 ;
        RECT 43.840 166.640 44.160 166.960 ;
        RECT 44.240 166.640 44.560 166.960 ;
        RECT 44.640 166.640 44.960 166.960 ;
        RECT 70.560 166.640 70.880 166.960 ;
        RECT 70.960 166.640 71.280 166.960 ;
        RECT 71.360 166.640 71.680 166.960 ;
        RECT 71.760 166.640 72.080 166.960 ;
        RECT 120.560 166.640 120.880 166.960 ;
        RECT 120.960 166.640 121.280 166.960 ;
        RECT 121.360 166.640 121.680 166.960 ;
        RECT 121.760 166.640 122.080 166.960 ;
        RECT 160.720 166.640 161.040 166.960 ;
        RECT 161.120 166.640 161.440 166.960 ;
        RECT 161.520 166.640 161.840 166.960 ;
        RECT 161.920 166.640 162.240 166.960 ;
        RECT 162.320 166.640 162.640 166.960 ;
        RECT 162.720 166.640 163.040 166.960 ;
        RECT 163.120 166.640 163.440 166.960 ;
        RECT 163.520 166.640 163.840 166.960 ;
        RECT 163.920 166.640 164.240 166.960 ;
        RECT 164.320 166.640 164.640 166.960 ;
        RECT 164.720 166.640 165.040 166.960 ;
        RECT 165.120 166.640 165.440 166.960 ;
        RECT 165.520 166.640 165.840 166.960 ;
        RECT 165.920 166.640 166.240 166.960 ;
        RECT 166.320 166.640 166.640 166.960 ;
        RECT 166.720 166.640 167.040 166.960 ;
        RECT 167.120 166.640 167.440 166.960 ;
        RECT 167.520 166.640 167.840 166.960 ;
        RECT 167.920 166.640 168.240 166.960 ;
        RECT 168.320 166.640 168.640 166.960 ;
        RECT 168.720 166.640 169.040 166.960 ;
        RECT 169.120 166.640 169.440 166.960 ;
        RECT 169.520 166.640 169.840 166.960 ;
        RECT 169.920 166.640 170.240 166.960 ;
        RECT 170.320 166.640 170.640 166.960 ;
        RECT 170.720 166.640 171.040 166.960 ;
        RECT 171.120 166.640 171.440 166.960 ;
        RECT 171.520 166.640 171.840 166.960 ;
        RECT 171.920 166.640 172.240 166.960 ;
        RECT 172.320 166.640 172.640 166.960 ;
        RECT 172.720 166.640 173.040 166.960 ;
        RECT 173.120 166.640 173.440 166.960 ;
        RECT 173.520 166.640 173.840 166.960 ;
        RECT 173.920 166.640 174.240 166.960 ;
        RECT 174.320 166.640 174.640 166.960 ;
        RECT 174.720 166.640 175.040 166.960 ;
        RECT 175.120 166.640 175.440 166.960 ;
        RECT 175.520 166.640 175.840 166.960 ;
        RECT 175.920 166.640 176.240 166.960 ;
        RECT 176.320 166.640 176.640 166.960 ;
        RECT 176.720 166.640 177.040 166.960 ;
        RECT 177.120 166.640 177.440 166.960 ;
        RECT 177.520 166.640 177.840 166.960 ;
        RECT 177.920 166.640 178.240 166.960 ;
        RECT 178.320 166.640 178.640 166.960 ;
        RECT 178.720 166.640 179.040 166.960 ;
        RECT 179.120 166.640 179.440 166.960 ;
        RECT 179.520 166.640 179.840 166.960 ;
        RECT 179.920 166.640 180.240 166.960 ;
        RECT 180.320 166.640 180.640 166.960 ;
        RECT 25.040 166.240 25.360 166.560 ;
        RECT 25.440 166.240 25.760 166.560 ;
        RECT 25.840 166.240 26.160 166.560 ;
        RECT 26.240 166.240 26.560 166.560 ;
        RECT 26.640 166.240 26.960 166.560 ;
        RECT 27.040 166.240 27.360 166.560 ;
        RECT 27.440 166.240 27.760 166.560 ;
        RECT 27.840 166.240 28.160 166.560 ;
        RECT 28.240 166.240 28.560 166.560 ;
        RECT 28.640 166.240 28.960 166.560 ;
        RECT 29.040 166.240 29.360 166.560 ;
        RECT 29.440 166.240 29.760 166.560 ;
        RECT 29.840 166.240 30.160 166.560 ;
        RECT 30.240 166.240 30.560 166.560 ;
        RECT 30.640 166.240 30.960 166.560 ;
        RECT 31.040 166.240 31.360 166.560 ;
        RECT 31.440 166.240 31.760 166.560 ;
        RECT 31.840 166.240 32.160 166.560 ;
        RECT 32.240 166.240 32.560 166.560 ;
        RECT 32.640 166.240 32.960 166.560 ;
        RECT 33.040 166.240 33.360 166.560 ;
        RECT 33.440 166.240 33.760 166.560 ;
        RECT 33.840 166.240 34.160 166.560 ;
        RECT 34.240 166.240 34.560 166.560 ;
        RECT 34.640 166.240 34.960 166.560 ;
        RECT 35.040 166.240 35.360 166.560 ;
        RECT 35.440 166.240 35.760 166.560 ;
        RECT 35.840 166.240 36.160 166.560 ;
        RECT 36.240 166.240 36.560 166.560 ;
        RECT 36.640 166.240 36.960 166.560 ;
        RECT 37.040 166.240 37.360 166.560 ;
        RECT 37.440 166.240 37.760 166.560 ;
        RECT 37.840 166.240 38.160 166.560 ;
        RECT 38.240 166.240 38.560 166.560 ;
        RECT 38.640 166.240 38.960 166.560 ;
        RECT 39.040 166.240 39.360 166.560 ;
        RECT 39.440 166.240 39.760 166.560 ;
        RECT 39.840 166.240 40.160 166.560 ;
        RECT 40.240 166.240 40.560 166.560 ;
        RECT 40.640 166.240 40.960 166.560 ;
        RECT 41.040 166.240 41.360 166.560 ;
        RECT 41.440 166.240 41.760 166.560 ;
        RECT 41.840 166.240 42.160 166.560 ;
        RECT 42.240 166.240 42.560 166.560 ;
        RECT 42.640 166.240 42.960 166.560 ;
        RECT 43.040 166.240 43.360 166.560 ;
        RECT 43.440 166.240 43.760 166.560 ;
        RECT 43.840 166.240 44.160 166.560 ;
        RECT 44.240 166.240 44.560 166.560 ;
        RECT 44.640 166.240 44.960 166.560 ;
        RECT 70.560 166.240 70.880 166.560 ;
        RECT 70.960 166.240 71.280 166.560 ;
        RECT 71.360 166.240 71.680 166.560 ;
        RECT 71.760 166.240 72.080 166.560 ;
        RECT 120.560 166.240 120.880 166.560 ;
        RECT 120.960 166.240 121.280 166.560 ;
        RECT 121.360 166.240 121.680 166.560 ;
        RECT 121.760 166.240 122.080 166.560 ;
        RECT 160.720 166.240 161.040 166.560 ;
        RECT 161.120 166.240 161.440 166.560 ;
        RECT 161.520 166.240 161.840 166.560 ;
        RECT 161.920 166.240 162.240 166.560 ;
        RECT 162.320 166.240 162.640 166.560 ;
        RECT 162.720 166.240 163.040 166.560 ;
        RECT 163.120 166.240 163.440 166.560 ;
        RECT 163.520 166.240 163.840 166.560 ;
        RECT 163.920 166.240 164.240 166.560 ;
        RECT 164.320 166.240 164.640 166.560 ;
        RECT 164.720 166.240 165.040 166.560 ;
        RECT 165.120 166.240 165.440 166.560 ;
        RECT 165.520 166.240 165.840 166.560 ;
        RECT 165.920 166.240 166.240 166.560 ;
        RECT 166.320 166.240 166.640 166.560 ;
        RECT 166.720 166.240 167.040 166.560 ;
        RECT 167.120 166.240 167.440 166.560 ;
        RECT 167.520 166.240 167.840 166.560 ;
        RECT 167.920 166.240 168.240 166.560 ;
        RECT 168.320 166.240 168.640 166.560 ;
        RECT 168.720 166.240 169.040 166.560 ;
        RECT 169.120 166.240 169.440 166.560 ;
        RECT 169.520 166.240 169.840 166.560 ;
        RECT 169.920 166.240 170.240 166.560 ;
        RECT 170.320 166.240 170.640 166.560 ;
        RECT 170.720 166.240 171.040 166.560 ;
        RECT 171.120 166.240 171.440 166.560 ;
        RECT 171.520 166.240 171.840 166.560 ;
        RECT 171.920 166.240 172.240 166.560 ;
        RECT 172.320 166.240 172.640 166.560 ;
        RECT 172.720 166.240 173.040 166.560 ;
        RECT 173.120 166.240 173.440 166.560 ;
        RECT 173.520 166.240 173.840 166.560 ;
        RECT 173.920 166.240 174.240 166.560 ;
        RECT 174.320 166.240 174.640 166.560 ;
        RECT 174.720 166.240 175.040 166.560 ;
        RECT 175.120 166.240 175.440 166.560 ;
        RECT 175.520 166.240 175.840 166.560 ;
        RECT 175.920 166.240 176.240 166.560 ;
        RECT 176.320 166.240 176.640 166.560 ;
        RECT 176.720 166.240 177.040 166.560 ;
        RECT 177.120 166.240 177.440 166.560 ;
        RECT 177.520 166.240 177.840 166.560 ;
        RECT 177.920 166.240 178.240 166.560 ;
        RECT 178.320 166.240 178.640 166.560 ;
        RECT 178.720 166.240 179.040 166.560 ;
        RECT 179.120 166.240 179.440 166.560 ;
        RECT 179.520 166.240 179.840 166.560 ;
        RECT 179.920 166.240 180.240 166.560 ;
        RECT 180.320 166.240 180.640 166.560 ;
        RECT 25.040 165.840 25.360 166.160 ;
        RECT 25.440 165.840 25.760 166.160 ;
        RECT 25.840 165.840 26.160 166.160 ;
        RECT 26.240 165.840 26.560 166.160 ;
        RECT 26.640 165.840 26.960 166.160 ;
        RECT 27.040 165.840 27.360 166.160 ;
        RECT 27.440 165.840 27.760 166.160 ;
        RECT 27.840 165.840 28.160 166.160 ;
        RECT 28.240 165.840 28.560 166.160 ;
        RECT 28.640 165.840 28.960 166.160 ;
        RECT 29.040 165.840 29.360 166.160 ;
        RECT 29.440 165.840 29.760 166.160 ;
        RECT 29.840 165.840 30.160 166.160 ;
        RECT 30.240 165.840 30.560 166.160 ;
        RECT 30.640 165.840 30.960 166.160 ;
        RECT 31.040 165.840 31.360 166.160 ;
        RECT 31.440 165.840 31.760 166.160 ;
        RECT 31.840 165.840 32.160 166.160 ;
        RECT 32.240 165.840 32.560 166.160 ;
        RECT 32.640 165.840 32.960 166.160 ;
        RECT 33.040 165.840 33.360 166.160 ;
        RECT 33.440 165.840 33.760 166.160 ;
        RECT 33.840 165.840 34.160 166.160 ;
        RECT 34.240 165.840 34.560 166.160 ;
        RECT 34.640 165.840 34.960 166.160 ;
        RECT 35.040 165.840 35.360 166.160 ;
        RECT 35.440 165.840 35.760 166.160 ;
        RECT 35.840 165.840 36.160 166.160 ;
        RECT 36.240 165.840 36.560 166.160 ;
        RECT 36.640 165.840 36.960 166.160 ;
        RECT 37.040 165.840 37.360 166.160 ;
        RECT 37.440 165.840 37.760 166.160 ;
        RECT 37.840 165.840 38.160 166.160 ;
        RECT 38.240 165.840 38.560 166.160 ;
        RECT 38.640 165.840 38.960 166.160 ;
        RECT 39.040 165.840 39.360 166.160 ;
        RECT 39.440 165.840 39.760 166.160 ;
        RECT 39.840 165.840 40.160 166.160 ;
        RECT 40.240 165.840 40.560 166.160 ;
        RECT 40.640 165.840 40.960 166.160 ;
        RECT 41.040 165.840 41.360 166.160 ;
        RECT 41.440 165.840 41.760 166.160 ;
        RECT 41.840 165.840 42.160 166.160 ;
        RECT 42.240 165.840 42.560 166.160 ;
        RECT 42.640 165.840 42.960 166.160 ;
        RECT 43.040 165.840 43.360 166.160 ;
        RECT 43.440 165.840 43.760 166.160 ;
        RECT 43.840 165.840 44.160 166.160 ;
        RECT 44.240 165.840 44.560 166.160 ;
        RECT 44.640 165.840 44.960 166.160 ;
        RECT 70.560 165.840 70.880 166.160 ;
        RECT 70.960 165.840 71.280 166.160 ;
        RECT 71.360 165.840 71.680 166.160 ;
        RECT 71.760 165.840 72.080 166.160 ;
        RECT 120.560 165.840 120.880 166.160 ;
        RECT 120.960 165.840 121.280 166.160 ;
        RECT 121.360 165.840 121.680 166.160 ;
        RECT 121.760 165.840 122.080 166.160 ;
        RECT 160.720 165.840 161.040 166.160 ;
        RECT 161.120 165.840 161.440 166.160 ;
        RECT 161.520 165.840 161.840 166.160 ;
        RECT 161.920 165.840 162.240 166.160 ;
        RECT 162.320 165.840 162.640 166.160 ;
        RECT 162.720 165.840 163.040 166.160 ;
        RECT 163.120 165.840 163.440 166.160 ;
        RECT 163.520 165.840 163.840 166.160 ;
        RECT 163.920 165.840 164.240 166.160 ;
        RECT 164.320 165.840 164.640 166.160 ;
        RECT 164.720 165.840 165.040 166.160 ;
        RECT 165.120 165.840 165.440 166.160 ;
        RECT 165.520 165.840 165.840 166.160 ;
        RECT 165.920 165.840 166.240 166.160 ;
        RECT 166.320 165.840 166.640 166.160 ;
        RECT 166.720 165.840 167.040 166.160 ;
        RECT 167.120 165.840 167.440 166.160 ;
        RECT 167.520 165.840 167.840 166.160 ;
        RECT 167.920 165.840 168.240 166.160 ;
        RECT 168.320 165.840 168.640 166.160 ;
        RECT 168.720 165.840 169.040 166.160 ;
        RECT 169.120 165.840 169.440 166.160 ;
        RECT 169.520 165.840 169.840 166.160 ;
        RECT 169.920 165.840 170.240 166.160 ;
        RECT 170.320 165.840 170.640 166.160 ;
        RECT 170.720 165.840 171.040 166.160 ;
        RECT 171.120 165.840 171.440 166.160 ;
        RECT 171.520 165.840 171.840 166.160 ;
        RECT 171.920 165.840 172.240 166.160 ;
        RECT 172.320 165.840 172.640 166.160 ;
        RECT 172.720 165.840 173.040 166.160 ;
        RECT 173.120 165.840 173.440 166.160 ;
        RECT 173.520 165.840 173.840 166.160 ;
        RECT 173.920 165.840 174.240 166.160 ;
        RECT 174.320 165.840 174.640 166.160 ;
        RECT 174.720 165.840 175.040 166.160 ;
        RECT 175.120 165.840 175.440 166.160 ;
        RECT 175.520 165.840 175.840 166.160 ;
        RECT 175.920 165.840 176.240 166.160 ;
        RECT 176.320 165.840 176.640 166.160 ;
        RECT 176.720 165.840 177.040 166.160 ;
        RECT 177.120 165.840 177.440 166.160 ;
        RECT 177.520 165.840 177.840 166.160 ;
        RECT 177.920 165.840 178.240 166.160 ;
        RECT 178.320 165.840 178.640 166.160 ;
        RECT 178.720 165.840 179.040 166.160 ;
        RECT 179.120 165.840 179.440 166.160 ;
        RECT 179.520 165.840 179.840 166.160 ;
        RECT 179.920 165.840 180.240 166.160 ;
        RECT 180.320 165.840 180.640 166.160 ;
        RECT 25.040 165.440 25.360 165.760 ;
        RECT 25.440 165.440 25.760 165.760 ;
        RECT 25.840 165.440 26.160 165.760 ;
        RECT 26.240 165.440 26.560 165.760 ;
        RECT 26.640 165.440 26.960 165.760 ;
        RECT 27.040 165.440 27.360 165.760 ;
        RECT 27.440 165.440 27.760 165.760 ;
        RECT 27.840 165.440 28.160 165.760 ;
        RECT 28.240 165.440 28.560 165.760 ;
        RECT 28.640 165.440 28.960 165.760 ;
        RECT 29.040 165.440 29.360 165.760 ;
        RECT 29.440 165.440 29.760 165.760 ;
        RECT 29.840 165.440 30.160 165.760 ;
        RECT 30.240 165.440 30.560 165.760 ;
        RECT 30.640 165.440 30.960 165.760 ;
        RECT 31.040 165.440 31.360 165.760 ;
        RECT 31.440 165.440 31.760 165.760 ;
        RECT 31.840 165.440 32.160 165.760 ;
        RECT 32.240 165.440 32.560 165.760 ;
        RECT 32.640 165.440 32.960 165.760 ;
        RECT 33.040 165.440 33.360 165.760 ;
        RECT 33.440 165.440 33.760 165.760 ;
        RECT 33.840 165.440 34.160 165.760 ;
        RECT 34.240 165.440 34.560 165.760 ;
        RECT 34.640 165.440 34.960 165.760 ;
        RECT 35.040 165.440 35.360 165.760 ;
        RECT 35.440 165.440 35.760 165.760 ;
        RECT 35.840 165.440 36.160 165.760 ;
        RECT 36.240 165.440 36.560 165.760 ;
        RECT 36.640 165.440 36.960 165.760 ;
        RECT 37.040 165.440 37.360 165.760 ;
        RECT 37.440 165.440 37.760 165.760 ;
        RECT 37.840 165.440 38.160 165.760 ;
        RECT 38.240 165.440 38.560 165.760 ;
        RECT 38.640 165.440 38.960 165.760 ;
        RECT 39.040 165.440 39.360 165.760 ;
        RECT 39.440 165.440 39.760 165.760 ;
        RECT 39.840 165.440 40.160 165.760 ;
        RECT 40.240 165.440 40.560 165.760 ;
        RECT 40.640 165.440 40.960 165.760 ;
        RECT 41.040 165.440 41.360 165.760 ;
        RECT 41.440 165.440 41.760 165.760 ;
        RECT 41.840 165.440 42.160 165.760 ;
        RECT 42.240 165.440 42.560 165.760 ;
        RECT 42.640 165.440 42.960 165.760 ;
        RECT 43.040 165.440 43.360 165.760 ;
        RECT 43.440 165.440 43.760 165.760 ;
        RECT 43.840 165.440 44.160 165.760 ;
        RECT 44.240 165.440 44.560 165.760 ;
        RECT 44.640 165.440 44.960 165.760 ;
        RECT 70.560 165.440 70.880 165.760 ;
        RECT 70.960 165.440 71.280 165.760 ;
        RECT 71.360 165.440 71.680 165.760 ;
        RECT 71.760 165.440 72.080 165.760 ;
        RECT 120.560 165.440 120.880 165.760 ;
        RECT 120.960 165.440 121.280 165.760 ;
        RECT 121.360 165.440 121.680 165.760 ;
        RECT 121.760 165.440 122.080 165.760 ;
        RECT 160.720 165.440 161.040 165.760 ;
        RECT 161.120 165.440 161.440 165.760 ;
        RECT 161.520 165.440 161.840 165.760 ;
        RECT 161.920 165.440 162.240 165.760 ;
        RECT 162.320 165.440 162.640 165.760 ;
        RECT 162.720 165.440 163.040 165.760 ;
        RECT 163.120 165.440 163.440 165.760 ;
        RECT 163.520 165.440 163.840 165.760 ;
        RECT 163.920 165.440 164.240 165.760 ;
        RECT 164.320 165.440 164.640 165.760 ;
        RECT 164.720 165.440 165.040 165.760 ;
        RECT 165.120 165.440 165.440 165.760 ;
        RECT 165.520 165.440 165.840 165.760 ;
        RECT 165.920 165.440 166.240 165.760 ;
        RECT 166.320 165.440 166.640 165.760 ;
        RECT 166.720 165.440 167.040 165.760 ;
        RECT 167.120 165.440 167.440 165.760 ;
        RECT 167.520 165.440 167.840 165.760 ;
        RECT 167.920 165.440 168.240 165.760 ;
        RECT 168.320 165.440 168.640 165.760 ;
        RECT 168.720 165.440 169.040 165.760 ;
        RECT 169.120 165.440 169.440 165.760 ;
        RECT 169.520 165.440 169.840 165.760 ;
        RECT 169.920 165.440 170.240 165.760 ;
        RECT 170.320 165.440 170.640 165.760 ;
        RECT 170.720 165.440 171.040 165.760 ;
        RECT 171.120 165.440 171.440 165.760 ;
        RECT 171.520 165.440 171.840 165.760 ;
        RECT 171.920 165.440 172.240 165.760 ;
        RECT 172.320 165.440 172.640 165.760 ;
        RECT 172.720 165.440 173.040 165.760 ;
        RECT 173.120 165.440 173.440 165.760 ;
        RECT 173.520 165.440 173.840 165.760 ;
        RECT 173.920 165.440 174.240 165.760 ;
        RECT 174.320 165.440 174.640 165.760 ;
        RECT 174.720 165.440 175.040 165.760 ;
        RECT 175.120 165.440 175.440 165.760 ;
        RECT 175.520 165.440 175.840 165.760 ;
        RECT 175.920 165.440 176.240 165.760 ;
        RECT 176.320 165.440 176.640 165.760 ;
        RECT 176.720 165.440 177.040 165.760 ;
        RECT 177.120 165.440 177.440 165.760 ;
        RECT 177.520 165.440 177.840 165.760 ;
        RECT 177.920 165.440 178.240 165.760 ;
        RECT 178.320 165.440 178.640 165.760 ;
        RECT 178.720 165.440 179.040 165.760 ;
        RECT 179.120 165.440 179.440 165.760 ;
        RECT 179.520 165.440 179.840 165.760 ;
        RECT 179.920 165.440 180.240 165.760 ;
        RECT 180.320 165.440 180.640 165.760 ;
        RECT 25.040 165.040 25.360 165.360 ;
        RECT 25.440 165.040 25.760 165.360 ;
        RECT 25.840 165.040 26.160 165.360 ;
        RECT 26.240 165.040 26.560 165.360 ;
        RECT 26.640 165.040 26.960 165.360 ;
        RECT 27.040 165.040 27.360 165.360 ;
        RECT 27.440 165.040 27.760 165.360 ;
        RECT 27.840 165.040 28.160 165.360 ;
        RECT 28.240 165.040 28.560 165.360 ;
        RECT 28.640 165.040 28.960 165.360 ;
        RECT 29.040 165.040 29.360 165.360 ;
        RECT 29.440 165.040 29.760 165.360 ;
        RECT 29.840 165.040 30.160 165.360 ;
        RECT 30.240 165.040 30.560 165.360 ;
        RECT 30.640 165.040 30.960 165.360 ;
        RECT 31.040 165.040 31.360 165.360 ;
        RECT 31.440 165.040 31.760 165.360 ;
        RECT 31.840 165.040 32.160 165.360 ;
        RECT 32.240 165.040 32.560 165.360 ;
        RECT 32.640 165.040 32.960 165.360 ;
        RECT 33.040 165.040 33.360 165.360 ;
        RECT 33.440 165.040 33.760 165.360 ;
        RECT 33.840 165.040 34.160 165.360 ;
        RECT 34.240 165.040 34.560 165.360 ;
        RECT 34.640 165.040 34.960 165.360 ;
        RECT 35.040 165.040 35.360 165.360 ;
        RECT 35.440 165.040 35.760 165.360 ;
        RECT 35.840 165.040 36.160 165.360 ;
        RECT 36.240 165.040 36.560 165.360 ;
        RECT 36.640 165.040 36.960 165.360 ;
        RECT 37.040 165.040 37.360 165.360 ;
        RECT 37.440 165.040 37.760 165.360 ;
        RECT 37.840 165.040 38.160 165.360 ;
        RECT 38.240 165.040 38.560 165.360 ;
        RECT 38.640 165.040 38.960 165.360 ;
        RECT 39.040 165.040 39.360 165.360 ;
        RECT 39.440 165.040 39.760 165.360 ;
        RECT 39.840 165.040 40.160 165.360 ;
        RECT 40.240 165.040 40.560 165.360 ;
        RECT 40.640 165.040 40.960 165.360 ;
        RECT 41.040 165.040 41.360 165.360 ;
        RECT 41.440 165.040 41.760 165.360 ;
        RECT 41.840 165.040 42.160 165.360 ;
        RECT 42.240 165.040 42.560 165.360 ;
        RECT 42.640 165.040 42.960 165.360 ;
        RECT 43.040 165.040 43.360 165.360 ;
        RECT 43.440 165.040 43.760 165.360 ;
        RECT 43.840 165.040 44.160 165.360 ;
        RECT 44.240 165.040 44.560 165.360 ;
        RECT 44.640 165.040 44.960 165.360 ;
        RECT 70.560 165.040 70.880 165.360 ;
        RECT 70.960 165.040 71.280 165.360 ;
        RECT 71.360 165.040 71.680 165.360 ;
        RECT 71.760 165.040 72.080 165.360 ;
        RECT 120.560 165.040 120.880 165.360 ;
        RECT 120.960 165.040 121.280 165.360 ;
        RECT 121.360 165.040 121.680 165.360 ;
        RECT 121.760 165.040 122.080 165.360 ;
        RECT 160.720 165.040 161.040 165.360 ;
        RECT 161.120 165.040 161.440 165.360 ;
        RECT 161.520 165.040 161.840 165.360 ;
        RECT 161.920 165.040 162.240 165.360 ;
        RECT 162.320 165.040 162.640 165.360 ;
        RECT 162.720 165.040 163.040 165.360 ;
        RECT 163.120 165.040 163.440 165.360 ;
        RECT 163.520 165.040 163.840 165.360 ;
        RECT 163.920 165.040 164.240 165.360 ;
        RECT 164.320 165.040 164.640 165.360 ;
        RECT 164.720 165.040 165.040 165.360 ;
        RECT 165.120 165.040 165.440 165.360 ;
        RECT 165.520 165.040 165.840 165.360 ;
        RECT 165.920 165.040 166.240 165.360 ;
        RECT 166.320 165.040 166.640 165.360 ;
        RECT 166.720 165.040 167.040 165.360 ;
        RECT 167.120 165.040 167.440 165.360 ;
        RECT 167.520 165.040 167.840 165.360 ;
        RECT 167.920 165.040 168.240 165.360 ;
        RECT 168.320 165.040 168.640 165.360 ;
        RECT 168.720 165.040 169.040 165.360 ;
        RECT 169.120 165.040 169.440 165.360 ;
        RECT 169.520 165.040 169.840 165.360 ;
        RECT 169.920 165.040 170.240 165.360 ;
        RECT 170.320 165.040 170.640 165.360 ;
        RECT 170.720 165.040 171.040 165.360 ;
        RECT 171.120 165.040 171.440 165.360 ;
        RECT 171.520 165.040 171.840 165.360 ;
        RECT 171.920 165.040 172.240 165.360 ;
        RECT 172.320 165.040 172.640 165.360 ;
        RECT 172.720 165.040 173.040 165.360 ;
        RECT 173.120 165.040 173.440 165.360 ;
        RECT 173.520 165.040 173.840 165.360 ;
        RECT 173.920 165.040 174.240 165.360 ;
        RECT 174.320 165.040 174.640 165.360 ;
        RECT 174.720 165.040 175.040 165.360 ;
        RECT 175.120 165.040 175.440 165.360 ;
        RECT 175.520 165.040 175.840 165.360 ;
        RECT 175.920 165.040 176.240 165.360 ;
        RECT 176.320 165.040 176.640 165.360 ;
        RECT 176.720 165.040 177.040 165.360 ;
        RECT 177.120 165.040 177.440 165.360 ;
        RECT 177.520 165.040 177.840 165.360 ;
        RECT 177.920 165.040 178.240 165.360 ;
        RECT 178.320 165.040 178.640 165.360 ;
        RECT 178.720 165.040 179.040 165.360 ;
        RECT 179.120 165.040 179.440 165.360 ;
        RECT 179.520 165.040 179.840 165.360 ;
        RECT 179.920 165.040 180.240 165.360 ;
        RECT 180.320 165.040 180.640 165.360 ;
        RECT 25.040 164.640 25.360 164.960 ;
        RECT 25.440 164.640 25.760 164.960 ;
        RECT 25.840 164.640 26.160 164.960 ;
        RECT 26.240 164.640 26.560 164.960 ;
        RECT 26.640 164.640 26.960 164.960 ;
        RECT 27.040 164.640 27.360 164.960 ;
        RECT 27.440 164.640 27.760 164.960 ;
        RECT 27.840 164.640 28.160 164.960 ;
        RECT 28.240 164.640 28.560 164.960 ;
        RECT 28.640 164.640 28.960 164.960 ;
        RECT 29.040 164.640 29.360 164.960 ;
        RECT 29.440 164.640 29.760 164.960 ;
        RECT 29.840 164.640 30.160 164.960 ;
        RECT 30.240 164.640 30.560 164.960 ;
        RECT 30.640 164.640 30.960 164.960 ;
        RECT 31.040 164.640 31.360 164.960 ;
        RECT 31.440 164.640 31.760 164.960 ;
        RECT 31.840 164.640 32.160 164.960 ;
        RECT 32.240 164.640 32.560 164.960 ;
        RECT 32.640 164.640 32.960 164.960 ;
        RECT 33.040 164.640 33.360 164.960 ;
        RECT 33.440 164.640 33.760 164.960 ;
        RECT 33.840 164.640 34.160 164.960 ;
        RECT 34.240 164.640 34.560 164.960 ;
        RECT 34.640 164.640 34.960 164.960 ;
        RECT 35.040 164.640 35.360 164.960 ;
        RECT 35.440 164.640 35.760 164.960 ;
        RECT 35.840 164.640 36.160 164.960 ;
        RECT 36.240 164.640 36.560 164.960 ;
        RECT 36.640 164.640 36.960 164.960 ;
        RECT 37.040 164.640 37.360 164.960 ;
        RECT 37.440 164.640 37.760 164.960 ;
        RECT 37.840 164.640 38.160 164.960 ;
        RECT 38.240 164.640 38.560 164.960 ;
        RECT 38.640 164.640 38.960 164.960 ;
        RECT 39.040 164.640 39.360 164.960 ;
        RECT 39.440 164.640 39.760 164.960 ;
        RECT 39.840 164.640 40.160 164.960 ;
        RECT 40.240 164.640 40.560 164.960 ;
        RECT 40.640 164.640 40.960 164.960 ;
        RECT 41.040 164.640 41.360 164.960 ;
        RECT 41.440 164.640 41.760 164.960 ;
        RECT 41.840 164.640 42.160 164.960 ;
        RECT 42.240 164.640 42.560 164.960 ;
        RECT 42.640 164.640 42.960 164.960 ;
        RECT 43.040 164.640 43.360 164.960 ;
        RECT 43.440 164.640 43.760 164.960 ;
        RECT 43.840 164.640 44.160 164.960 ;
        RECT 44.240 164.640 44.560 164.960 ;
        RECT 44.640 164.640 44.960 164.960 ;
        RECT 70.560 164.640 70.880 164.960 ;
        RECT 70.960 164.640 71.280 164.960 ;
        RECT 71.360 164.640 71.680 164.960 ;
        RECT 71.760 164.640 72.080 164.960 ;
        RECT 120.560 164.640 120.880 164.960 ;
        RECT 120.960 164.640 121.280 164.960 ;
        RECT 121.360 164.640 121.680 164.960 ;
        RECT 121.760 164.640 122.080 164.960 ;
        RECT 160.720 164.640 161.040 164.960 ;
        RECT 161.120 164.640 161.440 164.960 ;
        RECT 161.520 164.640 161.840 164.960 ;
        RECT 161.920 164.640 162.240 164.960 ;
        RECT 162.320 164.640 162.640 164.960 ;
        RECT 162.720 164.640 163.040 164.960 ;
        RECT 163.120 164.640 163.440 164.960 ;
        RECT 163.520 164.640 163.840 164.960 ;
        RECT 163.920 164.640 164.240 164.960 ;
        RECT 164.320 164.640 164.640 164.960 ;
        RECT 164.720 164.640 165.040 164.960 ;
        RECT 165.120 164.640 165.440 164.960 ;
        RECT 165.520 164.640 165.840 164.960 ;
        RECT 165.920 164.640 166.240 164.960 ;
        RECT 166.320 164.640 166.640 164.960 ;
        RECT 166.720 164.640 167.040 164.960 ;
        RECT 167.120 164.640 167.440 164.960 ;
        RECT 167.520 164.640 167.840 164.960 ;
        RECT 167.920 164.640 168.240 164.960 ;
        RECT 168.320 164.640 168.640 164.960 ;
        RECT 168.720 164.640 169.040 164.960 ;
        RECT 169.120 164.640 169.440 164.960 ;
        RECT 169.520 164.640 169.840 164.960 ;
        RECT 169.920 164.640 170.240 164.960 ;
        RECT 170.320 164.640 170.640 164.960 ;
        RECT 170.720 164.640 171.040 164.960 ;
        RECT 171.120 164.640 171.440 164.960 ;
        RECT 171.520 164.640 171.840 164.960 ;
        RECT 171.920 164.640 172.240 164.960 ;
        RECT 172.320 164.640 172.640 164.960 ;
        RECT 172.720 164.640 173.040 164.960 ;
        RECT 173.120 164.640 173.440 164.960 ;
        RECT 173.520 164.640 173.840 164.960 ;
        RECT 173.920 164.640 174.240 164.960 ;
        RECT 174.320 164.640 174.640 164.960 ;
        RECT 174.720 164.640 175.040 164.960 ;
        RECT 175.120 164.640 175.440 164.960 ;
        RECT 175.520 164.640 175.840 164.960 ;
        RECT 175.920 164.640 176.240 164.960 ;
        RECT 176.320 164.640 176.640 164.960 ;
        RECT 176.720 164.640 177.040 164.960 ;
        RECT 177.120 164.640 177.440 164.960 ;
        RECT 177.520 164.640 177.840 164.960 ;
        RECT 177.920 164.640 178.240 164.960 ;
        RECT 178.320 164.640 178.640 164.960 ;
        RECT 178.720 164.640 179.040 164.960 ;
        RECT 179.120 164.640 179.440 164.960 ;
        RECT 179.520 164.640 179.840 164.960 ;
        RECT 179.920 164.640 180.240 164.960 ;
        RECT 180.320 164.640 180.640 164.960 ;
        RECT 25.040 164.240 25.360 164.560 ;
        RECT 25.440 164.240 25.760 164.560 ;
        RECT 25.840 164.240 26.160 164.560 ;
        RECT 26.240 164.240 26.560 164.560 ;
        RECT 26.640 164.240 26.960 164.560 ;
        RECT 27.040 164.240 27.360 164.560 ;
        RECT 27.440 164.240 27.760 164.560 ;
        RECT 27.840 164.240 28.160 164.560 ;
        RECT 28.240 164.240 28.560 164.560 ;
        RECT 28.640 164.240 28.960 164.560 ;
        RECT 29.040 164.240 29.360 164.560 ;
        RECT 29.440 164.240 29.760 164.560 ;
        RECT 29.840 164.240 30.160 164.560 ;
        RECT 30.240 164.240 30.560 164.560 ;
        RECT 30.640 164.240 30.960 164.560 ;
        RECT 31.040 164.240 31.360 164.560 ;
        RECT 31.440 164.240 31.760 164.560 ;
        RECT 31.840 164.240 32.160 164.560 ;
        RECT 32.240 164.240 32.560 164.560 ;
        RECT 32.640 164.240 32.960 164.560 ;
        RECT 33.040 164.240 33.360 164.560 ;
        RECT 33.440 164.240 33.760 164.560 ;
        RECT 33.840 164.240 34.160 164.560 ;
        RECT 34.240 164.240 34.560 164.560 ;
        RECT 34.640 164.240 34.960 164.560 ;
        RECT 35.040 164.240 35.360 164.560 ;
        RECT 35.440 164.240 35.760 164.560 ;
        RECT 35.840 164.240 36.160 164.560 ;
        RECT 36.240 164.240 36.560 164.560 ;
        RECT 36.640 164.240 36.960 164.560 ;
        RECT 37.040 164.240 37.360 164.560 ;
        RECT 37.440 164.240 37.760 164.560 ;
        RECT 37.840 164.240 38.160 164.560 ;
        RECT 38.240 164.240 38.560 164.560 ;
        RECT 38.640 164.240 38.960 164.560 ;
        RECT 39.040 164.240 39.360 164.560 ;
        RECT 39.440 164.240 39.760 164.560 ;
        RECT 39.840 164.240 40.160 164.560 ;
        RECT 40.240 164.240 40.560 164.560 ;
        RECT 40.640 164.240 40.960 164.560 ;
        RECT 41.040 164.240 41.360 164.560 ;
        RECT 41.440 164.240 41.760 164.560 ;
        RECT 41.840 164.240 42.160 164.560 ;
        RECT 42.240 164.240 42.560 164.560 ;
        RECT 42.640 164.240 42.960 164.560 ;
        RECT 43.040 164.240 43.360 164.560 ;
        RECT 43.440 164.240 43.760 164.560 ;
        RECT 43.840 164.240 44.160 164.560 ;
        RECT 44.240 164.240 44.560 164.560 ;
        RECT 44.640 164.240 44.960 164.560 ;
        RECT 70.560 164.240 70.880 164.560 ;
        RECT 70.960 164.240 71.280 164.560 ;
        RECT 71.360 164.240 71.680 164.560 ;
        RECT 71.760 164.240 72.080 164.560 ;
        RECT 120.560 164.240 120.880 164.560 ;
        RECT 120.960 164.240 121.280 164.560 ;
        RECT 121.360 164.240 121.680 164.560 ;
        RECT 121.760 164.240 122.080 164.560 ;
        RECT 160.720 164.240 161.040 164.560 ;
        RECT 161.120 164.240 161.440 164.560 ;
        RECT 161.520 164.240 161.840 164.560 ;
        RECT 161.920 164.240 162.240 164.560 ;
        RECT 162.320 164.240 162.640 164.560 ;
        RECT 162.720 164.240 163.040 164.560 ;
        RECT 163.120 164.240 163.440 164.560 ;
        RECT 163.520 164.240 163.840 164.560 ;
        RECT 163.920 164.240 164.240 164.560 ;
        RECT 164.320 164.240 164.640 164.560 ;
        RECT 164.720 164.240 165.040 164.560 ;
        RECT 165.120 164.240 165.440 164.560 ;
        RECT 165.520 164.240 165.840 164.560 ;
        RECT 165.920 164.240 166.240 164.560 ;
        RECT 166.320 164.240 166.640 164.560 ;
        RECT 166.720 164.240 167.040 164.560 ;
        RECT 167.120 164.240 167.440 164.560 ;
        RECT 167.520 164.240 167.840 164.560 ;
        RECT 167.920 164.240 168.240 164.560 ;
        RECT 168.320 164.240 168.640 164.560 ;
        RECT 168.720 164.240 169.040 164.560 ;
        RECT 169.120 164.240 169.440 164.560 ;
        RECT 169.520 164.240 169.840 164.560 ;
        RECT 169.920 164.240 170.240 164.560 ;
        RECT 170.320 164.240 170.640 164.560 ;
        RECT 170.720 164.240 171.040 164.560 ;
        RECT 171.120 164.240 171.440 164.560 ;
        RECT 171.520 164.240 171.840 164.560 ;
        RECT 171.920 164.240 172.240 164.560 ;
        RECT 172.320 164.240 172.640 164.560 ;
        RECT 172.720 164.240 173.040 164.560 ;
        RECT 173.120 164.240 173.440 164.560 ;
        RECT 173.520 164.240 173.840 164.560 ;
        RECT 173.920 164.240 174.240 164.560 ;
        RECT 174.320 164.240 174.640 164.560 ;
        RECT 174.720 164.240 175.040 164.560 ;
        RECT 175.120 164.240 175.440 164.560 ;
        RECT 175.520 164.240 175.840 164.560 ;
        RECT 175.920 164.240 176.240 164.560 ;
        RECT 176.320 164.240 176.640 164.560 ;
        RECT 176.720 164.240 177.040 164.560 ;
        RECT 177.120 164.240 177.440 164.560 ;
        RECT 177.520 164.240 177.840 164.560 ;
        RECT 177.920 164.240 178.240 164.560 ;
        RECT 178.320 164.240 178.640 164.560 ;
        RECT 178.720 164.240 179.040 164.560 ;
        RECT 179.120 164.240 179.440 164.560 ;
        RECT 179.520 164.240 179.840 164.560 ;
        RECT 179.920 164.240 180.240 164.560 ;
        RECT 180.320 164.240 180.640 164.560 ;
        RECT 25.040 163.840 25.360 164.160 ;
        RECT 25.440 163.840 25.760 164.160 ;
        RECT 25.840 163.840 26.160 164.160 ;
        RECT 26.240 163.840 26.560 164.160 ;
        RECT 26.640 163.840 26.960 164.160 ;
        RECT 27.040 163.840 27.360 164.160 ;
        RECT 27.440 163.840 27.760 164.160 ;
        RECT 27.840 163.840 28.160 164.160 ;
        RECT 28.240 163.840 28.560 164.160 ;
        RECT 28.640 163.840 28.960 164.160 ;
        RECT 29.040 163.840 29.360 164.160 ;
        RECT 29.440 163.840 29.760 164.160 ;
        RECT 29.840 163.840 30.160 164.160 ;
        RECT 30.240 163.840 30.560 164.160 ;
        RECT 30.640 163.840 30.960 164.160 ;
        RECT 31.040 163.840 31.360 164.160 ;
        RECT 31.440 163.840 31.760 164.160 ;
        RECT 31.840 163.840 32.160 164.160 ;
        RECT 32.240 163.840 32.560 164.160 ;
        RECT 32.640 163.840 32.960 164.160 ;
        RECT 33.040 163.840 33.360 164.160 ;
        RECT 33.440 163.840 33.760 164.160 ;
        RECT 33.840 163.840 34.160 164.160 ;
        RECT 34.240 163.840 34.560 164.160 ;
        RECT 34.640 163.840 34.960 164.160 ;
        RECT 35.040 163.840 35.360 164.160 ;
        RECT 35.440 163.840 35.760 164.160 ;
        RECT 35.840 163.840 36.160 164.160 ;
        RECT 36.240 163.840 36.560 164.160 ;
        RECT 36.640 163.840 36.960 164.160 ;
        RECT 37.040 163.840 37.360 164.160 ;
        RECT 37.440 163.840 37.760 164.160 ;
        RECT 37.840 163.840 38.160 164.160 ;
        RECT 38.240 163.840 38.560 164.160 ;
        RECT 38.640 163.840 38.960 164.160 ;
        RECT 39.040 163.840 39.360 164.160 ;
        RECT 39.440 163.840 39.760 164.160 ;
        RECT 39.840 163.840 40.160 164.160 ;
        RECT 40.240 163.840 40.560 164.160 ;
        RECT 40.640 163.840 40.960 164.160 ;
        RECT 41.040 163.840 41.360 164.160 ;
        RECT 41.440 163.840 41.760 164.160 ;
        RECT 41.840 163.840 42.160 164.160 ;
        RECT 42.240 163.840 42.560 164.160 ;
        RECT 42.640 163.840 42.960 164.160 ;
        RECT 43.040 163.840 43.360 164.160 ;
        RECT 43.440 163.840 43.760 164.160 ;
        RECT 43.840 163.840 44.160 164.160 ;
        RECT 44.240 163.840 44.560 164.160 ;
        RECT 44.640 163.840 44.960 164.160 ;
        RECT 70.560 163.840 70.880 164.160 ;
        RECT 70.960 163.840 71.280 164.160 ;
        RECT 71.360 163.840 71.680 164.160 ;
        RECT 71.760 163.840 72.080 164.160 ;
        RECT 120.560 163.840 120.880 164.160 ;
        RECT 120.960 163.840 121.280 164.160 ;
        RECT 121.360 163.840 121.680 164.160 ;
        RECT 121.760 163.840 122.080 164.160 ;
        RECT 160.720 163.840 161.040 164.160 ;
        RECT 161.120 163.840 161.440 164.160 ;
        RECT 161.520 163.840 161.840 164.160 ;
        RECT 161.920 163.840 162.240 164.160 ;
        RECT 162.320 163.840 162.640 164.160 ;
        RECT 162.720 163.840 163.040 164.160 ;
        RECT 163.120 163.840 163.440 164.160 ;
        RECT 163.520 163.840 163.840 164.160 ;
        RECT 163.920 163.840 164.240 164.160 ;
        RECT 164.320 163.840 164.640 164.160 ;
        RECT 164.720 163.840 165.040 164.160 ;
        RECT 165.120 163.840 165.440 164.160 ;
        RECT 165.520 163.840 165.840 164.160 ;
        RECT 165.920 163.840 166.240 164.160 ;
        RECT 166.320 163.840 166.640 164.160 ;
        RECT 166.720 163.840 167.040 164.160 ;
        RECT 167.120 163.840 167.440 164.160 ;
        RECT 167.520 163.840 167.840 164.160 ;
        RECT 167.920 163.840 168.240 164.160 ;
        RECT 168.320 163.840 168.640 164.160 ;
        RECT 168.720 163.840 169.040 164.160 ;
        RECT 169.120 163.840 169.440 164.160 ;
        RECT 169.520 163.840 169.840 164.160 ;
        RECT 169.920 163.840 170.240 164.160 ;
        RECT 170.320 163.840 170.640 164.160 ;
        RECT 170.720 163.840 171.040 164.160 ;
        RECT 171.120 163.840 171.440 164.160 ;
        RECT 171.520 163.840 171.840 164.160 ;
        RECT 171.920 163.840 172.240 164.160 ;
        RECT 172.320 163.840 172.640 164.160 ;
        RECT 172.720 163.840 173.040 164.160 ;
        RECT 173.120 163.840 173.440 164.160 ;
        RECT 173.520 163.840 173.840 164.160 ;
        RECT 173.920 163.840 174.240 164.160 ;
        RECT 174.320 163.840 174.640 164.160 ;
        RECT 174.720 163.840 175.040 164.160 ;
        RECT 175.120 163.840 175.440 164.160 ;
        RECT 175.520 163.840 175.840 164.160 ;
        RECT 175.920 163.840 176.240 164.160 ;
        RECT 176.320 163.840 176.640 164.160 ;
        RECT 176.720 163.840 177.040 164.160 ;
        RECT 177.120 163.840 177.440 164.160 ;
        RECT 177.520 163.840 177.840 164.160 ;
        RECT 177.920 163.840 178.240 164.160 ;
        RECT 178.320 163.840 178.640 164.160 ;
        RECT 178.720 163.840 179.040 164.160 ;
        RECT 179.120 163.840 179.440 164.160 ;
        RECT 179.520 163.840 179.840 164.160 ;
        RECT 179.920 163.840 180.240 164.160 ;
        RECT 180.320 163.840 180.640 164.160 ;
        RECT 25.040 163.440 25.360 163.760 ;
        RECT 25.440 163.440 25.760 163.760 ;
        RECT 25.840 163.440 26.160 163.760 ;
        RECT 26.240 163.440 26.560 163.760 ;
        RECT 26.640 163.440 26.960 163.760 ;
        RECT 27.040 163.440 27.360 163.760 ;
        RECT 27.440 163.440 27.760 163.760 ;
        RECT 27.840 163.440 28.160 163.760 ;
        RECT 28.240 163.440 28.560 163.760 ;
        RECT 28.640 163.440 28.960 163.760 ;
        RECT 29.040 163.440 29.360 163.760 ;
        RECT 29.440 163.440 29.760 163.760 ;
        RECT 29.840 163.440 30.160 163.760 ;
        RECT 30.240 163.440 30.560 163.760 ;
        RECT 30.640 163.440 30.960 163.760 ;
        RECT 31.040 163.440 31.360 163.760 ;
        RECT 31.440 163.440 31.760 163.760 ;
        RECT 31.840 163.440 32.160 163.760 ;
        RECT 32.240 163.440 32.560 163.760 ;
        RECT 32.640 163.440 32.960 163.760 ;
        RECT 33.040 163.440 33.360 163.760 ;
        RECT 33.440 163.440 33.760 163.760 ;
        RECT 33.840 163.440 34.160 163.760 ;
        RECT 34.240 163.440 34.560 163.760 ;
        RECT 34.640 163.440 34.960 163.760 ;
        RECT 35.040 163.440 35.360 163.760 ;
        RECT 35.440 163.440 35.760 163.760 ;
        RECT 35.840 163.440 36.160 163.760 ;
        RECT 36.240 163.440 36.560 163.760 ;
        RECT 36.640 163.440 36.960 163.760 ;
        RECT 37.040 163.440 37.360 163.760 ;
        RECT 37.440 163.440 37.760 163.760 ;
        RECT 37.840 163.440 38.160 163.760 ;
        RECT 38.240 163.440 38.560 163.760 ;
        RECT 38.640 163.440 38.960 163.760 ;
        RECT 39.040 163.440 39.360 163.760 ;
        RECT 39.440 163.440 39.760 163.760 ;
        RECT 39.840 163.440 40.160 163.760 ;
        RECT 40.240 163.440 40.560 163.760 ;
        RECT 40.640 163.440 40.960 163.760 ;
        RECT 41.040 163.440 41.360 163.760 ;
        RECT 41.440 163.440 41.760 163.760 ;
        RECT 41.840 163.440 42.160 163.760 ;
        RECT 42.240 163.440 42.560 163.760 ;
        RECT 42.640 163.440 42.960 163.760 ;
        RECT 43.040 163.440 43.360 163.760 ;
        RECT 43.440 163.440 43.760 163.760 ;
        RECT 43.840 163.440 44.160 163.760 ;
        RECT 44.240 163.440 44.560 163.760 ;
        RECT 44.640 163.440 44.960 163.760 ;
        RECT 70.560 163.440 70.880 163.760 ;
        RECT 70.960 163.440 71.280 163.760 ;
        RECT 71.360 163.440 71.680 163.760 ;
        RECT 71.760 163.440 72.080 163.760 ;
        RECT 120.560 163.440 120.880 163.760 ;
        RECT 120.960 163.440 121.280 163.760 ;
        RECT 121.360 163.440 121.680 163.760 ;
        RECT 121.760 163.440 122.080 163.760 ;
        RECT 160.720 163.440 161.040 163.760 ;
        RECT 161.120 163.440 161.440 163.760 ;
        RECT 161.520 163.440 161.840 163.760 ;
        RECT 161.920 163.440 162.240 163.760 ;
        RECT 162.320 163.440 162.640 163.760 ;
        RECT 162.720 163.440 163.040 163.760 ;
        RECT 163.120 163.440 163.440 163.760 ;
        RECT 163.520 163.440 163.840 163.760 ;
        RECT 163.920 163.440 164.240 163.760 ;
        RECT 164.320 163.440 164.640 163.760 ;
        RECT 164.720 163.440 165.040 163.760 ;
        RECT 165.120 163.440 165.440 163.760 ;
        RECT 165.520 163.440 165.840 163.760 ;
        RECT 165.920 163.440 166.240 163.760 ;
        RECT 166.320 163.440 166.640 163.760 ;
        RECT 166.720 163.440 167.040 163.760 ;
        RECT 167.120 163.440 167.440 163.760 ;
        RECT 167.520 163.440 167.840 163.760 ;
        RECT 167.920 163.440 168.240 163.760 ;
        RECT 168.320 163.440 168.640 163.760 ;
        RECT 168.720 163.440 169.040 163.760 ;
        RECT 169.120 163.440 169.440 163.760 ;
        RECT 169.520 163.440 169.840 163.760 ;
        RECT 169.920 163.440 170.240 163.760 ;
        RECT 170.320 163.440 170.640 163.760 ;
        RECT 170.720 163.440 171.040 163.760 ;
        RECT 171.120 163.440 171.440 163.760 ;
        RECT 171.520 163.440 171.840 163.760 ;
        RECT 171.920 163.440 172.240 163.760 ;
        RECT 172.320 163.440 172.640 163.760 ;
        RECT 172.720 163.440 173.040 163.760 ;
        RECT 173.120 163.440 173.440 163.760 ;
        RECT 173.520 163.440 173.840 163.760 ;
        RECT 173.920 163.440 174.240 163.760 ;
        RECT 174.320 163.440 174.640 163.760 ;
        RECT 174.720 163.440 175.040 163.760 ;
        RECT 175.120 163.440 175.440 163.760 ;
        RECT 175.520 163.440 175.840 163.760 ;
        RECT 175.920 163.440 176.240 163.760 ;
        RECT 176.320 163.440 176.640 163.760 ;
        RECT 176.720 163.440 177.040 163.760 ;
        RECT 177.120 163.440 177.440 163.760 ;
        RECT 177.520 163.440 177.840 163.760 ;
        RECT 177.920 163.440 178.240 163.760 ;
        RECT 178.320 163.440 178.640 163.760 ;
        RECT 178.720 163.440 179.040 163.760 ;
        RECT 179.120 163.440 179.440 163.760 ;
        RECT 179.520 163.440 179.840 163.760 ;
        RECT 179.920 163.440 180.240 163.760 ;
        RECT 180.320 163.440 180.640 163.760 ;
        RECT 25.040 163.040 25.360 163.360 ;
        RECT 25.440 163.040 25.760 163.360 ;
        RECT 25.840 163.040 26.160 163.360 ;
        RECT 26.240 163.040 26.560 163.360 ;
        RECT 26.640 163.040 26.960 163.360 ;
        RECT 27.040 163.040 27.360 163.360 ;
        RECT 27.440 163.040 27.760 163.360 ;
        RECT 27.840 163.040 28.160 163.360 ;
        RECT 28.240 163.040 28.560 163.360 ;
        RECT 28.640 163.040 28.960 163.360 ;
        RECT 29.040 163.040 29.360 163.360 ;
        RECT 29.440 163.040 29.760 163.360 ;
        RECT 29.840 163.040 30.160 163.360 ;
        RECT 30.240 163.040 30.560 163.360 ;
        RECT 30.640 163.040 30.960 163.360 ;
        RECT 31.040 163.040 31.360 163.360 ;
        RECT 31.440 163.040 31.760 163.360 ;
        RECT 31.840 163.040 32.160 163.360 ;
        RECT 32.240 163.040 32.560 163.360 ;
        RECT 32.640 163.040 32.960 163.360 ;
        RECT 33.040 163.040 33.360 163.360 ;
        RECT 33.440 163.040 33.760 163.360 ;
        RECT 33.840 163.040 34.160 163.360 ;
        RECT 34.240 163.040 34.560 163.360 ;
        RECT 34.640 163.040 34.960 163.360 ;
        RECT 35.040 163.040 35.360 163.360 ;
        RECT 35.440 163.040 35.760 163.360 ;
        RECT 35.840 163.040 36.160 163.360 ;
        RECT 36.240 163.040 36.560 163.360 ;
        RECT 36.640 163.040 36.960 163.360 ;
        RECT 37.040 163.040 37.360 163.360 ;
        RECT 37.440 163.040 37.760 163.360 ;
        RECT 37.840 163.040 38.160 163.360 ;
        RECT 38.240 163.040 38.560 163.360 ;
        RECT 38.640 163.040 38.960 163.360 ;
        RECT 39.040 163.040 39.360 163.360 ;
        RECT 39.440 163.040 39.760 163.360 ;
        RECT 39.840 163.040 40.160 163.360 ;
        RECT 40.240 163.040 40.560 163.360 ;
        RECT 40.640 163.040 40.960 163.360 ;
        RECT 41.040 163.040 41.360 163.360 ;
        RECT 41.440 163.040 41.760 163.360 ;
        RECT 41.840 163.040 42.160 163.360 ;
        RECT 42.240 163.040 42.560 163.360 ;
        RECT 42.640 163.040 42.960 163.360 ;
        RECT 43.040 163.040 43.360 163.360 ;
        RECT 43.440 163.040 43.760 163.360 ;
        RECT 43.840 163.040 44.160 163.360 ;
        RECT 44.240 163.040 44.560 163.360 ;
        RECT 44.640 163.040 44.960 163.360 ;
        RECT 70.560 163.040 70.880 163.360 ;
        RECT 70.960 163.040 71.280 163.360 ;
        RECT 71.360 163.040 71.680 163.360 ;
        RECT 71.760 163.040 72.080 163.360 ;
        RECT 120.560 163.040 120.880 163.360 ;
        RECT 120.960 163.040 121.280 163.360 ;
        RECT 121.360 163.040 121.680 163.360 ;
        RECT 121.760 163.040 122.080 163.360 ;
        RECT 160.720 163.040 161.040 163.360 ;
        RECT 161.120 163.040 161.440 163.360 ;
        RECT 161.520 163.040 161.840 163.360 ;
        RECT 161.920 163.040 162.240 163.360 ;
        RECT 162.320 163.040 162.640 163.360 ;
        RECT 162.720 163.040 163.040 163.360 ;
        RECT 163.120 163.040 163.440 163.360 ;
        RECT 163.520 163.040 163.840 163.360 ;
        RECT 163.920 163.040 164.240 163.360 ;
        RECT 164.320 163.040 164.640 163.360 ;
        RECT 164.720 163.040 165.040 163.360 ;
        RECT 165.120 163.040 165.440 163.360 ;
        RECT 165.520 163.040 165.840 163.360 ;
        RECT 165.920 163.040 166.240 163.360 ;
        RECT 166.320 163.040 166.640 163.360 ;
        RECT 166.720 163.040 167.040 163.360 ;
        RECT 167.120 163.040 167.440 163.360 ;
        RECT 167.520 163.040 167.840 163.360 ;
        RECT 167.920 163.040 168.240 163.360 ;
        RECT 168.320 163.040 168.640 163.360 ;
        RECT 168.720 163.040 169.040 163.360 ;
        RECT 169.120 163.040 169.440 163.360 ;
        RECT 169.520 163.040 169.840 163.360 ;
        RECT 169.920 163.040 170.240 163.360 ;
        RECT 170.320 163.040 170.640 163.360 ;
        RECT 170.720 163.040 171.040 163.360 ;
        RECT 171.120 163.040 171.440 163.360 ;
        RECT 171.520 163.040 171.840 163.360 ;
        RECT 171.920 163.040 172.240 163.360 ;
        RECT 172.320 163.040 172.640 163.360 ;
        RECT 172.720 163.040 173.040 163.360 ;
        RECT 173.120 163.040 173.440 163.360 ;
        RECT 173.520 163.040 173.840 163.360 ;
        RECT 173.920 163.040 174.240 163.360 ;
        RECT 174.320 163.040 174.640 163.360 ;
        RECT 174.720 163.040 175.040 163.360 ;
        RECT 175.120 163.040 175.440 163.360 ;
        RECT 175.520 163.040 175.840 163.360 ;
        RECT 175.920 163.040 176.240 163.360 ;
        RECT 176.320 163.040 176.640 163.360 ;
        RECT 176.720 163.040 177.040 163.360 ;
        RECT 177.120 163.040 177.440 163.360 ;
        RECT 177.520 163.040 177.840 163.360 ;
        RECT 177.920 163.040 178.240 163.360 ;
        RECT 178.320 163.040 178.640 163.360 ;
        RECT 178.720 163.040 179.040 163.360 ;
        RECT 179.120 163.040 179.440 163.360 ;
        RECT 179.520 163.040 179.840 163.360 ;
        RECT 179.920 163.040 180.240 163.360 ;
        RECT 180.320 163.040 180.640 163.360 ;
        RECT 25.040 162.640 25.360 162.960 ;
        RECT 25.440 162.640 25.760 162.960 ;
        RECT 25.840 162.640 26.160 162.960 ;
        RECT 26.240 162.640 26.560 162.960 ;
        RECT 26.640 162.640 26.960 162.960 ;
        RECT 27.040 162.640 27.360 162.960 ;
        RECT 27.440 162.640 27.760 162.960 ;
        RECT 27.840 162.640 28.160 162.960 ;
        RECT 28.240 162.640 28.560 162.960 ;
        RECT 28.640 162.640 28.960 162.960 ;
        RECT 29.040 162.640 29.360 162.960 ;
        RECT 29.440 162.640 29.760 162.960 ;
        RECT 29.840 162.640 30.160 162.960 ;
        RECT 30.240 162.640 30.560 162.960 ;
        RECT 30.640 162.640 30.960 162.960 ;
        RECT 31.040 162.640 31.360 162.960 ;
        RECT 31.440 162.640 31.760 162.960 ;
        RECT 31.840 162.640 32.160 162.960 ;
        RECT 32.240 162.640 32.560 162.960 ;
        RECT 32.640 162.640 32.960 162.960 ;
        RECT 33.040 162.640 33.360 162.960 ;
        RECT 33.440 162.640 33.760 162.960 ;
        RECT 33.840 162.640 34.160 162.960 ;
        RECT 34.240 162.640 34.560 162.960 ;
        RECT 34.640 162.640 34.960 162.960 ;
        RECT 35.040 162.640 35.360 162.960 ;
        RECT 35.440 162.640 35.760 162.960 ;
        RECT 35.840 162.640 36.160 162.960 ;
        RECT 36.240 162.640 36.560 162.960 ;
        RECT 36.640 162.640 36.960 162.960 ;
        RECT 37.040 162.640 37.360 162.960 ;
        RECT 37.440 162.640 37.760 162.960 ;
        RECT 37.840 162.640 38.160 162.960 ;
        RECT 38.240 162.640 38.560 162.960 ;
        RECT 38.640 162.640 38.960 162.960 ;
        RECT 39.040 162.640 39.360 162.960 ;
        RECT 39.440 162.640 39.760 162.960 ;
        RECT 39.840 162.640 40.160 162.960 ;
        RECT 40.240 162.640 40.560 162.960 ;
        RECT 40.640 162.640 40.960 162.960 ;
        RECT 41.040 162.640 41.360 162.960 ;
        RECT 41.440 162.640 41.760 162.960 ;
        RECT 41.840 162.640 42.160 162.960 ;
        RECT 42.240 162.640 42.560 162.960 ;
        RECT 42.640 162.640 42.960 162.960 ;
        RECT 43.040 162.640 43.360 162.960 ;
        RECT 43.440 162.640 43.760 162.960 ;
        RECT 43.840 162.640 44.160 162.960 ;
        RECT 44.240 162.640 44.560 162.960 ;
        RECT 44.640 162.640 44.960 162.960 ;
        RECT 70.560 162.640 70.880 162.960 ;
        RECT 70.960 162.640 71.280 162.960 ;
        RECT 71.360 162.640 71.680 162.960 ;
        RECT 71.760 162.640 72.080 162.960 ;
        RECT 120.560 162.640 120.880 162.960 ;
        RECT 120.960 162.640 121.280 162.960 ;
        RECT 121.360 162.640 121.680 162.960 ;
        RECT 121.760 162.640 122.080 162.960 ;
        RECT 160.720 162.640 161.040 162.960 ;
        RECT 161.120 162.640 161.440 162.960 ;
        RECT 161.520 162.640 161.840 162.960 ;
        RECT 161.920 162.640 162.240 162.960 ;
        RECT 162.320 162.640 162.640 162.960 ;
        RECT 162.720 162.640 163.040 162.960 ;
        RECT 163.120 162.640 163.440 162.960 ;
        RECT 163.520 162.640 163.840 162.960 ;
        RECT 163.920 162.640 164.240 162.960 ;
        RECT 164.320 162.640 164.640 162.960 ;
        RECT 164.720 162.640 165.040 162.960 ;
        RECT 165.120 162.640 165.440 162.960 ;
        RECT 165.520 162.640 165.840 162.960 ;
        RECT 165.920 162.640 166.240 162.960 ;
        RECT 166.320 162.640 166.640 162.960 ;
        RECT 166.720 162.640 167.040 162.960 ;
        RECT 167.120 162.640 167.440 162.960 ;
        RECT 167.520 162.640 167.840 162.960 ;
        RECT 167.920 162.640 168.240 162.960 ;
        RECT 168.320 162.640 168.640 162.960 ;
        RECT 168.720 162.640 169.040 162.960 ;
        RECT 169.120 162.640 169.440 162.960 ;
        RECT 169.520 162.640 169.840 162.960 ;
        RECT 169.920 162.640 170.240 162.960 ;
        RECT 170.320 162.640 170.640 162.960 ;
        RECT 170.720 162.640 171.040 162.960 ;
        RECT 171.120 162.640 171.440 162.960 ;
        RECT 171.520 162.640 171.840 162.960 ;
        RECT 171.920 162.640 172.240 162.960 ;
        RECT 172.320 162.640 172.640 162.960 ;
        RECT 172.720 162.640 173.040 162.960 ;
        RECT 173.120 162.640 173.440 162.960 ;
        RECT 173.520 162.640 173.840 162.960 ;
        RECT 173.920 162.640 174.240 162.960 ;
        RECT 174.320 162.640 174.640 162.960 ;
        RECT 174.720 162.640 175.040 162.960 ;
        RECT 175.120 162.640 175.440 162.960 ;
        RECT 175.520 162.640 175.840 162.960 ;
        RECT 175.920 162.640 176.240 162.960 ;
        RECT 176.320 162.640 176.640 162.960 ;
        RECT 176.720 162.640 177.040 162.960 ;
        RECT 177.120 162.640 177.440 162.960 ;
        RECT 177.520 162.640 177.840 162.960 ;
        RECT 177.920 162.640 178.240 162.960 ;
        RECT 178.320 162.640 178.640 162.960 ;
        RECT 178.720 162.640 179.040 162.960 ;
        RECT 179.120 162.640 179.440 162.960 ;
        RECT 179.520 162.640 179.840 162.960 ;
        RECT 179.920 162.640 180.240 162.960 ;
        RECT 180.320 162.640 180.640 162.960 ;
        RECT 25.040 162.240 25.360 162.560 ;
        RECT 25.440 162.240 25.760 162.560 ;
        RECT 25.840 162.240 26.160 162.560 ;
        RECT 26.240 162.240 26.560 162.560 ;
        RECT 26.640 162.240 26.960 162.560 ;
        RECT 27.040 162.240 27.360 162.560 ;
        RECT 27.440 162.240 27.760 162.560 ;
        RECT 27.840 162.240 28.160 162.560 ;
        RECT 28.240 162.240 28.560 162.560 ;
        RECT 28.640 162.240 28.960 162.560 ;
        RECT 29.040 162.240 29.360 162.560 ;
        RECT 29.440 162.240 29.760 162.560 ;
        RECT 29.840 162.240 30.160 162.560 ;
        RECT 30.240 162.240 30.560 162.560 ;
        RECT 30.640 162.240 30.960 162.560 ;
        RECT 31.040 162.240 31.360 162.560 ;
        RECT 31.440 162.240 31.760 162.560 ;
        RECT 31.840 162.240 32.160 162.560 ;
        RECT 32.240 162.240 32.560 162.560 ;
        RECT 32.640 162.240 32.960 162.560 ;
        RECT 33.040 162.240 33.360 162.560 ;
        RECT 33.440 162.240 33.760 162.560 ;
        RECT 33.840 162.240 34.160 162.560 ;
        RECT 34.240 162.240 34.560 162.560 ;
        RECT 34.640 162.240 34.960 162.560 ;
        RECT 35.040 162.240 35.360 162.560 ;
        RECT 35.440 162.240 35.760 162.560 ;
        RECT 35.840 162.240 36.160 162.560 ;
        RECT 36.240 162.240 36.560 162.560 ;
        RECT 36.640 162.240 36.960 162.560 ;
        RECT 37.040 162.240 37.360 162.560 ;
        RECT 37.440 162.240 37.760 162.560 ;
        RECT 37.840 162.240 38.160 162.560 ;
        RECT 38.240 162.240 38.560 162.560 ;
        RECT 38.640 162.240 38.960 162.560 ;
        RECT 39.040 162.240 39.360 162.560 ;
        RECT 39.440 162.240 39.760 162.560 ;
        RECT 39.840 162.240 40.160 162.560 ;
        RECT 40.240 162.240 40.560 162.560 ;
        RECT 40.640 162.240 40.960 162.560 ;
        RECT 41.040 162.240 41.360 162.560 ;
        RECT 41.440 162.240 41.760 162.560 ;
        RECT 41.840 162.240 42.160 162.560 ;
        RECT 42.240 162.240 42.560 162.560 ;
        RECT 42.640 162.240 42.960 162.560 ;
        RECT 43.040 162.240 43.360 162.560 ;
        RECT 43.440 162.240 43.760 162.560 ;
        RECT 43.840 162.240 44.160 162.560 ;
        RECT 44.240 162.240 44.560 162.560 ;
        RECT 44.640 162.240 44.960 162.560 ;
        RECT 70.560 162.240 70.880 162.560 ;
        RECT 70.960 162.240 71.280 162.560 ;
        RECT 71.360 162.240 71.680 162.560 ;
        RECT 71.760 162.240 72.080 162.560 ;
        RECT 120.560 162.240 120.880 162.560 ;
        RECT 120.960 162.240 121.280 162.560 ;
        RECT 121.360 162.240 121.680 162.560 ;
        RECT 121.760 162.240 122.080 162.560 ;
        RECT 160.720 162.240 161.040 162.560 ;
        RECT 161.120 162.240 161.440 162.560 ;
        RECT 161.520 162.240 161.840 162.560 ;
        RECT 161.920 162.240 162.240 162.560 ;
        RECT 162.320 162.240 162.640 162.560 ;
        RECT 162.720 162.240 163.040 162.560 ;
        RECT 163.120 162.240 163.440 162.560 ;
        RECT 163.520 162.240 163.840 162.560 ;
        RECT 163.920 162.240 164.240 162.560 ;
        RECT 164.320 162.240 164.640 162.560 ;
        RECT 164.720 162.240 165.040 162.560 ;
        RECT 165.120 162.240 165.440 162.560 ;
        RECT 165.520 162.240 165.840 162.560 ;
        RECT 165.920 162.240 166.240 162.560 ;
        RECT 166.320 162.240 166.640 162.560 ;
        RECT 166.720 162.240 167.040 162.560 ;
        RECT 167.120 162.240 167.440 162.560 ;
        RECT 167.520 162.240 167.840 162.560 ;
        RECT 167.920 162.240 168.240 162.560 ;
        RECT 168.320 162.240 168.640 162.560 ;
        RECT 168.720 162.240 169.040 162.560 ;
        RECT 169.120 162.240 169.440 162.560 ;
        RECT 169.520 162.240 169.840 162.560 ;
        RECT 169.920 162.240 170.240 162.560 ;
        RECT 170.320 162.240 170.640 162.560 ;
        RECT 170.720 162.240 171.040 162.560 ;
        RECT 171.120 162.240 171.440 162.560 ;
        RECT 171.520 162.240 171.840 162.560 ;
        RECT 171.920 162.240 172.240 162.560 ;
        RECT 172.320 162.240 172.640 162.560 ;
        RECT 172.720 162.240 173.040 162.560 ;
        RECT 173.120 162.240 173.440 162.560 ;
        RECT 173.520 162.240 173.840 162.560 ;
        RECT 173.920 162.240 174.240 162.560 ;
        RECT 174.320 162.240 174.640 162.560 ;
        RECT 174.720 162.240 175.040 162.560 ;
        RECT 175.120 162.240 175.440 162.560 ;
        RECT 175.520 162.240 175.840 162.560 ;
        RECT 175.920 162.240 176.240 162.560 ;
        RECT 176.320 162.240 176.640 162.560 ;
        RECT 176.720 162.240 177.040 162.560 ;
        RECT 177.120 162.240 177.440 162.560 ;
        RECT 177.520 162.240 177.840 162.560 ;
        RECT 177.920 162.240 178.240 162.560 ;
        RECT 178.320 162.240 178.640 162.560 ;
        RECT 178.720 162.240 179.040 162.560 ;
        RECT 179.120 162.240 179.440 162.560 ;
        RECT 179.520 162.240 179.840 162.560 ;
        RECT 179.920 162.240 180.240 162.560 ;
        RECT 180.320 162.240 180.640 162.560 ;
        RECT 25.040 161.840 25.360 162.160 ;
        RECT 25.440 161.840 25.760 162.160 ;
        RECT 25.840 161.840 26.160 162.160 ;
        RECT 26.240 161.840 26.560 162.160 ;
        RECT 26.640 161.840 26.960 162.160 ;
        RECT 27.040 161.840 27.360 162.160 ;
        RECT 27.440 161.840 27.760 162.160 ;
        RECT 27.840 161.840 28.160 162.160 ;
        RECT 28.240 161.840 28.560 162.160 ;
        RECT 28.640 161.840 28.960 162.160 ;
        RECT 29.040 161.840 29.360 162.160 ;
        RECT 29.440 161.840 29.760 162.160 ;
        RECT 29.840 161.840 30.160 162.160 ;
        RECT 30.240 161.840 30.560 162.160 ;
        RECT 30.640 161.840 30.960 162.160 ;
        RECT 31.040 161.840 31.360 162.160 ;
        RECT 31.440 161.840 31.760 162.160 ;
        RECT 31.840 161.840 32.160 162.160 ;
        RECT 32.240 161.840 32.560 162.160 ;
        RECT 32.640 161.840 32.960 162.160 ;
        RECT 33.040 161.840 33.360 162.160 ;
        RECT 33.440 161.840 33.760 162.160 ;
        RECT 33.840 161.840 34.160 162.160 ;
        RECT 34.240 161.840 34.560 162.160 ;
        RECT 34.640 161.840 34.960 162.160 ;
        RECT 35.040 161.840 35.360 162.160 ;
        RECT 35.440 161.840 35.760 162.160 ;
        RECT 35.840 161.840 36.160 162.160 ;
        RECT 36.240 161.840 36.560 162.160 ;
        RECT 36.640 161.840 36.960 162.160 ;
        RECT 37.040 161.840 37.360 162.160 ;
        RECT 37.440 161.840 37.760 162.160 ;
        RECT 37.840 161.840 38.160 162.160 ;
        RECT 38.240 161.840 38.560 162.160 ;
        RECT 38.640 161.840 38.960 162.160 ;
        RECT 39.040 161.840 39.360 162.160 ;
        RECT 39.440 161.840 39.760 162.160 ;
        RECT 39.840 161.840 40.160 162.160 ;
        RECT 40.240 161.840 40.560 162.160 ;
        RECT 40.640 161.840 40.960 162.160 ;
        RECT 41.040 161.840 41.360 162.160 ;
        RECT 41.440 161.840 41.760 162.160 ;
        RECT 41.840 161.840 42.160 162.160 ;
        RECT 42.240 161.840 42.560 162.160 ;
        RECT 42.640 161.840 42.960 162.160 ;
        RECT 43.040 161.840 43.360 162.160 ;
        RECT 43.440 161.840 43.760 162.160 ;
        RECT 43.840 161.840 44.160 162.160 ;
        RECT 44.240 161.840 44.560 162.160 ;
        RECT 44.640 161.840 44.960 162.160 ;
        RECT 70.560 161.840 70.880 162.160 ;
        RECT 70.960 161.840 71.280 162.160 ;
        RECT 71.360 161.840 71.680 162.160 ;
        RECT 71.760 161.840 72.080 162.160 ;
        RECT 120.560 161.840 120.880 162.160 ;
        RECT 120.960 161.840 121.280 162.160 ;
        RECT 121.360 161.840 121.680 162.160 ;
        RECT 121.760 161.840 122.080 162.160 ;
        RECT 160.720 161.840 161.040 162.160 ;
        RECT 161.120 161.840 161.440 162.160 ;
        RECT 161.520 161.840 161.840 162.160 ;
        RECT 161.920 161.840 162.240 162.160 ;
        RECT 162.320 161.840 162.640 162.160 ;
        RECT 162.720 161.840 163.040 162.160 ;
        RECT 163.120 161.840 163.440 162.160 ;
        RECT 163.520 161.840 163.840 162.160 ;
        RECT 163.920 161.840 164.240 162.160 ;
        RECT 164.320 161.840 164.640 162.160 ;
        RECT 164.720 161.840 165.040 162.160 ;
        RECT 165.120 161.840 165.440 162.160 ;
        RECT 165.520 161.840 165.840 162.160 ;
        RECT 165.920 161.840 166.240 162.160 ;
        RECT 166.320 161.840 166.640 162.160 ;
        RECT 166.720 161.840 167.040 162.160 ;
        RECT 167.120 161.840 167.440 162.160 ;
        RECT 167.520 161.840 167.840 162.160 ;
        RECT 167.920 161.840 168.240 162.160 ;
        RECT 168.320 161.840 168.640 162.160 ;
        RECT 168.720 161.840 169.040 162.160 ;
        RECT 169.120 161.840 169.440 162.160 ;
        RECT 169.520 161.840 169.840 162.160 ;
        RECT 169.920 161.840 170.240 162.160 ;
        RECT 170.320 161.840 170.640 162.160 ;
        RECT 170.720 161.840 171.040 162.160 ;
        RECT 171.120 161.840 171.440 162.160 ;
        RECT 171.520 161.840 171.840 162.160 ;
        RECT 171.920 161.840 172.240 162.160 ;
        RECT 172.320 161.840 172.640 162.160 ;
        RECT 172.720 161.840 173.040 162.160 ;
        RECT 173.120 161.840 173.440 162.160 ;
        RECT 173.520 161.840 173.840 162.160 ;
        RECT 173.920 161.840 174.240 162.160 ;
        RECT 174.320 161.840 174.640 162.160 ;
        RECT 174.720 161.840 175.040 162.160 ;
        RECT 175.120 161.840 175.440 162.160 ;
        RECT 175.520 161.840 175.840 162.160 ;
        RECT 175.920 161.840 176.240 162.160 ;
        RECT 176.320 161.840 176.640 162.160 ;
        RECT 176.720 161.840 177.040 162.160 ;
        RECT 177.120 161.840 177.440 162.160 ;
        RECT 177.520 161.840 177.840 162.160 ;
        RECT 177.920 161.840 178.240 162.160 ;
        RECT 178.320 161.840 178.640 162.160 ;
        RECT 178.720 161.840 179.040 162.160 ;
        RECT 179.120 161.840 179.440 162.160 ;
        RECT 179.520 161.840 179.840 162.160 ;
        RECT 179.920 161.840 180.240 162.160 ;
        RECT 180.320 161.840 180.640 162.160 ;
        RECT 25.040 161.440 25.360 161.760 ;
        RECT 25.440 161.440 25.760 161.760 ;
        RECT 25.840 161.440 26.160 161.760 ;
        RECT 26.240 161.440 26.560 161.760 ;
        RECT 26.640 161.440 26.960 161.760 ;
        RECT 27.040 161.440 27.360 161.760 ;
        RECT 27.440 161.440 27.760 161.760 ;
        RECT 27.840 161.440 28.160 161.760 ;
        RECT 28.240 161.440 28.560 161.760 ;
        RECT 28.640 161.440 28.960 161.760 ;
        RECT 29.040 161.440 29.360 161.760 ;
        RECT 29.440 161.440 29.760 161.760 ;
        RECT 29.840 161.440 30.160 161.760 ;
        RECT 30.240 161.440 30.560 161.760 ;
        RECT 30.640 161.440 30.960 161.760 ;
        RECT 31.040 161.440 31.360 161.760 ;
        RECT 31.440 161.440 31.760 161.760 ;
        RECT 31.840 161.440 32.160 161.760 ;
        RECT 32.240 161.440 32.560 161.760 ;
        RECT 32.640 161.440 32.960 161.760 ;
        RECT 33.040 161.440 33.360 161.760 ;
        RECT 33.440 161.440 33.760 161.760 ;
        RECT 33.840 161.440 34.160 161.760 ;
        RECT 34.240 161.440 34.560 161.760 ;
        RECT 34.640 161.440 34.960 161.760 ;
        RECT 35.040 161.440 35.360 161.760 ;
        RECT 35.440 161.440 35.760 161.760 ;
        RECT 35.840 161.440 36.160 161.760 ;
        RECT 36.240 161.440 36.560 161.760 ;
        RECT 36.640 161.440 36.960 161.760 ;
        RECT 37.040 161.440 37.360 161.760 ;
        RECT 37.440 161.440 37.760 161.760 ;
        RECT 37.840 161.440 38.160 161.760 ;
        RECT 38.240 161.440 38.560 161.760 ;
        RECT 38.640 161.440 38.960 161.760 ;
        RECT 39.040 161.440 39.360 161.760 ;
        RECT 39.440 161.440 39.760 161.760 ;
        RECT 39.840 161.440 40.160 161.760 ;
        RECT 40.240 161.440 40.560 161.760 ;
        RECT 40.640 161.440 40.960 161.760 ;
        RECT 41.040 161.440 41.360 161.760 ;
        RECT 41.440 161.440 41.760 161.760 ;
        RECT 41.840 161.440 42.160 161.760 ;
        RECT 42.240 161.440 42.560 161.760 ;
        RECT 42.640 161.440 42.960 161.760 ;
        RECT 43.040 161.440 43.360 161.760 ;
        RECT 43.440 161.440 43.760 161.760 ;
        RECT 43.840 161.440 44.160 161.760 ;
        RECT 44.240 161.440 44.560 161.760 ;
        RECT 44.640 161.440 44.960 161.760 ;
        RECT 70.560 161.440 70.880 161.760 ;
        RECT 70.960 161.440 71.280 161.760 ;
        RECT 71.360 161.440 71.680 161.760 ;
        RECT 71.760 161.440 72.080 161.760 ;
        RECT 120.560 161.440 120.880 161.760 ;
        RECT 120.960 161.440 121.280 161.760 ;
        RECT 121.360 161.440 121.680 161.760 ;
        RECT 121.760 161.440 122.080 161.760 ;
        RECT 160.720 161.440 161.040 161.760 ;
        RECT 161.120 161.440 161.440 161.760 ;
        RECT 161.520 161.440 161.840 161.760 ;
        RECT 161.920 161.440 162.240 161.760 ;
        RECT 162.320 161.440 162.640 161.760 ;
        RECT 162.720 161.440 163.040 161.760 ;
        RECT 163.120 161.440 163.440 161.760 ;
        RECT 163.520 161.440 163.840 161.760 ;
        RECT 163.920 161.440 164.240 161.760 ;
        RECT 164.320 161.440 164.640 161.760 ;
        RECT 164.720 161.440 165.040 161.760 ;
        RECT 165.120 161.440 165.440 161.760 ;
        RECT 165.520 161.440 165.840 161.760 ;
        RECT 165.920 161.440 166.240 161.760 ;
        RECT 166.320 161.440 166.640 161.760 ;
        RECT 166.720 161.440 167.040 161.760 ;
        RECT 167.120 161.440 167.440 161.760 ;
        RECT 167.520 161.440 167.840 161.760 ;
        RECT 167.920 161.440 168.240 161.760 ;
        RECT 168.320 161.440 168.640 161.760 ;
        RECT 168.720 161.440 169.040 161.760 ;
        RECT 169.120 161.440 169.440 161.760 ;
        RECT 169.520 161.440 169.840 161.760 ;
        RECT 169.920 161.440 170.240 161.760 ;
        RECT 170.320 161.440 170.640 161.760 ;
        RECT 170.720 161.440 171.040 161.760 ;
        RECT 171.120 161.440 171.440 161.760 ;
        RECT 171.520 161.440 171.840 161.760 ;
        RECT 171.920 161.440 172.240 161.760 ;
        RECT 172.320 161.440 172.640 161.760 ;
        RECT 172.720 161.440 173.040 161.760 ;
        RECT 173.120 161.440 173.440 161.760 ;
        RECT 173.520 161.440 173.840 161.760 ;
        RECT 173.920 161.440 174.240 161.760 ;
        RECT 174.320 161.440 174.640 161.760 ;
        RECT 174.720 161.440 175.040 161.760 ;
        RECT 175.120 161.440 175.440 161.760 ;
        RECT 175.520 161.440 175.840 161.760 ;
        RECT 175.920 161.440 176.240 161.760 ;
        RECT 176.320 161.440 176.640 161.760 ;
        RECT 176.720 161.440 177.040 161.760 ;
        RECT 177.120 161.440 177.440 161.760 ;
        RECT 177.520 161.440 177.840 161.760 ;
        RECT 177.920 161.440 178.240 161.760 ;
        RECT 178.320 161.440 178.640 161.760 ;
        RECT 178.720 161.440 179.040 161.760 ;
        RECT 179.120 161.440 179.440 161.760 ;
        RECT 179.520 161.440 179.840 161.760 ;
        RECT 179.920 161.440 180.240 161.760 ;
        RECT 180.320 161.440 180.640 161.760 ;
        RECT 25.040 161.040 25.360 161.360 ;
        RECT 25.440 161.040 25.760 161.360 ;
        RECT 25.840 161.040 26.160 161.360 ;
        RECT 26.240 161.040 26.560 161.360 ;
        RECT 26.640 161.040 26.960 161.360 ;
        RECT 27.040 161.040 27.360 161.360 ;
        RECT 27.440 161.040 27.760 161.360 ;
        RECT 27.840 161.040 28.160 161.360 ;
        RECT 28.240 161.040 28.560 161.360 ;
        RECT 28.640 161.040 28.960 161.360 ;
        RECT 29.040 161.040 29.360 161.360 ;
        RECT 29.440 161.040 29.760 161.360 ;
        RECT 29.840 161.040 30.160 161.360 ;
        RECT 30.240 161.040 30.560 161.360 ;
        RECT 30.640 161.040 30.960 161.360 ;
        RECT 31.040 161.040 31.360 161.360 ;
        RECT 31.440 161.040 31.760 161.360 ;
        RECT 31.840 161.040 32.160 161.360 ;
        RECT 32.240 161.040 32.560 161.360 ;
        RECT 32.640 161.040 32.960 161.360 ;
        RECT 33.040 161.040 33.360 161.360 ;
        RECT 33.440 161.040 33.760 161.360 ;
        RECT 33.840 161.040 34.160 161.360 ;
        RECT 34.240 161.040 34.560 161.360 ;
        RECT 34.640 161.040 34.960 161.360 ;
        RECT 35.040 161.040 35.360 161.360 ;
        RECT 35.440 161.040 35.760 161.360 ;
        RECT 35.840 161.040 36.160 161.360 ;
        RECT 36.240 161.040 36.560 161.360 ;
        RECT 36.640 161.040 36.960 161.360 ;
        RECT 37.040 161.040 37.360 161.360 ;
        RECT 37.440 161.040 37.760 161.360 ;
        RECT 37.840 161.040 38.160 161.360 ;
        RECT 38.240 161.040 38.560 161.360 ;
        RECT 38.640 161.040 38.960 161.360 ;
        RECT 39.040 161.040 39.360 161.360 ;
        RECT 39.440 161.040 39.760 161.360 ;
        RECT 39.840 161.040 40.160 161.360 ;
        RECT 40.240 161.040 40.560 161.360 ;
        RECT 40.640 161.040 40.960 161.360 ;
        RECT 41.040 161.040 41.360 161.360 ;
        RECT 41.440 161.040 41.760 161.360 ;
        RECT 41.840 161.040 42.160 161.360 ;
        RECT 42.240 161.040 42.560 161.360 ;
        RECT 42.640 161.040 42.960 161.360 ;
        RECT 43.040 161.040 43.360 161.360 ;
        RECT 43.440 161.040 43.760 161.360 ;
        RECT 43.840 161.040 44.160 161.360 ;
        RECT 44.240 161.040 44.560 161.360 ;
        RECT 44.640 161.040 44.960 161.360 ;
        RECT 70.560 161.040 70.880 161.360 ;
        RECT 70.960 161.040 71.280 161.360 ;
        RECT 71.360 161.040 71.680 161.360 ;
        RECT 71.760 161.040 72.080 161.360 ;
        RECT 120.560 161.040 120.880 161.360 ;
        RECT 120.960 161.040 121.280 161.360 ;
        RECT 121.360 161.040 121.680 161.360 ;
        RECT 121.760 161.040 122.080 161.360 ;
        RECT 160.720 161.040 161.040 161.360 ;
        RECT 161.120 161.040 161.440 161.360 ;
        RECT 161.520 161.040 161.840 161.360 ;
        RECT 161.920 161.040 162.240 161.360 ;
        RECT 162.320 161.040 162.640 161.360 ;
        RECT 162.720 161.040 163.040 161.360 ;
        RECT 163.120 161.040 163.440 161.360 ;
        RECT 163.520 161.040 163.840 161.360 ;
        RECT 163.920 161.040 164.240 161.360 ;
        RECT 164.320 161.040 164.640 161.360 ;
        RECT 164.720 161.040 165.040 161.360 ;
        RECT 165.120 161.040 165.440 161.360 ;
        RECT 165.520 161.040 165.840 161.360 ;
        RECT 165.920 161.040 166.240 161.360 ;
        RECT 166.320 161.040 166.640 161.360 ;
        RECT 166.720 161.040 167.040 161.360 ;
        RECT 167.120 161.040 167.440 161.360 ;
        RECT 167.520 161.040 167.840 161.360 ;
        RECT 167.920 161.040 168.240 161.360 ;
        RECT 168.320 161.040 168.640 161.360 ;
        RECT 168.720 161.040 169.040 161.360 ;
        RECT 169.120 161.040 169.440 161.360 ;
        RECT 169.520 161.040 169.840 161.360 ;
        RECT 169.920 161.040 170.240 161.360 ;
        RECT 170.320 161.040 170.640 161.360 ;
        RECT 170.720 161.040 171.040 161.360 ;
        RECT 171.120 161.040 171.440 161.360 ;
        RECT 171.520 161.040 171.840 161.360 ;
        RECT 171.920 161.040 172.240 161.360 ;
        RECT 172.320 161.040 172.640 161.360 ;
        RECT 172.720 161.040 173.040 161.360 ;
        RECT 173.120 161.040 173.440 161.360 ;
        RECT 173.520 161.040 173.840 161.360 ;
        RECT 173.920 161.040 174.240 161.360 ;
        RECT 174.320 161.040 174.640 161.360 ;
        RECT 174.720 161.040 175.040 161.360 ;
        RECT 175.120 161.040 175.440 161.360 ;
        RECT 175.520 161.040 175.840 161.360 ;
        RECT 175.920 161.040 176.240 161.360 ;
        RECT 176.320 161.040 176.640 161.360 ;
        RECT 176.720 161.040 177.040 161.360 ;
        RECT 177.120 161.040 177.440 161.360 ;
        RECT 177.520 161.040 177.840 161.360 ;
        RECT 177.920 161.040 178.240 161.360 ;
        RECT 178.320 161.040 178.640 161.360 ;
        RECT 178.720 161.040 179.040 161.360 ;
        RECT 179.120 161.040 179.440 161.360 ;
        RECT 179.520 161.040 179.840 161.360 ;
        RECT 179.920 161.040 180.240 161.360 ;
        RECT 180.320 161.040 180.640 161.360 ;
        RECT 25.040 160.640 25.360 160.960 ;
        RECT 25.440 160.640 25.760 160.960 ;
        RECT 25.840 160.640 26.160 160.960 ;
        RECT 26.240 160.640 26.560 160.960 ;
        RECT 26.640 160.640 26.960 160.960 ;
        RECT 27.040 160.640 27.360 160.960 ;
        RECT 27.440 160.640 27.760 160.960 ;
        RECT 27.840 160.640 28.160 160.960 ;
        RECT 28.240 160.640 28.560 160.960 ;
        RECT 28.640 160.640 28.960 160.960 ;
        RECT 29.040 160.640 29.360 160.960 ;
        RECT 29.440 160.640 29.760 160.960 ;
        RECT 29.840 160.640 30.160 160.960 ;
        RECT 30.240 160.640 30.560 160.960 ;
        RECT 30.640 160.640 30.960 160.960 ;
        RECT 31.040 160.640 31.360 160.960 ;
        RECT 31.440 160.640 31.760 160.960 ;
        RECT 31.840 160.640 32.160 160.960 ;
        RECT 32.240 160.640 32.560 160.960 ;
        RECT 32.640 160.640 32.960 160.960 ;
        RECT 33.040 160.640 33.360 160.960 ;
        RECT 33.440 160.640 33.760 160.960 ;
        RECT 33.840 160.640 34.160 160.960 ;
        RECT 34.240 160.640 34.560 160.960 ;
        RECT 34.640 160.640 34.960 160.960 ;
        RECT 35.040 160.640 35.360 160.960 ;
        RECT 35.440 160.640 35.760 160.960 ;
        RECT 35.840 160.640 36.160 160.960 ;
        RECT 36.240 160.640 36.560 160.960 ;
        RECT 36.640 160.640 36.960 160.960 ;
        RECT 37.040 160.640 37.360 160.960 ;
        RECT 37.440 160.640 37.760 160.960 ;
        RECT 37.840 160.640 38.160 160.960 ;
        RECT 38.240 160.640 38.560 160.960 ;
        RECT 38.640 160.640 38.960 160.960 ;
        RECT 39.040 160.640 39.360 160.960 ;
        RECT 39.440 160.640 39.760 160.960 ;
        RECT 39.840 160.640 40.160 160.960 ;
        RECT 40.240 160.640 40.560 160.960 ;
        RECT 40.640 160.640 40.960 160.960 ;
        RECT 41.040 160.640 41.360 160.960 ;
        RECT 41.440 160.640 41.760 160.960 ;
        RECT 41.840 160.640 42.160 160.960 ;
        RECT 42.240 160.640 42.560 160.960 ;
        RECT 42.640 160.640 42.960 160.960 ;
        RECT 43.040 160.640 43.360 160.960 ;
        RECT 43.440 160.640 43.760 160.960 ;
        RECT 43.840 160.640 44.160 160.960 ;
        RECT 44.240 160.640 44.560 160.960 ;
        RECT 44.640 160.640 44.960 160.960 ;
        RECT 70.560 160.640 70.880 160.960 ;
        RECT 70.960 160.640 71.280 160.960 ;
        RECT 71.360 160.640 71.680 160.960 ;
        RECT 71.760 160.640 72.080 160.960 ;
        RECT 120.560 160.640 120.880 160.960 ;
        RECT 120.960 160.640 121.280 160.960 ;
        RECT 121.360 160.640 121.680 160.960 ;
        RECT 121.760 160.640 122.080 160.960 ;
        RECT 160.720 160.640 161.040 160.960 ;
        RECT 161.120 160.640 161.440 160.960 ;
        RECT 161.520 160.640 161.840 160.960 ;
        RECT 161.920 160.640 162.240 160.960 ;
        RECT 162.320 160.640 162.640 160.960 ;
        RECT 162.720 160.640 163.040 160.960 ;
        RECT 163.120 160.640 163.440 160.960 ;
        RECT 163.520 160.640 163.840 160.960 ;
        RECT 163.920 160.640 164.240 160.960 ;
        RECT 164.320 160.640 164.640 160.960 ;
        RECT 164.720 160.640 165.040 160.960 ;
        RECT 165.120 160.640 165.440 160.960 ;
        RECT 165.520 160.640 165.840 160.960 ;
        RECT 165.920 160.640 166.240 160.960 ;
        RECT 166.320 160.640 166.640 160.960 ;
        RECT 166.720 160.640 167.040 160.960 ;
        RECT 167.120 160.640 167.440 160.960 ;
        RECT 167.520 160.640 167.840 160.960 ;
        RECT 167.920 160.640 168.240 160.960 ;
        RECT 168.320 160.640 168.640 160.960 ;
        RECT 168.720 160.640 169.040 160.960 ;
        RECT 169.120 160.640 169.440 160.960 ;
        RECT 169.520 160.640 169.840 160.960 ;
        RECT 169.920 160.640 170.240 160.960 ;
        RECT 170.320 160.640 170.640 160.960 ;
        RECT 170.720 160.640 171.040 160.960 ;
        RECT 171.120 160.640 171.440 160.960 ;
        RECT 171.520 160.640 171.840 160.960 ;
        RECT 171.920 160.640 172.240 160.960 ;
        RECT 172.320 160.640 172.640 160.960 ;
        RECT 172.720 160.640 173.040 160.960 ;
        RECT 173.120 160.640 173.440 160.960 ;
        RECT 173.520 160.640 173.840 160.960 ;
        RECT 173.920 160.640 174.240 160.960 ;
        RECT 174.320 160.640 174.640 160.960 ;
        RECT 174.720 160.640 175.040 160.960 ;
        RECT 175.120 160.640 175.440 160.960 ;
        RECT 175.520 160.640 175.840 160.960 ;
        RECT 175.920 160.640 176.240 160.960 ;
        RECT 176.320 160.640 176.640 160.960 ;
        RECT 176.720 160.640 177.040 160.960 ;
        RECT 177.120 160.640 177.440 160.960 ;
        RECT 177.520 160.640 177.840 160.960 ;
        RECT 177.920 160.640 178.240 160.960 ;
        RECT 178.320 160.640 178.640 160.960 ;
        RECT 178.720 160.640 179.040 160.960 ;
        RECT 179.120 160.640 179.440 160.960 ;
        RECT 179.520 160.640 179.840 160.960 ;
        RECT 179.920 160.640 180.240 160.960 ;
        RECT 180.320 160.640 180.640 160.960 ;
        RECT 25.040 160.240 25.360 160.560 ;
        RECT 25.440 160.240 25.760 160.560 ;
        RECT 25.840 160.240 26.160 160.560 ;
        RECT 26.240 160.240 26.560 160.560 ;
        RECT 26.640 160.240 26.960 160.560 ;
        RECT 27.040 160.240 27.360 160.560 ;
        RECT 27.440 160.240 27.760 160.560 ;
        RECT 27.840 160.240 28.160 160.560 ;
        RECT 28.240 160.240 28.560 160.560 ;
        RECT 28.640 160.240 28.960 160.560 ;
        RECT 29.040 160.240 29.360 160.560 ;
        RECT 29.440 160.240 29.760 160.560 ;
        RECT 29.840 160.240 30.160 160.560 ;
        RECT 30.240 160.240 30.560 160.560 ;
        RECT 30.640 160.240 30.960 160.560 ;
        RECT 31.040 160.240 31.360 160.560 ;
        RECT 31.440 160.240 31.760 160.560 ;
        RECT 31.840 160.240 32.160 160.560 ;
        RECT 32.240 160.240 32.560 160.560 ;
        RECT 32.640 160.240 32.960 160.560 ;
        RECT 33.040 160.240 33.360 160.560 ;
        RECT 33.440 160.240 33.760 160.560 ;
        RECT 33.840 160.240 34.160 160.560 ;
        RECT 34.240 160.240 34.560 160.560 ;
        RECT 34.640 160.240 34.960 160.560 ;
        RECT 35.040 160.240 35.360 160.560 ;
        RECT 35.440 160.240 35.760 160.560 ;
        RECT 35.840 160.240 36.160 160.560 ;
        RECT 36.240 160.240 36.560 160.560 ;
        RECT 36.640 160.240 36.960 160.560 ;
        RECT 37.040 160.240 37.360 160.560 ;
        RECT 37.440 160.240 37.760 160.560 ;
        RECT 37.840 160.240 38.160 160.560 ;
        RECT 38.240 160.240 38.560 160.560 ;
        RECT 38.640 160.240 38.960 160.560 ;
        RECT 39.040 160.240 39.360 160.560 ;
        RECT 39.440 160.240 39.760 160.560 ;
        RECT 39.840 160.240 40.160 160.560 ;
        RECT 40.240 160.240 40.560 160.560 ;
        RECT 40.640 160.240 40.960 160.560 ;
        RECT 41.040 160.240 41.360 160.560 ;
        RECT 41.440 160.240 41.760 160.560 ;
        RECT 41.840 160.240 42.160 160.560 ;
        RECT 42.240 160.240 42.560 160.560 ;
        RECT 42.640 160.240 42.960 160.560 ;
        RECT 43.040 160.240 43.360 160.560 ;
        RECT 43.440 160.240 43.760 160.560 ;
        RECT 43.840 160.240 44.160 160.560 ;
        RECT 44.240 160.240 44.560 160.560 ;
        RECT 44.640 160.240 44.960 160.560 ;
        RECT 70.560 160.240 70.880 160.560 ;
        RECT 70.960 160.240 71.280 160.560 ;
        RECT 71.360 160.240 71.680 160.560 ;
        RECT 71.760 160.240 72.080 160.560 ;
        RECT 120.560 160.240 120.880 160.560 ;
        RECT 120.960 160.240 121.280 160.560 ;
        RECT 121.360 160.240 121.680 160.560 ;
        RECT 121.760 160.240 122.080 160.560 ;
        RECT 160.720 160.240 161.040 160.560 ;
        RECT 161.120 160.240 161.440 160.560 ;
        RECT 161.520 160.240 161.840 160.560 ;
        RECT 161.920 160.240 162.240 160.560 ;
        RECT 162.320 160.240 162.640 160.560 ;
        RECT 162.720 160.240 163.040 160.560 ;
        RECT 163.120 160.240 163.440 160.560 ;
        RECT 163.520 160.240 163.840 160.560 ;
        RECT 163.920 160.240 164.240 160.560 ;
        RECT 164.320 160.240 164.640 160.560 ;
        RECT 164.720 160.240 165.040 160.560 ;
        RECT 165.120 160.240 165.440 160.560 ;
        RECT 165.520 160.240 165.840 160.560 ;
        RECT 165.920 160.240 166.240 160.560 ;
        RECT 166.320 160.240 166.640 160.560 ;
        RECT 166.720 160.240 167.040 160.560 ;
        RECT 167.120 160.240 167.440 160.560 ;
        RECT 167.520 160.240 167.840 160.560 ;
        RECT 167.920 160.240 168.240 160.560 ;
        RECT 168.320 160.240 168.640 160.560 ;
        RECT 168.720 160.240 169.040 160.560 ;
        RECT 169.120 160.240 169.440 160.560 ;
        RECT 169.520 160.240 169.840 160.560 ;
        RECT 169.920 160.240 170.240 160.560 ;
        RECT 170.320 160.240 170.640 160.560 ;
        RECT 170.720 160.240 171.040 160.560 ;
        RECT 171.120 160.240 171.440 160.560 ;
        RECT 171.520 160.240 171.840 160.560 ;
        RECT 171.920 160.240 172.240 160.560 ;
        RECT 172.320 160.240 172.640 160.560 ;
        RECT 172.720 160.240 173.040 160.560 ;
        RECT 173.120 160.240 173.440 160.560 ;
        RECT 173.520 160.240 173.840 160.560 ;
        RECT 173.920 160.240 174.240 160.560 ;
        RECT 174.320 160.240 174.640 160.560 ;
        RECT 174.720 160.240 175.040 160.560 ;
        RECT 175.120 160.240 175.440 160.560 ;
        RECT 175.520 160.240 175.840 160.560 ;
        RECT 175.920 160.240 176.240 160.560 ;
        RECT 176.320 160.240 176.640 160.560 ;
        RECT 176.720 160.240 177.040 160.560 ;
        RECT 177.120 160.240 177.440 160.560 ;
        RECT 177.520 160.240 177.840 160.560 ;
        RECT 177.920 160.240 178.240 160.560 ;
        RECT 178.320 160.240 178.640 160.560 ;
        RECT 178.720 160.240 179.040 160.560 ;
        RECT 179.120 160.240 179.440 160.560 ;
        RECT 179.520 160.240 179.840 160.560 ;
        RECT 179.920 160.240 180.240 160.560 ;
        RECT 180.320 160.240 180.640 160.560 ;
        RECT 25.040 44.640 25.360 44.960 ;
        RECT 25.440 44.640 25.760 44.960 ;
        RECT 25.840 44.640 26.160 44.960 ;
        RECT 26.240 44.640 26.560 44.960 ;
        RECT 26.640 44.640 26.960 44.960 ;
        RECT 27.040 44.640 27.360 44.960 ;
        RECT 27.440 44.640 27.760 44.960 ;
        RECT 27.840 44.640 28.160 44.960 ;
        RECT 28.240 44.640 28.560 44.960 ;
        RECT 28.640 44.640 28.960 44.960 ;
        RECT 29.040 44.640 29.360 44.960 ;
        RECT 29.440 44.640 29.760 44.960 ;
        RECT 29.840 44.640 30.160 44.960 ;
        RECT 30.240 44.640 30.560 44.960 ;
        RECT 30.640 44.640 30.960 44.960 ;
        RECT 31.040 44.640 31.360 44.960 ;
        RECT 31.440 44.640 31.760 44.960 ;
        RECT 31.840 44.640 32.160 44.960 ;
        RECT 32.240 44.640 32.560 44.960 ;
        RECT 32.640 44.640 32.960 44.960 ;
        RECT 33.040 44.640 33.360 44.960 ;
        RECT 33.440 44.640 33.760 44.960 ;
        RECT 33.840 44.640 34.160 44.960 ;
        RECT 34.240 44.640 34.560 44.960 ;
        RECT 34.640 44.640 34.960 44.960 ;
        RECT 35.040 44.640 35.360 44.960 ;
        RECT 35.440 44.640 35.760 44.960 ;
        RECT 35.840 44.640 36.160 44.960 ;
        RECT 36.240 44.640 36.560 44.960 ;
        RECT 36.640 44.640 36.960 44.960 ;
        RECT 37.040 44.640 37.360 44.960 ;
        RECT 37.440 44.640 37.760 44.960 ;
        RECT 37.840 44.640 38.160 44.960 ;
        RECT 38.240 44.640 38.560 44.960 ;
        RECT 38.640 44.640 38.960 44.960 ;
        RECT 39.040 44.640 39.360 44.960 ;
        RECT 39.440 44.640 39.760 44.960 ;
        RECT 39.840 44.640 40.160 44.960 ;
        RECT 40.240 44.640 40.560 44.960 ;
        RECT 40.640 44.640 40.960 44.960 ;
        RECT 41.040 44.640 41.360 44.960 ;
        RECT 41.440 44.640 41.760 44.960 ;
        RECT 41.840 44.640 42.160 44.960 ;
        RECT 42.240 44.640 42.560 44.960 ;
        RECT 42.640 44.640 42.960 44.960 ;
        RECT 43.040 44.640 43.360 44.960 ;
        RECT 43.440 44.640 43.760 44.960 ;
        RECT 43.840 44.640 44.160 44.960 ;
        RECT 44.240 44.640 44.560 44.960 ;
        RECT 44.640 44.640 44.960 44.960 ;
        RECT 70.560 44.640 70.880 44.960 ;
        RECT 70.960 44.640 71.280 44.960 ;
        RECT 71.360 44.640 71.680 44.960 ;
        RECT 71.760 44.640 72.080 44.960 ;
        RECT 120.560 44.640 120.880 44.960 ;
        RECT 120.960 44.640 121.280 44.960 ;
        RECT 121.360 44.640 121.680 44.960 ;
        RECT 121.760 44.640 122.080 44.960 ;
        RECT 160.720 44.640 161.040 44.960 ;
        RECT 161.120 44.640 161.440 44.960 ;
        RECT 161.520 44.640 161.840 44.960 ;
        RECT 161.920 44.640 162.240 44.960 ;
        RECT 162.320 44.640 162.640 44.960 ;
        RECT 162.720 44.640 163.040 44.960 ;
        RECT 163.120 44.640 163.440 44.960 ;
        RECT 163.520 44.640 163.840 44.960 ;
        RECT 163.920 44.640 164.240 44.960 ;
        RECT 164.320 44.640 164.640 44.960 ;
        RECT 164.720 44.640 165.040 44.960 ;
        RECT 165.120 44.640 165.440 44.960 ;
        RECT 165.520 44.640 165.840 44.960 ;
        RECT 165.920 44.640 166.240 44.960 ;
        RECT 166.320 44.640 166.640 44.960 ;
        RECT 166.720 44.640 167.040 44.960 ;
        RECT 167.120 44.640 167.440 44.960 ;
        RECT 167.520 44.640 167.840 44.960 ;
        RECT 167.920 44.640 168.240 44.960 ;
        RECT 168.320 44.640 168.640 44.960 ;
        RECT 168.720 44.640 169.040 44.960 ;
        RECT 169.120 44.640 169.440 44.960 ;
        RECT 169.520 44.640 169.840 44.960 ;
        RECT 169.920 44.640 170.240 44.960 ;
        RECT 170.320 44.640 170.640 44.960 ;
        RECT 170.720 44.640 171.040 44.960 ;
        RECT 171.120 44.640 171.440 44.960 ;
        RECT 171.520 44.640 171.840 44.960 ;
        RECT 171.920 44.640 172.240 44.960 ;
        RECT 172.320 44.640 172.640 44.960 ;
        RECT 172.720 44.640 173.040 44.960 ;
        RECT 173.120 44.640 173.440 44.960 ;
        RECT 173.520 44.640 173.840 44.960 ;
        RECT 173.920 44.640 174.240 44.960 ;
        RECT 174.320 44.640 174.640 44.960 ;
        RECT 174.720 44.640 175.040 44.960 ;
        RECT 175.120 44.640 175.440 44.960 ;
        RECT 175.520 44.640 175.840 44.960 ;
        RECT 175.920 44.640 176.240 44.960 ;
        RECT 176.320 44.640 176.640 44.960 ;
        RECT 176.720 44.640 177.040 44.960 ;
        RECT 177.120 44.640 177.440 44.960 ;
        RECT 177.520 44.640 177.840 44.960 ;
        RECT 177.920 44.640 178.240 44.960 ;
        RECT 178.320 44.640 178.640 44.960 ;
        RECT 178.720 44.640 179.040 44.960 ;
        RECT 179.120 44.640 179.440 44.960 ;
        RECT 179.520 44.640 179.840 44.960 ;
        RECT 179.920 44.640 180.240 44.960 ;
        RECT 180.320 44.640 180.640 44.960 ;
        RECT 25.040 44.240 25.360 44.560 ;
        RECT 25.440 44.240 25.760 44.560 ;
        RECT 25.840 44.240 26.160 44.560 ;
        RECT 26.240 44.240 26.560 44.560 ;
        RECT 26.640 44.240 26.960 44.560 ;
        RECT 27.040 44.240 27.360 44.560 ;
        RECT 27.440 44.240 27.760 44.560 ;
        RECT 27.840 44.240 28.160 44.560 ;
        RECT 28.240 44.240 28.560 44.560 ;
        RECT 28.640 44.240 28.960 44.560 ;
        RECT 29.040 44.240 29.360 44.560 ;
        RECT 29.440 44.240 29.760 44.560 ;
        RECT 29.840 44.240 30.160 44.560 ;
        RECT 30.240 44.240 30.560 44.560 ;
        RECT 30.640 44.240 30.960 44.560 ;
        RECT 31.040 44.240 31.360 44.560 ;
        RECT 31.440 44.240 31.760 44.560 ;
        RECT 31.840 44.240 32.160 44.560 ;
        RECT 32.240 44.240 32.560 44.560 ;
        RECT 32.640 44.240 32.960 44.560 ;
        RECT 33.040 44.240 33.360 44.560 ;
        RECT 33.440 44.240 33.760 44.560 ;
        RECT 33.840 44.240 34.160 44.560 ;
        RECT 34.240 44.240 34.560 44.560 ;
        RECT 34.640 44.240 34.960 44.560 ;
        RECT 35.040 44.240 35.360 44.560 ;
        RECT 35.440 44.240 35.760 44.560 ;
        RECT 35.840 44.240 36.160 44.560 ;
        RECT 36.240 44.240 36.560 44.560 ;
        RECT 36.640 44.240 36.960 44.560 ;
        RECT 37.040 44.240 37.360 44.560 ;
        RECT 37.440 44.240 37.760 44.560 ;
        RECT 37.840 44.240 38.160 44.560 ;
        RECT 38.240 44.240 38.560 44.560 ;
        RECT 38.640 44.240 38.960 44.560 ;
        RECT 39.040 44.240 39.360 44.560 ;
        RECT 39.440 44.240 39.760 44.560 ;
        RECT 39.840 44.240 40.160 44.560 ;
        RECT 40.240 44.240 40.560 44.560 ;
        RECT 40.640 44.240 40.960 44.560 ;
        RECT 41.040 44.240 41.360 44.560 ;
        RECT 41.440 44.240 41.760 44.560 ;
        RECT 41.840 44.240 42.160 44.560 ;
        RECT 42.240 44.240 42.560 44.560 ;
        RECT 42.640 44.240 42.960 44.560 ;
        RECT 43.040 44.240 43.360 44.560 ;
        RECT 43.440 44.240 43.760 44.560 ;
        RECT 43.840 44.240 44.160 44.560 ;
        RECT 44.240 44.240 44.560 44.560 ;
        RECT 44.640 44.240 44.960 44.560 ;
        RECT 70.560 44.240 70.880 44.560 ;
        RECT 70.960 44.240 71.280 44.560 ;
        RECT 71.360 44.240 71.680 44.560 ;
        RECT 71.760 44.240 72.080 44.560 ;
        RECT 120.560 44.240 120.880 44.560 ;
        RECT 120.960 44.240 121.280 44.560 ;
        RECT 121.360 44.240 121.680 44.560 ;
        RECT 121.760 44.240 122.080 44.560 ;
        RECT 160.720 44.240 161.040 44.560 ;
        RECT 161.120 44.240 161.440 44.560 ;
        RECT 161.520 44.240 161.840 44.560 ;
        RECT 161.920 44.240 162.240 44.560 ;
        RECT 162.320 44.240 162.640 44.560 ;
        RECT 162.720 44.240 163.040 44.560 ;
        RECT 163.120 44.240 163.440 44.560 ;
        RECT 163.520 44.240 163.840 44.560 ;
        RECT 163.920 44.240 164.240 44.560 ;
        RECT 164.320 44.240 164.640 44.560 ;
        RECT 164.720 44.240 165.040 44.560 ;
        RECT 165.120 44.240 165.440 44.560 ;
        RECT 165.520 44.240 165.840 44.560 ;
        RECT 165.920 44.240 166.240 44.560 ;
        RECT 166.320 44.240 166.640 44.560 ;
        RECT 166.720 44.240 167.040 44.560 ;
        RECT 167.120 44.240 167.440 44.560 ;
        RECT 167.520 44.240 167.840 44.560 ;
        RECT 167.920 44.240 168.240 44.560 ;
        RECT 168.320 44.240 168.640 44.560 ;
        RECT 168.720 44.240 169.040 44.560 ;
        RECT 169.120 44.240 169.440 44.560 ;
        RECT 169.520 44.240 169.840 44.560 ;
        RECT 169.920 44.240 170.240 44.560 ;
        RECT 170.320 44.240 170.640 44.560 ;
        RECT 170.720 44.240 171.040 44.560 ;
        RECT 171.120 44.240 171.440 44.560 ;
        RECT 171.520 44.240 171.840 44.560 ;
        RECT 171.920 44.240 172.240 44.560 ;
        RECT 172.320 44.240 172.640 44.560 ;
        RECT 172.720 44.240 173.040 44.560 ;
        RECT 173.120 44.240 173.440 44.560 ;
        RECT 173.520 44.240 173.840 44.560 ;
        RECT 173.920 44.240 174.240 44.560 ;
        RECT 174.320 44.240 174.640 44.560 ;
        RECT 174.720 44.240 175.040 44.560 ;
        RECT 175.120 44.240 175.440 44.560 ;
        RECT 175.520 44.240 175.840 44.560 ;
        RECT 175.920 44.240 176.240 44.560 ;
        RECT 176.320 44.240 176.640 44.560 ;
        RECT 176.720 44.240 177.040 44.560 ;
        RECT 177.120 44.240 177.440 44.560 ;
        RECT 177.520 44.240 177.840 44.560 ;
        RECT 177.920 44.240 178.240 44.560 ;
        RECT 178.320 44.240 178.640 44.560 ;
        RECT 178.720 44.240 179.040 44.560 ;
        RECT 179.120 44.240 179.440 44.560 ;
        RECT 179.520 44.240 179.840 44.560 ;
        RECT 179.920 44.240 180.240 44.560 ;
        RECT 180.320 44.240 180.640 44.560 ;
        RECT 25.040 43.840 25.360 44.160 ;
        RECT 25.440 43.840 25.760 44.160 ;
        RECT 25.840 43.840 26.160 44.160 ;
        RECT 26.240 43.840 26.560 44.160 ;
        RECT 26.640 43.840 26.960 44.160 ;
        RECT 27.040 43.840 27.360 44.160 ;
        RECT 27.440 43.840 27.760 44.160 ;
        RECT 27.840 43.840 28.160 44.160 ;
        RECT 28.240 43.840 28.560 44.160 ;
        RECT 28.640 43.840 28.960 44.160 ;
        RECT 29.040 43.840 29.360 44.160 ;
        RECT 29.440 43.840 29.760 44.160 ;
        RECT 29.840 43.840 30.160 44.160 ;
        RECT 30.240 43.840 30.560 44.160 ;
        RECT 30.640 43.840 30.960 44.160 ;
        RECT 31.040 43.840 31.360 44.160 ;
        RECT 31.440 43.840 31.760 44.160 ;
        RECT 31.840 43.840 32.160 44.160 ;
        RECT 32.240 43.840 32.560 44.160 ;
        RECT 32.640 43.840 32.960 44.160 ;
        RECT 33.040 43.840 33.360 44.160 ;
        RECT 33.440 43.840 33.760 44.160 ;
        RECT 33.840 43.840 34.160 44.160 ;
        RECT 34.240 43.840 34.560 44.160 ;
        RECT 34.640 43.840 34.960 44.160 ;
        RECT 35.040 43.840 35.360 44.160 ;
        RECT 35.440 43.840 35.760 44.160 ;
        RECT 35.840 43.840 36.160 44.160 ;
        RECT 36.240 43.840 36.560 44.160 ;
        RECT 36.640 43.840 36.960 44.160 ;
        RECT 37.040 43.840 37.360 44.160 ;
        RECT 37.440 43.840 37.760 44.160 ;
        RECT 37.840 43.840 38.160 44.160 ;
        RECT 38.240 43.840 38.560 44.160 ;
        RECT 38.640 43.840 38.960 44.160 ;
        RECT 39.040 43.840 39.360 44.160 ;
        RECT 39.440 43.840 39.760 44.160 ;
        RECT 39.840 43.840 40.160 44.160 ;
        RECT 40.240 43.840 40.560 44.160 ;
        RECT 40.640 43.840 40.960 44.160 ;
        RECT 41.040 43.840 41.360 44.160 ;
        RECT 41.440 43.840 41.760 44.160 ;
        RECT 41.840 43.840 42.160 44.160 ;
        RECT 42.240 43.840 42.560 44.160 ;
        RECT 42.640 43.840 42.960 44.160 ;
        RECT 43.040 43.840 43.360 44.160 ;
        RECT 43.440 43.840 43.760 44.160 ;
        RECT 43.840 43.840 44.160 44.160 ;
        RECT 44.240 43.840 44.560 44.160 ;
        RECT 44.640 43.840 44.960 44.160 ;
        RECT 70.560 43.840 70.880 44.160 ;
        RECT 70.960 43.840 71.280 44.160 ;
        RECT 71.360 43.840 71.680 44.160 ;
        RECT 71.760 43.840 72.080 44.160 ;
        RECT 120.560 43.840 120.880 44.160 ;
        RECT 120.960 43.840 121.280 44.160 ;
        RECT 121.360 43.840 121.680 44.160 ;
        RECT 121.760 43.840 122.080 44.160 ;
        RECT 160.720 43.840 161.040 44.160 ;
        RECT 161.120 43.840 161.440 44.160 ;
        RECT 161.520 43.840 161.840 44.160 ;
        RECT 161.920 43.840 162.240 44.160 ;
        RECT 162.320 43.840 162.640 44.160 ;
        RECT 162.720 43.840 163.040 44.160 ;
        RECT 163.120 43.840 163.440 44.160 ;
        RECT 163.520 43.840 163.840 44.160 ;
        RECT 163.920 43.840 164.240 44.160 ;
        RECT 164.320 43.840 164.640 44.160 ;
        RECT 164.720 43.840 165.040 44.160 ;
        RECT 165.120 43.840 165.440 44.160 ;
        RECT 165.520 43.840 165.840 44.160 ;
        RECT 165.920 43.840 166.240 44.160 ;
        RECT 166.320 43.840 166.640 44.160 ;
        RECT 166.720 43.840 167.040 44.160 ;
        RECT 167.120 43.840 167.440 44.160 ;
        RECT 167.520 43.840 167.840 44.160 ;
        RECT 167.920 43.840 168.240 44.160 ;
        RECT 168.320 43.840 168.640 44.160 ;
        RECT 168.720 43.840 169.040 44.160 ;
        RECT 169.120 43.840 169.440 44.160 ;
        RECT 169.520 43.840 169.840 44.160 ;
        RECT 169.920 43.840 170.240 44.160 ;
        RECT 170.320 43.840 170.640 44.160 ;
        RECT 170.720 43.840 171.040 44.160 ;
        RECT 171.120 43.840 171.440 44.160 ;
        RECT 171.520 43.840 171.840 44.160 ;
        RECT 171.920 43.840 172.240 44.160 ;
        RECT 172.320 43.840 172.640 44.160 ;
        RECT 172.720 43.840 173.040 44.160 ;
        RECT 173.120 43.840 173.440 44.160 ;
        RECT 173.520 43.840 173.840 44.160 ;
        RECT 173.920 43.840 174.240 44.160 ;
        RECT 174.320 43.840 174.640 44.160 ;
        RECT 174.720 43.840 175.040 44.160 ;
        RECT 175.120 43.840 175.440 44.160 ;
        RECT 175.520 43.840 175.840 44.160 ;
        RECT 175.920 43.840 176.240 44.160 ;
        RECT 176.320 43.840 176.640 44.160 ;
        RECT 176.720 43.840 177.040 44.160 ;
        RECT 177.120 43.840 177.440 44.160 ;
        RECT 177.520 43.840 177.840 44.160 ;
        RECT 177.920 43.840 178.240 44.160 ;
        RECT 178.320 43.840 178.640 44.160 ;
        RECT 178.720 43.840 179.040 44.160 ;
        RECT 179.120 43.840 179.440 44.160 ;
        RECT 179.520 43.840 179.840 44.160 ;
        RECT 179.920 43.840 180.240 44.160 ;
        RECT 180.320 43.840 180.640 44.160 ;
        RECT 25.040 43.440 25.360 43.760 ;
        RECT 25.440 43.440 25.760 43.760 ;
        RECT 25.840 43.440 26.160 43.760 ;
        RECT 26.240 43.440 26.560 43.760 ;
        RECT 26.640 43.440 26.960 43.760 ;
        RECT 27.040 43.440 27.360 43.760 ;
        RECT 27.440 43.440 27.760 43.760 ;
        RECT 27.840 43.440 28.160 43.760 ;
        RECT 28.240 43.440 28.560 43.760 ;
        RECT 28.640 43.440 28.960 43.760 ;
        RECT 29.040 43.440 29.360 43.760 ;
        RECT 29.440 43.440 29.760 43.760 ;
        RECT 29.840 43.440 30.160 43.760 ;
        RECT 30.240 43.440 30.560 43.760 ;
        RECT 30.640 43.440 30.960 43.760 ;
        RECT 31.040 43.440 31.360 43.760 ;
        RECT 31.440 43.440 31.760 43.760 ;
        RECT 31.840 43.440 32.160 43.760 ;
        RECT 32.240 43.440 32.560 43.760 ;
        RECT 32.640 43.440 32.960 43.760 ;
        RECT 33.040 43.440 33.360 43.760 ;
        RECT 33.440 43.440 33.760 43.760 ;
        RECT 33.840 43.440 34.160 43.760 ;
        RECT 34.240 43.440 34.560 43.760 ;
        RECT 34.640 43.440 34.960 43.760 ;
        RECT 35.040 43.440 35.360 43.760 ;
        RECT 35.440 43.440 35.760 43.760 ;
        RECT 35.840 43.440 36.160 43.760 ;
        RECT 36.240 43.440 36.560 43.760 ;
        RECT 36.640 43.440 36.960 43.760 ;
        RECT 37.040 43.440 37.360 43.760 ;
        RECT 37.440 43.440 37.760 43.760 ;
        RECT 37.840 43.440 38.160 43.760 ;
        RECT 38.240 43.440 38.560 43.760 ;
        RECT 38.640 43.440 38.960 43.760 ;
        RECT 39.040 43.440 39.360 43.760 ;
        RECT 39.440 43.440 39.760 43.760 ;
        RECT 39.840 43.440 40.160 43.760 ;
        RECT 40.240 43.440 40.560 43.760 ;
        RECT 40.640 43.440 40.960 43.760 ;
        RECT 41.040 43.440 41.360 43.760 ;
        RECT 41.440 43.440 41.760 43.760 ;
        RECT 41.840 43.440 42.160 43.760 ;
        RECT 42.240 43.440 42.560 43.760 ;
        RECT 42.640 43.440 42.960 43.760 ;
        RECT 43.040 43.440 43.360 43.760 ;
        RECT 43.440 43.440 43.760 43.760 ;
        RECT 43.840 43.440 44.160 43.760 ;
        RECT 44.240 43.440 44.560 43.760 ;
        RECT 44.640 43.440 44.960 43.760 ;
        RECT 70.560 43.440 70.880 43.760 ;
        RECT 70.960 43.440 71.280 43.760 ;
        RECT 71.360 43.440 71.680 43.760 ;
        RECT 71.760 43.440 72.080 43.760 ;
        RECT 120.560 43.440 120.880 43.760 ;
        RECT 120.960 43.440 121.280 43.760 ;
        RECT 121.360 43.440 121.680 43.760 ;
        RECT 121.760 43.440 122.080 43.760 ;
        RECT 160.720 43.440 161.040 43.760 ;
        RECT 161.120 43.440 161.440 43.760 ;
        RECT 161.520 43.440 161.840 43.760 ;
        RECT 161.920 43.440 162.240 43.760 ;
        RECT 162.320 43.440 162.640 43.760 ;
        RECT 162.720 43.440 163.040 43.760 ;
        RECT 163.120 43.440 163.440 43.760 ;
        RECT 163.520 43.440 163.840 43.760 ;
        RECT 163.920 43.440 164.240 43.760 ;
        RECT 164.320 43.440 164.640 43.760 ;
        RECT 164.720 43.440 165.040 43.760 ;
        RECT 165.120 43.440 165.440 43.760 ;
        RECT 165.520 43.440 165.840 43.760 ;
        RECT 165.920 43.440 166.240 43.760 ;
        RECT 166.320 43.440 166.640 43.760 ;
        RECT 166.720 43.440 167.040 43.760 ;
        RECT 167.120 43.440 167.440 43.760 ;
        RECT 167.520 43.440 167.840 43.760 ;
        RECT 167.920 43.440 168.240 43.760 ;
        RECT 168.320 43.440 168.640 43.760 ;
        RECT 168.720 43.440 169.040 43.760 ;
        RECT 169.120 43.440 169.440 43.760 ;
        RECT 169.520 43.440 169.840 43.760 ;
        RECT 169.920 43.440 170.240 43.760 ;
        RECT 170.320 43.440 170.640 43.760 ;
        RECT 170.720 43.440 171.040 43.760 ;
        RECT 171.120 43.440 171.440 43.760 ;
        RECT 171.520 43.440 171.840 43.760 ;
        RECT 171.920 43.440 172.240 43.760 ;
        RECT 172.320 43.440 172.640 43.760 ;
        RECT 172.720 43.440 173.040 43.760 ;
        RECT 173.120 43.440 173.440 43.760 ;
        RECT 173.520 43.440 173.840 43.760 ;
        RECT 173.920 43.440 174.240 43.760 ;
        RECT 174.320 43.440 174.640 43.760 ;
        RECT 174.720 43.440 175.040 43.760 ;
        RECT 175.120 43.440 175.440 43.760 ;
        RECT 175.520 43.440 175.840 43.760 ;
        RECT 175.920 43.440 176.240 43.760 ;
        RECT 176.320 43.440 176.640 43.760 ;
        RECT 176.720 43.440 177.040 43.760 ;
        RECT 177.120 43.440 177.440 43.760 ;
        RECT 177.520 43.440 177.840 43.760 ;
        RECT 177.920 43.440 178.240 43.760 ;
        RECT 178.320 43.440 178.640 43.760 ;
        RECT 178.720 43.440 179.040 43.760 ;
        RECT 179.120 43.440 179.440 43.760 ;
        RECT 179.520 43.440 179.840 43.760 ;
        RECT 179.920 43.440 180.240 43.760 ;
        RECT 180.320 43.440 180.640 43.760 ;
        RECT 25.040 43.040 25.360 43.360 ;
        RECT 25.440 43.040 25.760 43.360 ;
        RECT 25.840 43.040 26.160 43.360 ;
        RECT 26.240 43.040 26.560 43.360 ;
        RECT 26.640 43.040 26.960 43.360 ;
        RECT 27.040 43.040 27.360 43.360 ;
        RECT 27.440 43.040 27.760 43.360 ;
        RECT 27.840 43.040 28.160 43.360 ;
        RECT 28.240 43.040 28.560 43.360 ;
        RECT 28.640 43.040 28.960 43.360 ;
        RECT 29.040 43.040 29.360 43.360 ;
        RECT 29.440 43.040 29.760 43.360 ;
        RECT 29.840 43.040 30.160 43.360 ;
        RECT 30.240 43.040 30.560 43.360 ;
        RECT 30.640 43.040 30.960 43.360 ;
        RECT 31.040 43.040 31.360 43.360 ;
        RECT 31.440 43.040 31.760 43.360 ;
        RECT 31.840 43.040 32.160 43.360 ;
        RECT 32.240 43.040 32.560 43.360 ;
        RECT 32.640 43.040 32.960 43.360 ;
        RECT 33.040 43.040 33.360 43.360 ;
        RECT 33.440 43.040 33.760 43.360 ;
        RECT 33.840 43.040 34.160 43.360 ;
        RECT 34.240 43.040 34.560 43.360 ;
        RECT 34.640 43.040 34.960 43.360 ;
        RECT 35.040 43.040 35.360 43.360 ;
        RECT 35.440 43.040 35.760 43.360 ;
        RECT 35.840 43.040 36.160 43.360 ;
        RECT 36.240 43.040 36.560 43.360 ;
        RECT 36.640 43.040 36.960 43.360 ;
        RECT 37.040 43.040 37.360 43.360 ;
        RECT 37.440 43.040 37.760 43.360 ;
        RECT 37.840 43.040 38.160 43.360 ;
        RECT 38.240 43.040 38.560 43.360 ;
        RECT 38.640 43.040 38.960 43.360 ;
        RECT 39.040 43.040 39.360 43.360 ;
        RECT 39.440 43.040 39.760 43.360 ;
        RECT 39.840 43.040 40.160 43.360 ;
        RECT 40.240 43.040 40.560 43.360 ;
        RECT 40.640 43.040 40.960 43.360 ;
        RECT 41.040 43.040 41.360 43.360 ;
        RECT 41.440 43.040 41.760 43.360 ;
        RECT 41.840 43.040 42.160 43.360 ;
        RECT 42.240 43.040 42.560 43.360 ;
        RECT 42.640 43.040 42.960 43.360 ;
        RECT 43.040 43.040 43.360 43.360 ;
        RECT 43.440 43.040 43.760 43.360 ;
        RECT 43.840 43.040 44.160 43.360 ;
        RECT 44.240 43.040 44.560 43.360 ;
        RECT 44.640 43.040 44.960 43.360 ;
        RECT 70.560 43.040 70.880 43.360 ;
        RECT 70.960 43.040 71.280 43.360 ;
        RECT 71.360 43.040 71.680 43.360 ;
        RECT 71.760 43.040 72.080 43.360 ;
        RECT 120.560 43.040 120.880 43.360 ;
        RECT 120.960 43.040 121.280 43.360 ;
        RECT 121.360 43.040 121.680 43.360 ;
        RECT 121.760 43.040 122.080 43.360 ;
        RECT 160.720 43.040 161.040 43.360 ;
        RECT 161.120 43.040 161.440 43.360 ;
        RECT 161.520 43.040 161.840 43.360 ;
        RECT 161.920 43.040 162.240 43.360 ;
        RECT 162.320 43.040 162.640 43.360 ;
        RECT 162.720 43.040 163.040 43.360 ;
        RECT 163.120 43.040 163.440 43.360 ;
        RECT 163.520 43.040 163.840 43.360 ;
        RECT 163.920 43.040 164.240 43.360 ;
        RECT 164.320 43.040 164.640 43.360 ;
        RECT 164.720 43.040 165.040 43.360 ;
        RECT 165.120 43.040 165.440 43.360 ;
        RECT 165.520 43.040 165.840 43.360 ;
        RECT 165.920 43.040 166.240 43.360 ;
        RECT 166.320 43.040 166.640 43.360 ;
        RECT 166.720 43.040 167.040 43.360 ;
        RECT 167.120 43.040 167.440 43.360 ;
        RECT 167.520 43.040 167.840 43.360 ;
        RECT 167.920 43.040 168.240 43.360 ;
        RECT 168.320 43.040 168.640 43.360 ;
        RECT 168.720 43.040 169.040 43.360 ;
        RECT 169.120 43.040 169.440 43.360 ;
        RECT 169.520 43.040 169.840 43.360 ;
        RECT 169.920 43.040 170.240 43.360 ;
        RECT 170.320 43.040 170.640 43.360 ;
        RECT 170.720 43.040 171.040 43.360 ;
        RECT 171.120 43.040 171.440 43.360 ;
        RECT 171.520 43.040 171.840 43.360 ;
        RECT 171.920 43.040 172.240 43.360 ;
        RECT 172.320 43.040 172.640 43.360 ;
        RECT 172.720 43.040 173.040 43.360 ;
        RECT 173.120 43.040 173.440 43.360 ;
        RECT 173.520 43.040 173.840 43.360 ;
        RECT 173.920 43.040 174.240 43.360 ;
        RECT 174.320 43.040 174.640 43.360 ;
        RECT 174.720 43.040 175.040 43.360 ;
        RECT 175.120 43.040 175.440 43.360 ;
        RECT 175.520 43.040 175.840 43.360 ;
        RECT 175.920 43.040 176.240 43.360 ;
        RECT 176.320 43.040 176.640 43.360 ;
        RECT 176.720 43.040 177.040 43.360 ;
        RECT 177.120 43.040 177.440 43.360 ;
        RECT 177.520 43.040 177.840 43.360 ;
        RECT 177.920 43.040 178.240 43.360 ;
        RECT 178.320 43.040 178.640 43.360 ;
        RECT 178.720 43.040 179.040 43.360 ;
        RECT 179.120 43.040 179.440 43.360 ;
        RECT 179.520 43.040 179.840 43.360 ;
        RECT 179.920 43.040 180.240 43.360 ;
        RECT 180.320 43.040 180.640 43.360 ;
        RECT 25.040 42.640 25.360 42.960 ;
        RECT 25.440 42.640 25.760 42.960 ;
        RECT 25.840 42.640 26.160 42.960 ;
        RECT 26.240 42.640 26.560 42.960 ;
        RECT 26.640 42.640 26.960 42.960 ;
        RECT 27.040 42.640 27.360 42.960 ;
        RECT 27.440 42.640 27.760 42.960 ;
        RECT 27.840 42.640 28.160 42.960 ;
        RECT 28.240 42.640 28.560 42.960 ;
        RECT 28.640 42.640 28.960 42.960 ;
        RECT 29.040 42.640 29.360 42.960 ;
        RECT 29.440 42.640 29.760 42.960 ;
        RECT 29.840 42.640 30.160 42.960 ;
        RECT 30.240 42.640 30.560 42.960 ;
        RECT 30.640 42.640 30.960 42.960 ;
        RECT 31.040 42.640 31.360 42.960 ;
        RECT 31.440 42.640 31.760 42.960 ;
        RECT 31.840 42.640 32.160 42.960 ;
        RECT 32.240 42.640 32.560 42.960 ;
        RECT 32.640 42.640 32.960 42.960 ;
        RECT 33.040 42.640 33.360 42.960 ;
        RECT 33.440 42.640 33.760 42.960 ;
        RECT 33.840 42.640 34.160 42.960 ;
        RECT 34.240 42.640 34.560 42.960 ;
        RECT 34.640 42.640 34.960 42.960 ;
        RECT 35.040 42.640 35.360 42.960 ;
        RECT 35.440 42.640 35.760 42.960 ;
        RECT 35.840 42.640 36.160 42.960 ;
        RECT 36.240 42.640 36.560 42.960 ;
        RECT 36.640 42.640 36.960 42.960 ;
        RECT 37.040 42.640 37.360 42.960 ;
        RECT 37.440 42.640 37.760 42.960 ;
        RECT 37.840 42.640 38.160 42.960 ;
        RECT 38.240 42.640 38.560 42.960 ;
        RECT 38.640 42.640 38.960 42.960 ;
        RECT 39.040 42.640 39.360 42.960 ;
        RECT 39.440 42.640 39.760 42.960 ;
        RECT 39.840 42.640 40.160 42.960 ;
        RECT 40.240 42.640 40.560 42.960 ;
        RECT 40.640 42.640 40.960 42.960 ;
        RECT 41.040 42.640 41.360 42.960 ;
        RECT 41.440 42.640 41.760 42.960 ;
        RECT 41.840 42.640 42.160 42.960 ;
        RECT 42.240 42.640 42.560 42.960 ;
        RECT 42.640 42.640 42.960 42.960 ;
        RECT 43.040 42.640 43.360 42.960 ;
        RECT 43.440 42.640 43.760 42.960 ;
        RECT 43.840 42.640 44.160 42.960 ;
        RECT 44.240 42.640 44.560 42.960 ;
        RECT 44.640 42.640 44.960 42.960 ;
        RECT 70.560 42.640 70.880 42.960 ;
        RECT 70.960 42.640 71.280 42.960 ;
        RECT 71.360 42.640 71.680 42.960 ;
        RECT 71.760 42.640 72.080 42.960 ;
        RECT 120.560 42.640 120.880 42.960 ;
        RECT 120.960 42.640 121.280 42.960 ;
        RECT 121.360 42.640 121.680 42.960 ;
        RECT 121.760 42.640 122.080 42.960 ;
        RECT 160.720 42.640 161.040 42.960 ;
        RECT 161.120 42.640 161.440 42.960 ;
        RECT 161.520 42.640 161.840 42.960 ;
        RECT 161.920 42.640 162.240 42.960 ;
        RECT 162.320 42.640 162.640 42.960 ;
        RECT 162.720 42.640 163.040 42.960 ;
        RECT 163.120 42.640 163.440 42.960 ;
        RECT 163.520 42.640 163.840 42.960 ;
        RECT 163.920 42.640 164.240 42.960 ;
        RECT 164.320 42.640 164.640 42.960 ;
        RECT 164.720 42.640 165.040 42.960 ;
        RECT 165.120 42.640 165.440 42.960 ;
        RECT 165.520 42.640 165.840 42.960 ;
        RECT 165.920 42.640 166.240 42.960 ;
        RECT 166.320 42.640 166.640 42.960 ;
        RECT 166.720 42.640 167.040 42.960 ;
        RECT 167.120 42.640 167.440 42.960 ;
        RECT 167.520 42.640 167.840 42.960 ;
        RECT 167.920 42.640 168.240 42.960 ;
        RECT 168.320 42.640 168.640 42.960 ;
        RECT 168.720 42.640 169.040 42.960 ;
        RECT 169.120 42.640 169.440 42.960 ;
        RECT 169.520 42.640 169.840 42.960 ;
        RECT 169.920 42.640 170.240 42.960 ;
        RECT 170.320 42.640 170.640 42.960 ;
        RECT 170.720 42.640 171.040 42.960 ;
        RECT 171.120 42.640 171.440 42.960 ;
        RECT 171.520 42.640 171.840 42.960 ;
        RECT 171.920 42.640 172.240 42.960 ;
        RECT 172.320 42.640 172.640 42.960 ;
        RECT 172.720 42.640 173.040 42.960 ;
        RECT 173.120 42.640 173.440 42.960 ;
        RECT 173.520 42.640 173.840 42.960 ;
        RECT 173.920 42.640 174.240 42.960 ;
        RECT 174.320 42.640 174.640 42.960 ;
        RECT 174.720 42.640 175.040 42.960 ;
        RECT 175.120 42.640 175.440 42.960 ;
        RECT 175.520 42.640 175.840 42.960 ;
        RECT 175.920 42.640 176.240 42.960 ;
        RECT 176.320 42.640 176.640 42.960 ;
        RECT 176.720 42.640 177.040 42.960 ;
        RECT 177.120 42.640 177.440 42.960 ;
        RECT 177.520 42.640 177.840 42.960 ;
        RECT 177.920 42.640 178.240 42.960 ;
        RECT 178.320 42.640 178.640 42.960 ;
        RECT 178.720 42.640 179.040 42.960 ;
        RECT 179.120 42.640 179.440 42.960 ;
        RECT 179.520 42.640 179.840 42.960 ;
        RECT 179.920 42.640 180.240 42.960 ;
        RECT 180.320 42.640 180.640 42.960 ;
        RECT 25.040 42.240 25.360 42.560 ;
        RECT 25.440 42.240 25.760 42.560 ;
        RECT 25.840 42.240 26.160 42.560 ;
        RECT 26.240 42.240 26.560 42.560 ;
        RECT 26.640 42.240 26.960 42.560 ;
        RECT 27.040 42.240 27.360 42.560 ;
        RECT 27.440 42.240 27.760 42.560 ;
        RECT 27.840 42.240 28.160 42.560 ;
        RECT 28.240 42.240 28.560 42.560 ;
        RECT 28.640 42.240 28.960 42.560 ;
        RECT 29.040 42.240 29.360 42.560 ;
        RECT 29.440 42.240 29.760 42.560 ;
        RECT 29.840 42.240 30.160 42.560 ;
        RECT 30.240 42.240 30.560 42.560 ;
        RECT 30.640 42.240 30.960 42.560 ;
        RECT 31.040 42.240 31.360 42.560 ;
        RECT 31.440 42.240 31.760 42.560 ;
        RECT 31.840 42.240 32.160 42.560 ;
        RECT 32.240 42.240 32.560 42.560 ;
        RECT 32.640 42.240 32.960 42.560 ;
        RECT 33.040 42.240 33.360 42.560 ;
        RECT 33.440 42.240 33.760 42.560 ;
        RECT 33.840 42.240 34.160 42.560 ;
        RECT 34.240 42.240 34.560 42.560 ;
        RECT 34.640 42.240 34.960 42.560 ;
        RECT 35.040 42.240 35.360 42.560 ;
        RECT 35.440 42.240 35.760 42.560 ;
        RECT 35.840 42.240 36.160 42.560 ;
        RECT 36.240 42.240 36.560 42.560 ;
        RECT 36.640 42.240 36.960 42.560 ;
        RECT 37.040 42.240 37.360 42.560 ;
        RECT 37.440 42.240 37.760 42.560 ;
        RECT 37.840 42.240 38.160 42.560 ;
        RECT 38.240 42.240 38.560 42.560 ;
        RECT 38.640 42.240 38.960 42.560 ;
        RECT 39.040 42.240 39.360 42.560 ;
        RECT 39.440 42.240 39.760 42.560 ;
        RECT 39.840 42.240 40.160 42.560 ;
        RECT 40.240 42.240 40.560 42.560 ;
        RECT 40.640 42.240 40.960 42.560 ;
        RECT 41.040 42.240 41.360 42.560 ;
        RECT 41.440 42.240 41.760 42.560 ;
        RECT 41.840 42.240 42.160 42.560 ;
        RECT 42.240 42.240 42.560 42.560 ;
        RECT 42.640 42.240 42.960 42.560 ;
        RECT 43.040 42.240 43.360 42.560 ;
        RECT 43.440 42.240 43.760 42.560 ;
        RECT 43.840 42.240 44.160 42.560 ;
        RECT 44.240 42.240 44.560 42.560 ;
        RECT 44.640 42.240 44.960 42.560 ;
        RECT 70.560 42.240 70.880 42.560 ;
        RECT 70.960 42.240 71.280 42.560 ;
        RECT 71.360 42.240 71.680 42.560 ;
        RECT 71.760 42.240 72.080 42.560 ;
        RECT 120.560 42.240 120.880 42.560 ;
        RECT 120.960 42.240 121.280 42.560 ;
        RECT 121.360 42.240 121.680 42.560 ;
        RECT 121.760 42.240 122.080 42.560 ;
        RECT 160.720 42.240 161.040 42.560 ;
        RECT 161.120 42.240 161.440 42.560 ;
        RECT 161.520 42.240 161.840 42.560 ;
        RECT 161.920 42.240 162.240 42.560 ;
        RECT 162.320 42.240 162.640 42.560 ;
        RECT 162.720 42.240 163.040 42.560 ;
        RECT 163.120 42.240 163.440 42.560 ;
        RECT 163.520 42.240 163.840 42.560 ;
        RECT 163.920 42.240 164.240 42.560 ;
        RECT 164.320 42.240 164.640 42.560 ;
        RECT 164.720 42.240 165.040 42.560 ;
        RECT 165.120 42.240 165.440 42.560 ;
        RECT 165.520 42.240 165.840 42.560 ;
        RECT 165.920 42.240 166.240 42.560 ;
        RECT 166.320 42.240 166.640 42.560 ;
        RECT 166.720 42.240 167.040 42.560 ;
        RECT 167.120 42.240 167.440 42.560 ;
        RECT 167.520 42.240 167.840 42.560 ;
        RECT 167.920 42.240 168.240 42.560 ;
        RECT 168.320 42.240 168.640 42.560 ;
        RECT 168.720 42.240 169.040 42.560 ;
        RECT 169.120 42.240 169.440 42.560 ;
        RECT 169.520 42.240 169.840 42.560 ;
        RECT 169.920 42.240 170.240 42.560 ;
        RECT 170.320 42.240 170.640 42.560 ;
        RECT 170.720 42.240 171.040 42.560 ;
        RECT 171.120 42.240 171.440 42.560 ;
        RECT 171.520 42.240 171.840 42.560 ;
        RECT 171.920 42.240 172.240 42.560 ;
        RECT 172.320 42.240 172.640 42.560 ;
        RECT 172.720 42.240 173.040 42.560 ;
        RECT 173.120 42.240 173.440 42.560 ;
        RECT 173.520 42.240 173.840 42.560 ;
        RECT 173.920 42.240 174.240 42.560 ;
        RECT 174.320 42.240 174.640 42.560 ;
        RECT 174.720 42.240 175.040 42.560 ;
        RECT 175.120 42.240 175.440 42.560 ;
        RECT 175.520 42.240 175.840 42.560 ;
        RECT 175.920 42.240 176.240 42.560 ;
        RECT 176.320 42.240 176.640 42.560 ;
        RECT 176.720 42.240 177.040 42.560 ;
        RECT 177.120 42.240 177.440 42.560 ;
        RECT 177.520 42.240 177.840 42.560 ;
        RECT 177.920 42.240 178.240 42.560 ;
        RECT 178.320 42.240 178.640 42.560 ;
        RECT 178.720 42.240 179.040 42.560 ;
        RECT 179.120 42.240 179.440 42.560 ;
        RECT 179.520 42.240 179.840 42.560 ;
        RECT 179.920 42.240 180.240 42.560 ;
        RECT 180.320 42.240 180.640 42.560 ;
        RECT 25.040 41.840 25.360 42.160 ;
        RECT 25.440 41.840 25.760 42.160 ;
        RECT 25.840 41.840 26.160 42.160 ;
        RECT 26.240 41.840 26.560 42.160 ;
        RECT 26.640 41.840 26.960 42.160 ;
        RECT 27.040 41.840 27.360 42.160 ;
        RECT 27.440 41.840 27.760 42.160 ;
        RECT 27.840 41.840 28.160 42.160 ;
        RECT 28.240 41.840 28.560 42.160 ;
        RECT 28.640 41.840 28.960 42.160 ;
        RECT 29.040 41.840 29.360 42.160 ;
        RECT 29.440 41.840 29.760 42.160 ;
        RECT 29.840 41.840 30.160 42.160 ;
        RECT 30.240 41.840 30.560 42.160 ;
        RECT 30.640 41.840 30.960 42.160 ;
        RECT 31.040 41.840 31.360 42.160 ;
        RECT 31.440 41.840 31.760 42.160 ;
        RECT 31.840 41.840 32.160 42.160 ;
        RECT 32.240 41.840 32.560 42.160 ;
        RECT 32.640 41.840 32.960 42.160 ;
        RECT 33.040 41.840 33.360 42.160 ;
        RECT 33.440 41.840 33.760 42.160 ;
        RECT 33.840 41.840 34.160 42.160 ;
        RECT 34.240 41.840 34.560 42.160 ;
        RECT 34.640 41.840 34.960 42.160 ;
        RECT 35.040 41.840 35.360 42.160 ;
        RECT 35.440 41.840 35.760 42.160 ;
        RECT 35.840 41.840 36.160 42.160 ;
        RECT 36.240 41.840 36.560 42.160 ;
        RECT 36.640 41.840 36.960 42.160 ;
        RECT 37.040 41.840 37.360 42.160 ;
        RECT 37.440 41.840 37.760 42.160 ;
        RECT 37.840 41.840 38.160 42.160 ;
        RECT 38.240 41.840 38.560 42.160 ;
        RECT 38.640 41.840 38.960 42.160 ;
        RECT 39.040 41.840 39.360 42.160 ;
        RECT 39.440 41.840 39.760 42.160 ;
        RECT 39.840 41.840 40.160 42.160 ;
        RECT 40.240 41.840 40.560 42.160 ;
        RECT 40.640 41.840 40.960 42.160 ;
        RECT 41.040 41.840 41.360 42.160 ;
        RECT 41.440 41.840 41.760 42.160 ;
        RECT 41.840 41.840 42.160 42.160 ;
        RECT 42.240 41.840 42.560 42.160 ;
        RECT 42.640 41.840 42.960 42.160 ;
        RECT 43.040 41.840 43.360 42.160 ;
        RECT 43.440 41.840 43.760 42.160 ;
        RECT 43.840 41.840 44.160 42.160 ;
        RECT 44.240 41.840 44.560 42.160 ;
        RECT 44.640 41.840 44.960 42.160 ;
        RECT 70.560 41.840 70.880 42.160 ;
        RECT 70.960 41.840 71.280 42.160 ;
        RECT 71.360 41.840 71.680 42.160 ;
        RECT 71.760 41.840 72.080 42.160 ;
        RECT 120.560 41.840 120.880 42.160 ;
        RECT 120.960 41.840 121.280 42.160 ;
        RECT 121.360 41.840 121.680 42.160 ;
        RECT 121.760 41.840 122.080 42.160 ;
        RECT 160.720 41.840 161.040 42.160 ;
        RECT 161.120 41.840 161.440 42.160 ;
        RECT 161.520 41.840 161.840 42.160 ;
        RECT 161.920 41.840 162.240 42.160 ;
        RECT 162.320 41.840 162.640 42.160 ;
        RECT 162.720 41.840 163.040 42.160 ;
        RECT 163.120 41.840 163.440 42.160 ;
        RECT 163.520 41.840 163.840 42.160 ;
        RECT 163.920 41.840 164.240 42.160 ;
        RECT 164.320 41.840 164.640 42.160 ;
        RECT 164.720 41.840 165.040 42.160 ;
        RECT 165.120 41.840 165.440 42.160 ;
        RECT 165.520 41.840 165.840 42.160 ;
        RECT 165.920 41.840 166.240 42.160 ;
        RECT 166.320 41.840 166.640 42.160 ;
        RECT 166.720 41.840 167.040 42.160 ;
        RECT 167.120 41.840 167.440 42.160 ;
        RECT 167.520 41.840 167.840 42.160 ;
        RECT 167.920 41.840 168.240 42.160 ;
        RECT 168.320 41.840 168.640 42.160 ;
        RECT 168.720 41.840 169.040 42.160 ;
        RECT 169.120 41.840 169.440 42.160 ;
        RECT 169.520 41.840 169.840 42.160 ;
        RECT 169.920 41.840 170.240 42.160 ;
        RECT 170.320 41.840 170.640 42.160 ;
        RECT 170.720 41.840 171.040 42.160 ;
        RECT 171.120 41.840 171.440 42.160 ;
        RECT 171.520 41.840 171.840 42.160 ;
        RECT 171.920 41.840 172.240 42.160 ;
        RECT 172.320 41.840 172.640 42.160 ;
        RECT 172.720 41.840 173.040 42.160 ;
        RECT 173.120 41.840 173.440 42.160 ;
        RECT 173.520 41.840 173.840 42.160 ;
        RECT 173.920 41.840 174.240 42.160 ;
        RECT 174.320 41.840 174.640 42.160 ;
        RECT 174.720 41.840 175.040 42.160 ;
        RECT 175.120 41.840 175.440 42.160 ;
        RECT 175.520 41.840 175.840 42.160 ;
        RECT 175.920 41.840 176.240 42.160 ;
        RECT 176.320 41.840 176.640 42.160 ;
        RECT 176.720 41.840 177.040 42.160 ;
        RECT 177.120 41.840 177.440 42.160 ;
        RECT 177.520 41.840 177.840 42.160 ;
        RECT 177.920 41.840 178.240 42.160 ;
        RECT 178.320 41.840 178.640 42.160 ;
        RECT 178.720 41.840 179.040 42.160 ;
        RECT 179.120 41.840 179.440 42.160 ;
        RECT 179.520 41.840 179.840 42.160 ;
        RECT 179.920 41.840 180.240 42.160 ;
        RECT 180.320 41.840 180.640 42.160 ;
        RECT 25.040 41.440 25.360 41.760 ;
        RECT 25.440 41.440 25.760 41.760 ;
        RECT 25.840 41.440 26.160 41.760 ;
        RECT 26.240 41.440 26.560 41.760 ;
        RECT 26.640 41.440 26.960 41.760 ;
        RECT 27.040 41.440 27.360 41.760 ;
        RECT 27.440 41.440 27.760 41.760 ;
        RECT 27.840 41.440 28.160 41.760 ;
        RECT 28.240 41.440 28.560 41.760 ;
        RECT 28.640 41.440 28.960 41.760 ;
        RECT 29.040 41.440 29.360 41.760 ;
        RECT 29.440 41.440 29.760 41.760 ;
        RECT 29.840 41.440 30.160 41.760 ;
        RECT 30.240 41.440 30.560 41.760 ;
        RECT 30.640 41.440 30.960 41.760 ;
        RECT 31.040 41.440 31.360 41.760 ;
        RECT 31.440 41.440 31.760 41.760 ;
        RECT 31.840 41.440 32.160 41.760 ;
        RECT 32.240 41.440 32.560 41.760 ;
        RECT 32.640 41.440 32.960 41.760 ;
        RECT 33.040 41.440 33.360 41.760 ;
        RECT 33.440 41.440 33.760 41.760 ;
        RECT 33.840 41.440 34.160 41.760 ;
        RECT 34.240 41.440 34.560 41.760 ;
        RECT 34.640 41.440 34.960 41.760 ;
        RECT 35.040 41.440 35.360 41.760 ;
        RECT 35.440 41.440 35.760 41.760 ;
        RECT 35.840 41.440 36.160 41.760 ;
        RECT 36.240 41.440 36.560 41.760 ;
        RECT 36.640 41.440 36.960 41.760 ;
        RECT 37.040 41.440 37.360 41.760 ;
        RECT 37.440 41.440 37.760 41.760 ;
        RECT 37.840 41.440 38.160 41.760 ;
        RECT 38.240 41.440 38.560 41.760 ;
        RECT 38.640 41.440 38.960 41.760 ;
        RECT 39.040 41.440 39.360 41.760 ;
        RECT 39.440 41.440 39.760 41.760 ;
        RECT 39.840 41.440 40.160 41.760 ;
        RECT 40.240 41.440 40.560 41.760 ;
        RECT 40.640 41.440 40.960 41.760 ;
        RECT 41.040 41.440 41.360 41.760 ;
        RECT 41.440 41.440 41.760 41.760 ;
        RECT 41.840 41.440 42.160 41.760 ;
        RECT 42.240 41.440 42.560 41.760 ;
        RECT 42.640 41.440 42.960 41.760 ;
        RECT 43.040 41.440 43.360 41.760 ;
        RECT 43.440 41.440 43.760 41.760 ;
        RECT 43.840 41.440 44.160 41.760 ;
        RECT 44.240 41.440 44.560 41.760 ;
        RECT 44.640 41.440 44.960 41.760 ;
        RECT 70.560 41.440 70.880 41.760 ;
        RECT 70.960 41.440 71.280 41.760 ;
        RECT 71.360 41.440 71.680 41.760 ;
        RECT 71.760 41.440 72.080 41.760 ;
        RECT 120.560 41.440 120.880 41.760 ;
        RECT 120.960 41.440 121.280 41.760 ;
        RECT 121.360 41.440 121.680 41.760 ;
        RECT 121.760 41.440 122.080 41.760 ;
        RECT 160.720 41.440 161.040 41.760 ;
        RECT 161.120 41.440 161.440 41.760 ;
        RECT 161.520 41.440 161.840 41.760 ;
        RECT 161.920 41.440 162.240 41.760 ;
        RECT 162.320 41.440 162.640 41.760 ;
        RECT 162.720 41.440 163.040 41.760 ;
        RECT 163.120 41.440 163.440 41.760 ;
        RECT 163.520 41.440 163.840 41.760 ;
        RECT 163.920 41.440 164.240 41.760 ;
        RECT 164.320 41.440 164.640 41.760 ;
        RECT 164.720 41.440 165.040 41.760 ;
        RECT 165.120 41.440 165.440 41.760 ;
        RECT 165.520 41.440 165.840 41.760 ;
        RECT 165.920 41.440 166.240 41.760 ;
        RECT 166.320 41.440 166.640 41.760 ;
        RECT 166.720 41.440 167.040 41.760 ;
        RECT 167.120 41.440 167.440 41.760 ;
        RECT 167.520 41.440 167.840 41.760 ;
        RECT 167.920 41.440 168.240 41.760 ;
        RECT 168.320 41.440 168.640 41.760 ;
        RECT 168.720 41.440 169.040 41.760 ;
        RECT 169.120 41.440 169.440 41.760 ;
        RECT 169.520 41.440 169.840 41.760 ;
        RECT 169.920 41.440 170.240 41.760 ;
        RECT 170.320 41.440 170.640 41.760 ;
        RECT 170.720 41.440 171.040 41.760 ;
        RECT 171.120 41.440 171.440 41.760 ;
        RECT 171.520 41.440 171.840 41.760 ;
        RECT 171.920 41.440 172.240 41.760 ;
        RECT 172.320 41.440 172.640 41.760 ;
        RECT 172.720 41.440 173.040 41.760 ;
        RECT 173.120 41.440 173.440 41.760 ;
        RECT 173.520 41.440 173.840 41.760 ;
        RECT 173.920 41.440 174.240 41.760 ;
        RECT 174.320 41.440 174.640 41.760 ;
        RECT 174.720 41.440 175.040 41.760 ;
        RECT 175.120 41.440 175.440 41.760 ;
        RECT 175.520 41.440 175.840 41.760 ;
        RECT 175.920 41.440 176.240 41.760 ;
        RECT 176.320 41.440 176.640 41.760 ;
        RECT 176.720 41.440 177.040 41.760 ;
        RECT 177.120 41.440 177.440 41.760 ;
        RECT 177.520 41.440 177.840 41.760 ;
        RECT 177.920 41.440 178.240 41.760 ;
        RECT 178.320 41.440 178.640 41.760 ;
        RECT 178.720 41.440 179.040 41.760 ;
        RECT 179.120 41.440 179.440 41.760 ;
        RECT 179.520 41.440 179.840 41.760 ;
        RECT 179.920 41.440 180.240 41.760 ;
        RECT 180.320 41.440 180.640 41.760 ;
        RECT 25.040 41.040 25.360 41.360 ;
        RECT 25.440 41.040 25.760 41.360 ;
        RECT 25.840 41.040 26.160 41.360 ;
        RECT 26.240 41.040 26.560 41.360 ;
        RECT 26.640 41.040 26.960 41.360 ;
        RECT 27.040 41.040 27.360 41.360 ;
        RECT 27.440 41.040 27.760 41.360 ;
        RECT 27.840 41.040 28.160 41.360 ;
        RECT 28.240 41.040 28.560 41.360 ;
        RECT 28.640 41.040 28.960 41.360 ;
        RECT 29.040 41.040 29.360 41.360 ;
        RECT 29.440 41.040 29.760 41.360 ;
        RECT 29.840 41.040 30.160 41.360 ;
        RECT 30.240 41.040 30.560 41.360 ;
        RECT 30.640 41.040 30.960 41.360 ;
        RECT 31.040 41.040 31.360 41.360 ;
        RECT 31.440 41.040 31.760 41.360 ;
        RECT 31.840 41.040 32.160 41.360 ;
        RECT 32.240 41.040 32.560 41.360 ;
        RECT 32.640 41.040 32.960 41.360 ;
        RECT 33.040 41.040 33.360 41.360 ;
        RECT 33.440 41.040 33.760 41.360 ;
        RECT 33.840 41.040 34.160 41.360 ;
        RECT 34.240 41.040 34.560 41.360 ;
        RECT 34.640 41.040 34.960 41.360 ;
        RECT 35.040 41.040 35.360 41.360 ;
        RECT 35.440 41.040 35.760 41.360 ;
        RECT 35.840 41.040 36.160 41.360 ;
        RECT 36.240 41.040 36.560 41.360 ;
        RECT 36.640 41.040 36.960 41.360 ;
        RECT 37.040 41.040 37.360 41.360 ;
        RECT 37.440 41.040 37.760 41.360 ;
        RECT 37.840 41.040 38.160 41.360 ;
        RECT 38.240 41.040 38.560 41.360 ;
        RECT 38.640 41.040 38.960 41.360 ;
        RECT 39.040 41.040 39.360 41.360 ;
        RECT 39.440 41.040 39.760 41.360 ;
        RECT 39.840 41.040 40.160 41.360 ;
        RECT 40.240 41.040 40.560 41.360 ;
        RECT 40.640 41.040 40.960 41.360 ;
        RECT 41.040 41.040 41.360 41.360 ;
        RECT 41.440 41.040 41.760 41.360 ;
        RECT 41.840 41.040 42.160 41.360 ;
        RECT 42.240 41.040 42.560 41.360 ;
        RECT 42.640 41.040 42.960 41.360 ;
        RECT 43.040 41.040 43.360 41.360 ;
        RECT 43.440 41.040 43.760 41.360 ;
        RECT 43.840 41.040 44.160 41.360 ;
        RECT 44.240 41.040 44.560 41.360 ;
        RECT 44.640 41.040 44.960 41.360 ;
        RECT 70.560 41.040 70.880 41.360 ;
        RECT 70.960 41.040 71.280 41.360 ;
        RECT 71.360 41.040 71.680 41.360 ;
        RECT 71.760 41.040 72.080 41.360 ;
        RECT 120.560 41.040 120.880 41.360 ;
        RECT 120.960 41.040 121.280 41.360 ;
        RECT 121.360 41.040 121.680 41.360 ;
        RECT 121.760 41.040 122.080 41.360 ;
        RECT 160.720 41.040 161.040 41.360 ;
        RECT 161.120 41.040 161.440 41.360 ;
        RECT 161.520 41.040 161.840 41.360 ;
        RECT 161.920 41.040 162.240 41.360 ;
        RECT 162.320 41.040 162.640 41.360 ;
        RECT 162.720 41.040 163.040 41.360 ;
        RECT 163.120 41.040 163.440 41.360 ;
        RECT 163.520 41.040 163.840 41.360 ;
        RECT 163.920 41.040 164.240 41.360 ;
        RECT 164.320 41.040 164.640 41.360 ;
        RECT 164.720 41.040 165.040 41.360 ;
        RECT 165.120 41.040 165.440 41.360 ;
        RECT 165.520 41.040 165.840 41.360 ;
        RECT 165.920 41.040 166.240 41.360 ;
        RECT 166.320 41.040 166.640 41.360 ;
        RECT 166.720 41.040 167.040 41.360 ;
        RECT 167.120 41.040 167.440 41.360 ;
        RECT 167.520 41.040 167.840 41.360 ;
        RECT 167.920 41.040 168.240 41.360 ;
        RECT 168.320 41.040 168.640 41.360 ;
        RECT 168.720 41.040 169.040 41.360 ;
        RECT 169.120 41.040 169.440 41.360 ;
        RECT 169.520 41.040 169.840 41.360 ;
        RECT 169.920 41.040 170.240 41.360 ;
        RECT 170.320 41.040 170.640 41.360 ;
        RECT 170.720 41.040 171.040 41.360 ;
        RECT 171.120 41.040 171.440 41.360 ;
        RECT 171.520 41.040 171.840 41.360 ;
        RECT 171.920 41.040 172.240 41.360 ;
        RECT 172.320 41.040 172.640 41.360 ;
        RECT 172.720 41.040 173.040 41.360 ;
        RECT 173.120 41.040 173.440 41.360 ;
        RECT 173.520 41.040 173.840 41.360 ;
        RECT 173.920 41.040 174.240 41.360 ;
        RECT 174.320 41.040 174.640 41.360 ;
        RECT 174.720 41.040 175.040 41.360 ;
        RECT 175.120 41.040 175.440 41.360 ;
        RECT 175.520 41.040 175.840 41.360 ;
        RECT 175.920 41.040 176.240 41.360 ;
        RECT 176.320 41.040 176.640 41.360 ;
        RECT 176.720 41.040 177.040 41.360 ;
        RECT 177.120 41.040 177.440 41.360 ;
        RECT 177.520 41.040 177.840 41.360 ;
        RECT 177.920 41.040 178.240 41.360 ;
        RECT 178.320 41.040 178.640 41.360 ;
        RECT 178.720 41.040 179.040 41.360 ;
        RECT 179.120 41.040 179.440 41.360 ;
        RECT 179.520 41.040 179.840 41.360 ;
        RECT 179.920 41.040 180.240 41.360 ;
        RECT 180.320 41.040 180.640 41.360 ;
        RECT 25.040 40.640 25.360 40.960 ;
        RECT 25.440 40.640 25.760 40.960 ;
        RECT 25.840 40.640 26.160 40.960 ;
        RECT 26.240 40.640 26.560 40.960 ;
        RECT 26.640 40.640 26.960 40.960 ;
        RECT 27.040 40.640 27.360 40.960 ;
        RECT 27.440 40.640 27.760 40.960 ;
        RECT 27.840 40.640 28.160 40.960 ;
        RECT 28.240 40.640 28.560 40.960 ;
        RECT 28.640 40.640 28.960 40.960 ;
        RECT 29.040 40.640 29.360 40.960 ;
        RECT 29.440 40.640 29.760 40.960 ;
        RECT 29.840 40.640 30.160 40.960 ;
        RECT 30.240 40.640 30.560 40.960 ;
        RECT 30.640 40.640 30.960 40.960 ;
        RECT 31.040 40.640 31.360 40.960 ;
        RECT 31.440 40.640 31.760 40.960 ;
        RECT 31.840 40.640 32.160 40.960 ;
        RECT 32.240 40.640 32.560 40.960 ;
        RECT 32.640 40.640 32.960 40.960 ;
        RECT 33.040 40.640 33.360 40.960 ;
        RECT 33.440 40.640 33.760 40.960 ;
        RECT 33.840 40.640 34.160 40.960 ;
        RECT 34.240 40.640 34.560 40.960 ;
        RECT 34.640 40.640 34.960 40.960 ;
        RECT 35.040 40.640 35.360 40.960 ;
        RECT 35.440 40.640 35.760 40.960 ;
        RECT 35.840 40.640 36.160 40.960 ;
        RECT 36.240 40.640 36.560 40.960 ;
        RECT 36.640 40.640 36.960 40.960 ;
        RECT 37.040 40.640 37.360 40.960 ;
        RECT 37.440 40.640 37.760 40.960 ;
        RECT 37.840 40.640 38.160 40.960 ;
        RECT 38.240 40.640 38.560 40.960 ;
        RECT 38.640 40.640 38.960 40.960 ;
        RECT 39.040 40.640 39.360 40.960 ;
        RECT 39.440 40.640 39.760 40.960 ;
        RECT 39.840 40.640 40.160 40.960 ;
        RECT 40.240 40.640 40.560 40.960 ;
        RECT 40.640 40.640 40.960 40.960 ;
        RECT 41.040 40.640 41.360 40.960 ;
        RECT 41.440 40.640 41.760 40.960 ;
        RECT 41.840 40.640 42.160 40.960 ;
        RECT 42.240 40.640 42.560 40.960 ;
        RECT 42.640 40.640 42.960 40.960 ;
        RECT 43.040 40.640 43.360 40.960 ;
        RECT 43.440 40.640 43.760 40.960 ;
        RECT 43.840 40.640 44.160 40.960 ;
        RECT 44.240 40.640 44.560 40.960 ;
        RECT 44.640 40.640 44.960 40.960 ;
        RECT 70.560 40.640 70.880 40.960 ;
        RECT 70.960 40.640 71.280 40.960 ;
        RECT 71.360 40.640 71.680 40.960 ;
        RECT 71.760 40.640 72.080 40.960 ;
        RECT 120.560 40.640 120.880 40.960 ;
        RECT 120.960 40.640 121.280 40.960 ;
        RECT 121.360 40.640 121.680 40.960 ;
        RECT 121.760 40.640 122.080 40.960 ;
        RECT 160.720 40.640 161.040 40.960 ;
        RECT 161.120 40.640 161.440 40.960 ;
        RECT 161.520 40.640 161.840 40.960 ;
        RECT 161.920 40.640 162.240 40.960 ;
        RECT 162.320 40.640 162.640 40.960 ;
        RECT 162.720 40.640 163.040 40.960 ;
        RECT 163.120 40.640 163.440 40.960 ;
        RECT 163.520 40.640 163.840 40.960 ;
        RECT 163.920 40.640 164.240 40.960 ;
        RECT 164.320 40.640 164.640 40.960 ;
        RECT 164.720 40.640 165.040 40.960 ;
        RECT 165.120 40.640 165.440 40.960 ;
        RECT 165.520 40.640 165.840 40.960 ;
        RECT 165.920 40.640 166.240 40.960 ;
        RECT 166.320 40.640 166.640 40.960 ;
        RECT 166.720 40.640 167.040 40.960 ;
        RECT 167.120 40.640 167.440 40.960 ;
        RECT 167.520 40.640 167.840 40.960 ;
        RECT 167.920 40.640 168.240 40.960 ;
        RECT 168.320 40.640 168.640 40.960 ;
        RECT 168.720 40.640 169.040 40.960 ;
        RECT 169.120 40.640 169.440 40.960 ;
        RECT 169.520 40.640 169.840 40.960 ;
        RECT 169.920 40.640 170.240 40.960 ;
        RECT 170.320 40.640 170.640 40.960 ;
        RECT 170.720 40.640 171.040 40.960 ;
        RECT 171.120 40.640 171.440 40.960 ;
        RECT 171.520 40.640 171.840 40.960 ;
        RECT 171.920 40.640 172.240 40.960 ;
        RECT 172.320 40.640 172.640 40.960 ;
        RECT 172.720 40.640 173.040 40.960 ;
        RECT 173.120 40.640 173.440 40.960 ;
        RECT 173.520 40.640 173.840 40.960 ;
        RECT 173.920 40.640 174.240 40.960 ;
        RECT 174.320 40.640 174.640 40.960 ;
        RECT 174.720 40.640 175.040 40.960 ;
        RECT 175.120 40.640 175.440 40.960 ;
        RECT 175.520 40.640 175.840 40.960 ;
        RECT 175.920 40.640 176.240 40.960 ;
        RECT 176.320 40.640 176.640 40.960 ;
        RECT 176.720 40.640 177.040 40.960 ;
        RECT 177.120 40.640 177.440 40.960 ;
        RECT 177.520 40.640 177.840 40.960 ;
        RECT 177.920 40.640 178.240 40.960 ;
        RECT 178.320 40.640 178.640 40.960 ;
        RECT 178.720 40.640 179.040 40.960 ;
        RECT 179.120 40.640 179.440 40.960 ;
        RECT 179.520 40.640 179.840 40.960 ;
        RECT 179.920 40.640 180.240 40.960 ;
        RECT 180.320 40.640 180.640 40.960 ;
        RECT 25.040 40.240 25.360 40.560 ;
        RECT 25.440 40.240 25.760 40.560 ;
        RECT 25.840 40.240 26.160 40.560 ;
        RECT 26.240 40.240 26.560 40.560 ;
        RECT 26.640 40.240 26.960 40.560 ;
        RECT 27.040 40.240 27.360 40.560 ;
        RECT 27.440 40.240 27.760 40.560 ;
        RECT 27.840 40.240 28.160 40.560 ;
        RECT 28.240 40.240 28.560 40.560 ;
        RECT 28.640 40.240 28.960 40.560 ;
        RECT 29.040 40.240 29.360 40.560 ;
        RECT 29.440 40.240 29.760 40.560 ;
        RECT 29.840 40.240 30.160 40.560 ;
        RECT 30.240 40.240 30.560 40.560 ;
        RECT 30.640 40.240 30.960 40.560 ;
        RECT 31.040 40.240 31.360 40.560 ;
        RECT 31.440 40.240 31.760 40.560 ;
        RECT 31.840 40.240 32.160 40.560 ;
        RECT 32.240 40.240 32.560 40.560 ;
        RECT 32.640 40.240 32.960 40.560 ;
        RECT 33.040 40.240 33.360 40.560 ;
        RECT 33.440 40.240 33.760 40.560 ;
        RECT 33.840 40.240 34.160 40.560 ;
        RECT 34.240 40.240 34.560 40.560 ;
        RECT 34.640 40.240 34.960 40.560 ;
        RECT 35.040 40.240 35.360 40.560 ;
        RECT 35.440 40.240 35.760 40.560 ;
        RECT 35.840 40.240 36.160 40.560 ;
        RECT 36.240 40.240 36.560 40.560 ;
        RECT 36.640 40.240 36.960 40.560 ;
        RECT 37.040 40.240 37.360 40.560 ;
        RECT 37.440 40.240 37.760 40.560 ;
        RECT 37.840 40.240 38.160 40.560 ;
        RECT 38.240 40.240 38.560 40.560 ;
        RECT 38.640 40.240 38.960 40.560 ;
        RECT 39.040 40.240 39.360 40.560 ;
        RECT 39.440 40.240 39.760 40.560 ;
        RECT 39.840 40.240 40.160 40.560 ;
        RECT 40.240 40.240 40.560 40.560 ;
        RECT 40.640 40.240 40.960 40.560 ;
        RECT 41.040 40.240 41.360 40.560 ;
        RECT 41.440 40.240 41.760 40.560 ;
        RECT 41.840 40.240 42.160 40.560 ;
        RECT 42.240 40.240 42.560 40.560 ;
        RECT 42.640 40.240 42.960 40.560 ;
        RECT 43.040 40.240 43.360 40.560 ;
        RECT 43.440 40.240 43.760 40.560 ;
        RECT 43.840 40.240 44.160 40.560 ;
        RECT 44.240 40.240 44.560 40.560 ;
        RECT 44.640 40.240 44.960 40.560 ;
        RECT 70.560 40.240 70.880 40.560 ;
        RECT 70.960 40.240 71.280 40.560 ;
        RECT 71.360 40.240 71.680 40.560 ;
        RECT 71.760 40.240 72.080 40.560 ;
        RECT 120.560 40.240 120.880 40.560 ;
        RECT 120.960 40.240 121.280 40.560 ;
        RECT 121.360 40.240 121.680 40.560 ;
        RECT 121.760 40.240 122.080 40.560 ;
        RECT 160.720 40.240 161.040 40.560 ;
        RECT 161.120 40.240 161.440 40.560 ;
        RECT 161.520 40.240 161.840 40.560 ;
        RECT 161.920 40.240 162.240 40.560 ;
        RECT 162.320 40.240 162.640 40.560 ;
        RECT 162.720 40.240 163.040 40.560 ;
        RECT 163.120 40.240 163.440 40.560 ;
        RECT 163.520 40.240 163.840 40.560 ;
        RECT 163.920 40.240 164.240 40.560 ;
        RECT 164.320 40.240 164.640 40.560 ;
        RECT 164.720 40.240 165.040 40.560 ;
        RECT 165.120 40.240 165.440 40.560 ;
        RECT 165.520 40.240 165.840 40.560 ;
        RECT 165.920 40.240 166.240 40.560 ;
        RECT 166.320 40.240 166.640 40.560 ;
        RECT 166.720 40.240 167.040 40.560 ;
        RECT 167.120 40.240 167.440 40.560 ;
        RECT 167.520 40.240 167.840 40.560 ;
        RECT 167.920 40.240 168.240 40.560 ;
        RECT 168.320 40.240 168.640 40.560 ;
        RECT 168.720 40.240 169.040 40.560 ;
        RECT 169.120 40.240 169.440 40.560 ;
        RECT 169.520 40.240 169.840 40.560 ;
        RECT 169.920 40.240 170.240 40.560 ;
        RECT 170.320 40.240 170.640 40.560 ;
        RECT 170.720 40.240 171.040 40.560 ;
        RECT 171.120 40.240 171.440 40.560 ;
        RECT 171.520 40.240 171.840 40.560 ;
        RECT 171.920 40.240 172.240 40.560 ;
        RECT 172.320 40.240 172.640 40.560 ;
        RECT 172.720 40.240 173.040 40.560 ;
        RECT 173.120 40.240 173.440 40.560 ;
        RECT 173.520 40.240 173.840 40.560 ;
        RECT 173.920 40.240 174.240 40.560 ;
        RECT 174.320 40.240 174.640 40.560 ;
        RECT 174.720 40.240 175.040 40.560 ;
        RECT 175.120 40.240 175.440 40.560 ;
        RECT 175.520 40.240 175.840 40.560 ;
        RECT 175.920 40.240 176.240 40.560 ;
        RECT 176.320 40.240 176.640 40.560 ;
        RECT 176.720 40.240 177.040 40.560 ;
        RECT 177.120 40.240 177.440 40.560 ;
        RECT 177.520 40.240 177.840 40.560 ;
        RECT 177.920 40.240 178.240 40.560 ;
        RECT 178.320 40.240 178.640 40.560 ;
        RECT 178.720 40.240 179.040 40.560 ;
        RECT 179.120 40.240 179.440 40.560 ;
        RECT 179.520 40.240 179.840 40.560 ;
        RECT 179.920 40.240 180.240 40.560 ;
        RECT 180.320 40.240 180.640 40.560 ;
        RECT 25.040 39.840 25.360 40.160 ;
        RECT 25.440 39.840 25.760 40.160 ;
        RECT 25.840 39.840 26.160 40.160 ;
        RECT 26.240 39.840 26.560 40.160 ;
        RECT 26.640 39.840 26.960 40.160 ;
        RECT 27.040 39.840 27.360 40.160 ;
        RECT 27.440 39.840 27.760 40.160 ;
        RECT 27.840 39.840 28.160 40.160 ;
        RECT 28.240 39.840 28.560 40.160 ;
        RECT 28.640 39.840 28.960 40.160 ;
        RECT 29.040 39.840 29.360 40.160 ;
        RECT 29.440 39.840 29.760 40.160 ;
        RECT 29.840 39.840 30.160 40.160 ;
        RECT 30.240 39.840 30.560 40.160 ;
        RECT 30.640 39.840 30.960 40.160 ;
        RECT 31.040 39.840 31.360 40.160 ;
        RECT 31.440 39.840 31.760 40.160 ;
        RECT 31.840 39.840 32.160 40.160 ;
        RECT 32.240 39.840 32.560 40.160 ;
        RECT 32.640 39.840 32.960 40.160 ;
        RECT 33.040 39.840 33.360 40.160 ;
        RECT 33.440 39.840 33.760 40.160 ;
        RECT 33.840 39.840 34.160 40.160 ;
        RECT 34.240 39.840 34.560 40.160 ;
        RECT 34.640 39.840 34.960 40.160 ;
        RECT 35.040 39.840 35.360 40.160 ;
        RECT 35.440 39.840 35.760 40.160 ;
        RECT 35.840 39.840 36.160 40.160 ;
        RECT 36.240 39.840 36.560 40.160 ;
        RECT 36.640 39.840 36.960 40.160 ;
        RECT 37.040 39.840 37.360 40.160 ;
        RECT 37.440 39.840 37.760 40.160 ;
        RECT 37.840 39.840 38.160 40.160 ;
        RECT 38.240 39.840 38.560 40.160 ;
        RECT 38.640 39.840 38.960 40.160 ;
        RECT 39.040 39.840 39.360 40.160 ;
        RECT 39.440 39.840 39.760 40.160 ;
        RECT 39.840 39.840 40.160 40.160 ;
        RECT 40.240 39.840 40.560 40.160 ;
        RECT 40.640 39.840 40.960 40.160 ;
        RECT 41.040 39.840 41.360 40.160 ;
        RECT 41.440 39.840 41.760 40.160 ;
        RECT 41.840 39.840 42.160 40.160 ;
        RECT 42.240 39.840 42.560 40.160 ;
        RECT 42.640 39.840 42.960 40.160 ;
        RECT 43.040 39.840 43.360 40.160 ;
        RECT 43.440 39.840 43.760 40.160 ;
        RECT 43.840 39.840 44.160 40.160 ;
        RECT 44.240 39.840 44.560 40.160 ;
        RECT 44.640 39.840 44.960 40.160 ;
        RECT 70.560 39.840 70.880 40.160 ;
        RECT 70.960 39.840 71.280 40.160 ;
        RECT 71.360 39.840 71.680 40.160 ;
        RECT 71.760 39.840 72.080 40.160 ;
        RECT 120.560 39.840 120.880 40.160 ;
        RECT 120.960 39.840 121.280 40.160 ;
        RECT 121.360 39.840 121.680 40.160 ;
        RECT 121.760 39.840 122.080 40.160 ;
        RECT 160.720 39.840 161.040 40.160 ;
        RECT 161.120 39.840 161.440 40.160 ;
        RECT 161.520 39.840 161.840 40.160 ;
        RECT 161.920 39.840 162.240 40.160 ;
        RECT 162.320 39.840 162.640 40.160 ;
        RECT 162.720 39.840 163.040 40.160 ;
        RECT 163.120 39.840 163.440 40.160 ;
        RECT 163.520 39.840 163.840 40.160 ;
        RECT 163.920 39.840 164.240 40.160 ;
        RECT 164.320 39.840 164.640 40.160 ;
        RECT 164.720 39.840 165.040 40.160 ;
        RECT 165.120 39.840 165.440 40.160 ;
        RECT 165.520 39.840 165.840 40.160 ;
        RECT 165.920 39.840 166.240 40.160 ;
        RECT 166.320 39.840 166.640 40.160 ;
        RECT 166.720 39.840 167.040 40.160 ;
        RECT 167.120 39.840 167.440 40.160 ;
        RECT 167.520 39.840 167.840 40.160 ;
        RECT 167.920 39.840 168.240 40.160 ;
        RECT 168.320 39.840 168.640 40.160 ;
        RECT 168.720 39.840 169.040 40.160 ;
        RECT 169.120 39.840 169.440 40.160 ;
        RECT 169.520 39.840 169.840 40.160 ;
        RECT 169.920 39.840 170.240 40.160 ;
        RECT 170.320 39.840 170.640 40.160 ;
        RECT 170.720 39.840 171.040 40.160 ;
        RECT 171.120 39.840 171.440 40.160 ;
        RECT 171.520 39.840 171.840 40.160 ;
        RECT 171.920 39.840 172.240 40.160 ;
        RECT 172.320 39.840 172.640 40.160 ;
        RECT 172.720 39.840 173.040 40.160 ;
        RECT 173.120 39.840 173.440 40.160 ;
        RECT 173.520 39.840 173.840 40.160 ;
        RECT 173.920 39.840 174.240 40.160 ;
        RECT 174.320 39.840 174.640 40.160 ;
        RECT 174.720 39.840 175.040 40.160 ;
        RECT 175.120 39.840 175.440 40.160 ;
        RECT 175.520 39.840 175.840 40.160 ;
        RECT 175.920 39.840 176.240 40.160 ;
        RECT 176.320 39.840 176.640 40.160 ;
        RECT 176.720 39.840 177.040 40.160 ;
        RECT 177.120 39.840 177.440 40.160 ;
        RECT 177.520 39.840 177.840 40.160 ;
        RECT 177.920 39.840 178.240 40.160 ;
        RECT 178.320 39.840 178.640 40.160 ;
        RECT 178.720 39.840 179.040 40.160 ;
        RECT 179.120 39.840 179.440 40.160 ;
        RECT 179.520 39.840 179.840 40.160 ;
        RECT 179.920 39.840 180.240 40.160 ;
        RECT 180.320 39.840 180.640 40.160 ;
        RECT 25.040 39.440 25.360 39.760 ;
        RECT 25.440 39.440 25.760 39.760 ;
        RECT 25.840 39.440 26.160 39.760 ;
        RECT 26.240 39.440 26.560 39.760 ;
        RECT 26.640 39.440 26.960 39.760 ;
        RECT 27.040 39.440 27.360 39.760 ;
        RECT 27.440 39.440 27.760 39.760 ;
        RECT 27.840 39.440 28.160 39.760 ;
        RECT 28.240 39.440 28.560 39.760 ;
        RECT 28.640 39.440 28.960 39.760 ;
        RECT 29.040 39.440 29.360 39.760 ;
        RECT 29.440 39.440 29.760 39.760 ;
        RECT 29.840 39.440 30.160 39.760 ;
        RECT 30.240 39.440 30.560 39.760 ;
        RECT 30.640 39.440 30.960 39.760 ;
        RECT 31.040 39.440 31.360 39.760 ;
        RECT 31.440 39.440 31.760 39.760 ;
        RECT 31.840 39.440 32.160 39.760 ;
        RECT 32.240 39.440 32.560 39.760 ;
        RECT 32.640 39.440 32.960 39.760 ;
        RECT 33.040 39.440 33.360 39.760 ;
        RECT 33.440 39.440 33.760 39.760 ;
        RECT 33.840 39.440 34.160 39.760 ;
        RECT 34.240 39.440 34.560 39.760 ;
        RECT 34.640 39.440 34.960 39.760 ;
        RECT 35.040 39.440 35.360 39.760 ;
        RECT 35.440 39.440 35.760 39.760 ;
        RECT 35.840 39.440 36.160 39.760 ;
        RECT 36.240 39.440 36.560 39.760 ;
        RECT 36.640 39.440 36.960 39.760 ;
        RECT 37.040 39.440 37.360 39.760 ;
        RECT 37.440 39.440 37.760 39.760 ;
        RECT 37.840 39.440 38.160 39.760 ;
        RECT 38.240 39.440 38.560 39.760 ;
        RECT 38.640 39.440 38.960 39.760 ;
        RECT 39.040 39.440 39.360 39.760 ;
        RECT 39.440 39.440 39.760 39.760 ;
        RECT 39.840 39.440 40.160 39.760 ;
        RECT 40.240 39.440 40.560 39.760 ;
        RECT 40.640 39.440 40.960 39.760 ;
        RECT 41.040 39.440 41.360 39.760 ;
        RECT 41.440 39.440 41.760 39.760 ;
        RECT 41.840 39.440 42.160 39.760 ;
        RECT 42.240 39.440 42.560 39.760 ;
        RECT 42.640 39.440 42.960 39.760 ;
        RECT 43.040 39.440 43.360 39.760 ;
        RECT 43.440 39.440 43.760 39.760 ;
        RECT 43.840 39.440 44.160 39.760 ;
        RECT 44.240 39.440 44.560 39.760 ;
        RECT 44.640 39.440 44.960 39.760 ;
        RECT 70.560 39.440 70.880 39.760 ;
        RECT 70.960 39.440 71.280 39.760 ;
        RECT 71.360 39.440 71.680 39.760 ;
        RECT 71.760 39.440 72.080 39.760 ;
        RECT 120.560 39.440 120.880 39.760 ;
        RECT 120.960 39.440 121.280 39.760 ;
        RECT 121.360 39.440 121.680 39.760 ;
        RECT 121.760 39.440 122.080 39.760 ;
        RECT 160.720 39.440 161.040 39.760 ;
        RECT 161.120 39.440 161.440 39.760 ;
        RECT 161.520 39.440 161.840 39.760 ;
        RECT 161.920 39.440 162.240 39.760 ;
        RECT 162.320 39.440 162.640 39.760 ;
        RECT 162.720 39.440 163.040 39.760 ;
        RECT 163.120 39.440 163.440 39.760 ;
        RECT 163.520 39.440 163.840 39.760 ;
        RECT 163.920 39.440 164.240 39.760 ;
        RECT 164.320 39.440 164.640 39.760 ;
        RECT 164.720 39.440 165.040 39.760 ;
        RECT 165.120 39.440 165.440 39.760 ;
        RECT 165.520 39.440 165.840 39.760 ;
        RECT 165.920 39.440 166.240 39.760 ;
        RECT 166.320 39.440 166.640 39.760 ;
        RECT 166.720 39.440 167.040 39.760 ;
        RECT 167.120 39.440 167.440 39.760 ;
        RECT 167.520 39.440 167.840 39.760 ;
        RECT 167.920 39.440 168.240 39.760 ;
        RECT 168.320 39.440 168.640 39.760 ;
        RECT 168.720 39.440 169.040 39.760 ;
        RECT 169.120 39.440 169.440 39.760 ;
        RECT 169.520 39.440 169.840 39.760 ;
        RECT 169.920 39.440 170.240 39.760 ;
        RECT 170.320 39.440 170.640 39.760 ;
        RECT 170.720 39.440 171.040 39.760 ;
        RECT 171.120 39.440 171.440 39.760 ;
        RECT 171.520 39.440 171.840 39.760 ;
        RECT 171.920 39.440 172.240 39.760 ;
        RECT 172.320 39.440 172.640 39.760 ;
        RECT 172.720 39.440 173.040 39.760 ;
        RECT 173.120 39.440 173.440 39.760 ;
        RECT 173.520 39.440 173.840 39.760 ;
        RECT 173.920 39.440 174.240 39.760 ;
        RECT 174.320 39.440 174.640 39.760 ;
        RECT 174.720 39.440 175.040 39.760 ;
        RECT 175.120 39.440 175.440 39.760 ;
        RECT 175.520 39.440 175.840 39.760 ;
        RECT 175.920 39.440 176.240 39.760 ;
        RECT 176.320 39.440 176.640 39.760 ;
        RECT 176.720 39.440 177.040 39.760 ;
        RECT 177.120 39.440 177.440 39.760 ;
        RECT 177.520 39.440 177.840 39.760 ;
        RECT 177.920 39.440 178.240 39.760 ;
        RECT 178.320 39.440 178.640 39.760 ;
        RECT 178.720 39.440 179.040 39.760 ;
        RECT 179.120 39.440 179.440 39.760 ;
        RECT 179.520 39.440 179.840 39.760 ;
        RECT 179.920 39.440 180.240 39.760 ;
        RECT 180.320 39.440 180.640 39.760 ;
        RECT 25.040 39.040 25.360 39.360 ;
        RECT 25.440 39.040 25.760 39.360 ;
        RECT 25.840 39.040 26.160 39.360 ;
        RECT 26.240 39.040 26.560 39.360 ;
        RECT 26.640 39.040 26.960 39.360 ;
        RECT 27.040 39.040 27.360 39.360 ;
        RECT 27.440 39.040 27.760 39.360 ;
        RECT 27.840 39.040 28.160 39.360 ;
        RECT 28.240 39.040 28.560 39.360 ;
        RECT 28.640 39.040 28.960 39.360 ;
        RECT 29.040 39.040 29.360 39.360 ;
        RECT 29.440 39.040 29.760 39.360 ;
        RECT 29.840 39.040 30.160 39.360 ;
        RECT 30.240 39.040 30.560 39.360 ;
        RECT 30.640 39.040 30.960 39.360 ;
        RECT 31.040 39.040 31.360 39.360 ;
        RECT 31.440 39.040 31.760 39.360 ;
        RECT 31.840 39.040 32.160 39.360 ;
        RECT 32.240 39.040 32.560 39.360 ;
        RECT 32.640 39.040 32.960 39.360 ;
        RECT 33.040 39.040 33.360 39.360 ;
        RECT 33.440 39.040 33.760 39.360 ;
        RECT 33.840 39.040 34.160 39.360 ;
        RECT 34.240 39.040 34.560 39.360 ;
        RECT 34.640 39.040 34.960 39.360 ;
        RECT 35.040 39.040 35.360 39.360 ;
        RECT 35.440 39.040 35.760 39.360 ;
        RECT 35.840 39.040 36.160 39.360 ;
        RECT 36.240 39.040 36.560 39.360 ;
        RECT 36.640 39.040 36.960 39.360 ;
        RECT 37.040 39.040 37.360 39.360 ;
        RECT 37.440 39.040 37.760 39.360 ;
        RECT 37.840 39.040 38.160 39.360 ;
        RECT 38.240 39.040 38.560 39.360 ;
        RECT 38.640 39.040 38.960 39.360 ;
        RECT 39.040 39.040 39.360 39.360 ;
        RECT 39.440 39.040 39.760 39.360 ;
        RECT 39.840 39.040 40.160 39.360 ;
        RECT 40.240 39.040 40.560 39.360 ;
        RECT 40.640 39.040 40.960 39.360 ;
        RECT 41.040 39.040 41.360 39.360 ;
        RECT 41.440 39.040 41.760 39.360 ;
        RECT 41.840 39.040 42.160 39.360 ;
        RECT 42.240 39.040 42.560 39.360 ;
        RECT 42.640 39.040 42.960 39.360 ;
        RECT 43.040 39.040 43.360 39.360 ;
        RECT 43.440 39.040 43.760 39.360 ;
        RECT 43.840 39.040 44.160 39.360 ;
        RECT 44.240 39.040 44.560 39.360 ;
        RECT 44.640 39.040 44.960 39.360 ;
        RECT 70.560 39.040 70.880 39.360 ;
        RECT 70.960 39.040 71.280 39.360 ;
        RECT 71.360 39.040 71.680 39.360 ;
        RECT 71.760 39.040 72.080 39.360 ;
        RECT 120.560 39.040 120.880 39.360 ;
        RECT 120.960 39.040 121.280 39.360 ;
        RECT 121.360 39.040 121.680 39.360 ;
        RECT 121.760 39.040 122.080 39.360 ;
        RECT 160.720 39.040 161.040 39.360 ;
        RECT 161.120 39.040 161.440 39.360 ;
        RECT 161.520 39.040 161.840 39.360 ;
        RECT 161.920 39.040 162.240 39.360 ;
        RECT 162.320 39.040 162.640 39.360 ;
        RECT 162.720 39.040 163.040 39.360 ;
        RECT 163.120 39.040 163.440 39.360 ;
        RECT 163.520 39.040 163.840 39.360 ;
        RECT 163.920 39.040 164.240 39.360 ;
        RECT 164.320 39.040 164.640 39.360 ;
        RECT 164.720 39.040 165.040 39.360 ;
        RECT 165.120 39.040 165.440 39.360 ;
        RECT 165.520 39.040 165.840 39.360 ;
        RECT 165.920 39.040 166.240 39.360 ;
        RECT 166.320 39.040 166.640 39.360 ;
        RECT 166.720 39.040 167.040 39.360 ;
        RECT 167.120 39.040 167.440 39.360 ;
        RECT 167.520 39.040 167.840 39.360 ;
        RECT 167.920 39.040 168.240 39.360 ;
        RECT 168.320 39.040 168.640 39.360 ;
        RECT 168.720 39.040 169.040 39.360 ;
        RECT 169.120 39.040 169.440 39.360 ;
        RECT 169.520 39.040 169.840 39.360 ;
        RECT 169.920 39.040 170.240 39.360 ;
        RECT 170.320 39.040 170.640 39.360 ;
        RECT 170.720 39.040 171.040 39.360 ;
        RECT 171.120 39.040 171.440 39.360 ;
        RECT 171.520 39.040 171.840 39.360 ;
        RECT 171.920 39.040 172.240 39.360 ;
        RECT 172.320 39.040 172.640 39.360 ;
        RECT 172.720 39.040 173.040 39.360 ;
        RECT 173.120 39.040 173.440 39.360 ;
        RECT 173.520 39.040 173.840 39.360 ;
        RECT 173.920 39.040 174.240 39.360 ;
        RECT 174.320 39.040 174.640 39.360 ;
        RECT 174.720 39.040 175.040 39.360 ;
        RECT 175.120 39.040 175.440 39.360 ;
        RECT 175.520 39.040 175.840 39.360 ;
        RECT 175.920 39.040 176.240 39.360 ;
        RECT 176.320 39.040 176.640 39.360 ;
        RECT 176.720 39.040 177.040 39.360 ;
        RECT 177.120 39.040 177.440 39.360 ;
        RECT 177.520 39.040 177.840 39.360 ;
        RECT 177.920 39.040 178.240 39.360 ;
        RECT 178.320 39.040 178.640 39.360 ;
        RECT 178.720 39.040 179.040 39.360 ;
        RECT 179.120 39.040 179.440 39.360 ;
        RECT 179.520 39.040 179.840 39.360 ;
        RECT 179.920 39.040 180.240 39.360 ;
        RECT 180.320 39.040 180.640 39.360 ;
        RECT 25.040 38.640 25.360 38.960 ;
        RECT 25.440 38.640 25.760 38.960 ;
        RECT 25.840 38.640 26.160 38.960 ;
        RECT 26.240 38.640 26.560 38.960 ;
        RECT 26.640 38.640 26.960 38.960 ;
        RECT 27.040 38.640 27.360 38.960 ;
        RECT 27.440 38.640 27.760 38.960 ;
        RECT 27.840 38.640 28.160 38.960 ;
        RECT 28.240 38.640 28.560 38.960 ;
        RECT 28.640 38.640 28.960 38.960 ;
        RECT 29.040 38.640 29.360 38.960 ;
        RECT 29.440 38.640 29.760 38.960 ;
        RECT 29.840 38.640 30.160 38.960 ;
        RECT 30.240 38.640 30.560 38.960 ;
        RECT 30.640 38.640 30.960 38.960 ;
        RECT 31.040 38.640 31.360 38.960 ;
        RECT 31.440 38.640 31.760 38.960 ;
        RECT 31.840 38.640 32.160 38.960 ;
        RECT 32.240 38.640 32.560 38.960 ;
        RECT 32.640 38.640 32.960 38.960 ;
        RECT 33.040 38.640 33.360 38.960 ;
        RECT 33.440 38.640 33.760 38.960 ;
        RECT 33.840 38.640 34.160 38.960 ;
        RECT 34.240 38.640 34.560 38.960 ;
        RECT 34.640 38.640 34.960 38.960 ;
        RECT 35.040 38.640 35.360 38.960 ;
        RECT 35.440 38.640 35.760 38.960 ;
        RECT 35.840 38.640 36.160 38.960 ;
        RECT 36.240 38.640 36.560 38.960 ;
        RECT 36.640 38.640 36.960 38.960 ;
        RECT 37.040 38.640 37.360 38.960 ;
        RECT 37.440 38.640 37.760 38.960 ;
        RECT 37.840 38.640 38.160 38.960 ;
        RECT 38.240 38.640 38.560 38.960 ;
        RECT 38.640 38.640 38.960 38.960 ;
        RECT 39.040 38.640 39.360 38.960 ;
        RECT 39.440 38.640 39.760 38.960 ;
        RECT 39.840 38.640 40.160 38.960 ;
        RECT 40.240 38.640 40.560 38.960 ;
        RECT 40.640 38.640 40.960 38.960 ;
        RECT 41.040 38.640 41.360 38.960 ;
        RECT 41.440 38.640 41.760 38.960 ;
        RECT 41.840 38.640 42.160 38.960 ;
        RECT 42.240 38.640 42.560 38.960 ;
        RECT 42.640 38.640 42.960 38.960 ;
        RECT 43.040 38.640 43.360 38.960 ;
        RECT 43.440 38.640 43.760 38.960 ;
        RECT 43.840 38.640 44.160 38.960 ;
        RECT 44.240 38.640 44.560 38.960 ;
        RECT 44.640 38.640 44.960 38.960 ;
        RECT 70.560 38.640 70.880 38.960 ;
        RECT 70.960 38.640 71.280 38.960 ;
        RECT 71.360 38.640 71.680 38.960 ;
        RECT 71.760 38.640 72.080 38.960 ;
        RECT 120.560 38.640 120.880 38.960 ;
        RECT 120.960 38.640 121.280 38.960 ;
        RECT 121.360 38.640 121.680 38.960 ;
        RECT 121.760 38.640 122.080 38.960 ;
        RECT 160.720 38.640 161.040 38.960 ;
        RECT 161.120 38.640 161.440 38.960 ;
        RECT 161.520 38.640 161.840 38.960 ;
        RECT 161.920 38.640 162.240 38.960 ;
        RECT 162.320 38.640 162.640 38.960 ;
        RECT 162.720 38.640 163.040 38.960 ;
        RECT 163.120 38.640 163.440 38.960 ;
        RECT 163.520 38.640 163.840 38.960 ;
        RECT 163.920 38.640 164.240 38.960 ;
        RECT 164.320 38.640 164.640 38.960 ;
        RECT 164.720 38.640 165.040 38.960 ;
        RECT 165.120 38.640 165.440 38.960 ;
        RECT 165.520 38.640 165.840 38.960 ;
        RECT 165.920 38.640 166.240 38.960 ;
        RECT 166.320 38.640 166.640 38.960 ;
        RECT 166.720 38.640 167.040 38.960 ;
        RECT 167.120 38.640 167.440 38.960 ;
        RECT 167.520 38.640 167.840 38.960 ;
        RECT 167.920 38.640 168.240 38.960 ;
        RECT 168.320 38.640 168.640 38.960 ;
        RECT 168.720 38.640 169.040 38.960 ;
        RECT 169.120 38.640 169.440 38.960 ;
        RECT 169.520 38.640 169.840 38.960 ;
        RECT 169.920 38.640 170.240 38.960 ;
        RECT 170.320 38.640 170.640 38.960 ;
        RECT 170.720 38.640 171.040 38.960 ;
        RECT 171.120 38.640 171.440 38.960 ;
        RECT 171.520 38.640 171.840 38.960 ;
        RECT 171.920 38.640 172.240 38.960 ;
        RECT 172.320 38.640 172.640 38.960 ;
        RECT 172.720 38.640 173.040 38.960 ;
        RECT 173.120 38.640 173.440 38.960 ;
        RECT 173.520 38.640 173.840 38.960 ;
        RECT 173.920 38.640 174.240 38.960 ;
        RECT 174.320 38.640 174.640 38.960 ;
        RECT 174.720 38.640 175.040 38.960 ;
        RECT 175.120 38.640 175.440 38.960 ;
        RECT 175.520 38.640 175.840 38.960 ;
        RECT 175.920 38.640 176.240 38.960 ;
        RECT 176.320 38.640 176.640 38.960 ;
        RECT 176.720 38.640 177.040 38.960 ;
        RECT 177.120 38.640 177.440 38.960 ;
        RECT 177.520 38.640 177.840 38.960 ;
        RECT 177.920 38.640 178.240 38.960 ;
        RECT 178.320 38.640 178.640 38.960 ;
        RECT 178.720 38.640 179.040 38.960 ;
        RECT 179.120 38.640 179.440 38.960 ;
        RECT 179.520 38.640 179.840 38.960 ;
        RECT 179.920 38.640 180.240 38.960 ;
        RECT 180.320 38.640 180.640 38.960 ;
        RECT 25.040 38.240 25.360 38.560 ;
        RECT 25.440 38.240 25.760 38.560 ;
        RECT 25.840 38.240 26.160 38.560 ;
        RECT 26.240 38.240 26.560 38.560 ;
        RECT 26.640 38.240 26.960 38.560 ;
        RECT 27.040 38.240 27.360 38.560 ;
        RECT 27.440 38.240 27.760 38.560 ;
        RECT 27.840 38.240 28.160 38.560 ;
        RECT 28.240 38.240 28.560 38.560 ;
        RECT 28.640 38.240 28.960 38.560 ;
        RECT 29.040 38.240 29.360 38.560 ;
        RECT 29.440 38.240 29.760 38.560 ;
        RECT 29.840 38.240 30.160 38.560 ;
        RECT 30.240 38.240 30.560 38.560 ;
        RECT 30.640 38.240 30.960 38.560 ;
        RECT 31.040 38.240 31.360 38.560 ;
        RECT 31.440 38.240 31.760 38.560 ;
        RECT 31.840 38.240 32.160 38.560 ;
        RECT 32.240 38.240 32.560 38.560 ;
        RECT 32.640 38.240 32.960 38.560 ;
        RECT 33.040 38.240 33.360 38.560 ;
        RECT 33.440 38.240 33.760 38.560 ;
        RECT 33.840 38.240 34.160 38.560 ;
        RECT 34.240 38.240 34.560 38.560 ;
        RECT 34.640 38.240 34.960 38.560 ;
        RECT 35.040 38.240 35.360 38.560 ;
        RECT 35.440 38.240 35.760 38.560 ;
        RECT 35.840 38.240 36.160 38.560 ;
        RECT 36.240 38.240 36.560 38.560 ;
        RECT 36.640 38.240 36.960 38.560 ;
        RECT 37.040 38.240 37.360 38.560 ;
        RECT 37.440 38.240 37.760 38.560 ;
        RECT 37.840 38.240 38.160 38.560 ;
        RECT 38.240 38.240 38.560 38.560 ;
        RECT 38.640 38.240 38.960 38.560 ;
        RECT 39.040 38.240 39.360 38.560 ;
        RECT 39.440 38.240 39.760 38.560 ;
        RECT 39.840 38.240 40.160 38.560 ;
        RECT 40.240 38.240 40.560 38.560 ;
        RECT 40.640 38.240 40.960 38.560 ;
        RECT 41.040 38.240 41.360 38.560 ;
        RECT 41.440 38.240 41.760 38.560 ;
        RECT 41.840 38.240 42.160 38.560 ;
        RECT 42.240 38.240 42.560 38.560 ;
        RECT 42.640 38.240 42.960 38.560 ;
        RECT 43.040 38.240 43.360 38.560 ;
        RECT 43.440 38.240 43.760 38.560 ;
        RECT 43.840 38.240 44.160 38.560 ;
        RECT 44.240 38.240 44.560 38.560 ;
        RECT 44.640 38.240 44.960 38.560 ;
        RECT 70.560 38.240 70.880 38.560 ;
        RECT 70.960 38.240 71.280 38.560 ;
        RECT 71.360 38.240 71.680 38.560 ;
        RECT 71.760 38.240 72.080 38.560 ;
        RECT 120.560 38.240 120.880 38.560 ;
        RECT 120.960 38.240 121.280 38.560 ;
        RECT 121.360 38.240 121.680 38.560 ;
        RECT 121.760 38.240 122.080 38.560 ;
        RECT 160.720 38.240 161.040 38.560 ;
        RECT 161.120 38.240 161.440 38.560 ;
        RECT 161.520 38.240 161.840 38.560 ;
        RECT 161.920 38.240 162.240 38.560 ;
        RECT 162.320 38.240 162.640 38.560 ;
        RECT 162.720 38.240 163.040 38.560 ;
        RECT 163.120 38.240 163.440 38.560 ;
        RECT 163.520 38.240 163.840 38.560 ;
        RECT 163.920 38.240 164.240 38.560 ;
        RECT 164.320 38.240 164.640 38.560 ;
        RECT 164.720 38.240 165.040 38.560 ;
        RECT 165.120 38.240 165.440 38.560 ;
        RECT 165.520 38.240 165.840 38.560 ;
        RECT 165.920 38.240 166.240 38.560 ;
        RECT 166.320 38.240 166.640 38.560 ;
        RECT 166.720 38.240 167.040 38.560 ;
        RECT 167.120 38.240 167.440 38.560 ;
        RECT 167.520 38.240 167.840 38.560 ;
        RECT 167.920 38.240 168.240 38.560 ;
        RECT 168.320 38.240 168.640 38.560 ;
        RECT 168.720 38.240 169.040 38.560 ;
        RECT 169.120 38.240 169.440 38.560 ;
        RECT 169.520 38.240 169.840 38.560 ;
        RECT 169.920 38.240 170.240 38.560 ;
        RECT 170.320 38.240 170.640 38.560 ;
        RECT 170.720 38.240 171.040 38.560 ;
        RECT 171.120 38.240 171.440 38.560 ;
        RECT 171.520 38.240 171.840 38.560 ;
        RECT 171.920 38.240 172.240 38.560 ;
        RECT 172.320 38.240 172.640 38.560 ;
        RECT 172.720 38.240 173.040 38.560 ;
        RECT 173.120 38.240 173.440 38.560 ;
        RECT 173.520 38.240 173.840 38.560 ;
        RECT 173.920 38.240 174.240 38.560 ;
        RECT 174.320 38.240 174.640 38.560 ;
        RECT 174.720 38.240 175.040 38.560 ;
        RECT 175.120 38.240 175.440 38.560 ;
        RECT 175.520 38.240 175.840 38.560 ;
        RECT 175.920 38.240 176.240 38.560 ;
        RECT 176.320 38.240 176.640 38.560 ;
        RECT 176.720 38.240 177.040 38.560 ;
        RECT 177.120 38.240 177.440 38.560 ;
        RECT 177.520 38.240 177.840 38.560 ;
        RECT 177.920 38.240 178.240 38.560 ;
        RECT 178.320 38.240 178.640 38.560 ;
        RECT 178.720 38.240 179.040 38.560 ;
        RECT 179.120 38.240 179.440 38.560 ;
        RECT 179.520 38.240 179.840 38.560 ;
        RECT 179.920 38.240 180.240 38.560 ;
        RECT 180.320 38.240 180.640 38.560 ;
        RECT 25.040 37.840 25.360 38.160 ;
        RECT 25.440 37.840 25.760 38.160 ;
        RECT 25.840 37.840 26.160 38.160 ;
        RECT 26.240 37.840 26.560 38.160 ;
        RECT 26.640 37.840 26.960 38.160 ;
        RECT 27.040 37.840 27.360 38.160 ;
        RECT 27.440 37.840 27.760 38.160 ;
        RECT 27.840 37.840 28.160 38.160 ;
        RECT 28.240 37.840 28.560 38.160 ;
        RECT 28.640 37.840 28.960 38.160 ;
        RECT 29.040 37.840 29.360 38.160 ;
        RECT 29.440 37.840 29.760 38.160 ;
        RECT 29.840 37.840 30.160 38.160 ;
        RECT 30.240 37.840 30.560 38.160 ;
        RECT 30.640 37.840 30.960 38.160 ;
        RECT 31.040 37.840 31.360 38.160 ;
        RECT 31.440 37.840 31.760 38.160 ;
        RECT 31.840 37.840 32.160 38.160 ;
        RECT 32.240 37.840 32.560 38.160 ;
        RECT 32.640 37.840 32.960 38.160 ;
        RECT 33.040 37.840 33.360 38.160 ;
        RECT 33.440 37.840 33.760 38.160 ;
        RECT 33.840 37.840 34.160 38.160 ;
        RECT 34.240 37.840 34.560 38.160 ;
        RECT 34.640 37.840 34.960 38.160 ;
        RECT 35.040 37.840 35.360 38.160 ;
        RECT 35.440 37.840 35.760 38.160 ;
        RECT 35.840 37.840 36.160 38.160 ;
        RECT 36.240 37.840 36.560 38.160 ;
        RECT 36.640 37.840 36.960 38.160 ;
        RECT 37.040 37.840 37.360 38.160 ;
        RECT 37.440 37.840 37.760 38.160 ;
        RECT 37.840 37.840 38.160 38.160 ;
        RECT 38.240 37.840 38.560 38.160 ;
        RECT 38.640 37.840 38.960 38.160 ;
        RECT 39.040 37.840 39.360 38.160 ;
        RECT 39.440 37.840 39.760 38.160 ;
        RECT 39.840 37.840 40.160 38.160 ;
        RECT 40.240 37.840 40.560 38.160 ;
        RECT 40.640 37.840 40.960 38.160 ;
        RECT 41.040 37.840 41.360 38.160 ;
        RECT 41.440 37.840 41.760 38.160 ;
        RECT 41.840 37.840 42.160 38.160 ;
        RECT 42.240 37.840 42.560 38.160 ;
        RECT 42.640 37.840 42.960 38.160 ;
        RECT 43.040 37.840 43.360 38.160 ;
        RECT 43.440 37.840 43.760 38.160 ;
        RECT 43.840 37.840 44.160 38.160 ;
        RECT 44.240 37.840 44.560 38.160 ;
        RECT 44.640 37.840 44.960 38.160 ;
        RECT 70.560 37.840 70.880 38.160 ;
        RECT 70.960 37.840 71.280 38.160 ;
        RECT 71.360 37.840 71.680 38.160 ;
        RECT 71.760 37.840 72.080 38.160 ;
        RECT 120.560 37.840 120.880 38.160 ;
        RECT 120.960 37.840 121.280 38.160 ;
        RECT 121.360 37.840 121.680 38.160 ;
        RECT 121.760 37.840 122.080 38.160 ;
        RECT 160.720 37.840 161.040 38.160 ;
        RECT 161.120 37.840 161.440 38.160 ;
        RECT 161.520 37.840 161.840 38.160 ;
        RECT 161.920 37.840 162.240 38.160 ;
        RECT 162.320 37.840 162.640 38.160 ;
        RECT 162.720 37.840 163.040 38.160 ;
        RECT 163.120 37.840 163.440 38.160 ;
        RECT 163.520 37.840 163.840 38.160 ;
        RECT 163.920 37.840 164.240 38.160 ;
        RECT 164.320 37.840 164.640 38.160 ;
        RECT 164.720 37.840 165.040 38.160 ;
        RECT 165.120 37.840 165.440 38.160 ;
        RECT 165.520 37.840 165.840 38.160 ;
        RECT 165.920 37.840 166.240 38.160 ;
        RECT 166.320 37.840 166.640 38.160 ;
        RECT 166.720 37.840 167.040 38.160 ;
        RECT 167.120 37.840 167.440 38.160 ;
        RECT 167.520 37.840 167.840 38.160 ;
        RECT 167.920 37.840 168.240 38.160 ;
        RECT 168.320 37.840 168.640 38.160 ;
        RECT 168.720 37.840 169.040 38.160 ;
        RECT 169.120 37.840 169.440 38.160 ;
        RECT 169.520 37.840 169.840 38.160 ;
        RECT 169.920 37.840 170.240 38.160 ;
        RECT 170.320 37.840 170.640 38.160 ;
        RECT 170.720 37.840 171.040 38.160 ;
        RECT 171.120 37.840 171.440 38.160 ;
        RECT 171.520 37.840 171.840 38.160 ;
        RECT 171.920 37.840 172.240 38.160 ;
        RECT 172.320 37.840 172.640 38.160 ;
        RECT 172.720 37.840 173.040 38.160 ;
        RECT 173.120 37.840 173.440 38.160 ;
        RECT 173.520 37.840 173.840 38.160 ;
        RECT 173.920 37.840 174.240 38.160 ;
        RECT 174.320 37.840 174.640 38.160 ;
        RECT 174.720 37.840 175.040 38.160 ;
        RECT 175.120 37.840 175.440 38.160 ;
        RECT 175.520 37.840 175.840 38.160 ;
        RECT 175.920 37.840 176.240 38.160 ;
        RECT 176.320 37.840 176.640 38.160 ;
        RECT 176.720 37.840 177.040 38.160 ;
        RECT 177.120 37.840 177.440 38.160 ;
        RECT 177.520 37.840 177.840 38.160 ;
        RECT 177.920 37.840 178.240 38.160 ;
        RECT 178.320 37.840 178.640 38.160 ;
        RECT 178.720 37.840 179.040 38.160 ;
        RECT 179.120 37.840 179.440 38.160 ;
        RECT 179.520 37.840 179.840 38.160 ;
        RECT 179.920 37.840 180.240 38.160 ;
        RECT 180.320 37.840 180.640 38.160 ;
        RECT 25.040 37.440 25.360 37.760 ;
        RECT 25.440 37.440 25.760 37.760 ;
        RECT 25.840 37.440 26.160 37.760 ;
        RECT 26.240 37.440 26.560 37.760 ;
        RECT 26.640 37.440 26.960 37.760 ;
        RECT 27.040 37.440 27.360 37.760 ;
        RECT 27.440 37.440 27.760 37.760 ;
        RECT 27.840 37.440 28.160 37.760 ;
        RECT 28.240 37.440 28.560 37.760 ;
        RECT 28.640 37.440 28.960 37.760 ;
        RECT 29.040 37.440 29.360 37.760 ;
        RECT 29.440 37.440 29.760 37.760 ;
        RECT 29.840 37.440 30.160 37.760 ;
        RECT 30.240 37.440 30.560 37.760 ;
        RECT 30.640 37.440 30.960 37.760 ;
        RECT 31.040 37.440 31.360 37.760 ;
        RECT 31.440 37.440 31.760 37.760 ;
        RECT 31.840 37.440 32.160 37.760 ;
        RECT 32.240 37.440 32.560 37.760 ;
        RECT 32.640 37.440 32.960 37.760 ;
        RECT 33.040 37.440 33.360 37.760 ;
        RECT 33.440 37.440 33.760 37.760 ;
        RECT 33.840 37.440 34.160 37.760 ;
        RECT 34.240 37.440 34.560 37.760 ;
        RECT 34.640 37.440 34.960 37.760 ;
        RECT 35.040 37.440 35.360 37.760 ;
        RECT 35.440 37.440 35.760 37.760 ;
        RECT 35.840 37.440 36.160 37.760 ;
        RECT 36.240 37.440 36.560 37.760 ;
        RECT 36.640 37.440 36.960 37.760 ;
        RECT 37.040 37.440 37.360 37.760 ;
        RECT 37.440 37.440 37.760 37.760 ;
        RECT 37.840 37.440 38.160 37.760 ;
        RECT 38.240 37.440 38.560 37.760 ;
        RECT 38.640 37.440 38.960 37.760 ;
        RECT 39.040 37.440 39.360 37.760 ;
        RECT 39.440 37.440 39.760 37.760 ;
        RECT 39.840 37.440 40.160 37.760 ;
        RECT 40.240 37.440 40.560 37.760 ;
        RECT 40.640 37.440 40.960 37.760 ;
        RECT 41.040 37.440 41.360 37.760 ;
        RECT 41.440 37.440 41.760 37.760 ;
        RECT 41.840 37.440 42.160 37.760 ;
        RECT 42.240 37.440 42.560 37.760 ;
        RECT 42.640 37.440 42.960 37.760 ;
        RECT 43.040 37.440 43.360 37.760 ;
        RECT 43.440 37.440 43.760 37.760 ;
        RECT 43.840 37.440 44.160 37.760 ;
        RECT 44.240 37.440 44.560 37.760 ;
        RECT 44.640 37.440 44.960 37.760 ;
        RECT 70.560 37.440 70.880 37.760 ;
        RECT 70.960 37.440 71.280 37.760 ;
        RECT 71.360 37.440 71.680 37.760 ;
        RECT 71.760 37.440 72.080 37.760 ;
        RECT 120.560 37.440 120.880 37.760 ;
        RECT 120.960 37.440 121.280 37.760 ;
        RECT 121.360 37.440 121.680 37.760 ;
        RECT 121.760 37.440 122.080 37.760 ;
        RECT 160.720 37.440 161.040 37.760 ;
        RECT 161.120 37.440 161.440 37.760 ;
        RECT 161.520 37.440 161.840 37.760 ;
        RECT 161.920 37.440 162.240 37.760 ;
        RECT 162.320 37.440 162.640 37.760 ;
        RECT 162.720 37.440 163.040 37.760 ;
        RECT 163.120 37.440 163.440 37.760 ;
        RECT 163.520 37.440 163.840 37.760 ;
        RECT 163.920 37.440 164.240 37.760 ;
        RECT 164.320 37.440 164.640 37.760 ;
        RECT 164.720 37.440 165.040 37.760 ;
        RECT 165.120 37.440 165.440 37.760 ;
        RECT 165.520 37.440 165.840 37.760 ;
        RECT 165.920 37.440 166.240 37.760 ;
        RECT 166.320 37.440 166.640 37.760 ;
        RECT 166.720 37.440 167.040 37.760 ;
        RECT 167.120 37.440 167.440 37.760 ;
        RECT 167.520 37.440 167.840 37.760 ;
        RECT 167.920 37.440 168.240 37.760 ;
        RECT 168.320 37.440 168.640 37.760 ;
        RECT 168.720 37.440 169.040 37.760 ;
        RECT 169.120 37.440 169.440 37.760 ;
        RECT 169.520 37.440 169.840 37.760 ;
        RECT 169.920 37.440 170.240 37.760 ;
        RECT 170.320 37.440 170.640 37.760 ;
        RECT 170.720 37.440 171.040 37.760 ;
        RECT 171.120 37.440 171.440 37.760 ;
        RECT 171.520 37.440 171.840 37.760 ;
        RECT 171.920 37.440 172.240 37.760 ;
        RECT 172.320 37.440 172.640 37.760 ;
        RECT 172.720 37.440 173.040 37.760 ;
        RECT 173.120 37.440 173.440 37.760 ;
        RECT 173.520 37.440 173.840 37.760 ;
        RECT 173.920 37.440 174.240 37.760 ;
        RECT 174.320 37.440 174.640 37.760 ;
        RECT 174.720 37.440 175.040 37.760 ;
        RECT 175.120 37.440 175.440 37.760 ;
        RECT 175.520 37.440 175.840 37.760 ;
        RECT 175.920 37.440 176.240 37.760 ;
        RECT 176.320 37.440 176.640 37.760 ;
        RECT 176.720 37.440 177.040 37.760 ;
        RECT 177.120 37.440 177.440 37.760 ;
        RECT 177.520 37.440 177.840 37.760 ;
        RECT 177.920 37.440 178.240 37.760 ;
        RECT 178.320 37.440 178.640 37.760 ;
        RECT 178.720 37.440 179.040 37.760 ;
        RECT 179.120 37.440 179.440 37.760 ;
        RECT 179.520 37.440 179.840 37.760 ;
        RECT 179.920 37.440 180.240 37.760 ;
        RECT 180.320 37.440 180.640 37.760 ;
        RECT 25.040 37.040 25.360 37.360 ;
        RECT 25.440 37.040 25.760 37.360 ;
        RECT 25.840 37.040 26.160 37.360 ;
        RECT 26.240 37.040 26.560 37.360 ;
        RECT 26.640 37.040 26.960 37.360 ;
        RECT 27.040 37.040 27.360 37.360 ;
        RECT 27.440 37.040 27.760 37.360 ;
        RECT 27.840 37.040 28.160 37.360 ;
        RECT 28.240 37.040 28.560 37.360 ;
        RECT 28.640 37.040 28.960 37.360 ;
        RECT 29.040 37.040 29.360 37.360 ;
        RECT 29.440 37.040 29.760 37.360 ;
        RECT 29.840 37.040 30.160 37.360 ;
        RECT 30.240 37.040 30.560 37.360 ;
        RECT 30.640 37.040 30.960 37.360 ;
        RECT 31.040 37.040 31.360 37.360 ;
        RECT 31.440 37.040 31.760 37.360 ;
        RECT 31.840 37.040 32.160 37.360 ;
        RECT 32.240 37.040 32.560 37.360 ;
        RECT 32.640 37.040 32.960 37.360 ;
        RECT 33.040 37.040 33.360 37.360 ;
        RECT 33.440 37.040 33.760 37.360 ;
        RECT 33.840 37.040 34.160 37.360 ;
        RECT 34.240 37.040 34.560 37.360 ;
        RECT 34.640 37.040 34.960 37.360 ;
        RECT 35.040 37.040 35.360 37.360 ;
        RECT 35.440 37.040 35.760 37.360 ;
        RECT 35.840 37.040 36.160 37.360 ;
        RECT 36.240 37.040 36.560 37.360 ;
        RECT 36.640 37.040 36.960 37.360 ;
        RECT 37.040 37.040 37.360 37.360 ;
        RECT 37.440 37.040 37.760 37.360 ;
        RECT 37.840 37.040 38.160 37.360 ;
        RECT 38.240 37.040 38.560 37.360 ;
        RECT 38.640 37.040 38.960 37.360 ;
        RECT 39.040 37.040 39.360 37.360 ;
        RECT 39.440 37.040 39.760 37.360 ;
        RECT 39.840 37.040 40.160 37.360 ;
        RECT 40.240 37.040 40.560 37.360 ;
        RECT 40.640 37.040 40.960 37.360 ;
        RECT 41.040 37.040 41.360 37.360 ;
        RECT 41.440 37.040 41.760 37.360 ;
        RECT 41.840 37.040 42.160 37.360 ;
        RECT 42.240 37.040 42.560 37.360 ;
        RECT 42.640 37.040 42.960 37.360 ;
        RECT 43.040 37.040 43.360 37.360 ;
        RECT 43.440 37.040 43.760 37.360 ;
        RECT 43.840 37.040 44.160 37.360 ;
        RECT 44.240 37.040 44.560 37.360 ;
        RECT 44.640 37.040 44.960 37.360 ;
        RECT 70.560 37.040 70.880 37.360 ;
        RECT 70.960 37.040 71.280 37.360 ;
        RECT 71.360 37.040 71.680 37.360 ;
        RECT 71.760 37.040 72.080 37.360 ;
        RECT 120.560 37.040 120.880 37.360 ;
        RECT 120.960 37.040 121.280 37.360 ;
        RECT 121.360 37.040 121.680 37.360 ;
        RECT 121.760 37.040 122.080 37.360 ;
        RECT 160.720 37.040 161.040 37.360 ;
        RECT 161.120 37.040 161.440 37.360 ;
        RECT 161.520 37.040 161.840 37.360 ;
        RECT 161.920 37.040 162.240 37.360 ;
        RECT 162.320 37.040 162.640 37.360 ;
        RECT 162.720 37.040 163.040 37.360 ;
        RECT 163.120 37.040 163.440 37.360 ;
        RECT 163.520 37.040 163.840 37.360 ;
        RECT 163.920 37.040 164.240 37.360 ;
        RECT 164.320 37.040 164.640 37.360 ;
        RECT 164.720 37.040 165.040 37.360 ;
        RECT 165.120 37.040 165.440 37.360 ;
        RECT 165.520 37.040 165.840 37.360 ;
        RECT 165.920 37.040 166.240 37.360 ;
        RECT 166.320 37.040 166.640 37.360 ;
        RECT 166.720 37.040 167.040 37.360 ;
        RECT 167.120 37.040 167.440 37.360 ;
        RECT 167.520 37.040 167.840 37.360 ;
        RECT 167.920 37.040 168.240 37.360 ;
        RECT 168.320 37.040 168.640 37.360 ;
        RECT 168.720 37.040 169.040 37.360 ;
        RECT 169.120 37.040 169.440 37.360 ;
        RECT 169.520 37.040 169.840 37.360 ;
        RECT 169.920 37.040 170.240 37.360 ;
        RECT 170.320 37.040 170.640 37.360 ;
        RECT 170.720 37.040 171.040 37.360 ;
        RECT 171.120 37.040 171.440 37.360 ;
        RECT 171.520 37.040 171.840 37.360 ;
        RECT 171.920 37.040 172.240 37.360 ;
        RECT 172.320 37.040 172.640 37.360 ;
        RECT 172.720 37.040 173.040 37.360 ;
        RECT 173.120 37.040 173.440 37.360 ;
        RECT 173.520 37.040 173.840 37.360 ;
        RECT 173.920 37.040 174.240 37.360 ;
        RECT 174.320 37.040 174.640 37.360 ;
        RECT 174.720 37.040 175.040 37.360 ;
        RECT 175.120 37.040 175.440 37.360 ;
        RECT 175.520 37.040 175.840 37.360 ;
        RECT 175.920 37.040 176.240 37.360 ;
        RECT 176.320 37.040 176.640 37.360 ;
        RECT 176.720 37.040 177.040 37.360 ;
        RECT 177.120 37.040 177.440 37.360 ;
        RECT 177.520 37.040 177.840 37.360 ;
        RECT 177.920 37.040 178.240 37.360 ;
        RECT 178.320 37.040 178.640 37.360 ;
        RECT 178.720 37.040 179.040 37.360 ;
        RECT 179.120 37.040 179.440 37.360 ;
        RECT 179.520 37.040 179.840 37.360 ;
        RECT 179.920 37.040 180.240 37.360 ;
        RECT 180.320 37.040 180.640 37.360 ;
        RECT 25.040 36.640 25.360 36.960 ;
        RECT 25.440 36.640 25.760 36.960 ;
        RECT 25.840 36.640 26.160 36.960 ;
        RECT 26.240 36.640 26.560 36.960 ;
        RECT 26.640 36.640 26.960 36.960 ;
        RECT 27.040 36.640 27.360 36.960 ;
        RECT 27.440 36.640 27.760 36.960 ;
        RECT 27.840 36.640 28.160 36.960 ;
        RECT 28.240 36.640 28.560 36.960 ;
        RECT 28.640 36.640 28.960 36.960 ;
        RECT 29.040 36.640 29.360 36.960 ;
        RECT 29.440 36.640 29.760 36.960 ;
        RECT 29.840 36.640 30.160 36.960 ;
        RECT 30.240 36.640 30.560 36.960 ;
        RECT 30.640 36.640 30.960 36.960 ;
        RECT 31.040 36.640 31.360 36.960 ;
        RECT 31.440 36.640 31.760 36.960 ;
        RECT 31.840 36.640 32.160 36.960 ;
        RECT 32.240 36.640 32.560 36.960 ;
        RECT 32.640 36.640 32.960 36.960 ;
        RECT 33.040 36.640 33.360 36.960 ;
        RECT 33.440 36.640 33.760 36.960 ;
        RECT 33.840 36.640 34.160 36.960 ;
        RECT 34.240 36.640 34.560 36.960 ;
        RECT 34.640 36.640 34.960 36.960 ;
        RECT 35.040 36.640 35.360 36.960 ;
        RECT 35.440 36.640 35.760 36.960 ;
        RECT 35.840 36.640 36.160 36.960 ;
        RECT 36.240 36.640 36.560 36.960 ;
        RECT 36.640 36.640 36.960 36.960 ;
        RECT 37.040 36.640 37.360 36.960 ;
        RECT 37.440 36.640 37.760 36.960 ;
        RECT 37.840 36.640 38.160 36.960 ;
        RECT 38.240 36.640 38.560 36.960 ;
        RECT 38.640 36.640 38.960 36.960 ;
        RECT 39.040 36.640 39.360 36.960 ;
        RECT 39.440 36.640 39.760 36.960 ;
        RECT 39.840 36.640 40.160 36.960 ;
        RECT 40.240 36.640 40.560 36.960 ;
        RECT 40.640 36.640 40.960 36.960 ;
        RECT 41.040 36.640 41.360 36.960 ;
        RECT 41.440 36.640 41.760 36.960 ;
        RECT 41.840 36.640 42.160 36.960 ;
        RECT 42.240 36.640 42.560 36.960 ;
        RECT 42.640 36.640 42.960 36.960 ;
        RECT 43.040 36.640 43.360 36.960 ;
        RECT 43.440 36.640 43.760 36.960 ;
        RECT 43.840 36.640 44.160 36.960 ;
        RECT 44.240 36.640 44.560 36.960 ;
        RECT 44.640 36.640 44.960 36.960 ;
        RECT 70.560 36.640 70.880 36.960 ;
        RECT 70.960 36.640 71.280 36.960 ;
        RECT 71.360 36.640 71.680 36.960 ;
        RECT 71.760 36.640 72.080 36.960 ;
        RECT 120.560 36.640 120.880 36.960 ;
        RECT 120.960 36.640 121.280 36.960 ;
        RECT 121.360 36.640 121.680 36.960 ;
        RECT 121.760 36.640 122.080 36.960 ;
        RECT 160.720 36.640 161.040 36.960 ;
        RECT 161.120 36.640 161.440 36.960 ;
        RECT 161.520 36.640 161.840 36.960 ;
        RECT 161.920 36.640 162.240 36.960 ;
        RECT 162.320 36.640 162.640 36.960 ;
        RECT 162.720 36.640 163.040 36.960 ;
        RECT 163.120 36.640 163.440 36.960 ;
        RECT 163.520 36.640 163.840 36.960 ;
        RECT 163.920 36.640 164.240 36.960 ;
        RECT 164.320 36.640 164.640 36.960 ;
        RECT 164.720 36.640 165.040 36.960 ;
        RECT 165.120 36.640 165.440 36.960 ;
        RECT 165.520 36.640 165.840 36.960 ;
        RECT 165.920 36.640 166.240 36.960 ;
        RECT 166.320 36.640 166.640 36.960 ;
        RECT 166.720 36.640 167.040 36.960 ;
        RECT 167.120 36.640 167.440 36.960 ;
        RECT 167.520 36.640 167.840 36.960 ;
        RECT 167.920 36.640 168.240 36.960 ;
        RECT 168.320 36.640 168.640 36.960 ;
        RECT 168.720 36.640 169.040 36.960 ;
        RECT 169.120 36.640 169.440 36.960 ;
        RECT 169.520 36.640 169.840 36.960 ;
        RECT 169.920 36.640 170.240 36.960 ;
        RECT 170.320 36.640 170.640 36.960 ;
        RECT 170.720 36.640 171.040 36.960 ;
        RECT 171.120 36.640 171.440 36.960 ;
        RECT 171.520 36.640 171.840 36.960 ;
        RECT 171.920 36.640 172.240 36.960 ;
        RECT 172.320 36.640 172.640 36.960 ;
        RECT 172.720 36.640 173.040 36.960 ;
        RECT 173.120 36.640 173.440 36.960 ;
        RECT 173.520 36.640 173.840 36.960 ;
        RECT 173.920 36.640 174.240 36.960 ;
        RECT 174.320 36.640 174.640 36.960 ;
        RECT 174.720 36.640 175.040 36.960 ;
        RECT 175.120 36.640 175.440 36.960 ;
        RECT 175.520 36.640 175.840 36.960 ;
        RECT 175.920 36.640 176.240 36.960 ;
        RECT 176.320 36.640 176.640 36.960 ;
        RECT 176.720 36.640 177.040 36.960 ;
        RECT 177.120 36.640 177.440 36.960 ;
        RECT 177.520 36.640 177.840 36.960 ;
        RECT 177.920 36.640 178.240 36.960 ;
        RECT 178.320 36.640 178.640 36.960 ;
        RECT 178.720 36.640 179.040 36.960 ;
        RECT 179.120 36.640 179.440 36.960 ;
        RECT 179.520 36.640 179.840 36.960 ;
        RECT 179.920 36.640 180.240 36.960 ;
        RECT 180.320 36.640 180.640 36.960 ;
        RECT 25.040 36.240 25.360 36.560 ;
        RECT 25.440 36.240 25.760 36.560 ;
        RECT 25.840 36.240 26.160 36.560 ;
        RECT 26.240 36.240 26.560 36.560 ;
        RECT 26.640 36.240 26.960 36.560 ;
        RECT 27.040 36.240 27.360 36.560 ;
        RECT 27.440 36.240 27.760 36.560 ;
        RECT 27.840 36.240 28.160 36.560 ;
        RECT 28.240 36.240 28.560 36.560 ;
        RECT 28.640 36.240 28.960 36.560 ;
        RECT 29.040 36.240 29.360 36.560 ;
        RECT 29.440 36.240 29.760 36.560 ;
        RECT 29.840 36.240 30.160 36.560 ;
        RECT 30.240 36.240 30.560 36.560 ;
        RECT 30.640 36.240 30.960 36.560 ;
        RECT 31.040 36.240 31.360 36.560 ;
        RECT 31.440 36.240 31.760 36.560 ;
        RECT 31.840 36.240 32.160 36.560 ;
        RECT 32.240 36.240 32.560 36.560 ;
        RECT 32.640 36.240 32.960 36.560 ;
        RECT 33.040 36.240 33.360 36.560 ;
        RECT 33.440 36.240 33.760 36.560 ;
        RECT 33.840 36.240 34.160 36.560 ;
        RECT 34.240 36.240 34.560 36.560 ;
        RECT 34.640 36.240 34.960 36.560 ;
        RECT 35.040 36.240 35.360 36.560 ;
        RECT 35.440 36.240 35.760 36.560 ;
        RECT 35.840 36.240 36.160 36.560 ;
        RECT 36.240 36.240 36.560 36.560 ;
        RECT 36.640 36.240 36.960 36.560 ;
        RECT 37.040 36.240 37.360 36.560 ;
        RECT 37.440 36.240 37.760 36.560 ;
        RECT 37.840 36.240 38.160 36.560 ;
        RECT 38.240 36.240 38.560 36.560 ;
        RECT 38.640 36.240 38.960 36.560 ;
        RECT 39.040 36.240 39.360 36.560 ;
        RECT 39.440 36.240 39.760 36.560 ;
        RECT 39.840 36.240 40.160 36.560 ;
        RECT 40.240 36.240 40.560 36.560 ;
        RECT 40.640 36.240 40.960 36.560 ;
        RECT 41.040 36.240 41.360 36.560 ;
        RECT 41.440 36.240 41.760 36.560 ;
        RECT 41.840 36.240 42.160 36.560 ;
        RECT 42.240 36.240 42.560 36.560 ;
        RECT 42.640 36.240 42.960 36.560 ;
        RECT 43.040 36.240 43.360 36.560 ;
        RECT 43.440 36.240 43.760 36.560 ;
        RECT 43.840 36.240 44.160 36.560 ;
        RECT 44.240 36.240 44.560 36.560 ;
        RECT 44.640 36.240 44.960 36.560 ;
        RECT 70.560 36.240 70.880 36.560 ;
        RECT 70.960 36.240 71.280 36.560 ;
        RECT 71.360 36.240 71.680 36.560 ;
        RECT 71.760 36.240 72.080 36.560 ;
        RECT 120.560 36.240 120.880 36.560 ;
        RECT 120.960 36.240 121.280 36.560 ;
        RECT 121.360 36.240 121.680 36.560 ;
        RECT 121.760 36.240 122.080 36.560 ;
        RECT 160.720 36.240 161.040 36.560 ;
        RECT 161.120 36.240 161.440 36.560 ;
        RECT 161.520 36.240 161.840 36.560 ;
        RECT 161.920 36.240 162.240 36.560 ;
        RECT 162.320 36.240 162.640 36.560 ;
        RECT 162.720 36.240 163.040 36.560 ;
        RECT 163.120 36.240 163.440 36.560 ;
        RECT 163.520 36.240 163.840 36.560 ;
        RECT 163.920 36.240 164.240 36.560 ;
        RECT 164.320 36.240 164.640 36.560 ;
        RECT 164.720 36.240 165.040 36.560 ;
        RECT 165.120 36.240 165.440 36.560 ;
        RECT 165.520 36.240 165.840 36.560 ;
        RECT 165.920 36.240 166.240 36.560 ;
        RECT 166.320 36.240 166.640 36.560 ;
        RECT 166.720 36.240 167.040 36.560 ;
        RECT 167.120 36.240 167.440 36.560 ;
        RECT 167.520 36.240 167.840 36.560 ;
        RECT 167.920 36.240 168.240 36.560 ;
        RECT 168.320 36.240 168.640 36.560 ;
        RECT 168.720 36.240 169.040 36.560 ;
        RECT 169.120 36.240 169.440 36.560 ;
        RECT 169.520 36.240 169.840 36.560 ;
        RECT 169.920 36.240 170.240 36.560 ;
        RECT 170.320 36.240 170.640 36.560 ;
        RECT 170.720 36.240 171.040 36.560 ;
        RECT 171.120 36.240 171.440 36.560 ;
        RECT 171.520 36.240 171.840 36.560 ;
        RECT 171.920 36.240 172.240 36.560 ;
        RECT 172.320 36.240 172.640 36.560 ;
        RECT 172.720 36.240 173.040 36.560 ;
        RECT 173.120 36.240 173.440 36.560 ;
        RECT 173.520 36.240 173.840 36.560 ;
        RECT 173.920 36.240 174.240 36.560 ;
        RECT 174.320 36.240 174.640 36.560 ;
        RECT 174.720 36.240 175.040 36.560 ;
        RECT 175.120 36.240 175.440 36.560 ;
        RECT 175.520 36.240 175.840 36.560 ;
        RECT 175.920 36.240 176.240 36.560 ;
        RECT 176.320 36.240 176.640 36.560 ;
        RECT 176.720 36.240 177.040 36.560 ;
        RECT 177.120 36.240 177.440 36.560 ;
        RECT 177.520 36.240 177.840 36.560 ;
        RECT 177.920 36.240 178.240 36.560 ;
        RECT 178.320 36.240 178.640 36.560 ;
        RECT 178.720 36.240 179.040 36.560 ;
        RECT 179.120 36.240 179.440 36.560 ;
        RECT 179.520 36.240 179.840 36.560 ;
        RECT 179.920 36.240 180.240 36.560 ;
        RECT 180.320 36.240 180.640 36.560 ;
        RECT 25.040 35.840 25.360 36.160 ;
        RECT 25.440 35.840 25.760 36.160 ;
        RECT 25.840 35.840 26.160 36.160 ;
        RECT 26.240 35.840 26.560 36.160 ;
        RECT 26.640 35.840 26.960 36.160 ;
        RECT 27.040 35.840 27.360 36.160 ;
        RECT 27.440 35.840 27.760 36.160 ;
        RECT 27.840 35.840 28.160 36.160 ;
        RECT 28.240 35.840 28.560 36.160 ;
        RECT 28.640 35.840 28.960 36.160 ;
        RECT 29.040 35.840 29.360 36.160 ;
        RECT 29.440 35.840 29.760 36.160 ;
        RECT 29.840 35.840 30.160 36.160 ;
        RECT 30.240 35.840 30.560 36.160 ;
        RECT 30.640 35.840 30.960 36.160 ;
        RECT 31.040 35.840 31.360 36.160 ;
        RECT 31.440 35.840 31.760 36.160 ;
        RECT 31.840 35.840 32.160 36.160 ;
        RECT 32.240 35.840 32.560 36.160 ;
        RECT 32.640 35.840 32.960 36.160 ;
        RECT 33.040 35.840 33.360 36.160 ;
        RECT 33.440 35.840 33.760 36.160 ;
        RECT 33.840 35.840 34.160 36.160 ;
        RECT 34.240 35.840 34.560 36.160 ;
        RECT 34.640 35.840 34.960 36.160 ;
        RECT 35.040 35.840 35.360 36.160 ;
        RECT 35.440 35.840 35.760 36.160 ;
        RECT 35.840 35.840 36.160 36.160 ;
        RECT 36.240 35.840 36.560 36.160 ;
        RECT 36.640 35.840 36.960 36.160 ;
        RECT 37.040 35.840 37.360 36.160 ;
        RECT 37.440 35.840 37.760 36.160 ;
        RECT 37.840 35.840 38.160 36.160 ;
        RECT 38.240 35.840 38.560 36.160 ;
        RECT 38.640 35.840 38.960 36.160 ;
        RECT 39.040 35.840 39.360 36.160 ;
        RECT 39.440 35.840 39.760 36.160 ;
        RECT 39.840 35.840 40.160 36.160 ;
        RECT 40.240 35.840 40.560 36.160 ;
        RECT 40.640 35.840 40.960 36.160 ;
        RECT 41.040 35.840 41.360 36.160 ;
        RECT 41.440 35.840 41.760 36.160 ;
        RECT 41.840 35.840 42.160 36.160 ;
        RECT 42.240 35.840 42.560 36.160 ;
        RECT 42.640 35.840 42.960 36.160 ;
        RECT 43.040 35.840 43.360 36.160 ;
        RECT 43.440 35.840 43.760 36.160 ;
        RECT 43.840 35.840 44.160 36.160 ;
        RECT 44.240 35.840 44.560 36.160 ;
        RECT 44.640 35.840 44.960 36.160 ;
        RECT 70.560 35.840 70.880 36.160 ;
        RECT 70.960 35.840 71.280 36.160 ;
        RECT 71.360 35.840 71.680 36.160 ;
        RECT 71.760 35.840 72.080 36.160 ;
        RECT 120.560 35.840 120.880 36.160 ;
        RECT 120.960 35.840 121.280 36.160 ;
        RECT 121.360 35.840 121.680 36.160 ;
        RECT 121.760 35.840 122.080 36.160 ;
        RECT 160.720 35.840 161.040 36.160 ;
        RECT 161.120 35.840 161.440 36.160 ;
        RECT 161.520 35.840 161.840 36.160 ;
        RECT 161.920 35.840 162.240 36.160 ;
        RECT 162.320 35.840 162.640 36.160 ;
        RECT 162.720 35.840 163.040 36.160 ;
        RECT 163.120 35.840 163.440 36.160 ;
        RECT 163.520 35.840 163.840 36.160 ;
        RECT 163.920 35.840 164.240 36.160 ;
        RECT 164.320 35.840 164.640 36.160 ;
        RECT 164.720 35.840 165.040 36.160 ;
        RECT 165.120 35.840 165.440 36.160 ;
        RECT 165.520 35.840 165.840 36.160 ;
        RECT 165.920 35.840 166.240 36.160 ;
        RECT 166.320 35.840 166.640 36.160 ;
        RECT 166.720 35.840 167.040 36.160 ;
        RECT 167.120 35.840 167.440 36.160 ;
        RECT 167.520 35.840 167.840 36.160 ;
        RECT 167.920 35.840 168.240 36.160 ;
        RECT 168.320 35.840 168.640 36.160 ;
        RECT 168.720 35.840 169.040 36.160 ;
        RECT 169.120 35.840 169.440 36.160 ;
        RECT 169.520 35.840 169.840 36.160 ;
        RECT 169.920 35.840 170.240 36.160 ;
        RECT 170.320 35.840 170.640 36.160 ;
        RECT 170.720 35.840 171.040 36.160 ;
        RECT 171.120 35.840 171.440 36.160 ;
        RECT 171.520 35.840 171.840 36.160 ;
        RECT 171.920 35.840 172.240 36.160 ;
        RECT 172.320 35.840 172.640 36.160 ;
        RECT 172.720 35.840 173.040 36.160 ;
        RECT 173.120 35.840 173.440 36.160 ;
        RECT 173.520 35.840 173.840 36.160 ;
        RECT 173.920 35.840 174.240 36.160 ;
        RECT 174.320 35.840 174.640 36.160 ;
        RECT 174.720 35.840 175.040 36.160 ;
        RECT 175.120 35.840 175.440 36.160 ;
        RECT 175.520 35.840 175.840 36.160 ;
        RECT 175.920 35.840 176.240 36.160 ;
        RECT 176.320 35.840 176.640 36.160 ;
        RECT 176.720 35.840 177.040 36.160 ;
        RECT 177.120 35.840 177.440 36.160 ;
        RECT 177.520 35.840 177.840 36.160 ;
        RECT 177.920 35.840 178.240 36.160 ;
        RECT 178.320 35.840 178.640 36.160 ;
        RECT 178.720 35.840 179.040 36.160 ;
        RECT 179.120 35.840 179.440 36.160 ;
        RECT 179.520 35.840 179.840 36.160 ;
        RECT 179.920 35.840 180.240 36.160 ;
        RECT 180.320 35.840 180.640 36.160 ;
        RECT 25.040 35.440 25.360 35.760 ;
        RECT 25.440 35.440 25.760 35.760 ;
        RECT 25.840 35.440 26.160 35.760 ;
        RECT 26.240 35.440 26.560 35.760 ;
        RECT 26.640 35.440 26.960 35.760 ;
        RECT 27.040 35.440 27.360 35.760 ;
        RECT 27.440 35.440 27.760 35.760 ;
        RECT 27.840 35.440 28.160 35.760 ;
        RECT 28.240 35.440 28.560 35.760 ;
        RECT 28.640 35.440 28.960 35.760 ;
        RECT 29.040 35.440 29.360 35.760 ;
        RECT 29.440 35.440 29.760 35.760 ;
        RECT 29.840 35.440 30.160 35.760 ;
        RECT 30.240 35.440 30.560 35.760 ;
        RECT 30.640 35.440 30.960 35.760 ;
        RECT 31.040 35.440 31.360 35.760 ;
        RECT 31.440 35.440 31.760 35.760 ;
        RECT 31.840 35.440 32.160 35.760 ;
        RECT 32.240 35.440 32.560 35.760 ;
        RECT 32.640 35.440 32.960 35.760 ;
        RECT 33.040 35.440 33.360 35.760 ;
        RECT 33.440 35.440 33.760 35.760 ;
        RECT 33.840 35.440 34.160 35.760 ;
        RECT 34.240 35.440 34.560 35.760 ;
        RECT 34.640 35.440 34.960 35.760 ;
        RECT 35.040 35.440 35.360 35.760 ;
        RECT 35.440 35.440 35.760 35.760 ;
        RECT 35.840 35.440 36.160 35.760 ;
        RECT 36.240 35.440 36.560 35.760 ;
        RECT 36.640 35.440 36.960 35.760 ;
        RECT 37.040 35.440 37.360 35.760 ;
        RECT 37.440 35.440 37.760 35.760 ;
        RECT 37.840 35.440 38.160 35.760 ;
        RECT 38.240 35.440 38.560 35.760 ;
        RECT 38.640 35.440 38.960 35.760 ;
        RECT 39.040 35.440 39.360 35.760 ;
        RECT 39.440 35.440 39.760 35.760 ;
        RECT 39.840 35.440 40.160 35.760 ;
        RECT 40.240 35.440 40.560 35.760 ;
        RECT 40.640 35.440 40.960 35.760 ;
        RECT 41.040 35.440 41.360 35.760 ;
        RECT 41.440 35.440 41.760 35.760 ;
        RECT 41.840 35.440 42.160 35.760 ;
        RECT 42.240 35.440 42.560 35.760 ;
        RECT 42.640 35.440 42.960 35.760 ;
        RECT 43.040 35.440 43.360 35.760 ;
        RECT 43.440 35.440 43.760 35.760 ;
        RECT 43.840 35.440 44.160 35.760 ;
        RECT 44.240 35.440 44.560 35.760 ;
        RECT 44.640 35.440 44.960 35.760 ;
        RECT 70.560 35.440 70.880 35.760 ;
        RECT 70.960 35.440 71.280 35.760 ;
        RECT 71.360 35.440 71.680 35.760 ;
        RECT 71.760 35.440 72.080 35.760 ;
        RECT 120.560 35.440 120.880 35.760 ;
        RECT 120.960 35.440 121.280 35.760 ;
        RECT 121.360 35.440 121.680 35.760 ;
        RECT 121.760 35.440 122.080 35.760 ;
        RECT 160.720 35.440 161.040 35.760 ;
        RECT 161.120 35.440 161.440 35.760 ;
        RECT 161.520 35.440 161.840 35.760 ;
        RECT 161.920 35.440 162.240 35.760 ;
        RECT 162.320 35.440 162.640 35.760 ;
        RECT 162.720 35.440 163.040 35.760 ;
        RECT 163.120 35.440 163.440 35.760 ;
        RECT 163.520 35.440 163.840 35.760 ;
        RECT 163.920 35.440 164.240 35.760 ;
        RECT 164.320 35.440 164.640 35.760 ;
        RECT 164.720 35.440 165.040 35.760 ;
        RECT 165.120 35.440 165.440 35.760 ;
        RECT 165.520 35.440 165.840 35.760 ;
        RECT 165.920 35.440 166.240 35.760 ;
        RECT 166.320 35.440 166.640 35.760 ;
        RECT 166.720 35.440 167.040 35.760 ;
        RECT 167.120 35.440 167.440 35.760 ;
        RECT 167.520 35.440 167.840 35.760 ;
        RECT 167.920 35.440 168.240 35.760 ;
        RECT 168.320 35.440 168.640 35.760 ;
        RECT 168.720 35.440 169.040 35.760 ;
        RECT 169.120 35.440 169.440 35.760 ;
        RECT 169.520 35.440 169.840 35.760 ;
        RECT 169.920 35.440 170.240 35.760 ;
        RECT 170.320 35.440 170.640 35.760 ;
        RECT 170.720 35.440 171.040 35.760 ;
        RECT 171.120 35.440 171.440 35.760 ;
        RECT 171.520 35.440 171.840 35.760 ;
        RECT 171.920 35.440 172.240 35.760 ;
        RECT 172.320 35.440 172.640 35.760 ;
        RECT 172.720 35.440 173.040 35.760 ;
        RECT 173.120 35.440 173.440 35.760 ;
        RECT 173.520 35.440 173.840 35.760 ;
        RECT 173.920 35.440 174.240 35.760 ;
        RECT 174.320 35.440 174.640 35.760 ;
        RECT 174.720 35.440 175.040 35.760 ;
        RECT 175.120 35.440 175.440 35.760 ;
        RECT 175.520 35.440 175.840 35.760 ;
        RECT 175.920 35.440 176.240 35.760 ;
        RECT 176.320 35.440 176.640 35.760 ;
        RECT 176.720 35.440 177.040 35.760 ;
        RECT 177.120 35.440 177.440 35.760 ;
        RECT 177.520 35.440 177.840 35.760 ;
        RECT 177.920 35.440 178.240 35.760 ;
        RECT 178.320 35.440 178.640 35.760 ;
        RECT 178.720 35.440 179.040 35.760 ;
        RECT 179.120 35.440 179.440 35.760 ;
        RECT 179.520 35.440 179.840 35.760 ;
        RECT 179.920 35.440 180.240 35.760 ;
        RECT 180.320 35.440 180.640 35.760 ;
        RECT 25.040 35.040 25.360 35.360 ;
        RECT 25.440 35.040 25.760 35.360 ;
        RECT 25.840 35.040 26.160 35.360 ;
        RECT 26.240 35.040 26.560 35.360 ;
        RECT 26.640 35.040 26.960 35.360 ;
        RECT 27.040 35.040 27.360 35.360 ;
        RECT 27.440 35.040 27.760 35.360 ;
        RECT 27.840 35.040 28.160 35.360 ;
        RECT 28.240 35.040 28.560 35.360 ;
        RECT 28.640 35.040 28.960 35.360 ;
        RECT 29.040 35.040 29.360 35.360 ;
        RECT 29.440 35.040 29.760 35.360 ;
        RECT 29.840 35.040 30.160 35.360 ;
        RECT 30.240 35.040 30.560 35.360 ;
        RECT 30.640 35.040 30.960 35.360 ;
        RECT 31.040 35.040 31.360 35.360 ;
        RECT 31.440 35.040 31.760 35.360 ;
        RECT 31.840 35.040 32.160 35.360 ;
        RECT 32.240 35.040 32.560 35.360 ;
        RECT 32.640 35.040 32.960 35.360 ;
        RECT 33.040 35.040 33.360 35.360 ;
        RECT 33.440 35.040 33.760 35.360 ;
        RECT 33.840 35.040 34.160 35.360 ;
        RECT 34.240 35.040 34.560 35.360 ;
        RECT 34.640 35.040 34.960 35.360 ;
        RECT 35.040 35.040 35.360 35.360 ;
        RECT 35.440 35.040 35.760 35.360 ;
        RECT 35.840 35.040 36.160 35.360 ;
        RECT 36.240 35.040 36.560 35.360 ;
        RECT 36.640 35.040 36.960 35.360 ;
        RECT 37.040 35.040 37.360 35.360 ;
        RECT 37.440 35.040 37.760 35.360 ;
        RECT 37.840 35.040 38.160 35.360 ;
        RECT 38.240 35.040 38.560 35.360 ;
        RECT 38.640 35.040 38.960 35.360 ;
        RECT 39.040 35.040 39.360 35.360 ;
        RECT 39.440 35.040 39.760 35.360 ;
        RECT 39.840 35.040 40.160 35.360 ;
        RECT 40.240 35.040 40.560 35.360 ;
        RECT 40.640 35.040 40.960 35.360 ;
        RECT 41.040 35.040 41.360 35.360 ;
        RECT 41.440 35.040 41.760 35.360 ;
        RECT 41.840 35.040 42.160 35.360 ;
        RECT 42.240 35.040 42.560 35.360 ;
        RECT 42.640 35.040 42.960 35.360 ;
        RECT 43.040 35.040 43.360 35.360 ;
        RECT 43.440 35.040 43.760 35.360 ;
        RECT 43.840 35.040 44.160 35.360 ;
        RECT 44.240 35.040 44.560 35.360 ;
        RECT 44.640 35.040 44.960 35.360 ;
        RECT 70.560 35.040 70.880 35.360 ;
        RECT 70.960 35.040 71.280 35.360 ;
        RECT 71.360 35.040 71.680 35.360 ;
        RECT 71.760 35.040 72.080 35.360 ;
        RECT 120.560 35.040 120.880 35.360 ;
        RECT 120.960 35.040 121.280 35.360 ;
        RECT 121.360 35.040 121.680 35.360 ;
        RECT 121.760 35.040 122.080 35.360 ;
        RECT 160.720 35.040 161.040 35.360 ;
        RECT 161.120 35.040 161.440 35.360 ;
        RECT 161.520 35.040 161.840 35.360 ;
        RECT 161.920 35.040 162.240 35.360 ;
        RECT 162.320 35.040 162.640 35.360 ;
        RECT 162.720 35.040 163.040 35.360 ;
        RECT 163.120 35.040 163.440 35.360 ;
        RECT 163.520 35.040 163.840 35.360 ;
        RECT 163.920 35.040 164.240 35.360 ;
        RECT 164.320 35.040 164.640 35.360 ;
        RECT 164.720 35.040 165.040 35.360 ;
        RECT 165.120 35.040 165.440 35.360 ;
        RECT 165.520 35.040 165.840 35.360 ;
        RECT 165.920 35.040 166.240 35.360 ;
        RECT 166.320 35.040 166.640 35.360 ;
        RECT 166.720 35.040 167.040 35.360 ;
        RECT 167.120 35.040 167.440 35.360 ;
        RECT 167.520 35.040 167.840 35.360 ;
        RECT 167.920 35.040 168.240 35.360 ;
        RECT 168.320 35.040 168.640 35.360 ;
        RECT 168.720 35.040 169.040 35.360 ;
        RECT 169.120 35.040 169.440 35.360 ;
        RECT 169.520 35.040 169.840 35.360 ;
        RECT 169.920 35.040 170.240 35.360 ;
        RECT 170.320 35.040 170.640 35.360 ;
        RECT 170.720 35.040 171.040 35.360 ;
        RECT 171.120 35.040 171.440 35.360 ;
        RECT 171.520 35.040 171.840 35.360 ;
        RECT 171.920 35.040 172.240 35.360 ;
        RECT 172.320 35.040 172.640 35.360 ;
        RECT 172.720 35.040 173.040 35.360 ;
        RECT 173.120 35.040 173.440 35.360 ;
        RECT 173.520 35.040 173.840 35.360 ;
        RECT 173.920 35.040 174.240 35.360 ;
        RECT 174.320 35.040 174.640 35.360 ;
        RECT 174.720 35.040 175.040 35.360 ;
        RECT 175.120 35.040 175.440 35.360 ;
        RECT 175.520 35.040 175.840 35.360 ;
        RECT 175.920 35.040 176.240 35.360 ;
        RECT 176.320 35.040 176.640 35.360 ;
        RECT 176.720 35.040 177.040 35.360 ;
        RECT 177.120 35.040 177.440 35.360 ;
        RECT 177.520 35.040 177.840 35.360 ;
        RECT 177.920 35.040 178.240 35.360 ;
        RECT 178.320 35.040 178.640 35.360 ;
        RECT 178.720 35.040 179.040 35.360 ;
        RECT 179.120 35.040 179.440 35.360 ;
        RECT 179.520 35.040 179.840 35.360 ;
        RECT 179.920 35.040 180.240 35.360 ;
        RECT 180.320 35.040 180.640 35.360 ;
        RECT 25.040 34.640 25.360 34.960 ;
        RECT 25.440 34.640 25.760 34.960 ;
        RECT 25.840 34.640 26.160 34.960 ;
        RECT 26.240 34.640 26.560 34.960 ;
        RECT 26.640 34.640 26.960 34.960 ;
        RECT 27.040 34.640 27.360 34.960 ;
        RECT 27.440 34.640 27.760 34.960 ;
        RECT 27.840 34.640 28.160 34.960 ;
        RECT 28.240 34.640 28.560 34.960 ;
        RECT 28.640 34.640 28.960 34.960 ;
        RECT 29.040 34.640 29.360 34.960 ;
        RECT 29.440 34.640 29.760 34.960 ;
        RECT 29.840 34.640 30.160 34.960 ;
        RECT 30.240 34.640 30.560 34.960 ;
        RECT 30.640 34.640 30.960 34.960 ;
        RECT 31.040 34.640 31.360 34.960 ;
        RECT 31.440 34.640 31.760 34.960 ;
        RECT 31.840 34.640 32.160 34.960 ;
        RECT 32.240 34.640 32.560 34.960 ;
        RECT 32.640 34.640 32.960 34.960 ;
        RECT 33.040 34.640 33.360 34.960 ;
        RECT 33.440 34.640 33.760 34.960 ;
        RECT 33.840 34.640 34.160 34.960 ;
        RECT 34.240 34.640 34.560 34.960 ;
        RECT 34.640 34.640 34.960 34.960 ;
        RECT 35.040 34.640 35.360 34.960 ;
        RECT 35.440 34.640 35.760 34.960 ;
        RECT 35.840 34.640 36.160 34.960 ;
        RECT 36.240 34.640 36.560 34.960 ;
        RECT 36.640 34.640 36.960 34.960 ;
        RECT 37.040 34.640 37.360 34.960 ;
        RECT 37.440 34.640 37.760 34.960 ;
        RECT 37.840 34.640 38.160 34.960 ;
        RECT 38.240 34.640 38.560 34.960 ;
        RECT 38.640 34.640 38.960 34.960 ;
        RECT 39.040 34.640 39.360 34.960 ;
        RECT 39.440 34.640 39.760 34.960 ;
        RECT 39.840 34.640 40.160 34.960 ;
        RECT 40.240 34.640 40.560 34.960 ;
        RECT 40.640 34.640 40.960 34.960 ;
        RECT 41.040 34.640 41.360 34.960 ;
        RECT 41.440 34.640 41.760 34.960 ;
        RECT 41.840 34.640 42.160 34.960 ;
        RECT 42.240 34.640 42.560 34.960 ;
        RECT 42.640 34.640 42.960 34.960 ;
        RECT 43.040 34.640 43.360 34.960 ;
        RECT 43.440 34.640 43.760 34.960 ;
        RECT 43.840 34.640 44.160 34.960 ;
        RECT 44.240 34.640 44.560 34.960 ;
        RECT 44.640 34.640 44.960 34.960 ;
        RECT 70.560 34.640 70.880 34.960 ;
        RECT 70.960 34.640 71.280 34.960 ;
        RECT 71.360 34.640 71.680 34.960 ;
        RECT 71.760 34.640 72.080 34.960 ;
        RECT 120.560 34.640 120.880 34.960 ;
        RECT 120.960 34.640 121.280 34.960 ;
        RECT 121.360 34.640 121.680 34.960 ;
        RECT 121.760 34.640 122.080 34.960 ;
        RECT 160.720 34.640 161.040 34.960 ;
        RECT 161.120 34.640 161.440 34.960 ;
        RECT 161.520 34.640 161.840 34.960 ;
        RECT 161.920 34.640 162.240 34.960 ;
        RECT 162.320 34.640 162.640 34.960 ;
        RECT 162.720 34.640 163.040 34.960 ;
        RECT 163.120 34.640 163.440 34.960 ;
        RECT 163.520 34.640 163.840 34.960 ;
        RECT 163.920 34.640 164.240 34.960 ;
        RECT 164.320 34.640 164.640 34.960 ;
        RECT 164.720 34.640 165.040 34.960 ;
        RECT 165.120 34.640 165.440 34.960 ;
        RECT 165.520 34.640 165.840 34.960 ;
        RECT 165.920 34.640 166.240 34.960 ;
        RECT 166.320 34.640 166.640 34.960 ;
        RECT 166.720 34.640 167.040 34.960 ;
        RECT 167.120 34.640 167.440 34.960 ;
        RECT 167.520 34.640 167.840 34.960 ;
        RECT 167.920 34.640 168.240 34.960 ;
        RECT 168.320 34.640 168.640 34.960 ;
        RECT 168.720 34.640 169.040 34.960 ;
        RECT 169.120 34.640 169.440 34.960 ;
        RECT 169.520 34.640 169.840 34.960 ;
        RECT 169.920 34.640 170.240 34.960 ;
        RECT 170.320 34.640 170.640 34.960 ;
        RECT 170.720 34.640 171.040 34.960 ;
        RECT 171.120 34.640 171.440 34.960 ;
        RECT 171.520 34.640 171.840 34.960 ;
        RECT 171.920 34.640 172.240 34.960 ;
        RECT 172.320 34.640 172.640 34.960 ;
        RECT 172.720 34.640 173.040 34.960 ;
        RECT 173.120 34.640 173.440 34.960 ;
        RECT 173.520 34.640 173.840 34.960 ;
        RECT 173.920 34.640 174.240 34.960 ;
        RECT 174.320 34.640 174.640 34.960 ;
        RECT 174.720 34.640 175.040 34.960 ;
        RECT 175.120 34.640 175.440 34.960 ;
        RECT 175.520 34.640 175.840 34.960 ;
        RECT 175.920 34.640 176.240 34.960 ;
        RECT 176.320 34.640 176.640 34.960 ;
        RECT 176.720 34.640 177.040 34.960 ;
        RECT 177.120 34.640 177.440 34.960 ;
        RECT 177.520 34.640 177.840 34.960 ;
        RECT 177.920 34.640 178.240 34.960 ;
        RECT 178.320 34.640 178.640 34.960 ;
        RECT 178.720 34.640 179.040 34.960 ;
        RECT 179.120 34.640 179.440 34.960 ;
        RECT 179.520 34.640 179.840 34.960 ;
        RECT 179.920 34.640 180.240 34.960 ;
        RECT 180.320 34.640 180.640 34.960 ;
        RECT 25.040 34.240 25.360 34.560 ;
        RECT 25.440 34.240 25.760 34.560 ;
        RECT 25.840 34.240 26.160 34.560 ;
        RECT 26.240 34.240 26.560 34.560 ;
        RECT 26.640 34.240 26.960 34.560 ;
        RECT 27.040 34.240 27.360 34.560 ;
        RECT 27.440 34.240 27.760 34.560 ;
        RECT 27.840 34.240 28.160 34.560 ;
        RECT 28.240 34.240 28.560 34.560 ;
        RECT 28.640 34.240 28.960 34.560 ;
        RECT 29.040 34.240 29.360 34.560 ;
        RECT 29.440 34.240 29.760 34.560 ;
        RECT 29.840 34.240 30.160 34.560 ;
        RECT 30.240 34.240 30.560 34.560 ;
        RECT 30.640 34.240 30.960 34.560 ;
        RECT 31.040 34.240 31.360 34.560 ;
        RECT 31.440 34.240 31.760 34.560 ;
        RECT 31.840 34.240 32.160 34.560 ;
        RECT 32.240 34.240 32.560 34.560 ;
        RECT 32.640 34.240 32.960 34.560 ;
        RECT 33.040 34.240 33.360 34.560 ;
        RECT 33.440 34.240 33.760 34.560 ;
        RECT 33.840 34.240 34.160 34.560 ;
        RECT 34.240 34.240 34.560 34.560 ;
        RECT 34.640 34.240 34.960 34.560 ;
        RECT 35.040 34.240 35.360 34.560 ;
        RECT 35.440 34.240 35.760 34.560 ;
        RECT 35.840 34.240 36.160 34.560 ;
        RECT 36.240 34.240 36.560 34.560 ;
        RECT 36.640 34.240 36.960 34.560 ;
        RECT 37.040 34.240 37.360 34.560 ;
        RECT 37.440 34.240 37.760 34.560 ;
        RECT 37.840 34.240 38.160 34.560 ;
        RECT 38.240 34.240 38.560 34.560 ;
        RECT 38.640 34.240 38.960 34.560 ;
        RECT 39.040 34.240 39.360 34.560 ;
        RECT 39.440 34.240 39.760 34.560 ;
        RECT 39.840 34.240 40.160 34.560 ;
        RECT 40.240 34.240 40.560 34.560 ;
        RECT 40.640 34.240 40.960 34.560 ;
        RECT 41.040 34.240 41.360 34.560 ;
        RECT 41.440 34.240 41.760 34.560 ;
        RECT 41.840 34.240 42.160 34.560 ;
        RECT 42.240 34.240 42.560 34.560 ;
        RECT 42.640 34.240 42.960 34.560 ;
        RECT 43.040 34.240 43.360 34.560 ;
        RECT 43.440 34.240 43.760 34.560 ;
        RECT 43.840 34.240 44.160 34.560 ;
        RECT 44.240 34.240 44.560 34.560 ;
        RECT 44.640 34.240 44.960 34.560 ;
        RECT 70.560 34.240 70.880 34.560 ;
        RECT 70.960 34.240 71.280 34.560 ;
        RECT 71.360 34.240 71.680 34.560 ;
        RECT 71.760 34.240 72.080 34.560 ;
        RECT 120.560 34.240 120.880 34.560 ;
        RECT 120.960 34.240 121.280 34.560 ;
        RECT 121.360 34.240 121.680 34.560 ;
        RECT 121.760 34.240 122.080 34.560 ;
        RECT 160.720 34.240 161.040 34.560 ;
        RECT 161.120 34.240 161.440 34.560 ;
        RECT 161.520 34.240 161.840 34.560 ;
        RECT 161.920 34.240 162.240 34.560 ;
        RECT 162.320 34.240 162.640 34.560 ;
        RECT 162.720 34.240 163.040 34.560 ;
        RECT 163.120 34.240 163.440 34.560 ;
        RECT 163.520 34.240 163.840 34.560 ;
        RECT 163.920 34.240 164.240 34.560 ;
        RECT 164.320 34.240 164.640 34.560 ;
        RECT 164.720 34.240 165.040 34.560 ;
        RECT 165.120 34.240 165.440 34.560 ;
        RECT 165.520 34.240 165.840 34.560 ;
        RECT 165.920 34.240 166.240 34.560 ;
        RECT 166.320 34.240 166.640 34.560 ;
        RECT 166.720 34.240 167.040 34.560 ;
        RECT 167.120 34.240 167.440 34.560 ;
        RECT 167.520 34.240 167.840 34.560 ;
        RECT 167.920 34.240 168.240 34.560 ;
        RECT 168.320 34.240 168.640 34.560 ;
        RECT 168.720 34.240 169.040 34.560 ;
        RECT 169.120 34.240 169.440 34.560 ;
        RECT 169.520 34.240 169.840 34.560 ;
        RECT 169.920 34.240 170.240 34.560 ;
        RECT 170.320 34.240 170.640 34.560 ;
        RECT 170.720 34.240 171.040 34.560 ;
        RECT 171.120 34.240 171.440 34.560 ;
        RECT 171.520 34.240 171.840 34.560 ;
        RECT 171.920 34.240 172.240 34.560 ;
        RECT 172.320 34.240 172.640 34.560 ;
        RECT 172.720 34.240 173.040 34.560 ;
        RECT 173.120 34.240 173.440 34.560 ;
        RECT 173.520 34.240 173.840 34.560 ;
        RECT 173.920 34.240 174.240 34.560 ;
        RECT 174.320 34.240 174.640 34.560 ;
        RECT 174.720 34.240 175.040 34.560 ;
        RECT 175.120 34.240 175.440 34.560 ;
        RECT 175.520 34.240 175.840 34.560 ;
        RECT 175.920 34.240 176.240 34.560 ;
        RECT 176.320 34.240 176.640 34.560 ;
        RECT 176.720 34.240 177.040 34.560 ;
        RECT 177.120 34.240 177.440 34.560 ;
        RECT 177.520 34.240 177.840 34.560 ;
        RECT 177.920 34.240 178.240 34.560 ;
        RECT 178.320 34.240 178.640 34.560 ;
        RECT 178.720 34.240 179.040 34.560 ;
        RECT 179.120 34.240 179.440 34.560 ;
        RECT 179.520 34.240 179.840 34.560 ;
        RECT 179.920 34.240 180.240 34.560 ;
        RECT 180.320 34.240 180.640 34.560 ;
        RECT 25.040 33.840 25.360 34.160 ;
        RECT 25.440 33.840 25.760 34.160 ;
        RECT 25.840 33.840 26.160 34.160 ;
        RECT 26.240 33.840 26.560 34.160 ;
        RECT 26.640 33.840 26.960 34.160 ;
        RECT 27.040 33.840 27.360 34.160 ;
        RECT 27.440 33.840 27.760 34.160 ;
        RECT 27.840 33.840 28.160 34.160 ;
        RECT 28.240 33.840 28.560 34.160 ;
        RECT 28.640 33.840 28.960 34.160 ;
        RECT 29.040 33.840 29.360 34.160 ;
        RECT 29.440 33.840 29.760 34.160 ;
        RECT 29.840 33.840 30.160 34.160 ;
        RECT 30.240 33.840 30.560 34.160 ;
        RECT 30.640 33.840 30.960 34.160 ;
        RECT 31.040 33.840 31.360 34.160 ;
        RECT 31.440 33.840 31.760 34.160 ;
        RECT 31.840 33.840 32.160 34.160 ;
        RECT 32.240 33.840 32.560 34.160 ;
        RECT 32.640 33.840 32.960 34.160 ;
        RECT 33.040 33.840 33.360 34.160 ;
        RECT 33.440 33.840 33.760 34.160 ;
        RECT 33.840 33.840 34.160 34.160 ;
        RECT 34.240 33.840 34.560 34.160 ;
        RECT 34.640 33.840 34.960 34.160 ;
        RECT 35.040 33.840 35.360 34.160 ;
        RECT 35.440 33.840 35.760 34.160 ;
        RECT 35.840 33.840 36.160 34.160 ;
        RECT 36.240 33.840 36.560 34.160 ;
        RECT 36.640 33.840 36.960 34.160 ;
        RECT 37.040 33.840 37.360 34.160 ;
        RECT 37.440 33.840 37.760 34.160 ;
        RECT 37.840 33.840 38.160 34.160 ;
        RECT 38.240 33.840 38.560 34.160 ;
        RECT 38.640 33.840 38.960 34.160 ;
        RECT 39.040 33.840 39.360 34.160 ;
        RECT 39.440 33.840 39.760 34.160 ;
        RECT 39.840 33.840 40.160 34.160 ;
        RECT 40.240 33.840 40.560 34.160 ;
        RECT 40.640 33.840 40.960 34.160 ;
        RECT 41.040 33.840 41.360 34.160 ;
        RECT 41.440 33.840 41.760 34.160 ;
        RECT 41.840 33.840 42.160 34.160 ;
        RECT 42.240 33.840 42.560 34.160 ;
        RECT 42.640 33.840 42.960 34.160 ;
        RECT 43.040 33.840 43.360 34.160 ;
        RECT 43.440 33.840 43.760 34.160 ;
        RECT 43.840 33.840 44.160 34.160 ;
        RECT 44.240 33.840 44.560 34.160 ;
        RECT 44.640 33.840 44.960 34.160 ;
        RECT 70.560 33.840 70.880 34.160 ;
        RECT 70.960 33.840 71.280 34.160 ;
        RECT 71.360 33.840 71.680 34.160 ;
        RECT 71.760 33.840 72.080 34.160 ;
        RECT 120.560 33.840 120.880 34.160 ;
        RECT 120.960 33.840 121.280 34.160 ;
        RECT 121.360 33.840 121.680 34.160 ;
        RECT 121.760 33.840 122.080 34.160 ;
        RECT 160.720 33.840 161.040 34.160 ;
        RECT 161.120 33.840 161.440 34.160 ;
        RECT 161.520 33.840 161.840 34.160 ;
        RECT 161.920 33.840 162.240 34.160 ;
        RECT 162.320 33.840 162.640 34.160 ;
        RECT 162.720 33.840 163.040 34.160 ;
        RECT 163.120 33.840 163.440 34.160 ;
        RECT 163.520 33.840 163.840 34.160 ;
        RECT 163.920 33.840 164.240 34.160 ;
        RECT 164.320 33.840 164.640 34.160 ;
        RECT 164.720 33.840 165.040 34.160 ;
        RECT 165.120 33.840 165.440 34.160 ;
        RECT 165.520 33.840 165.840 34.160 ;
        RECT 165.920 33.840 166.240 34.160 ;
        RECT 166.320 33.840 166.640 34.160 ;
        RECT 166.720 33.840 167.040 34.160 ;
        RECT 167.120 33.840 167.440 34.160 ;
        RECT 167.520 33.840 167.840 34.160 ;
        RECT 167.920 33.840 168.240 34.160 ;
        RECT 168.320 33.840 168.640 34.160 ;
        RECT 168.720 33.840 169.040 34.160 ;
        RECT 169.120 33.840 169.440 34.160 ;
        RECT 169.520 33.840 169.840 34.160 ;
        RECT 169.920 33.840 170.240 34.160 ;
        RECT 170.320 33.840 170.640 34.160 ;
        RECT 170.720 33.840 171.040 34.160 ;
        RECT 171.120 33.840 171.440 34.160 ;
        RECT 171.520 33.840 171.840 34.160 ;
        RECT 171.920 33.840 172.240 34.160 ;
        RECT 172.320 33.840 172.640 34.160 ;
        RECT 172.720 33.840 173.040 34.160 ;
        RECT 173.120 33.840 173.440 34.160 ;
        RECT 173.520 33.840 173.840 34.160 ;
        RECT 173.920 33.840 174.240 34.160 ;
        RECT 174.320 33.840 174.640 34.160 ;
        RECT 174.720 33.840 175.040 34.160 ;
        RECT 175.120 33.840 175.440 34.160 ;
        RECT 175.520 33.840 175.840 34.160 ;
        RECT 175.920 33.840 176.240 34.160 ;
        RECT 176.320 33.840 176.640 34.160 ;
        RECT 176.720 33.840 177.040 34.160 ;
        RECT 177.120 33.840 177.440 34.160 ;
        RECT 177.520 33.840 177.840 34.160 ;
        RECT 177.920 33.840 178.240 34.160 ;
        RECT 178.320 33.840 178.640 34.160 ;
        RECT 178.720 33.840 179.040 34.160 ;
        RECT 179.120 33.840 179.440 34.160 ;
        RECT 179.520 33.840 179.840 34.160 ;
        RECT 179.920 33.840 180.240 34.160 ;
        RECT 180.320 33.840 180.640 34.160 ;
        RECT 25.040 33.440 25.360 33.760 ;
        RECT 25.440 33.440 25.760 33.760 ;
        RECT 25.840 33.440 26.160 33.760 ;
        RECT 26.240 33.440 26.560 33.760 ;
        RECT 26.640 33.440 26.960 33.760 ;
        RECT 27.040 33.440 27.360 33.760 ;
        RECT 27.440 33.440 27.760 33.760 ;
        RECT 27.840 33.440 28.160 33.760 ;
        RECT 28.240 33.440 28.560 33.760 ;
        RECT 28.640 33.440 28.960 33.760 ;
        RECT 29.040 33.440 29.360 33.760 ;
        RECT 29.440 33.440 29.760 33.760 ;
        RECT 29.840 33.440 30.160 33.760 ;
        RECT 30.240 33.440 30.560 33.760 ;
        RECT 30.640 33.440 30.960 33.760 ;
        RECT 31.040 33.440 31.360 33.760 ;
        RECT 31.440 33.440 31.760 33.760 ;
        RECT 31.840 33.440 32.160 33.760 ;
        RECT 32.240 33.440 32.560 33.760 ;
        RECT 32.640 33.440 32.960 33.760 ;
        RECT 33.040 33.440 33.360 33.760 ;
        RECT 33.440 33.440 33.760 33.760 ;
        RECT 33.840 33.440 34.160 33.760 ;
        RECT 34.240 33.440 34.560 33.760 ;
        RECT 34.640 33.440 34.960 33.760 ;
        RECT 35.040 33.440 35.360 33.760 ;
        RECT 35.440 33.440 35.760 33.760 ;
        RECT 35.840 33.440 36.160 33.760 ;
        RECT 36.240 33.440 36.560 33.760 ;
        RECT 36.640 33.440 36.960 33.760 ;
        RECT 37.040 33.440 37.360 33.760 ;
        RECT 37.440 33.440 37.760 33.760 ;
        RECT 37.840 33.440 38.160 33.760 ;
        RECT 38.240 33.440 38.560 33.760 ;
        RECT 38.640 33.440 38.960 33.760 ;
        RECT 39.040 33.440 39.360 33.760 ;
        RECT 39.440 33.440 39.760 33.760 ;
        RECT 39.840 33.440 40.160 33.760 ;
        RECT 40.240 33.440 40.560 33.760 ;
        RECT 40.640 33.440 40.960 33.760 ;
        RECT 41.040 33.440 41.360 33.760 ;
        RECT 41.440 33.440 41.760 33.760 ;
        RECT 41.840 33.440 42.160 33.760 ;
        RECT 42.240 33.440 42.560 33.760 ;
        RECT 42.640 33.440 42.960 33.760 ;
        RECT 43.040 33.440 43.360 33.760 ;
        RECT 43.440 33.440 43.760 33.760 ;
        RECT 43.840 33.440 44.160 33.760 ;
        RECT 44.240 33.440 44.560 33.760 ;
        RECT 44.640 33.440 44.960 33.760 ;
        RECT 70.560 33.440 70.880 33.760 ;
        RECT 70.960 33.440 71.280 33.760 ;
        RECT 71.360 33.440 71.680 33.760 ;
        RECT 71.760 33.440 72.080 33.760 ;
        RECT 120.560 33.440 120.880 33.760 ;
        RECT 120.960 33.440 121.280 33.760 ;
        RECT 121.360 33.440 121.680 33.760 ;
        RECT 121.760 33.440 122.080 33.760 ;
        RECT 160.720 33.440 161.040 33.760 ;
        RECT 161.120 33.440 161.440 33.760 ;
        RECT 161.520 33.440 161.840 33.760 ;
        RECT 161.920 33.440 162.240 33.760 ;
        RECT 162.320 33.440 162.640 33.760 ;
        RECT 162.720 33.440 163.040 33.760 ;
        RECT 163.120 33.440 163.440 33.760 ;
        RECT 163.520 33.440 163.840 33.760 ;
        RECT 163.920 33.440 164.240 33.760 ;
        RECT 164.320 33.440 164.640 33.760 ;
        RECT 164.720 33.440 165.040 33.760 ;
        RECT 165.120 33.440 165.440 33.760 ;
        RECT 165.520 33.440 165.840 33.760 ;
        RECT 165.920 33.440 166.240 33.760 ;
        RECT 166.320 33.440 166.640 33.760 ;
        RECT 166.720 33.440 167.040 33.760 ;
        RECT 167.120 33.440 167.440 33.760 ;
        RECT 167.520 33.440 167.840 33.760 ;
        RECT 167.920 33.440 168.240 33.760 ;
        RECT 168.320 33.440 168.640 33.760 ;
        RECT 168.720 33.440 169.040 33.760 ;
        RECT 169.120 33.440 169.440 33.760 ;
        RECT 169.520 33.440 169.840 33.760 ;
        RECT 169.920 33.440 170.240 33.760 ;
        RECT 170.320 33.440 170.640 33.760 ;
        RECT 170.720 33.440 171.040 33.760 ;
        RECT 171.120 33.440 171.440 33.760 ;
        RECT 171.520 33.440 171.840 33.760 ;
        RECT 171.920 33.440 172.240 33.760 ;
        RECT 172.320 33.440 172.640 33.760 ;
        RECT 172.720 33.440 173.040 33.760 ;
        RECT 173.120 33.440 173.440 33.760 ;
        RECT 173.520 33.440 173.840 33.760 ;
        RECT 173.920 33.440 174.240 33.760 ;
        RECT 174.320 33.440 174.640 33.760 ;
        RECT 174.720 33.440 175.040 33.760 ;
        RECT 175.120 33.440 175.440 33.760 ;
        RECT 175.520 33.440 175.840 33.760 ;
        RECT 175.920 33.440 176.240 33.760 ;
        RECT 176.320 33.440 176.640 33.760 ;
        RECT 176.720 33.440 177.040 33.760 ;
        RECT 177.120 33.440 177.440 33.760 ;
        RECT 177.520 33.440 177.840 33.760 ;
        RECT 177.920 33.440 178.240 33.760 ;
        RECT 178.320 33.440 178.640 33.760 ;
        RECT 178.720 33.440 179.040 33.760 ;
        RECT 179.120 33.440 179.440 33.760 ;
        RECT 179.520 33.440 179.840 33.760 ;
        RECT 179.920 33.440 180.240 33.760 ;
        RECT 180.320 33.440 180.640 33.760 ;
        RECT 25.040 33.040 25.360 33.360 ;
        RECT 25.440 33.040 25.760 33.360 ;
        RECT 25.840 33.040 26.160 33.360 ;
        RECT 26.240 33.040 26.560 33.360 ;
        RECT 26.640 33.040 26.960 33.360 ;
        RECT 27.040 33.040 27.360 33.360 ;
        RECT 27.440 33.040 27.760 33.360 ;
        RECT 27.840 33.040 28.160 33.360 ;
        RECT 28.240 33.040 28.560 33.360 ;
        RECT 28.640 33.040 28.960 33.360 ;
        RECT 29.040 33.040 29.360 33.360 ;
        RECT 29.440 33.040 29.760 33.360 ;
        RECT 29.840 33.040 30.160 33.360 ;
        RECT 30.240 33.040 30.560 33.360 ;
        RECT 30.640 33.040 30.960 33.360 ;
        RECT 31.040 33.040 31.360 33.360 ;
        RECT 31.440 33.040 31.760 33.360 ;
        RECT 31.840 33.040 32.160 33.360 ;
        RECT 32.240 33.040 32.560 33.360 ;
        RECT 32.640 33.040 32.960 33.360 ;
        RECT 33.040 33.040 33.360 33.360 ;
        RECT 33.440 33.040 33.760 33.360 ;
        RECT 33.840 33.040 34.160 33.360 ;
        RECT 34.240 33.040 34.560 33.360 ;
        RECT 34.640 33.040 34.960 33.360 ;
        RECT 35.040 33.040 35.360 33.360 ;
        RECT 35.440 33.040 35.760 33.360 ;
        RECT 35.840 33.040 36.160 33.360 ;
        RECT 36.240 33.040 36.560 33.360 ;
        RECT 36.640 33.040 36.960 33.360 ;
        RECT 37.040 33.040 37.360 33.360 ;
        RECT 37.440 33.040 37.760 33.360 ;
        RECT 37.840 33.040 38.160 33.360 ;
        RECT 38.240 33.040 38.560 33.360 ;
        RECT 38.640 33.040 38.960 33.360 ;
        RECT 39.040 33.040 39.360 33.360 ;
        RECT 39.440 33.040 39.760 33.360 ;
        RECT 39.840 33.040 40.160 33.360 ;
        RECT 40.240 33.040 40.560 33.360 ;
        RECT 40.640 33.040 40.960 33.360 ;
        RECT 41.040 33.040 41.360 33.360 ;
        RECT 41.440 33.040 41.760 33.360 ;
        RECT 41.840 33.040 42.160 33.360 ;
        RECT 42.240 33.040 42.560 33.360 ;
        RECT 42.640 33.040 42.960 33.360 ;
        RECT 43.040 33.040 43.360 33.360 ;
        RECT 43.440 33.040 43.760 33.360 ;
        RECT 43.840 33.040 44.160 33.360 ;
        RECT 44.240 33.040 44.560 33.360 ;
        RECT 44.640 33.040 44.960 33.360 ;
        RECT 70.560 33.040 70.880 33.360 ;
        RECT 70.960 33.040 71.280 33.360 ;
        RECT 71.360 33.040 71.680 33.360 ;
        RECT 71.760 33.040 72.080 33.360 ;
        RECT 120.560 33.040 120.880 33.360 ;
        RECT 120.960 33.040 121.280 33.360 ;
        RECT 121.360 33.040 121.680 33.360 ;
        RECT 121.760 33.040 122.080 33.360 ;
        RECT 160.720 33.040 161.040 33.360 ;
        RECT 161.120 33.040 161.440 33.360 ;
        RECT 161.520 33.040 161.840 33.360 ;
        RECT 161.920 33.040 162.240 33.360 ;
        RECT 162.320 33.040 162.640 33.360 ;
        RECT 162.720 33.040 163.040 33.360 ;
        RECT 163.120 33.040 163.440 33.360 ;
        RECT 163.520 33.040 163.840 33.360 ;
        RECT 163.920 33.040 164.240 33.360 ;
        RECT 164.320 33.040 164.640 33.360 ;
        RECT 164.720 33.040 165.040 33.360 ;
        RECT 165.120 33.040 165.440 33.360 ;
        RECT 165.520 33.040 165.840 33.360 ;
        RECT 165.920 33.040 166.240 33.360 ;
        RECT 166.320 33.040 166.640 33.360 ;
        RECT 166.720 33.040 167.040 33.360 ;
        RECT 167.120 33.040 167.440 33.360 ;
        RECT 167.520 33.040 167.840 33.360 ;
        RECT 167.920 33.040 168.240 33.360 ;
        RECT 168.320 33.040 168.640 33.360 ;
        RECT 168.720 33.040 169.040 33.360 ;
        RECT 169.120 33.040 169.440 33.360 ;
        RECT 169.520 33.040 169.840 33.360 ;
        RECT 169.920 33.040 170.240 33.360 ;
        RECT 170.320 33.040 170.640 33.360 ;
        RECT 170.720 33.040 171.040 33.360 ;
        RECT 171.120 33.040 171.440 33.360 ;
        RECT 171.520 33.040 171.840 33.360 ;
        RECT 171.920 33.040 172.240 33.360 ;
        RECT 172.320 33.040 172.640 33.360 ;
        RECT 172.720 33.040 173.040 33.360 ;
        RECT 173.120 33.040 173.440 33.360 ;
        RECT 173.520 33.040 173.840 33.360 ;
        RECT 173.920 33.040 174.240 33.360 ;
        RECT 174.320 33.040 174.640 33.360 ;
        RECT 174.720 33.040 175.040 33.360 ;
        RECT 175.120 33.040 175.440 33.360 ;
        RECT 175.520 33.040 175.840 33.360 ;
        RECT 175.920 33.040 176.240 33.360 ;
        RECT 176.320 33.040 176.640 33.360 ;
        RECT 176.720 33.040 177.040 33.360 ;
        RECT 177.120 33.040 177.440 33.360 ;
        RECT 177.520 33.040 177.840 33.360 ;
        RECT 177.920 33.040 178.240 33.360 ;
        RECT 178.320 33.040 178.640 33.360 ;
        RECT 178.720 33.040 179.040 33.360 ;
        RECT 179.120 33.040 179.440 33.360 ;
        RECT 179.520 33.040 179.840 33.360 ;
        RECT 179.920 33.040 180.240 33.360 ;
        RECT 180.320 33.040 180.640 33.360 ;
        RECT 25.040 32.640 25.360 32.960 ;
        RECT 25.440 32.640 25.760 32.960 ;
        RECT 25.840 32.640 26.160 32.960 ;
        RECT 26.240 32.640 26.560 32.960 ;
        RECT 26.640 32.640 26.960 32.960 ;
        RECT 27.040 32.640 27.360 32.960 ;
        RECT 27.440 32.640 27.760 32.960 ;
        RECT 27.840 32.640 28.160 32.960 ;
        RECT 28.240 32.640 28.560 32.960 ;
        RECT 28.640 32.640 28.960 32.960 ;
        RECT 29.040 32.640 29.360 32.960 ;
        RECT 29.440 32.640 29.760 32.960 ;
        RECT 29.840 32.640 30.160 32.960 ;
        RECT 30.240 32.640 30.560 32.960 ;
        RECT 30.640 32.640 30.960 32.960 ;
        RECT 31.040 32.640 31.360 32.960 ;
        RECT 31.440 32.640 31.760 32.960 ;
        RECT 31.840 32.640 32.160 32.960 ;
        RECT 32.240 32.640 32.560 32.960 ;
        RECT 32.640 32.640 32.960 32.960 ;
        RECT 33.040 32.640 33.360 32.960 ;
        RECT 33.440 32.640 33.760 32.960 ;
        RECT 33.840 32.640 34.160 32.960 ;
        RECT 34.240 32.640 34.560 32.960 ;
        RECT 34.640 32.640 34.960 32.960 ;
        RECT 35.040 32.640 35.360 32.960 ;
        RECT 35.440 32.640 35.760 32.960 ;
        RECT 35.840 32.640 36.160 32.960 ;
        RECT 36.240 32.640 36.560 32.960 ;
        RECT 36.640 32.640 36.960 32.960 ;
        RECT 37.040 32.640 37.360 32.960 ;
        RECT 37.440 32.640 37.760 32.960 ;
        RECT 37.840 32.640 38.160 32.960 ;
        RECT 38.240 32.640 38.560 32.960 ;
        RECT 38.640 32.640 38.960 32.960 ;
        RECT 39.040 32.640 39.360 32.960 ;
        RECT 39.440 32.640 39.760 32.960 ;
        RECT 39.840 32.640 40.160 32.960 ;
        RECT 40.240 32.640 40.560 32.960 ;
        RECT 40.640 32.640 40.960 32.960 ;
        RECT 41.040 32.640 41.360 32.960 ;
        RECT 41.440 32.640 41.760 32.960 ;
        RECT 41.840 32.640 42.160 32.960 ;
        RECT 42.240 32.640 42.560 32.960 ;
        RECT 42.640 32.640 42.960 32.960 ;
        RECT 43.040 32.640 43.360 32.960 ;
        RECT 43.440 32.640 43.760 32.960 ;
        RECT 43.840 32.640 44.160 32.960 ;
        RECT 44.240 32.640 44.560 32.960 ;
        RECT 44.640 32.640 44.960 32.960 ;
        RECT 70.560 32.640 70.880 32.960 ;
        RECT 70.960 32.640 71.280 32.960 ;
        RECT 71.360 32.640 71.680 32.960 ;
        RECT 71.760 32.640 72.080 32.960 ;
        RECT 120.560 32.640 120.880 32.960 ;
        RECT 120.960 32.640 121.280 32.960 ;
        RECT 121.360 32.640 121.680 32.960 ;
        RECT 121.760 32.640 122.080 32.960 ;
        RECT 160.720 32.640 161.040 32.960 ;
        RECT 161.120 32.640 161.440 32.960 ;
        RECT 161.520 32.640 161.840 32.960 ;
        RECT 161.920 32.640 162.240 32.960 ;
        RECT 162.320 32.640 162.640 32.960 ;
        RECT 162.720 32.640 163.040 32.960 ;
        RECT 163.120 32.640 163.440 32.960 ;
        RECT 163.520 32.640 163.840 32.960 ;
        RECT 163.920 32.640 164.240 32.960 ;
        RECT 164.320 32.640 164.640 32.960 ;
        RECT 164.720 32.640 165.040 32.960 ;
        RECT 165.120 32.640 165.440 32.960 ;
        RECT 165.520 32.640 165.840 32.960 ;
        RECT 165.920 32.640 166.240 32.960 ;
        RECT 166.320 32.640 166.640 32.960 ;
        RECT 166.720 32.640 167.040 32.960 ;
        RECT 167.120 32.640 167.440 32.960 ;
        RECT 167.520 32.640 167.840 32.960 ;
        RECT 167.920 32.640 168.240 32.960 ;
        RECT 168.320 32.640 168.640 32.960 ;
        RECT 168.720 32.640 169.040 32.960 ;
        RECT 169.120 32.640 169.440 32.960 ;
        RECT 169.520 32.640 169.840 32.960 ;
        RECT 169.920 32.640 170.240 32.960 ;
        RECT 170.320 32.640 170.640 32.960 ;
        RECT 170.720 32.640 171.040 32.960 ;
        RECT 171.120 32.640 171.440 32.960 ;
        RECT 171.520 32.640 171.840 32.960 ;
        RECT 171.920 32.640 172.240 32.960 ;
        RECT 172.320 32.640 172.640 32.960 ;
        RECT 172.720 32.640 173.040 32.960 ;
        RECT 173.120 32.640 173.440 32.960 ;
        RECT 173.520 32.640 173.840 32.960 ;
        RECT 173.920 32.640 174.240 32.960 ;
        RECT 174.320 32.640 174.640 32.960 ;
        RECT 174.720 32.640 175.040 32.960 ;
        RECT 175.120 32.640 175.440 32.960 ;
        RECT 175.520 32.640 175.840 32.960 ;
        RECT 175.920 32.640 176.240 32.960 ;
        RECT 176.320 32.640 176.640 32.960 ;
        RECT 176.720 32.640 177.040 32.960 ;
        RECT 177.120 32.640 177.440 32.960 ;
        RECT 177.520 32.640 177.840 32.960 ;
        RECT 177.920 32.640 178.240 32.960 ;
        RECT 178.320 32.640 178.640 32.960 ;
        RECT 178.720 32.640 179.040 32.960 ;
        RECT 179.120 32.640 179.440 32.960 ;
        RECT 179.520 32.640 179.840 32.960 ;
        RECT 179.920 32.640 180.240 32.960 ;
        RECT 180.320 32.640 180.640 32.960 ;
        RECT 25.040 32.240 25.360 32.560 ;
        RECT 25.440 32.240 25.760 32.560 ;
        RECT 25.840 32.240 26.160 32.560 ;
        RECT 26.240 32.240 26.560 32.560 ;
        RECT 26.640 32.240 26.960 32.560 ;
        RECT 27.040 32.240 27.360 32.560 ;
        RECT 27.440 32.240 27.760 32.560 ;
        RECT 27.840 32.240 28.160 32.560 ;
        RECT 28.240 32.240 28.560 32.560 ;
        RECT 28.640 32.240 28.960 32.560 ;
        RECT 29.040 32.240 29.360 32.560 ;
        RECT 29.440 32.240 29.760 32.560 ;
        RECT 29.840 32.240 30.160 32.560 ;
        RECT 30.240 32.240 30.560 32.560 ;
        RECT 30.640 32.240 30.960 32.560 ;
        RECT 31.040 32.240 31.360 32.560 ;
        RECT 31.440 32.240 31.760 32.560 ;
        RECT 31.840 32.240 32.160 32.560 ;
        RECT 32.240 32.240 32.560 32.560 ;
        RECT 32.640 32.240 32.960 32.560 ;
        RECT 33.040 32.240 33.360 32.560 ;
        RECT 33.440 32.240 33.760 32.560 ;
        RECT 33.840 32.240 34.160 32.560 ;
        RECT 34.240 32.240 34.560 32.560 ;
        RECT 34.640 32.240 34.960 32.560 ;
        RECT 35.040 32.240 35.360 32.560 ;
        RECT 35.440 32.240 35.760 32.560 ;
        RECT 35.840 32.240 36.160 32.560 ;
        RECT 36.240 32.240 36.560 32.560 ;
        RECT 36.640 32.240 36.960 32.560 ;
        RECT 37.040 32.240 37.360 32.560 ;
        RECT 37.440 32.240 37.760 32.560 ;
        RECT 37.840 32.240 38.160 32.560 ;
        RECT 38.240 32.240 38.560 32.560 ;
        RECT 38.640 32.240 38.960 32.560 ;
        RECT 39.040 32.240 39.360 32.560 ;
        RECT 39.440 32.240 39.760 32.560 ;
        RECT 39.840 32.240 40.160 32.560 ;
        RECT 40.240 32.240 40.560 32.560 ;
        RECT 40.640 32.240 40.960 32.560 ;
        RECT 41.040 32.240 41.360 32.560 ;
        RECT 41.440 32.240 41.760 32.560 ;
        RECT 41.840 32.240 42.160 32.560 ;
        RECT 42.240 32.240 42.560 32.560 ;
        RECT 42.640 32.240 42.960 32.560 ;
        RECT 43.040 32.240 43.360 32.560 ;
        RECT 43.440 32.240 43.760 32.560 ;
        RECT 43.840 32.240 44.160 32.560 ;
        RECT 44.240 32.240 44.560 32.560 ;
        RECT 44.640 32.240 44.960 32.560 ;
        RECT 70.560 32.240 70.880 32.560 ;
        RECT 70.960 32.240 71.280 32.560 ;
        RECT 71.360 32.240 71.680 32.560 ;
        RECT 71.760 32.240 72.080 32.560 ;
        RECT 120.560 32.240 120.880 32.560 ;
        RECT 120.960 32.240 121.280 32.560 ;
        RECT 121.360 32.240 121.680 32.560 ;
        RECT 121.760 32.240 122.080 32.560 ;
        RECT 160.720 32.240 161.040 32.560 ;
        RECT 161.120 32.240 161.440 32.560 ;
        RECT 161.520 32.240 161.840 32.560 ;
        RECT 161.920 32.240 162.240 32.560 ;
        RECT 162.320 32.240 162.640 32.560 ;
        RECT 162.720 32.240 163.040 32.560 ;
        RECT 163.120 32.240 163.440 32.560 ;
        RECT 163.520 32.240 163.840 32.560 ;
        RECT 163.920 32.240 164.240 32.560 ;
        RECT 164.320 32.240 164.640 32.560 ;
        RECT 164.720 32.240 165.040 32.560 ;
        RECT 165.120 32.240 165.440 32.560 ;
        RECT 165.520 32.240 165.840 32.560 ;
        RECT 165.920 32.240 166.240 32.560 ;
        RECT 166.320 32.240 166.640 32.560 ;
        RECT 166.720 32.240 167.040 32.560 ;
        RECT 167.120 32.240 167.440 32.560 ;
        RECT 167.520 32.240 167.840 32.560 ;
        RECT 167.920 32.240 168.240 32.560 ;
        RECT 168.320 32.240 168.640 32.560 ;
        RECT 168.720 32.240 169.040 32.560 ;
        RECT 169.120 32.240 169.440 32.560 ;
        RECT 169.520 32.240 169.840 32.560 ;
        RECT 169.920 32.240 170.240 32.560 ;
        RECT 170.320 32.240 170.640 32.560 ;
        RECT 170.720 32.240 171.040 32.560 ;
        RECT 171.120 32.240 171.440 32.560 ;
        RECT 171.520 32.240 171.840 32.560 ;
        RECT 171.920 32.240 172.240 32.560 ;
        RECT 172.320 32.240 172.640 32.560 ;
        RECT 172.720 32.240 173.040 32.560 ;
        RECT 173.120 32.240 173.440 32.560 ;
        RECT 173.520 32.240 173.840 32.560 ;
        RECT 173.920 32.240 174.240 32.560 ;
        RECT 174.320 32.240 174.640 32.560 ;
        RECT 174.720 32.240 175.040 32.560 ;
        RECT 175.120 32.240 175.440 32.560 ;
        RECT 175.520 32.240 175.840 32.560 ;
        RECT 175.920 32.240 176.240 32.560 ;
        RECT 176.320 32.240 176.640 32.560 ;
        RECT 176.720 32.240 177.040 32.560 ;
        RECT 177.120 32.240 177.440 32.560 ;
        RECT 177.520 32.240 177.840 32.560 ;
        RECT 177.920 32.240 178.240 32.560 ;
        RECT 178.320 32.240 178.640 32.560 ;
        RECT 178.720 32.240 179.040 32.560 ;
        RECT 179.120 32.240 179.440 32.560 ;
        RECT 179.520 32.240 179.840 32.560 ;
        RECT 179.920 32.240 180.240 32.560 ;
        RECT 180.320 32.240 180.640 32.560 ;
        RECT 25.040 31.840 25.360 32.160 ;
        RECT 25.440 31.840 25.760 32.160 ;
        RECT 25.840 31.840 26.160 32.160 ;
        RECT 26.240 31.840 26.560 32.160 ;
        RECT 26.640 31.840 26.960 32.160 ;
        RECT 27.040 31.840 27.360 32.160 ;
        RECT 27.440 31.840 27.760 32.160 ;
        RECT 27.840 31.840 28.160 32.160 ;
        RECT 28.240 31.840 28.560 32.160 ;
        RECT 28.640 31.840 28.960 32.160 ;
        RECT 29.040 31.840 29.360 32.160 ;
        RECT 29.440 31.840 29.760 32.160 ;
        RECT 29.840 31.840 30.160 32.160 ;
        RECT 30.240 31.840 30.560 32.160 ;
        RECT 30.640 31.840 30.960 32.160 ;
        RECT 31.040 31.840 31.360 32.160 ;
        RECT 31.440 31.840 31.760 32.160 ;
        RECT 31.840 31.840 32.160 32.160 ;
        RECT 32.240 31.840 32.560 32.160 ;
        RECT 32.640 31.840 32.960 32.160 ;
        RECT 33.040 31.840 33.360 32.160 ;
        RECT 33.440 31.840 33.760 32.160 ;
        RECT 33.840 31.840 34.160 32.160 ;
        RECT 34.240 31.840 34.560 32.160 ;
        RECT 34.640 31.840 34.960 32.160 ;
        RECT 35.040 31.840 35.360 32.160 ;
        RECT 35.440 31.840 35.760 32.160 ;
        RECT 35.840 31.840 36.160 32.160 ;
        RECT 36.240 31.840 36.560 32.160 ;
        RECT 36.640 31.840 36.960 32.160 ;
        RECT 37.040 31.840 37.360 32.160 ;
        RECT 37.440 31.840 37.760 32.160 ;
        RECT 37.840 31.840 38.160 32.160 ;
        RECT 38.240 31.840 38.560 32.160 ;
        RECT 38.640 31.840 38.960 32.160 ;
        RECT 39.040 31.840 39.360 32.160 ;
        RECT 39.440 31.840 39.760 32.160 ;
        RECT 39.840 31.840 40.160 32.160 ;
        RECT 40.240 31.840 40.560 32.160 ;
        RECT 40.640 31.840 40.960 32.160 ;
        RECT 41.040 31.840 41.360 32.160 ;
        RECT 41.440 31.840 41.760 32.160 ;
        RECT 41.840 31.840 42.160 32.160 ;
        RECT 42.240 31.840 42.560 32.160 ;
        RECT 42.640 31.840 42.960 32.160 ;
        RECT 43.040 31.840 43.360 32.160 ;
        RECT 43.440 31.840 43.760 32.160 ;
        RECT 43.840 31.840 44.160 32.160 ;
        RECT 44.240 31.840 44.560 32.160 ;
        RECT 44.640 31.840 44.960 32.160 ;
        RECT 70.560 31.840 70.880 32.160 ;
        RECT 70.960 31.840 71.280 32.160 ;
        RECT 71.360 31.840 71.680 32.160 ;
        RECT 71.760 31.840 72.080 32.160 ;
        RECT 120.560 31.840 120.880 32.160 ;
        RECT 120.960 31.840 121.280 32.160 ;
        RECT 121.360 31.840 121.680 32.160 ;
        RECT 121.760 31.840 122.080 32.160 ;
        RECT 160.720 31.840 161.040 32.160 ;
        RECT 161.120 31.840 161.440 32.160 ;
        RECT 161.520 31.840 161.840 32.160 ;
        RECT 161.920 31.840 162.240 32.160 ;
        RECT 162.320 31.840 162.640 32.160 ;
        RECT 162.720 31.840 163.040 32.160 ;
        RECT 163.120 31.840 163.440 32.160 ;
        RECT 163.520 31.840 163.840 32.160 ;
        RECT 163.920 31.840 164.240 32.160 ;
        RECT 164.320 31.840 164.640 32.160 ;
        RECT 164.720 31.840 165.040 32.160 ;
        RECT 165.120 31.840 165.440 32.160 ;
        RECT 165.520 31.840 165.840 32.160 ;
        RECT 165.920 31.840 166.240 32.160 ;
        RECT 166.320 31.840 166.640 32.160 ;
        RECT 166.720 31.840 167.040 32.160 ;
        RECT 167.120 31.840 167.440 32.160 ;
        RECT 167.520 31.840 167.840 32.160 ;
        RECT 167.920 31.840 168.240 32.160 ;
        RECT 168.320 31.840 168.640 32.160 ;
        RECT 168.720 31.840 169.040 32.160 ;
        RECT 169.120 31.840 169.440 32.160 ;
        RECT 169.520 31.840 169.840 32.160 ;
        RECT 169.920 31.840 170.240 32.160 ;
        RECT 170.320 31.840 170.640 32.160 ;
        RECT 170.720 31.840 171.040 32.160 ;
        RECT 171.120 31.840 171.440 32.160 ;
        RECT 171.520 31.840 171.840 32.160 ;
        RECT 171.920 31.840 172.240 32.160 ;
        RECT 172.320 31.840 172.640 32.160 ;
        RECT 172.720 31.840 173.040 32.160 ;
        RECT 173.120 31.840 173.440 32.160 ;
        RECT 173.520 31.840 173.840 32.160 ;
        RECT 173.920 31.840 174.240 32.160 ;
        RECT 174.320 31.840 174.640 32.160 ;
        RECT 174.720 31.840 175.040 32.160 ;
        RECT 175.120 31.840 175.440 32.160 ;
        RECT 175.520 31.840 175.840 32.160 ;
        RECT 175.920 31.840 176.240 32.160 ;
        RECT 176.320 31.840 176.640 32.160 ;
        RECT 176.720 31.840 177.040 32.160 ;
        RECT 177.120 31.840 177.440 32.160 ;
        RECT 177.520 31.840 177.840 32.160 ;
        RECT 177.920 31.840 178.240 32.160 ;
        RECT 178.320 31.840 178.640 32.160 ;
        RECT 178.720 31.840 179.040 32.160 ;
        RECT 179.120 31.840 179.440 32.160 ;
        RECT 179.520 31.840 179.840 32.160 ;
        RECT 179.920 31.840 180.240 32.160 ;
        RECT 180.320 31.840 180.640 32.160 ;
        RECT 25.040 31.440 25.360 31.760 ;
        RECT 25.440 31.440 25.760 31.760 ;
        RECT 25.840 31.440 26.160 31.760 ;
        RECT 26.240 31.440 26.560 31.760 ;
        RECT 26.640 31.440 26.960 31.760 ;
        RECT 27.040 31.440 27.360 31.760 ;
        RECT 27.440 31.440 27.760 31.760 ;
        RECT 27.840 31.440 28.160 31.760 ;
        RECT 28.240 31.440 28.560 31.760 ;
        RECT 28.640 31.440 28.960 31.760 ;
        RECT 29.040 31.440 29.360 31.760 ;
        RECT 29.440 31.440 29.760 31.760 ;
        RECT 29.840 31.440 30.160 31.760 ;
        RECT 30.240 31.440 30.560 31.760 ;
        RECT 30.640 31.440 30.960 31.760 ;
        RECT 31.040 31.440 31.360 31.760 ;
        RECT 31.440 31.440 31.760 31.760 ;
        RECT 31.840 31.440 32.160 31.760 ;
        RECT 32.240 31.440 32.560 31.760 ;
        RECT 32.640 31.440 32.960 31.760 ;
        RECT 33.040 31.440 33.360 31.760 ;
        RECT 33.440 31.440 33.760 31.760 ;
        RECT 33.840 31.440 34.160 31.760 ;
        RECT 34.240 31.440 34.560 31.760 ;
        RECT 34.640 31.440 34.960 31.760 ;
        RECT 35.040 31.440 35.360 31.760 ;
        RECT 35.440 31.440 35.760 31.760 ;
        RECT 35.840 31.440 36.160 31.760 ;
        RECT 36.240 31.440 36.560 31.760 ;
        RECT 36.640 31.440 36.960 31.760 ;
        RECT 37.040 31.440 37.360 31.760 ;
        RECT 37.440 31.440 37.760 31.760 ;
        RECT 37.840 31.440 38.160 31.760 ;
        RECT 38.240 31.440 38.560 31.760 ;
        RECT 38.640 31.440 38.960 31.760 ;
        RECT 39.040 31.440 39.360 31.760 ;
        RECT 39.440 31.440 39.760 31.760 ;
        RECT 39.840 31.440 40.160 31.760 ;
        RECT 40.240 31.440 40.560 31.760 ;
        RECT 40.640 31.440 40.960 31.760 ;
        RECT 41.040 31.440 41.360 31.760 ;
        RECT 41.440 31.440 41.760 31.760 ;
        RECT 41.840 31.440 42.160 31.760 ;
        RECT 42.240 31.440 42.560 31.760 ;
        RECT 42.640 31.440 42.960 31.760 ;
        RECT 43.040 31.440 43.360 31.760 ;
        RECT 43.440 31.440 43.760 31.760 ;
        RECT 43.840 31.440 44.160 31.760 ;
        RECT 44.240 31.440 44.560 31.760 ;
        RECT 44.640 31.440 44.960 31.760 ;
        RECT 70.560 31.440 70.880 31.760 ;
        RECT 70.960 31.440 71.280 31.760 ;
        RECT 71.360 31.440 71.680 31.760 ;
        RECT 71.760 31.440 72.080 31.760 ;
        RECT 120.560 31.440 120.880 31.760 ;
        RECT 120.960 31.440 121.280 31.760 ;
        RECT 121.360 31.440 121.680 31.760 ;
        RECT 121.760 31.440 122.080 31.760 ;
        RECT 160.720 31.440 161.040 31.760 ;
        RECT 161.120 31.440 161.440 31.760 ;
        RECT 161.520 31.440 161.840 31.760 ;
        RECT 161.920 31.440 162.240 31.760 ;
        RECT 162.320 31.440 162.640 31.760 ;
        RECT 162.720 31.440 163.040 31.760 ;
        RECT 163.120 31.440 163.440 31.760 ;
        RECT 163.520 31.440 163.840 31.760 ;
        RECT 163.920 31.440 164.240 31.760 ;
        RECT 164.320 31.440 164.640 31.760 ;
        RECT 164.720 31.440 165.040 31.760 ;
        RECT 165.120 31.440 165.440 31.760 ;
        RECT 165.520 31.440 165.840 31.760 ;
        RECT 165.920 31.440 166.240 31.760 ;
        RECT 166.320 31.440 166.640 31.760 ;
        RECT 166.720 31.440 167.040 31.760 ;
        RECT 167.120 31.440 167.440 31.760 ;
        RECT 167.520 31.440 167.840 31.760 ;
        RECT 167.920 31.440 168.240 31.760 ;
        RECT 168.320 31.440 168.640 31.760 ;
        RECT 168.720 31.440 169.040 31.760 ;
        RECT 169.120 31.440 169.440 31.760 ;
        RECT 169.520 31.440 169.840 31.760 ;
        RECT 169.920 31.440 170.240 31.760 ;
        RECT 170.320 31.440 170.640 31.760 ;
        RECT 170.720 31.440 171.040 31.760 ;
        RECT 171.120 31.440 171.440 31.760 ;
        RECT 171.520 31.440 171.840 31.760 ;
        RECT 171.920 31.440 172.240 31.760 ;
        RECT 172.320 31.440 172.640 31.760 ;
        RECT 172.720 31.440 173.040 31.760 ;
        RECT 173.120 31.440 173.440 31.760 ;
        RECT 173.520 31.440 173.840 31.760 ;
        RECT 173.920 31.440 174.240 31.760 ;
        RECT 174.320 31.440 174.640 31.760 ;
        RECT 174.720 31.440 175.040 31.760 ;
        RECT 175.120 31.440 175.440 31.760 ;
        RECT 175.520 31.440 175.840 31.760 ;
        RECT 175.920 31.440 176.240 31.760 ;
        RECT 176.320 31.440 176.640 31.760 ;
        RECT 176.720 31.440 177.040 31.760 ;
        RECT 177.120 31.440 177.440 31.760 ;
        RECT 177.520 31.440 177.840 31.760 ;
        RECT 177.920 31.440 178.240 31.760 ;
        RECT 178.320 31.440 178.640 31.760 ;
        RECT 178.720 31.440 179.040 31.760 ;
        RECT 179.120 31.440 179.440 31.760 ;
        RECT 179.520 31.440 179.840 31.760 ;
        RECT 179.920 31.440 180.240 31.760 ;
        RECT 180.320 31.440 180.640 31.760 ;
        RECT 25.040 31.040 25.360 31.360 ;
        RECT 25.440 31.040 25.760 31.360 ;
        RECT 25.840 31.040 26.160 31.360 ;
        RECT 26.240 31.040 26.560 31.360 ;
        RECT 26.640 31.040 26.960 31.360 ;
        RECT 27.040 31.040 27.360 31.360 ;
        RECT 27.440 31.040 27.760 31.360 ;
        RECT 27.840 31.040 28.160 31.360 ;
        RECT 28.240 31.040 28.560 31.360 ;
        RECT 28.640 31.040 28.960 31.360 ;
        RECT 29.040 31.040 29.360 31.360 ;
        RECT 29.440 31.040 29.760 31.360 ;
        RECT 29.840 31.040 30.160 31.360 ;
        RECT 30.240 31.040 30.560 31.360 ;
        RECT 30.640 31.040 30.960 31.360 ;
        RECT 31.040 31.040 31.360 31.360 ;
        RECT 31.440 31.040 31.760 31.360 ;
        RECT 31.840 31.040 32.160 31.360 ;
        RECT 32.240 31.040 32.560 31.360 ;
        RECT 32.640 31.040 32.960 31.360 ;
        RECT 33.040 31.040 33.360 31.360 ;
        RECT 33.440 31.040 33.760 31.360 ;
        RECT 33.840 31.040 34.160 31.360 ;
        RECT 34.240 31.040 34.560 31.360 ;
        RECT 34.640 31.040 34.960 31.360 ;
        RECT 35.040 31.040 35.360 31.360 ;
        RECT 35.440 31.040 35.760 31.360 ;
        RECT 35.840 31.040 36.160 31.360 ;
        RECT 36.240 31.040 36.560 31.360 ;
        RECT 36.640 31.040 36.960 31.360 ;
        RECT 37.040 31.040 37.360 31.360 ;
        RECT 37.440 31.040 37.760 31.360 ;
        RECT 37.840 31.040 38.160 31.360 ;
        RECT 38.240 31.040 38.560 31.360 ;
        RECT 38.640 31.040 38.960 31.360 ;
        RECT 39.040 31.040 39.360 31.360 ;
        RECT 39.440 31.040 39.760 31.360 ;
        RECT 39.840 31.040 40.160 31.360 ;
        RECT 40.240 31.040 40.560 31.360 ;
        RECT 40.640 31.040 40.960 31.360 ;
        RECT 41.040 31.040 41.360 31.360 ;
        RECT 41.440 31.040 41.760 31.360 ;
        RECT 41.840 31.040 42.160 31.360 ;
        RECT 42.240 31.040 42.560 31.360 ;
        RECT 42.640 31.040 42.960 31.360 ;
        RECT 43.040 31.040 43.360 31.360 ;
        RECT 43.440 31.040 43.760 31.360 ;
        RECT 43.840 31.040 44.160 31.360 ;
        RECT 44.240 31.040 44.560 31.360 ;
        RECT 44.640 31.040 44.960 31.360 ;
        RECT 70.560 31.040 70.880 31.360 ;
        RECT 70.960 31.040 71.280 31.360 ;
        RECT 71.360 31.040 71.680 31.360 ;
        RECT 71.760 31.040 72.080 31.360 ;
        RECT 120.560 31.040 120.880 31.360 ;
        RECT 120.960 31.040 121.280 31.360 ;
        RECT 121.360 31.040 121.680 31.360 ;
        RECT 121.760 31.040 122.080 31.360 ;
        RECT 160.720 31.040 161.040 31.360 ;
        RECT 161.120 31.040 161.440 31.360 ;
        RECT 161.520 31.040 161.840 31.360 ;
        RECT 161.920 31.040 162.240 31.360 ;
        RECT 162.320 31.040 162.640 31.360 ;
        RECT 162.720 31.040 163.040 31.360 ;
        RECT 163.120 31.040 163.440 31.360 ;
        RECT 163.520 31.040 163.840 31.360 ;
        RECT 163.920 31.040 164.240 31.360 ;
        RECT 164.320 31.040 164.640 31.360 ;
        RECT 164.720 31.040 165.040 31.360 ;
        RECT 165.120 31.040 165.440 31.360 ;
        RECT 165.520 31.040 165.840 31.360 ;
        RECT 165.920 31.040 166.240 31.360 ;
        RECT 166.320 31.040 166.640 31.360 ;
        RECT 166.720 31.040 167.040 31.360 ;
        RECT 167.120 31.040 167.440 31.360 ;
        RECT 167.520 31.040 167.840 31.360 ;
        RECT 167.920 31.040 168.240 31.360 ;
        RECT 168.320 31.040 168.640 31.360 ;
        RECT 168.720 31.040 169.040 31.360 ;
        RECT 169.120 31.040 169.440 31.360 ;
        RECT 169.520 31.040 169.840 31.360 ;
        RECT 169.920 31.040 170.240 31.360 ;
        RECT 170.320 31.040 170.640 31.360 ;
        RECT 170.720 31.040 171.040 31.360 ;
        RECT 171.120 31.040 171.440 31.360 ;
        RECT 171.520 31.040 171.840 31.360 ;
        RECT 171.920 31.040 172.240 31.360 ;
        RECT 172.320 31.040 172.640 31.360 ;
        RECT 172.720 31.040 173.040 31.360 ;
        RECT 173.120 31.040 173.440 31.360 ;
        RECT 173.520 31.040 173.840 31.360 ;
        RECT 173.920 31.040 174.240 31.360 ;
        RECT 174.320 31.040 174.640 31.360 ;
        RECT 174.720 31.040 175.040 31.360 ;
        RECT 175.120 31.040 175.440 31.360 ;
        RECT 175.520 31.040 175.840 31.360 ;
        RECT 175.920 31.040 176.240 31.360 ;
        RECT 176.320 31.040 176.640 31.360 ;
        RECT 176.720 31.040 177.040 31.360 ;
        RECT 177.120 31.040 177.440 31.360 ;
        RECT 177.520 31.040 177.840 31.360 ;
        RECT 177.920 31.040 178.240 31.360 ;
        RECT 178.320 31.040 178.640 31.360 ;
        RECT 178.720 31.040 179.040 31.360 ;
        RECT 179.120 31.040 179.440 31.360 ;
        RECT 179.520 31.040 179.840 31.360 ;
        RECT 179.920 31.040 180.240 31.360 ;
        RECT 180.320 31.040 180.640 31.360 ;
        RECT 25.040 30.640 25.360 30.960 ;
        RECT 25.440 30.640 25.760 30.960 ;
        RECT 25.840 30.640 26.160 30.960 ;
        RECT 26.240 30.640 26.560 30.960 ;
        RECT 26.640 30.640 26.960 30.960 ;
        RECT 27.040 30.640 27.360 30.960 ;
        RECT 27.440 30.640 27.760 30.960 ;
        RECT 27.840 30.640 28.160 30.960 ;
        RECT 28.240 30.640 28.560 30.960 ;
        RECT 28.640 30.640 28.960 30.960 ;
        RECT 29.040 30.640 29.360 30.960 ;
        RECT 29.440 30.640 29.760 30.960 ;
        RECT 29.840 30.640 30.160 30.960 ;
        RECT 30.240 30.640 30.560 30.960 ;
        RECT 30.640 30.640 30.960 30.960 ;
        RECT 31.040 30.640 31.360 30.960 ;
        RECT 31.440 30.640 31.760 30.960 ;
        RECT 31.840 30.640 32.160 30.960 ;
        RECT 32.240 30.640 32.560 30.960 ;
        RECT 32.640 30.640 32.960 30.960 ;
        RECT 33.040 30.640 33.360 30.960 ;
        RECT 33.440 30.640 33.760 30.960 ;
        RECT 33.840 30.640 34.160 30.960 ;
        RECT 34.240 30.640 34.560 30.960 ;
        RECT 34.640 30.640 34.960 30.960 ;
        RECT 35.040 30.640 35.360 30.960 ;
        RECT 35.440 30.640 35.760 30.960 ;
        RECT 35.840 30.640 36.160 30.960 ;
        RECT 36.240 30.640 36.560 30.960 ;
        RECT 36.640 30.640 36.960 30.960 ;
        RECT 37.040 30.640 37.360 30.960 ;
        RECT 37.440 30.640 37.760 30.960 ;
        RECT 37.840 30.640 38.160 30.960 ;
        RECT 38.240 30.640 38.560 30.960 ;
        RECT 38.640 30.640 38.960 30.960 ;
        RECT 39.040 30.640 39.360 30.960 ;
        RECT 39.440 30.640 39.760 30.960 ;
        RECT 39.840 30.640 40.160 30.960 ;
        RECT 40.240 30.640 40.560 30.960 ;
        RECT 40.640 30.640 40.960 30.960 ;
        RECT 41.040 30.640 41.360 30.960 ;
        RECT 41.440 30.640 41.760 30.960 ;
        RECT 41.840 30.640 42.160 30.960 ;
        RECT 42.240 30.640 42.560 30.960 ;
        RECT 42.640 30.640 42.960 30.960 ;
        RECT 43.040 30.640 43.360 30.960 ;
        RECT 43.440 30.640 43.760 30.960 ;
        RECT 43.840 30.640 44.160 30.960 ;
        RECT 44.240 30.640 44.560 30.960 ;
        RECT 44.640 30.640 44.960 30.960 ;
        RECT 70.560 30.640 70.880 30.960 ;
        RECT 70.960 30.640 71.280 30.960 ;
        RECT 71.360 30.640 71.680 30.960 ;
        RECT 71.760 30.640 72.080 30.960 ;
        RECT 120.560 30.640 120.880 30.960 ;
        RECT 120.960 30.640 121.280 30.960 ;
        RECT 121.360 30.640 121.680 30.960 ;
        RECT 121.760 30.640 122.080 30.960 ;
        RECT 160.720 30.640 161.040 30.960 ;
        RECT 161.120 30.640 161.440 30.960 ;
        RECT 161.520 30.640 161.840 30.960 ;
        RECT 161.920 30.640 162.240 30.960 ;
        RECT 162.320 30.640 162.640 30.960 ;
        RECT 162.720 30.640 163.040 30.960 ;
        RECT 163.120 30.640 163.440 30.960 ;
        RECT 163.520 30.640 163.840 30.960 ;
        RECT 163.920 30.640 164.240 30.960 ;
        RECT 164.320 30.640 164.640 30.960 ;
        RECT 164.720 30.640 165.040 30.960 ;
        RECT 165.120 30.640 165.440 30.960 ;
        RECT 165.520 30.640 165.840 30.960 ;
        RECT 165.920 30.640 166.240 30.960 ;
        RECT 166.320 30.640 166.640 30.960 ;
        RECT 166.720 30.640 167.040 30.960 ;
        RECT 167.120 30.640 167.440 30.960 ;
        RECT 167.520 30.640 167.840 30.960 ;
        RECT 167.920 30.640 168.240 30.960 ;
        RECT 168.320 30.640 168.640 30.960 ;
        RECT 168.720 30.640 169.040 30.960 ;
        RECT 169.120 30.640 169.440 30.960 ;
        RECT 169.520 30.640 169.840 30.960 ;
        RECT 169.920 30.640 170.240 30.960 ;
        RECT 170.320 30.640 170.640 30.960 ;
        RECT 170.720 30.640 171.040 30.960 ;
        RECT 171.120 30.640 171.440 30.960 ;
        RECT 171.520 30.640 171.840 30.960 ;
        RECT 171.920 30.640 172.240 30.960 ;
        RECT 172.320 30.640 172.640 30.960 ;
        RECT 172.720 30.640 173.040 30.960 ;
        RECT 173.120 30.640 173.440 30.960 ;
        RECT 173.520 30.640 173.840 30.960 ;
        RECT 173.920 30.640 174.240 30.960 ;
        RECT 174.320 30.640 174.640 30.960 ;
        RECT 174.720 30.640 175.040 30.960 ;
        RECT 175.120 30.640 175.440 30.960 ;
        RECT 175.520 30.640 175.840 30.960 ;
        RECT 175.920 30.640 176.240 30.960 ;
        RECT 176.320 30.640 176.640 30.960 ;
        RECT 176.720 30.640 177.040 30.960 ;
        RECT 177.120 30.640 177.440 30.960 ;
        RECT 177.520 30.640 177.840 30.960 ;
        RECT 177.920 30.640 178.240 30.960 ;
        RECT 178.320 30.640 178.640 30.960 ;
        RECT 178.720 30.640 179.040 30.960 ;
        RECT 179.120 30.640 179.440 30.960 ;
        RECT 179.520 30.640 179.840 30.960 ;
        RECT 179.920 30.640 180.240 30.960 ;
        RECT 180.320 30.640 180.640 30.960 ;
        RECT 25.040 30.240 25.360 30.560 ;
        RECT 25.440 30.240 25.760 30.560 ;
        RECT 25.840 30.240 26.160 30.560 ;
        RECT 26.240 30.240 26.560 30.560 ;
        RECT 26.640 30.240 26.960 30.560 ;
        RECT 27.040 30.240 27.360 30.560 ;
        RECT 27.440 30.240 27.760 30.560 ;
        RECT 27.840 30.240 28.160 30.560 ;
        RECT 28.240 30.240 28.560 30.560 ;
        RECT 28.640 30.240 28.960 30.560 ;
        RECT 29.040 30.240 29.360 30.560 ;
        RECT 29.440 30.240 29.760 30.560 ;
        RECT 29.840 30.240 30.160 30.560 ;
        RECT 30.240 30.240 30.560 30.560 ;
        RECT 30.640 30.240 30.960 30.560 ;
        RECT 31.040 30.240 31.360 30.560 ;
        RECT 31.440 30.240 31.760 30.560 ;
        RECT 31.840 30.240 32.160 30.560 ;
        RECT 32.240 30.240 32.560 30.560 ;
        RECT 32.640 30.240 32.960 30.560 ;
        RECT 33.040 30.240 33.360 30.560 ;
        RECT 33.440 30.240 33.760 30.560 ;
        RECT 33.840 30.240 34.160 30.560 ;
        RECT 34.240 30.240 34.560 30.560 ;
        RECT 34.640 30.240 34.960 30.560 ;
        RECT 35.040 30.240 35.360 30.560 ;
        RECT 35.440 30.240 35.760 30.560 ;
        RECT 35.840 30.240 36.160 30.560 ;
        RECT 36.240 30.240 36.560 30.560 ;
        RECT 36.640 30.240 36.960 30.560 ;
        RECT 37.040 30.240 37.360 30.560 ;
        RECT 37.440 30.240 37.760 30.560 ;
        RECT 37.840 30.240 38.160 30.560 ;
        RECT 38.240 30.240 38.560 30.560 ;
        RECT 38.640 30.240 38.960 30.560 ;
        RECT 39.040 30.240 39.360 30.560 ;
        RECT 39.440 30.240 39.760 30.560 ;
        RECT 39.840 30.240 40.160 30.560 ;
        RECT 40.240 30.240 40.560 30.560 ;
        RECT 40.640 30.240 40.960 30.560 ;
        RECT 41.040 30.240 41.360 30.560 ;
        RECT 41.440 30.240 41.760 30.560 ;
        RECT 41.840 30.240 42.160 30.560 ;
        RECT 42.240 30.240 42.560 30.560 ;
        RECT 42.640 30.240 42.960 30.560 ;
        RECT 43.040 30.240 43.360 30.560 ;
        RECT 43.440 30.240 43.760 30.560 ;
        RECT 43.840 30.240 44.160 30.560 ;
        RECT 44.240 30.240 44.560 30.560 ;
        RECT 44.640 30.240 44.960 30.560 ;
        RECT 70.560 30.240 70.880 30.560 ;
        RECT 70.960 30.240 71.280 30.560 ;
        RECT 71.360 30.240 71.680 30.560 ;
        RECT 71.760 30.240 72.080 30.560 ;
        RECT 120.560 30.240 120.880 30.560 ;
        RECT 120.960 30.240 121.280 30.560 ;
        RECT 121.360 30.240 121.680 30.560 ;
        RECT 121.760 30.240 122.080 30.560 ;
        RECT 160.720 30.240 161.040 30.560 ;
        RECT 161.120 30.240 161.440 30.560 ;
        RECT 161.520 30.240 161.840 30.560 ;
        RECT 161.920 30.240 162.240 30.560 ;
        RECT 162.320 30.240 162.640 30.560 ;
        RECT 162.720 30.240 163.040 30.560 ;
        RECT 163.120 30.240 163.440 30.560 ;
        RECT 163.520 30.240 163.840 30.560 ;
        RECT 163.920 30.240 164.240 30.560 ;
        RECT 164.320 30.240 164.640 30.560 ;
        RECT 164.720 30.240 165.040 30.560 ;
        RECT 165.120 30.240 165.440 30.560 ;
        RECT 165.520 30.240 165.840 30.560 ;
        RECT 165.920 30.240 166.240 30.560 ;
        RECT 166.320 30.240 166.640 30.560 ;
        RECT 166.720 30.240 167.040 30.560 ;
        RECT 167.120 30.240 167.440 30.560 ;
        RECT 167.520 30.240 167.840 30.560 ;
        RECT 167.920 30.240 168.240 30.560 ;
        RECT 168.320 30.240 168.640 30.560 ;
        RECT 168.720 30.240 169.040 30.560 ;
        RECT 169.120 30.240 169.440 30.560 ;
        RECT 169.520 30.240 169.840 30.560 ;
        RECT 169.920 30.240 170.240 30.560 ;
        RECT 170.320 30.240 170.640 30.560 ;
        RECT 170.720 30.240 171.040 30.560 ;
        RECT 171.120 30.240 171.440 30.560 ;
        RECT 171.520 30.240 171.840 30.560 ;
        RECT 171.920 30.240 172.240 30.560 ;
        RECT 172.320 30.240 172.640 30.560 ;
        RECT 172.720 30.240 173.040 30.560 ;
        RECT 173.120 30.240 173.440 30.560 ;
        RECT 173.520 30.240 173.840 30.560 ;
        RECT 173.920 30.240 174.240 30.560 ;
        RECT 174.320 30.240 174.640 30.560 ;
        RECT 174.720 30.240 175.040 30.560 ;
        RECT 175.120 30.240 175.440 30.560 ;
        RECT 175.520 30.240 175.840 30.560 ;
        RECT 175.920 30.240 176.240 30.560 ;
        RECT 176.320 30.240 176.640 30.560 ;
        RECT 176.720 30.240 177.040 30.560 ;
        RECT 177.120 30.240 177.440 30.560 ;
        RECT 177.520 30.240 177.840 30.560 ;
        RECT 177.920 30.240 178.240 30.560 ;
        RECT 178.320 30.240 178.640 30.560 ;
        RECT 178.720 30.240 179.040 30.560 ;
        RECT 179.120 30.240 179.440 30.560 ;
        RECT 179.520 30.240 179.840 30.560 ;
        RECT 179.920 30.240 180.240 30.560 ;
        RECT 180.320 30.240 180.640 30.560 ;
        RECT 25.040 29.840 25.360 30.160 ;
        RECT 25.440 29.840 25.760 30.160 ;
        RECT 25.840 29.840 26.160 30.160 ;
        RECT 26.240 29.840 26.560 30.160 ;
        RECT 26.640 29.840 26.960 30.160 ;
        RECT 27.040 29.840 27.360 30.160 ;
        RECT 27.440 29.840 27.760 30.160 ;
        RECT 27.840 29.840 28.160 30.160 ;
        RECT 28.240 29.840 28.560 30.160 ;
        RECT 28.640 29.840 28.960 30.160 ;
        RECT 29.040 29.840 29.360 30.160 ;
        RECT 29.440 29.840 29.760 30.160 ;
        RECT 29.840 29.840 30.160 30.160 ;
        RECT 30.240 29.840 30.560 30.160 ;
        RECT 30.640 29.840 30.960 30.160 ;
        RECT 31.040 29.840 31.360 30.160 ;
        RECT 31.440 29.840 31.760 30.160 ;
        RECT 31.840 29.840 32.160 30.160 ;
        RECT 32.240 29.840 32.560 30.160 ;
        RECT 32.640 29.840 32.960 30.160 ;
        RECT 33.040 29.840 33.360 30.160 ;
        RECT 33.440 29.840 33.760 30.160 ;
        RECT 33.840 29.840 34.160 30.160 ;
        RECT 34.240 29.840 34.560 30.160 ;
        RECT 34.640 29.840 34.960 30.160 ;
        RECT 35.040 29.840 35.360 30.160 ;
        RECT 35.440 29.840 35.760 30.160 ;
        RECT 35.840 29.840 36.160 30.160 ;
        RECT 36.240 29.840 36.560 30.160 ;
        RECT 36.640 29.840 36.960 30.160 ;
        RECT 37.040 29.840 37.360 30.160 ;
        RECT 37.440 29.840 37.760 30.160 ;
        RECT 37.840 29.840 38.160 30.160 ;
        RECT 38.240 29.840 38.560 30.160 ;
        RECT 38.640 29.840 38.960 30.160 ;
        RECT 39.040 29.840 39.360 30.160 ;
        RECT 39.440 29.840 39.760 30.160 ;
        RECT 39.840 29.840 40.160 30.160 ;
        RECT 40.240 29.840 40.560 30.160 ;
        RECT 40.640 29.840 40.960 30.160 ;
        RECT 41.040 29.840 41.360 30.160 ;
        RECT 41.440 29.840 41.760 30.160 ;
        RECT 41.840 29.840 42.160 30.160 ;
        RECT 42.240 29.840 42.560 30.160 ;
        RECT 42.640 29.840 42.960 30.160 ;
        RECT 43.040 29.840 43.360 30.160 ;
        RECT 43.440 29.840 43.760 30.160 ;
        RECT 43.840 29.840 44.160 30.160 ;
        RECT 44.240 29.840 44.560 30.160 ;
        RECT 44.640 29.840 44.960 30.160 ;
        RECT 70.560 29.840 70.880 30.160 ;
        RECT 70.960 29.840 71.280 30.160 ;
        RECT 71.360 29.840 71.680 30.160 ;
        RECT 71.760 29.840 72.080 30.160 ;
        RECT 120.560 29.840 120.880 30.160 ;
        RECT 120.960 29.840 121.280 30.160 ;
        RECT 121.360 29.840 121.680 30.160 ;
        RECT 121.760 29.840 122.080 30.160 ;
        RECT 160.720 29.840 161.040 30.160 ;
        RECT 161.120 29.840 161.440 30.160 ;
        RECT 161.520 29.840 161.840 30.160 ;
        RECT 161.920 29.840 162.240 30.160 ;
        RECT 162.320 29.840 162.640 30.160 ;
        RECT 162.720 29.840 163.040 30.160 ;
        RECT 163.120 29.840 163.440 30.160 ;
        RECT 163.520 29.840 163.840 30.160 ;
        RECT 163.920 29.840 164.240 30.160 ;
        RECT 164.320 29.840 164.640 30.160 ;
        RECT 164.720 29.840 165.040 30.160 ;
        RECT 165.120 29.840 165.440 30.160 ;
        RECT 165.520 29.840 165.840 30.160 ;
        RECT 165.920 29.840 166.240 30.160 ;
        RECT 166.320 29.840 166.640 30.160 ;
        RECT 166.720 29.840 167.040 30.160 ;
        RECT 167.120 29.840 167.440 30.160 ;
        RECT 167.520 29.840 167.840 30.160 ;
        RECT 167.920 29.840 168.240 30.160 ;
        RECT 168.320 29.840 168.640 30.160 ;
        RECT 168.720 29.840 169.040 30.160 ;
        RECT 169.120 29.840 169.440 30.160 ;
        RECT 169.520 29.840 169.840 30.160 ;
        RECT 169.920 29.840 170.240 30.160 ;
        RECT 170.320 29.840 170.640 30.160 ;
        RECT 170.720 29.840 171.040 30.160 ;
        RECT 171.120 29.840 171.440 30.160 ;
        RECT 171.520 29.840 171.840 30.160 ;
        RECT 171.920 29.840 172.240 30.160 ;
        RECT 172.320 29.840 172.640 30.160 ;
        RECT 172.720 29.840 173.040 30.160 ;
        RECT 173.120 29.840 173.440 30.160 ;
        RECT 173.520 29.840 173.840 30.160 ;
        RECT 173.920 29.840 174.240 30.160 ;
        RECT 174.320 29.840 174.640 30.160 ;
        RECT 174.720 29.840 175.040 30.160 ;
        RECT 175.120 29.840 175.440 30.160 ;
        RECT 175.520 29.840 175.840 30.160 ;
        RECT 175.920 29.840 176.240 30.160 ;
        RECT 176.320 29.840 176.640 30.160 ;
        RECT 176.720 29.840 177.040 30.160 ;
        RECT 177.120 29.840 177.440 30.160 ;
        RECT 177.520 29.840 177.840 30.160 ;
        RECT 177.920 29.840 178.240 30.160 ;
        RECT 178.320 29.840 178.640 30.160 ;
        RECT 178.720 29.840 179.040 30.160 ;
        RECT 179.120 29.840 179.440 30.160 ;
        RECT 179.520 29.840 179.840 30.160 ;
        RECT 179.920 29.840 180.240 30.160 ;
        RECT 180.320 29.840 180.640 30.160 ;
        RECT 25.040 29.440 25.360 29.760 ;
        RECT 25.440 29.440 25.760 29.760 ;
        RECT 25.840 29.440 26.160 29.760 ;
        RECT 26.240 29.440 26.560 29.760 ;
        RECT 26.640 29.440 26.960 29.760 ;
        RECT 27.040 29.440 27.360 29.760 ;
        RECT 27.440 29.440 27.760 29.760 ;
        RECT 27.840 29.440 28.160 29.760 ;
        RECT 28.240 29.440 28.560 29.760 ;
        RECT 28.640 29.440 28.960 29.760 ;
        RECT 29.040 29.440 29.360 29.760 ;
        RECT 29.440 29.440 29.760 29.760 ;
        RECT 29.840 29.440 30.160 29.760 ;
        RECT 30.240 29.440 30.560 29.760 ;
        RECT 30.640 29.440 30.960 29.760 ;
        RECT 31.040 29.440 31.360 29.760 ;
        RECT 31.440 29.440 31.760 29.760 ;
        RECT 31.840 29.440 32.160 29.760 ;
        RECT 32.240 29.440 32.560 29.760 ;
        RECT 32.640 29.440 32.960 29.760 ;
        RECT 33.040 29.440 33.360 29.760 ;
        RECT 33.440 29.440 33.760 29.760 ;
        RECT 33.840 29.440 34.160 29.760 ;
        RECT 34.240 29.440 34.560 29.760 ;
        RECT 34.640 29.440 34.960 29.760 ;
        RECT 35.040 29.440 35.360 29.760 ;
        RECT 35.440 29.440 35.760 29.760 ;
        RECT 35.840 29.440 36.160 29.760 ;
        RECT 36.240 29.440 36.560 29.760 ;
        RECT 36.640 29.440 36.960 29.760 ;
        RECT 37.040 29.440 37.360 29.760 ;
        RECT 37.440 29.440 37.760 29.760 ;
        RECT 37.840 29.440 38.160 29.760 ;
        RECT 38.240 29.440 38.560 29.760 ;
        RECT 38.640 29.440 38.960 29.760 ;
        RECT 39.040 29.440 39.360 29.760 ;
        RECT 39.440 29.440 39.760 29.760 ;
        RECT 39.840 29.440 40.160 29.760 ;
        RECT 40.240 29.440 40.560 29.760 ;
        RECT 40.640 29.440 40.960 29.760 ;
        RECT 41.040 29.440 41.360 29.760 ;
        RECT 41.440 29.440 41.760 29.760 ;
        RECT 41.840 29.440 42.160 29.760 ;
        RECT 42.240 29.440 42.560 29.760 ;
        RECT 42.640 29.440 42.960 29.760 ;
        RECT 43.040 29.440 43.360 29.760 ;
        RECT 43.440 29.440 43.760 29.760 ;
        RECT 43.840 29.440 44.160 29.760 ;
        RECT 44.240 29.440 44.560 29.760 ;
        RECT 44.640 29.440 44.960 29.760 ;
        RECT 70.560 29.440 70.880 29.760 ;
        RECT 70.960 29.440 71.280 29.760 ;
        RECT 71.360 29.440 71.680 29.760 ;
        RECT 71.760 29.440 72.080 29.760 ;
        RECT 120.560 29.440 120.880 29.760 ;
        RECT 120.960 29.440 121.280 29.760 ;
        RECT 121.360 29.440 121.680 29.760 ;
        RECT 121.760 29.440 122.080 29.760 ;
        RECT 160.720 29.440 161.040 29.760 ;
        RECT 161.120 29.440 161.440 29.760 ;
        RECT 161.520 29.440 161.840 29.760 ;
        RECT 161.920 29.440 162.240 29.760 ;
        RECT 162.320 29.440 162.640 29.760 ;
        RECT 162.720 29.440 163.040 29.760 ;
        RECT 163.120 29.440 163.440 29.760 ;
        RECT 163.520 29.440 163.840 29.760 ;
        RECT 163.920 29.440 164.240 29.760 ;
        RECT 164.320 29.440 164.640 29.760 ;
        RECT 164.720 29.440 165.040 29.760 ;
        RECT 165.120 29.440 165.440 29.760 ;
        RECT 165.520 29.440 165.840 29.760 ;
        RECT 165.920 29.440 166.240 29.760 ;
        RECT 166.320 29.440 166.640 29.760 ;
        RECT 166.720 29.440 167.040 29.760 ;
        RECT 167.120 29.440 167.440 29.760 ;
        RECT 167.520 29.440 167.840 29.760 ;
        RECT 167.920 29.440 168.240 29.760 ;
        RECT 168.320 29.440 168.640 29.760 ;
        RECT 168.720 29.440 169.040 29.760 ;
        RECT 169.120 29.440 169.440 29.760 ;
        RECT 169.520 29.440 169.840 29.760 ;
        RECT 169.920 29.440 170.240 29.760 ;
        RECT 170.320 29.440 170.640 29.760 ;
        RECT 170.720 29.440 171.040 29.760 ;
        RECT 171.120 29.440 171.440 29.760 ;
        RECT 171.520 29.440 171.840 29.760 ;
        RECT 171.920 29.440 172.240 29.760 ;
        RECT 172.320 29.440 172.640 29.760 ;
        RECT 172.720 29.440 173.040 29.760 ;
        RECT 173.120 29.440 173.440 29.760 ;
        RECT 173.520 29.440 173.840 29.760 ;
        RECT 173.920 29.440 174.240 29.760 ;
        RECT 174.320 29.440 174.640 29.760 ;
        RECT 174.720 29.440 175.040 29.760 ;
        RECT 175.120 29.440 175.440 29.760 ;
        RECT 175.520 29.440 175.840 29.760 ;
        RECT 175.920 29.440 176.240 29.760 ;
        RECT 176.320 29.440 176.640 29.760 ;
        RECT 176.720 29.440 177.040 29.760 ;
        RECT 177.120 29.440 177.440 29.760 ;
        RECT 177.520 29.440 177.840 29.760 ;
        RECT 177.920 29.440 178.240 29.760 ;
        RECT 178.320 29.440 178.640 29.760 ;
        RECT 178.720 29.440 179.040 29.760 ;
        RECT 179.120 29.440 179.440 29.760 ;
        RECT 179.520 29.440 179.840 29.760 ;
        RECT 179.920 29.440 180.240 29.760 ;
        RECT 180.320 29.440 180.640 29.760 ;
        RECT 25.040 29.040 25.360 29.360 ;
        RECT 25.440 29.040 25.760 29.360 ;
        RECT 25.840 29.040 26.160 29.360 ;
        RECT 26.240 29.040 26.560 29.360 ;
        RECT 26.640 29.040 26.960 29.360 ;
        RECT 27.040 29.040 27.360 29.360 ;
        RECT 27.440 29.040 27.760 29.360 ;
        RECT 27.840 29.040 28.160 29.360 ;
        RECT 28.240 29.040 28.560 29.360 ;
        RECT 28.640 29.040 28.960 29.360 ;
        RECT 29.040 29.040 29.360 29.360 ;
        RECT 29.440 29.040 29.760 29.360 ;
        RECT 29.840 29.040 30.160 29.360 ;
        RECT 30.240 29.040 30.560 29.360 ;
        RECT 30.640 29.040 30.960 29.360 ;
        RECT 31.040 29.040 31.360 29.360 ;
        RECT 31.440 29.040 31.760 29.360 ;
        RECT 31.840 29.040 32.160 29.360 ;
        RECT 32.240 29.040 32.560 29.360 ;
        RECT 32.640 29.040 32.960 29.360 ;
        RECT 33.040 29.040 33.360 29.360 ;
        RECT 33.440 29.040 33.760 29.360 ;
        RECT 33.840 29.040 34.160 29.360 ;
        RECT 34.240 29.040 34.560 29.360 ;
        RECT 34.640 29.040 34.960 29.360 ;
        RECT 35.040 29.040 35.360 29.360 ;
        RECT 35.440 29.040 35.760 29.360 ;
        RECT 35.840 29.040 36.160 29.360 ;
        RECT 36.240 29.040 36.560 29.360 ;
        RECT 36.640 29.040 36.960 29.360 ;
        RECT 37.040 29.040 37.360 29.360 ;
        RECT 37.440 29.040 37.760 29.360 ;
        RECT 37.840 29.040 38.160 29.360 ;
        RECT 38.240 29.040 38.560 29.360 ;
        RECT 38.640 29.040 38.960 29.360 ;
        RECT 39.040 29.040 39.360 29.360 ;
        RECT 39.440 29.040 39.760 29.360 ;
        RECT 39.840 29.040 40.160 29.360 ;
        RECT 40.240 29.040 40.560 29.360 ;
        RECT 40.640 29.040 40.960 29.360 ;
        RECT 41.040 29.040 41.360 29.360 ;
        RECT 41.440 29.040 41.760 29.360 ;
        RECT 41.840 29.040 42.160 29.360 ;
        RECT 42.240 29.040 42.560 29.360 ;
        RECT 42.640 29.040 42.960 29.360 ;
        RECT 43.040 29.040 43.360 29.360 ;
        RECT 43.440 29.040 43.760 29.360 ;
        RECT 43.840 29.040 44.160 29.360 ;
        RECT 44.240 29.040 44.560 29.360 ;
        RECT 44.640 29.040 44.960 29.360 ;
        RECT 70.560 29.040 70.880 29.360 ;
        RECT 70.960 29.040 71.280 29.360 ;
        RECT 71.360 29.040 71.680 29.360 ;
        RECT 71.760 29.040 72.080 29.360 ;
        RECT 120.560 29.040 120.880 29.360 ;
        RECT 120.960 29.040 121.280 29.360 ;
        RECT 121.360 29.040 121.680 29.360 ;
        RECT 121.760 29.040 122.080 29.360 ;
        RECT 160.720 29.040 161.040 29.360 ;
        RECT 161.120 29.040 161.440 29.360 ;
        RECT 161.520 29.040 161.840 29.360 ;
        RECT 161.920 29.040 162.240 29.360 ;
        RECT 162.320 29.040 162.640 29.360 ;
        RECT 162.720 29.040 163.040 29.360 ;
        RECT 163.120 29.040 163.440 29.360 ;
        RECT 163.520 29.040 163.840 29.360 ;
        RECT 163.920 29.040 164.240 29.360 ;
        RECT 164.320 29.040 164.640 29.360 ;
        RECT 164.720 29.040 165.040 29.360 ;
        RECT 165.120 29.040 165.440 29.360 ;
        RECT 165.520 29.040 165.840 29.360 ;
        RECT 165.920 29.040 166.240 29.360 ;
        RECT 166.320 29.040 166.640 29.360 ;
        RECT 166.720 29.040 167.040 29.360 ;
        RECT 167.120 29.040 167.440 29.360 ;
        RECT 167.520 29.040 167.840 29.360 ;
        RECT 167.920 29.040 168.240 29.360 ;
        RECT 168.320 29.040 168.640 29.360 ;
        RECT 168.720 29.040 169.040 29.360 ;
        RECT 169.120 29.040 169.440 29.360 ;
        RECT 169.520 29.040 169.840 29.360 ;
        RECT 169.920 29.040 170.240 29.360 ;
        RECT 170.320 29.040 170.640 29.360 ;
        RECT 170.720 29.040 171.040 29.360 ;
        RECT 171.120 29.040 171.440 29.360 ;
        RECT 171.520 29.040 171.840 29.360 ;
        RECT 171.920 29.040 172.240 29.360 ;
        RECT 172.320 29.040 172.640 29.360 ;
        RECT 172.720 29.040 173.040 29.360 ;
        RECT 173.120 29.040 173.440 29.360 ;
        RECT 173.520 29.040 173.840 29.360 ;
        RECT 173.920 29.040 174.240 29.360 ;
        RECT 174.320 29.040 174.640 29.360 ;
        RECT 174.720 29.040 175.040 29.360 ;
        RECT 175.120 29.040 175.440 29.360 ;
        RECT 175.520 29.040 175.840 29.360 ;
        RECT 175.920 29.040 176.240 29.360 ;
        RECT 176.320 29.040 176.640 29.360 ;
        RECT 176.720 29.040 177.040 29.360 ;
        RECT 177.120 29.040 177.440 29.360 ;
        RECT 177.520 29.040 177.840 29.360 ;
        RECT 177.920 29.040 178.240 29.360 ;
        RECT 178.320 29.040 178.640 29.360 ;
        RECT 178.720 29.040 179.040 29.360 ;
        RECT 179.120 29.040 179.440 29.360 ;
        RECT 179.520 29.040 179.840 29.360 ;
        RECT 179.920 29.040 180.240 29.360 ;
        RECT 180.320 29.040 180.640 29.360 ;
        RECT 25.040 28.640 25.360 28.960 ;
        RECT 25.440 28.640 25.760 28.960 ;
        RECT 25.840 28.640 26.160 28.960 ;
        RECT 26.240 28.640 26.560 28.960 ;
        RECT 26.640 28.640 26.960 28.960 ;
        RECT 27.040 28.640 27.360 28.960 ;
        RECT 27.440 28.640 27.760 28.960 ;
        RECT 27.840 28.640 28.160 28.960 ;
        RECT 28.240 28.640 28.560 28.960 ;
        RECT 28.640 28.640 28.960 28.960 ;
        RECT 29.040 28.640 29.360 28.960 ;
        RECT 29.440 28.640 29.760 28.960 ;
        RECT 29.840 28.640 30.160 28.960 ;
        RECT 30.240 28.640 30.560 28.960 ;
        RECT 30.640 28.640 30.960 28.960 ;
        RECT 31.040 28.640 31.360 28.960 ;
        RECT 31.440 28.640 31.760 28.960 ;
        RECT 31.840 28.640 32.160 28.960 ;
        RECT 32.240 28.640 32.560 28.960 ;
        RECT 32.640 28.640 32.960 28.960 ;
        RECT 33.040 28.640 33.360 28.960 ;
        RECT 33.440 28.640 33.760 28.960 ;
        RECT 33.840 28.640 34.160 28.960 ;
        RECT 34.240 28.640 34.560 28.960 ;
        RECT 34.640 28.640 34.960 28.960 ;
        RECT 35.040 28.640 35.360 28.960 ;
        RECT 35.440 28.640 35.760 28.960 ;
        RECT 35.840 28.640 36.160 28.960 ;
        RECT 36.240 28.640 36.560 28.960 ;
        RECT 36.640 28.640 36.960 28.960 ;
        RECT 37.040 28.640 37.360 28.960 ;
        RECT 37.440 28.640 37.760 28.960 ;
        RECT 37.840 28.640 38.160 28.960 ;
        RECT 38.240 28.640 38.560 28.960 ;
        RECT 38.640 28.640 38.960 28.960 ;
        RECT 39.040 28.640 39.360 28.960 ;
        RECT 39.440 28.640 39.760 28.960 ;
        RECT 39.840 28.640 40.160 28.960 ;
        RECT 40.240 28.640 40.560 28.960 ;
        RECT 40.640 28.640 40.960 28.960 ;
        RECT 41.040 28.640 41.360 28.960 ;
        RECT 41.440 28.640 41.760 28.960 ;
        RECT 41.840 28.640 42.160 28.960 ;
        RECT 42.240 28.640 42.560 28.960 ;
        RECT 42.640 28.640 42.960 28.960 ;
        RECT 43.040 28.640 43.360 28.960 ;
        RECT 43.440 28.640 43.760 28.960 ;
        RECT 43.840 28.640 44.160 28.960 ;
        RECT 44.240 28.640 44.560 28.960 ;
        RECT 44.640 28.640 44.960 28.960 ;
        RECT 70.560 28.640 70.880 28.960 ;
        RECT 70.960 28.640 71.280 28.960 ;
        RECT 71.360 28.640 71.680 28.960 ;
        RECT 71.760 28.640 72.080 28.960 ;
        RECT 120.560 28.640 120.880 28.960 ;
        RECT 120.960 28.640 121.280 28.960 ;
        RECT 121.360 28.640 121.680 28.960 ;
        RECT 121.760 28.640 122.080 28.960 ;
        RECT 160.720 28.640 161.040 28.960 ;
        RECT 161.120 28.640 161.440 28.960 ;
        RECT 161.520 28.640 161.840 28.960 ;
        RECT 161.920 28.640 162.240 28.960 ;
        RECT 162.320 28.640 162.640 28.960 ;
        RECT 162.720 28.640 163.040 28.960 ;
        RECT 163.120 28.640 163.440 28.960 ;
        RECT 163.520 28.640 163.840 28.960 ;
        RECT 163.920 28.640 164.240 28.960 ;
        RECT 164.320 28.640 164.640 28.960 ;
        RECT 164.720 28.640 165.040 28.960 ;
        RECT 165.120 28.640 165.440 28.960 ;
        RECT 165.520 28.640 165.840 28.960 ;
        RECT 165.920 28.640 166.240 28.960 ;
        RECT 166.320 28.640 166.640 28.960 ;
        RECT 166.720 28.640 167.040 28.960 ;
        RECT 167.120 28.640 167.440 28.960 ;
        RECT 167.520 28.640 167.840 28.960 ;
        RECT 167.920 28.640 168.240 28.960 ;
        RECT 168.320 28.640 168.640 28.960 ;
        RECT 168.720 28.640 169.040 28.960 ;
        RECT 169.120 28.640 169.440 28.960 ;
        RECT 169.520 28.640 169.840 28.960 ;
        RECT 169.920 28.640 170.240 28.960 ;
        RECT 170.320 28.640 170.640 28.960 ;
        RECT 170.720 28.640 171.040 28.960 ;
        RECT 171.120 28.640 171.440 28.960 ;
        RECT 171.520 28.640 171.840 28.960 ;
        RECT 171.920 28.640 172.240 28.960 ;
        RECT 172.320 28.640 172.640 28.960 ;
        RECT 172.720 28.640 173.040 28.960 ;
        RECT 173.120 28.640 173.440 28.960 ;
        RECT 173.520 28.640 173.840 28.960 ;
        RECT 173.920 28.640 174.240 28.960 ;
        RECT 174.320 28.640 174.640 28.960 ;
        RECT 174.720 28.640 175.040 28.960 ;
        RECT 175.120 28.640 175.440 28.960 ;
        RECT 175.520 28.640 175.840 28.960 ;
        RECT 175.920 28.640 176.240 28.960 ;
        RECT 176.320 28.640 176.640 28.960 ;
        RECT 176.720 28.640 177.040 28.960 ;
        RECT 177.120 28.640 177.440 28.960 ;
        RECT 177.520 28.640 177.840 28.960 ;
        RECT 177.920 28.640 178.240 28.960 ;
        RECT 178.320 28.640 178.640 28.960 ;
        RECT 178.720 28.640 179.040 28.960 ;
        RECT 179.120 28.640 179.440 28.960 ;
        RECT 179.520 28.640 179.840 28.960 ;
        RECT 179.920 28.640 180.240 28.960 ;
        RECT 180.320 28.640 180.640 28.960 ;
        RECT 25.040 28.240 25.360 28.560 ;
        RECT 25.440 28.240 25.760 28.560 ;
        RECT 25.840 28.240 26.160 28.560 ;
        RECT 26.240 28.240 26.560 28.560 ;
        RECT 26.640 28.240 26.960 28.560 ;
        RECT 27.040 28.240 27.360 28.560 ;
        RECT 27.440 28.240 27.760 28.560 ;
        RECT 27.840 28.240 28.160 28.560 ;
        RECT 28.240 28.240 28.560 28.560 ;
        RECT 28.640 28.240 28.960 28.560 ;
        RECT 29.040 28.240 29.360 28.560 ;
        RECT 29.440 28.240 29.760 28.560 ;
        RECT 29.840 28.240 30.160 28.560 ;
        RECT 30.240 28.240 30.560 28.560 ;
        RECT 30.640 28.240 30.960 28.560 ;
        RECT 31.040 28.240 31.360 28.560 ;
        RECT 31.440 28.240 31.760 28.560 ;
        RECT 31.840 28.240 32.160 28.560 ;
        RECT 32.240 28.240 32.560 28.560 ;
        RECT 32.640 28.240 32.960 28.560 ;
        RECT 33.040 28.240 33.360 28.560 ;
        RECT 33.440 28.240 33.760 28.560 ;
        RECT 33.840 28.240 34.160 28.560 ;
        RECT 34.240 28.240 34.560 28.560 ;
        RECT 34.640 28.240 34.960 28.560 ;
        RECT 35.040 28.240 35.360 28.560 ;
        RECT 35.440 28.240 35.760 28.560 ;
        RECT 35.840 28.240 36.160 28.560 ;
        RECT 36.240 28.240 36.560 28.560 ;
        RECT 36.640 28.240 36.960 28.560 ;
        RECT 37.040 28.240 37.360 28.560 ;
        RECT 37.440 28.240 37.760 28.560 ;
        RECT 37.840 28.240 38.160 28.560 ;
        RECT 38.240 28.240 38.560 28.560 ;
        RECT 38.640 28.240 38.960 28.560 ;
        RECT 39.040 28.240 39.360 28.560 ;
        RECT 39.440 28.240 39.760 28.560 ;
        RECT 39.840 28.240 40.160 28.560 ;
        RECT 40.240 28.240 40.560 28.560 ;
        RECT 40.640 28.240 40.960 28.560 ;
        RECT 41.040 28.240 41.360 28.560 ;
        RECT 41.440 28.240 41.760 28.560 ;
        RECT 41.840 28.240 42.160 28.560 ;
        RECT 42.240 28.240 42.560 28.560 ;
        RECT 42.640 28.240 42.960 28.560 ;
        RECT 43.040 28.240 43.360 28.560 ;
        RECT 43.440 28.240 43.760 28.560 ;
        RECT 43.840 28.240 44.160 28.560 ;
        RECT 44.240 28.240 44.560 28.560 ;
        RECT 44.640 28.240 44.960 28.560 ;
        RECT 70.560 28.240 70.880 28.560 ;
        RECT 70.960 28.240 71.280 28.560 ;
        RECT 71.360 28.240 71.680 28.560 ;
        RECT 71.760 28.240 72.080 28.560 ;
        RECT 120.560 28.240 120.880 28.560 ;
        RECT 120.960 28.240 121.280 28.560 ;
        RECT 121.360 28.240 121.680 28.560 ;
        RECT 121.760 28.240 122.080 28.560 ;
        RECT 160.720 28.240 161.040 28.560 ;
        RECT 161.120 28.240 161.440 28.560 ;
        RECT 161.520 28.240 161.840 28.560 ;
        RECT 161.920 28.240 162.240 28.560 ;
        RECT 162.320 28.240 162.640 28.560 ;
        RECT 162.720 28.240 163.040 28.560 ;
        RECT 163.120 28.240 163.440 28.560 ;
        RECT 163.520 28.240 163.840 28.560 ;
        RECT 163.920 28.240 164.240 28.560 ;
        RECT 164.320 28.240 164.640 28.560 ;
        RECT 164.720 28.240 165.040 28.560 ;
        RECT 165.120 28.240 165.440 28.560 ;
        RECT 165.520 28.240 165.840 28.560 ;
        RECT 165.920 28.240 166.240 28.560 ;
        RECT 166.320 28.240 166.640 28.560 ;
        RECT 166.720 28.240 167.040 28.560 ;
        RECT 167.120 28.240 167.440 28.560 ;
        RECT 167.520 28.240 167.840 28.560 ;
        RECT 167.920 28.240 168.240 28.560 ;
        RECT 168.320 28.240 168.640 28.560 ;
        RECT 168.720 28.240 169.040 28.560 ;
        RECT 169.120 28.240 169.440 28.560 ;
        RECT 169.520 28.240 169.840 28.560 ;
        RECT 169.920 28.240 170.240 28.560 ;
        RECT 170.320 28.240 170.640 28.560 ;
        RECT 170.720 28.240 171.040 28.560 ;
        RECT 171.120 28.240 171.440 28.560 ;
        RECT 171.520 28.240 171.840 28.560 ;
        RECT 171.920 28.240 172.240 28.560 ;
        RECT 172.320 28.240 172.640 28.560 ;
        RECT 172.720 28.240 173.040 28.560 ;
        RECT 173.120 28.240 173.440 28.560 ;
        RECT 173.520 28.240 173.840 28.560 ;
        RECT 173.920 28.240 174.240 28.560 ;
        RECT 174.320 28.240 174.640 28.560 ;
        RECT 174.720 28.240 175.040 28.560 ;
        RECT 175.120 28.240 175.440 28.560 ;
        RECT 175.520 28.240 175.840 28.560 ;
        RECT 175.920 28.240 176.240 28.560 ;
        RECT 176.320 28.240 176.640 28.560 ;
        RECT 176.720 28.240 177.040 28.560 ;
        RECT 177.120 28.240 177.440 28.560 ;
        RECT 177.520 28.240 177.840 28.560 ;
        RECT 177.920 28.240 178.240 28.560 ;
        RECT 178.320 28.240 178.640 28.560 ;
        RECT 178.720 28.240 179.040 28.560 ;
        RECT 179.120 28.240 179.440 28.560 ;
        RECT 179.520 28.240 179.840 28.560 ;
        RECT 179.920 28.240 180.240 28.560 ;
        RECT 180.320 28.240 180.640 28.560 ;
        RECT 25.040 27.840 25.360 28.160 ;
        RECT 25.440 27.840 25.760 28.160 ;
        RECT 25.840 27.840 26.160 28.160 ;
        RECT 26.240 27.840 26.560 28.160 ;
        RECT 26.640 27.840 26.960 28.160 ;
        RECT 27.040 27.840 27.360 28.160 ;
        RECT 27.440 27.840 27.760 28.160 ;
        RECT 27.840 27.840 28.160 28.160 ;
        RECT 28.240 27.840 28.560 28.160 ;
        RECT 28.640 27.840 28.960 28.160 ;
        RECT 29.040 27.840 29.360 28.160 ;
        RECT 29.440 27.840 29.760 28.160 ;
        RECT 29.840 27.840 30.160 28.160 ;
        RECT 30.240 27.840 30.560 28.160 ;
        RECT 30.640 27.840 30.960 28.160 ;
        RECT 31.040 27.840 31.360 28.160 ;
        RECT 31.440 27.840 31.760 28.160 ;
        RECT 31.840 27.840 32.160 28.160 ;
        RECT 32.240 27.840 32.560 28.160 ;
        RECT 32.640 27.840 32.960 28.160 ;
        RECT 33.040 27.840 33.360 28.160 ;
        RECT 33.440 27.840 33.760 28.160 ;
        RECT 33.840 27.840 34.160 28.160 ;
        RECT 34.240 27.840 34.560 28.160 ;
        RECT 34.640 27.840 34.960 28.160 ;
        RECT 35.040 27.840 35.360 28.160 ;
        RECT 35.440 27.840 35.760 28.160 ;
        RECT 35.840 27.840 36.160 28.160 ;
        RECT 36.240 27.840 36.560 28.160 ;
        RECT 36.640 27.840 36.960 28.160 ;
        RECT 37.040 27.840 37.360 28.160 ;
        RECT 37.440 27.840 37.760 28.160 ;
        RECT 37.840 27.840 38.160 28.160 ;
        RECT 38.240 27.840 38.560 28.160 ;
        RECT 38.640 27.840 38.960 28.160 ;
        RECT 39.040 27.840 39.360 28.160 ;
        RECT 39.440 27.840 39.760 28.160 ;
        RECT 39.840 27.840 40.160 28.160 ;
        RECT 40.240 27.840 40.560 28.160 ;
        RECT 40.640 27.840 40.960 28.160 ;
        RECT 41.040 27.840 41.360 28.160 ;
        RECT 41.440 27.840 41.760 28.160 ;
        RECT 41.840 27.840 42.160 28.160 ;
        RECT 42.240 27.840 42.560 28.160 ;
        RECT 42.640 27.840 42.960 28.160 ;
        RECT 43.040 27.840 43.360 28.160 ;
        RECT 43.440 27.840 43.760 28.160 ;
        RECT 43.840 27.840 44.160 28.160 ;
        RECT 44.240 27.840 44.560 28.160 ;
        RECT 44.640 27.840 44.960 28.160 ;
        RECT 70.560 27.840 70.880 28.160 ;
        RECT 70.960 27.840 71.280 28.160 ;
        RECT 71.360 27.840 71.680 28.160 ;
        RECT 71.760 27.840 72.080 28.160 ;
        RECT 120.560 27.840 120.880 28.160 ;
        RECT 120.960 27.840 121.280 28.160 ;
        RECT 121.360 27.840 121.680 28.160 ;
        RECT 121.760 27.840 122.080 28.160 ;
        RECT 160.720 27.840 161.040 28.160 ;
        RECT 161.120 27.840 161.440 28.160 ;
        RECT 161.520 27.840 161.840 28.160 ;
        RECT 161.920 27.840 162.240 28.160 ;
        RECT 162.320 27.840 162.640 28.160 ;
        RECT 162.720 27.840 163.040 28.160 ;
        RECT 163.120 27.840 163.440 28.160 ;
        RECT 163.520 27.840 163.840 28.160 ;
        RECT 163.920 27.840 164.240 28.160 ;
        RECT 164.320 27.840 164.640 28.160 ;
        RECT 164.720 27.840 165.040 28.160 ;
        RECT 165.120 27.840 165.440 28.160 ;
        RECT 165.520 27.840 165.840 28.160 ;
        RECT 165.920 27.840 166.240 28.160 ;
        RECT 166.320 27.840 166.640 28.160 ;
        RECT 166.720 27.840 167.040 28.160 ;
        RECT 167.120 27.840 167.440 28.160 ;
        RECT 167.520 27.840 167.840 28.160 ;
        RECT 167.920 27.840 168.240 28.160 ;
        RECT 168.320 27.840 168.640 28.160 ;
        RECT 168.720 27.840 169.040 28.160 ;
        RECT 169.120 27.840 169.440 28.160 ;
        RECT 169.520 27.840 169.840 28.160 ;
        RECT 169.920 27.840 170.240 28.160 ;
        RECT 170.320 27.840 170.640 28.160 ;
        RECT 170.720 27.840 171.040 28.160 ;
        RECT 171.120 27.840 171.440 28.160 ;
        RECT 171.520 27.840 171.840 28.160 ;
        RECT 171.920 27.840 172.240 28.160 ;
        RECT 172.320 27.840 172.640 28.160 ;
        RECT 172.720 27.840 173.040 28.160 ;
        RECT 173.120 27.840 173.440 28.160 ;
        RECT 173.520 27.840 173.840 28.160 ;
        RECT 173.920 27.840 174.240 28.160 ;
        RECT 174.320 27.840 174.640 28.160 ;
        RECT 174.720 27.840 175.040 28.160 ;
        RECT 175.120 27.840 175.440 28.160 ;
        RECT 175.520 27.840 175.840 28.160 ;
        RECT 175.920 27.840 176.240 28.160 ;
        RECT 176.320 27.840 176.640 28.160 ;
        RECT 176.720 27.840 177.040 28.160 ;
        RECT 177.120 27.840 177.440 28.160 ;
        RECT 177.520 27.840 177.840 28.160 ;
        RECT 177.920 27.840 178.240 28.160 ;
        RECT 178.320 27.840 178.640 28.160 ;
        RECT 178.720 27.840 179.040 28.160 ;
        RECT 179.120 27.840 179.440 28.160 ;
        RECT 179.520 27.840 179.840 28.160 ;
        RECT 179.920 27.840 180.240 28.160 ;
        RECT 180.320 27.840 180.640 28.160 ;
        RECT 25.040 27.440 25.360 27.760 ;
        RECT 25.440 27.440 25.760 27.760 ;
        RECT 25.840 27.440 26.160 27.760 ;
        RECT 26.240 27.440 26.560 27.760 ;
        RECT 26.640 27.440 26.960 27.760 ;
        RECT 27.040 27.440 27.360 27.760 ;
        RECT 27.440 27.440 27.760 27.760 ;
        RECT 27.840 27.440 28.160 27.760 ;
        RECT 28.240 27.440 28.560 27.760 ;
        RECT 28.640 27.440 28.960 27.760 ;
        RECT 29.040 27.440 29.360 27.760 ;
        RECT 29.440 27.440 29.760 27.760 ;
        RECT 29.840 27.440 30.160 27.760 ;
        RECT 30.240 27.440 30.560 27.760 ;
        RECT 30.640 27.440 30.960 27.760 ;
        RECT 31.040 27.440 31.360 27.760 ;
        RECT 31.440 27.440 31.760 27.760 ;
        RECT 31.840 27.440 32.160 27.760 ;
        RECT 32.240 27.440 32.560 27.760 ;
        RECT 32.640 27.440 32.960 27.760 ;
        RECT 33.040 27.440 33.360 27.760 ;
        RECT 33.440 27.440 33.760 27.760 ;
        RECT 33.840 27.440 34.160 27.760 ;
        RECT 34.240 27.440 34.560 27.760 ;
        RECT 34.640 27.440 34.960 27.760 ;
        RECT 35.040 27.440 35.360 27.760 ;
        RECT 35.440 27.440 35.760 27.760 ;
        RECT 35.840 27.440 36.160 27.760 ;
        RECT 36.240 27.440 36.560 27.760 ;
        RECT 36.640 27.440 36.960 27.760 ;
        RECT 37.040 27.440 37.360 27.760 ;
        RECT 37.440 27.440 37.760 27.760 ;
        RECT 37.840 27.440 38.160 27.760 ;
        RECT 38.240 27.440 38.560 27.760 ;
        RECT 38.640 27.440 38.960 27.760 ;
        RECT 39.040 27.440 39.360 27.760 ;
        RECT 39.440 27.440 39.760 27.760 ;
        RECT 39.840 27.440 40.160 27.760 ;
        RECT 40.240 27.440 40.560 27.760 ;
        RECT 40.640 27.440 40.960 27.760 ;
        RECT 41.040 27.440 41.360 27.760 ;
        RECT 41.440 27.440 41.760 27.760 ;
        RECT 41.840 27.440 42.160 27.760 ;
        RECT 42.240 27.440 42.560 27.760 ;
        RECT 42.640 27.440 42.960 27.760 ;
        RECT 43.040 27.440 43.360 27.760 ;
        RECT 43.440 27.440 43.760 27.760 ;
        RECT 43.840 27.440 44.160 27.760 ;
        RECT 44.240 27.440 44.560 27.760 ;
        RECT 44.640 27.440 44.960 27.760 ;
        RECT 70.560 27.440 70.880 27.760 ;
        RECT 70.960 27.440 71.280 27.760 ;
        RECT 71.360 27.440 71.680 27.760 ;
        RECT 71.760 27.440 72.080 27.760 ;
        RECT 120.560 27.440 120.880 27.760 ;
        RECT 120.960 27.440 121.280 27.760 ;
        RECT 121.360 27.440 121.680 27.760 ;
        RECT 121.760 27.440 122.080 27.760 ;
        RECT 160.720 27.440 161.040 27.760 ;
        RECT 161.120 27.440 161.440 27.760 ;
        RECT 161.520 27.440 161.840 27.760 ;
        RECT 161.920 27.440 162.240 27.760 ;
        RECT 162.320 27.440 162.640 27.760 ;
        RECT 162.720 27.440 163.040 27.760 ;
        RECT 163.120 27.440 163.440 27.760 ;
        RECT 163.520 27.440 163.840 27.760 ;
        RECT 163.920 27.440 164.240 27.760 ;
        RECT 164.320 27.440 164.640 27.760 ;
        RECT 164.720 27.440 165.040 27.760 ;
        RECT 165.120 27.440 165.440 27.760 ;
        RECT 165.520 27.440 165.840 27.760 ;
        RECT 165.920 27.440 166.240 27.760 ;
        RECT 166.320 27.440 166.640 27.760 ;
        RECT 166.720 27.440 167.040 27.760 ;
        RECT 167.120 27.440 167.440 27.760 ;
        RECT 167.520 27.440 167.840 27.760 ;
        RECT 167.920 27.440 168.240 27.760 ;
        RECT 168.320 27.440 168.640 27.760 ;
        RECT 168.720 27.440 169.040 27.760 ;
        RECT 169.120 27.440 169.440 27.760 ;
        RECT 169.520 27.440 169.840 27.760 ;
        RECT 169.920 27.440 170.240 27.760 ;
        RECT 170.320 27.440 170.640 27.760 ;
        RECT 170.720 27.440 171.040 27.760 ;
        RECT 171.120 27.440 171.440 27.760 ;
        RECT 171.520 27.440 171.840 27.760 ;
        RECT 171.920 27.440 172.240 27.760 ;
        RECT 172.320 27.440 172.640 27.760 ;
        RECT 172.720 27.440 173.040 27.760 ;
        RECT 173.120 27.440 173.440 27.760 ;
        RECT 173.520 27.440 173.840 27.760 ;
        RECT 173.920 27.440 174.240 27.760 ;
        RECT 174.320 27.440 174.640 27.760 ;
        RECT 174.720 27.440 175.040 27.760 ;
        RECT 175.120 27.440 175.440 27.760 ;
        RECT 175.520 27.440 175.840 27.760 ;
        RECT 175.920 27.440 176.240 27.760 ;
        RECT 176.320 27.440 176.640 27.760 ;
        RECT 176.720 27.440 177.040 27.760 ;
        RECT 177.120 27.440 177.440 27.760 ;
        RECT 177.520 27.440 177.840 27.760 ;
        RECT 177.920 27.440 178.240 27.760 ;
        RECT 178.320 27.440 178.640 27.760 ;
        RECT 178.720 27.440 179.040 27.760 ;
        RECT 179.120 27.440 179.440 27.760 ;
        RECT 179.520 27.440 179.840 27.760 ;
        RECT 179.920 27.440 180.240 27.760 ;
        RECT 180.320 27.440 180.640 27.760 ;
        RECT 25.040 27.040 25.360 27.360 ;
        RECT 25.440 27.040 25.760 27.360 ;
        RECT 25.840 27.040 26.160 27.360 ;
        RECT 26.240 27.040 26.560 27.360 ;
        RECT 26.640 27.040 26.960 27.360 ;
        RECT 27.040 27.040 27.360 27.360 ;
        RECT 27.440 27.040 27.760 27.360 ;
        RECT 27.840 27.040 28.160 27.360 ;
        RECT 28.240 27.040 28.560 27.360 ;
        RECT 28.640 27.040 28.960 27.360 ;
        RECT 29.040 27.040 29.360 27.360 ;
        RECT 29.440 27.040 29.760 27.360 ;
        RECT 29.840 27.040 30.160 27.360 ;
        RECT 30.240 27.040 30.560 27.360 ;
        RECT 30.640 27.040 30.960 27.360 ;
        RECT 31.040 27.040 31.360 27.360 ;
        RECT 31.440 27.040 31.760 27.360 ;
        RECT 31.840 27.040 32.160 27.360 ;
        RECT 32.240 27.040 32.560 27.360 ;
        RECT 32.640 27.040 32.960 27.360 ;
        RECT 33.040 27.040 33.360 27.360 ;
        RECT 33.440 27.040 33.760 27.360 ;
        RECT 33.840 27.040 34.160 27.360 ;
        RECT 34.240 27.040 34.560 27.360 ;
        RECT 34.640 27.040 34.960 27.360 ;
        RECT 35.040 27.040 35.360 27.360 ;
        RECT 35.440 27.040 35.760 27.360 ;
        RECT 35.840 27.040 36.160 27.360 ;
        RECT 36.240 27.040 36.560 27.360 ;
        RECT 36.640 27.040 36.960 27.360 ;
        RECT 37.040 27.040 37.360 27.360 ;
        RECT 37.440 27.040 37.760 27.360 ;
        RECT 37.840 27.040 38.160 27.360 ;
        RECT 38.240 27.040 38.560 27.360 ;
        RECT 38.640 27.040 38.960 27.360 ;
        RECT 39.040 27.040 39.360 27.360 ;
        RECT 39.440 27.040 39.760 27.360 ;
        RECT 39.840 27.040 40.160 27.360 ;
        RECT 40.240 27.040 40.560 27.360 ;
        RECT 40.640 27.040 40.960 27.360 ;
        RECT 41.040 27.040 41.360 27.360 ;
        RECT 41.440 27.040 41.760 27.360 ;
        RECT 41.840 27.040 42.160 27.360 ;
        RECT 42.240 27.040 42.560 27.360 ;
        RECT 42.640 27.040 42.960 27.360 ;
        RECT 43.040 27.040 43.360 27.360 ;
        RECT 43.440 27.040 43.760 27.360 ;
        RECT 43.840 27.040 44.160 27.360 ;
        RECT 44.240 27.040 44.560 27.360 ;
        RECT 44.640 27.040 44.960 27.360 ;
        RECT 70.560 27.040 70.880 27.360 ;
        RECT 70.960 27.040 71.280 27.360 ;
        RECT 71.360 27.040 71.680 27.360 ;
        RECT 71.760 27.040 72.080 27.360 ;
        RECT 120.560 27.040 120.880 27.360 ;
        RECT 120.960 27.040 121.280 27.360 ;
        RECT 121.360 27.040 121.680 27.360 ;
        RECT 121.760 27.040 122.080 27.360 ;
        RECT 160.720 27.040 161.040 27.360 ;
        RECT 161.120 27.040 161.440 27.360 ;
        RECT 161.520 27.040 161.840 27.360 ;
        RECT 161.920 27.040 162.240 27.360 ;
        RECT 162.320 27.040 162.640 27.360 ;
        RECT 162.720 27.040 163.040 27.360 ;
        RECT 163.120 27.040 163.440 27.360 ;
        RECT 163.520 27.040 163.840 27.360 ;
        RECT 163.920 27.040 164.240 27.360 ;
        RECT 164.320 27.040 164.640 27.360 ;
        RECT 164.720 27.040 165.040 27.360 ;
        RECT 165.120 27.040 165.440 27.360 ;
        RECT 165.520 27.040 165.840 27.360 ;
        RECT 165.920 27.040 166.240 27.360 ;
        RECT 166.320 27.040 166.640 27.360 ;
        RECT 166.720 27.040 167.040 27.360 ;
        RECT 167.120 27.040 167.440 27.360 ;
        RECT 167.520 27.040 167.840 27.360 ;
        RECT 167.920 27.040 168.240 27.360 ;
        RECT 168.320 27.040 168.640 27.360 ;
        RECT 168.720 27.040 169.040 27.360 ;
        RECT 169.120 27.040 169.440 27.360 ;
        RECT 169.520 27.040 169.840 27.360 ;
        RECT 169.920 27.040 170.240 27.360 ;
        RECT 170.320 27.040 170.640 27.360 ;
        RECT 170.720 27.040 171.040 27.360 ;
        RECT 171.120 27.040 171.440 27.360 ;
        RECT 171.520 27.040 171.840 27.360 ;
        RECT 171.920 27.040 172.240 27.360 ;
        RECT 172.320 27.040 172.640 27.360 ;
        RECT 172.720 27.040 173.040 27.360 ;
        RECT 173.120 27.040 173.440 27.360 ;
        RECT 173.520 27.040 173.840 27.360 ;
        RECT 173.920 27.040 174.240 27.360 ;
        RECT 174.320 27.040 174.640 27.360 ;
        RECT 174.720 27.040 175.040 27.360 ;
        RECT 175.120 27.040 175.440 27.360 ;
        RECT 175.520 27.040 175.840 27.360 ;
        RECT 175.920 27.040 176.240 27.360 ;
        RECT 176.320 27.040 176.640 27.360 ;
        RECT 176.720 27.040 177.040 27.360 ;
        RECT 177.120 27.040 177.440 27.360 ;
        RECT 177.520 27.040 177.840 27.360 ;
        RECT 177.920 27.040 178.240 27.360 ;
        RECT 178.320 27.040 178.640 27.360 ;
        RECT 178.720 27.040 179.040 27.360 ;
        RECT 179.120 27.040 179.440 27.360 ;
        RECT 179.520 27.040 179.840 27.360 ;
        RECT 179.920 27.040 180.240 27.360 ;
        RECT 180.320 27.040 180.640 27.360 ;
        RECT 25.040 26.640 25.360 26.960 ;
        RECT 25.440 26.640 25.760 26.960 ;
        RECT 25.840 26.640 26.160 26.960 ;
        RECT 26.240 26.640 26.560 26.960 ;
        RECT 26.640 26.640 26.960 26.960 ;
        RECT 27.040 26.640 27.360 26.960 ;
        RECT 27.440 26.640 27.760 26.960 ;
        RECT 27.840 26.640 28.160 26.960 ;
        RECT 28.240 26.640 28.560 26.960 ;
        RECT 28.640 26.640 28.960 26.960 ;
        RECT 29.040 26.640 29.360 26.960 ;
        RECT 29.440 26.640 29.760 26.960 ;
        RECT 29.840 26.640 30.160 26.960 ;
        RECT 30.240 26.640 30.560 26.960 ;
        RECT 30.640 26.640 30.960 26.960 ;
        RECT 31.040 26.640 31.360 26.960 ;
        RECT 31.440 26.640 31.760 26.960 ;
        RECT 31.840 26.640 32.160 26.960 ;
        RECT 32.240 26.640 32.560 26.960 ;
        RECT 32.640 26.640 32.960 26.960 ;
        RECT 33.040 26.640 33.360 26.960 ;
        RECT 33.440 26.640 33.760 26.960 ;
        RECT 33.840 26.640 34.160 26.960 ;
        RECT 34.240 26.640 34.560 26.960 ;
        RECT 34.640 26.640 34.960 26.960 ;
        RECT 35.040 26.640 35.360 26.960 ;
        RECT 35.440 26.640 35.760 26.960 ;
        RECT 35.840 26.640 36.160 26.960 ;
        RECT 36.240 26.640 36.560 26.960 ;
        RECT 36.640 26.640 36.960 26.960 ;
        RECT 37.040 26.640 37.360 26.960 ;
        RECT 37.440 26.640 37.760 26.960 ;
        RECT 37.840 26.640 38.160 26.960 ;
        RECT 38.240 26.640 38.560 26.960 ;
        RECT 38.640 26.640 38.960 26.960 ;
        RECT 39.040 26.640 39.360 26.960 ;
        RECT 39.440 26.640 39.760 26.960 ;
        RECT 39.840 26.640 40.160 26.960 ;
        RECT 40.240 26.640 40.560 26.960 ;
        RECT 40.640 26.640 40.960 26.960 ;
        RECT 41.040 26.640 41.360 26.960 ;
        RECT 41.440 26.640 41.760 26.960 ;
        RECT 41.840 26.640 42.160 26.960 ;
        RECT 42.240 26.640 42.560 26.960 ;
        RECT 42.640 26.640 42.960 26.960 ;
        RECT 43.040 26.640 43.360 26.960 ;
        RECT 43.440 26.640 43.760 26.960 ;
        RECT 43.840 26.640 44.160 26.960 ;
        RECT 44.240 26.640 44.560 26.960 ;
        RECT 44.640 26.640 44.960 26.960 ;
        RECT 70.560 26.640 70.880 26.960 ;
        RECT 70.960 26.640 71.280 26.960 ;
        RECT 71.360 26.640 71.680 26.960 ;
        RECT 71.760 26.640 72.080 26.960 ;
        RECT 120.560 26.640 120.880 26.960 ;
        RECT 120.960 26.640 121.280 26.960 ;
        RECT 121.360 26.640 121.680 26.960 ;
        RECT 121.760 26.640 122.080 26.960 ;
        RECT 160.720 26.640 161.040 26.960 ;
        RECT 161.120 26.640 161.440 26.960 ;
        RECT 161.520 26.640 161.840 26.960 ;
        RECT 161.920 26.640 162.240 26.960 ;
        RECT 162.320 26.640 162.640 26.960 ;
        RECT 162.720 26.640 163.040 26.960 ;
        RECT 163.120 26.640 163.440 26.960 ;
        RECT 163.520 26.640 163.840 26.960 ;
        RECT 163.920 26.640 164.240 26.960 ;
        RECT 164.320 26.640 164.640 26.960 ;
        RECT 164.720 26.640 165.040 26.960 ;
        RECT 165.120 26.640 165.440 26.960 ;
        RECT 165.520 26.640 165.840 26.960 ;
        RECT 165.920 26.640 166.240 26.960 ;
        RECT 166.320 26.640 166.640 26.960 ;
        RECT 166.720 26.640 167.040 26.960 ;
        RECT 167.120 26.640 167.440 26.960 ;
        RECT 167.520 26.640 167.840 26.960 ;
        RECT 167.920 26.640 168.240 26.960 ;
        RECT 168.320 26.640 168.640 26.960 ;
        RECT 168.720 26.640 169.040 26.960 ;
        RECT 169.120 26.640 169.440 26.960 ;
        RECT 169.520 26.640 169.840 26.960 ;
        RECT 169.920 26.640 170.240 26.960 ;
        RECT 170.320 26.640 170.640 26.960 ;
        RECT 170.720 26.640 171.040 26.960 ;
        RECT 171.120 26.640 171.440 26.960 ;
        RECT 171.520 26.640 171.840 26.960 ;
        RECT 171.920 26.640 172.240 26.960 ;
        RECT 172.320 26.640 172.640 26.960 ;
        RECT 172.720 26.640 173.040 26.960 ;
        RECT 173.120 26.640 173.440 26.960 ;
        RECT 173.520 26.640 173.840 26.960 ;
        RECT 173.920 26.640 174.240 26.960 ;
        RECT 174.320 26.640 174.640 26.960 ;
        RECT 174.720 26.640 175.040 26.960 ;
        RECT 175.120 26.640 175.440 26.960 ;
        RECT 175.520 26.640 175.840 26.960 ;
        RECT 175.920 26.640 176.240 26.960 ;
        RECT 176.320 26.640 176.640 26.960 ;
        RECT 176.720 26.640 177.040 26.960 ;
        RECT 177.120 26.640 177.440 26.960 ;
        RECT 177.520 26.640 177.840 26.960 ;
        RECT 177.920 26.640 178.240 26.960 ;
        RECT 178.320 26.640 178.640 26.960 ;
        RECT 178.720 26.640 179.040 26.960 ;
        RECT 179.120 26.640 179.440 26.960 ;
        RECT 179.520 26.640 179.840 26.960 ;
        RECT 179.920 26.640 180.240 26.960 ;
        RECT 180.320 26.640 180.640 26.960 ;
        RECT 25.040 26.240 25.360 26.560 ;
        RECT 25.440 26.240 25.760 26.560 ;
        RECT 25.840 26.240 26.160 26.560 ;
        RECT 26.240 26.240 26.560 26.560 ;
        RECT 26.640 26.240 26.960 26.560 ;
        RECT 27.040 26.240 27.360 26.560 ;
        RECT 27.440 26.240 27.760 26.560 ;
        RECT 27.840 26.240 28.160 26.560 ;
        RECT 28.240 26.240 28.560 26.560 ;
        RECT 28.640 26.240 28.960 26.560 ;
        RECT 29.040 26.240 29.360 26.560 ;
        RECT 29.440 26.240 29.760 26.560 ;
        RECT 29.840 26.240 30.160 26.560 ;
        RECT 30.240 26.240 30.560 26.560 ;
        RECT 30.640 26.240 30.960 26.560 ;
        RECT 31.040 26.240 31.360 26.560 ;
        RECT 31.440 26.240 31.760 26.560 ;
        RECT 31.840 26.240 32.160 26.560 ;
        RECT 32.240 26.240 32.560 26.560 ;
        RECT 32.640 26.240 32.960 26.560 ;
        RECT 33.040 26.240 33.360 26.560 ;
        RECT 33.440 26.240 33.760 26.560 ;
        RECT 33.840 26.240 34.160 26.560 ;
        RECT 34.240 26.240 34.560 26.560 ;
        RECT 34.640 26.240 34.960 26.560 ;
        RECT 35.040 26.240 35.360 26.560 ;
        RECT 35.440 26.240 35.760 26.560 ;
        RECT 35.840 26.240 36.160 26.560 ;
        RECT 36.240 26.240 36.560 26.560 ;
        RECT 36.640 26.240 36.960 26.560 ;
        RECT 37.040 26.240 37.360 26.560 ;
        RECT 37.440 26.240 37.760 26.560 ;
        RECT 37.840 26.240 38.160 26.560 ;
        RECT 38.240 26.240 38.560 26.560 ;
        RECT 38.640 26.240 38.960 26.560 ;
        RECT 39.040 26.240 39.360 26.560 ;
        RECT 39.440 26.240 39.760 26.560 ;
        RECT 39.840 26.240 40.160 26.560 ;
        RECT 40.240 26.240 40.560 26.560 ;
        RECT 40.640 26.240 40.960 26.560 ;
        RECT 41.040 26.240 41.360 26.560 ;
        RECT 41.440 26.240 41.760 26.560 ;
        RECT 41.840 26.240 42.160 26.560 ;
        RECT 42.240 26.240 42.560 26.560 ;
        RECT 42.640 26.240 42.960 26.560 ;
        RECT 43.040 26.240 43.360 26.560 ;
        RECT 43.440 26.240 43.760 26.560 ;
        RECT 43.840 26.240 44.160 26.560 ;
        RECT 44.240 26.240 44.560 26.560 ;
        RECT 44.640 26.240 44.960 26.560 ;
        RECT 70.560 26.240 70.880 26.560 ;
        RECT 70.960 26.240 71.280 26.560 ;
        RECT 71.360 26.240 71.680 26.560 ;
        RECT 71.760 26.240 72.080 26.560 ;
        RECT 120.560 26.240 120.880 26.560 ;
        RECT 120.960 26.240 121.280 26.560 ;
        RECT 121.360 26.240 121.680 26.560 ;
        RECT 121.760 26.240 122.080 26.560 ;
        RECT 160.720 26.240 161.040 26.560 ;
        RECT 161.120 26.240 161.440 26.560 ;
        RECT 161.520 26.240 161.840 26.560 ;
        RECT 161.920 26.240 162.240 26.560 ;
        RECT 162.320 26.240 162.640 26.560 ;
        RECT 162.720 26.240 163.040 26.560 ;
        RECT 163.120 26.240 163.440 26.560 ;
        RECT 163.520 26.240 163.840 26.560 ;
        RECT 163.920 26.240 164.240 26.560 ;
        RECT 164.320 26.240 164.640 26.560 ;
        RECT 164.720 26.240 165.040 26.560 ;
        RECT 165.120 26.240 165.440 26.560 ;
        RECT 165.520 26.240 165.840 26.560 ;
        RECT 165.920 26.240 166.240 26.560 ;
        RECT 166.320 26.240 166.640 26.560 ;
        RECT 166.720 26.240 167.040 26.560 ;
        RECT 167.120 26.240 167.440 26.560 ;
        RECT 167.520 26.240 167.840 26.560 ;
        RECT 167.920 26.240 168.240 26.560 ;
        RECT 168.320 26.240 168.640 26.560 ;
        RECT 168.720 26.240 169.040 26.560 ;
        RECT 169.120 26.240 169.440 26.560 ;
        RECT 169.520 26.240 169.840 26.560 ;
        RECT 169.920 26.240 170.240 26.560 ;
        RECT 170.320 26.240 170.640 26.560 ;
        RECT 170.720 26.240 171.040 26.560 ;
        RECT 171.120 26.240 171.440 26.560 ;
        RECT 171.520 26.240 171.840 26.560 ;
        RECT 171.920 26.240 172.240 26.560 ;
        RECT 172.320 26.240 172.640 26.560 ;
        RECT 172.720 26.240 173.040 26.560 ;
        RECT 173.120 26.240 173.440 26.560 ;
        RECT 173.520 26.240 173.840 26.560 ;
        RECT 173.920 26.240 174.240 26.560 ;
        RECT 174.320 26.240 174.640 26.560 ;
        RECT 174.720 26.240 175.040 26.560 ;
        RECT 175.120 26.240 175.440 26.560 ;
        RECT 175.520 26.240 175.840 26.560 ;
        RECT 175.920 26.240 176.240 26.560 ;
        RECT 176.320 26.240 176.640 26.560 ;
        RECT 176.720 26.240 177.040 26.560 ;
        RECT 177.120 26.240 177.440 26.560 ;
        RECT 177.520 26.240 177.840 26.560 ;
        RECT 177.920 26.240 178.240 26.560 ;
        RECT 178.320 26.240 178.640 26.560 ;
        RECT 178.720 26.240 179.040 26.560 ;
        RECT 179.120 26.240 179.440 26.560 ;
        RECT 179.520 26.240 179.840 26.560 ;
        RECT 179.920 26.240 180.240 26.560 ;
        RECT 180.320 26.240 180.640 26.560 ;
        RECT 25.040 25.840 25.360 26.160 ;
        RECT 25.440 25.840 25.760 26.160 ;
        RECT 25.840 25.840 26.160 26.160 ;
        RECT 26.240 25.840 26.560 26.160 ;
        RECT 26.640 25.840 26.960 26.160 ;
        RECT 27.040 25.840 27.360 26.160 ;
        RECT 27.440 25.840 27.760 26.160 ;
        RECT 27.840 25.840 28.160 26.160 ;
        RECT 28.240 25.840 28.560 26.160 ;
        RECT 28.640 25.840 28.960 26.160 ;
        RECT 29.040 25.840 29.360 26.160 ;
        RECT 29.440 25.840 29.760 26.160 ;
        RECT 29.840 25.840 30.160 26.160 ;
        RECT 30.240 25.840 30.560 26.160 ;
        RECT 30.640 25.840 30.960 26.160 ;
        RECT 31.040 25.840 31.360 26.160 ;
        RECT 31.440 25.840 31.760 26.160 ;
        RECT 31.840 25.840 32.160 26.160 ;
        RECT 32.240 25.840 32.560 26.160 ;
        RECT 32.640 25.840 32.960 26.160 ;
        RECT 33.040 25.840 33.360 26.160 ;
        RECT 33.440 25.840 33.760 26.160 ;
        RECT 33.840 25.840 34.160 26.160 ;
        RECT 34.240 25.840 34.560 26.160 ;
        RECT 34.640 25.840 34.960 26.160 ;
        RECT 35.040 25.840 35.360 26.160 ;
        RECT 35.440 25.840 35.760 26.160 ;
        RECT 35.840 25.840 36.160 26.160 ;
        RECT 36.240 25.840 36.560 26.160 ;
        RECT 36.640 25.840 36.960 26.160 ;
        RECT 37.040 25.840 37.360 26.160 ;
        RECT 37.440 25.840 37.760 26.160 ;
        RECT 37.840 25.840 38.160 26.160 ;
        RECT 38.240 25.840 38.560 26.160 ;
        RECT 38.640 25.840 38.960 26.160 ;
        RECT 39.040 25.840 39.360 26.160 ;
        RECT 39.440 25.840 39.760 26.160 ;
        RECT 39.840 25.840 40.160 26.160 ;
        RECT 40.240 25.840 40.560 26.160 ;
        RECT 40.640 25.840 40.960 26.160 ;
        RECT 41.040 25.840 41.360 26.160 ;
        RECT 41.440 25.840 41.760 26.160 ;
        RECT 41.840 25.840 42.160 26.160 ;
        RECT 42.240 25.840 42.560 26.160 ;
        RECT 42.640 25.840 42.960 26.160 ;
        RECT 43.040 25.840 43.360 26.160 ;
        RECT 43.440 25.840 43.760 26.160 ;
        RECT 43.840 25.840 44.160 26.160 ;
        RECT 44.240 25.840 44.560 26.160 ;
        RECT 44.640 25.840 44.960 26.160 ;
        RECT 70.560 25.840 70.880 26.160 ;
        RECT 70.960 25.840 71.280 26.160 ;
        RECT 71.360 25.840 71.680 26.160 ;
        RECT 71.760 25.840 72.080 26.160 ;
        RECT 120.560 25.840 120.880 26.160 ;
        RECT 120.960 25.840 121.280 26.160 ;
        RECT 121.360 25.840 121.680 26.160 ;
        RECT 121.760 25.840 122.080 26.160 ;
        RECT 160.720 25.840 161.040 26.160 ;
        RECT 161.120 25.840 161.440 26.160 ;
        RECT 161.520 25.840 161.840 26.160 ;
        RECT 161.920 25.840 162.240 26.160 ;
        RECT 162.320 25.840 162.640 26.160 ;
        RECT 162.720 25.840 163.040 26.160 ;
        RECT 163.120 25.840 163.440 26.160 ;
        RECT 163.520 25.840 163.840 26.160 ;
        RECT 163.920 25.840 164.240 26.160 ;
        RECT 164.320 25.840 164.640 26.160 ;
        RECT 164.720 25.840 165.040 26.160 ;
        RECT 165.120 25.840 165.440 26.160 ;
        RECT 165.520 25.840 165.840 26.160 ;
        RECT 165.920 25.840 166.240 26.160 ;
        RECT 166.320 25.840 166.640 26.160 ;
        RECT 166.720 25.840 167.040 26.160 ;
        RECT 167.120 25.840 167.440 26.160 ;
        RECT 167.520 25.840 167.840 26.160 ;
        RECT 167.920 25.840 168.240 26.160 ;
        RECT 168.320 25.840 168.640 26.160 ;
        RECT 168.720 25.840 169.040 26.160 ;
        RECT 169.120 25.840 169.440 26.160 ;
        RECT 169.520 25.840 169.840 26.160 ;
        RECT 169.920 25.840 170.240 26.160 ;
        RECT 170.320 25.840 170.640 26.160 ;
        RECT 170.720 25.840 171.040 26.160 ;
        RECT 171.120 25.840 171.440 26.160 ;
        RECT 171.520 25.840 171.840 26.160 ;
        RECT 171.920 25.840 172.240 26.160 ;
        RECT 172.320 25.840 172.640 26.160 ;
        RECT 172.720 25.840 173.040 26.160 ;
        RECT 173.120 25.840 173.440 26.160 ;
        RECT 173.520 25.840 173.840 26.160 ;
        RECT 173.920 25.840 174.240 26.160 ;
        RECT 174.320 25.840 174.640 26.160 ;
        RECT 174.720 25.840 175.040 26.160 ;
        RECT 175.120 25.840 175.440 26.160 ;
        RECT 175.520 25.840 175.840 26.160 ;
        RECT 175.920 25.840 176.240 26.160 ;
        RECT 176.320 25.840 176.640 26.160 ;
        RECT 176.720 25.840 177.040 26.160 ;
        RECT 177.120 25.840 177.440 26.160 ;
        RECT 177.520 25.840 177.840 26.160 ;
        RECT 177.920 25.840 178.240 26.160 ;
        RECT 178.320 25.840 178.640 26.160 ;
        RECT 178.720 25.840 179.040 26.160 ;
        RECT 179.120 25.840 179.440 26.160 ;
        RECT 179.520 25.840 179.840 26.160 ;
        RECT 179.920 25.840 180.240 26.160 ;
        RECT 180.320 25.840 180.640 26.160 ;
        RECT 25.040 25.440 25.360 25.760 ;
        RECT 25.440 25.440 25.760 25.760 ;
        RECT 25.840 25.440 26.160 25.760 ;
        RECT 26.240 25.440 26.560 25.760 ;
        RECT 26.640 25.440 26.960 25.760 ;
        RECT 27.040 25.440 27.360 25.760 ;
        RECT 27.440 25.440 27.760 25.760 ;
        RECT 27.840 25.440 28.160 25.760 ;
        RECT 28.240 25.440 28.560 25.760 ;
        RECT 28.640 25.440 28.960 25.760 ;
        RECT 29.040 25.440 29.360 25.760 ;
        RECT 29.440 25.440 29.760 25.760 ;
        RECT 29.840 25.440 30.160 25.760 ;
        RECT 30.240 25.440 30.560 25.760 ;
        RECT 30.640 25.440 30.960 25.760 ;
        RECT 31.040 25.440 31.360 25.760 ;
        RECT 31.440 25.440 31.760 25.760 ;
        RECT 31.840 25.440 32.160 25.760 ;
        RECT 32.240 25.440 32.560 25.760 ;
        RECT 32.640 25.440 32.960 25.760 ;
        RECT 33.040 25.440 33.360 25.760 ;
        RECT 33.440 25.440 33.760 25.760 ;
        RECT 33.840 25.440 34.160 25.760 ;
        RECT 34.240 25.440 34.560 25.760 ;
        RECT 34.640 25.440 34.960 25.760 ;
        RECT 35.040 25.440 35.360 25.760 ;
        RECT 35.440 25.440 35.760 25.760 ;
        RECT 35.840 25.440 36.160 25.760 ;
        RECT 36.240 25.440 36.560 25.760 ;
        RECT 36.640 25.440 36.960 25.760 ;
        RECT 37.040 25.440 37.360 25.760 ;
        RECT 37.440 25.440 37.760 25.760 ;
        RECT 37.840 25.440 38.160 25.760 ;
        RECT 38.240 25.440 38.560 25.760 ;
        RECT 38.640 25.440 38.960 25.760 ;
        RECT 39.040 25.440 39.360 25.760 ;
        RECT 39.440 25.440 39.760 25.760 ;
        RECT 39.840 25.440 40.160 25.760 ;
        RECT 40.240 25.440 40.560 25.760 ;
        RECT 40.640 25.440 40.960 25.760 ;
        RECT 41.040 25.440 41.360 25.760 ;
        RECT 41.440 25.440 41.760 25.760 ;
        RECT 41.840 25.440 42.160 25.760 ;
        RECT 42.240 25.440 42.560 25.760 ;
        RECT 42.640 25.440 42.960 25.760 ;
        RECT 43.040 25.440 43.360 25.760 ;
        RECT 43.440 25.440 43.760 25.760 ;
        RECT 43.840 25.440 44.160 25.760 ;
        RECT 44.240 25.440 44.560 25.760 ;
        RECT 44.640 25.440 44.960 25.760 ;
        RECT 70.560 25.440 70.880 25.760 ;
        RECT 70.960 25.440 71.280 25.760 ;
        RECT 71.360 25.440 71.680 25.760 ;
        RECT 71.760 25.440 72.080 25.760 ;
        RECT 120.560 25.440 120.880 25.760 ;
        RECT 120.960 25.440 121.280 25.760 ;
        RECT 121.360 25.440 121.680 25.760 ;
        RECT 121.760 25.440 122.080 25.760 ;
        RECT 160.720 25.440 161.040 25.760 ;
        RECT 161.120 25.440 161.440 25.760 ;
        RECT 161.520 25.440 161.840 25.760 ;
        RECT 161.920 25.440 162.240 25.760 ;
        RECT 162.320 25.440 162.640 25.760 ;
        RECT 162.720 25.440 163.040 25.760 ;
        RECT 163.120 25.440 163.440 25.760 ;
        RECT 163.520 25.440 163.840 25.760 ;
        RECT 163.920 25.440 164.240 25.760 ;
        RECT 164.320 25.440 164.640 25.760 ;
        RECT 164.720 25.440 165.040 25.760 ;
        RECT 165.120 25.440 165.440 25.760 ;
        RECT 165.520 25.440 165.840 25.760 ;
        RECT 165.920 25.440 166.240 25.760 ;
        RECT 166.320 25.440 166.640 25.760 ;
        RECT 166.720 25.440 167.040 25.760 ;
        RECT 167.120 25.440 167.440 25.760 ;
        RECT 167.520 25.440 167.840 25.760 ;
        RECT 167.920 25.440 168.240 25.760 ;
        RECT 168.320 25.440 168.640 25.760 ;
        RECT 168.720 25.440 169.040 25.760 ;
        RECT 169.120 25.440 169.440 25.760 ;
        RECT 169.520 25.440 169.840 25.760 ;
        RECT 169.920 25.440 170.240 25.760 ;
        RECT 170.320 25.440 170.640 25.760 ;
        RECT 170.720 25.440 171.040 25.760 ;
        RECT 171.120 25.440 171.440 25.760 ;
        RECT 171.520 25.440 171.840 25.760 ;
        RECT 171.920 25.440 172.240 25.760 ;
        RECT 172.320 25.440 172.640 25.760 ;
        RECT 172.720 25.440 173.040 25.760 ;
        RECT 173.120 25.440 173.440 25.760 ;
        RECT 173.520 25.440 173.840 25.760 ;
        RECT 173.920 25.440 174.240 25.760 ;
        RECT 174.320 25.440 174.640 25.760 ;
        RECT 174.720 25.440 175.040 25.760 ;
        RECT 175.120 25.440 175.440 25.760 ;
        RECT 175.520 25.440 175.840 25.760 ;
        RECT 175.920 25.440 176.240 25.760 ;
        RECT 176.320 25.440 176.640 25.760 ;
        RECT 176.720 25.440 177.040 25.760 ;
        RECT 177.120 25.440 177.440 25.760 ;
        RECT 177.520 25.440 177.840 25.760 ;
        RECT 177.920 25.440 178.240 25.760 ;
        RECT 178.320 25.440 178.640 25.760 ;
        RECT 178.720 25.440 179.040 25.760 ;
        RECT 179.120 25.440 179.440 25.760 ;
        RECT 179.520 25.440 179.840 25.760 ;
        RECT 179.920 25.440 180.240 25.760 ;
        RECT 180.320 25.440 180.640 25.760 ;
        RECT 25.040 25.040 25.360 25.360 ;
        RECT 25.440 25.040 25.760 25.360 ;
        RECT 25.840 25.040 26.160 25.360 ;
        RECT 26.240 25.040 26.560 25.360 ;
        RECT 26.640 25.040 26.960 25.360 ;
        RECT 27.040 25.040 27.360 25.360 ;
        RECT 27.440 25.040 27.760 25.360 ;
        RECT 27.840 25.040 28.160 25.360 ;
        RECT 28.240 25.040 28.560 25.360 ;
        RECT 28.640 25.040 28.960 25.360 ;
        RECT 29.040 25.040 29.360 25.360 ;
        RECT 29.440 25.040 29.760 25.360 ;
        RECT 29.840 25.040 30.160 25.360 ;
        RECT 30.240 25.040 30.560 25.360 ;
        RECT 30.640 25.040 30.960 25.360 ;
        RECT 31.040 25.040 31.360 25.360 ;
        RECT 31.440 25.040 31.760 25.360 ;
        RECT 31.840 25.040 32.160 25.360 ;
        RECT 32.240 25.040 32.560 25.360 ;
        RECT 32.640 25.040 32.960 25.360 ;
        RECT 33.040 25.040 33.360 25.360 ;
        RECT 33.440 25.040 33.760 25.360 ;
        RECT 33.840 25.040 34.160 25.360 ;
        RECT 34.240 25.040 34.560 25.360 ;
        RECT 34.640 25.040 34.960 25.360 ;
        RECT 35.040 25.040 35.360 25.360 ;
        RECT 35.440 25.040 35.760 25.360 ;
        RECT 35.840 25.040 36.160 25.360 ;
        RECT 36.240 25.040 36.560 25.360 ;
        RECT 36.640 25.040 36.960 25.360 ;
        RECT 37.040 25.040 37.360 25.360 ;
        RECT 37.440 25.040 37.760 25.360 ;
        RECT 37.840 25.040 38.160 25.360 ;
        RECT 38.240 25.040 38.560 25.360 ;
        RECT 38.640 25.040 38.960 25.360 ;
        RECT 39.040 25.040 39.360 25.360 ;
        RECT 39.440 25.040 39.760 25.360 ;
        RECT 39.840 25.040 40.160 25.360 ;
        RECT 40.240 25.040 40.560 25.360 ;
        RECT 40.640 25.040 40.960 25.360 ;
        RECT 41.040 25.040 41.360 25.360 ;
        RECT 41.440 25.040 41.760 25.360 ;
        RECT 41.840 25.040 42.160 25.360 ;
        RECT 42.240 25.040 42.560 25.360 ;
        RECT 42.640 25.040 42.960 25.360 ;
        RECT 43.040 25.040 43.360 25.360 ;
        RECT 43.440 25.040 43.760 25.360 ;
        RECT 43.840 25.040 44.160 25.360 ;
        RECT 44.240 25.040 44.560 25.360 ;
        RECT 44.640 25.040 44.960 25.360 ;
        RECT 70.560 25.040 70.880 25.360 ;
        RECT 70.960 25.040 71.280 25.360 ;
        RECT 71.360 25.040 71.680 25.360 ;
        RECT 71.760 25.040 72.080 25.360 ;
        RECT 120.560 25.040 120.880 25.360 ;
        RECT 120.960 25.040 121.280 25.360 ;
        RECT 121.360 25.040 121.680 25.360 ;
        RECT 121.760 25.040 122.080 25.360 ;
        RECT 160.720 25.040 161.040 25.360 ;
        RECT 161.120 25.040 161.440 25.360 ;
        RECT 161.520 25.040 161.840 25.360 ;
        RECT 161.920 25.040 162.240 25.360 ;
        RECT 162.320 25.040 162.640 25.360 ;
        RECT 162.720 25.040 163.040 25.360 ;
        RECT 163.120 25.040 163.440 25.360 ;
        RECT 163.520 25.040 163.840 25.360 ;
        RECT 163.920 25.040 164.240 25.360 ;
        RECT 164.320 25.040 164.640 25.360 ;
        RECT 164.720 25.040 165.040 25.360 ;
        RECT 165.120 25.040 165.440 25.360 ;
        RECT 165.520 25.040 165.840 25.360 ;
        RECT 165.920 25.040 166.240 25.360 ;
        RECT 166.320 25.040 166.640 25.360 ;
        RECT 166.720 25.040 167.040 25.360 ;
        RECT 167.120 25.040 167.440 25.360 ;
        RECT 167.520 25.040 167.840 25.360 ;
        RECT 167.920 25.040 168.240 25.360 ;
        RECT 168.320 25.040 168.640 25.360 ;
        RECT 168.720 25.040 169.040 25.360 ;
        RECT 169.120 25.040 169.440 25.360 ;
        RECT 169.520 25.040 169.840 25.360 ;
        RECT 169.920 25.040 170.240 25.360 ;
        RECT 170.320 25.040 170.640 25.360 ;
        RECT 170.720 25.040 171.040 25.360 ;
        RECT 171.120 25.040 171.440 25.360 ;
        RECT 171.520 25.040 171.840 25.360 ;
        RECT 171.920 25.040 172.240 25.360 ;
        RECT 172.320 25.040 172.640 25.360 ;
        RECT 172.720 25.040 173.040 25.360 ;
        RECT 173.120 25.040 173.440 25.360 ;
        RECT 173.520 25.040 173.840 25.360 ;
        RECT 173.920 25.040 174.240 25.360 ;
        RECT 174.320 25.040 174.640 25.360 ;
        RECT 174.720 25.040 175.040 25.360 ;
        RECT 175.120 25.040 175.440 25.360 ;
        RECT 175.520 25.040 175.840 25.360 ;
        RECT 175.920 25.040 176.240 25.360 ;
        RECT 176.320 25.040 176.640 25.360 ;
        RECT 176.720 25.040 177.040 25.360 ;
        RECT 177.120 25.040 177.440 25.360 ;
        RECT 177.520 25.040 177.840 25.360 ;
        RECT 177.920 25.040 178.240 25.360 ;
        RECT 178.320 25.040 178.640 25.360 ;
        RECT 178.720 25.040 179.040 25.360 ;
        RECT 179.120 25.040 179.440 25.360 ;
        RECT 179.520 25.040 179.840 25.360 ;
        RECT 179.920 25.040 180.240 25.360 ;
        RECT 180.320 25.040 180.640 25.360 ;
      LAYER met4 ;
        RECT 25.000 25.000 45.000 180.200 ;
        RECT 70.520 151.200 72.120 205.200 ;
        RECT 120.520 151.200 122.120 205.200 ;
        RECT 70.520 0.000 72.120 54.000 ;
        RECT 120.520 0.000 122.120 54.000 ;
        RECT 160.680 25.000 180.680 180.200 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.200 205.680 205.200 ;
        RECT 0.000 0.000 205.680 20.000 ;
      LAYER via3 ;
        RECT 0.040 204.840 0.360 205.160 ;
        RECT 0.440 204.840 0.760 205.160 ;
        RECT 0.840 204.840 1.160 205.160 ;
        RECT 1.240 204.840 1.560 205.160 ;
        RECT 1.640 204.840 1.960 205.160 ;
        RECT 2.040 204.840 2.360 205.160 ;
        RECT 2.440 204.840 2.760 205.160 ;
        RECT 2.840 204.840 3.160 205.160 ;
        RECT 3.240 204.840 3.560 205.160 ;
        RECT 3.640 204.840 3.960 205.160 ;
        RECT 4.040 204.840 4.360 205.160 ;
        RECT 4.440 204.840 4.760 205.160 ;
        RECT 4.840 204.840 5.160 205.160 ;
        RECT 5.240 204.840 5.560 205.160 ;
        RECT 5.640 204.840 5.960 205.160 ;
        RECT 6.040 204.840 6.360 205.160 ;
        RECT 6.440 204.840 6.760 205.160 ;
        RECT 6.840 204.840 7.160 205.160 ;
        RECT 7.240 204.840 7.560 205.160 ;
        RECT 7.640 204.840 7.960 205.160 ;
        RECT 8.040 204.840 8.360 205.160 ;
        RECT 8.440 204.840 8.760 205.160 ;
        RECT 8.840 204.840 9.160 205.160 ;
        RECT 9.240 204.840 9.560 205.160 ;
        RECT 9.640 204.840 9.960 205.160 ;
        RECT 10.040 204.840 10.360 205.160 ;
        RECT 10.440 204.840 10.760 205.160 ;
        RECT 10.840 204.840 11.160 205.160 ;
        RECT 11.240 204.840 11.560 205.160 ;
        RECT 11.640 204.840 11.960 205.160 ;
        RECT 12.040 204.840 12.360 205.160 ;
        RECT 12.440 204.840 12.760 205.160 ;
        RECT 12.840 204.840 13.160 205.160 ;
        RECT 13.240 204.840 13.560 205.160 ;
        RECT 13.640 204.840 13.960 205.160 ;
        RECT 14.040 204.840 14.360 205.160 ;
        RECT 14.440 204.840 14.760 205.160 ;
        RECT 14.840 204.840 15.160 205.160 ;
        RECT 15.240 204.840 15.560 205.160 ;
        RECT 15.640 204.840 15.960 205.160 ;
        RECT 16.040 204.840 16.360 205.160 ;
        RECT 16.440 204.840 16.760 205.160 ;
        RECT 16.840 204.840 17.160 205.160 ;
        RECT 17.240 204.840 17.560 205.160 ;
        RECT 17.640 204.840 17.960 205.160 ;
        RECT 18.040 204.840 18.360 205.160 ;
        RECT 18.440 204.840 18.760 205.160 ;
        RECT 18.840 204.840 19.160 205.160 ;
        RECT 19.240 204.840 19.560 205.160 ;
        RECT 19.640 204.840 19.960 205.160 ;
        RECT 95.560 204.840 95.880 205.160 ;
        RECT 95.960 204.840 96.280 205.160 ;
        RECT 96.360 204.840 96.680 205.160 ;
        RECT 96.760 204.840 97.080 205.160 ;
        RECT 145.560 204.840 145.880 205.160 ;
        RECT 145.960 204.840 146.280 205.160 ;
        RECT 146.360 204.840 146.680 205.160 ;
        RECT 146.760 204.840 147.080 205.160 ;
        RECT 185.720 204.840 186.040 205.160 ;
        RECT 186.120 204.840 186.440 205.160 ;
        RECT 186.520 204.840 186.840 205.160 ;
        RECT 186.920 204.840 187.240 205.160 ;
        RECT 187.320 204.840 187.640 205.160 ;
        RECT 187.720 204.840 188.040 205.160 ;
        RECT 188.120 204.840 188.440 205.160 ;
        RECT 188.520 204.840 188.840 205.160 ;
        RECT 188.920 204.840 189.240 205.160 ;
        RECT 189.320 204.840 189.640 205.160 ;
        RECT 189.720 204.840 190.040 205.160 ;
        RECT 190.120 204.840 190.440 205.160 ;
        RECT 190.520 204.840 190.840 205.160 ;
        RECT 190.920 204.840 191.240 205.160 ;
        RECT 191.320 204.840 191.640 205.160 ;
        RECT 191.720 204.840 192.040 205.160 ;
        RECT 192.120 204.840 192.440 205.160 ;
        RECT 192.520 204.840 192.840 205.160 ;
        RECT 192.920 204.840 193.240 205.160 ;
        RECT 193.320 204.840 193.640 205.160 ;
        RECT 193.720 204.840 194.040 205.160 ;
        RECT 194.120 204.840 194.440 205.160 ;
        RECT 194.520 204.840 194.840 205.160 ;
        RECT 194.920 204.840 195.240 205.160 ;
        RECT 195.320 204.840 195.640 205.160 ;
        RECT 195.720 204.840 196.040 205.160 ;
        RECT 196.120 204.840 196.440 205.160 ;
        RECT 196.520 204.840 196.840 205.160 ;
        RECT 196.920 204.840 197.240 205.160 ;
        RECT 197.320 204.840 197.640 205.160 ;
        RECT 197.720 204.840 198.040 205.160 ;
        RECT 198.120 204.840 198.440 205.160 ;
        RECT 198.520 204.840 198.840 205.160 ;
        RECT 198.920 204.840 199.240 205.160 ;
        RECT 199.320 204.840 199.640 205.160 ;
        RECT 199.720 204.840 200.040 205.160 ;
        RECT 200.120 204.840 200.440 205.160 ;
        RECT 200.520 204.840 200.840 205.160 ;
        RECT 200.920 204.840 201.240 205.160 ;
        RECT 201.320 204.840 201.640 205.160 ;
        RECT 201.720 204.840 202.040 205.160 ;
        RECT 202.120 204.840 202.440 205.160 ;
        RECT 202.520 204.840 202.840 205.160 ;
        RECT 202.920 204.840 203.240 205.160 ;
        RECT 203.320 204.840 203.640 205.160 ;
        RECT 203.720 204.840 204.040 205.160 ;
        RECT 204.120 204.840 204.440 205.160 ;
        RECT 204.520 204.840 204.840 205.160 ;
        RECT 204.920 204.840 205.240 205.160 ;
        RECT 205.320 204.840 205.640 205.160 ;
        RECT 0.040 204.440 0.360 204.760 ;
        RECT 0.440 204.440 0.760 204.760 ;
        RECT 0.840 204.440 1.160 204.760 ;
        RECT 1.240 204.440 1.560 204.760 ;
        RECT 1.640 204.440 1.960 204.760 ;
        RECT 2.040 204.440 2.360 204.760 ;
        RECT 2.440 204.440 2.760 204.760 ;
        RECT 2.840 204.440 3.160 204.760 ;
        RECT 3.240 204.440 3.560 204.760 ;
        RECT 3.640 204.440 3.960 204.760 ;
        RECT 4.040 204.440 4.360 204.760 ;
        RECT 4.440 204.440 4.760 204.760 ;
        RECT 4.840 204.440 5.160 204.760 ;
        RECT 5.240 204.440 5.560 204.760 ;
        RECT 5.640 204.440 5.960 204.760 ;
        RECT 6.040 204.440 6.360 204.760 ;
        RECT 6.440 204.440 6.760 204.760 ;
        RECT 6.840 204.440 7.160 204.760 ;
        RECT 7.240 204.440 7.560 204.760 ;
        RECT 7.640 204.440 7.960 204.760 ;
        RECT 8.040 204.440 8.360 204.760 ;
        RECT 8.440 204.440 8.760 204.760 ;
        RECT 8.840 204.440 9.160 204.760 ;
        RECT 9.240 204.440 9.560 204.760 ;
        RECT 9.640 204.440 9.960 204.760 ;
        RECT 10.040 204.440 10.360 204.760 ;
        RECT 10.440 204.440 10.760 204.760 ;
        RECT 10.840 204.440 11.160 204.760 ;
        RECT 11.240 204.440 11.560 204.760 ;
        RECT 11.640 204.440 11.960 204.760 ;
        RECT 12.040 204.440 12.360 204.760 ;
        RECT 12.440 204.440 12.760 204.760 ;
        RECT 12.840 204.440 13.160 204.760 ;
        RECT 13.240 204.440 13.560 204.760 ;
        RECT 13.640 204.440 13.960 204.760 ;
        RECT 14.040 204.440 14.360 204.760 ;
        RECT 14.440 204.440 14.760 204.760 ;
        RECT 14.840 204.440 15.160 204.760 ;
        RECT 15.240 204.440 15.560 204.760 ;
        RECT 15.640 204.440 15.960 204.760 ;
        RECT 16.040 204.440 16.360 204.760 ;
        RECT 16.440 204.440 16.760 204.760 ;
        RECT 16.840 204.440 17.160 204.760 ;
        RECT 17.240 204.440 17.560 204.760 ;
        RECT 17.640 204.440 17.960 204.760 ;
        RECT 18.040 204.440 18.360 204.760 ;
        RECT 18.440 204.440 18.760 204.760 ;
        RECT 18.840 204.440 19.160 204.760 ;
        RECT 19.240 204.440 19.560 204.760 ;
        RECT 19.640 204.440 19.960 204.760 ;
        RECT 95.560 204.440 95.880 204.760 ;
        RECT 95.960 204.440 96.280 204.760 ;
        RECT 96.360 204.440 96.680 204.760 ;
        RECT 96.760 204.440 97.080 204.760 ;
        RECT 145.560 204.440 145.880 204.760 ;
        RECT 145.960 204.440 146.280 204.760 ;
        RECT 146.360 204.440 146.680 204.760 ;
        RECT 146.760 204.440 147.080 204.760 ;
        RECT 185.720 204.440 186.040 204.760 ;
        RECT 186.120 204.440 186.440 204.760 ;
        RECT 186.520 204.440 186.840 204.760 ;
        RECT 186.920 204.440 187.240 204.760 ;
        RECT 187.320 204.440 187.640 204.760 ;
        RECT 187.720 204.440 188.040 204.760 ;
        RECT 188.120 204.440 188.440 204.760 ;
        RECT 188.520 204.440 188.840 204.760 ;
        RECT 188.920 204.440 189.240 204.760 ;
        RECT 189.320 204.440 189.640 204.760 ;
        RECT 189.720 204.440 190.040 204.760 ;
        RECT 190.120 204.440 190.440 204.760 ;
        RECT 190.520 204.440 190.840 204.760 ;
        RECT 190.920 204.440 191.240 204.760 ;
        RECT 191.320 204.440 191.640 204.760 ;
        RECT 191.720 204.440 192.040 204.760 ;
        RECT 192.120 204.440 192.440 204.760 ;
        RECT 192.520 204.440 192.840 204.760 ;
        RECT 192.920 204.440 193.240 204.760 ;
        RECT 193.320 204.440 193.640 204.760 ;
        RECT 193.720 204.440 194.040 204.760 ;
        RECT 194.120 204.440 194.440 204.760 ;
        RECT 194.520 204.440 194.840 204.760 ;
        RECT 194.920 204.440 195.240 204.760 ;
        RECT 195.320 204.440 195.640 204.760 ;
        RECT 195.720 204.440 196.040 204.760 ;
        RECT 196.120 204.440 196.440 204.760 ;
        RECT 196.520 204.440 196.840 204.760 ;
        RECT 196.920 204.440 197.240 204.760 ;
        RECT 197.320 204.440 197.640 204.760 ;
        RECT 197.720 204.440 198.040 204.760 ;
        RECT 198.120 204.440 198.440 204.760 ;
        RECT 198.520 204.440 198.840 204.760 ;
        RECT 198.920 204.440 199.240 204.760 ;
        RECT 199.320 204.440 199.640 204.760 ;
        RECT 199.720 204.440 200.040 204.760 ;
        RECT 200.120 204.440 200.440 204.760 ;
        RECT 200.520 204.440 200.840 204.760 ;
        RECT 200.920 204.440 201.240 204.760 ;
        RECT 201.320 204.440 201.640 204.760 ;
        RECT 201.720 204.440 202.040 204.760 ;
        RECT 202.120 204.440 202.440 204.760 ;
        RECT 202.520 204.440 202.840 204.760 ;
        RECT 202.920 204.440 203.240 204.760 ;
        RECT 203.320 204.440 203.640 204.760 ;
        RECT 203.720 204.440 204.040 204.760 ;
        RECT 204.120 204.440 204.440 204.760 ;
        RECT 204.520 204.440 204.840 204.760 ;
        RECT 204.920 204.440 205.240 204.760 ;
        RECT 205.320 204.440 205.640 204.760 ;
        RECT 0.040 204.040 0.360 204.360 ;
        RECT 0.440 204.040 0.760 204.360 ;
        RECT 0.840 204.040 1.160 204.360 ;
        RECT 1.240 204.040 1.560 204.360 ;
        RECT 1.640 204.040 1.960 204.360 ;
        RECT 2.040 204.040 2.360 204.360 ;
        RECT 2.440 204.040 2.760 204.360 ;
        RECT 2.840 204.040 3.160 204.360 ;
        RECT 3.240 204.040 3.560 204.360 ;
        RECT 3.640 204.040 3.960 204.360 ;
        RECT 4.040 204.040 4.360 204.360 ;
        RECT 4.440 204.040 4.760 204.360 ;
        RECT 4.840 204.040 5.160 204.360 ;
        RECT 5.240 204.040 5.560 204.360 ;
        RECT 5.640 204.040 5.960 204.360 ;
        RECT 6.040 204.040 6.360 204.360 ;
        RECT 6.440 204.040 6.760 204.360 ;
        RECT 6.840 204.040 7.160 204.360 ;
        RECT 7.240 204.040 7.560 204.360 ;
        RECT 7.640 204.040 7.960 204.360 ;
        RECT 8.040 204.040 8.360 204.360 ;
        RECT 8.440 204.040 8.760 204.360 ;
        RECT 8.840 204.040 9.160 204.360 ;
        RECT 9.240 204.040 9.560 204.360 ;
        RECT 9.640 204.040 9.960 204.360 ;
        RECT 10.040 204.040 10.360 204.360 ;
        RECT 10.440 204.040 10.760 204.360 ;
        RECT 10.840 204.040 11.160 204.360 ;
        RECT 11.240 204.040 11.560 204.360 ;
        RECT 11.640 204.040 11.960 204.360 ;
        RECT 12.040 204.040 12.360 204.360 ;
        RECT 12.440 204.040 12.760 204.360 ;
        RECT 12.840 204.040 13.160 204.360 ;
        RECT 13.240 204.040 13.560 204.360 ;
        RECT 13.640 204.040 13.960 204.360 ;
        RECT 14.040 204.040 14.360 204.360 ;
        RECT 14.440 204.040 14.760 204.360 ;
        RECT 14.840 204.040 15.160 204.360 ;
        RECT 15.240 204.040 15.560 204.360 ;
        RECT 15.640 204.040 15.960 204.360 ;
        RECT 16.040 204.040 16.360 204.360 ;
        RECT 16.440 204.040 16.760 204.360 ;
        RECT 16.840 204.040 17.160 204.360 ;
        RECT 17.240 204.040 17.560 204.360 ;
        RECT 17.640 204.040 17.960 204.360 ;
        RECT 18.040 204.040 18.360 204.360 ;
        RECT 18.440 204.040 18.760 204.360 ;
        RECT 18.840 204.040 19.160 204.360 ;
        RECT 19.240 204.040 19.560 204.360 ;
        RECT 19.640 204.040 19.960 204.360 ;
        RECT 95.560 204.040 95.880 204.360 ;
        RECT 95.960 204.040 96.280 204.360 ;
        RECT 96.360 204.040 96.680 204.360 ;
        RECT 96.760 204.040 97.080 204.360 ;
        RECT 145.560 204.040 145.880 204.360 ;
        RECT 145.960 204.040 146.280 204.360 ;
        RECT 146.360 204.040 146.680 204.360 ;
        RECT 146.760 204.040 147.080 204.360 ;
        RECT 185.720 204.040 186.040 204.360 ;
        RECT 186.120 204.040 186.440 204.360 ;
        RECT 186.520 204.040 186.840 204.360 ;
        RECT 186.920 204.040 187.240 204.360 ;
        RECT 187.320 204.040 187.640 204.360 ;
        RECT 187.720 204.040 188.040 204.360 ;
        RECT 188.120 204.040 188.440 204.360 ;
        RECT 188.520 204.040 188.840 204.360 ;
        RECT 188.920 204.040 189.240 204.360 ;
        RECT 189.320 204.040 189.640 204.360 ;
        RECT 189.720 204.040 190.040 204.360 ;
        RECT 190.120 204.040 190.440 204.360 ;
        RECT 190.520 204.040 190.840 204.360 ;
        RECT 190.920 204.040 191.240 204.360 ;
        RECT 191.320 204.040 191.640 204.360 ;
        RECT 191.720 204.040 192.040 204.360 ;
        RECT 192.120 204.040 192.440 204.360 ;
        RECT 192.520 204.040 192.840 204.360 ;
        RECT 192.920 204.040 193.240 204.360 ;
        RECT 193.320 204.040 193.640 204.360 ;
        RECT 193.720 204.040 194.040 204.360 ;
        RECT 194.120 204.040 194.440 204.360 ;
        RECT 194.520 204.040 194.840 204.360 ;
        RECT 194.920 204.040 195.240 204.360 ;
        RECT 195.320 204.040 195.640 204.360 ;
        RECT 195.720 204.040 196.040 204.360 ;
        RECT 196.120 204.040 196.440 204.360 ;
        RECT 196.520 204.040 196.840 204.360 ;
        RECT 196.920 204.040 197.240 204.360 ;
        RECT 197.320 204.040 197.640 204.360 ;
        RECT 197.720 204.040 198.040 204.360 ;
        RECT 198.120 204.040 198.440 204.360 ;
        RECT 198.520 204.040 198.840 204.360 ;
        RECT 198.920 204.040 199.240 204.360 ;
        RECT 199.320 204.040 199.640 204.360 ;
        RECT 199.720 204.040 200.040 204.360 ;
        RECT 200.120 204.040 200.440 204.360 ;
        RECT 200.520 204.040 200.840 204.360 ;
        RECT 200.920 204.040 201.240 204.360 ;
        RECT 201.320 204.040 201.640 204.360 ;
        RECT 201.720 204.040 202.040 204.360 ;
        RECT 202.120 204.040 202.440 204.360 ;
        RECT 202.520 204.040 202.840 204.360 ;
        RECT 202.920 204.040 203.240 204.360 ;
        RECT 203.320 204.040 203.640 204.360 ;
        RECT 203.720 204.040 204.040 204.360 ;
        RECT 204.120 204.040 204.440 204.360 ;
        RECT 204.520 204.040 204.840 204.360 ;
        RECT 204.920 204.040 205.240 204.360 ;
        RECT 205.320 204.040 205.640 204.360 ;
        RECT 0.040 203.640 0.360 203.960 ;
        RECT 0.440 203.640 0.760 203.960 ;
        RECT 0.840 203.640 1.160 203.960 ;
        RECT 1.240 203.640 1.560 203.960 ;
        RECT 1.640 203.640 1.960 203.960 ;
        RECT 2.040 203.640 2.360 203.960 ;
        RECT 2.440 203.640 2.760 203.960 ;
        RECT 2.840 203.640 3.160 203.960 ;
        RECT 3.240 203.640 3.560 203.960 ;
        RECT 3.640 203.640 3.960 203.960 ;
        RECT 4.040 203.640 4.360 203.960 ;
        RECT 4.440 203.640 4.760 203.960 ;
        RECT 4.840 203.640 5.160 203.960 ;
        RECT 5.240 203.640 5.560 203.960 ;
        RECT 5.640 203.640 5.960 203.960 ;
        RECT 6.040 203.640 6.360 203.960 ;
        RECT 6.440 203.640 6.760 203.960 ;
        RECT 6.840 203.640 7.160 203.960 ;
        RECT 7.240 203.640 7.560 203.960 ;
        RECT 7.640 203.640 7.960 203.960 ;
        RECT 8.040 203.640 8.360 203.960 ;
        RECT 8.440 203.640 8.760 203.960 ;
        RECT 8.840 203.640 9.160 203.960 ;
        RECT 9.240 203.640 9.560 203.960 ;
        RECT 9.640 203.640 9.960 203.960 ;
        RECT 10.040 203.640 10.360 203.960 ;
        RECT 10.440 203.640 10.760 203.960 ;
        RECT 10.840 203.640 11.160 203.960 ;
        RECT 11.240 203.640 11.560 203.960 ;
        RECT 11.640 203.640 11.960 203.960 ;
        RECT 12.040 203.640 12.360 203.960 ;
        RECT 12.440 203.640 12.760 203.960 ;
        RECT 12.840 203.640 13.160 203.960 ;
        RECT 13.240 203.640 13.560 203.960 ;
        RECT 13.640 203.640 13.960 203.960 ;
        RECT 14.040 203.640 14.360 203.960 ;
        RECT 14.440 203.640 14.760 203.960 ;
        RECT 14.840 203.640 15.160 203.960 ;
        RECT 15.240 203.640 15.560 203.960 ;
        RECT 15.640 203.640 15.960 203.960 ;
        RECT 16.040 203.640 16.360 203.960 ;
        RECT 16.440 203.640 16.760 203.960 ;
        RECT 16.840 203.640 17.160 203.960 ;
        RECT 17.240 203.640 17.560 203.960 ;
        RECT 17.640 203.640 17.960 203.960 ;
        RECT 18.040 203.640 18.360 203.960 ;
        RECT 18.440 203.640 18.760 203.960 ;
        RECT 18.840 203.640 19.160 203.960 ;
        RECT 19.240 203.640 19.560 203.960 ;
        RECT 19.640 203.640 19.960 203.960 ;
        RECT 95.560 203.640 95.880 203.960 ;
        RECT 95.960 203.640 96.280 203.960 ;
        RECT 96.360 203.640 96.680 203.960 ;
        RECT 96.760 203.640 97.080 203.960 ;
        RECT 145.560 203.640 145.880 203.960 ;
        RECT 145.960 203.640 146.280 203.960 ;
        RECT 146.360 203.640 146.680 203.960 ;
        RECT 146.760 203.640 147.080 203.960 ;
        RECT 185.720 203.640 186.040 203.960 ;
        RECT 186.120 203.640 186.440 203.960 ;
        RECT 186.520 203.640 186.840 203.960 ;
        RECT 186.920 203.640 187.240 203.960 ;
        RECT 187.320 203.640 187.640 203.960 ;
        RECT 187.720 203.640 188.040 203.960 ;
        RECT 188.120 203.640 188.440 203.960 ;
        RECT 188.520 203.640 188.840 203.960 ;
        RECT 188.920 203.640 189.240 203.960 ;
        RECT 189.320 203.640 189.640 203.960 ;
        RECT 189.720 203.640 190.040 203.960 ;
        RECT 190.120 203.640 190.440 203.960 ;
        RECT 190.520 203.640 190.840 203.960 ;
        RECT 190.920 203.640 191.240 203.960 ;
        RECT 191.320 203.640 191.640 203.960 ;
        RECT 191.720 203.640 192.040 203.960 ;
        RECT 192.120 203.640 192.440 203.960 ;
        RECT 192.520 203.640 192.840 203.960 ;
        RECT 192.920 203.640 193.240 203.960 ;
        RECT 193.320 203.640 193.640 203.960 ;
        RECT 193.720 203.640 194.040 203.960 ;
        RECT 194.120 203.640 194.440 203.960 ;
        RECT 194.520 203.640 194.840 203.960 ;
        RECT 194.920 203.640 195.240 203.960 ;
        RECT 195.320 203.640 195.640 203.960 ;
        RECT 195.720 203.640 196.040 203.960 ;
        RECT 196.120 203.640 196.440 203.960 ;
        RECT 196.520 203.640 196.840 203.960 ;
        RECT 196.920 203.640 197.240 203.960 ;
        RECT 197.320 203.640 197.640 203.960 ;
        RECT 197.720 203.640 198.040 203.960 ;
        RECT 198.120 203.640 198.440 203.960 ;
        RECT 198.520 203.640 198.840 203.960 ;
        RECT 198.920 203.640 199.240 203.960 ;
        RECT 199.320 203.640 199.640 203.960 ;
        RECT 199.720 203.640 200.040 203.960 ;
        RECT 200.120 203.640 200.440 203.960 ;
        RECT 200.520 203.640 200.840 203.960 ;
        RECT 200.920 203.640 201.240 203.960 ;
        RECT 201.320 203.640 201.640 203.960 ;
        RECT 201.720 203.640 202.040 203.960 ;
        RECT 202.120 203.640 202.440 203.960 ;
        RECT 202.520 203.640 202.840 203.960 ;
        RECT 202.920 203.640 203.240 203.960 ;
        RECT 203.320 203.640 203.640 203.960 ;
        RECT 203.720 203.640 204.040 203.960 ;
        RECT 204.120 203.640 204.440 203.960 ;
        RECT 204.520 203.640 204.840 203.960 ;
        RECT 204.920 203.640 205.240 203.960 ;
        RECT 205.320 203.640 205.640 203.960 ;
        RECT 0.040 203.240 0.360 203.560 ;
        RECT 0.440 203.240 0.760 203.560 ;
        RECT 0.840 203.240 1.160 203.560 ;
        RECT 1.240 203.240 1.560 203.560 ;
        RECT 1.640 203.240 1.960 203.560 ;
        RECT 2.040 203.240 2.360 203.560 ;
        RECT 2.440 203.240 2.760 203.560 ;
        RECT 2.840 203.240 3.160 203.560 ;
        RECT 3.240 203.240 3.560 203.560 ;
        RECT 3.640 203.240 3.960 203.560 ;
        RECT 4.040 203.240 4.360 203.560 ;
        RECT 4.440 203.240 4.760 203.560 ;
        RECT 4.840 203.240 5.160 203.560 ;
        RECT 5.240 203.240 5.560 203.560 ;
        RECT 5.640 203.240 5.960 203.560 ;
        RECT 6.040 203.240 6.360 203.560 ;
        RECT 6.440 203.240 6.760 203.560 ;
        RECT 6.840 203.240 7.160 203.560 ;
        RECT 7.240 203.240 7.560 203.560 ;
        RECT 7.640 203.240 7.960 203.560 ;
        RECT 8.040 203.240 8.360 203.560 ;
        RECT 8.440 203.240 8.760 203.560 ;
        RECT 8.840 203.240 9.160 203.560 ;
        RECT 9.240 203.240 9.560 203.560 ;
        RECT 9.640 203.240 9.960 203.560 ;
        RECT 10.040 203.240 10.360 203.560 ;
        RECT 10.440 203.240 10.760 203.560 ;
        RECT 10.840 203.240 11.160 203.560 ;
        RECT 11.240 203.240 11.560 203.560 ;
        RECT 11.640 203.240 11.960 203.560 ;
        RECT 12.040 203.240 12.360 203.560 ;
        RECT 12.440 203.240 12.760 203.560 ;
        RECT 12.840 203.240 13.160 203.560 ;
        RECT 13.240 203.240 13.560 203.560 ;
        RECT 13.640 203.240 13.960 203.560 ;
        RECT 14.040 203.240 14.360 203.560 ;
        RECT 14.440 203.240 14.760 203.560 ;
        RECT 14.840 203.240 15.160 203.560 ;
        RECT 15.240 203.240 15.560 203.560 ;
        RECT 15.640 203.240 15.960 203.560 ;
        RECT 16.040 203.240 16.360 203.560 ;
        RECT 16.440 203.240 16.760 203.560 ;
        RECT 16.840 203.240 17.160 203.560 ;
        RECT 17.240 203.240 17.560 203.560 ;
        RECT 17.640 203.240 17.960 203.560 ;
        RECT 18.040 203.240 18.360 203.560 ;
        RECT 18.440 203.240 18.760 203.560 ;
        RECT 18.840 203.240 19.160 203.560 ;
        RECT 19.240 203.240 19.560 203.560 ;
        RECT 19.640 203.240 19.960 203.560 ;
        RECT 95.560 203.240 95.880 203.560 ;
        RECT 95.960 203.240 96.280 203.560 ;
        RECT 96.360 203.240 96.680 203.560 ;
        RECT 96.760 203.240 97.080 203.560 ;
        RECT 145.560 203.240 145.880 203.560 ;
        RECT 145.960 203.240 146.280 203.560 ;
        RECT 146.360 203.240 146.680 203.560 ;
        RECT 146.760 203.240 147.080 203.560 ;
        RECT 185.720 203.240 186.040 203.560 ;
        RECT 186.120 203.240 186.440 203.560 ;
        RECT 186.520 203.240 186.840 203.560 ;
        RECT 186.920 203.240 187.240 203.560 ;
        RECT 187.320 203.240 187.640 203.560 ;
        RECT 187.720 203.240 188.040 203.560 ;
        RECT 188.120 203.240 188.440 203.560 ;
        RECT 188.520 203.240 188.840 203.560 ;
        RECT 188.920 203.240 189.240 203.560 ;
        RECT 189.320 203.240 189.640 203.560 ;
        RECT 189.720 203.240 190.040 203.560 ;
        RECT 190.120 203.240 190.440 203.560 ;
        RECT 190.520 203.240 190.840 203.560 ;
        RECT 190.920 203.240 191.240 203.560 ;
        RECT 191.320 203.240 191.640 203.560 ;
        RECT 191.720 203.240 192.040 203.560 ;
        RECT 192.120 203.240 192.440 203.560 ;
        RECT 192.520 203.240 192.840 203.560 ;
        RECT 192.920 203.240 193.240 203.560 ;
        RECT 193.320 203.240 193.640 203.560 ;
        RECT 193.720 203.240 194.040 203.560 ;
        RECT 194.120 203.240 194.440 203.560 ;
        RECT 194.520 203.240 194.840 203.560 ;
        RECT 194.920 203.240 195.240 203.560 ;
        RECT 195.320 203.240 195.640 203.560 ;
        RECT 195.720 203.240 196.040 203.560 ;
        RECT 196.120 203.240 196.440 203.560 ;
        RECT 196.520 203.240 196.840 203.560 ;
        RECT 196.920 203.240 197.240 203.560 ;
        RECT 197.320 203.240 197.640 203.560 ;
        RECT 197.720 203.240 198.040 203.560 ;
        RECT 198.120 203.240 198.440 203.560 ;
        RECT 198.520 203.240 198.840 203.560 ;
        RECT 198.920 203.240 199.240 203.560 ;
        RECT 199.320 203.240 199.640 203.560 ;
        RECT 199.720 203.240 200.040 203.560 ;
        RECT 200.120 203.240 200.440 203.560 ;
        RECT 200.520 203.240 200.840 203.560 ;
        RECT 200.920 203.240 201.240 203.560 ;
        RECT 201.320 203.240 201.640 203.560 ;
        RECT 201.720 203.240 202.040 203.560 ;
        RECT 202.120 203.240 202.440 203.560 ;
        RECT 202.520 203.240 202.840 203.560 ;
        RECT 202.920 203.240 203.240 203.560 ;
        RECT 203.320 203.240 203.640 203.560 ;
        RECT 203.720 203.240 204.040 203.560 ;
        RECT 204.120 203.240 204.440 203.560 ;
        RECT 204.520 203.240 204.840 203.560 ;
        RECT 204.920 203.240 205.240 203.560 ;
        RECT 205.320 203.240 205.640 203.560 ;
        RECT 0.040 202.840 0.360 203.160 ;
        RECT 0.440 202.840 0.760 203.160 ;
        RECT 0.840 202.840 1.160 203.160 ;
        RECT 1.240 202.840 1.560 203.160 ;
        RECT 1.640 202.840 1.960 203.160 ;
        RECT 2.040 202.840 2.360 203.160 ;
        RECT 2.440 202.840 2.760 203.160 ;
        RECT 2.840 202.840 3.160 203.160 ;
        RECT 3.240 202.840 3.560 203.160 ;
        RECT 3.640 202.840 3.960 203.160 ;
        RECT 4.040 202.840 4.360 203.160 ;
        RECT 4.440 202.840 4.760 203.160 ;
        RECT 4.840 202.840 5.160 203.160 ;
        RECT 5.240 202.840 5.560 203.160 ;
        RECT 5.640 202.840 5.960 203.160 ;
        RECT 6.040 202.840 6.360 203.160 ;
        RECT 6.440 202.840 6.760 203.160 ;
        RECT 6.840 202.840 7.160 203.160 ;
        RECT 7.240 202.840 7.560 203.160 ;
        RECT 7.640 202.840 7.960 203.160 ;
        RECT 8.040 202.840 8.360 203.160 ;
        RECT 8.440 202.840 8.760 203.160 ;
        RECT 8.840 202.840 9.160 203.160 ;
        RECT 9.240 202.840 9.560 203.160 ;
        RECT 9.640 202.840 9.960 203.160 ;
        RECT 10.040 202.840 10.360 203.160 ;
        RECT 10.440 202.840 10.760 203.160 ;
        RECT 10.840 202.840 11.160 203.160 ;
        RECT 11.240 202.840 11.560 203.160 ;
        RECT 11.640 202.840 11.960 203.160 ;
        RECT 12.040 202.840 12.360 203.160 ;
        RECT 12.440 202.840 12.760 203.160 ;
        RECT 12.840 202.840 13.160 203.160 ;
        RECT 13.240 202.840 13.560 203.160 ;
        RECT 13.640 202.840 13.960 203.160 ;
        RECT 14.040 202.840 14.360 203.160 ;
        RECT 14.440 202.840 14.760 203.160 ;
        RECT 14.840 202.840 15.160 203.160 ;
        RECT 15.240 202.840 15.560 203.160 ;
        RECT 15.640 202.840 15.960 203.160 ;
        RECT 16.040 202.840 16.360 203.160 ;
        RECT 16.440 202.840 16.760 203.160 ;
        RECT 16.840 202.840 17.160 203.160 ;
        RECT 17.240 202.840 17.560 203.160 ;
        RECT 17.640 202.840 17.960 203.160 ;
        RECT 18.040 202.840 18.360 203.160 ;
        RECT 18.440 202.840 18.760 203.160 ;
        RECT 18.840 202.840 19.160 203.160 ;
        RECT 19.240 202.840 19.560 203.160 ;
        RECT 19.640 202.840 19.960 203.160 ;
        RECT 95.560 202.840 95.880 203.160 ;
        RECT 95.960 202.840 96.280 203.160 ;
        RECT 96.360 202.840 96.680 203.160 ;
        RECT 96.760 202.840 97.080 203.160 ;
        RECT 145.560 202.840 145.880 203.160 ;
        RECT 145.960 202.840 146.280 203.160 ;
        RECT 146.360 202.840 146.680 203.160 ;
        RECT 146.760 202.840 147.080 203.160 ;
        RECT 185.720 202.840 186.040 203.160 ;
        RECT 186.120 202.840 186.440 203.160 ;
        RECT 186.520 202.840 186.840 203.160 ;
        RECT 186.920 202.840 187.240 203.160 ;
        RECT 187.320 202.840 187.640 203.160 ;
        RECT 187.720 202.840 188.040 203.160 ;
        RECT 188.120 202.840 188.440 203.160 ;
        RECT 188.520 202.840 188.840 203.160 ;
        RECT 188.920 202.840 189.240 203.160 ;
        RECT 189.320 202.840 189.640 203.160 ;
        RECT 189.720 202.840 190.040 203.160 ;
        RECT 190.120 202.840 190.440 203.160 ;
        RECT 190.520 202.840 190.840 203.160 ;
        RECT 190.920 202.840 191.240 203.160 ;
        RECT 191.320 202.840 191.640 203.160 ;
        RECT 191.720 202.840 192.040 203.160 ;
        RECT 192.120 202.840 192.440 203.160 ;
        RECT 192.520 202.840 192.840 203.160 ;
        RECT 192.920 202.840 193.240 203.160 ;
        RECT 193.320 202.840 193.640 203.160 ;
        RECT 193.720 202.840 194.040 203.160 ;
        RECT 194.120 202.840 194.440 203.160 ;
        RECT 194.520 202.840 194.840 203.160 ;
        RECT 194.920 202.840 195.240 203.160 ;
        RECT 195.320 202.840 195.640 203.160 ;
        RECT 195.720 202.840 196.040 203.160 ;
        RECT 196.120 202.840 196.440 203.160 ;
        RECT 196.520 202.840 196.840 203.160 ;
        RECT 196.920 202.840 197.240 203.160 ;
        RECT 197.320 202.840 197.640 203.160 ;
        RECT 197.720 202.840 198.040 203.160 ;
        RECT 198.120 202.840 198.440 203.160 ;
        RECT 198.520 202.840 198.840 203.160 ;
        RECT 198.920 202.840 199.240 203.160 ;
        RECT 199.320 202.840 199.640 203.160 ;
        RECT 199.720 202.840 200.040 203.160 ;
        RECT 200.120 202.840 200.440 203.160 ;
        RECT 200.520 202.840 200.840 203.160 ;
        RECT 200.920 202.840 201.240 203.160 ;
        RECT 201.320 202.840 201.640 203.160 ;
        RECT 201.720 202.840 202.040 203.160 ;
        RECT 202.120 202.840 202.440 203.160 ;
        RECT 202.520 202.840 202.840 203.160 ;
        RECT 202.920 202.840 203.240 203.160 ;
        RECT 203.320 202.840 203.640 203.160 ;
        RECT 203.720 202.840 204.040 203.160 ;
        RECT 204.120 202.840 204.440 203.160 ;
        RECT 204.520 202.840 204.840 203.160 ;
        RECT 204.920 202.840 205.240 203.160 ;
        RECT 205.320 202.840 205.640 203.160 ;
        RECT 0.040 202.440 0.360 202.760 ;
        RECT 0.440 202.440 0.760 202.760 ;
        RECT 0.840 202.440 1.160 202.760 ;
        RECT 1.240 202.440 1.560 202.760 ;
        RECT 1.640 202.440 1.960 202.760 ;
        RECT 2.040 202.440 2.360 202.760 ;
        RECT 2.440 202.440 2.760 202.760 ;
        RECT 2.840 202.440 3.160 202.760 ;
        RECT 3.240 202.440 3.560 202.760 ;
        RECT 3.640 202.440 3.960 202.760 ;
        RECT 4.040 202.440 4.360 202.760 ;
        RECT 4.440 202.440 4.760 202.760 ;
        RECT 4.840 202.440 5.160 202.760 ;
        RECT 5.240 202.440 5.560 202.760 ;
        RECT 5.640 202.440 5.960 202.760 ;
        RECT 6.040 202.440 6.360 202.760 ;
        RECT 6.440 202.440 6.760 202.760 ;
        RECT 6.840 202.440 7.160 202.760 ;
        RECT 7.240 202.440 7.560 202.760 ;
        RECT 7.640 202.440 7.960 202.760 ;
        RECT 8.040 202.440 8.360 202.760 ;
        RECT 8.440 202.440 8.760 202.760 ;
        RECT 8.840 202.440 9.160 202.760 ;
        RECT 9.240 202.440 9.560 202.760 ;
        RECT 9.640 202.440 9.960 202.760 ;
        RECT 10.040 202.440 10.360 202.760 ;
        RECT 10.440 202.440 10.760 202.760 ;
        RECT 10.840 202.440 11.160 202.760 ;
        RECT 11.240 202.440 11.560 202.760 ;
        RECT 11.640 202.440 11.960 202.760 ;
        RECT 12.040 202.440 12.360 202.760 ;
        RECT 12.440 202.440 12.760 202.760 ;
        RECT 12.840 202.440 13.160 202.760 ;
        RECT 13.240 202.440 13.560 202.760 ;
        RECT 13.640 202.440 13.960 202.760 ;
        RECT 14.040 202.440 14.360 202.760 ;
        RECT 14.440 202.440 14.760 202.760 ;
        RECT 14.840 202.440 15.160 202.760 ;
        RECT 15.240 202.440 15.560 202.760 ;
        RECT 15.640 202.440 15.960 202.760 ;
        RECT 16.040 202.440 16.360 202.760 ;
        RECT 16.440 202.440 16.760 202.760 ;
        RECT 16.840 202.440 17.160 202.760 ;
        RECT 17.240 202.440 17.560 202.760 ;
        RECT 17.640 202.440 17.960 202.760 ;
        RECT 18.040 202.440 18.360 202.760 ;
        RECT 18.440 202.440 18.760 202.760 ;
        RECT 18.840 202.440 19.160 202.760 ;
        RECT 19.240 202.440 19.560 202.760 ;
        RECT 19.640 202.440 19.960 202.760 ;
        RECT 95.560 202.440 95.880 202.760 ;
        RECT 95.960 202.440 96.280 202.760 ;
        RECT 96.360 202.440 96.680 202.760 ;
        RECT 96.760 202.440 97.080 202.760 ;
        RECT 145.560 202.440 145.880 202.760 ;
        RECT 145.960 202.440 146.280 202.760 ;
        RECT 146.360 202.440 146.680 202.760 ;
        RECT 146.760 202.440 147.080 202.760 ;
        RECT 185.720 202.440 186.040 202.760 ;
        RECT 186.120 202.440 186.440 202.760 ;
        RECT 186.520 202.440 186.840 202.760 ;
        RECT 186.920 202.440 187.240 202.760 ;
        RECT 187.320 202.440 187.640 202.760 ;
        RECT 187.720 202.440 188.040 202.760 ;
        RECT 188.120 202.440 188.440 202.760 ;
        RECT 188.520 202.440 188.840 202.760 ;
        RECT 188.920 202.440 189.240 202.760 ;
        RECT 189.320 202.440 189.640 202.760 ;
        RECT 189.720 202.440 190.040 202.760 ;
        RECT 190.120 202.440 190.440 202.760 ;
        RECT 190.520 202.440 190.840 202.760 ;
        RECT 190.920 202.440 191.240 202.760 ;
        RECT 191.320 202.440 191.640 202.760 ;
        RECT 191.720 202.440 192.040 202.760 ;
        RECT 192.120 202.440 192.440 202.760 ;
        RECT 192.520 202.440 192.840 202.760 ;
        RECT 192.920 202.440 193.240 202.760 ;
        RECT 193.320 202.440 193.640 202.760 ;
        RECT 193.720 202.440 194.040 202.760 ;
        RECT 194.120 202.440 194.440 202.760 ;
        RECT 194.520 202.440 194.840 202.760 ;
        RECT 194.920 202.440 195.240 202.760 ;
        RECT 195.320 202.440 195.640 202.760 ;
        RECT 195.720 202.440 196.040 202.760 ;
        RECT 196.120 202.440 196.440 202.760 ;
        RECT 196.520 202.440 196.840 202.760 ;
        RECT 196.920 202.440 197.240 202.760 ;
        RECT 197.320 202.440 197.640 202.760 ;
        RECT 197.720 202.440 198.040 202.760 ;
        RECT 198.120 202.440 198.440 202.760 ;
        RECT 198.520 202.440 198.840 202.760 ;
        RECT 198.920 202.440 199.240 202.760 ;
        RECT 199.320 202.440 199.640 202.760 ;
        RECT 199.720 202.440 200.040 202.760 ;
        RECT 200.120 202.440 200.440 202.760 ;
        RECT 200.520 202.440 200.840 202.760 ;
        RECT 200.920 202.440 201.240 202.760 ;
        RECT 201.320 202.440 201.640 202.760 ;
        RECT 201.720 202.440 202.040 202.760 ;
        RECT 202.120 202.440 202.440 202.760 ;
        RECT 202.520 202.440 202.840 202.760 ;
        RECT 202.920 202.440 203.240 202.760 ;
        RECT 203.320 202.440 203.640 202.760 ;
        RECT 203.720 202.440 204.040 202.760 ;
        RECT 204.120 202.440 204.440 202.760 ;
        RECT 204.520 202.440 204.840 202.760 ;
        RECT 204.920 202.440 205.240 202.760 ;
        RECT 205.320 202.440 205.640 202.760 ;
        RECT 0.040 202.040 0.360 202.360 ;
        RECT 0.440 202.040 0.760 202.360 ;
        RECT 0.840 202.040 1.160 202.360 ;
        RECT 1.240 202.040 1.560 202.360 ;
        RECT 1.640 202.040 1.960 202.360 ;
        RECT 2.040 202.040 2.360 202.360 ;
        RECT 2.440 202.040 2.760 202.360 ;
        RECT 2.840 202.040 3.160 202.360 ;
        RECT 3.240 202.040 3.560 202.360 ;
        RECT 3.640 202.040 3.960 202.360 ;
        RECT 4.040 202.040 4.360 202.360 ;
        RECT 4.440 202.040 4.760 202.360 ;
        RECT 4.840 202.040 5.160 202.360 ;
        RECT 5.240 202.040 5.560 202.360 ;
        RECT 5.640 202.040 5.960 202.360 ;
        RECT 6.040 202.040 6.360 202.360 ;
        RECT 6.440 202.040 6.760 202.360 ;
        RECT 6.840 202.040 7.160 202.360 ;
        RECT 7.240 202.040 7.560 202.360 ;
        RECT 7.640 202.040 7.960 202.360 ;
        RECT 8.040 202.040 8.360 202.360 ;
        RECT 8.440 202.040 8.760 202.360 ;
        RECT 8.840 202.040 9.160 202.360 ;
        RECT 9.240 202.040 9.560 202.360 ;
        RECT 9.640 202.040 9.960 202.360 ;
        RECT 10.040 202.040 10.360 202.360 ;
        RECT 10.440 202.040 10.760 202.360 ;
        RECT 10.840 202.040 11.160 202.360 ;
        RECT 11.240 202.040 11.560 202.360 ;
        RECT 11.640 202.040 11.960 202.360 ;
        RECT 12.040 202.040 12.360 202.360 ;
        RECT 12.440 202.040 12.760 202.360 ;
        RECT 12.840 202.040 13.160 202.360 ;
        RECT 13.240 202.040 13.560 202.360 ;
        RECT 13.640 202.040 13.960 202.360 ;
        RECT 14.040 202.040 14.360 202.360 ;
        RECT 14.440 202.040 14.760 202.360 ;
        RECT 14.840 202.040 15.160 202.360 ;
        RECT 15.240 202.040 15.560 202.360 ;
        RECT 15.640 202.040 15.960 202.360 ;
        RECT 16.040 202.040 16.360 202.360 ;
        RECT 16.440 202.040 16.760 202.360 ;
        RECT 16.840 202.040 17.160 202.360 ;
        RECT 17.240 202.040 17.560 202.360 ;
        RECT 17.640 202.040 17.960 202.360 ;
        RECT 18.040 202.040 18.360 202.360 ;
        RECT 18.440 202.040 18.760 202.360 ;
        RECT 18.840 202.040 19.160 202.360 ;
        RECT 19.240 202.040 19.560 202.360 ;
        RECT 19.640 202.040 19.960 202.360 ;
        RECT 95.560 202.040 95.880 202.360 ;
        RECT 95.960 202.040 96.280 202.360 ;
        RECT 96.360 202.040 96.680 202.360 ;
        RECT 96.760 202.040 97.080 202.360 ;
        RECT 145.560 202.040 145.880 202.360 ;
        RECT 145.960 202.040 146.280 202.360 ;
        RECT 146.360 202.040 146.680 202.360 ;
        RECT 146.760 202.040 147.080 202.360 ;
        RECT 185.720 202.040 186.040 202.360 ;
        RECT 186.120 202.040 186.440 202.360 ;
        RECT 186.520 202.040 186.840 202.360 ;
        RECT 186.920 202.040 187.240 202.360 ;
        RECT 187.320 202.040 187.640 202.360 ;
        RECT 187.720 202.040 188.040 202.360 ;
        RECT 188.120 202.040 188.440 202.360 ;
        RECT 188.520 202.040 188.840 202.360 ;
        RECT 188.920 202.040 189.240 202.360 ;
        RECT 189.320 202.040 189.640 202.360 ;
        RECT 189.720 202.040 190.040 202.360 ;
        RECT 190.120 202.040 190.440 202.360 ;
        RECT 190.520 202.040 190.840 202.360 ;
        RECT 190.920 202.040 191.240 202.360 ;
        RECT 191.320 202.040 191.640 202.360 ;
        RECT 191.720 202.040 192.040 202.360 ;
        RECT 192.120 202.040 192.440 202.360 ;
        RECT 192.520 202.040 192.840 202.360 ;
        RECT 192.920 202.040 193.240 202.360 ;
        RECT 193.320 202.040 193.640 202.360 ;
        RECT 193.720 202.040 194.040 202.360 ;
        RECT 194.120 202.040 194.440 202.360 ;
        RECT 194.520 202.040 194.840 202.360 ;
        RECT 194.920 202.040 195.240 202.360 ;
        RECT 195.320 202.040 195.640 202.360 ;
        RECT 195.720 202.040 196.040 202.360 ;
        RECT 196.120 202.040 196.440 202.360 ;
        RECT 196.520 202.040 196.840 202.360 ;
        RECT 196.920 202.040 197.240 202.360 ;
        RECT 197.320 202.040 197.640 202.360 ;
        RECT 197.720 202.040 198.040 202.360 ;
        RECT 198.120 202.040 198.440 202.360 ;
        RECT 198.520 202.040 198.840 202.360 ;
        RECT 198.920 202.040 199.240 202.360 ;
        RECT 199.320 202.040 199.640 202.360 ;
        RECT 199.720 202.040 200.040 202.360 ;
        RECT 200.120 202.040 200.440 202.360 ;
        RECT 200.520 202.040 200.840 202.360 ;
        RECT 200.920 202.040 201.240 202.360 ;
        RECT 201.320 202.040 201.640 202.360 ;
        RECT 201.720 202.040 202.040 202.360 ;
        RECT 202.120 202.040 202.440 202.360 ;
        RECT 202.520 202.040 202.840 202.360 ;
        RECT 202.920 202.040 203.240 202.360 ;
        RECT 203.320 202.040 203.640 202.360 ;
        RECT 203.720 202.040 204.040 202.360 ;
        RECT 204.120 202.040 204.440 202.360 ;
        RECT 204.520 202.040 204.840 202.360 ;
        RECT 204.920 202.040 205.240 202.360 ;
        RECT 205.320 202.040 205.640 202.360 ;
        RECT 0.040 201.640 0.360 201.960 ;
        RECT 0.440 201.640 0.760 201.960 ;
        RECT 0.840 201.640 1.160 201.960 ;
        RECT 1.240 201.640 1.560 201.960 ;
        RECT 1.640 201.640 1.960 201.960 ;
        RECT 2.040 201.640 2.360 201.960 ;
        RECT 2.440 201.640 2.760 201.960 ;
        RECT 2.840 201.640 3.160 201.960 ;
        RECT 3.240 201.640 3.560 201.960 ;
        RECT 3.640 201.640 3.960 201.960 ;
        RECT 4.040 201.640 4.360 201.960 ;
        RECT 4.440 201.640 4.760 201.960 ;
        RECT 4.840 201.640 5.160 201.960 ;
        RECT 5.240 201.640 5.560 201.960 ;
        RECT 5.640 201.640 5.960 201.960 ;
        RECT 6.040 201.640 6.360 201.960 ;
        RECT 6.440 201.640 6.760 201.960 ;
        RECT 6.840 201.640 7.160 201.960 ;
        RECT 7.240 201.640 7.560 201.960 ;
        RECT 7.640 201.640 7.960 201.960 ;
        RECT 8.040 201.640 8.360 201.960 ;
        RECT 8.440 201.640 8.760 201.960 ;
        RECT 8.840 201.640 9.160 201.960 ;
        RECT 9.240 201.640 9.560 201.960 ;
        RECT 9.640 201.640 9.960 201.960 ;
        RECT 10.040 201.640 10.360 201.960 ;
        RECT 10.440 201.640 10.760 201.960 ;
        RECT 10.840 201.640 11.160 201.960 ;
        RECT 11.240 201.640 11.560 201.960 ;
        RECT 11.640 201.640 11.960 201.960 ;
        RECT 12.040 201.640 12.360 201.960 ;
        RECT 12.440 201.640 12.760 201.960 ;
        RECT 12.840 201.640 13.160 201.960 ;
        RECT 13.240 201.640 13.560 201.960 ;
        RECT 13.640 201.640 13.960 201.960 ;
        RECT 14.040 201.640 14.360 201.960 ;
        RECT 14.440 201.640 14.760 201.960 ;
        RECT 14.840 201.640 15.160 201.960 ;
        RECT 15.240 201.640 15.560 201.960 ;
        RECT 15.640 201.640 15.960 201.960 ;
        RECT 16.040 201.640 16.360 201.960 ;
        RECT 16.440 201.640 16.760 201.960 ;
        RECT 16.840 201.640 17.160 201.960 ;
        RECT 17.240 201.640 17.560 201.960 ;
        RECT 17.640 201.640 17.960 201.960 ;
        RECT 18.040 201.640 18.360 201.960 ;
        RECT 18.440 201.640 18.760 201.960 ;
        RECT 18.840 201.640 19.160 201.960 ;
        RECT 19.240 201.640 19.560 201.960 ;
        RECT 19.640 201.640 19.960 201.960 ;
        RECT 95.560 201.640 95.880 201.960 ;
        RECT 95.960 201.640 96.280 201.960 ;
        RECT 96.360 201.640 96.680 201.960 ;
        RECT 96.760 201.640 97.080 201.960 ;
        RECT 145.560 201.640 145.880 201.960 ;
        RECT 145.960 201.640 146.280 201.960 ;
        RECT 146.360 201.640 146.680 201.960 ;
        RECT 146.760 201.640 147.080 201.960 ;
        RECT 185.720 201.640 186.040 201.960 ;
        RECT 186.120 201.640 186.440 201.960 ;
        RECT 186.520 201.640 186.840 201.960 ;
        RECT 186.920 201.640 187.240 201.960 ;
        RECT 187.320 201.640 187.640 201.960 ;
        RECT 187.720 201.640 188.040 201.960 ;
        RECT 188.120 201.640 188.440 201.960 ;
        RECT 188.520 201.640 188.840 201.960 ;
        RECT 188.920 201.640 189.240 201.960 ;
        RECT 189.320 201.640 189.640 201.960 ;
        RECT 189.720 201.640 190.040 201.960 ;
        RECT 190.120 201.640 190.440 201.960 ;
        RECT 190.520 201.640 190.840 201.960 ;
        RECT 190.920 201.640 191.240 201.960 ;
        RECT 191.320 201.640 191.640 201.960 ;
        RECT 191.720 201.640 192.040 201.960 ;
        RECT 192.120 201.640 192.440 201.960 ;
        RECT 192.520 201.640 192.840 201.960 ;
        RECT 192.920 201.640 193.240 201.960 ;
        RECT 193.320 201.640 193.640 201.960 ;
        RECT 193.720 201.640 194.040 201.960 ;
        RECT 194.120 201.640 194.440 201.960 ;
        RECT 194.520 201.640 194.840 201.960 ;
        RECT 194.920 201.640 195.240 201.960 ;
        RECT 195.320 201.640 195.640 201.960 ;
        RECT 195.720 201.640 196.040 201.960 ;
        RECT 196.120 201.640 196.440 201.960 ;
        RECT 196.520 201.640 196.840 201.960 ;
        RECT 196.920 201.640 197.240 201.960 ;
        RECT 197.320 201.640 197.640 201.960 ;
        RECT 197.720 201.640 198.040 201.960 ;
        RECT 198.120 201.640 198.440 201.960 ;
        RECT 198.520 201.640 198.840 201.960 ;
        RECT 198.920 201.640 199.240 201.960 ;
        RECT 199.320 201.640 199.640 201.960 ;
        RECT 199.720 201.640 200.040 201.960 ;
        RECT 200.120 201.640 200.440 201.960 ;
        RECT 200.520 201.640 200.840 201.960 ;
        RECT 200.920 201.640 201.240 201.960 ;
        RECT 201.320 201.640 201.640 201.960 ;
        RECT 201.720 201.640 202.040 201.960 ;
        RECT 202.120 201.640 202.440 201.960 ;
        RECT 202.520 201.640 202.840 201.960 ;
        RECT 202.920 201.640 203.240 201.960 ;
        RECT 203.320 201.640 203.640 201.960 ;
        RECT 203.720 201.640 204.040 201.960 ;
        RECT 204.120 201.640 204.440 201.960 ;
        RECT 204.520 201.640 204.840 201.960 ;
        RECT 204.920 201.640 205.240 201.960 ;
        RECT 205.320 201.640 205.640 201.960 ;
        RECT 0.040 201.240 0.360 201.560 ;
        RECT 0.440 201.240 0.760 201.560 ;
        RECT 0.840 201.240 1.160 201.560 ;
        RECT 1.240 201.240 1.560 201.560 ;
        RECT 1.640 201.240 1.960 201.560 ;
        RECT 2.040 201.240 2.360 201.560 ;
        RECT 2.440 201.240 2.760 201.560 ;
        RECT 2.840 201.240 3.160 201.560 ;
        RECT 3.240 201.240 3.560 201.560 ;
        RECT 3.640 201.240 3.960 201.560 ;
        RECT 4.040 201.240 4.360 201.560 ;
        RECT 4.440 201.240 4.760 201.560 ;
        RECT 4.840 201.240 5.160 201.560 ;
        RECT 5.240 201.240 5.560 201.560 ;
        RECT 5.640 201.240 5.960 201.560 ;
        RECT 6.040 201.240 6.360 201.560 ;
        RECT 6.440 201.240 6.760 201.560 ;
        RECT 6.840 201.240 7.160 201.560 ;
        RECT 7.240 201.240 7.560 201.560 ;
        RECT 7.640 201.240 7.960 201.560 ;
        RECT 8.040 201.240 8.360 201.560 ;
        RECT 8.440 201.240 8.760 201.560 ;
        RECT 8.840 201.240 9.160 201.560 ;
        RECT 9.240 201.240 9.560 201.560 ;
        RECT 9.640 201.240 9.960 201.560 ;
        RECT 10.040 201.240 10.360 201.560 ;
        RECT 10.440 201.240 10.760 201.560 ;
        RECT 10.840 201.240 11.160 201.560 ;
        RECT 11.240 201.240 11.560 201.560 ;
        RECT 11.640 201.240 11.960 201.560 ;
        RECT 12.040 201.240 12.360 201.560 ;
        RECT 12.440 201.240 12.760 201.560 ;
        RECT 12.840 201.240 13.160 201.560 ;
        RECT 13.240 201.240 13.560 201.560 ;
        RECT 13.640 201.240 13.960 201.560 ;
        RECT 14.040 201.240 14.360 201.560 ;
        RECT 14.440 201.240 14.760 201.560 ;
        RECT 14.840 201.240 15.160 201.560 ;
        RECT 15.240 201.240 15.560 201.560 ;
        RECT 15.640 201.240 15.960 201.560 ;
        RECT 16.040 201.240 16.360 201.560 ;
        RECT 16.440 201.240 16.760 201.560 ;
        RECT 16.840 201.240 17.160 201.560 ;
        RECT 17.240 201.240 17.560 201.560 ;
        RECT 17.640 201.240 17.960 201.560 ;
        RECT 18.040 201.240 18.360 201.560 ;
        RECT 18.440 201.240 18.760 201.560 ;
        RECT 18.840 201.240 19.160 201.560 ;
        RECT 19.240 201.240 19.560 201.560 ;
        RECT 19.640 201.240 19.960 201.560 ;
        RECT 95.560 201.240 95.880 201.560 ;
        RECT 95.960 201.240 96.280 201.560 ;
        RECT 96.360 201.240 96.680 201.560 ;
        RECT 96.760 201.240 97.080 201.560 ;
        RECT 145.560 201.240 145.880 201.560 ;
        RECT 145.960 201.240 146.280 201.560 ;
        RECT 146.360 201.240 146.680 201.560 ;
        RECT 146.760 201.240 147.080 201.560 ;
        RECT 185.720 201.240 186.040 201.560 ;
        RECT 186.120 201.240 186.440 201.560 ;
        RECT 186.520 201.240 186.840 201.560 ;
        RECT 186.920 201.240 187.240 201.560 ;
        RECT 187.320 201.240 187.640 201.560 ;
        RECT 187.720 201.240 188.040 201.560 ;
        RECT 188.120 201.240 188.440 201.560 ;
        RECT 188.520 201.240 188.840 201.560 ;
        RECT 188.920 201.240 189.240 201.560 ;
        RECT 189.320 201.240 189.640 201.560 ;
        RECT 189.720 201.240 190.040 201.560 ;
        RECT 190.120 201.240 190.440 201.560 ;
        RECT 190.520 201.240 190.840 201.560 ;
        RECT 190.920 201.240 191.240 201.560 ;
        RECT 191.320 201.240 191.640 201.560 ;
        RECT 191.720 201.240 192.040 201.560 ;
        RECT 192.120 201.240 192.440 201.560 ;
        RECT 192.520 201.240 192.840 201.560 ;
        RECT 192.920 201.240 193.240 201.560 ;
        RECT 193.320 201.240 193.640 201.560 ;
        RECT 193.720 201.240 194.040 201.560 ;
        RECT 194.120 201.240 194.440 201.560 ;
        RECT 194.520 201.240 194.840 201.560 ;
        RECT 194.920 201.240 195.240 201.560 ;
        RECT 195.320 201.240 195.640 201.560 ;
        RECT 195.720 201.240 196.040 201.560 ;
        RECT 196.120 201.240 196.440 201.560 ;
        RECT 196.520 201.240 196.840 201.560 ;
        RECT 196.920 201.240 197.240 201.560 ;
        RECT 197.320 201.240 197.640 201.560 ;
        RECT 197.720 201.240 198.040 201.560 ;
        RECT 198.120 201.240 198.440 201.560 ;
        RECT 198.520 201.240 198.840 201.560 ;
        RECT 198.920 201.240 199.240 201.560 ;
        RECT 199.320 201.240 199.640 201.560 ;
        RECT 199.720 201.240 200.040 201.560 ;
        RECT 200.120 201.240 200.440 201.560 ;
        RECT 200.520 201.240 200.840 201.560 ;
        RECT 200.920 201.240 201.240 201.560 ;
        RECT 201.320 201.240 201.640 201.560 ;
        RECT 201.720 201.240 202.040 201.560 ;
        RECT 202.120 201.240 202.440 201.560 ;
        RECT 202.520 201.240 202.840 201.560 ;
        RECT 202.920 201.240 203.240 201.560 ;
        RECT 203.320 201.240 203.640 201.560 ;
        RECT 203.720 201.240 204.040 201.560 ;
        RECT 204.120 201.240 204.440 201.560 ;
        RECT 204.520 201.240 204.840 201.560 ;
        RECT 204.920 201.240 205.240 201.560 ;
        RECT 205.320 201.240 205.640 201.560 ;
        RECT 0.040 200.840 0.360 201.160 ;
        RECT 0.440 200.840 0.760 201.160 ;
        RECT 0.840 200.840 1.160 201.160 ;
        RECT 1.240 200.840 1.560 201.160 ;
        RECT 1.640 200.840 1.960 201.160 ;
        RECT 2.040 200.840 2.360 201.160 ;
        RECT 2.440 200.840 2.760 201.160 ;
        RECT 2.840 200.840 3.160 201.160 ;
        RECT 3.240 200.840 3.560 201.160 ;
        RECT 3.640 200.840 3.960 201.160 ;
        RECT 4.040 200.840 4.360 201.160 ;
        RECT 4.440 200.840 4.760 201.160 ;
        RECT 4.840 200.840 5.160 201.160 ;
        RECT 5.240 200.840 5.560 201.160 ;
        RECT 5.640 200.840 5.960 201.160 ;
        RECT 6.040 200.840 6.360 201.160 ;
        RECT 6.440 200.840 6.760 201.160 ;
        RECT 6.840 200.840 7.160 201.160 ;
        RECT 7.240 200.840 7.560 201.160 ;
        RECT 7.640 200.840 7.960 201.160 ;
        RECT 8.040 200.840 8.360 201.160 ;
        RECT 8.440 200.840 8.760 201.160 ;
        RECT 8.840 200.840 9.160 201.160 ;
        RECT 9.240 200.840 9.560 201.160 ;
        RECT 9.640 200.840 9.960 201.160 ;
        RECT 10.040 200.840 10.360 201.160 ;
        RECT 10.440 200.840 10.760 201.160 ;
        RECT 10.840 200.840 11.160 201.160 ;
        RECT 11.240 200.840 11.560 201.160 ;
        RECT 11.640 200.840 11.960 201.160 ;
        RECT 12.040 200.840 12.360 201.160 ;
        RECT 12.440 200.840 12.760 201.160 ;
        RECT 12.840 200.840 13.160 201.160 ;
        RECT 13.240 200.840 13.560 201.160 ;
        RECT 13.640 200.840 13.960 201.160 ;
        RECT 14.040 200.840 14.360 201.160 ;
        RECT 14.440 200.840 14.760 201.160 ;
        RECT 14.840 200.840 15.160 201.160 ;
        RECT 15.240 200.840 15.560 201.160 ;
        RECT 15.640 200.840 15.960 201.160 ;
        RECT 16.040 200.840 16.360 201.160 ;
        RECT 16.440 200.840 16.760 201.160 ;
        RECT 16.840 200.840 17.160 201.160 ;
        RECT 17.240 200.840 17.560 201.160 ;
        RECT 17.640 200.840 17.960 201.160 ;
        RECT 18.040 200.840 18.360 201.160 ;
        RECT 18.440 200.840 18.760 201.160 ;
        RECT 18.840 200.840 19.160 201.160 ;
        RECT 19.240 200.840 19.560 201.160 ;
        RECT 19.640 200.840 19.960 201.160 ;
        RECT 95.560 200.840 95.880 201.160 ;
        RECT 95.960 200.840 96.280 201.160 ;
        RECT 96.360 200.840 96.680 201.160 ;
        RECT 96.760 200.840 97.080 201.160 ;
        RECT 145.560 200.840 145.880 201.160 ;
        RECT 145.960 200.840 146.280 201.160 ;
        RECT 146.360 200.840 146.680 201.160 ;
        RECT 146.760 200.840 147.080 201.160 ;
        RECT 185.720 200.840 186.040 201.160 ;
        RECT 186.120 200.840 186.440 201.160 ;
        RECT 186.520 200.840 186.840 201.160 ;
        RECT 186.920 200.840 187.240 201.160 ;
        RECT 187.320 200.840 187.640 201.160 ;
        RECT 187.720 200.840 188.040 201.160 ;
        RECT 188.120 200.840 188.440 201.160 ;
        RECT 188.520 200.840 188.840 201.160 ;
        RECT 188.920 200.840 189.240 201.160 ;
        RECT 189.320 200.840 189.640 201.160 ;
        RECT 189.720 200.840 190.040 201.160 ;
        RECT 190.120 200.840 190.440 201.160 ;
        RECT 190.520 200.840 190.840 201.160 ;
        RECT 190.920 200.840 191.240 201.160 ;
        RECT 191.320 200.840 191.640 201.160 ;
        RECT 191.720 200.840 192.040 201.160 ;
        RECT 192.120 200.840 192.440 201.160 ;
        RECT 192.520 200.840 192.840 201.160 ;
        RECT 192.920 200.840 193.240 201.160 ;
        RECT 193.320 200.840 193.640 201.160 ;
        RECT 193.720 200.840 194.040 201.160 ;
        RECT 194.120 200.840 194.440 201.160 ;
        RECT 194.520 200.840 194.840 201.160 ;
        RECT 194.920 200.840 195.240 201.160 ;
        RECT 195.320 200.840 195.640 201.160 ;
        RECT 195.720 200.840 196.040 201.160 ;
        RECT 196.120 200.840 196.440 201.160 ;
        RECT 196.520 200.840 196.840 201.160 ;
        RECT 196.920 200.840 197.240 201.160 ;
        RECT 197.320 200.840 197.640 201.160 ;
        RECT 197.720 200.840 198.040 201.160 ;
        RECT 198.120 200.840 198.440 201.160 ;
        RECT 198.520 200.840 198.840 201.160 ;
        RECT 198.920 200.840 199.240 201.160 ;
        RECT 199.320 200.840 199.640 201.160 ;
        RECT 199.720 200.840 200.040 201.160 ;
        RECT 200.120 200.840 200.440 201.160 ;
        RECT 200.520 200.840 200.840 201.160 ;
        RECT 200.920 200.840 201.240 201.160 ;
        RECT 201.320 200.840 201.640 201.160 ;
        RECT 201.720 200.840 202.040 201.160 ;
        RECT 202.120 200.840 202.440 201.160 ;
        RECT 202.520 200.840 202.840 201.160 ;
        RECT 202.920 200.840 203.240 201.160 ;
        RECT 203.320 200.840 203.640 201.160 ;
        RECT 203.720 200.840 204.040 201.160 ;
        RECT 204.120 200.840 204.440 201.160 ;
        RECT 204.520 200.840 204.840 201.160 ;
        RECT 204.920 200.840 205.240 201.160 ;
        RECT 205.320 200.840 205.640 201.160 ;
        RECT 0.040 200.440 0.360 200.760 ;
        RECT 0.440 200.440 0.760 200.760 ;
        RECT 0.840 200.440 1.160 200.760 ;
        RECT 1.240 200.440 1.560 200.760 ;
        RECT 1.640 200.440 1.960 200.760 ;
        RECT 2.040 200.440 2.360 200.760 ;
        RECT 2.440 200.440 2.760 200.760 ;
        RECT 2.840 200.440 3.160 200.760 ;
        RECT 3.240 200.440 3.560 200.760 ;
        RECT 3.640 200.440 3.960 200.760 ;
        RECT 4.040 200.440 4.360 200.760 ;
        RECT 4.440 200.440 4.760 200.760 ;
        RECT 4.840 200.440 5.160 200.760 ;
        RECT 5.240 200.440 5.560 200.760 ;
        RECT 5.640 200.440 5.960 200.760 ;
        RECT 6.040 200.440 6.360 200.760 ;
        RECT 6.440 200.440 6.760 200.760 ;
        RECT 6.840 200.440 7.160 200.760 ;
        RECT 7.240 200.440 7.560 200.760 ;
        RECT 7.640 200.440 7.960 200.760 ;
        RECT 8.040 200.440 8.360 200.760 ;
        RECT 8.440 200.440 8.760 200.760 ;
        RECT 8.840 200.440 9.160 200.760 ;
        RECT 9.240 200.440 9.560 200.760 ;
        RECT 9.640 200.440 9.960 200.760 ;
        RECT 10.040 200.440 10.360 200.760 ;
        RECT 10.440 200.440 10.760 200.760 ;
        RECT 10.840 200.440 11.160 200.760 ;
        RECT 11.240 200.440 11.560 200.760 ;
        RECT 11.640 200.440 11.960 200.760 ;
        RECT 12.040 200.440 12.360 200.760 ;
        RECT 12.440 200.440 12.760 200.760 ;
        RECT 12.840 200.440 13.160 200.760 ;
        RECT 13.240 200.440 13.560 200.760 ;
        RECT 13.640 200.440 13.960 200.760 ;
        RECT 14.040 200.440 14.360 200.760 ;
        RECT 14.440 200.440 14.760 200.760 ;
        RECT 14.840 200.440 15.160 200.760 ;
        RECT 15.240 200.440 15.560 200.760 ;
        RECT 15.640 200.440 15.960 200.760 ;
        RECT 16.040 200.440 16.360 200.760 ;
        RECT 16.440 200.440 16.760 200.760 ;
        RECT 16.840 200.440 17.160 200.760 ;
        RECT 17.240 200.440 17.560 200.760 ;
        RECT 17.640 200.440 17.960 200.760 ;
        RECT 18.040 200.440 18.360 200.760 ;
        RECT 18.440 200.440 18.760 200.760 ;
        RECT 18.840 200.440 19.160 200.760 ;
        RECT 19.240 200.440 19.560 200.760 ;
        RECT 19.640 200.440 19.960 200.760 ;
        RECT 95.560 200.440 95.880 200.760 ;
        RECT 95.960 200.440 96.280 200.760 ;
        RECT 96.360 200.440 96.680 200.760 ;
        RECT 96.760 200.440 97.080 200.760 ;
        RECT 145.560 200.440 145.880 200.760 ;
        RECT 145.960 200.440 146.280 200.760 ;
        RECT 146.360 200.440 146.680 200.760 ;
        RECT 146.760 200.440 147.080 200.760 ;
        RECT 185.720 200.440 186.040 200.760 ;
        RECT 186.120 200.440 186.440 200.760 ;
        RECT 186.520 200.440 186.840 200.760 ;
        RECT 186.920 200.440 187.240 200.760 ;
        RECT 187.320 200.440 187.640 200.760 ;
        RECT 187.720 200.440 188.040 200.760 ;
        RECT 188.120 200.440 188.440 200.760 ;
        RECT 188.520 200.440 188.840 200.760 ;
        RECT 188.920 200.440 189.240 200.760 ;
        RECT 189.320 200.440 189.640 200.760 ;
        RECT 189.720 200.440 190.040 200.760 ;
        RECT 190.120 200.440 190.440 200.760 ;
        RECT 190.520 200.440 190.840 200.760 ;
        RECT 190.920 200.440 191.240 200.760 ;
        RECT 191.320 200.440 191.640 200.760 ;
        RECT 191.720 200.440 192.040 200.760 ;
        RECT 192.120 200.440 192.440 200.760 ;
        RECT 192.520 200.440 192.840 200.760 ;
        RECT 192.920 200.440 193.240 200.760 ;
        RECT 193.320 200.440 193.640 200.760 ;
        RECT 193.720 200.440 194.040 200.760 ;
        RECT 194.120 200.440 194.440 200.760 ;
        RECT 194.520 200.440 194.840 200.760 ;
        RECT 194.920 200.440 195.240 200.760 ;
        RECT 195.320 200.440 195.640 200.760 ;
        RECT 195.720 200.440 196.040 200.760 ;
        RECT 196.120 200.440 196.440 200.760 ;
        RECT 196.520 200.440 196.840 200.760 ;
        RECT 196.920 200.440 197.240 200.760 ;
        RECT 197.320 200.440 197.640 200.760 ;
        RECT 197.720 200.440 198.040 200.760 ;
        RECT 198.120 200.440 198.440 200.760 ;
        RECT 198.520 200.440 198.840 200.760 ;
        RECT 198.920 200.440 199.240 200.760 ;
        RECT 199.320 200.440 199.640 200.760 ;
        RECT 199.720 200.440 200.040 200.760 ;
        RECT 200.120 200.440 200.440 200.760 ;
        RECT 200.520 200.440 200.840 200.760 ;
        RECT 200.920 200.440 201.240 200.760 ;
        RECT 201.320 200.440 201.640 200.760 ;
        RECT 201.720 200.440 202.040 200.760 ;
        RECT 202.120 200.440 202.440 200.760 ;
        RECT 202.520 200.440 202.840 200.760 ;
        RECT 202.920 200.440 203.240 200.760 ;
        RECT 203.320 200.440 203.640 200.760 ;
        RECT 203.720 200.440 204.040 200.760 ;
        RECT 204.120 200.440 204.440 200.760 ;
        RECT 204.520 200.440 204.840 200.760 ;
        RECT 204.920 200.440 205.240 200.760 ;
        RECT 205.320 200.440 205.640 200.760 ;
        RECT 0.040 200.040 0.360 200.360 ;
        RECT 0.440 200.040 0.760 200.360 ;
        RECT 0.840 200.040 1.160 200.360 ;
        RECT 1.240 200.040 1.560 200.360 ;
        RECT 1.640 200.040 1.960 200.360 ;
        RECT 2.040 200.040 2.360 200.360 ;
        RECT 2.440 200.040 2.760 200.360 ;
        RECT 2.840 200.040 3.160 200.360 ;
        RECT 3.240 200.040 3.560 200.360 ;
        RECT 3.640 200.040 3.960 200.360 ;
        RECT 4.040 200.040 4.360 200.360 ;
        RECT 4.440 200.040 4.760 200.360 ;
        RECT 4.840 200.040 5.160 200.360 ;
        RECT 5.240 200.040 5.560 200.360 ;
        RECT 5.640 200.040 5.960 200.360 ;
        RECT 6.040 200.040 6.360 200.360 ;
        RECT 6.440 200.040 6.760 200.360 ;
        RECT 6.840 200.040 7.160 200.360 ;
        RECT 7.240 200.040 7.560 200.360 ;
        RECT 7.640 200.040 7.960 200.360 ;
        RECT 8.040 200.040 8.360 200.360 ;
        RECT 8.440 200.040 8.760 200.360 ;
        RECT 8.840 200.040 9.160 200.360 ;
        RECT 9.240 200.040 9.560 200.360 ;
        RECT 9.640 200.040 9.960 200.360 ;
        RECT 10.040 200.040 10.360 200.360 ;
        RECT 10.440 200.040 10.760 200.360 ;
        RECT 10.840 200.040 11.160 200.360 ;
        RECT 11.240 200.040 11.560 200.360 ;
        RECT 11.640 200.040 11.960 200.360 ;
        RECT 12.040 200.040 12.360 200.360 ;
        RECT 12.440 200.040 12.760 200.360 ;
        RECT 12.840 200.040 13.160 200.360 ;
        RECT 13.240 200.040 13.560 200.360 ;
        RECT 13.640 200.040 13.960 200.360 ;
        RECT 14.040 200.040 14.360 200.360 ;
        RECT 14.440 200.040 14.760 200.360 ;
        RECT 14.840 200.040 15.160 200.360 ;
        RECT 15.240 200.040 15.560 200.360 ;
        RECT 15.640 200.040 15.960 200.360 ;
        RECT 16.040 200.040 16.360 200.360 ;
        RECT 16.440 200.040 16.760 200.360 ;
        RECT 16.840 200.040 17.160 200.360 ;
        RECT 17.240 200.040 17.560 200.360 ;
        RECT 17.640 200.040 17.960 200.360 ;
        RECT 18.040 200.040 18.360 200.360 ;
        RECT 18.440 200.040 18.760 200.360 ;
        RECT 18.840 200.040 19.160 200.360 ;
        RECT 19.240 200.040 19.560 200.360 ;
        RECT 19.640 200.040 19.960 200.360 ;
        RECT 95.560 200.040 95.880 200.360 ;
        RECT 95.960 200.040 96.280 200.360 ;
        RECT 96.360 200.040 96.680 200.360 ;
        RECT 96.760 200.040 97.080 200.360 ;
        RECT 145.560 200.040 145.880 200.360 ;
        RECT 145.960 200.040 146.280 200.360 ;
        RECT 146.360 200.040 146.680 200.360 ;
        RECT 146.760 200.040 147.080 200.360 ;
        RECT 185.720 200.040 186.040 200.360 ;
        RECT 186.120 200.040 186.440 200.360 ;
        RECT 186.520 200.040 186.840 200.360 ;
        RECT 186.920 200.040 187.240 200.360 ;
        RECT 187.320 200.040 187.640 200.360 ;
        RECT 187.720 200.040 188.040 200.360 ;
        RECT 188.120 200.040 188.440 200.360 ;
        RECT 188.520 200.040 188.840 200.360 ;
        RECT 188.920 200.040 189.240 200.360 ;
        RECT 189.320 200.040 189.640 200.360 ;
        RECT 189.720 200.040 190.040 200.360 ;
        RECT 190.120 200.040 190.440 200.360 ;
        RECT 190.520 200.040 190.840 200.360 ;
        RECT 190.920 200.040 191.240 200.360 ;
        RECT 191.320 200.040 191.640 200.360 ;
        RECT 191.720 200.040 192.040 200.360 ;
        RECT 192.120 200.040 192.440 200.360 ;
        RECT 192.520 200.040 192.840 200.360 ;
        RECT 192.920 200.040 193.240 200.360 ;
        RECT 193.320 200.040 193.640 200.360 ;
        RECT 193.720 200.040 194.040 200.360 ;
        RECT 194.120 200.040 194.440 200.360 ;
        RECT 194.520 200.040 194.840 200.360 ;
        RECT 194.920 200.040 195.240 200.360 ;
        RECT 195.320 200.040 195.640 200.360 ;
        RECT 195.720 200.040 196.040 200.360 ;
        RECT 196.120 200.040 196.440 200.360 ;
        RECT 196.520 200.040 196.840 200.360 ;
        RECT 196.920 200.040 197.240 200.360 ;
        RECT 197.320 200.040 197.640 200.360 ;
        RECT 197.720 200.040 198.040 200.360 ;
        RECT 198.120 200.040 198.440 200.360 ;
        RECT 198.520 200.040 198.840 200.360 ;
        RECT 198.920 200.040 199.240 200.360 ;
        RECT 199.320 200.040 199.640 200.360 ;
        RECT 199.720 200.040 200.040 200.360 ;
        RECT 200.120 200.040 200.440 200.360 ;
        RECT 200.520 200.040 200.840 200.360 ;
        RECT 200.920 200.040 201.240 200.360 ;
        RECT 201.320 200.040 201.640 200.360 ;
        RECT 201.720 200.040 202.040 200.360 ;
        RECT 202.120 200.040 202.440 200.360 ;
        RECT 202.520 200.040 202.840 200.360 ;
        RECT 202.920 200.040 203.240 200.360 ;
        RECT 203.320 200.040 203.640 200.360 ;
        RECT 203.720 200.040 204.040 200.360 ;
        RECT 204.120 200.040 204.440 200.360 ;
        RECT 204.520 200.040 204.840 200.360 ;
        RECT 204.920 200.040 205.240 200.360 ;
        RECT 205.320 200.040 205.640 200.360 ;
        RECT 0.040 199.640 0.360 199.960 ;
        RECT 0.440 199.640 0.760 199.960 ;
        RECT 0.840 199.640 1.160 199.960 ;
        RECT 1.240 199.640 1.560 199.960 ;
        RECT 1.640 199.640 1.960 199.960 ;
        RECT 2.040 199.640 2.360 199.960 ;
        RECT 2.440 199.640 2.760 199.960 ;
        RECT 2.840 199.640 3.160 199.960 ;
        RECT 3.240 199.640 3.560 199.960 ;
        RECT 3.640 199.640 3.960 199.960 ;
        RECT 4.040 199.640 4.360 199.960 ;
        RECT 4.440 199.640 4.760 199.960 ;
        RECT 4.840 199.640 5.160 199.960 ;
        RECT 5.240 199.640 5.560 199.960 ;
        RECT 5.640 199.640 5.960 199.960 ;
        RECT 6.040 199.640 6.360 199.960 ;
        RECT 6.440 199.640 6.760 199.960 ;
        RECT 6.840 199.640 7.160 199.960 ;
        RECT 7.240 199.640 7.560 199.960 ;
        RECT 7.640 199.640 7.960 199.960 ;
        RECT 8.040 199.640 8.360 199.960 ;
        RECT 8.440 199.640 8.760 199.960 ;
        RECT 8.840 199.640 9.160 199.960 ;
        RECT 9.240 199.640 9.560 199.960 ;
        RECT 9.640 199.640 9.960 199.960 ;
        RECT 10.040 199.640 10.360 199.960 ;
        RECT 10.440 199.640 10.760 199.960 ;
        RECT 10.840 199.640 11.160 199.960 ;
        RECT 11.240 199.640 11.560 199.960 ;
        RECT 11.640 199.640 11.960 199.960 ;
        RECT 12.040 199.640 12.360 199.960 ;
        RECT 12.440 199.640 12.760 199.960 ;
        RECT 12.840 199.640 13.160 199.960 ;
        RECT 13.240 199.640 13.560 199.960 ;
        RECT 13.640 199.640 13.960 199.960 ;
        RECT 14.040 199.640 14.360 199.960 ;
        RECT 14.440 199.640 14.760 199.960 ;
        RECT 14.840 199.640 15.160 199.960 ;
        RECT 15.240 199.640 15.560 199.960 ;
        RECT 15.640 199.640 15.960 199.960 ;
        RECT 16.040 199.640 16.360 199.960 ;
        RECT 16.440 199.640 16.760 199.960 ;
        RECT 16.840 199.640 17.160 199.960 ;
        RECT 17.240 199.640 17.560 199.960 ;
        RECT 17.640 199.640 17.960 199.960 ;
        RECT 18.040 199.640 18.360 199.960 ;
        RECT 18.440 199.640 18.760 199.960 ;
        RECT 18.840 199.640 19.160 199.960 ;
        RECT 19.240 199.640 19.560 199.960 ;
        RECT 19.640 199.640 19.960 199.960 ;
        RECT 95.560 199.640 95.880 199.960 ;
        RECT 95.960 199.640 96.280 199.960 ;
        RECT 96.360 199.640 96.680 199.960 ;
        RECT 96.760 199.640 97.080 199.960 ;
        RECT 145.560 199.640 145.880 199.960 ;
        RECT 145.960 199.640 146.280 199.960 ;
        RECT 146.360 199.640 146.680 199.960 ;
        RECT 146.760 199.640 147.080 199.960 ;
        RECT 185.720 199.640 186.040 199.960 ;
        RECT 186.120 199.640 186.440 199.960 ;
        RECT 186.520 199.640 186.840 199.960 ;
        RECT 186.920 199.640 187.240 199.960 ;
        RECT 187.320 199.640 187.640 199.960 ;
        RECT 187.720 199.640 188.040 199.960 ;
        RECT 188.120 199.640 188.440 199.960 ;
        RECT 188.520 199.640 188.840 199.960 ;
        RECT 188.920 199.640 189.240 199.960 ;
        RECT 189.320 199.640 189.640 199.960 ;
        RECT 189.720 199.640 190.040 199.960 ;
        RECT 190.120 199.640 190.440 199.960 ;
        RECT 190.520 199.640 190.840 199.960 ;
        RECT 190.920 199.640 191.240 199.960 ;
        RECT 191.320 199.640 191.640 199.960 ;
        RECT 191.720 199.640 192.040 199.960 ;
        RECT 192.120 199.640 192.440 199.960 ;
        RECT 192.520 199.640 192.840 199.960 ;
        RECT 192.920 199.640 193.240 199.960 ;
        RECT 193.320 199.640 193.640 199.960 ;
        RECT 193.720 199.640 194.040 199.960 ;
        RECT 194.120 199.640 194.440 199.960 ;
        RECT 194.520 199.640 194.840 199.960 ;
        RECT 194.920 199.640 195.240 199.960 ;
        RECT 195.320 199.640 195.640 199.960 ;
        RECT 195.720 199.640 196.040 199.960 ;
        RECT 196.120 199.640 196.440 199.960 ;
        RECT 196.520 199.640 196.840 199.960 ;
        RECT 196.920 199.640 197.240 199.960 ;
        RECT 197.320 199.640 197.640 199.960 ;
        RECT 197.720 199.640 198.040 199.960 ;
        RECT 198.120 199.640 198.440 199.960 ;
        RECT 198.520 199.640 198.840 199.960 ;
        RECT 198.920 199.640 199.240 199.960 ;
        RECT 199.320 199.640 199.640 199.960 ;
        RECT 199.720 199.640 200.040 199.960 ;
        RECT 200.120 199.640 200.440 199.960 ;
        RECT 200.520 199.640 200.840 199.960 ;
        RECT 200.920 199.640 201.240 199.960 ;
        RECT 201.320 199.640 201.640 199.960 ;
        RECT 201.720 199.640 202.040 199.960 ;
        RECT 202.120 199.640 202.440 199.960 ;
        RECT 202.520 199.640 202.840 199.960 ;
        RECT 202.920 199.640 203.240 199.960 ;
        RECT 203.320 199.640 203.640 199.960 ;
        RECT 203.720 199.640 204.040 199.960 ;
        RECT 204.120 199.640 204.440 199.960 ;
        RECT 204.520 199.640 204.840 199.960 ;
        RECT 204.920 199.640 205.240 199.960 ;
        RECT 205.320 199.640 205.640 199.960 ;
        RECT 0.040 199.240 0.360 199.560 ;
        RECT 0.440 199.240 0.760 199.560 ;
        RECT 0.840 199.240 1.160 199.560 ;
        RECT 1.240 199.240 1.560 199.560 ;
        RECT 1.640 199.240 1.960 199.560 ;
        RECT 2.040 199.240 2.360 199.560 ;
        RECT 2.440 199.240 2.760 199.560 ;
        RECT 2.840 199.240 3.160 199.560 ;
        RECT 3.240 199.240 3.560 199.560 ;
        RECT 3.640 199.240 3.960 199.560 ;
        RECT 4.040 199.240 4.360 199.560 ;
        RECT 4.440 199.240 4.760 199.560 ;
        RECT 4.840 199.240 5.160 199.560 ;
        RECT 5.240 199.240 5.560 199.560 ;
        RECT 5.640 199.240 5.960 199.560 ;
        RECT 6.040 199.240 6.360 199.560 ;
        RECT 6.440 199.240 6.760 199.560 ;
        RECT 6.840 199.240 7.160 199.560 ;
        RECT 7.240 199.240 7.560 199.560 ;
        RECT 7.640 199.240 7.960 199.560 ;
        RECT 8.040 199.240 8.360 199.560 ;
        RECT 8.440 199.240 8.760 199.560 ;
        RECT 8.840 199.240 9.160 199.560 ;
        RECT 9.240 199.240 9.560 199.560 ;
        RECT 9.640 199.240 9.960 199.560 ;
        RECT 10.040 199.240 10.360 199.560 ;
        RECT 10.440 199.240 10.760 199.560 ;
        RECT 10.840 199.240 11.160 199.560 ;
        RECT 11.240 199.240 11.560 199.560 ;
        RECT 11.640 199.240 11.960 199.560 ;
        RECT 12.040 199.240 12.360 199.560 ;
        RECT 12.440 199.240 12.760 199.560 ;
        RECT 12.840 199.240 13.160 199.560 ;
        RECT 13.240 199.240 13.560 199.560 ;
        RECT 13.640 199.240 13.960 199.560 ;
        RECT 14.040 199.240 14.360 199.560 ;
        RECT 14.440 199.240 14.760 199.560 ;
        RECT 14.840 199.240 15.160 199.560 ;
        RECT 15.240 199.240 15.560 199.560 ;
        RECT 15.640 199.240 15.960 199.560 ;
        RECT 16.040 199.240 16.360 199.560 ;
        RECT 16.440 199.240 16.760 199.560 ;
        RECT 16.840 199.240 17.160 199.560 ;
        RECT 17.240 199.240 17.560 199.560 ;
        RECT 17.640 199.240 17.960 199.560 ;
        RECT 18.040 199.240 18.360 199.560 ;
        RECT 18.440 199.240 18.760 199.560 ;
        RECT 18.840 199.240 19.160 199.560 ;
        RECT 19.240 199.240 19.560 199.560 ;
        RECT 19.640 199.240 19.960 199.560 ;
        RECT 95.560 199.240 95.880 199.560 ;
        RECT 95.960 199.240 96.280 199.560 ;
        RECT 96.360 199.240 96.680 199.560 ;
        RECT 96.760 199.240 97.080 199.560 ;
        RECT 145.560 199.240 145.880 199.560 ;
        RECT 145.960 199.240 146.280 199.560 ;
        RECT 146.360 199.240 146.680 199.560 ;
        RECT 146.760 199.240 147.080 199.560 ;
        RECT 185.720 199.240 186.040 199.560 ;
        RECT 186.120 199.240 186.440 199.560 ;
        RECT 186.520 199.240 186.840 199.560 ;
        RECT 186.920 199.240 187.240 199.560 ;
        RECT 187.320 199.240 187.640 199.560 ;
        RECT 187.720 199.240 188.040 199.560 ;
        RECT 188.120 199.240 188.440 199.560 ;
        RECT 188.520 199.240 188.840 199.560 ;
        RECT 188.920 199.240 189.240 199.560 ;
        RECT 189.320 199.240 189.640 199.560 ;
        RECT 189.720 199.240 190.040 199.560 ;
        RECT 190.120 199.240 190.440 199.560 ;
        RECT 190.520 199.240 190.840 199.560 ;
        RECT 190.920 199.240 191.240 199.560 ;
        RECT 191.320 199.240 191.640 199.560 ;
        RECT 191.720 199.240 192.040 199.560 ;
        RECT 192.120 199.240 192.440 199.560 ;
        RECT 192.520 199.240 192.840 199.560 ;
        RECT 192.920 199.240 193.240 199.560 ;
        RECT 193.320 199.240 193.640 199.560 ;
        RECT 193.720 199.240 194.040 199.560 ;
        RECT 194.120 199.240 194.440 199.560 ;
        RECT 194.520 199.240 194.840 199.560 ;
        RECT 194.920 199.240 195.240 199.560 ;
        RECT 195.320 199.240 195.640 199.560 ;
        RECT 195.720 199.240 196.040 199.560 ;
        RECT 196.120 199.240 196.440 199.560 ;
        RECT 196.520 199.240 196.840 199.560 ;
        RECT 196.920 199.240 197.240 199.560 ;
        RECT 197.320 199.240 197.640 199.560 ;
        RECT 197.720 199.240 198.040 199.560 ;
        RECT 198.120 199.240 198.440 199.560 ;
        RECT 198.520 199.240 198.840 199.560 ;
        RECT 198.920 199.240 199.240 199.560 ;
        RECT 199.320 199.240 199.640 199.560 ;
        RECT 199.720 199.240 200.040 199.560 ;
        RECT 200.120 199.240 200.440 199.560 ;
        RECT 200.520 199.240 200.840 199.560 ;
        RECT 200.920 199.240 201.240 199.560 ;
        RECT 201.320 199.240 201.640 199.560 ;
        RECT 201.720 199.240 202.040 199.560 ;
        RECT 202.120 199.240 202.440 199.560 ;
        RECT 202.520 199.240 202.840 199.560 ;
        RECT 202.920 199.240 203.240 199.560 ;
        RECT 203.320 199.240 203.640 199.560 ;
        RECT 203.720 199.240 204.040 199.560 ;
        RECT 204.120 199.240 204.440 199.560 ;
        RECT 204.520 199.240 204.840 199.560 ;
        RECT 204.920 199.240 205.240 199.560 ;
        RECT 205.320 199.240 205.640 199.560 ;
        RECT 0.040 198.840 0.360 199.160 ;
        RECT 0.440 198.840 0.760 199.160 ;
        RECT 0.840 198.840 1.160 199.160 ;
        RECT 1.240 198.840 1.560 199.160 ;
        RECT 1.640 198.840 1.960 199.160 ;
        RECT 2.040 198.840 2.360 199.160 ;
        RECT 2.440 198.840 2.760 199.160 ;
        RECT 2.840 198.840 3.160 199.160 ;
        RECT 3.240 198.840 3.560 199.160 ;
        RECT 3.640 198.840 3.960 199.160 ;
        RECT 4.040 198.840 4.360 199.160 ;
        RECT 4.440 198.840 4.760 199.160 ;
        RECT 4.840 198.840 5.160 199.160 ;
        RECT 5.240 198.840 5.560 199.160 ;
        RECT 5.640 198.840 5.960 199.160 ;
        RECT 6.040 198.840 6.360 199.160 ;
        RECT 6.440 198.840 6.760 199.160 ;
        RECT 6.840 198.840 7.160 199.160 ;
        RECT 7.240 198.840 7.560 199.160 ;
        RECT 7.640 198.840 7.960 199.160 ;
        RECT 8.040 198.840 8.360 199.160 ;
        RECT 8.440 198.840 8.760 199.160 ;
        RECT 8.840 198.840 9.160 199.160 ;
        RECT 9.240 198.840 9.560 199.160 ;
        RECT 9.640 198.840 9.960 199.160 ;
        RECT 10.040 198.840 10.360 199.160 ;
        RECT 10.440 198.840 10.760 199.160 ;
        RECT 10.840 198.840 11.160 199.160 ;
        RECT 11.240 198.840 11.560 199.160 ;
        RECT 11.640 198.840 11.960 199.160 ;
        RECT 12.040 198.840 12.360 199.160 ;
        RECT 12.440 198.840 12.760 199.160 ;
        RECT 12.840 198.840 13.160 199.160 ;
        RECT 13.240 198.840 13.560 199.160 ;
        RECT 13.640 198.840 13.960 199.160 ;
        RECT 14.040 198.840 14.360 199.160 ;
        RECT 14.440 198.840 14.760 199.160 ;
        RECT 14.840 198.840 15.160 199.160 ;
        RECT 15.240 198.840 15.560 199.160 ;
        RECT 15.640 198.840 15.960 199.160 ;
        RECT 16.040 198.840 16.360 199.160 ;
        RECT 16.440 198.840 16.760 199.160 ;
        RECT 16.840 198.840 17.160 199.160 ;
        RECT 17.240 198.840 17.560 199.160 ;
        RECT 17.640 198.840 17.960 199.160 ;
        RECT 18.040 198.840 18.360 199.160 ;
        RECT 18.440 198.840 18.760 199.160 ;
        RECT 18.840 198.840 19.160 199.160 ;
        RECT 19.240 198.840 19.560 199.160 ;
        RECT 19.640 198.840 19.960 199.160 ;
        RECT 95.560 198.840 95.880 199.160 ;
        RECT 95.960 198.840 96.280 199.160 ;
        RECT 96.360 198.840 96.680 199.160 ;
        RECT 96.760 198.840 97.080 199.160 ;
        RECT 145.560 198.840 145.880 199.160 ;
        RECT 145.960 198.840 146.280 199.160 ;
        RECT 146.360 198.840 146.680 199.160 ;
        RECT 146.760 198.840 147.080 199.160 ;
        RECT 185.720 198.840 186.040 199.160 ;
        RECT 186.120 198.840 186.440 199.160 ;
        RECT 186.520 198.840 186.840 199.160 ;
        RECT 186.920 198.840 187.240 199.160 ;
        RECT 187.320 198.840 187.640 199.160 ;
        RECT 187.720 198.840 188.040 199.160 ;
        RECT 188.120 198.840 188.440 199.160 ;
        RECT 188.520 198.840 188.840 199.160 ;
        RECT 188.920 198.840 189.240 199.160 ;
        RECT 189.320 198.840 189.640 199.160 ;
        RECT 189.720 198.840 190.040 199.160 ;
        RECT 190.120 198.840 190.440 199.160 ;
        RECT 190.520 198.840 190.840 199.160 ;
        RECT 190.920 198.840 191.240 199.160 ;
        RECT 191.320 198.840 191.640 199.160 ;
        RECT 191.720 198.840 192.040 199.160 ;
        RECT 192.120 198.840 192.440 199.160 ;
        RECT 192.520 198.840 192.840 199.160 ;
        RECT 192.920 198.840 193.240 199.160 ;
        RECT 193.320 198.840 193.640 199.160 ;
        RECT 193.720 198.840 194.040 199.160 ;
        RECT 194.120 198.840 194.440 199.160 ;
        RECT 194.520 198.840 194.840 199.160 ;
        RECT 194.920 198.840 195.240 199.160 ;
        RECT 195.320 198.840 195.640 199.160 ;
        RECT 195.720 198.840 196.040 199.160 ;
        RECT 196.120 198.840 196.440 199.160 ;
        RECT 196.520 198.840 196.840 199.160 ;
        RECT 196.920 198.840 197.240 199.160 ;
        RECT 197.320 198.840 197.640 199.160 ;
        RECT 197.720 198.840 198.040 199.160 ;
        RECT 198.120 198.840 198.440 199.160 ;
        RECT 198.520 198.840 198.840 199.160 ;
        RECT 198.920 198.840 199.240 199.160 ;
        RECT 199.320 198.840 199.640 199.160 ;
        RECT 199.720 198.840 200.040 199.160 ;
        RECT 200.120 198.840 200.440 199.160 ;
        RECT 200.520 198.840 200.840 199.160 ;
        RECT 200.920 198.840 201.240 199.160 ;
        RECT 201.320 198.840 201.640 199.160 ;
        RECT 201.720 198.840 202.040 199.160 ;
        RECT 202.120 198.840 202.440 199.160 ;
        RECT 202.520 198.840 202.840 199.160 ;
        RECT 202.920 198.840 203.240 199.160 ;
        RECT 203.320 198.840 203.640 199.160 ;
        RECT 203.720 198.840 204.040 199.160 ;
        RECT 204.120 198.840 204.440 199.160 ;
        RECT 204.520 198.840 204.840 199.160 ;
        RECT 204.920 198.840 205.240 199.160 ;
        RECT 205.320 198.840 205.640 199.160 ;
        RECT 0.040 198.440 0.360 198.760 ;
        RECT 0.440 198.440 0.760 198.760 ;
        RECT 0.840 198.440 1.160 198.760 ;
        RECT 1.240 198.440 1.560 198.760 ;
        RECT 1.640 198.440 1.960 198.760 ;
        RECT 2.040 198.440 2.360 198.760 ;
        RECT 2.440 198.440 2.760 198.760 ;
        RECT 2.840 198.440 3.160 198.760 ;
        RECT 3.240 198.440 3.560 198.760 ;
        RECT 3.640 198.440 3.960 198.760 ;
        RECT 4.040 198.440 4.360 198.760 ;
        RECT 4.440 198.440 4.760 198.760 ;
        RECT 4.840 198.440 5.160 198.760 ;
        RECT 5.240 198.440 5.560 198.760 ;
        RECT 5.640 198.440 5.960 198.760 ;
        RECT 6.040 198.440 6.360 198.760 ;
        RECT 6.440 198.440 6.760 198.760 ;
        RECT 6.840 198.440 7.160 198.760 ;
        RECT 7.240 198.440 7.560 198.760 ;
        RECT 7.640 198.440 7.960 198.760 ;
        RECT 8.040 198.440 8.360 198.760 ;
        RECT 8.440 198.440 8.760 198.760 ;
        RECT 8.840 198.440 9.160 198.760 ;
        RECT 9.240 198.440 9.560 198.760 ;
        RECT 9.640 198.440 9.960 198.760 ;
        RECT 10.040 198.440 10.360 198.760 ;
        RECT 10.440 198.440 10.760 198.760 ;
        RECT 10.840 198.440 11.160 198.760 ;
        RECT 11.240 198.440 11.560 198.760 ;
        RECT 11.640 198.440 11.960 198.760 ;
        RECT 12.040 198.440 12.360 198.760 ;
        RECT 12.440 198.440 12.760 198.760 ;
        RECT 12.840 198.440 13.160 198.760 ;
        RECT 13.240 198.440 13.560 198.760 ;
        RECT 13.640 198.440 13.960 198.760 ;
        RECT 14.040 198.440 14.360 198.760 ;
        RECT 14.440 198.440 14.760 198.760 ;
        RECT 14.840 198.440 15.160 198.760 ;
        RECT 15.240 198.440 15.560 198.760 ;
        RECT 15.640 198.440 15.960 198.760 ;
        RECT 16.040 198.440 16.360 198.760 ;
        RECT 16.440 198.440 16.760 198.760 ;
        RECT 16.840 198.440 17.160 198.760 ;
        RECT 17.240 198.440 17.560 198.760 ;
        RECT 17.640 198.440 17.960 198.760 ;
        RECT 18.040 198.440 18.360 198.760 ;
        RECT 18.440 198.440 18.760 198.760 ;
        RECT 18.840 198.440 19.160 198.760 ;
        RECT 19.240 198.440 19.560 198.760 ;
        RECT 19.640 198.440 19.960 198.760 ;
        RECT 95.560 198.440 95.880 198.760 ;
        RECT 95.960 198.440 96.280 198.760 ;
        RECT 96.360 198.440 96.680 198.760 ;
        RECT 96.760 198.440 97.080 198.760 ;
        RECT 145.560 198.440 145.880 198.760 ;
        RECT 145.960 198.440 146.280 198.760 ;
        RECT 146.360 198.440 146.680 198.760 ;
        RECT 146.760 198.440 147.080 198.760 ;
        RECT 185.720 198.440 186.040 198.760 ;
        RECT 186.120 198.440 186.440 198.760 ;
        RECT 186.520 198.440 186.840 198.760 ;
        RECT 186.920 198.440 187.240 198.760 ;
        RECT 187.320 198.440 187.640 198.760 ;
        RECT 187.720 198.440 188.040 198.760 ;
        RECT 188.120 198.440 188.440 198.760 ;
        RECT 188.520 198.440 188.840 198.760 ;
        RECT 188.920 198.440 189.240 198.760 ;
        RECT 189.320 198.440 189.640 198.760 ;
        RECT 189.720 198.440 190.040 198.760 ;
        RECT 190.120 198.440 190.440 198.760 ;
        RECT 190.520 198.440 190.840 198.760 ;
        RECT 190.920 198.440 191.240 198.760 ;
        RECT 191.320 198.440 191.640 198.760 ;
        RECT 191.720 198.440 192.040 198.760 ;
        RECT 192.120 198.440 192.440 198.760 ;
        RECT 192.520 198.440 192.840 198.760 ;
        RECT 192.920 198.440 193.240 198.760 ;
        RECT 193.320 198.440 193.640 198.760 ;
        RECT 193.720 198.440 194.040 198.760 ;
        RECT 194.120 198.440 194.440 198.760 ;
        RECT 194.520 198.440 194.840 198.760 ;
        RECT 194.920 198.440 195.240 198.760 ;
        RECT 195.320 198.440 195.640 198.760 ;
        RECT 195.720 198.440 196.040 198.760 ;
        RECT 196.120 198.440 196.440 198.760 ;
        RECT 196.520 198.440 196.840 198.760 ;
        RECT 196.920 198.440 197.240 198.760 ;
        RECT 197.320 198.440 197.640 198.760 ;
        RECT 197.720 198.440 198.040 198.760 ;
        RECT 198.120 198.440 198.440 198.760 ;
        RECT 198.520 198.440 198.840 198.760 ;
        RECT 198.920 198.440 199.240 198.760 ;
        RECT 199.320 198.440 199.640 198.760 ;
        RECT 199.720 198.440 200.040 198.760 ;
        RECT 200.120 198.440 200.440 198.760 ;
        RECT 200.520 198.440 200.840 198.760 ;
        RECT 200.920 198.440 201.240 198.760 ;
        RECT 201.320 198.440 201.640 198.760 ;
        RECT 201.720 198.440 202.040 198.760 ;
        RECT 202.120 198.440 202.440 198.760 ;
        RECT 202.520 198.440 202.840 198.760 ;
        RECT 202.920 198.440 203.240 198.760 ;
        RECT 203.320 198.440 203.640 198.760 ;
        RECT 203.720 198.440 204.040 198.760 ;
        RECT 204.120 198.440 204.440 198.760 ;
        RECT 204.520 198.440 204.840 198.760 ;
        RECT 204.920 198.440 205.240 198.760 ;
        RECT 205.320 198.440 205.640 198.760 ;
        RECT 0.040 198.040 0.360 198.360 ;
        RECT 0.440 198.040 0.760 198.360 ;
        RECT 0.840 198.040 1.160 198.360 ;
        RECT 1.240 198.040 1.560 198.360 ;
        RECT 1.640 198.040 1.960 198.360 ;
        RECT 2.040 198.040 2.360 198.360 ;
        RECT 2.440 198.040 2.760 198.360 ;
        RECT 2.840 198.040 3.160 198.360 ;
        RECT 3.240 198.040 3.560 198.360 ;
        RECT 3.640 198.040 3.960 198.360 ;
        RECT 4.040 198.040 4.360 198.360 ;
        RECT 4.440 198.040 4.760 198.360 ;
        RECT 4.840 198.040 5.160 198.360 ;
        RECT 5.240 198.040 5.560 198.360 ;
        RECT 5.640 198.040 5.960 198.360 ;
        RECT 6.040 198.040 6.360 198.360 ;
        RECT 6.440 198.040 6.760 198.360 ;
        RECT 6.840 198.040 7.160 198.360 ;
        RECT 7.240 198.040 7.560 198.360 ;
        RECT 7.640 198.040 7.960 198.360 ;
        RECT 8.040 198.040 8.360 198.360 ;
        RECT 8.440 198.040 8.760 198.360 ;
        RECT 8.840 198.040 9.160 198.360 ;
        RECT 9.240 198.040 9.560 198.360 ;
        RECT 9.640 198.040 9.960 198.360 ;
        RECT 10.040 198.040 10.360 198.360 ;
        RECT 10.440 198.040 10.760 198.360 ;
        RECT 10.840 198.040 11.160 198.360 ;
        RECT 11.240 198.040 11.560 198.360 ;
        RECT 11.640 198.040 11.960 198.360 ;
        RECT 12.040 198.040 12.360 198.360 ;
        RECT 12.440 198.040 12.760 198.360 ;
        RECT 12.840 198.040 13.160 198.360 ;
        RECT 13.240 198.040 13.560 198.360 ;
        RECT 13.640 198.040 13.960 198.360 ;
        RECT 14.040 198.040 14.360 198.360 ;
        RECT 14.440 198.040 14.760 198.360 ;
        RECT 14.840 198.040 15.160 198.360 ;
        RECT 15.240 198.040 15.560 198.360 ;
        RECT 15.640 198.040 15.960 198.360 ;
        RECT 16.040 198.040 16.360 198.360 ;
        RECT 16.440 198.040 16.760 198.360 ;
        RECT 16.840 198.040 17.160 198.360 ;
        RECT 17.240 198.040 17.560 198.360 ;
        RECT 17.640 198.040 17.960 198.360 ;
        RECT 18.040 198.040 18.360 198.360 ;
        RECT 18.440 198.040 18.760 198.360 ;
        RECT 18.840 198.040 19.160 198.360 ;
        RECT 19.240 198.040 19.560 198.360 ;
        RECT 19.640 198.040 19.960 198.360 ;
        RECT 95.560 198.040 95.880 198.360 ;
        RECT 95.960 198.040 96.280 198.360 ;
        RECT 96.360 198.040 96.680 198.360 ;
        RECT 96.760 198.040 97.080 198.360 ;
        RECT 145.560 198.040 145.880 198.360 ;
        RECT 145.960 198.040 146.280 198.360 ;
        RECT 146.360 198.040 146.680 198.360 ;
        RECT 146.760 198.040 147.080 198.360 ;
        RECT 185.720 198.040 186.040 198.360 ;
        RECT 186.120 198.040 186.440 198.360 ;
        RECT 186.520 198.040 186.840 198.360 ;
        RECT 186.920 198.040 187.240 198.360 ;
        RECT 187.320 198.040 187.640 198.360 ;
        RECT 187.720 198.040 188.040 198.360 ;
        RECT 188.120 198.040 188.440 198.360 ;
        RECT 188.520 198.040 188.840 198.360 ;
        RECT 188.920 198.040 189.240 198.360 ;
        RECT 189.320 198.040 189.640 198.360 ;
        RECT 189.720 198.040 190.040 198.360 ;
        RECT 190.120 198.040 190.440 198.360 ;
        RECT 190.520 198.040 190.840 198.360 ;
        RECT 190.920 198.040 191.240 198.360 ;
        RECT 191.320 198.040 191.640 198.360 ;
        RECT 191.720 198.040 192.040 198.360 ;
        RECT 192.120 198.040 192.440 198.360 ;
        RECT 192.520 198.040 192.840 198.360 ;
        RECT 192.920 198.040 193.240 198.360 ;
        RECT 193.320 198.040 193.640 198.360 ;
        RECT 193.720 198.040 194.040 198.360 ;
        RECT 194.120 198.040 194.440 198.360 ;
        RECT 194.520 198.040 194.840 198.360 ;
        RECT 194.920 198.040 195.240 198.360 ;
        RECT 195.320 198.040 195.640 198.360 ;
        RECT 195.720 198.040 196.040 198.360 ;
        RECT 196.120 198.040 196.440 198.360 ;
        RECT 196.520 198.040 196.840 198.360 ;
        RECT 196.920 198.040 197.240 198.360 ;
        RECT 197.320 198.040 197.640 198.360 ;
        RECT 197.720 198.040 198.040 198.360 ;
        RECT 198.120 198.040 198.440 198.360 ;
        RECT 198.520 198.040 198.840 198.360 ;
        RECT 198.920 198.040 199.240 198.360 ;
        RECT 199.320 198.040 199.640 198.360 ;
        RECT 199.720 198.040 200.040 198.360 ;
        RECT 200.120 198.040 200.440 198.360 ;
        RECT 200.520 198.040 200.840 198.360 ;
        RECT 200.920 198.040 201.240 198.360 ;
        RECT 201.320 198.040 201.640 198.360 ;
        RECT 201.720 198.040 202.040 198.360 ;
        RECT 202.120 198.040 202.440 198.360 ;
        RECT 202.520 198.040 202.840 198.360 ;
        RECT 202.920 198.040 203.240 198.360 ;
        RECT 203.320 198.040 203.640 198.360 ;
        RECT 203.720 198.040 204.040 198.360 ;
        RECT 204.120 198.040 204.440 198.360 ;
        RECT 204.520 198.040 204.840 198.360 ;
        RECT 204.920 198.040 205.240 198.360 ;
        RECT 205.320 198.040 205.640 198.360 ;
        RECT 0.040 197.640 0.360 197.960 ;
        RECT 0.440 197.640 0.760 197.960 ;
        RECT 0.840 197.640 1.160 197.960 ;
        RECT 1.240 197.640 1.560 197.960 ;
        RECT 1.640 197.640 1.960 197.960 ;
        RECT 2.040 197.640 2.360 197.960 ;
        RECT 2.440 197.640 2.760 197.960 ;
        RECT 2.840 197.640 3.160 197.960 ;
        RECT 3.240 197.640 3.560 197.960 ;
        RECT 3.640 197.640 3.960 197.960 ;
        RECT 4.040 197.640 4.360 197.960 ;
        RECT 4.440 197.640 4.760 197.960 ;
        RECT 4.840 197.640 5.160 197.960 ;
        RECT 5.240 197.640 5.560 197.960 ;
        RECT 5.640 197.640 5.960 197.960 ;
        RECT 6.040 197.640 6.360 197.960 ;
        RECT 6.440 197.640 6.760 197.960 ;
        RECT 6.840 197.640 7.160 197.960 ;
        RECT 7.240 197.640 7.560 197.960 ;
        RECT 7.640 197.640 7.960 197.960 ;
        RECT 8.040 197.640 8.360 197.960 ;
        RECT 8.440 197.640 8.760 197.960 ;
        RECT 8.840 197.640 9.160 197.960 ;
        RECT 9.240 197.640 9.560 197.960 ;
        RECT 9.640 197.640 9.960 197.960 ;
        RECT 10.040 197.640 10.360 197.960 ;
        RECT 10.440 197.640 10.760 197.960 ;
        RECT 10.840 197.640 11.160 197.960 ;
        RECT 11.240 197.640 11.560 197.960 ;
        RECT 11.640 197.640 11.960 197.960 ;
        RECT 12.040 197.640 12.360 197.960 ;
        RECT 12.440 197.640 12.760 197.960 ;
        RECT 12.840 197.640 13.160 197.960 ;
        RECT 13.240 197.640 13.560 197.960 ;
        RECT 13.640 197.640 13.960 197.960 ;
        RECT 14.040 197.640 14.360 197.960 ;
        RECT 14.440 197.640 14.760 197.960 ;
        RECT 14.840 197.640 15.160 197.960 ;
        RECT 15.240 197.640 15.560 197.960 ;
        RECT 15.640 197.640 15.960 197.960 ;
        RECT 16.040 197.640 16.360 197.960 ;
        RECT 16.440 197.640 16.760 197.960 ;
        RECT 16.840 197.640 17.160 197.960 ;
        RECT 17.240 197.640 17.560 197.960 ;
        RECT 17.640 197.640 17.960 197.960 ;
        RECT 18.040 197.640 18.360 197.960 ;
        RECT 18.440 197.640 18.760 197.960 ;
        RECT 18.840 197.640 19.160 197.960 ;
        RECT 19.240 197.640 19.560 197.960 ;
        RECT 19.640 197.640 19.960 197.960 ;
        RECT 95.560 197.640 95.880 197.960 ;
        RECT 95.960 197.640 96.280 197.960 ;
        RECT 96.360 197.640 96.680 197.960 ;
        RECT 96.760 197.640 97.080 197.960 ;
        RECT 145.560 197.640 145.880 197.960 ;
        RECT 145.960 197.640 146.280 197.960 ;
        RECT 146.360 197.640 146.680 197.960 ;
        RECT 146.760 197.640 147.080 197.960 ;
        RECT 185.720 197.640 186.040 197.960 ;
        RECT 186.120 197.640 186.440 197.960 ;
        RECT 186.520 197.640 186.840 197.960 ;
        RECT 186.920 197.640 187.240 197.960 ;
        RECT 187.320 197.640 187.640 197.960 ;
        RECT 187.720 197.640 188.040 197.960 ;
        RECT 188.120 197.640 188.440 197.960 ;
        RECT 188.520 197.640 188.840 197.960 ;
        RECT 188.920 197.640 189.240 197.960 ;
        RECT 189.320 197.640 189.640 197.960 ;
        RECT 189.720 197.640 190.040 197.960 ;
        RECT 190.120 197.640 190.440 197.960 ;
        RECT 190.520 197.640 190.840 197.960 ;
        RECT 190.920 197.640 191.240 197.960 ;
        RECT 191.320 197.640 191.640 197.960 ;
        RECT 191.720 197.640 192.040 197.960 ;
        RECT 192.120 197.640 192.440 197.960 ;
        RECT 192.520 197.640 192.840 197.960 ;
        RECT 192.920 197.640 193.240 197.960 ;
        RECT 193.320 197.640 193.640 197.960 ;
        RECT 193.720 197.640 194.040 197.960 ;
        RECT 194.120 197.640 194.440 197.960 ;
        RECT 194.520 197.640 194.840 197.960 ;
        RECT 194.920 197.640 195.240 197.960 ;
        RECT 195.320 197.640 195.640 197.960 ;
        RECT 195.720 197.640 196.040 197.960 ;
        RECT 196.120 197.640 196.440 197.960 ;
        RECT 196.520 197.640 196.840 197.960 ;
        RECT 196.920 197.640 197.240 197.960 ;
        RECT 197.320 197.640 197.640 197.960 ;
        RECT 197.720 197.640 198.040 197.960 ;
        RECT 198.120 197.640 198.440 197.960 ;
        RECT 198.520 197.640 198.840 197.960 ;
        RECT 198.920 197.640 199.240 197.960 ;
        RECT 199.320 197.640 199.640 197.960 ;
        RECT 199.720 197.640 200.040 197.960 ;
        RECT 200.120 197.640 200.440 197.960 ;
        RECT 200.520 197.640 200.840 197.960 ;
        RECT 200.920 197.640 201.240 197.960 ;
        RECT 201.320 197.640 201.640 197.960 ;
        RECT 201.720 197.640 202.040 197.960 ;
        RECT 202.120 197.640 202.440 197.960 ;
        RECT 202.520 197.640 202.840 197.960 ;
        RECT 202.920 197.640 203.240 197.960 ;
        RECT 203.320 197.640 203.640 197.960 ;
        RECT 203.720 197.640 204.040 197.960 ;
        RECT 204.120 197.640 204.440 197.960 ;
        RECT 204.520 197.640 204.840 197.960 ;
        RECT 204.920 197.640 205.240 197.960 ;
        RECT 205.320 197.640 205.640 197.960 ;
        RECT 0.040 197.240 0.360 197.560 ;
        RECT 0.440 197.240 0.760 197.560 ;
        RECT 0.840 197.240 1.160 197.560 ;
        RECT 1.240 197.240 1.560 197.560 ;
        RECT 1.640 197.240 1.960 197.560 ;
        RECT 2.040 197.240 2.360 197.560 ;
        RECT 2.440 197.240 2.760 197.560 ;
        RECT 2.840 197.240 3.160 197.560 ;
        RECT 3.240 197.240 3.560 197.560 ;
        RECT 3.640 197.240 3.960 197.560 ;
        RECT 4.040 197.240 4.360 197.560 ;
        RECT 4.440 197.240 4.760 197.560 ;
        RECT 4.840 197.240 5.160 197.560 ;
        RECT 5.240 197.240 5.560 197.560 ;
        RECT 5.640 197.240 5.960 197.560 ;
        RECT 6.040 197.240 6.360 197.560 ;
        RECT 6.440 197.240 6.760 197.560 ;
        RECT 6.840 197.240 7.160 197.560 ;
        RECT 7.240 197.240 7.560 197.560 ;
        RECT 7.640 197.240 7.960 197.560 ;
        RECT 8.040 197.240 8.360 197.560 ;
        RECT 8.440 197.240 8.760 197.560 ;
        RECT 8.840 197.240 9.160 197.560 ;
        RECT 9.240 197.240 9.560 197.560 ;
        RECT 9.640 197.240 9.960 197.560 ;
        RECT 10.040 197.240 10.360 197.560 ;
        RECT 10.440 197.240 10.760 197.560 ;
        RECT 10.840 197.240 11.160 197.560 ;
        RECT 11.240 197.240 11.560 197.560 ;
        RECT 11.640 197.240 11.960 197.560 ;
        RECT 12.040 197.240 12.360 197.560 ;
        RECT 12.440 197.240 12.760 197.560 ;
        RECT 12.840 197.240 13.160 197.560 ;
        RECT 13.240 197.240 13.560 197.560 ;
        RECT 13.640 197.240 13.960 197.560 ;
        RECT 14.040 197.240 14.360 197.560 ;
        RECT 14.440 197.240 14.760 197.560 ;
        RECT 14.840 197.240 15.160 197.560 ;
        RECT 15.240 197.240 15.560 197.560 ;
        RECT 15.640 197.240 15.960 197.560 ;
        RECT 16.040 197.240 16.360 197.560 ;
        RECT 16.440 197.240 16.760 197.560 ;
        RECT 16.840 197.240 17.160 197.560 ;
        RECT 17.240 197.240 17.560 197.560 ;
        RECT 17.640 197.240 17.960 197.560 ;
        RECT 18.040 197.240 18.360 197.560 ;
        RECT 18.440 197.240 18.760 197.560 ;
        RECT 18.840 197.240 19.160 197.560 ;
        RECT 19.240 197.240 19.560 197.560 ;
        RECT 19.640 197.240 19.960 197.560 ;
        RECT 95.560 197.240 95.880 197.560 ;
        RECT 95.960 197.240 96.280 197.560 ;
        RECT 96.360 197.240 96.680 197.560 ;
        RECT 96.760 197.240 97.080 197.560 ;
        RECT 145.560 197.240 145.880 197.560 ;
        RECT 145.960 197.240 146.280 197.560 ;
        RECT 146.360 197.240 146.680 197.560 ;
        RECT 146.760 197.240 147.080 197.560 ;
        RECT 185.720 197.240 186.040 197.560 ;
        RECT 186.120 197.240 186.440 197.560 ;
        RECT 186.520 197.240 186.840 197.560 ;
        RECT 186.920 197.240 187.240 197.560 ;
        RECT 187.320 197.240 187.640 197.560 ;
        RECT 187.720 197.240 188.040 197.560 ;
        RECT 188.120 197.240 188.440 197.560 ;
        RECT 188.520 197.240 188.840 197.560 ;
        RECT 188.920 197.240 189.240 197.560 ;
        RECT 189.320 197.240 189.640 197.560 ;
        RECT 189.720 197.240 190.040 197.560 ;
        RECT 190.120 197.240 190.440 197.560 ;
        RECT 190.520 197.240 190.840 197.560 ;
        RECT 190.920 197.240 191.240 197.560 ;
        RECT 191.320 197.240 191.640 197.560 ;
        RECT 191.720 197.240 192.040 197.560 ;
        RECT 192.120 197.240 192.440 197.560 ;
        RECT 192.520 197.240 192.840 197.560 ;
        RECT 192.920 197.240 193.240 197.560 ;
        RECT 193.320 197.240 193.640 197.560 ;
        RECT 193.720 197.240 194.040 197.560 ;
        RECT 194.120 197.240 194.440 197.560 ;
        RECT 194.520 197.240 194.840 197.560 ;
        RECT 194.920 197.240 195.240 197.560 ;
        RECT 195.320 197.240 195.640 197.560 ;
        RECT 195.720 197.240 196.040 197.560 ;
        RECT 196.120 197.240 196.440 197.560 ;
        RECT 196.520 197.240 196.840 197.560 ;
        RECT 196.920 197.240 197.240 197.560 ;
        RECT 197.320 197.240 197.640 197.560 ;
        RECT 197.720 197.240 198.040 197.560 ;
        RECT 198.120 197.240 198.440 197.560 ;
        RECT 198.520 197.240 198.840 197.560 ;
        RECT 198.920 197.240 199.240 197.560 ;
        RECT 199.320 197.240 199.640 197.560 ;
        RECT 199.720 197.240 200.040 197.560 ;
        RECT 200.120 197.240 200.440 197.560 ;
        RECT 200.520 197.240 200.840 197.560 ;
        RECT 200.920 197.240 201.240 197.560 ;
        RECT 201.320 197.240 201.640 197.560 ;
        RECT 201.720 197.240 202.040 197.560 ;
        RECT 202.120 197.240 202.440 197.560 ;
        RECT 202.520 197.240 202.840 197.560 ;
        RECT 202.920 197.240 203.240 197.560 ;
        RECT 203.320 197.240 203.640 197.560 ;
        RECT 203.720 197.240 204.040 197.560 ;
        RECT 204.120 197.240 204.440 197.560 ;
        RECT 204.520 197.240 204.840 197.560 ;
        RECT 204.920 197.240 205.240 197.560 ;
        RECT 205.320 197.240 205.640 197.560 ;
        RECT 0.040 196.840 0.360 197.160 ;
        RECT 0.440 196.840 0.760 197.160 ;
        RECT 0.840 196.840 1.160 197.160 ;
        RECT 1.240 196.840 1.560 197.160 ;
        RECT 1.640 196.840 1.960 197.160 ;
        RECT 2.040 196.840 2.360 197.160 ;
        RECT 2.440 196.840 2.760 197.160 ;
        RECT 2.840 196.840 3.160 197.160 ;
        RECT 3.240 196.840 3.560 197.160 ;
        RECT 3.640 196.840 3.960 197.160 ;
        RECT 4.040 196.840 4.360 197.160 ;
        RECT 4.440 196.840 4.760 197.160 ;
        RECT 4.840 196.840 5.160 197.160 ;
        RECT 5.240 196.840 5.560 197.160 ;
        RECT 5.640 196.840 5.960 197.160 ;
        RECT 6.040 196.840 6.360 197.160 ;
        RECT 6.440 196.840 6.760 197.160 ;
        RECT 6.840 196.840 7.160 197.160 ;
        RECT 7.240 196.840 7.560 197.160 ;
        RECT 7.640 196.840 7.960 197.160 ;
        RECT 8.040 196.840 8.360 197.160 ;
        RECT 8.440 196.840 8.760 197.160 ;
        RECT 8.840 196.840 9.160 197.160 ;
        RECT 9.240 196.840 9.560 197.160 ;
        RECT 9.640 196.840 9.960 197.160 ;
        RECT 10.040 196.840 10.360 197.160 ;
        RECT 10.440 196.840 10.760 197.160 ;
        RECT 10.840 196.840 11.160 197.160 ;
        RECT 11.240 196.840 11.560 197.160 ;
        RECT 11.640 196.840 11.960 197.160 ;
        RECT 12.040 196.840 12.360 197.160 ;
        RECT 12.440 196.840 12.760 197.160 ;
        RECT 12.840 196.840 13.160 197.160 ;
        RECT 13.240 196.840 13.560 197.160 ;
        RECT 13.640 196.840 13.960 197.160 ;
        RECT 14.040 196.840 14.360 197.160 ;
        RECT 14.440 196.840 14.760 197.160 ;
        RECT 14.840 196.840 15.160 197.160 ;
        RECT 15.240 196.840 15.560 197.160 ;
        RECT 15.640 196.840 15.960 197.160 ;
        RECT 16.040 196.840 16.360 197.160 ;
        RECT 16.440 196.840 16.760 197.160 ;
        RECT 16.840 196.840 17.160 197.160 ;
        RECT 17.240 196.840 17.560 197.160 ;
        RECT 17.640 196.840 17.960 197.160 ;
        RECT 18.040 196.840 18.360 197.160 ;
        RECT 18.440 196.840 18.760 197.160 ;
        RECT 18.840 196.840 19.160 197.160 ;
        RECT 19.240 196.840 19.560 197.160 ;
        RECT 19.640 196.840 19.960 197.160 ;
        RECT 95.560 196.840 95.880 197.160 ;
        RECT 95.960 196.840 96.280 197.160 ;
        RECT 96.360 196.840 96.680 197.160 ;
        RECT 96.760 196.840 97.080 197.160 ;
        RECT 145.560 196.840 145.880 197.160 ;
        RECT 145.960 196.840 146.280 197.160 ;
        RECT 146.360 196.840 146.680 197.160 ;
        RECT 146.760 196.840 147.080 197.160 ;
        RECT 185.720 196.840 186.040 197.160 ;
        RECT 186.120 196.840 186.440 197.160 ;
        RECT 186.520 196.840 186.840 197.160 ;
        RECT 186.920 196.840 187.240 197.160 ;
        RECT 187.320 196.840 187.640 197.160 ;
        RECT 187.720 196.840 188.040 197.160 ;
        RECT 188.120 196.840 188.440 197.160 ;
        RECT 188.520 196.840 188.840 197.160 ;
        RECT 188.920 196.840 189.240 197.160 ;
        RECT 189.320 196.840 189.640 197.160 ;
        RECT 189.720 196.840 190.040 197.160 ;
        RECT 190.120 196.840 190.440 197.160 ;
        RECT 190.520 196.840 190.840 197.160 ;
        RECT 190.920 196.840 191.240 197.160 ;
        RECT 191.320 196.840 191.640 197.160 ;
        RECT 191.720 196.840 192.040 197.160 ;
        RECT 192.120 196.840 192.440 197.160 ;
        RECT 192.520 196.840 192.840 197.160 ;
        RECT 192.920 196.840 193.240 197.160 ;
        RECT 193.320 196.840 193.640 197.160 ;
        RECT 193.720 196.840 194.040 197.160 ;
        RECT 194.120 196.840 194.440 197.160 ;
        RECT 194.520 196.840 194.840 197.160 ;
        RECT 194.920 196.840 195.240 197.160 ;
        RECT 195.320 196.840 195.640 197.160 ;
        RECT 195.720 196.840 196.040 197.160 ;
        RECT 196.120 196.840 196.440 197.160 ;
        RECT 196.520 196.840 196.840 197.160 ;
        RECT 196.920 196.840 197.240 197.160 ;
        RECT 197.320 196.840 197.640 197.160 ;
        RECT 197.720 196.840 198.040 197.160 ;
        RECT 198.120 196.840 198.440 197.160 ;
        RECT 198.520 196.840 198.840 197.160 ;
        RECT 198.920 196.840 199.240 197.160 ;
        RECT 199.320 196.840 199.640 197.160 ;
        RECT 199.720 196.840 200.040 197.160 ;
        RECT 200.120 196.840 200.440 197.160 ;
        RECT 200.520 196.840 200.840 197.160 ;
        RECT 200.920 196.840 201.240 197.160 ;
        RECT 201.320 196.840 201.640 197.160 ;
        RECT 201.720 196.840 202.040 197.160 ;
        RECT 202.120 196.840 202.440 197.160 ;
        RECT 202.520 196.840 202.840 197.160 ;
        RECT 202.920 196.840 203.240 197.160 ;
        RECT 203.320 196.840 203.640 197.160 ;
        RECT 203.720 196.840 204.040 197.160 ;
        RECT 204.120 196.840 204.440 197.160 ;
        RECT 204.520 196.840 204.840 197.160 ;
        RECT 204.920 196.840 205.240 197.160 ;
        RECT 205.320 196.840 205.640 197.160 ;
        RECT 0.040 196.440 0.360 196.760 ;
        RECT 0.440 196.440 0.760 196.760 ;
        RECT 0.840 196.440 1.160 196.760 ;
        RECT 1.240 196.440 1.560 196.760 ;
        RECT 1.640 196.440 1.960 196.760 ;
        RECT 2.040 196.440 2.360 196.760 ;
        RECT 2.440 196.440 2.760 196.760 ;
        RECT 2.840 196.440 3.160 196.760 ;
        RECT 3.240 196.440 3.560 196.760 ;
        RECT 3.640 196.440 3.960 196.760 ;
        RECT 4.040 196.440 4.360 196.760 ;
        RECT 4.440 196.440 4.760 196.760 ;
        RECT 4.840 196.440 5.160 196.760 ;
        RECT 5.240 196.440 5.560 196.760 ;
        RECT 5.640 196.440 5.960 196.760 ;
        RECT 6.040 196.440 6.360 196.760 ;
        RECT 6.440 196.440 6.760 196.760 ;
        RECT 6.840 196.440 7.160 196.760 ;
        RECT 7.240 196.440 7.560 196.760 ;
        RECT 7.640 196.440 7.960 196.760 ;
        RECT 8.040 196.440 8.360 196.760 ;
        RECT 8.440 196.440 8.760 196.760 ;
        RECT 8.840 196.440 9.160 196.760 ;
        RECT 9.240 196.440 9.560 196.760 ;
        RECT 9.640 196.440 9.960 196.760 ;
        RECT 10.040 196.440 10.360 196.760 ;
        RECT 10.440 196.440 10.760 196.760 ;
        RECT 10.840 196.440 11.160 196.760 ;
        RECT 11.240 196.440 11.560 196.760 ;
        RECT 11.640 196.440 11.960 196.760 ;
        RECT 12.040 196.440 12.360 196.760 ;
        RECT 12.440 196.440 12.760 196.760 ;
        RECT 12.840 196.440 13.160 196.760 ;
        RECT 13.240 196.440 13.560 196.760 ;
        RECT 13.640 196.440 13.960 196.760 ;
        RECT 14.040 196.440 14.360 196.760 ;
        RECT 14.440 196.440 14.760 196.760 ;
        RECT 14.840 196.440 15.160 196.760 ;
        RECT 15.240 196.440 15.560 196.760 ;
        RECT 15.640 196.440 15.960 196.760 ;
        RECT 16.040 196.440 16.360 196.760 ;
        RECT 16.440 196.440 16.760 196.760 ;
        RECT 16.840 196.440 17.160 196.760 ;
        RECT 17.240 196.440 17.560 196.760 ;
        RECT 17.640 196.440 17.960 196.760 ;
        RECT 18.040 196.440 18.360 196.760 ;
        RECT 18.440 196.440 18.760 196.760 ;
        RECT 18.840 196.440 19.160 196.760 ;
        RECT 19.240 196.440 19.560 196.760 ;
        RECT 19.640 196.440 19.960 196.760 ;
        RECT 95.560 196.440 95.880 196.760 ;
        RECT 95.960 196.440 96.280 196.760 ;
        RECT 96.360 196.440 96.680 196.760 ;
        RECT 96.760 196.440 97.080 196.760 ;
        RECT 145.560 196.440 145.880 196.760 ;
        RECT 145.960 196.440 146.280 196.760 ;
        RECT 146.360 196.440 146.680 196.760 ;
        RECT 146.760 196.440 147.080 196.760 ;
        RECT 185.720 196.440 186.040 196.760 ;
        RECT 186.120 196.440 186.440 196.760 ;
        RECT 186.520 196.440 186.840 196.760 ;
        RECT 186.920 196.440 187.240 196.760 ;
        RECT 187.320 196.440 187.640 196.760 ;
        RECT 187.720 196.440 188.040 196.760 ;
        RECT 188.120 196.440 188.440 196.760 ;
        RECT 188.520 196.440 188.840 196.760 ;
        RECT 188.920 196.440 189.240 196.760 ;
        RECT 189.320 196.440 189.640 196.760 ;
        RECT 189.720 196.440 190.040 196.760 ;
        RECT 190.120 196.440 190.440 196.760 ;
        RECT 190.520 196.440 190.840 196.760 ;
        RECT 190.920 196.440 191.240 196.760 ;
        RECT 191.320 196.440 191.640 196.760 ;
        RECT 191.720 196.440 192.040 196.760 ;
        RECT 192.120 196.440 192.440 196.760 ;
        RECT 192.520 196.440 192.840 196.760 ;
        RECT 192.920 196.440 193.240 196.760 ;
        RECT 193.320 196.440 193.640 196.760 ;
        RECT 193.720 196.440 194.040 196.760 ;
        RECT 194.120 196.440 194.440 196.760 ;
        RECT 194.520 196.440 194.840 196.760 ;
        RECT 194.920 196.440 195.240 196.760 ;
        RECT 195.320 196.440 195.640 196.760 ;
        RECT 195.720 196.440 196.040 196.760 ;
        RECT 196.120 196.440 196.440 196.760 ;
        RECT 196.520 196.440 196.840 196.760 ;
        RECT 196.920 196.440 197.240 196.760 ;
        RECT 197.320 196.440 197.640 196.760 ;
        RECT 197.720 196.440 198.040 196.760 ;
        RECT 198.120 196.440 198.440 196.760 ;
        RECT 198.520 196.440 198.840 196.760 ;
        RECT 198.920 196.440 199.240 196.760 ;
        RECT 199.320 196.440 199.640 196.760 ;
        RECT 199.720 196.440 200.040 196.760 ;
        RECT 200.120 196.440 200.440 196.760 ;
        RECT 200.520 196.440 200.840 196.760 ;
        RECT 200.920 196.440 201.240 196.760 ;
        RECT 201.320 196.440 201.640 196.760 ;
        RECT 201.720 196.440 202.040 196.760 ;
        RECT 202.120 196.440 202.440 196.760 ;
        RECT 202.520 196.440 202.840 196.760 ;
        RECT 202.920 196.440 203.240 196.760 ;
        RECT 203.320 196.440 203.640 196.760 ;
        RECT 203.720 196.440 204.040 196.760 ;
        RECT 204.120 196.440 204.440 196.760 ;
        RECT 204.520 196.440 204.840 196.760 ;
        RECT 204.920 196.440 205.240 196.760 ;
        RECT 205.320 196.440 205.640 196.760 ;
        RECT 0.040 196.040 0.360 196.360 ;
        RECT 0.440 196.040 0.760 196.360 ;
        RECT 0.840 196.040 1.160 196.360 ;
        RECT 1.240 196.040 1.560 196.360 ;
        RECT 1.640 196.040 1.960 196.360 ;
        RECT 2.040 196.040 2.360 196.360 ;
        RECT 2.440 196.040 2.760 196.360 ;
        RECT 2.840 196.040 3.160 196.360 ;
        RECT 3.240 196.040 3.560 196.360 ;
        RECT 3.640 196.040 3.960 196.360 ;
        RECT 4.040 196.040 4.360 196.360 ;
        RECT 4.440 196.040 4.760 196.360 ;
        RECT 4.840 196.040 5.160 196.360 ;
        RECT 5.240 196.040 5.560 196.360 ;
        RECT 5.640 196.040 5.960 196.360 ;
        RECT 6.040 196.040 6.360 196.360 ;
        RECT 6.440 196.040 6.760 196.360 ;
        RECT 6.840 196.040 7.160 196.360 ;
        RECT 7.240 196.040 7.560 196.360 ;
        RECT 7.640 196.040 7.960 196.360 ;
        RECT 8.040 196.040 8.360 196.360 ;
        RECT 8.440 196.040 8.760 196.360 ;
        RECT 8.840 196.040 9.160 196.360 ;
        RECT 9.240 196.040 9.560 196.360 ;
        RECT 9.640 196.040 9.960 196.360 ;
        RECT 10.040 196.040 10.360 196.360 ;
        RECT 10.440 196.040 10.760 196.360 ;
        RECT 10.840 196.040 11.160 196.360 ;
        RECT 11.240 196.040 11.560 196.360 ;
        RECT 11.640 196.040 11.960 196.360 ;
        RECT 12.040 196.040 12.360 196.360 ;
        RECT 12.440 196.040 12.760 196.360 ;
        RECT 12.840 196.040 13.160 196.360 ;
        RECT 13.240 196.040 13.560 196.360 ;
        RECT 13.640 196.040 13.960 196.360 ;
        RECT 14.040 196.040 14.360 196.360 ;
        RECT 14.440 196.040 14.760 196.360 ;
        RECT 14.840 196.040 15.160 196.360 ;
        RECT 15.240 196.040 15.560 196.360 ;
        RECT 15.640 196.040 15.960 196.360 ;
        RECT 16.040 196.040 16.360 196.360 ;
        RECT 16.440 196.040 16.760 196.360 ;
        RECT 16.840 196.040 17.160 196.360 ;
        RECT 17.240 196.040 17.560 196.360 ;
        RECT 17.640 196.040 17.960 196.360 ;
        RECT 18.040 196.040 18.360 196.360 ;
        RECT 18.440 196.040 18.760 196.360 ;
        RECT 18.840 196.040 19.160 196.360 ;
        RECT 19.240 196.040 19.560 196.360 ;
        RECT 19.640 196.040 19.960 196.360 ;
        RECT 95.560 196.040 95.880 196.360 ;
        RECT 95.960 196.040 96.280 196.360 ;
        RECT 96.360 196.040 96.680 196.360 ;
        RECT 96.760 196.040 97.080 196.360 ;
        RECT 145.560 196.040 145.880 196.360 ;
        RECT 145.960 196.040 146.280 196.360 ;
        RECT 146.360 196.040 146.680 196.360 ;
        RECT 146.760 196.040 147.080 196.360 ;
        RECT 185.720 196.040 186.040 196.360 ;
        RECT 186.120 196.040 186.440 196.360 ;
        RECT 186.520 196.040 186.840 196.360 ;
        RECT 186.920 196.040 187.240 196.360 ;
        RECT 187.320 196.040 187.640 196.360 ;
        RECT 187.720 196.040 188.040 196.360 ;
        RECT 188.120 196.040 188.440 196.360 ;
        RECT 188.520 196.040 188.840 196.360 ;
        RECT 188.920 196.040 189.240 196.360 ;
        RECT 189.320 196.040 189.640 196.360 ;
        RECT 189.720 196.040 190.040 196.360 ;
        RECT 190.120 196.040 190.440 196.360 ;
        RECT 190.520 196.040 190.840 196.360 ;
        RECT 190.920 196.040 191.240 196.360 ;
        RECT 191.320 196.040 191.640 196.360 ;
        RECT 191.720 196.040 192.040 196.360 ;
        RECT 192.120 196.040 192.440 196.360 ;
        RECT 192.520 196.040 192.840 196.360 ;
        RECT 192.920 196.040 193.240 196.360 ;
        RECT 193.320 196.040 193.640 196.360 ;
        RECT 193.720 196.040 194.040 196.360 ;
        RECT 194.120 196.040 194.440 196.360 ;
        RECT 194.520 196.040 194.840 196.360 ;
        RECT 194.920 196.040 195.240 196.360 ;
        RECT 195.320 196.040 195.640 196.360 ;
        RECT 195.720 196.040 196.040 196.360 ;
        RECT 196.120 196.040 196.440 196.360 ;
        RECT 196.520 196.040 196.840 196.360 ;
        RECT 196.920 196.040 197.240 196.360 ;
        RECT 197.320 196.040 197.640 196.360 ;
        RECT 197.720 196.040 198.040 196.360 ;
        RECT 198.120 196.040 198.440 196.360 ;
        RECT 198.520 196.040 198.840 196.360 ;
        RECT 198.920 196.040 199.240 196.360 ;
        RECT 199.320 196.040 199.640 196.360 ;
        RECT 199.720 196.040 200.040 196.360 ;
        RECT 200.120 196.040 200.440 196.360 ;
        RECT 200.520 196.040 200.840 196.360 ;
        RECT 200.920 196.040 201.240 196.360 ;
        RECT 201.320 196.040 201.640 196.360 ;
        RECT 201.720 196.040 202.040 196.360 ;
        RECT 202.120 196.040 202.440 196.360 ;
        RECT 202.520 196.040 202.840 196.360 ;
        RECT 202.920 196.040 203.240 196.360 ;
        RECT 203.320 196.040 203.640 196.360 ;
        RECT 203.720 196.040 204.040 196.360 ;
        RECT 204.120 196.040 204.440 196.360 ;
        RECT 204.520 196.040 204.840 196.360 ;
        RECT 204.920 196.040 205.240 196.360 ;
        RECT 205.320 196.040 205.640 196.360 ;
        RECT 0.040 195.640 0.360 195.960 ;
        RECT 0.440 195.640 0.760 195.960 ;
        RECT 0.840 195.640 1.160 195.960 ;
        RECT 1.240 195.640 1.560 195.960 ;
        RECT 1.640 195.640 1.960 195.960 ;
        RECT 2.040 195.640 2.360 195.960 ;
        RECT 2.440 195.640 2.760 195.960 ;
        RECT 2.840 195.640 3.160 195.960 ;
        RECT 3.240 195.640 3.560 195.960 ;
        RECT 3.640 195.640 3.960 195.960 ;
        RECT 4.040 195.640 4.360 195.960 ;
        RECT 4.440 195.640 4.760 195.960 ;
        RECT 4.840 195.640 5.160 195.960 ;
        RECT 5.240 195.640 5.560 195.960 ;
        RECT 5.640 195.640 5.960 195.960 ;
        RECT 6.040 195.640 6.360 195.960 ;
        RECT 6.440 195.640 6.760 195.960 ;
        RECT 6.840 195.640 7.160 195.960 ;
        RECT 7.240 195.640 7.560 195.960 ;
        RECT 7.640 195.640 7.960 195.960 ;
        RECT 8.040 195.640 8.360 195.960 ;
        RECT 8.440 195.640 8.760 195.960 ;
        RECT 8.840 195.640 9.160 195.960 ;
        RECT 9.240 195.640 9.560 195.960 ;
        RECT 9.640 195.640 9.960 195.960 ;
        RECT 10.040 195.640 10.360 195.960 ;
        RECT 10.440 195.640 10.760 195.960 ;
        RECT 10.840 195.640 11.160 195.960 ;
        RECT 11.240 195.640 11.560 195.960 ;
        RECT 11.640 195.640 11.960 195.960 ;
        RECT 12.040 195.640 12.360 195.960 ;
        RECT 12.440 195.640 12.760 195.960 ;
        RECT 12.840 195.640 13.160 195.960 ;
        RECT 13.240 195.640 13.560 195.960 ;
        RECT 13.640 195.640 13.960 195.960 ;
        RECT 14.040 195.640 14.360 195.960 ;
        RECT 14.440 195.640 14.760 195.960 ;
        RECT 14.840 195.640 15.160 195.960 ;
        RECT 15.240 195.640 15.560 195.960 ;
        RECT 15.640 195.640 15.960 195.960 ;
        RECT 16.040 195.640 16.360 195.960 ;
        RECT 16.440 195.640 16.760 195.960 ;
        RECT 16.840 195.640 17.160 195.960 ;
        RECT 17.240 195.640 17.560 195.960 ;
        RECT 17.640 195.640 17.960 195.960 ;
        RECT 18.040 195.640 18.360 195.960 ;
        RECT 18.440 195.640 18.760 195.960 ;
        RECT 18.840 195.640 19.160 195.960 ;
        RECT 19.240 195.640 19.560 195.960 ;
        RECT 19.640 195.640 19.960 195.960 ;
        RECT 95.560 195.640 95.880 195.960 ;
        RECT 95.960 195.640 96.280 195.960 ;
        RECT 96.360 195.640 96.680 195.960 ;
        RECT 96.760 195.640 97.080 195.960 ;
        RECT 145.560 195.640 145.880 195.960 ;
        RECT 145.960 195.640 146.280 195.960 ;
        RECT 146.360 195.640 146.680 195.960 ;
        RECT 146.760 195.640 147.080 195.960 ;
        RECT 185.720 195.640 186.040 195.960 ;
        RECT 186.120 195.640 186.440 195.960 ;
        RECT 186.520 195.640 186.840 195.960 ;
        RECT 186.920 195.640 187.240 195.960 ;
        RECT 187.320 195.640 187.640 195.960 ;
        RECT 187.720 195.640 188.040 195.960 ;
        RECT 188.120 195.640 188.440 195.960 ;
        RECT 188.520 195.640 188.840 195.960 ;
        RECT 188.920 195.640 189.240 195.960 ;
        RECT 189.320 195.640 189.640 195.960 ;
        RECT 189.720 195.640 190.040 195.960 ;
        RECT 190.120 195.640 190.440 195.960 ;
        RECT 190.520 195.640 190.840 195.960 ;
        RECT 190.920 195.640 191.240 195.960 ;
        RECT 191.320 195.640 191.640 195.960 ;
        RECT 191.720 195.640 192.040 195.960 ;
        RECT 192.120 195.640 192.440 195.960 ;
        RECT 192.520 195.640 192.840 195.960 ;
        RECT 192.920 195.640 193.240 195.960 ;
        RECT 193.320 195.640 193.640 195.960 ;
        RECT 193.720 195.640 194.040 195.960 ;
        RECT 194.120 195.640 194.440 195.960 ;
        RECT 194.520 195.640 194.840 195.960 ;
        RECT 194.920 195.640 195.240 195.960 ;
        RECT 195.320 195.640 195.640 195.960 ;
        RECT 195.720 195.640 196.040 195.960 ;
        RECT 196.120 195.640 196.440 195.960 ;
        RECT 196.520 195.640 196.840 195.960 ;
        RECT 196.920 195.640 197.240 195.960 ;
        RECT 197.320 195.640 197.640 195.960 ;
        RECT 197.720 195.640 198.040 195.960 ;
        RECT 198.120 195.640 198.440 195.960 ;
        RECT 198.520 195.640 198.840 195.960 ;
        RECT 198.920 195.640 199.240 195.960 ;
        RECT 199.320 195.640 199.640 195.960 ;
        RECT 199.720 195.640 200.040 195.960 ;
        RECT 200.120 195.640 200.440 195.960 ;
        RECT 200.520 195.640 200.840 195.960 ;
        RECT 200.920 195.640 201.240 195.960 ;
        RECT 201.320 195.640 201.640 195.960 ;
        RECT 201.720 195.640 202.040 195.960 ;
        RECT 202.120 195.640 202.440 195.960 ;
        RECT 202.520 195.640 202.840 195.960 ;
        RECT 202.920 195.640 203.240 195.960 ;
        RECT 203.320 195.640 203.640 195.960 ;
        RECT 203.720 195.640 204.040 195.960 ;
        RECT 204.120 195.640 204.440 195.960 ;
        RECT 204.520 195.640 204.840 195.960 ;
        RECT 204.920 195.640 205.240 195.960 ;
        RECT 205.320 195.640 205.640 195.960 ;
        RECT 0.040 195.240 0.360 195.560 ;
        RECT 0.440 195.240 0.760 195.560 ;
        RECT 0.840 195.240 1.160 195.560 ;
        RECT 1.240 195.240 1.560 195.560 ;
        RECT 1.640 195.240 1.960 195.560 ;
        RECT 2.040 195.240 2.360 195.560 ;
        RECT 2.440 195.240 2.760 195.560 ;
        RECT 2.840 195.240 3.160 195.560 ;
        RECT 3.240 195.240 3.560 195.560 ;
        RECT 3.640 195.240 3.960 195.560 ;
        RECT 4.040 195.240 4.360 195.560 ;
        RECT 4.440 195.240 4.760 195.560 ;
        RECT 4.840 195.240 5.160 195.560 ;
        RECT 5.240 195.240 5.560 195.560 ;
        RECT 5.640 195.240 5.960 195.560 ;
        RECT 6.040 195.240 6.360 195.560 ;
        RECT 6.440 195.240 6.760 195.560 ;
        RECT 6.840 195.240 7.160 195.560 ;
        RECT 7.240 195.240 7.560 195.560 ;
        RECT 7.640 195.240 7.960 195.560 ;
        RECT 8.040 195.240 8.360 195.560 ;
        RECT 8.440 195.240 8.760 195.560 ;
        RECT 8.840 195.240 9.160 195.560 ;
        RECT 9.240 195.240 9.560 195.560 ;
        RECT 9.640 195.240 9.960 195.560 ;
        RECT 10.040 195.240 10.360 195.560 ;
        RECT 10.440 195.240 10.760 195.560 ;
        RECT 10.840 195.240 11.160 195.560 ;
        RECT 11.240 195.240 11.560 195.560 ;
        RECT 11.640 195.240 11.960 195.560 ;
        RECT 12.040 195.240 12.360 195.560 ;
        RECT 12.440 195.240 12.760 195.560 ;
        RECT 12.840 195.240 13.160 195.560 ;
        RECT 13.240 195.240 13.560 195.560 ;
        RECT 13.640 195.240 13.960 195.560 ;
        RECT 14.040 195.240 14.360 195.560 ;
        RECT 14.440 195.240 14.760 195.560 ;
        RECT 14.840 195.240 15.160 195.560 ;
        RECT 15.240 195.240 15.560 195.560 ;
        RECT 15.640 195.240 15.960 195.560 ;
        RECT 16.040 195.240 16.360 195.560 ;
        RECT 16.440 195.240 16.760 195.560 ;
        RECT 16.840 195.240 17.160 195.560 ;
        RECT 17.240 195.240 17.560 195.560 ;
        RECT 17.640 195.240 17.960 195.560 ;
        RECT 18.040 195.240 18.360 195.560 ;
        RECT 18.440 195.240 18.760 195.560 ;
        RECT 18.840 195.240 19.160 195.560 ;
        RECT 19.240 195.240 19.560 195.560 ;
        RECT 19.640 195.240 19.960 195.560 ;
        RECT 95.560 195.240 95.880 195.560 ;
        RECT 95.960 195.240 96.280 195.560 ;
        RECT 96.360 195.240 96.680 195.560 ;
        RECT 96.760 195.240 97.080 195.560 ;
        RECT 145.560 195.240 145.880 195.560 ;
        RECT 145.960 195.240 146.280 195.560 ;
        RECT 146.360 195.240 146.680 195.560 ;
        RECT 146.760 195.240 147.080 195.560 ;
        RECT 185.720 195.240 186.040 195.560 ;
        RECT 186.120 195.240 186.440 195.560 ;
        RECT 186.520 195.240 186.840 195.560 ;
        RECT 186.920 195.240 187.240 195.560 ;
        RECT 187.320 195.240 187.640 195.560 ;
        RECT 187.720 195.240 188.040 195.560 ;
        RECT 188.120 195.240 188.440 195.560 ;
        RECT 188.520 195.240 188.840 195.560 ;
        RECT 188.920 195.240 189.240 195.560 ;
        RECT 189.320 195.240 189.640 195.560 ;
        RECT 189.720 195.240 190.040 195.560 ;
        RECT 190.120 195.240 190.440 195.560 ;
        RECT 190.520 195.240 190.840 195.560 ;
        RECT 190.920 195.240 191.240 195.560 ;
        RECT 191.320 195.240 191.640 195.560 ;
        RECT 191.720 195.240 192.040 195.560 ;
        RECT 192.120 195.240 192.440 195.560 ;
        RECT 192.520 195.240 192.840 195.560 ;
        RECT 192.920 195.240 193.240 195.560 ;
        RECT 193.320 195.240 193.640 195.560 ;
        RECT 193.720 195.240 194.040 195.560 ;
        RECT 194.120 195.240 194.440 195.560 ;
        RECT 194.520 195.240 194.840 195.560 ;
        RECT 194.920 195.240 195.240 195.560 ;
        RECT 195.320 195.240 195.640 195.560 ;
        RECT 195.720 195.240 196.040 195.560 ;
        RECT 196.120 195.240 196.440 195.560 ;
        RECT 196.520 195.240 196.840 195.560 ;
        RECT 196.920 195.240 197.240 195.560 ;
        RECT 197.320 195.240 197.640 195.560 ;
        RECT 197.720 195.240 198.040 195.560 ;
        RECT 198.120 195.240 198.440 195.560 ;
        RECT 198.520 195.240 198.840 195.560 ;
        RECT 198.920 195.240 199.240 195.560 ;
        RECT 199.320 195.240 199.640 195.560 ;
        RECT 199.720 195.240 200.040 195.560 ;
        RECT 200.120 195.240 200.440 195.560 ;
        RECT 200.520 195.240 200.840 195.560 ;
        RECT 200.920 195.240 201.240 195.560 ;
        RECT 201.320 195.240 201.640 195.560 ;
        RECT 201.720 195.240 202.040 195.560 ;
        RECT 202.120 195.240 202.440 195.560 ;
        RECT 202.520 195.240 202.840 195.560 ;
        RECT 202.920 195.240 203.240 195.560 ;
        RECT 203.320 195.240 203.640 195.560 ;
        RECT 203.720 195.240 204.040 195.560 ;
        RECT 204.120 195.240 204.440 195.560 ;
        RECT 204.520 195.240 204.840 195.560 ;
        RECT 204.920 195.240 205.240 195.560 ;
        RECT 205.320 195.240 205.640 195.560 ;
        RECT 0.040 194.840 0.360 195.160 ;
        RECT 0.440 194.840 0.760 195.160 ;
        RECT 0.840 194.840 1.160 195.160 ;
        RECT 1.240 194.840 1.560 195.160 ;
        RECT 1.640 194.840 1.960 195.160 ;
        RECT 2.040 194.840 2.360 195.160 ;
        RECT 2.440 194.840 2.760 195.160 ;
        RECT 2.840 194.840 3.160 195.160 ;
        RECT 3.240 194.840 3.560 195.160 ;
        RECT 3.640 194.840 3.960 195.160 ;
        RECT 4.040 194.840 4.360 195.160 ;
        RECT 4.440 194.840 4.760 195.160 ;
        RECT 4.840 194.840 5.160 195.160 ;
        RECT 5.240 194.840 5.560 195.160 ;
        RECT 5.640 194.840 5.960 195.160 ;
        RECT 6.040 194.840 6.360 195.160 ;
        RECT 6.440 194.840 6.760 195.160 ;
        RECT 6.840 194.840 7.160 195.160 ;
        RECT 7.240 194.840 7.560 195.160 ;
        RECT 7.640 194.840 7.960 195.160 ;
        RECT 8.040 194.840 8.360 195.160 ;
        RECT 8.440 194.840 8.760 195.160 ;
        RECT 8.840 194.840 9.160 195.160 ;
        RECT 9.240 194.840 9.560 195.160 ;
        RECT 9.640 194.840 9.960 195.160 ;
        RECT 10.040 194.840 10.360 195.160 ;
        RECT 10.440 194.840 10.760 195.160 ;
        RECT 10.840 194.840 11.160 195.160 ;
        RECT 11.240 194.840 11.560 195.160 ;
        RECT 11.640 194.840 11.960 195.160 ;
        RECT 12.040 194.840 12.360 195.160 ;
        RECT 12.440 194.840 12.760 195.160 ;
        RECT 12.840 194.840 13.160 195.160 ;
        RECT 13.240 194.840 13.560 195.160 ;
        RECT 13.640 194.840 13.960 195.160 ;
        RECT 14.040 194.840 14.360 195.160 ;
        RECT 14.440 194.840 14.760 195.160 ;
        RECT 14.840 194.840 15.160 195.160 ;
        RECT 15.240 194.840 15.560 195.160 ;
        RECT 15.640 194.840 15.960 195.160 ;
        RECT 16.040 194.840 16.360 195.160 ;
        RECT 16.440 194.840 16.760 195.160 ;
        RECT 16.840 194.840 17.160 195.160 ;
        RECT 17.240 194.840 17.560 195.160 ;
        RECT 17.640 194.840 17.960 195.160 ;
        RECT 18.040 194.840 18.360 195.160 ;
        RECT 18.440 194.840 18.760 195.160 ;
        RECT 18.840 194.840 19.160 195.160 ;
        RECT 19.240 194.840 19.560 195.160 ;
        RECT 19.640 194.840 19.960 195.160 ;
        RECT 95.560 194.840 95.880 195.160 ;
        RECT 95.960 194.840 96.280 195.160 ;
        RECT 96.360 194.840 96.680 195.160 ;
        RECT 96.760 194.840 97.080 195.160 ;
        RECT 145.560 194.840 145.880 195.160 ;
        RECT 145.960 194.840 146.280 195.160 ;
        RECT 146.360 194.840 146.680 195.160 ;
        RECT 146.760 194.840 147.080 195.160 ;
        RECT 185.720 194.840 186.040 195.160 ;
        RECT 186.120 194.840 186.440 195.160 ;
        RECT 186.520 194.840 186.840 195.160 ;
        RECT 186.920 194.840 187.240 195.160 ;
        RECT 187.320 194.840 187.640 195.160 ;
        RECT 187.720 194.840 188.040 195.160 ;
        RECT 188.120 194.840 188.440 195.160 ;
        RECT 188.520 194.840 188.840 195.160 ;
        RECT 188.920 194.840 189.240 195.160 ;
        RECT 189.320 194.840 189.640 195.160 ;
        RECT 189.720 194.840 190.040 195.160 ;
        RECT 190.120 194.840 190.440 195.160 ;
        RECT 190.520 194.840 190.840 195.160 ;
        RECT 190.920 194.840 191.240 195.160 ;
        RECT 191.320 194.840 191.640 195.160 ;
        RECT 191.720 194.840 192.040 195.160 ;
        RECT 192.120 194.840 192.440 195.160 ;
        RECT 192.520 194.840 192.840 195.160 ;
        RECT 192.920 194.840 193.240 195.160 ;
        RECT 193.320 194.840 193.640 195.160 ;
        RECT 193.720 194.840 194.040 195.160 ;
        RECT 194.120 194.840 194.440 195.160 ;
        RECT 194.520 194.840 194.840 195.160 ;
        RECT 194.920 194.840 195.240 195.160 ;
        RECT 195.320 194.840 195.640 195.160 ;
        RECT 195.720 194.840 196.040 195.160 ;
        RECT 196.120 194.840 196.440 195.160 ;
        RECT 196.520 194.840 196.840 195.160 ;
        RECT 196.920 194.840 197.240 195.160 ;
        RECT 197.320 194.840 197.640 195.160 ;
        RECT 197.720 194.840 198.040 195.160 ;
        RECT 198.120 194.840 198.440 195.160 ;
        RECT 198.520 194.840 198.840 195.160 ;
        RECT 198.920 194.840 199.240 195.160 ;
        RECT 199.320 194.840 199.640 195.160 ;
        RECT 199.720 194.840 200.040 195.160 ;
        RECT 200.120 194.840 200.440 195.160 ;
        RECT 200.520 194.840 200.840 195.160 ;
        RECT 200.920 194.840 201.240 195.160 ;
        RECT 201.320 194.840 201.640 195.160 ;
        RECT 201.720 194.840 202.040 195.160 ;
        RECT 202.120 194.840 202.440 195.160 ;
        RECT 202.520 194.840 202.840 195.160 ;
        RECT 202.920 194.840 203.240 195.160 ;
        RECT 203.320 194.840 203.640 195.160 ;
        RECT 203.720 194.840 204.040 195.160 ;
        RECT 204.120 194.840 204.440 195.160 ;
        RECT 204.520 194.840 204.840 195.160 ;
        RECT 204.920 194.840 205.240 195.160 ;
        RECT 205.320 194.840 205.640 195.160 ;
        RECT 0.040 194.440 0.360 194.760 ;
        RECT 0.440 194.440 0.760 194.760 ;
        RECT 0.840 194.440 1.160 194.760 ;
        RECT 1.240 194.440 1.560 194.760 ;
        RECT 1.640 194.440 1.960 194.760 ;
        RECT 2.040 194.440 2.360 194.760 ;
        RECT 2.440 194.440 2.760 194.760 ;
        RECT 2.840 194.440 3.160 194.760 ;
        RECT 3.240 194.440 3.560 194.760 ;
        RECT 3.640 194.440 3.960 194.760 ;
        RECT 4.040 194.440 4.360 194.760 ;
        RECT 4.440 194.440 4.760 194.760 ;
        RECT 4.840 194.440 5.160 194.760 ;
        RECT 5.240 194.440 5.560 194.760 ;
        RECT 5.640 194.440 5.960 194.760 ;
        RECT 6.040 194.440 6.360 194.760 ;
        RECT 6.440 194.440 6.760 194.760 ;
        RECT 6.840 194.440 7.160 194.760 ;
        RECT 7.240 194.440 7.560 194.760 ;
        RECT 7.640 194.440 7.960 194.760 ;
        RECT 8.040 194.440 8.360 194.760 ;
        RECT 8.440 194.440 8.760 194.760 ;
        RECT 8.840 194.440 9.160 194.760 ;
        RECT 9.240 194.440 9.560 194.760 ;
        RECT 9.640 194.440 9.960 194.760 ;
        RECT 10.040 194.440 10.360 194.760 ;
        RECT 10.440 194.440 10.760 194.760 ;
        RECT 10.840 194.440 11.160 194.760 ;
        RECT 11.240 194.440 11.560 194.760 ;
        RECT 11.640 194.440 11.960 194.760 ;
        RECT 12.040 194.440 12.360 194.760 ;
        RECT 12.440 194.440 12.760 194.760 ;
        RECT 12.840 194.440 13.160 194.760 ;
        RECT 13.240 194.440 13.560 194.760 ;
        RECT 13.640 194.440 13.960 194.760 ;
        RECT 14.040 194.440 14.360 194.760 ;
        RECT 14.440 194.440 14.760 194.760 ;
        RECT 14.840 194.440 15.160 194.760 ;
        RECT 15.240 194.440 15.560 194.760 ;
        RECT 15.640 194.440 15.960 194.760 ;
        RECT 16.040 194.440 16.360 194.760 ;
        RECT 16.440 194.440 16.760 194.760 ;
        RECT 16.840 194.440 17.160 194.760 ;
        RECT 17.240 194.440 17.560 194.760 ;
        RECT 17.640 194.440 17.960 194.760 ;
        RECT 18.040 194.440 18.360 194.760 ;
        RECT 18.440 194.440 18.760 194.760 ;
        RECT 18.840 194.440 19.160 194.760 ;
        RECT 19.240 194.440 19.560 194.760 ;
        RECT 19.640 194.440 19.960 194.760 ;
        RECT 95.560 194.440 95.880 194.760 ;
        RECT 95.960 194.440 96.280 194.760 ;
        RECT 96.360 194.440 96.680 194.760 ;
        RECT 96.760 194.440 97.080 194.760 ;
        RECT 145.560 194.440 145.880 194.760 ;
        RECT 145.960 194.440 146.280 194.760 ;
        RECT 146.360 194.440 146.680 194.760 ;
        RECT 146.760 194.440 147.080 194.760 ;
        RECT 185.720 194.440 186.040 194.760 ;
        RECT 186.120 194.440 186.440 194.760 ;
        RECT 186.520 194.440 186.840 194.760 ;
        RECT 186.920 194.440 187.240 194.760 ;
        RECT 187.320 194.440 187.640 194.760 ;
        RECT 187.720 194.440 188.040 194.760 ;
        RECT 188.120 194.440 188.440 194.760 ;
        RECT 188.520 194.440 188.840 194.760 ;
        RECT 188.920 194.440 189.240 194.760 ;
        RECT 189.320 194.440 189.640 194.760 ;
        RECT 189.720 194.440 190.040 194.760 ;
        RECT 190.120 194.440 190.440 194.760 ;
        RECT 190.520 194.440 190.840 194.760 ;
        RECT 190.920 194.440 191.240 194.760 ;
        RECT 191.320 194.440 191.640 194.760 ;
        RECT 191.720 194.440 192.040 194.760 ;
        RECT 192.120 194.440 192.440 194.760 ;
        RECT 192.520 194.440 192.840 194.760 ;
        RECT 192.920 194.440 193.240 194.760 ;
        RECT 193.320 194.440 193.640 194.760 ;
        RECT 193.720 194.440 194.040 194.760 ;
        RECT 194.120 194.440 194.440 194.760 ;
        RECT 194.520 194.440 194.840 194.760 ;
        RECT 194.920 194.440 195.240 194.760 ;
        RECT 195.320 194.440 195.640 194.760 ;
        RECT 195.720 194.440 196.040 194.760 ;
        RECT 196.120 194.440 196.440 194.760 ;
        RECT 196.520 194.440 196.840 194.760 ;
        RECT 196.920 194.440 197.240 194.760 ;
        RECT 197.320 194.440 197.640 194.760 ;
        RECT 197.720 194.440 198.040 194.760 ;
        RECT 198.120 194.440 198.440 194.760 ;
        RECT 198.520 194.440 198.840 194.760 ;
        RECT 198.920 194.440 199.240 194.760 ;
        RECT 199.320 194.440 199.640 194.760 ;
        RECT 199.720 194.440 200.040 194.760 ;
        RECT 200.120 194.440 200.440 194.760 ;
        RECT 200.520 194.440 200.840 194.760 ;
        RECT 200.920 194.440 201.240 194.760 ;
        RECT 201.320 194.440 201.640 194.760 ;
        RECT 201.720 194.440 202.040 194.760 ;
        RECT 202.120 194.440 202.440 194.760 ;
        RECT 202.520 194.440 202.840 194.760 ;
        RECT 202.920 194.440 203.240 194.760 ;
        RECT 203.320 194.440 203.640 194.760 ;
        RECT 203.720 194.440 204.040 194.760 ;
        RECT 204.120 194.440 204.440 194.760 ;
        RECT 204.520 194.440 204.840 194.760 ;
        RECT 204.920 194.440 205.240 194.760 ;
        RECT 205.320 194.440 205.640 194.760 ;
        RECT 0.040 194.040 0.360 194.360 ;
        RECT 0.440 194.040 0.760 194.360 ;
        RECT 0.840 194.040 1.160 194.360 ;
        RECT 1.240 194.040 1.560 194.360 ;
        RECT 1.640 194.040 1.960 194.360 ;
        RECT 2.040 194.040 2.360 194.360 ;
        RECT 2.440 194.040 2.760 194.360 ;
        RECT 2.840 194.040 3.160 194.360 ;
        RECT 3.240 194.040 3.560 194.360 ;
        RECT 3.640 194.040 3.960 194.360 ;
        RECT 4.040 194.040 4.360 194.360 ;
        RECT 4.440 194.040 4.760 194.360 ;
        RECT 4.840 194.040 5.160 194.360 ;
        RECT 5.240 194.040 5.560 194.360 ;
        RECT 5.640 194.040 5.960 194.360 ;
        RECT 6.040 194.040 6.360 194.360 ;
        RECT 6.440 194.040 6.760 194.360 ;
        RECT 6.840 194.040 7.160 194.360 ;
        RECT 7.240 194.040 7.560 194.360 ;
        RECT 7.640 194.040 7.960 194.360 ;
        RECT 8.040 194.040 8.360 194.360 ;
        RECT 8.440 194.040 8.760 194.360 ;
        RECT 8.840 194.040 9.160 194.360 ;
        RECT 9.240 194.040 9.560 194.360 ;
        RECT 9.640 194.040 9.960 194.360 ;
        RECT 10.040 194.040 10.360 194.360 ;
        RECT 10.440 194.040 10.760 194.360 ;
        RECT 10.840 194.040 11.160 194.360 ;
        RECT 11.240 194.040 11.560 194.360 ;
        RECT 11.640 194.040 11.960 194.360 ;
        RECT 12.040 194.040 12.360 194.360 ;
        RECT 12.440 194.040 12.760 194.360 ;
        RECT 12.840 194.040 13.160 194.360 ;
        RECT 13.240 194.040 13.560 194.360 ;
        RECT 13.640 194.040 13.960 194.360 ;
        RECT 14.040 194.040 14.360 194.360 ;
        RECT 14.440 194.040 14.760 194.360 ;
        RECT 14.840 194.040 15.160 194.360 ;
        RECT 15.240 194.040 15.560 194.360 ;
        RECT 15.640 194.040 15.960 194.360 ;
        RECT 16.040 194.040 16.360 194.360 ;
        RECT 16.440 194.040 16.760 194.360 ;
        RECT 16.840 194.040 17.160 194.360 ;
        RECT 17.240 194.040 17.560 194.360 ;
        RECT 17.640 194.040 17.960 194.360 ;
        RECT 18.040 194.040 18.360 194.360 ;
        RECT 18.440 194.040 18.760 194.360 ;
        RECT 18.840 194.040 19.160 194.360 ;
        RECT 19.240 194.040 19.560 194.360 ;
        RECT 19.640 194.040 19.960 194.360 ;
        RECT 95.560 194.040 95.880 194.360 ;
        RECT 95.960 194.040 96.280 194.360 ;
        RECT 96.360 194.040 96.680 194.360 ;
        RECT 96.760 194.040 97.080 194.360 ;
        RECT 145.560 194.040 145.880 194.360 ;
        RECT 145.960 194.040 146.280 194.360 ;
        RECT 146.360 194.040 146.680 194.360 ;
        RECT 146.760 194.040 147.080 194.360 ;
        RECT 185.720 194.040 186.040 194.360 ;
        RECT 186.120 194.040 186.440 194.360 ;
        RECT 186.520 194.040 186.840 194.360 ;
        RECT 186.920 194.040 187.240 194.360 ;
        RECT 187.320 194.040 187.640 194.360 ;
        RECT 187.720 194.040 188.040 194.360 ;
        RECT 188.120 194.040 188.440 194.360 ;
        RECT 188.520 194.040 188.840 194.360 ;
        RECT 188.920 194.040 189.240 194.360 ;
        RECT 189.320 194.040 189.640 194.360 ;
        RECT 189.720 194.040 190.040 194.360 ;
        RECT 190.120 194.040 190.440 194.360 ;
        RECT 190.520 194.040 190.840 194.360 ;
        RECT 190.920 194.040 191.240 194.360 ;
        RECT 191.320 194.040 191.640 194.360 ;
        RECT 191.720 194.040 192.040 194.360 ;
        RECT 192.120 194.040 192.440 194.360 ;
        RECT 192.520 194.040 192.840 194.360 ;
        RECT 192.920 194.040 193.240 194.360 ;
        RECT 193.320 194.040 193.640 194.360 ;
        RECT 193.720 194.040 194.040 194.360 ;
        RECT 194.120 194.040 194.440 194.360 ;
        RECT 194.520 194.040 194.840 194.360 ;
        RECT 194.920 194.040 195.240 194.360 ;
        RECT 195.320 194.040 195.640 194.360 ;
        RECT 195.720 194.040 196.040 194.360 ;
        RECT 196.120 194.040 196.440 194.360 ;
        RECT 196.520 194.040 196.840 194.360 ;
        RECT 196.920 194.040 197.240 194.360 ;
        RECT 197.320 194.040 197.640 194.360 ;
        RECT 197.720 194.040 198.040 194.360 ;
        RECT 198.120 194.040 198.440 194.360 ;
        RECT 198.520 194.040 198.840 194.360 ;
        RECT 198.920 194.040 199.240 194.360 ;
        RECT 199.320 194.040 199.640 194.360 ;
        RECT 199.720 194.040 200.040 194.360 ;
        RECT 200.120 194.040 200.440 194.360 ;
        RECT 200.520 194.040 200.840 194.360 ;
        RECT 200.920 194.040 201.240 194.360 ;
        RECT 201.320 194.040 201.640 194.360 ;
        RECT 201.720 194.040 202.040 194.360 ;
        RECT 202.120 194.040 202.440 194.360 ;
        RECT 202.520 194.040 202.840 194.360 ;
        RECT 202.920 194.040 203.240 194.360 ;
        RECT 203.320 194.040 203.640 194.360 ;
        RECT 203.720 194.040 204.040 194.360 ;
        RECT 204.120 194.040 204.440 194.360 ;
        RECT 204.520 194.040 204.840 194.360 ;
        RECT 204.920 194.040 205.240 194.360 ;
        RECT 205.320 194.040 205.640 194.360 ;
        RECT 0.040 193.640 0.360 193.960 ;
        RECT 0.440 193.640 0.760 193.960 ;
        RECT 0.840 193.640 1.160 193.960 ;
        RECT 1.240 193.640 1.560 193.960 ;
        RECT 1.640 193.640 1.960 193.960 ;
        RECT 2.040 193.640 2.360 193.960 ;
        RECT 2.440 193.640 2.760 193.960 ;
        RECT 2.840 193.640 3.160 193.960 ;
        RECT 3.240 193.640 3.560 193.960 ;
        RECT 3.640 193.640 3.960 193.960 ;
        RECT 4.040 193.640 4.360 193.960 ;
        RECT 4.440 193.640 4.760 193.960 ;
        RECT 4.840 193.640 5.160 193.960 ;
        RECT 5.240 193.640 5.560 193.960 ;
        RECT 5.640 193.640 5.960 193.960 ;
        RECT 6.040 193.640 6.360 193.960 ;
        RECT 6.440 193.640 6.760 193.960 ;
        RECT 6.840 193.640 7.160 193.960 ;
        RECT 7.240 193.640 7.560 193.960 ;
        RECT 7.640 193.640 7.960 193.960 ;
        RECT 8.040 193.640 8.360 193.960 ;
        RECT 8.440 193.640 8.760 193.960 ;
        RECT 8.840 193.640 9.160 193.960 ;
        RECT 9.240 193.640 9.560 193.960 ;
        RECT 9.640 193.640 9.960 193.960 ;
        RECT 10.040 193.640 10.360 193.960 ;
        RECT 10.440 193.640 10.760 193.960 ;
        RECT 10.840 193.640 11.160 193.960 ;
        RECT 11.240 193.640 11.560 193.960 ;
        RECT 11.640 193.640 11.960 193.960 ;
        RECT 12.040 193.640 12.360 193.960 ;
        RECT 12.440 193.640 12.760 193.960 ;
        RECT 12.840 193.640 13.160 193.960 ;
        RECT 13.240 193.640 13.560 193.960 ;
        RECT 13.640 193.640 13.960 193.960 ;
        RECT 14.040 193.640 14.360 193.960 ;
        RECT 14.440 193.640 14.760 193.960 ;
        RECT 14.840 193.640 15.160 193.960 ;
        RECT 15.240 193.640 15.560 193.960 ;
        RECT 15.640 193.640 15.960 193.960 ;
        RECT 16.040 193.640 16.360 193.960 ;
        RECT 16.440 193.640 16.760 193.960 ;
        RECT 16.840 193.640 17.160 193.960 ;
        RECT 17.240 193.640 17.560 193.960 ;
        RECT 17.640 193.640 17.960 193.960 ;
        RECT 18.040 193.640 18.360 193.960 ;
        RECT 18.440 193.640 18.760 193.960 ;
        RECT 18.840 193.640 19.160 193.960 ;
        RECT 19.240 193.640 19.560 193.960 ;
        RECT 19.640 193.640 19.960 193.960 ;
        RECT 95.560 193.640 95.880 193.960 ;
        RECT 95.960 193.640 96.280 193.960 ;
        RECT 96.360 193.640 96.680 193.960 ;
        RECT 96.760 193.640 97.080 193.960 ;
        RECT 145.560 193.640 145.880 193.960 ;
        RECT 145.960 193.640 146.280 193.960 ;
        RECT 146.360 193.640 146.680 193.960 ;
        RECT 146.760 193.640 147.080 193.960 ;
        RECT 185.720 193.640 186.040 193.960 ;
        RECT 186.120 193.640 186.440 193.960 ;
        RECT 186.520 193.640 186.840 193.960 ;
        RECT 186.920 193.640 187.240 193.960 ;
        RECT 187.320 193.640 187.640 193.960 ;
        RECT 187.720 193.640 188.040 193.960 ;
        RECT 188.120 193.640 188.440 193.960 ;
        RECT 188.520 193.640 188.840 193.960 ;
        RECT 188.920 193.640 189.240 193.960 ;
        RECT 189.320 193.640 189.640 193.960 ;
        RECT 189.720 193.640 190.040 193.960 ;
        RECT 190.120 193.640 190.440 193.960 ;
        RECT 190.520 193.640 190.840 193.960 ;
        RECT 190.920 193.640 191.240 193.960 ;
        RECT 191.320 193.640 191.640 193.960 ;
        RECT 191.720 193.640 192.040 193.960 ;
        RECT 192.120 193.640 192.440 193.960 ;
        RECT 192.520 193.640 192.840 193.960 ;
        RECT 192.920 193.640 193.240 193.960 ;
        RECT 193.320 193.640 193.640 193.960 ;
        RECT 193.720 193.640 194.040 193.960 ;
        RECT 194.120 193.640 194.440 193.960 ;
        RECT 194.520 193.640 194.840 193.960 ;
        RECT 194.920 193.640 195.240 193.960 ;
        RECT 195.320 193.640 195.640 193.960 ;
        RECT 195.720 193.640 196.040 193.960 ;
        RECT 196.120 193.640 196.440 193.960 ;
        RECT 196.520 193.640 196.840 193.960 ;
        RECT 196.920 193.640 197.240 193.960 ;
        RECT 197.320 193.640 197.640 193.960 ;
        RECT 197.720 193.640 198.040 193.960 ;
        RECT 198.120 193.640 198.440 193.960 ;
        RECT 198.520 193.640 198.840 193.960 ;
        RECT 198.920 193.640 199.240 193.960 ;
        RECT 199.320 193.640 199.640 193.960 ;
        RECT 199.720 193.640 200.040 193.960 ;
        RECT 200.120 193.640 200.440 193.960 ;
        RECT 200.520 193.640 200.840 193.960 ;
        RECT 200.920 193.640 201.240 193.960 ;
        RECT 201.320 193.640 201.640 193.960 ;
        RECT 201.720 193.640 202.040 193.960 ;
        RECT 202.120 193.640 202.440 193.960 ;
        RECT 202.520 193.640 202.840 193.960 ;
        RECT 202.920 193.640 203.240 193.960 ;
        RECT 203.320 193.640 203.640 193.960 ;
        RECT 203.720 193.640 204.040 193.960 ;
        RECT 204.120 193.640 204.440 193.960 ;
        RECT 204.520 193.640 204.840 193.960 ;
        RECT 204.920 193.640 205.240 193.960 ;
        RECT 205.320 193.640 205.640 193.960 ;
        RECT 0.040 193.240 0.360 193.560 ;
        RECT 0.440 193.240 0.760 193.560 ;
        RECT 0.840 193.240 1.160 193.560 ;
        RECT 1.240 193.240 1.560 193.560 ;
        RECT 1.640 193.240 1.960 193.560 ;
        RECT 2.040 193.240 2.360 193.560 ;
        RECT 2.440 193.240 2.760 193.560 ;
        RECT 2.840 193.240 3.160 193.560 ;
        RECT 3.240 193.240 3.560 193.560 ;
        RECT 3.640 193.240 3.960 193.560 ;
        RECT 4.040 193.240 4.360 193.560 ;
        RECT 4.440 193.240 4.760 193.560 ;
        RECT 4.840 193.240 5.160 193.560 ;
        RECT 5.240 193.240 5.560 193.560 ;
        RECT 5.640 193.240 5.960 193.560 ;
        RECT 6.040 193.240 6.360 193.560 ;
        RECT 6.440 193.240 6.760 193.560 ;
        RECT 6.840 193.240 7.160 193.560 ;
        RECT 7.240 193.240 7.560 193.560 ;
        RECT 7.640 193.240 7.960 193.560 ;
        RECT 8.040 193.240 8.360 193.560 ;
        RECT 8.440 193.240 8.760 193.560 ;
        RECT 8.840 193.240 9.160 193.560 ;
        RECT 9.240 193.240 9.560 193.560 ;
        RECT 9.640 193.240 9.960 193.560 ;
        RECT 10.040 193.240 10.360 193.560 ;
        RECT 10.440 193.240 10.760 193.560 ;
        RECT 10.840 193.240 11.160 193.560 ;
        RECT 11.240 193.240 11.560 193.560 ;
        RECT 11.640 193.240 11.960 193.560 ;
        RECT 12.040 193.240 12.360 193.560 ;
        RECT 12.440 193.240 12.760 193.560 ;
        RECT 12.840 193.240 13.160 193.560 ;
        RECT 13.240 193.240 13.560 193.560 ;
        RECT 13.640 193.240 13.960 193.560 ;
        RECT 14.040 193.240 14.360 193.560 ;
        RECT 14.440 193.240 14.760 193.560 ;
        RECT 14.840 193.240 15.160 193.560 ;
        RECT 15.240 193.240 15.560 193.560 ;
        RECT 15.640 193.240 15.960 193.560 ;
        RECT 16.040 193.240 16.360 193.560 ;
        RECT 16.440 193.240 16.760 193.560 ;
        RECT 16.840 193.240 17.160 193.560 ;
        RECT 17.240 193.240 17.560 193.560 ;
        RECT 17.640 193.240 17.960 193.560 ;
        RECT 18.040 193.240 18.360 193.560 ;
        RECT 18.440 193.240 18.760 193.560 ;
        RECT 18.840 193.240 19.160 193.560 ;
        RECT 19.240 193.240 19.560 193.560 ;
        RECT 19.640 193.240 19.960 193.560 ;
        RECT 95.560 193.240 95.880 193.560 ;
        RECT 95.960 193.240 96.280 193.560 ;
        RECT 96.360 193.240 96.680 193.560 ;
        RECT 96.760 193.240 97.080 193.560 ;
        RECT 145.560 193.240 145.880 193.560 ;
        RECT 145.960 193.240 146.280 193.560 ;
        RECT 146.360 193.240 146.680 193.560 ;
        RECT 146.760 193.240 147.080 193.560 ;
        RECT 185.720 193.240 186.040 193.560 ;
        RECT 186.120 193.240 186.440 193.560 ;
        RECT 186.520 193.240 186.840 193.560 ;
        RECT 186.920 193.240 187.240 193.560 ;
        RECT 187.320 193.240 187.640 193.560 ;
        RECT 187.720 193.240 188.040 193.560 ;
        RECT 188.120 193.240 188.440 193.560 ;
        RECT 188.520 193.240 188.840 193.560 ;
        RECT 188.920 193.240 189.240 193.560 ;
        RECT 189.320 193.240 189.640 193.560 ;
        RECT 189.720 193.240 190.040 193.560 ;
        RECT 190.120 193.240 190.440 193.560 ;
        RECT 190.520 193.240 190.840 193.560 ;
        RECT 190.920 193.240 191.240 193.560 ;
        RECT 191.320 193.240 191.640 193.560 ;
        RECT 191.720 193.240 192.040 193.560 ;
        RECT 192.120 193.240 192.440 193.560 ;
        RECT 192.520 193.240 192.840 193.560 ;
        RECT 192.920 193.240 193.240 193.560 ;
        RECT 193.320 193.240 193.640 193.560 ;
        RECT 193.720 193.240 194.040 193.560 ;
        RECT 194.120 193.240 194.440 193.560 ;
        RECT 194.520 193.240 194.840 193.560 ;
        RECT 194.920 193.240 195.240 193.560 ;
        RECT 195.320 193.240 195.640 193.560 ;
        RECT 195.720 193.240 196.040 193.560 ;
        RECT 196.120 193.240 196.440 193.560 ;
        RECT 196.520 193.240 196.840 193.560 ;
        RECT 196.920 193.240 197.240 193.560 ;
        RECT 197.320 193.240 197.640 193.560 ;
        RECT 197.720 193.240 198.040 193.560 ;
        RECT 198.120 193.240 198.440 193.560 ;
        RECT 198.520 193.240 198.840 193.560 ;
        RECT 198.920 193.240 199.240 193.560 ;
        RECT 199.320 193.240 199.640 193.560 ;
        RECT 199.720 193.240 200.040 193.560 ;
        RECT 200.120 193.240 200.440 193.560 ;
        RECT 200.520 193.240 200.840 193.560 ;
        RECT 200.920 193.240 201.240 193.560 ;
        RECT 201.320 193.240 201.640 193.560 ;
        RECT 201.720 193.240 202.040 193.560 ;
        RECT 202.120 193.240 202.440 193.560 ;
        RECT 202.520 193.240 202.840 193.560 ;
        RECT 202.920 193.240 203.240 193.560 ;
        RECT 203.320 193.240 203.640 193.560 ;
        RECT 203.720 193.240 204.040 193.560 ;
        RECT 204.120 193.240 204.440 193.560 ;
        RECT 204.520 193.240 204.840 193.560 ;
        RECT 204.920 193.240 205.240 193.560 ;
        RECT 205.320 193.240 205.640 193.560 ;
        RECT 0.040 192.840 0.360 193.160 ;
        RECT 0.440 192.840 0.760 193.160 ;
        RECT 0.840 192.840 1.160 193.160 ;
        RECT 1.240 192.840 1.560 193.160 ;
        RECT 1.640 192.840 1.960 193.160 ;
        RECT 2.040 192.840 2.360 193.160 ;
        RECT 2.440 192.840 2.760 193.160 ;
        RECT 2.840 192.840 3.160 193.160 ;
        RECT 3.240 192.840 3.560 193.160 ;
        RECT 3.640 192.840 3.960 193.160 ;
        RECT 4.040 192.840 4.360 193.160 ;
        RECT 4.440 192.840 4.760 193.160 ;
        RECT 4.840 192.840 5.160 193.160 ;
        RECT 5.240 192.840 5.560 193.160 ;
        RECT 5.640 192.840 5.960 193.160 ;
        RECT 6.040 192.840 6.360 193.160 ;
        RECT 6.440 192.840 6.760 193.160 ;
        RECT 6.840 192.840 7.160 193.160 ;
        RECT 7.240 192.840 7.560 193.160 ;
        RECT 7.640 192.840 7.960 193.160 ;
        RECT 8.040 192.840 8.360 193.160 ;
        RECT 8.440 192.840 8.760 193.160 ;
        RECT 8.840 192.840 9.160 193.160 ;
        RECT 9.240 192.840 9.560 193.160 ;
        RECT 9.640 192.840 9.960 193.160 ;
        RECT 10.040 192.840 10.360 193.160 ;
        RECT 10.440 192.840 10.760 193.160 ;
        RECT 10.840 192.840 11.160 193.160 ;
        RECT 11.240 192.840 11.560 193.160 ;
        RECT 11.640 192.840 11.960 193.160 ;
        RECT 12.040 192.840 12.360 193.160 ;
        RECT 12.440 192.840 12.760 193.160 ;
        RECT 12.840 192.840 13.160 193.160 ;
        RECT 13.240 192.840 13.560 193.160 ;
        RECT 13.640 192.840 13.960 193.160 ;
        RECT 14.040 192.840 14.360 193.160 ;
        RECT 14.440 192.840 14.760 193.160 ;
        RECT 14.840 192.840 15.160 193.160 ;
        RECT 15.240 192.840 15.560 193.160 ;
        RECT 15.640 192.840 15.960 193.160 ;
        RECT 16.040 192.840 16.360 193.160 ;
        RECT 16.440 192.840 16.760 193.160 ;
        RECT 16.840 192.840 17.160 193.160 ;
        RECT 17.240 192.840 17.560 193.160 ;
        RECT 17.640 192.840 17.960 193.160 ;
        RECT 18.040 192.840 18.360 193.160 ;
        RECT 18.440 192.840 18.760 193.160 ;
        RECT 18.840 192.840 19.160 193.160 ;
        RECT 19.240 192.840 19.560 193.160 ;
        RECT 19.640 192.840 19.960 193.160 ;
        RECT 95.560 192.840 95.880 193.160 ;
        RECT 95.960 192.840 96.280 193.160 ;
        RECT 96.360 192.840 96.680 193.160 ;
        RECT 96.760 192.840 97.080 193.160 ;
        RECT 145.560 192.840 145.880 193.160 ;
        RECT 145.960 192.840 146.280 193.160 ;
        RECT 146.360 192.840 146.680 193.160 ;
        RECT 146.760 192.840 147.080 193.160 ;
        RECT 185.720 192.840 186.040 193.160 ;
        RECT 186.120 192.840 186.440 193.160 ;
        RECT 186.520 192.840 186.840 193.160 ;
        RECT 186.920 192.840 187.240 193.160 ;
        RECT 187.320 192.840 187.640 193.160 ;
        RECT 187.720 192.840 188.040 193.160 ;
        RECT 188.120 192.840 188.440 193.160 ;
        RECT 188.520 192.840 188.840 193.160 ;
        RECT 188.920 192.840 189.240 193.160 ;
        RECT 189.320 192.840 189.640 193.160 ;
        RECT 189.720 192.840 190.040 193.160 ;
        RECT 190.120 192.840 190.440 193.160 ;
        RECT 190.520 192.840 190.840 193.160 ;
        RECT 190.920 192.840 191.240 193.160 ;
        RECT 191.320 192.840 191.640 193.160 ;
        RECT 191.720 192.840 192.040 193.160 ;
        RECT 192.120 192.840 192.440 193.160 ;
        RECT 192.520 192.840 192.840 193.160 ;
        RECT 192.920 192.840 193.240 193.160 ;
        RECT 193.320 192.840 193.640 193.160 ;
        RECT 193.720 192.840 194.040 193.160 ;
        RECT 194.120 192.840 194.440 193.160 ;
        RECT 194.520 192.840 194.840 193.160 ;
        RECT 194.920 192.840 195.240 193.160 ;
        RECT 195.320 192.840 195.640 193.160 ;
        RECT 195.720 192.840 196.040 193.160 ;
        RECT 196.120 192.840 196.440 193.160 ;
        RECT 196.520 192.840 196.840 193.160 ;
        RECT 196.920 192.840 197.240 193.160 ;
        RECT 197.320 192.840 197.640 193.160 ;
        RECT 197.720 192.840 198.040 193.160 ;
        RECT 198.120 192.840 198.440 193.160 ;
        RECT 198.520 192.840 198.840 193.160 ;
        RECT 198.920 192.840 199.240 193.160 ;
        RECT 199.320 192.840 199.640 193.160 ;
        RECT 199.720 192.840 200.040 193.160 ;
        RECT 200.120 192.840 200.440 193.160 ;
        RECT 200.520 192.840 200.840 193.160 ;
        RECT 200.920 192.840 201.240 193.160 ;
        RECT 201.320 192.840 201.640 193.160 ;
        RECT 201.720 192.840 202.040 193.160 ;
        RECT 202.120 192.840 202.440 193.160 ;
        RECT 202.520 192.840 202.840 193.160 ;
        RECT 202.920 192.840 203.240 193.160 ;
        RECT 203.320 192.840 203.640 193.160 ;
        RECT 203.720 192.840 204.040 193.160 ;
        RECT 204.120 192.840 204.440 193.160 ;
        RECT 204.520 192.840 204.840 193.160 ;
        RECT 204.920 192.840 205.240 193.160 ;
        RECT 205.320 192.840 205.640 193.160 ;
        RECT 0.040 192.440 0.360 192.760 ;
        RECT 0.440 192.440 0.760 192.760 ;
        RECT 0.840 192.440 1.160 192.760 ;
        RECT 1.240 192.440 1.560 192.760 ;
        RECT 1.640 192.440 1.960 192.760 ;
        RECT 2.040 192.440 2.360 192.760 ;
        RECT 2.440 192.440 2.760 192.760 ;
        RECT 2.840 192.440 3.160 192.760 ;
        RECT 3.240 192.440 3.560 192.760 ;
        RECT 3.640 192.440 3.960 192.760 ;
        RECT 4.040 192.440 4.360 192.760 ;
        RECT 4.440 192.440 4.760 192.760 ;
        RECT 4.840 192.440 5.160 192.760 ;
        RECT 5.240 192.440 5.560 192.760 ;
        RECT 5.640 192.440 5.960 192.760 ;
        RECT 6.040 192.440 6.360 192.760 ;
        RECT 6.440 192.440 6.760 192.760 ;
        RECT 6.840 192.440 7.160 192.760 ;
        RECT 7.240 192.440 7.560 192.760 ;
        RECT 7.640 192.440 7.960 192.760 ;
        RECT 8.040 192.440 8.360 192.760 ;
        RECT 8.440 192.440 8.760 192.760 ;
        RECT 8.840 192.440 9.160 192.760 ;
        RECT 9.240 192.440 9.560 192.760 ;
        RECT 9.640 192.440 9.960 192.760 ;
        RECT 10.040 192.440 10.360 192.760 ;
        RECT 10.440 192.440 10.760 192.760 ;
        RECT 10.840 192.440 11.160 192.760 ;
        RECT 11.240 192.440 11.560 192.760 ;
        RECT 11.640 192.440 11.960 192.760 ;
        RECT 12.040 192.440 12.360 192.760 ;
        RECT 12.440 192.440 12.760 192.760 ;
        RECT 12.840 192.440 13.160 192.760 ;
        RECT 13.240 192.440 13.560 192.760 ;
        RECT 13.640 192.440 13.960 192.760 ;
        RECT 14.040 192.440 14.360 192.760 ;
        RECT 14.440 192.440 14.760 192.760 ;
        RECT 14.840 192.440 15.160 192.760 ;
        RECT 15.240 192.440 15.560 192.760 ;
        RECT 15.640 192.440 15.960 192.760 ;
        RECT 16.040 192.440 16.360 192.760 ;
        RECT 16.440 192.440 16.760 192.760 ;
        RECT 16.840 192.440 17.160 192.760 ;
        RECT 17.240 192.440 17.560 192.760 ;
        RECT 17.640 192.440 17.960 192.760 ;
        RECT 18.040 192.440 18.360 192.760 ;
        RECT 18.440 192.440 18.760 192.760 ;
        RECT 18.840 192.440 19.160 192.760 ;
        RECT 19.240 192.440 19.560 192.760 ;
        RECT 19.640 192.440 19.960 192.760 ;
        RECT 95.560 192.440 95.880 192.760 ;
        RECT 95.960 192.440 96.280 192.760 ;
        RECT 96.360 192.440 96.680 192.760 ;
        RECT 96.760 192.440 97.080 192.760 ;
        RECT 145.560 192.440 145.880 192.760 ;
        RECT 145.960 192.440 146.280 192.760 ;
        RECT 146.360 192.440 146.680 192.760 ;
        RECT 146.760 192.440 147.080 192.760 ;
        RECT 185.720 192.440 186.040 192.760 ;
        RECT 186.120 192.440 186.440 192.760 ;
        RECT 186.520 192.440 186.840 192.760 ;
        RECT 186.920 192.440 187.240 192.760 ;
        RECT 187.320 192.440 187.640 192.760 ;
        RECT 187.720 192.440 188.040 192.760 ;
        RECT 188.120 192.440 188.440 192.760 ;
        RECT 188.520 192.440 188.840 192.760 ;
        RECT 188.920 192.440 189.240 192.760 ;
        RECT 189.320 192.440 189.640 192.760 ;
        RECT 189.720 192.440 190.040 192.760 ;
        RECT 190.120 192.440 190.440 192.760 ;
        RECT 190.520 192.440 190.840 192.760 ;
        RECT 190.920 192.440 191.240 192.760 ;
        RECT 191.320 192.440 191.640 192.760 ;
        RECT 191.720 192.440 192.040 192.760 ;
        RECT 192.120 192.440 192.440 192.760 ;
        RECT 192.520 192.440 192.840 192.760 ;
        RECT 192.920 192.440 193.240 192.760 ;
        RECT 193.320 192.440 193.640 192.760 ;
        RECT 193.720 192.440 194.040 192.760 ;
        RECT 194.120 192.440 194.440 192.760 ;
        RECT 194.520 192.440 194.840 192.760 ;
        RECT 194.920 192.440 195.240 192.760 ;
        RECT 195.320 192.440 195.640 192.760 ;
        RECT 195.720 192.440 196.040 192.760 ;
        RECT 196.120 192.440 196.440 192.760 ;
        RECT 196.520 192.440 196.840 192.760 ;
        RECT 196.920 192.440 197.240 192.760 ;
        RECT 197.320 192.440 197.640 192.760 ;
        RECT 197.720 192.440 198.040 192.760 ;
        RECT 198.120 192.440 198.440 192.760 ;
        RECT 198.520 192.440 198.840 192.760 ;
        RECT 198.920 192.440 199.240 192.760 ;
        RECT 199.320 192.440 199.640 192.760 ;
        RECT 199.720 192.440 200.040 192.760 ;
        RECT 200.120 192.440 200.440 192.760 ;
        RECT 200.520 192.440 200.840 192.760 ;
        RECT 200.920 192.440 201.240 192.760 ;
        RECT 201.320 192.440 201.640 192.760 ;
        RECT 201.720 192.440 202.040 192.760 ;
        RECT 202.120 192.440 202.440 192.760 ;
        RECT 202.520 192.440 202.840 192.760 ;
        RECT 202.920 192.440 203.240 192.760 ;
        RECT 203.320 192.440 203.640 192.760 ;
        RECT 203.720 192.440 204.040 192.760 ;
        RECT 204.120 192.440 204.440 192.760 ;
        RECT 204.520 192.440 204.840 192.760 ;
        RECT 204.920 192.440 205.240 192.760 ;
        RECT 205.320 192.440 205.640 192.760 ;
        RECT 0.040 192.040 0.360 192.360 ;
        RECT 0.440 192.040 0.760 192.360 ;
        RECT 0.840 192.040 1.160 192.360 ;
        RECT 1.240 192.040 1.560 192.360 ;
        RECT 1.640 192.040 1.960 192.360 ;
        RECT 2.040 192.040 2.360 192.360 ;
        RECT 2.440 192.040 2.760 192.360 ;
        RECT 2.840 192.040 3.160 192.360 ;
        RECT 3.240 192.040 3.560 192.360 ;
        RECT 3.640 192.040 3.960 192.360 ;
        RECT 4.040 192.040 4.360 192.360 ;
        RECT 4.440 192.040 4.760 192.360 ;
        RECT 4.840 192.040 5.160 192.360 ;
        RECT 5.240 192.040 5.560 192.360 ;
        RECT 5.640 192.040 5.960 192.360 ;
        RECT 6.040 192.040 6.360 192.360 ;
        RECT 6.440 192.040 6.760 192.360 ;
        RECT 6.840 192.040 7.160 192.360 ;
        RECT 7.240 192.040 7.560 192.360 ;
        RECT 7.640 192.040 7.960 192.360 ;
        RECT 8.040 192.040 8.360 192.360 ;
        RECT 8.440 192.040 8.760 192.360 ;
        RECT 8.840 192.040 9.160 192.360 ;
        RECT 9.240 192.040 9.560 192.360 ;
        RECT 9.640 192.040 9.960 192.360 ;
        RECT 10.040 192.040 10.360 192.360 ;
        RECT 10.440 192.040 10.760 192.360 ;
        RECT 10.840 192.040 11.160 192.360 ;
        RECT 11.240 192.040 11.560 192.360 ;
        RECT 11.640 192.040 11.960 192.360 ;
        RECT 12.040 192.040 12.360 192.360 ;
        RECT 12.440 192.040 12.760 192.360 ;
        RECT 12.840 192.040 13.160 192.360 ;
        RECT 13.240 192.040 13.560 192.360 ;
        RECT 13.640 192.040 13.960 192.360 ;
        RECT 14.040 192.040 14.360 192.360 ;
        RECT 14.440 192.040 14.760 192.360 ;
        RECT 14.840 192.040 15.160 192.360 ;
        RECT 15.240 192.040 15.560 192.360 ;
        RECT 15.640 192.040 15.960 192.360 ;
        RECT 16.040 192.040 16.360 192.360 ;
        RECT 16.440 192.040 16.760 192.360 ;
        RECT 16.840 192.040 17.160 192.360 ;
        RECT 17.240 192.040 17.560 192.360 ;
        RECT 17.640 192.040 17.960 192.360 ;
        RECT 18.040 192.040 18.360 192.360 ;
        RECT 18.440 192.040 18.760 192.360 ;
        RECT 18.840 192.040 19.160 192.360 ;
        RECT 19.240 192.040 19.560 192.360 ;
        RECT 19.640 192.040 19.960 192.360 ;
        RECT 95.560 192.040 95.880 192.360 ;
        RECT 95.960 192.040 96.280 192.360 ;
        RECT 96.360 192.040 96.680 192.360 ;
        RECT 96.760 192.040 97.080 192.360 ;
        RECT 145.560 192.040 145.880 192.360 ;
        RECT 145.960 192.040 146.280 192.360 ;
        RECT 146.360 192.040 146.680 192.360 ;
        RECT 146.760 192.040 147.080 192.360 ;
        RECT 185.720 192.040 186.040 192.360 ;
        RECT 186.120 192.040 186.440 192.360 ;
        RECT 186.520 192.040 186.840 192.360 ;
        RECT 186.920 192.040 187.240 192.360 ;
        RECT 187.320 192.040 187.640 192.360 ;
        RECT 187.720 192.040 188.040 192.360 ;
        RECT 188.120 192.040 188.440 192.360 ;
        RECT 188.520 192.040 188.840 192.360 ;
        RECT 188.920 192.040 189.240 192.360 ;
        RECT 189.320 192.040 189.640 192.360 ;
        RECT 189.720 192.040 190.040 192.360 ;
        RECT 190.120 192.040 190.440 192.360 ;
        RECT 190.520 192.040 190.840 192.360 ;
        RECT 190.920 192.040 191.240 192.360 ;
        RECT 191.320 192.040 191.640 192.360 ;
        RECT 191.720 192.040 192.040 192.360 ;
        RECT 192.120 192.040 192.440 192.360 ;
        RECT 192.520 192.040 192.840 192.360 ;
        RECT 192.920 192.040 193.240 192.360 ;
        RECT 193.320 192.040 193.640 192.360 ;
        RECT 193.720 192.040 194.040 192.360 ;
        RECT 194.120 192.040 194.440 192.360 ;
        RECT 194.520 192.040 194.840 192.360 ;
        RECT 194.920 192.040 195.240 192.360 ;
        RECT 195.320 192.040 195.640 192.360 ;
        RECT 195.720 192.040 196.040 192.360 ;
        RECT 196.120 192.040 196.440 192.360 ;
        RECT 196.520 192.040 196.840 192.360 ;
        RECT 196.920 192.040 197.240 192.360 ;
        RECT 197.320 192.040 197.640 192.360 ;
        RECT 197.720 192.040 198.040 192.360 ;
        RECT 198.120 192.040 198.440 192.360 ;
        RECT 198.520 192.040 198.840 192.360 ;
        RECT 198.920 192.040 199.240 192.360 ;
        RECT 199.320 192.040 199.640 192.360 ;
        RECT 199.720 192.040 200.040 192.360 ;
        RECT 200.120 192.040 200.440 192.360 ;
        RECT 200.520 192.040 200.840 192.360 ;
        RECT 200.920 192.040 201.240 192.360 ;
        RECT 201.320 192.040 201.640 192.360 ;
        RECT 201.720 192.040 202.040 192.360 ;
        RECT 202.120 192.040 202.440 192.360 ;
        RECT 202.520 192.040 202.840 192.360 ;
        RECT 202.920 192.040 203.240 192.360 ;
        RECT 203.320 192.040 203.640 192.360 ;
        RECT 203.720 192.040 204.040 192.360 ;
        RECT 204.120 192.040 204.440 192.360 ;
        RECT 204.520 192.040 204.840 192.360 ;
        RECT 204.920 192.040 205.240 192.360 ;
        RECT 205.320 192.040 205.640 192.360 ;
        RECT 0.040 191.640 0.360 191.960 ;
        RECT 0.440 191.640 0.760 191.960 ;
        RECT 0.840 191.640 1.160 191.960 ;
        RECT 1.240 191.640 1.560 191.960 ;
        RECT 1.640 191.640 1.960 191.960 ;
        RECT 2.040 191.640 2.360 191.960 ;
        RECT 2.440 191.640 2.760 191.960 ;
        RECT 2.840 191.640 3.160 191.960 ;
        RECT 3.240 191.640 3.560 191.960 ;
        RECT 3.640 191.640 3.960 191.960 ;
        RECT 4.040 191.640 4.360 191.960 ;
        RECT 4.440 191.640 4.760 191.960 ;
        RECT 4.840 191.640 5.160 191.960 ;
        RECT 5.240 191.640 5.560 191.960 ;
        RECT 5.640 191.640 5.960 191.960 ;
        RECT 6.040 191.640 6.360 191.960 ;
        RECT 6.440 191.640 6.760 191.960 ;
        RECT 6.840 191.640 7.160 191.960 ;
        RECT 7.240 191.640 7.560 191.960 ;
        RECT 7.640 191.640 7.960 191.960 ;
        RECT 8.040 191.640 8.360 191.960 ;
        RECT 8.440 191.640 8.760 191.960 ;
        RECT 8.840 191.640 9.160 191.960 ;
        RECT 9.240 191.640 9.560 191.960 ;
        RECT 9.640 191.640 9.960 191.960 ;
        RECT 10.040 191.640 10.360 191.960 ;
        RECT 10.440 191.640 10.760 191.960 ;
        RECT 10.840 191.640 11.160 191.960 ;
        RECT 11.240 191.640 11.560 191.960 ;
        RECT 11.640 191.640 11.960 191.960 ;
        RECT 12.040 191.640 12.360 191.960 ;
        RECT 12.440 191.640 12.760 191.960 ;
        RECT 12.840 191.640 13.160 191.960 ;
        RECT 13.240 191.640 13.560 191.960 ;
        RECT 13.640 191.640 13.960 191.960 ;
        RECT 14.040 191.640 14.360 191.960 ;
        RECT 14.440 191.640 14.760 191.960 ;
        RECT 14.840 191.640 15.160 191.960 ;
        RECT 15.240 191.640 15.560 191.960 ;
        RECT 15.640 191.640 15.960 191.960 ;
        RECT 16.040 191.640 16.360 191.960 ;
        RECT 16.440 191.640 16.760 191.960 ;
        RECT 16.840 191.640 17.160 191.960 ;
        RECT 17.240 191.640 17.560 191.960 ;
        RECT 17.640 191.640 17.960 191.960 ;
        RECT 18.040 191.640 18.360 191.960 ;
        RECT 18.440 191.640 18.760 191.960 ;
        RECT 18.840 191.640 19.160 191.960 ;
        RECT 19.240 191.640 19.560 191.960 ;
        RECT 19.640 191.640 19.960 191.960 ;
        RECT 95.560 191.640 95.880 191.960 ;
        RECT 95.960 191.640 96.280 191.960 ;
        RECT 96.360 191.640 96.680 191.960 ;
        RECT 96.760 191.640 97.080 191.960 ;
        RECT 145.560 191.640 145.880 191.960 ;
        RECT 145.960 191.640 146.280 191.960 ;
        RECT 146.360 191.640 146.680 191.960 ;
        RECT 146.760 191.640 147.080 191.960 ;
        RECT 185.720 191.640 186.040 191.960 ;
        RECT 186.120 191.640 186.440 191.960 ;
        RECT 186.520 191.640 186.840 191.960 ;
        RECT 186.920 191.640 187.240 191.960 ;
        RECT 187.320 191.640 187.640 191.960 ;
        RECT 187.720 191.640 188.040 191.960 ;
        RECT 188.120 191.640 188.440 191.960 ;
        RECT 188.520 191.640 188.840 191.960 ;
        RECT 188.920 191.640 189.240 191.960 ;
        RECT 189.320 191.640 189.640 191.960 ;
        RECT 189.720 191.640 190.040 191.960 ;
        RECT 190.120 191.640 190.440 191.960 ;
        RECT 190.520 191.640 190.840 191.960 ;
        RECT 190.920 191.640 191.240 191.960 ;
        RECT 191.320 191.640 191.640 191.960 ;
        RECT 191.720 191.640 192.040 191.960 ;
        RECT 192.120 191.640 192.440 191.960 ;
        RECT 192.520 191.640 192.840 191.960 ;
        RECT 192.920 191.640 193.240 191.960 ;
        RECT 193.320 191.640 193.640 191.960 ;
        RECT 193.720 191.640 194.040 191.960 ;
        RECT 194.120 191.640 194.440 191.960 ;
        RECT 194.520 191.640 194.840 191.960 ;
        RECT 194.920 191.640 195.240 191.960 ;
        RECT 195.320 191.640 195.640 191.960 ;
        RECT 195.720 191.640 196.040 191.960 ;
        RECT 196.120 191.640 196.440 191.960 ;
        RECT 196.520 191.640 196.840 191.960 ;
        RECT 196.920 191.640 197.240 191.960 ;
        RECT 197.320 191.640 197.640 191.960 ;
        RECT 197.720 191.640 198.040 191.960 ;
        RECT 198.120 191.640 198.440 191.960 ;
        RECT 198.520 191.640 198.840 191.960 ;
        RECT 198.920 191.640 199.240 191.960 ;
        RECT 199.320 191.640 199.640 191.960 ;
        RECT 199.720 191.640 200.040 191.960 ;
        RECT 200.120 191.640 200.440 191.960 ;
        RECT 200.520 191.640 200.840 191.960 ;
        RECT 200.920 191.640 201.240 191.960 ;
        RECT 201.320 191.640 201.640 191.960 ;
        RECT 201.720 191.640 202.040 191.960 ;
        RECT 202.120 191.640 202.440 191.960 ;
        RECT 202.520 191.640 202.840 191.960 ;
        RECT 202.920 191.640 203.240 191.960 ;
        RECT 203.320 191.640 203.640 191.960 ;
        RECT 203.720 191.640 204.040 191.960 ;
        RECT 204.120 191.640 204.440 191.960 ;
        RECT 204.520 191.640 204.840 191.960 ;
        RECT 204.920 191.640 205.240 191.960 ;
        RECT 205.320 191.640 205.640 191.960 ;
        RECT 0.040 191.240 0.360 191.560 ;
        RECT 0.440 191.240 0.760 191.560 ;
        RECT 0.840 191.240 1.160 191.560 ;
        RECT 1.240 191.240 1.560 191.560 ;
        RECT 1.640 191.240 1.960 191.560 ;
        RECT 2.040 191.240 2.360 191.560 ;
        RECT 2.440 191.240 2.760 191.560 ;
        RECT 2.840 191.240 3.160 191.560 ;
        RECT 3.240 191.240 3.560 191.560 ;
        RECT 3.640 191.240 3.960 191.560 ;
        RECT 4.040 191.240 4.360 191.560 ;
        RECT 4.440 191.240 4.760 191.560 ;
        RECT 4.840 191.240 5.160 191.560 ;
        RECT 5.240 191.240 5.560 191.560 ;
        RECT 5.640 191.240 5.960 191.560 ;
        RECT 6.040 191.240 6.360 191.560 ;
        RECT 6.440 191.240 6.760 191.560 ;
        RECT 6.840 191.240 7.160 191.560 ;
        RECT 7.240 191.240 7.560 191.560 ;
        RECT 7.640 191.240 7.960 191.560 ;
        RECT 8.040 191.240 8.360 191.560 ;
        RECT 8.440 191.240 8.760 191.560 ;
        RECT 8.840 191.240 9.160 191.560 ;
        RECT 9.240 191.240 9.560 191.560 ;
        RECT 9.640 191.240 9.960 191.560 ;
        RECT 10.040 191.240 10.360 191.560 ;
        RECT 10.440 191.240 10.760 191.560 ;
        RECT 10.840 191.240 11.160 191.560 ;
        RECT 11.240 191.240 11.560 191.560 ;
        RECT 11.640 191.240 11.960 191.560 ;
        RECT 12.040 191.240 12.360 191.560 ;
        RECT 12.440 191.240 12.760 191.560 ;
        RECT 12.840 191.240 13.160 191.560 ;
        RECT 13.240 191.240 13.560 191.560 ;
        RECT 13.640 191.240 13.960 191.560 ;
        RECT 14.040 191.240 14.360 191.560 ;
        RECT 14.440 191.240 14.760 191.560 ;
        RECT 14.840 191.240 15.160 191.560 ;
        RECT 15.240 191.240 15.560 191.560 ;
        RECT 15.640 191.240 15.960 191.560 ;
        RECT 16.040 191.240 16.360 191.560 ;
        RECT 16.440 191.240 16.760 191.560 ;
        RECT 16.840 191.240 17.160 191.560 ;
        RECT 17.240 191.240 17.560 191.560 ;
        RECT 17.640 191.240 17.960 191.560 ;
        RECT 18.040 191.240 18.360 191.560 ;
        RECT 18.440 191.240 18.760 191.560 ;
        RECT 18.840 191.240 19.160 191.560 ;
        RECT 19.240 191.240 19.560 191.560 ;
        RECT 19.640 191.240 19.960 191.560 ;
        RECT 95.560 191.240 95.880 191.560 ;
        RECT 95.960 191.240 96.280 191.560 ;
        RECT 96.360 191.240 96.680 191.560 ;
        RECT 96.760 191.240 97.080 191.560 ;
        RECT 145.560 191.240 145.880 191.560 ;
        RECT 145.960 191.240 146.280 191.560 ;
        RECT 146.360 191.240 146.680 191.560 ;
        RECT 146.760 191.240 147.080 191.560 ;
        RECT 185.720 191.240 186.040 191.560 ;
        RECT 186.120 191.240 186.440 191.560 ;
        RECT 186.520 191.240 186.840 191.560 ;
        RECT 186.920 191.240 187.240 191.560 ;
        RECT 187.320 191.240 187.640 191.560 ;
        RECT 187.720 191.240 188.040 191.560 ;
        RECT 188.120 191.240 188.440 191.560 ;
        RECT 188.520 191.240 188.840 191.560 ;
        RECT 188.920 191.240 189.240 191.560 ;
        RECT 189.320 191.240 189.640 191.560 ;
        RECT 189.720 191.240 190.040 191.560 ;
        RECT 190.120 191.240 190.440 191.560 ;
        RECT 190.520 191.240 190.840 191.560 ;
        RECT 190.920 191.240 191.240 191.560 ;
        RECT 191.320 191.240 191.640 191.560 ;
        RECT 191.720 191.240 192.040 191.560 ;
        RECT 192.120 191.240 192.440 191.560 ;
        RECT 192.520 191.240 192.840 191.560 ;
        RECT 192.920 191.240 193.240 191.560 ;
        RECT 193.320 191.240 193.640 191.560 ;
        RECT 193.720 191.240 194.040 191.560 ;
        RECT 194.120 191.240 194.440 191.560 ;
        RECT 194.520 191.240 194.840 191.560 ;
        RECT 194.920 191.240 195.240 191.560 ;
        RECT 195.320 191.240 195.640 191.560 ;
        RECT 195.720 191.240 196.040 191.560 ;
        RECT 196.120 191.240 196.440 191.560 ;
        RECT 196.520 191.240 196.840 191.560 ;
        RECT 196.920 191.240 197.240 191.560 ;
        RECT 197.320 191.240 197.640 191.560 ;
        RECT 197.720 191.240 198.040 191.560 ;
        RECT 198.120 191.240 198.440 191.560 ;
        RECT 198.520 191.240 198.840 191.560 ;
        RECT 198.920 191.240 199.240 191.560 ;
        RECT 199.320 191.240 199.640 191.560 ;
        RECT 199.720 191.240 200.040 191.560 ;
        RECT 200.120 191.240 200.440 191.560 ;
        RECT 200.520 191.240 200.840 191.560 ;
        RECT 200.920 191.240 201.240 191.560 ;
        RECT 201.320 191.240 201.640 191.560 ;
        RECT 201.720 191.240 202.040 191.560 ;
        RECT 202.120 191.240 202.440 191.560 ;
        RECT 202.520 191.240 202.840 191.560 ;
        RECT 202.920 191.240 203.240 191.560 ;
        RECT 203.320 191.240 203.640 191.560 ;
        RECT 203.720 191.240 204.040 191.560 ;
        RECT 204.120 191.240 204.440 191.560 ;
        RECT 204.520 191.240 204.840 191.560 ;
        RECT 204.920 191.240 205.240 191.560 ;
        RECT 205.320 191.240 205.640 191.560 ;
        RECT 0.040 190.840 0.360 191.160 ;
        RECT 0.440 190.840 0.760 191.160 ;
        RECT 0.840 190.840 1.160 191.160 ;
        RECT 1.240 190.840 1.560 191.160 ;
        RECT 1.640 190.840 1.960 191.160 ;
        RECT 2.040 190.840 2.360 191.160 ;
        RECT 2.440 190.840 2.760 191.160 ;
        RECT 2.840 190.840 3.160 191.160 ;
        RECT 3.240 190.840 3.560 191.160 ;
        RECT 3.640 190.840 3.960 191.160 ;
        RECT 4.040 190.840 4.360 191.160 ;
        RECT 4.440 190.840 4.760 191.160 ;
        RECT 4.840 190.840 5.160 191.160 ;
        RECT 5.240 190.840 5.560 191.160 ;
        RECT 5.640 190.840 5.960 191.160 ;
        RECT 6.040 190.840 6.360 191.160 ;
        RECT 6.440 190.840 6.760 191.160 ;
        RECT 6.840 190.840 7.160 191.160 ;
        RECT 7.240 190.840 7.560 191.160 ;
        RECT 7.640 190.840 7.960 191.160 ;
        RECT 8.040 190.840 8.360 191.160 ;
        RECT 8.440 190.840 8.760 191.160 ;
        RECT 8.840 190.840 9.160 191.160 ;
        RECT 9.240 190.840 9.560 191.160 ;
        RECT 9.640 190.840 9.960 191.160 ;
        RECT 10.040 190.840 10.360 191.160 ;
        RECT 10.440 190.840 10.760 191.160 ;
        RECT 10.840 190.840 11.160 191.160 ;
        RECT 11.240 190.840 11.560 191.160 ;
        RECT 11.640 190.840 11.960 191.160 ;
        RECT 12.040 190.840 12.360 191.160 ;
        RECT 12.440 190.840 12.760 191.160 ;
        RECT 12.840 190.840 13.160 191.160 ;
        RECT 13.240 190.840 13.560 191.160 ;
        RECT 13.640 190.840 13.960 191.160 ;
        RECT 14.040 190.840 14.360 191.160 ;
        RECT 14.440 190.840 14.760 191.160 ;
        RECT 14.840 190.840 15.160 191.160 ;
        RECT 15.240 190.840 15.560 191.160 ;
        RECT 15.640 190.840 15.960 191.160 ;
        RECT 16.040 190.840 16.360 191.160 ;
        RECT 16.440 190.840 16.760 191.160 ;
        RECT 16.840 190.840 17.160 191.160 ;
        RECT 17.240 190.840 17.560 191.160 ;
        RECT 17.640 190.840 17.960 191.160 ;
        RECT 18.040 190.840 18.360 191.160 ;
        RECT 18.440 190.840 18.760 191.160 ;
        RECT 18.840 190.840 19.160 191.160 ;
        RECT 19.240 190.840 19.560 191.160 ;
        RECT 19.640 190.840 19.960 191.160 ;
        RECT 95.560 190.840 95.880 191.160 ;
        RECT 95.960 190.840 96.280 191.160 ;
        RECT 96.360 190.840 96.680 191.160 ;
        RECT 96.760 190.840 97.080 191.160 ;
        RECT 145.560 190.840 145.880 191.160 ;
        RECT 145.960 190.840 146.280 191.160 ;
        RECT 146.360 190.840 146.680 191.160 ;
        RECT 146.760 190.840 147.080 191.160 ;
        RECT 185.720 190.840 186.040 191.160 ;
        RECT 186.120 190.840 186.440 191.160 ;
        RECT 186.520 190.840 186.840 191.160 ;
        RECT 186.920 190.840 187.240 191.160 ;
        RECT 187.320 190.840 187.640 191.160 ;
        RECT 187.720 190.840 188.040 191.160 ;
        RECT 188.120 190.840 188.440 191.160 ;
        RECT 188.520 190.840 188.840 191.160 ;
        RECT 188.920 190.840 189.240 191.160 ;
        RECT 189.320 190.840 189.640 191.160 ;
        RECT 189.720 190.840 190.040 191.160 ;
        RECT 190.120 190.840 190.440 191.160 ;
        RECT 190.520 190.840 190.840 191.160 ;
        RECT 190.920 190.840 191.240 191.160 ;
        RECT 191.320 190.840 191.640 191.160 ;
        RECT 191.720 190.840 192.040 191.160 ;
        RECT 192.120 190.840 192.440 191.160 ;
        RECT 192.520 190.840 192.840 191.160 ;
        RECT 192.920 190.840 193.240 191.160 ;
        RECT 193.320 190.840 193.640 191.160 ;
        RECT 193.720 190.840 194.040 191.160 ;
        RECT 194.120 190.840 194.440 191.160 ;
        RECT 194.520 190.840 194.840 191.160 ;
        RECT 194.920 190.840 195.240 191.160 ;
        RECT 195.320 190.840 195.640 191.160 ;
        RECT 195.720 190.840 196.040 191.160 ;
        RECT 196.120 190.840 196.440 191.160 ;
        RECT 196.520 190.840 196.840 191.160 ;
        RECT 196.920 190.840 197.240 191.160 ;
        RECT 197.320 190.840 197.640 191.160 ;
        RECT 197.720 190.840 198.040 191.160 ;
        RECT 198.120 190.840 198.440 191.160 ;
        RECT 198.520 190.840 198.840 191.160 ;
        RECT 198.920 190.840 199.240 191.160 ;
        RECT 199.320 190.840 199.640 191.160 ;
        RECT 199.720 190.840 200.040 191.160 ;
        RECT 200.120 190.840 200.440 191.160 ;
        RECT 200.520 190.840 200.840 191.160 ;
        RECT 200.920 190.840 201.240 191.160 ;
        RECT 201.320 190.840 201.640 191.160 ;
        RECT 201.720 190.840 202.040 191.160 ;
        RECT 202.120 190.840 202.440 191.160 ;
        RECT 202.520 190.840 202.840 191.160 ;
        RECT 202.920 190.840 203.240 191.160 ;
        RECT 203.320 190.840 203.640 191.160 ;
        RECT 203.720 190.840 204.040 191.160 ;
        RECT 204.120 190.840 204.440 191.160 ;
        RECT 204.520 190.840 204.840 191.160 ;
        RECT 204.920 190.840 205.240 191.160 ;
        RECT 205.320 190.840 205.640 191.160 ;
        RECT 0.040 190.440 0.360 190.760 ;
        RECT 0.440 190.440 0.760 190.760 ;
        RECT 0.840 190.440 1.160 190.760 ;
        RECT 1.240 190.440 1.560 190.760 ;
        RECT 1.640 190.440 1.960 190.760 ;
        RECT 2.040 190.440 2.360 190.760 ;
        RECT 2.440 190.440 2.760 190.760 ;
        RECT 2.840 190.440 3.160 190.760 ;
        RECT 3.240 190.440 3.560 190.760 ;
        RECT 3.640 190.440 3.960 190.760 ;
        RECT 4.040 190.440 4.360 190.760 ;
        RECT 4.440 190.440 4.760 190.760 ;
        RECT 4.840 190.440 5.160 190.760 ;
        RECT 5.240 190.440 5.560 190.760 ;
        RECT 5.640 190.440 5.960 190.760 ;
        RECT 6.040 190.440 6.360 190.760 ;
        RECT 6.440 190.440 6.760 190.760 ;
        RECT 6.840 190.440 7.160 190.760 ;
        RECT 7.240 190.440 7.560 190.760 ;
        RECT 7.640 190.440 7.960 190.760 ;
        RECT 8.040 190.440 8.360 190.760 ;
        RECT 8.440 190.440 8.760 190.760 ;
        RECT 8.840 190.440 9.160 190.760 ;
        RECT 9.240 190.440 9.560 190.760 ;
        RECT 9.640 190.440 9.960 190.760 ;
        RECT 10.040 190.440 10.360 190.760 ;
        RECT 10.440 190.440 10.760 190.760 ;
        RECT 10.840 190.440 11.160 190.760 ;
        RECT 11.240 190.440 11.560 190.760 ;
        RECT 11.640 190.440 11.960 190.760 ;
        RECT 12.040 190.440 12.360 190.760 ;
        RECT 12.440 190.440 12.760 190.760 ;
        RECT 12.840 190.440 13.160 190.760 ;
        RECT 13.240 190.440 13.560 190.760 ;
        RECT 13.640 190.440 13.960 190.760 ;
        RECT 14.040 190.440 14.360 190.760 ;
        RECT 14.440 190.440 14.760 190.760 ;
        RECT 14.840 190.440 15.160 190.760 ;
        RECT 15.240 190.440 15.560 190.760 ;
        RECT 15.640 190.440 15.960 190.760 ;
        RECT 16.040 190.440 16.360 190.760 ;
        RECT 16.440 190.440 16.760 190.760 ;
        RECT 16.840 190.440 17.160 190.760 ;
        RECT 17.240 190.440 17.560 190.760 ;
        RECT 17.640 190.440 17.960 190.760 ;
        RECT 18.040 190.440 18.360 190.760 ;
        RECT 18.440 190.440 18.760 190.760 ;
        RECT 18.840 190.440 19.160 190.760 ;
        RECT 19.240 190.440 19.560 190.760 ;
        RECT 19.640 190.440 19.960 190.760 ;
        RECT 95.560 190.440 95.880 190.760 ;
        RECT 95.960 190.440 96.280 190.760 ;
        RECT 96.360 190.440 96.680 190.760 ;
        RECT 96.760 190.440 97.080 190.760 ;
        RECT 145.560 190.440 145.880 190.760 ;
        RECT 145.960 190.440 146.280 190.760 ;
        RECT 146.360 190.440 146.680 190.760 ;
        RECT 146.760 190.440 147.080 190.760 ;
        RECT 185.720 190.440 186.040 190.760 ;
        RECT 186.120 190.440 186.440 190.760 ;
        RECT 186.520 190.440 186.840 190.760 ;
        RECT 186.920 190.440 187.240 190.760 ;
        RECT 187.320 190.440 187.640 190.760 ;
        RECT 187.720 190.440 188.040 190.760 ;
        RECT 188.120 190.440 188.440 190.760 ;
        RECT 188.520 190.440 188.840 190.760 ;
        RECT 188.920 190.440 189.240 190.760 ;
        RECT 189.320 190.440 189.640 190.760 ;
        RECT 189.720 190.440 190.040 190.760 ;
        RECT 190.120 190.440 190.440 190.760 ;
        RECT 190.520 190.440 190.840 190.760 ;
        RECT 190.920 190.440 191.240 190.760 ;
        RECT 191.320 190.440 191.640 190.760 ;
        RECT 191.720 190.440 192.040 190.760 ;
        RECT 192.120 190.440 192.440 190.760 ;
        RECT 192.520 190.440 192.840 190.760 ;
        RECT 192.920 190.440 193.240 190.760 ;
        RECT 193.320 190.440 193.640 190.760 ;
        RECT 193.720 190.440 194.040 190.760 ;
        RECT 194.120 190.440 194.440 190.760 ;
        RECT 194.520 190.440 194.840 190.760 ;
        RECT 194.920 190.440 195.240 190.760 ;
        RECT 195.320 190.440 195.640 190.760 ;
        RECT 195.720 190.440 196.040 190.760 ;
        RECT 196.120 190.440 196.440 190.760 ;
        RECT 196.520 190.440 196.840 190.760 ;
        RECT 196.920 190.440 197.240 190.760 ;
        RECT 197.320 190.440 197.640 190.760 ;
        RECT 197.720 190.440 198.040 190.760 ;
        RECT 198.120 190.440 198.440 190.760 ;
        RECT 198.520 190.440 198.840 190.760 ;
        RECT 198.920 190.440 199.240 190.760 ;
        RECT 199.320 190.440 199.640 190.760 ;
        RECT 199.720 190.440 200.040 190.760 ;
        RECT 200.120 190.440 200.440 190.760 ;
        RECT 200.520 190.440 200.840 190.760 ;
        RECT 200.920 190.440 201.240 190.760 ;
        RECT 201.320 190.440 201.640 190.760 ;
        RECT 201.720 190.440 202.040 190.760 ;
        RECT 202.120 190.440 202.440 190.760 ;
        RECT 202.520 190.440 202.840 190.760 ;
        RECT 202.920 190.440 203.240 190.760 ;
        RECT 203.320 190.440 203.640 190.760 ;
        RECT 203.720 190.440 204.040 190.760 ;
        RECT 204.120 190.440 204.440 190.760 ;
        RECT 204.520 190.440 204.840 190.760 ;
        RECT 204.920 190.440 205.240 190.760 ;
        RECT 205.320 190.440 205.640 190.760 ;
        RECT 0.040 190.040 0.360 190.360 ;
        RECT 0.440 190.040 0.760 190.360 ;
        RECT 0.840 190.040 1.160 190.360 ;
        RECT 1.240 190.040 1.560 190.360 ;
        RECT 1.640 190.040 1.960 190.360 ;
        RECT 2.040 190.040 2.360 190.360 ;
        RECT 2.440 190.040 2.760 190.360 ;
        RECT 2.840 190.040 3.160 190.360 ;
        RECT 3.240 190.040 3.560 190.360 ;
        RECT 3.640 190.040 3.960 190.360 ;
        RECT 4.040 190.040 4.360 190.360 ;
        RECT 4.440 190.040 4.760 190.360 ;
        RECT 4.840 190.040 5.160 190.360 ;
        RECT 5.240 190.040 5.560 190.360 ;
        RECT 5.640 190.040 5.960 190.360 ;
        RECT 6.040 190.040 6.360 190.360 ;
        RECT 6.440 190.040 6.760 190.360 ;
        RECT 6.840 190.040 7.160 190.360 ;
        RECT 7.240 190.040 7.560 190.360 ;
        RECT 7.640 190.040 7.960 190.360 ;
        RECT 8.040 190.040 8.360 190.360 ;
        RECT 8.440 190.040 8.760 190.360 ;
        RECT 8.840 190.040 9.160 190.360 ;
        RECT 9.240 190.040 9.560 190.360 ;
        RECT 9.640 190.040 9.960 190.360 ;
        RECT 10.040 190.040 10.360 190.360 ;
        RECT 10.440 190.040 10.760 190.360 ;
        RECT 10.840 190.040 11.160 190.360 ;
        RECT 11.240 190.040 11.560 190.360 ;
        RECT 11.640 190.040 11.960 190.360 ;
        RECT 12.040 190.040 12.360 190.360 ;
        RECT 12.440 190.040 12.760 190.360 ;
        RECT 12.840 190.040 13.160 190.360 ;
        RECT 13.240 190.040 13.560 190.360 ;
        RECT 13.640 190.040 13.960 190.360 ;
        RECT 14.040 190.040 14.360 190.360 ;
        RECT 14.440 190.040 14.760 190.360 ;
        RECT 14.840 190.040 15.160 190.360 ;
        RECT 15.240 190.040 15.560 190.360 ;
        RECT 15.640 190.040 15.960 190.360 ;
        RECT 16.040 190.040 16.360 190.360 ;
        RECT 16.440 190.040 16.760 190.360 ;
        RECT 16.840 190.040 17.160 190.360 ;
        RECT 17.240 190.040 17.560 190.360 ;
        RECT 17.640 190.040 17.960 190.360 ;
        RECT 18.040 190.040 18.360 190.360 ;
        RECT 18.440 190.040 18.760 190.360 ;
        RECT 18.840 190.040 19.160 190.360 ;
        RECT 19.240 190.040 19.560 190.360 ;
        RECT 19.640 190.040 19.960 190.360 ;
        RECT 95.560 190.040 95.880 190.360 ;
        RECT 95.960 190.040 96.280 190.360 ;
        RECT 96.360 190.040 96.680 190.360 ;
        RECT 96.760 190.040 97.080 190.360 ;
        RECT 145.560 190.040 145.880 190.360 ;
        RECT 145.960 190.040 146.280 190.360 ;
        RECT 146.360 190.040 146.680 190.360 ;
        RECT 146.760 190.040 147.080 190.360 ;
        RECT 185.720 190.040 186.040 190.360 ;
        RECT 186.120 190.040 186.440 190.360 ;
        RECT 186.520 190.040 186.840 190.360 ;
        RECT 186.920 190.040 187.240 190.360 ;
        RECT 187.320 190.040 187.640 190.360 ;
        RECT 187.720 190.040 188.040 190.360 ;
        RECT 188.120 190.040 188.440 190.360 ;
        RECT 188.520 190.040 188.840 190.360 ;
        RECT 188.920 190.040 189.240 190.360 ;
        RECT 189.320 190.040 189.640 190.360 ;
        RECT 189.720 190.040 190.040 190.360 ;
        RECT 190.120 190.040 190.440 190.360 ;
        RECT 190.520 190.040 190.840 190.360 ;
        RECT 190.920 190.040 191.240 190.360 ;
        RECT 191.320 190.040 191.640 190.360 ;
        RECT 191.720 190.040 192.040 190.360 ;
        RECT 192.120 190.040 192.440 190.360 ;
        RECT 192.520 190.040 192.840 190.360 ;
        RECT 192.920 190.040 193.240 190.360 ;
        RECT 193.320 190.040 193.640 190.360 ;
        RECT 193.720 190.040 194.040 190.360 ;
        RECT 194.120 190.040 194.440 190.360 ;
        RECT 194.520 190.040 194.840 190.360 ;
        RECT 194.920 190.040 195.240 190.360 ;
        RECT 195.320 190.040 195.640 190.360 ;
        RECT 195.720 190.040 196.040 190.360 ;
        RECT 196.120 190.040 196.440 190.360 ;
        RECT 196.520 190.040 196.840 190.360 ;
        RECT 196.920 190.040 197.240 190.360 ;
        RECT 197.320 190.040 197.640 190.360 ;
        RECT 197.720 190.040 198.040 190.360 ;
        RECT 198.120 190.040 198.440 190.360 ;
        RECT 198.520 190.040 198.840 190.360 ;
        RECT 198.920 190.040 199.240 190.360 ;
        RECT 199.320 190.040 199.640 190.360 ;
        RECT 199.720 190.040 200.040 190.360 ;
        RECT 200.120 190.040 200.440 190.360 ;
        RECT 200.520 190.040 200.840 190.360 ;
        RECT 200.920 190.040 201.240 190.360 ;
        RECT 201.320 190.040 201.640 190.360 ;
        RECT 201.720 190.040 202.040 190.360 ;
        RECT 202.120 190.040 202.440 190.360 ;
        RECT 202.520 190.040 202.840 190.360 ;
        RECT 202.920 190.040 203.240 190.360 ;
        RECT 203.320 190.040 203.640 190.360 ;
        RECT 203.720 190.040 204.040 190.360 ;
        RECT 204.120 190.040 204.440 190.360 ;
        RECT 204.520 190.040 204.840 190.360 ;
        RECT 204.920 190.040 205.240 190.360 ;
        RECT 205.320 190.040 205.640 190.360 ;
        RECT 0.040 189.640 0.360 189.960 ;
        RECT 0.440 189.640 0.760 189.960 ;
        RECT 0.840 189.640 1.160 189.960 ;
        RECT 1.240 189.640 1.560 189.960 ;
        RECT 1.640 189.640 1.960 189.960 ;
        RECT 2.040 189.640 2.360 189.960 ;
        RECT 2.440 189.640 2.760 189.960 ;
        RECT 2.840 189.640 3.160 189.960 ;
        RECT 3.240 189.640 3.560 189.960 ;
        RECT 3.640 189.640 3.960 189.960 ;
        RECT 4.040 189.640 4.360 189.960 ;
        RECT 4.440 189.640 4.760 189.960 ;
        RECT 4.840 189.640 5.160 189.960 ;
        RECT 5.240 189.640 5.560 189.960 ;
        RECT 5.640 189.640 5.960 189.960 ;
        RECT 6.040 189.640 6.360 189.960 ;
        RECT 6.440 189.640 6.760 189.960 ;
        RECT 6.840 189.640 7.160 189.960 ;
        RECT 7.240 189.640 7.560 189.960 ;
        RECT 7.640 189.640 7.960 189.960 ;
        RECT 8.040 189.640 8.360 189.960 ;
        RECT 8.440 189.640 8.760 189.960 ;
        RECT 8.840 189.640 9.160 189.960 ;
        RECT 9.240 189.640 9.560 189.960 ;
        RECT 9.640 189.640 9.960 189.960 ;
        RECT 10.040 189.640 10.360 189.960 ;
        RECT 10.440 189.640 10.760 189.960 ;
        RECT 10.840 189.640 11.160 189.960 ;
        RECT 11.240 189.640 11.560 189.960 ;
        RECT 11.640 189.640 11.960 189.960 ;
        RECT 12.040 189.640 12.360 189.960 ;
        RECT 12.440 189.640 12.760 189.960 ;
        RECT 12.840 189.640 13.160 189.960 ;
        RECT 13.240 189.640 13.560 189.960 ;
        RECT 13.640 189.640 13.960 189.960 ;
        RECT 14.040 189.640 14.360 189.960 ;
        RECT 14.440 189.640 14.760 189.960 ;
        RECT 14.840 189.640 15.160 189.960 ;
        RECT 15.240 189.640 15.560 189.960 ;
        RECT 15.640 189.640 15.960 189.960 ;
        RECT 16.040 189.640 16.360 189.960 ;
        RECT 16.440 189.640 16.760 189.960 ;
        RECT 16.840 189.640 17.160 189.960 ;
        RECT 17.240 189.640 17.560 189.960 ;
        RECT 17.640 189.640 17.960 189.960 ;
        RECT 18.040 189.640 18.360 189.960 ;
        RECT 18.440 189.640 18.760 189.960 ;
        RECT 18.840 189.640 19.160 189.960 ;
        RECT 19.240 189.640 19.560 189.960 ;
        RECT 19.640 189.640 19.960 189.960 ;
        RECT 95.560 189.640 95.880 189.960 ;
        RECT 95.960 189.640 96.280 189.960 ;
        RECT 96.360 189.640 96.680 189.960 ;
        RECT 96.760 189.640 97.080 189.960 ;
        RECT 145.560 189.640 145.880 189.960 ;
        RECT 145.960 189.640 146.280 189.960 ;
        RECT 146.360 189.640 146.680 189.960 ;
        RECT 146.760 189.640 147.080 189.960 ;
        RECT 185.720 189.640 186.040 189.960 ;
        RECT 186.120 189.640 186.440 189.960 ;
        RECT 186.520 189.640 186.840 189.960 ;
        RECT 186.920 189.640 187.240 189.960 ;
        RECT 187.320 189.640 187.640 189.960 ;
        RECT 187.720 189.640 188.040 189.960 ;
        RECT 188.120 189.640 188.440 189.960 ;
        RECT 188.520 189.640 188.840 189.960 ;
        RECT 188.920 189.640 189.240 189.960 ;
        RECT 189.320 189.640 189.640 189.960 ;
        RECT 189.720 189.640 190.040 189.960 ;
        RECT 190.120 189.640 190.440 189.960 ;
        RECT 190.520 189.640 190.840 189.960 ;
        RECT 190.920 189.640 191.240 189.960 ;
        RECT 191.320 189.640 191.640 189.960 ;
        RECT 191.720 189.640 192.040 189.960 ;
        RECT 192.120 189.640 192.440 189.960 ;
        RECT 192.520 189.640 192.840 189.960 ;
        RECT 192.920 189.640 193.240 189.960 ;
        RECT 193.320 189.640 193.640 189.960 ;
        RECT 193.720 189.640 194.040 189.960 ;
        RECT 194.120 189.640 194.440 189.960 ;
        RECT 194.520 189.640 194.840 189.960 ;
        RECT 194.920 189.640 195.240 189.960 ;
        RECT 195.320 189.640 195.640 189.960 ;
        RECT 195.720 189.640 196.040 189.960 ;
        RECT 196.120 189.640 196.440 189.960 ;
        RECT 196.520 189.640 196.840 189.960 ;
        RECT 196.920 189.640 197.240 189.960 ;
        RECT 197.320 189.640 197.640 189.960 ;
        RECT 197.720 189.640 198.040 189.960 ;
        RECT 198.120 189.640 198.440 189.960 ;
        RECT 198.520 189.640 198.840 189.960 ;
        RECT 198.920 189.640 199.240 189.960 ;
        RECT 199.320 189.640 199.640 189.960 ;
        RECT 199.720 189.640 200.040 189.960 ;
        RECT 200.120 189.640 200.440 189.960 ;
        RECT 200.520 189.640 200.840 189.960 ;
        RECT 200.920 189.640 201.240 189.960 ;
        RECT 201.320 189.640 201.640 189.960 ;
        RECT 201.720 189.640 202.040 189.960 ;
        RECT 202.120 189.640 202.440 189.960 ;
        RECT 202.520 189.640 202.840 189.960 ;
        RECT 202.920 189.640 203.240 189.960 ;
        RECT 203.320 189.640 203.640 189.960 ;
        RECT 203.720 189.640 204.040 189.960 ;
        RECT 204.120 189.640 204.440 189.960 ;
        RECT 204.520 189.640 204.840 189.960 ;
        RECT 204.920 189.640 205.240 189.960 ;
        RECT 205.320 189.640 205.640 189.960 ;
        RECT 0.040 189.240 0.360 189.560 ;
        RECT 0.440 189.240 0.760 189.560 ;
        RECT 0.840 189.240 1.160 189.560 ;
        RECT 1.240 189.240 1.560 189.560 ;
        RECT 1.640 189.240 1.960 189.560 ;
        RECT 2.040 189.240 2.360 189.560 ;
        RECT 2.440 189.240 2.760 189.560 ;
        RECT 2.840 189.240 3.160 189.560 ;
        RECT 3.240 189.240 3.560 189.560 ;
        RECT 3.640 189.240 3.960 189.560 ;
        RECT 4.040 189.240 4.360 189.560 ;
        RECT 4.440 189.240 4.760 189.560 ;
        RECT 4.840 189.240 5.160 189.560 ;
        RECT 5.240 189.240 5.560 189.560 ;
        RECT 5.640 189.240 5.960 189.560 ;
        RECT 6.040 189.240 6.360 189.560 ;
        RECT 6.440 189.240 6.760 189.560 ;
        RECT 6.840 189.240 7.160 189.560 ;
        RECT 7.240 189.240 7.560 189.560 ;
        RECT 7.640 189.240 7.960 189.560 ;
        RECT 8.040 189.240 8.360 189.560 ;
        RECT 8.440 189.240 8.760 189.560 ;
        RECT 8.840 189.240 9.160 189.560 ;
        RECT 9.240 189.240 9.560 189.560 ;
        RECT 9.640 189.240 9.960 189.560 ;
        RECT 10.040 189.240 10.360 189.560 ;
        RECT 10.440 189.240 10.760 189.560 ;
        RECT 10.840 189.240 11.160 189.560 ;
        RECT 11.240 189.240 11.560 189.560 ;
        RECT 11.640 189.240 11.960 189.560 ;
        RECT 12.040 189.240 12.360 189.560 ;
        RECT 12.440 189.240 12.760 189.560 ;
        RECT 12.840 189.240 13.160 189.560 ;
        RECT 13.240 189.240 13.560 189.560 ;
        RECT 13.640 189.240 13.960 189.560 ;
        RECT 14.040 189.240 14.360 189.560 ;
        RECT 14.440 189.240 14.760 189.560 ;
        RECT 14.840 189.240 15.160 189.560 ;
        RECT 15.240 189.240 15.560 189.560 ;
        RECT 15.640 189.240 15.960 189.560 ;
        RECT 16.040 189.240 16.360 189.560 ;
        RECT 16.440 189.240 16.760 189.560 ;
        RECT 16.840 189.240 17.160 189.560 ;
        RECT 17.240 189.240 17.560 189.560 ;
        RECT 17.640 189.240 17.960 189.560 ;
        RECT 18.040 189.240 18.360 189.560 ;
        RECT 18.440 189.240 18.760 189.560 ;
        RECT 18.840 189.240 19.160 189.560 ;
        RECT 19.240 189.240 19.560 189.560 ;
        RECT 19.640 189.240 19.960 189.560 ;
        RECT 95.560 189.240 95.880 189.560 ;
        RECT 95.960 189.240 96.280 189.560 ;
        RECT 96.360 189.240 96.680 189.560 ;
        RECT 96.760 189.240 97.080 189.560 ;
        RECT 145.560 189.240 145.880 189.560 ;
        RECT 145.960 189.240 146.280 189.560 ;
        RECT 146.360 189.240 146.680 189.560 ;
        RECT 146.760 189.240 147.080 189.560 ;
        RECT 185.720 189.240 186.040 189.560 ;
        RECT 186.120 189.240 186.440 189.560 ;
        RECT 186.520 189.240 186.840 189.560 ;
        RECT 186.920 189.240 187.240 189.560 ;
        RECT 187.320 189.240 187.640 189.560 ;
        RECT 187.720 189.240 188.040 189.560 ;
        RECT 188.120 189.240 188.440 189.560 ;
        RECT 188.520 189.240 188.840 189.560 ;
        RECT 188.920 189.240 189.240 189.560 ;
        RECT 189.320 189.240 189.640 189.560 ;
        RECT 189.720 189.240 190.040 189.560 ;
        RECT 190.120 189.240 190.440 189.560 ;
        RECT 190.520 189.240 190.840 189.560 ;
        RECT 190.920 189.240 191.240 189.560 ;
        RECT 191.320 189.240 191.640 189.560 ;
        RECT 191.720 189.240 192.040 189.560 ;
        RECT 192.120 189.240 192.440 189.560 ;
        RECT 192.520 189.240 192.840 189.560 ;
        RECT 192.920 189.240 193.240 189.560 ;
        RECT 193.320 189.240 193.640 189.560 ;
        RECT 193.720 189.240 194.040 189.560 ;
        RECT 194.120 189.240 194.440 189.560 ;
        RECT 194.520 189.240 194.840 189.560 ;
        RECT 194.920 189.240 195.240 189.560 ;
        RECT 195.320 189.240 195.640 189.560 ;
        RECT 195.720 189.240 196.040 189.560 ;
        RECT 196.120 189.240 196.440 189.560 ;
        RECT 196.520 189.240 196.840 189.560 ;
        RECT 196.920 189.240 197.240 189.560 ;
        RECT 197.320 189.240 197.640 189.560 ;
        RECT 197.720 189.240 198.040 189.560 ;
        RECT 198.120 189.240 198.440 189.560 ;
        RECT 198.520 189.240 198.840 189.560 ;
        RECT 198.920 189.240 199.240 189.560 ;
        RECT 199.320 189.240 199.640 189.560 ;
        RECT 199.720 189.240 200.040 189.560 ;
        RECT 200.120 189.240 200.440 189.560 ;
        RECT 200.520 189.240 200.840 189.560 ;
        RECT 200.920 189.240 201.240 189.560 ;
        RECT 201.320 189.240 201.640 189.560 ;
        RECT 201.720 189.240 202.040 189.560 ;
        RECT 202.120 189.240 202.440 189.560 ;
        RECT 202.520 189.240 202.840 189.560 ;
        RECT 202.920 189.240 203.240 189.560 ;
        RECT 203.320 189.240 203.640 189.560 ;
        RECT 203.720 189.240 204.040 189.560 ;
        RECT 204.120 189.240 204.440 189.560 ;
        RECT 204.520 189.240 204.840 189.560 ;
        RECT 204.920 189.240 205.240 189.560 ;
        RECT 205.320 189.240 205.640 189.560 ;
        RECT 0.040 188.840 0.360 189.160 ;
        RECT 0.440 188.840 0.760 189.160 ;
        RECT 0.840 188.840 1.160 189.160 ;
        RECT 1.240 188.840 1.560 189.160 ;
        RECT 1.640 188.840 1.960 189.160 ;
        RECT 2.040 188.840 2.360 189.160 ;
        RECT 2.440 188.840 2.760 189.160 ;
        RECT 2.840 188.840 3.160 189.160 ;
        RECT 3.240 188.840 3.560 189.160 ;
        RECT 3.640 188.840 3.960 189.160 ;
        RECT 4.040 188.840 4.360 189.160 ;
        RECT 4.440 188.840 4.760 189.160 ;
        RECT 4.840 188.840 5.160 189.160 ;
        RECT 5.240 188.840 5.560 189.160 ;
        RECT 5.640 188.840 5.960 189.160 ;
        RECT 6.040 188.840 6.360 189.160 ;
        RECT 6.440 188.840 6.760 189.160 ;
        RECT 6.840 188.840 7.160 189.160 ;
        RECT 7.240 188.840 7.560 189.160 ;
        RECT 7.640 188.840 7.960 189.160 ;
        RECT 8.040 188.840 8.360 189.160 ;
        RECT 8.440 188.840 8.760 189.160 ;
        RECT 8.840 188.840 9.160 189.160 ;
        RECT 9.240 188.840 9.560 189.160 ;
        RECT 9.640 188.840 9.960 189.160 ;
        RECT 10.040 188.840 10.360 189.160 ;
        RECT 10.440 188.840 10.760 189.160 ;
        RECT 10.840 188.840 11.160 189.160 ;
        RECT 11.240 188.840 11.560 189.160 ;
        RECT 11.640 188.840 11.960 189.160 ;
        RECT 12.040 188.840 12.360 189.160 ;
        RECT 12.440 188.840 12.760 189.160 ;
        RECT 12.840 188.840 13.160 189.160 ;
        RECT 13.240 188.840 13.560 189.160 ;
        RECT 13.640 188.840 13.960 189.160 ;
        RECT 14.040 188.840 14.360 189.160 ;
        RECT 14.440 188.840 14.760 189.160 ;
        RECT 14.840 188.840 15.160 189.160 ;
        RECT 15.240 188.840 15.560 189.160 ;
        RECT 15.640 188.840 15.960 189.160 ;
        RECT 16.040 188.840 16.360 189.160 ;
        RECT 16.440 188.840 16.760 189.160 ;
        RECT 16.840 188.840 17.160 189.160 ;
        RECT 17.240 188.840 17.560 189.160 ;
        RECT 17.640 188.840 17.960 189.160 ;
        RECT 18.040 188.840 18.360 189.160 ;
        RECT 18.440 188.840 18.760 189.160 ;
        RECT 18.840 188.840 19.160 189.160 ;
        RECT 19.240 188.840 19.560 189.160 ;
        RECT 19.640 188.840 19.960 189.160 ;
        RECT 95.560 188.840 95.880 189.160 ;
        RECT 95.960 188.840 96.280 189.160 ;
        RECT 96.360 188.840 96.680 189.160 ;
        RECT 96.760 188.840 97.080 189.160 ;
        RECT 145.560 188.840 145.880 189.160 ;
        RECT 145.960 188.840 146.280 189.160 ;
        RECT 146.360 188.840 146.680 189.160 ;
        RECT 146.760 188.840 147.080 189.160 ;
        RECT 185.720 188.840 186.040 189.160 ;
        RECT 186.120 188.840 186.440 189.160 ;
        RECT 186.520 188.840 186.840 189.160 ;
        RECT 186.920 188.840 187.240 189.160 ;
        RECT 187.320 188.840 187.640 189.160 ;
        RECT 187.720 188.840 188.040 189.160 ;
        RECT 188.120 188.840 188.440 189.160 ;
        RECT 188.520 188.840 188.840 189.160 ;
        RECT 188.920 188.840 189.240 189.160 ;
        RECT 189.320 188.840 189.640 189.160 ;
        RECT 189.720 188.840 190.040 189.160 ;
        RECT 190.120 188.840 190.440 189.160 ;
        RECT 190.520 188.840 190.840 189.160 ;
        RECT 190.920 188.840 191.240 189.160 ;
        RECT 191.320 188.840 191.640 189.160 ;
        RECT 191.720 188.840 192.040 189.160 ;
        RECT 192.120 188.840 192.440 189.160 ;
        RECT 192.520 188.840 192.840 189.160 ;
        RECT 192.920 188.840 193.240 189.160 ;
        RECT 193.320 188.840 193.640 189.160 ;
        RECT 193.720 188.840 194.040 189.160 ;
        RECT 194.120 188.840 194.440 189.160 ;
        RECT 194.520 188.840 194.840 189.160 ;
        RECT 194.920 188.840 195.240 189.160 ;
        RECT 195.320 188.840 195.640 189.160 ;
        RECT 195.720 188.840 196.040 189.160 ;
        RECT 196.120 188.840 196.440 189.160 ;
        RECT 196.520 188.840 196.840 189.160 ;
        RECT 196.920 188.840 197.240 189.160 ;
        RECT 197.320 188.840 197.640 189.160 ;
        RECT 197.720 188.840 198.040 189.160 ;
        RECT 198.120 188.840 198.440 189.160 ;
        RECT 198.520 188.840 198.840 189.160 ;
        RECT 198.920 188.840 199.240 189.160 ;
        RECT 199.320 188.840 199.640 189.160 ;
        RECT 199.720 188.840 200.040 189.160 ;
        RECT 200.120 188.840 200.440 189.160 ;
        RECT 200.520 188.840 200.840 189.160 ;
        RECT 200.920 188.840 201.240 189.160 ;
        RECT 201.320 188.840 201.640 189.160 ;
        RECT 201.720 188.840 202.040 189.160 ;
        RECT 202.120 188.840 202.440 189.160 ;
        RECT 202.520 188.840 202.840 189.160 ;
        RECT 202.920 188.840 203.240 189.160 ;
        RECT 203.320 188.840 203.640 189.160 ;
        RECT 203.720 188.840 204.040 189.160 ;
        RECT 204.120 188.840 204.440 189.160 ;
        RECT 204.520 188.840 204.840 189.160 ;
        RECT 204.920 188.840 205.240 189.160 ;
        RECT 205.320 188.840 205.640 189.160 ;
        RECT 0.040 188.440 0.360 188.760 ;
        RECT 0.440 188.440 0.760 188.760 ;
        RECT 0.840 188.440 1.160 188.760 ;
        RECT 1.240 188.440 1.560 188.760 ;
        RECT 1.640 188.440 1.960 188.760 ;
        RECT 2.040 188.440 2.360 188.760 ;
        RECT 2.440 188.440 2.760 188.760 ;
        RECT 2.840 188.440 3.160 188.760 ;
        RECT 3.240 188.440 3.560 188.760 ;
        RECT 3.640 188.440 3.960 188.760 ;
        RECT 4.040 188.440 4.360 188.760 ;
        RECT 4.440 188.440 4.760 188.760 ;
        RECT 4.840 188.440 5.160 188.760 ;
        RECT 5.240 188.440 5.560 188.760 ;
        RECT 5.640 188.440 5.960 188.760 ;
        RECT 6.040 188.440 6.360 188.760 ;
        RECT 6.440 188.440 6.760 188.760 ;
        RECT 6.840 188.440 7.160 188.760 ;
        RECT 7.240 188.440 7.560 188.760 ;
        RECT 7.640 188.440 7.960 188.760 ;
        RECT 8.040 188.440 8.360 188.760 ;
        RECT 8.440 188.440 8.760 188.760 ;
        RECT 8.840 188.440 9.160 188.760 ;
        RECT 9.240 188.440 9.560 188.760 ;
        RECT 9.640 188.440 9.960 188.760 ;
        RECT 10.040 188.440 10.360 188.760 ;
        RECT 10.440 188.440 10.760 188.760 ;
        RECT 10.840 188.440 11.160 188.760 ;
        RECT 11.240 188.440 11.560 188.760 ;
        RECT 11.640 188.440 11.960 188.760 ;
        RECT 12.040 188.440 12.360 188.760 ;
        RECT 12.440 188.440 12.760 188.760 ;
        RECT 12.840 188.440 13.160 188.760 ;
        RECT 13.240 188.440 13.560 188.760 ;
        RECT 13.640 188.440 13.960 188.760 ;
        RECT 14.040 188.440 14.360 188.760 ;
        RECT 14.440 188.440 14.760 188.760 ;
        RECT 14.840 188.440 15.160 188.760 ;
        RECT 15.240 188.440 15.560 188.760 ;
        RECT 15.640 188.440 15.960 188.760 ;
        RECT 16.040 188.440 16.360 188.760 ;
        RECT 16.440 188.440 16.760 188.760 ;
        RECT 16.840 188.440 17.160 188.760 ;
        RECT 17.240 188.440 17.560 188.760 ;
        RECT 17.640 188.440 17.960 188.760 ;
        RECT 18.040 188.440 18.360 188.760 ;
        RECT 18.440 188.440 18.760 188.760 ;
        RECT 18.840 188.440 19.160 188.760 ;
        RECT 19.240 188.440 19.560 188.760 ;
        RECT 19.640 188.440 19.960 188.760 ;
        RECT 95.560 188.440 95.880 188.760 ;
        RECT 95.960 188.440 96.280 188.760 ;
        RECT 96.360 188.440 96.680 188.760 ;
        RECT 96.760 188.440 97.080 188.760 ;
        RECT 145.560 188.440 145.880 188.760 ;
        RECT 145.960 188.440 146.280 188.760 ;
        RECT 146.360 188.440 146.680 188.760 ;
        RECT 146.760 188.440 147.080 188.760 ;
        RECT 185.720 188.440 186.040 188.760 ;
        RECT 186.120 188.440 186.440 188.760 ;
        RECT 186.520 188.440 186.840 188.760 ;
        RECT 186.920 188.440 187.240 188.760 ;
        RECT 187.320 188.440 187.640 188.760 ;
        RECT 187.720 188.440 188.040 188.760 ;
        RECT 188.120 188.440 188.440 188.760 ;
        RECT 188.520 188.440 188.840 188.760 ;
        RECT 188.920 188.440 189.240 188.760 ;
        RECT 189.320 188.440 189.640 188.760 ;
        RECT 189.720 188.440 190.040 188.760 ;
        RECT 190.120 188.440 190.440 188.760 ;
        RECT 190.520 188.440 190.840 188.760 ;
        RECT 190.920 188.440 191.240 188.760 ;
        RECT 191.320 188.440 191.640 188.760 ;
        RECT 191.720 188.440 192.040 188.760 ;
        RECT 192.120 188.440 192.440 188.760 ;
        RECT 192.520 188.440 192.840 188.760 ;
        RECT 192.920 188.440 193.240 188.760 ;
        RECT 193.320 188.440 193.640 188.760 ;
        RECT 193.720 188.440 194.040 188.760 ;
        RECT 194.120 188.440 194.440 188.760 ;
        RECT 194.520 188.440 194.840 188.760 ;
        RECT 194.920 188.440 195.240 188.760 ;
        RECT 195.320 188.440 195.640 188.760 ;
        RECT 195.720 188.440 196.040 188.760 ;
        RECT 196.120 188.440 196.440 188.760 ;
        RECT 196.520 188.440 196.840 188.760 ;
        RECT 196.920 188.440 197.240 188.760 ;
        RECT 197.320 188.440 197.640 188.760 ;
        RECT 197.720 188.440 198.040 188.760 ;
        RECT 198.120 188.440 198.440 188.760 ;
        RECT 198.520 188.440 198.840 188.760 ;
        RECT 198.920 188.440 199.240 188.760 ;
        RECT 199.320 188.440 199.640 188.760 ;
        RECT 199.720 188.440 200.040 188.760 ;
        RECT 200.120 188.440 200.440 188.760 ;
        RECT 200.520 188.440 200.840 188.760 ;
        RECT 200.920 188.440 201.240 188.760 ;
        RECT 201.320 188.440 201.640 188.760 ;
        RECT 201.720 188.440 202.040 188.760 ;
        RECT 202.120 188.440 202.440 188.760 ;
        RECT 202.520 188.440 202.840 188.760 ;
        RECT 202.920 188.440 203.240 188.760 ;
        RECT 203.320 188.440 203.640 188.760 ;
        RECT 203.720 188.440 204.040 188.760 ;
        RECT 204.120 188.440 204.440 188.760 ;
        RECT 204.520 188.440 204.840 188.760 ;
        RECT 204.920 188.440 205.240 188.760 ;
        RECT 205.320 188.440 205.640 188.760 ;
        RECT 0.040 188.040 0.360 188.360 ;
        RECT 0.440 188.040 0.760 188.360 ;
        RECT 0.840 188.040 1.160 188.360 ;
        RECT 1.240 188.040 1.560 188.360 ;
        RECT 1.640 188.040 1.960 188.360 ;
        RECT 2.040 188.040 2.360 188.360 ;
        RECT 2.440 188.040 2.760 188.360 ;
        RECT 2.840 188.040 3.160 188.360 ;
        RECT 3.240 188.040 3.560 188.360 ;
        RECT 3.640 188.040 3.960 188.360 ;
        RECT 4.040 188.040 4.360 188.360 ;
        RECT 4.440 188.040 4.760 188.360 ;
        RECT 4.840 188.040 5.160 188.360 ;
        RECT 5.240 188.040 5.560 188.360 ;
        RECT 5.640 188.040 5.960 188.360 ;
        RECT 6.040 188.040 6.360 188.360 ;
        RECT 6.440 188.040 6.760 188.360 ;
        RECT 6.840 188.040 7.160 188.360 ;
        RECT 7.240 188.040 7.560 188.360 ;
        RECT 7.640 188.040 7.960 188.360 ;
        RECT 8.040 188.040 8.360 188.360 ;
        RECT 8.440 188.040 8.760 188.360 ;
        RECT 8.840 188.040 9.160 188.360 ;
        RECT 9.240 188.040 9.560 188.360 ;
        RECT 9.640 188.040 9.960 188.360 ;
        RECT 10.040 188.040 10.360 188.360 ;
        RECT 10.440 188.040 10.760 188.360 ;
        RECT 10.840 188.040 11.160 188.360 ;
        RECT 11.240 188.040 11.560 188.360 ;
        RECT 11.640 188.040 11.960 188.360 ;
        RECT 12.040 188.040 12.360 188.360 ;
        RECT 12.440 188.040 12.760 188.360 ;
        RECT 12.840 188.040 13.160 188.360 ;
        RECT 13.240 188.040 13.560 188.360 ;
        RECT 13.640 188.040 13.960 188.360 ;
        RECT 14.040 188.040 14.360 188.360 ;
        RECT 14.440 188.040 14.760 188.360 ;
        RECT 14.840 188.040 15.160 188.360 ;
        RECT 15.240 188.040 15.560 188.360 ;
        RECT 15.640 188.040 15.960 188.360 ;
        RECT 16.040 188.040 16.360 188.360 ;
        RECT 16.440 188.040 16.760 188.360 ;
        RECT 16.840 188.040 17.160 188.360 ;
        RECT 17.240 188.040 17.560 188.360 ;
        RECT 17.640 188.040 17.960 188.360 ;
        RECT 18.040 188.040 18.360 188.360 ;
        RECT 18.440 188.040 18.760 188.360 ;
        RECT 18.840 188.040 19.160 188.360 ;
        RECT 19.240 188.040 19.560 188.360 ;
        RECT 19.640 188.040 19.960 188.360 ;
        RECT 95.560 188.040 95.880 188.360 ;
        RECT 95.960 188.040 96.280 188.360 ;
        RECT 96.360 188.040 96.680 188.360 ;
        RECT 96.760 188.040 97.080 188.360 ;
        RECT 145.560 188.040 145.880 188.360 ;
        RECT 145.960 188.040 146.280 188.360 ;
        RECT 146.360 188.040 146.680 188.360 ;
        RECT 146.760 188.040 147.080 188.360 ;
        RECT 185.720 188.040 186.040 188.360 ;
        RECT 186.120 188.040 186.440 188.360 ;
        RECT 186.520 188.040 186.840 188.360 ;
        RECT 186.920 188.040 187.240 188.360 ;
        RECT 187.320 188.040 187.640 188.360 ;
        RECT 187.720 188.040 188.040 188.360 ;
        RECT 188.120 188.040 188.440 188.360 ;
        RECT 188.520 188.040 188.840 188.360 ;
        RECT 188.920 188.040 189.240 188.360 ;
        RECT 189.320 188.040 189.640 188.360 ;
        RECT 189.720 188.040 190.040 188.360 ;
        RECT 190.120 188.040 190.440 188.360 ;
        RECT 190.520 188.040 190.840 188.360 ;
        RECT 190.920 188.040 191.240 188.360 ;
        RECT 191.320 188.040 191.640 188.360 ;
        RECT 191.720 188.040 192.040 188.360 ;
        RECT 192.120 188.040 192.440 188.360 ;
        RECT 192.520 188.040 192.840 188.360 ;
        RECT 192.920 188.040 193.240 188.360 ;
        RECT 193.320 188.040 193.640 188.360 ;
        RECT 193.720 188.040 194.040 188.360 ;
        RECT 194.120 188.040 194.440 188.360 ;
        RECT 194.520 188.040 194.840 188.360 ;
        RECT 194.920 188.040 195.240 188.360 ;
        RECT 195.320 188.040 195.640 188.360 ;
        RECT 195.720 188.040 196.040 188.360 ;
        RECT 196.120 188.040 196.440 188.360 ;
        RECT 196.520 188.040 196.840 188.360 ;
        RECT 196.920 188.040 197.240 188.360 ;
        RECT 197.320 188.040 197.640 188.360 ;
        RECT 197.720 188.040 198.040 188.360 ;
        RECT 198.120 188.040 198.440 188.360 ;
        RECT 198.520 188.040 198.840 188.360 ;
        RECT 198.920 188.040 199.240 188.360 ;
        RECT 199.320 188.040 199.640 188.360 ;
        RECT 199.720 188.040 200.040 188.360 ;
        RECT 200.120 188.040 200.440 188.360 ;
        RECT 200.520 188.040 200.840 188.360 ;
        RECT 200.920 188.040 201.240 188.360 ;
        RECT 201.320 188.040 201.640 188.360 ;
        RECT 201.720 188.040 202.040 188.360 ;
        RECT 202.120 188.040 202.440 188.360 ;
        RECT 202.520 188.040 202.840 188.360 ;
        RECT 202.920 188.040 203.240 188.360 ;
        RECT 203.320 188.040 203.640 188.360 ;
        RECT 203.720 188.040 204.040 188.360 ;
        RECT 204.120 188.040 204.440 188.360 ;
        RECT 204.520 188.040 204.840 188.360 ;
        RECT 204.920 188.040 205.240 188.360 ;
        RECT 205.320 188.040 205.640 188.360 ;
        RECT 0.040 187.640 0.360 187.960 ;
        RECT 0.440 187.640 0.760 187.960 ;
        RECT 0.840 187.640 1.160 187.960 ;
        RECT 1.240 187.640 1.560 187.960 ;
        RECT 1.640 187.640 1.960 187.960 ;
        RECT 2.040 187.640 2.360 187.960 ;
        RECT 2.440 187.640 2.760 187.960 ;
        RECT 2.840 187.640 3.160 187.960 ;
        RECT 3.240 187.640 3.560 187.960 ;
        RECT 3.640 187.640 3.960 187.960 ;
        RECT 4.040 187.640 4.360 187.960 ;
        RECT 4.440 187.640 4.760 187.960 ;
        RECT 4.840 187.640 5.160 187.960 ;
        RECT 5.240 187.640 5.560 187.960 ;
        RECT 5.640 187.640 5.960 187.960 ;
        RECT 6.040 187.640 6.360 187.960 ;
        RECT 6.440 187.640 6.760 187.960 ;
        RECT 6.840 187.640 7.160 187.960 ;
        RECT 7.240 187.640 7.560 187.960 ;
        RECT 7.640 187.640 7.960 187.960 ;
        RECT 8.040 187.640 8.360 187.960 ;
        RECT 8.440 187.640 8.760 187.960 ;
        RECT 8.840 187.640 9.160 187.960 ;
        RECT 9.240 187.640 9.560 187.960 ;
        RECT 9.640 187.640 9.960 187.960 ;
        RECT 10.040 187.640 10.360 187.960 ;
        RECT 10.440 187.640 10.760 187.960 ;
        RECT 10.840 187.640 11.160 187.960 ;
        RECT 11.240 187.640 11.560 187.960 ;
        RECT 11.640 187.640 11.960 187.960 ;
        RECT 12.040 187.640 12.360 187.960 ;
        RECT 12.440 187.640 12.760 187.960 ;
        RECT 12.840 187.640 13.160 187.960 ;
        RECT 13.240 187.640 13.560 187.960 ;
        RECT 13.640 187.640 13.960 187.960 ;
        RECT 14.040 187.640 14.360 187.960 ;
        RECT 14.440 187.640 14.760 187.960 ;
        RECT 14.840 187.640 15.160 187.960 ;
        RECT 15.240 187.640 15.560 187.960 ;
        RECT 15.640 187.640 15.960 187.960 ;
        RECT 16.040 187.640 16.360 187.960 ;
        RECT 16.440 187.640 16.760 187.960 ;
        RECT 16.840 187.640 17.160 187.960 ;
        RECT 17.240 187.640 17.560 187.960 ;
        RECT 17.640 187.640 17.960 187.960 ;
        RECT 18.040 187.640 18.360 187.960 ;
        RECT 18.440 187.640 18.760 187.960 ;
        RECT 18.840 187.640 19.160 187.960 ;
        RECT 19.240 187.640 19.560 187.960 ;
        RECT 19.640 187.640 19.960 187.960 ;
        RECT 95.560 187.640 95.880 187.960 ;
        RECT 95.960 187.640 96.280 187.960 ;
        RECT 96.360 187.640 96.680 187.960 ;
        RECT 96.760 187.640 97.080 187.960 ;
        RECT 145.560 187.640 145.880 187.960 ;
        RECT 145.960 187.640 146.280 187.960 ;
        RECT 146.360 187.640 146.680 187.960 ;
        RECT 146.760 187.640 147.080 187.960 ;
        RECT 185.720 187.640 186.040 187.960 ;
        RECT 186.120 187.640 186.440 187.960 ;
        RECT 186.520 187.640 186.840 187.960 ;
        RECT 186.920 187.640 187.240 187.960 ;
        RECT 187.320 187.640 187.640 187.960 ;
        RECT 187.720 187.640 188.040 187.960 ;
        RECT 188.120 187.640 188.440 187.960 ;
        RECT 188.520 187.640 188.840 187.960 ;
        RECT 188.920 187.640 189.240 187.960 ;
        RECT 189.320 187.640 189.640 187.960 ;
        RECT 189.720 187.640 190.040 187.960 ;
        RECT 190.120 187.640 190.440 187.960 ;
        RECT 190.520 187.640 190.840 187.960 ;
        RECT 190.920 187.640 191.240 187.960 ;
        RECT 191.320 187.640 191.640 187.960 ;
        RECT 191.720 187.640 192.040 187.960 ;
        RECT 192.120 187.640 192.440 187.960 ;
        RECT 192.520 187.640 192.840 187.960 ;
        RECT 192.920 187.640 193.240 187.960 ;
        RECT 193.320 187.640 193.640 187.960 ;
        RECT 193.720 187.640 194.040 187.960 ;
        RECT 194.120 187.640 194.440 187.960 ;
        RECT 194.520 187.640 194.840 187.960 ;
        RECT 194.920 187.640 195.240 187.960 ;
        RECT 195.320 187.640 195.640 187.960 ;
        RECT 195.720 187.640 196.040 187.960 ;
        RECT 196.120 187.640 196.440 187.960 ;
        RECT 196.520 187.640 196.840 187.960 ;
        RECT 196.920 187.640 197.240 187.960 ;
        RECT 197.320 187.640 197.640 187.960 ;
        RECT 197.720 187.640 198.040 187.960 ;
        RECT 198.120 187.640 198.440 187.960 ;
        RECT 198.520 187.640 198.840 187.960 ;
        RECT 198.920 187.640 199.240 187.960 ;
        RECT 199.320 187.640 199.640 187.960 ;
        RECT 199.720 187.640 200.040 187.960 ;
        RECT 200.120 187.640 200.440 187.960 ;
        RECT 200.520 187.640 200.840 187.960 ;
        RECT 200.920 187.640 201.240 187.960 ;
        RECT 201.320 187.640 201.640 187.960 ;
        RECT 201.720 187.640 202.040 187.960 ;
        RECT 202.120 187.640 202.440 187.960 ;
        RECT 202.520 187.640 202.840 187.960 ;
        RECT 202.920 187.640 203.240 187.960 ;
        RECT 203.320 187.640 203.640 187.960 ;
        RECT 203.720 187.640 204.040 187.960 ;
        RECT 204.120 187.640 204.440 187.960 ;
        RECT 204.520 187.640 204.840 187.960 ;
        RECT 204.920 187.640 205.240 187.960 ;
        RECT 205.320 187.640 205.640 187.960 ;
        RECT 0.040 187.240 0.360 187.560 ;
        RECT 0.440 187.240 0.760 187.560 ;
        RECT 0.840 187.240 1.160 187.560 ;
        RECT 1.240 187.240 1.560 187.560 ;
        RECT 1.640 187.240 1.960 187.560 ;
        RECT 2.040 187.240 2.360 187.560 ;
        RECT 2.440 187.240 2.760 187.560 ;
        RECT 2.840 187.240 3.160 187.560 ;
        RECT 3.240 187.240 3.560 187.560 ;
        RECT 3.640 187.240 3.960 187.560 ;
        RECT 4.040 187.240 4.360 187.560 ;
        RECT 4.440 187.240 4.760 187.560 ;
        RECT 4.840 187.240 5.160 187.560 ;
        RECT 5.240 187.240 5.560 187.560 ;
        RECT 5.640 187.240 5.960 187.560 ;
        RECT 6.040 187.240 6.360 187.560 ;
        RECT 6.440 187.240 6.760 187.560 ;
        RECT 6.840 187.240 7.160 187.560 ;
        RECT 7.240 187.240 7.560 187.560 ;
        RECT 7.640 187.240 7.960 187.560 ;
        RECT 8.040 187.240 8.360 187.560 ;
        RECT 8.440 187.240 8.760 187.560 ;
        RECT 8.840 187.240 9.160 187.560 ;
        RECT 9.240 187.240 9.560 187.560 ;
        RECT 9.640 187.240 9.960 187.560 ;
        RECT 10.040 187.240 10.360 187.560 ;
        RECT 10.440 187.240 10.760 187.560 ;
        RECT 10.840 187.240 11.160 187.560 ;
        RECT 11.240 187.240 11.560 187.560 ;
        RECT 11.640 187.240 11.960 187.560 ;
        RECT 12.040 187.240 12.360 187.560 ;
        RECT 12.440 187.240 12.760 187.560 ;
        RECT 12.840 187.240 13.160 187.560 ;
        RECT 13.240 187.240 13.560 187.560 ;
        RECT 13.640 187.240 13.960 187.560 ;
        RECT 14.040 187.240 14.360 187.560 ;
        RECT 14.440 187.240 14.760 187.560 ;
        RECT 14.840 187.240 15.160 187.560 ;
        RECT 15.240 187.240 15.560 187.560 ;
        RECT 15.640 187.240 15.960 187.560 ;
        RECT 16.040 187.240 16.360 187.560 ;
        RECT 16.440 187.240 16.760 187.560 ;
        RECT 16.840 187.240 17.160 187.560 ;
        RECT 17.240 187.240 17.560 187.560 ;
        RECT 17.640 187.240 17.960 187.560 ;
        RECT 18.040 187.240 18.360 187.560 ;
        RECT 18.440 187.240 18.760 187.560 ;
        RECT 18.840 187.240 19.160 187.560 ;
        RECT 19.240 187.240 19.560 187.560 ;
        RECT 19.640 187.240 19.960 187.560 ;
        RECT 95.560 187.240 95.880 187.560 ;
        RECT 95.960 187.240 96.280 187.560 ;
        RECT 96.360 187.240 96.680 187.560 ;
        RECT 96.760 187.240 97.080 187.560 ;
        RECT 145.560 187.240 145.880 187.560 ;
        RECT 145.960 187.240 146.280 187.560 ;
        RECT 146.360 187.240 146.680 187.560 ;
        RECT 146.760 187.240 147.080 187.560 ;
        RECT 185.720 187.240 186.040 187.560 ;
        RECT 186.120 187.240 186.440 187.560 ;
        RECT 186.520 187.240 186.840 187.560 ;
        RECT 186.920 187.240 187.240 187.560 ;
        RECT 187.320 187.240 187.640 187.560 ;
        RECT 187.720 187.240 188.040 187.560 ;
        RECT 188.120 187.240 188.440 187.560 ;
        RECT 188.520 187.240 188.840 187.560 ;
        RECT 188.920 187.240 189.240 187.560 ;
        RECT 189.320 187.240 189.640 187.560 ;
        RECT 189.720 187.240 190.040 187.560 ;
        RECT 190.120 187.240 190.440 187.560 ;
        RECT 190.520 187.240 190.840 187.560 ;
        RECT 190.920 187.240 191.240 187.560 ;
        RECT 191.320 187.240 191.640 187.560 ;
        RECT 191.720 187.240 192.040 187.560 ;
        RECT 192.120 187.240 192.440 187.560 ;
        RECT 192.520 187.240 192.840 187.560 ;
        RECT 192.920 187.240 193.240 187.560 ;
        RECT 193.320 187.240 193.640 187.560 ;
        RECT 193.720 187.240 194.040 187.560 ;
        RECT 194.120 187.240 194.440 187.560 ;
        RECT 194.520 187.240 194.840 187.560 ;
        RECT 194.920 187.240 195.240 187.560 ;
        RECT 195.320 187.240 195.640 187.560 ;
        RECT 195.720 187.240 196.040 187.560 ;
        RECT 196.120 187.240 196.440 187.560 ;
        RECT 196.520 187.240 196.840 187.560 ;
        RECT 196.920 187.240 197.240 187.560 ;
        RECT 197.320 187.240 197.640 187.560 ;
        RECT 197.720 187.240 198.040 187.560 ;
        RECT 198.120 187.240 198.440 187.560 ;
        RECT 198.520 187.240 198.840 187.560 ;
        RECT 198.920 187.240 199.240 187.560 ;
        RECT 199.320 187.240 199.640 187.560 ;
        RECT 199.720 187.240 200.040 187.560 ;
        RECT 200.120 187.240 200.440 187.560 ;
        RECT 200.520 187.240 200.840 187.560 ;
        RECT 200.920 187.240 201.240 187.560 ;
        RECT 201.320 187.240 201.640 187.560 ;
        RECT 201.720 187.240 202.040 187.560 ;
        RECT 202.120 187.240 202.440 187.560 ;
        RECT 202.520 187.240 202.840 187.560 ;
        RECT 202.920 187.240 203.240 187.560 ;
        RECT 203.320 187.240 203.640 187.560 ;
        RECT 203.720 187.240 204.040 187.560 ;
        RECT 204.120 187.240 204.440 187.560 ;
        RECT 204.520 187.240 204.840 187.560 ;
        RECT 204.920 187.240 205.240 187.560 ;
        RECT 205.320 187.240 205.640 187.560 ;
        RECT 0.040 186.840 0.360 187.160 ;
        RECT 0.440 186.840 0.760 187.160 ;
        RECT 0.840 186.840 1.160 187.160 ;
        RECT 1.240 186.840 1.560 187.160 ;
        RECT 1.640 186.840 1.960 187.160 ;
        RECT 2.040 186.840 2.360 187.160 ;
        RECT 2.440 186.840 2.760 187.160 ;
        RECT 2.840 186.840 3.160 187.160 ;
        RECT 3.240 186.840 3.560 187.160 ;
        RECT 3.640 186.840 3.960 187.160 ;
        RECT 4.040 186.840 4.360 187.160 ;
        RECT 4.440 186.840 4.760 187.160 ;
        RECT 4.840 186.840 5.160 187.160 ;
        RECT 5.240 186.840 5.560 187.160 ;
        RECT 5.640 186.840 5.960 187.160 ;
        RECT 6.040 186.840 6.360 187.160 ;
        RECT 6.440 186.840 6.760 187.160 ;
        RECT 6.840 186.840 7.160 187.160 ;
        RECT 7.240 186.840 7.560 187.160 ;
        RECT 7.640 186.840 7.960 187.160 ;
        RECT 8.040 186.840 8.360 187.160 ;
        RECT 8.440 186.840 8.760 187.160 ;
        RECT 8.840 186.840 9.160 187.160 ;
        RECT 9.240 186.840 9.560 187.160 ;
        RECT 9.640 186.840 9.960 187.160 ;
        RECT 10.040 186.840 10.360 187.160 ;
        RECT 10.440 186.840 10.760 187.160 ;
        RECT 10.840 186.840 11.160 187.160 ;
        RECT 11.240 186.840 11.560 187.160 ;
        RECT 11.640 186.840 11.960 187.160 ;
        RECT 12.040 186.840 12.360 187.160 ;
        RECT 12.440 186.840 12.760 187.160 ;
        RECT 12.840 186.840 13.160 187.160 ;
        RECT 13.240 186.840 13.560 187.160 ;
        RECT 13.640 186.840 13.960 187.160 ;
        RECT 14.040 186.840 14.360 187.160 ;
        RECT 14.440 186.840 14.760 187.160 ;
        RECT 14.840 186.840 15.160 187.160 ;
        RECT 15.240 186.840 15.560 187.160 ;
        RECT 15.640 186.840 15.960 187.160 ;
        RECT 16.040 186.840 16.360 187.160 ;
        RECT 16.440 186.840 16.760 187.160 ;
        RECT 16.840 186.840 17.160 187.160 ;
        RECT 17.240 186.840 17.560 187.160 ;
        RECT 17.640 186.840 17.960 187.160 ;
        RECT 18.040 186.840 18.360 187.160 ;
        RECT 18.440 186.840 18.760 187.160 ;
        RECT 18.840 186.840 19.160 187.160 ;
        RECT 19.240 186.840 19.560 187.160 ;
        RECT 19.640 186.840 19.960 187.160 ;
        RECT 95.560 186.840 95.880 187.160 ;
        RECT 95.960 186.840 96.280 187.160 ;
        RECT 96.360 186.840 96.680 187.160 ;
        RECT 96.760 186.840 97.080 187.160 ;
        RECT 145.560 186.840 145.880 187.160 ;
        RECT 145.960 186.840 146.280 187.160 ;
        RECT 146.360 186.840 146.680 187.160 ;
        RECT 146.760 186.840 147.080 187.160 ;
        RECT 185.720 186.840 186.040 187.160 ;
        RECT 186.120 186.840 186.440 187.160 ;
        RECT 186.520 186.840 186.840 187.160 ;
        RECT 186.920 186.840 187.240 187.160 ;
        RECT 187.320 186.840 187.640 187.160 ;
        RECT 187.720 186.840 188.040 187.160 ;
        RECT 188.120 186.840 188.440 187.160 ;
        RECT 188.520 186.840 188.840 187.160 ;
        RECT 188.920 186.840 189.240 187.160 ;
        RECT 189.320 186.840 189.640 187.160 ;
        RECT 189.720 186.840 190.040 187.160 ;
        RECT 190.120 186.840 190.440 187.160 ;
        RECT 190.520 186.840 190.840 187.160 ;
        RECT 190.920 186.840 191.240 187.160 ;
        RECT 191.320 186.840 191.640 187.160 ;
        RECT 191.720 186.840 192.040 187.160 ;
        RECT 192.120 186.840 192.440 187.160 ;
        RECT 192.520 186.840 192.840 187.160 ;
        RECT 192.920 186.840 193.240 187.160 ;
        RECT 193.320 186.840 193.640 187.160 ;
        RECT 193.720 186.840 194.040 187.160 ;
        RECT 194.120 186.840 194.440 187.160 ;
        RECT 194.520 186.840 194.840 187.160 ;
        RECT 194.920 186.840 195.240 187.160 ;
        RECT 195.320 186.840 195.640 187.160 ;
        RECT 195.720 186.840 196.040 187.160 ;
        RECT 196.120 186.840 196.440 187.160 ;
        RECT 196.520 186.840 196.840 187.160 ;
        RECT 196.920 186.840 197.240 187.160 ;
        RECT 197.320 186.840 197.640 187.160 ;
        RECT 197.720 186.840 198.040 187.160 ;
        RECT 198.120 186.840 198.440 187.160 ;
        RECT 198.520 186.840 198.840 187.160 ;
        RECT 198.920 186.840 199.240 187.160 ;
        RECT 199.320 186.840 199.640 187.160 ;
        RECT 199.720 186.840 200.040 187.160 ;
        RECT 200.120 186.840 200.440 187.160 ;
        RECT 200.520 186.840 200.840 187.160 ;
        RECT 200.920 186.840 201.240 187.160 ;
        RECT 201.320 186.840 201.640 187.160 ;
        RECT 201.720 186.840 202.040 187.160 ;
        RECT 202.120 186.840 202.440 187.160 ;
        RECT 202.520 186.840 202.840 187.160 ;
        RECT 202.920 186.840 203.240 187.160 ;
        RECT 203.320 186.840 203.640 187.160 ;
        RECT 203.720 186.840 204.040 187.160 ;
        RECT 204.120 186.840 204.440 187.160 ;
        RECT 204.520 186.840 204.840 187.160 ;
        RECT 204.920 186.840 205.240 187.160 ;
        RECT 205.320 186.840 205.640 187.160 ;
        RECT 0.040 186.440 0.360 186.760 ;
        RECT 0.440 186.440 0.760 186.760 ;
        RECT 0.840 186.440 1.160 186.760 ;
        RECT 1.240 186.440 1.560 186.760 ;
        RECT 1.640 186.440 1.960 186.760 ;
        RECT 2.040 186.440 2.360 186.760 ;
        RECT 2.440 186.440 2.760 186.760 ;
        RECT 2.840 186.440 3.160 186.760 ;
        RECT 3.240 186.440 3.560 186.760 ;
        RECT 3.640 186.440 3.960 186.760 ;
        RECT 4.040 186.440 4.360 186.760 ;
        RECT 4.440 186.440 4.760 186.760 ;
        RECT 4.840 186.440 5.160 186.760 ;
        RECT 5.240 186.440 5.560 186.760 ;
        RECT 5.640 186.440 5.960 186.760 ;
        RECT 6.040 186.440 6.360 186.760 ;
        RECT 6.440 186.440 6.760 186.760 ;
        RECT 6.840 186.440 7.160 186.760 ;
        RECT 7.240 186.440 7.560 186.760 ;
        RECT 7.640 186.440 7.960 186.760 ;
        RECT 8.040 186.440 8.360 186.760 ;
        RECT 8.440 186.440 8.760 186.760 ;
        RECT 8.840 186.440 9.160 186.760 ;
        RECT 9.240 186.440 9.560 186.760 ;
        RECT 9.640 186.440 9.960 186.760 ;
        RECT 10.040 186.440 10.360 186.760 ;
        RECT 10.440 186.440 10.760 186.760 ;
        RECT 10.840 186.440 11.160 186.760 ;
        RECT 11.240 186.440 11.560 186.760 ;
        RECT 11.640 186.440 11.960 186.760 ;
        RECT 12.040 186.440 12.360 186.760 ;
        RECT 12.440 186.440 12.760 186.760 ;
        RECT 12.840 186.440 13.160 186.760 ;
        RECT 13.240 186.440 13.560 186.760 ;
        RECT 13.640 186.440 13.960 186.760 ;
        RECT 14.040 186.440 14.360 186.760 ;
        RECT 14.440 186.440 14.760 186.760 ;
        RECT 14.840 186.440 15.160 186.760 ;
        RECT 15.240 186.440 15.560 186.760 ;
        RECT 15.640 186.440 15.960 186.760 ;
        RECT 16.040 186.440 16.360 186.760 ;
        RECT 16.440 186.440 16.760 186.760 ;
        RECT 16.840 186.440 17.160 186.760 ;
        RECT 17.240 186.440 17.560 186.760 ;
        RECT 17.640 186.440 17.960 186.760 ;
        RECT 18.040 186.440 18.360 186.760 ;
        RECT 18.440 186.440 18.760 186.760 ;
        RECT 18.840 186.440 19.160 186.760 ;
        RECT 19.240 186.440 19.560 186.760 ;
        RECT 19.640 186.440 19.960 186.760 ;
        RECT 95.560 186.440 95.880 186.760 ;
        RECT 95.960 186.440 96.280 186.760 ;
        RECT 96.360 186.440 96.680 186.760 ;
        RECT 96.760 186.440 97.080 186.760 ;
        RECT 145.560 186.440 145.880 186.760 ;
        RECT 145.960 186.440 146.280 186.760 ;
        RECT 146.360 186.440 146.680 186.760 ;
        RECT 146.760 186.440 147.080 186.760 ;
        RECT 185.720 186.440 186.040 186.760 ;
        RECT 186.120 186.440 186.440 186.760 ;
        RECT 186.520 186.440 186.840 186.760 ;
        RECT 186.920 186.440 187.240 186.760 ;
        RECT 187.320 186.440 187.640 186.760 ;
        RECT 187.720 186.440 188.040 186.760 ;
        RECT 188.120 186.440 188.440 186.760 ;
        RECT 188.520 186.440 188.840 186.760 ;
        RECT 188.920 186.440 189.240 186.760 ;
        RECT 189.320 186.440 189.640 186.760 ;
        RECT 189.720 186.440 190.040 186.760 ;
        RECT 190.120 186.440 190.440 186.760 ;
        RECT 190.520 186.440 190.840 186.760 ;
        RECT 190.920 186.440 191.240 186.760 ;
        RECT 191.320 186.440 191.640 186.760 ;
        RECT 191.720 186.440 192.040 186.760 ;
        RECT 192.120 186.440 192.440 186.760 ;
        RECT 192.520 186.440 192.840 186.760 ;
        RECT 192.920 186.440 193.240 186.760 ;
        RECT 193.320 186.440 193.640 186.760 ;
        RECT 193.720 186.440 194.040 186.760 ;
        RECT 194.120 186.440 194.440 186.760 ;
        RECT 194.520 186.440 194.840 186.760 ;
        RECT 194.920 186.440 195.240 186.760 ;
        RECT 195.320 186.440 195.640 186.760 ;
        RECT 195.720 186.440 196.040 186.760 ;
        RECT 196.120 186.440 196.440 186.760 ;
        RECT 196.520 186.440 196.840 186.760 ;
        RECT 196.920 186.440 197.240 186.760 ;
        RECT 197.320 186.440 197.640 186.760 ;
        RECT 197.720 186.440 198.040 186.760 ;
        RECT 198.120 186.440 198.440 186.760 ;
        RECT 198.520 186.440 198.840 186.760 ;
        RECT 198.920 186.440 199.240 186.760 ;
        RECT 199.320 186.440 199.640 186.760 ;
        RECT 199.720 186.440 200.040 186.760 ;
        RECT 200.120 186.440 200.440 186.760 ;
        RECT 200.520 186.440 200.840 186.760 ;
        RECT 200.920 186.440 201.240 186.760 ;
        RECT 201.320 186.440 201.640 186.760 ;
        RECT 201.720 186.440 202.040 186.760 ;
        RECT 202.120 186.440 202.440 186.760 ;
        RECT 202.520 186.440 202.840 186.760 ;
        RECT 202.920 186.440 203.240 186.760 ;
        RECT 203.320 186.440 203.640 186.760 ;
        RECT 203.720 186.440 204.040 186.760 ;
        RECT 204.120 186.440 204.440 186.760 ;
        RECT 204.520 186.440 204.840 186.760 ;
        RECT 204.920 186.440 205.240 186.760 ;
        RECT 205.320 186.440 205.640 186.760 ;
        RECT 0.040 186.040 0.360 186.360 ;
        RECT 0.440 186.040 0.760 186.360 ;
        RECT 0.840 186.040 1.160 186.360 ;
        RECT 1.240 186.040 1.560 186.360 ;
        RECT 1.640 186.040 1.960 186.360 ;
        RECT 2.040 186.040 2.360 186.360 ;
        RECT 2.440 186.040 2.760 186.360 ;
        RECT 2.840 186.040 3.160 186.360 ;
        RECT 3.240 186.040 3.560 186.360 ;
        RECT 3.640 186.040 3.960 186.360 ;
        RECT 4.040 186.040 4.360 186.360 ;
        RECT 4.440 186.040 4.760 186.360 ;
        RECT 4.840 186.040 5.160 186.360 ;
        RECT 5.240 186.040 5.560 186.360 ;
        RECT 5.640 186.040 5.960 186.360 ;
        RECT 6.040 186.040 6.360 186.360 ;
        RECT 6.440 186.040 6.760 186.360 ;
        RECT 6.840 186.040 7.160 186.360 ;
        RECT 7.240 186.040 7.560 186.360 ;
        RECT 7.640 186.040 7.960 186.360 ;
        RECT 8.040 186.040 8.360 186.360 ;
        RECT 8.440 186.040 8.760 186.360 ;
        RECT 8.840 186.040 9.160 186.360 ;
        RECT 9.240 186.040 9.560 186.360 ;
        RECT 9.640 186.040 9.960 186.360 ;
        RECT 10.040 186.040 10.360 186.360 ;
        RECT 10.440 186.040 10.760 186.360 ;
        RECT 10.840 186.040 11.160 186.360 ;
        RECT 11.240 186.040 11.560 186.360 ;
        RECT 11.640 186.040 11.960 186.360 ;
        RECT 12.040 186.040 12.360 186.360 ;
        RECT 12.440 186.040 12.760 186.360 ;
        RECT 12.840 186.040 13.160 186.360 ;
        RECT 13.240 186.040 13.560 186.360 ;
        RECT 13.640 186.040 13.960 186.360 ;
        RECT 14.040 186.040 14.360 186.360 ;
        RECT 14.440 186.040 14.760 186.360 ;
        RECT 14.840 186.040 15.160 186.360 ;
        RECT 15.240 186.040 15.560 186.360 ;
        RECT 15.640 186.040 15.960 186.360 ;
        RECT 16.040 186.040 16.360 186.360 ;
        RECT 16.440 186.040 16.760 186.360 ;
        RECT 16.840 186.040 17.160 186.360 ;
        RECT 17.240 186.040 17.560 186.360 ;
        RECT 17.640 186.040 17.960 186.360 ;
        RECT 18.040 186.040 18.360 186.360 ;
        RECT 18.440 186.040 18.760 186.360 ;
        RECT 18.840 186.040 19.160 186.360 ;
        RECT 19.240 186.040 19.560 186.360 ;
        RECT 19.640 186.040 19.960 186.360 ;
        RECT 95.560 186.040 95.880 186.360 ;
        RECT 95.960 186.040 96.280 186.360 ;
        RECT 96.360 186.040 96.680 186.360 ;
        RECT 96.760 186.040 97.080 186.360 ;
        RECT 145.560 186.040 145.880 186.360 ;
        RECT 145.960 186.040 146.280 186.360 ;
        RECT 146.360 186.040 146.680 186.360 ;
        RECT 146.760 186.040 147.080 186.360 ;
        RECT 185.720 186.040 186.040 186.360 ;
        RECT 186.120 186.040 186.440 186.360 ;
        RECT 186.520 186.040 186.840 186.360 ;
        RECT 186.920 186.040 187.240 186.360 ;
        RECT 187.320 186.040 187.640 186.360 ;
        RECT 187.720 186.040 188.040 186.360 ;
        RECT 188.120 186.040 188.440 186.360 ;
        RECT 188.520 186.040 188.840 186.360 ;
        RECT 188.920 186.040 189.240 186.360 ;
        RECT 189.320 186.040 189.640 186.360 ;
        RECT 189.720 186.040 190.040 186.360 ;
        RECT 190.120 186.040 190.440 186.360 ;
        RECT 190.520 186.040 190.840 186.360 ;
        RECT 190.920 186.040 191.240 186.360 ;
        RECT 191.320 186.040 191.640 186.360 ;
        RECT 191.720 186.040 192.040 186.360 ;
        RECT 192.120 186.040 192.440 186.360 ;
        RECT 192.520 186.040 192.840 186.360 ;
        RECT 192.920 186.040 193.240 186.360 ;
        RECT 193.320 186.040 193.640 186.360 ;
        RECT 193.720 186.040 194.040 186.360 ;
        RECT 194.120 186.040 194.440 186.360 ;
        RECT 194.520 186.040 194.840 186.360 ;
        RECT 194.920 186.040 195.240 186.360 ;
        RECT 195.320 186.040 195.640 186.360 ;
        RECT 195.720 186.040 196.040 186.360 ;
        RECT 196.120 186.040 196.440 186.360 ;
        RECT 196.520 186.040 196.840 186.360 ;
        RECT 196.920 186.040 197.240 186.360 ;
        RECT 197.320 186.040 197.640 186.360 ;
        RECT 197.720 186.040 198.040 186.360 ;
        RECT 198.120 186.040 198.440 186.360 ;
        RECT 198.520 186.040 198.840 186.360 ;
        RECT 198.920 186.040 199.240 186.360 ;
        RECT 199.320 186.040 199.640 186.360 ;
        RECT 199.720 186.040 200.040 186.360 ;
        RECT 200.120 186.040 200.440 186.360 ;
        RECT 200.520 186.040 200.840 186.360 ;
        RECT 200.920 186.040 201.240 186.360 ;
        RECT 201.320 186.040 201.640 186.360 ;
        RECT 201.720 186.040 202.040 186.360 ;
        RECT 202.120 186.040 202.440 186.360 ;
        RECT 202.520 186.040 202.840 186.360 ;
        RECT 202.920 186.040 203.240 186.360 ;
        RECT 203.320 186.040 203.640 186.360 ;
        RECT 203.720 186.040 204.040 186.360 ;
        RECT 204.120 186.040 204.440 186.360 ;
        RECT 204.520 186.040 204.840 186.360 ;
        RECT 204.920 186.040 205.240 186.360 ;
        RECT 205.320 186.040 205.640 186.360 ;
        RECT 0.040 185.640 0.360 185.960 ;
        RECT 0.440 185.640 0.760 185.960 ;
        RECT 0.840 185.640 1.160 185.960 ;
        RECT 1.240 185.640 1.560 185.960 ;
        RECT 1.640 185.640 1.960 185.960 ;
        RECT 2.040 185.640 2.360 185.960 ;
        RECT 2.440 185.640 2.760 185.960 ;
        RECT 2.840 185.640 3.160 185.960 ;
        RECT 3.240 185.640 3.560 185.960 ;
        RECT 3.640 185.640 3.960 185.960 ;
        RECT 4.040 185.640 4.360 185.960 ;
        RECT 4.440 185.640 4.760 185.960 ;
        RECT 4.840 185.640 5.160 185.960 ;
        RECT 5.240 185.640 5.560 185.960 ;
        RECT 5.640 185.640 5.960 185.960 ;
        RECT 6.040 185.640 6.360 185.960 ;
        RECT 6.440 185.640 6.760 185.960 ;
        RECT 6.840 185.640 7.160 185.960 ;
        RECT 7.240 185.640 7.560 185.960 ;
        RECT 7.640 185.640 7.960 185.960 ;
        RECT 8.040 185.640 8.360 185.960 ;
        RECT 8.440 185.640 8.760 185.960 ;
        RECT 8.840 185.640 9.160 185.960 ;
        RECT 9.240 185.640 9.560 185.960 ;
        RECT 9.640 185.640 9.960 185.960 ;
        RECT 10.040 185.640 10.360 185.960 ;
        RECT 10.440 185.640 10.760 185.960 ;
        RECT 10.840 185.640 11.160 185.960 ;
        RECT 11.240 185.640 11.560 185.960 ;
        RECT 11.640 185.640 11.960 185.960 ;
        RECT 12.040 185.640 12.360 185.960 ;
        RECT 12.440 185.640 12.760 185.960 ;
        RECT 12.840 185.640 13.160 185.960 ;
        RECT 13.240 185.640 13.560 185.960 ;
        RECT 13.640 185.640 13.960 185.960 ;
        RECT 14.040 185.640 14.360 185.960 ;
        RECT 14.440 185.640 14.760 185.960 ;
        RECT 14.840 185.640 15.160 185.960 ;
        RECT 15.240 185.640 15.560 185.960 ;
        RECT 15.640 185.640 15.960 185.960 ;
        RECT 16.040 185.640 16.360 185.960 ;
        RECT 16.440 185.640 16.760 185.960 ;
        RECT 16.840 185.640 17.160 185.960 ;
        RECT 17.240 185.640 17.560 185.960 ;
        RECT 17.640 185.640 17.960 185.960 ;
        RECT 18.040 185.640 18.360 185.960 ;
        RECT 18.440 185.640 18.760 185.960 ;
        RECT 18.840 185.640 19.160 185.960 ;
        RECT 19.240 185.640 19.560 185.960 ;
        RECT 19.640 185.640 19.960 185.960 ;
        RECT 95.560 185.640 95.880 185.960 ;
        RECT 95.960 185.640 96.280 185.960 ;
        RECT 96.360 185.640 96.680 185.960 ;
        RECT 96.760 185.640 97.080 185.960 ;
        RECT 145.560 185.640 145.880 185.960 ;
        RECT 145.960 185.640 146.280 185.960 ;
        RECT 146.360 185.640 146.680 185.960 ;
        RECT 146.760 185.640 147.080 185.960 ;
        RECT 185.720 185.640 186.040 185.960 ;
        RECT 186.120 185.640 186.440 185.960 ;
        RECT 186.520 185.640 186.840 185.960 ;
        RECT 186.920 185.640 187.240 185.960 ;
        RECT 187.320 185.640 187.640 185.960 ;
        RECT 187.720 185.640 188.040 185.960 ;
        RECT 188.120 185.640 188.440 185.960 ;
        RECT 188.520 185.640 188.840 185.960 ;
        RECT 188.920 185.640 189.240 185.960 ;
        RECT 189.320 185.640 189.640 185.960 ;
        RECT 189.720 185.640 190.040 185.960 ;
        RECT 190.120 185.640 190.440 185.960 ;
        RECT 190.520 185.640 190.840 185.960 ;
        RECT 190.920 185.640 191.240 185.960 ;
        RECT 191.320 185.640 191.640 185.960 ;
        RECT 191.720 185.640 192.040 185.960 ;
        RECT 192.120 185.640 192.440 185.960 ;
        RECT 192.520 185.640 192.840 185.960 ;
        RECT 192.920 185.640 193.240 185.960 ;
        RECT 193.320 185.640 193.640 185.960 ;
        RECT 193.720 185.640 194.040 185.960 ;
        RECT 194.120 185.640 194.440 185.960 ;
        RECT 194.520 185.640 194.840 185.960 ;
        RECT 194.920 185.640 195.240 185.960 ;
        RECT 195.320 185.640 195.640 185.960 ;
        RECT 195.720 185.640 196.040 185.960 ;
        RECT 196.120 185.640 196.440 185.960 ;
        RECT 196.520 185.640 196.840 185.960 ;
        RECT 196.920 185.640 197.240 185.960 ;
        RECT 197.320 185.640 197.640 185.960 ;
        RECT 197.720 185.640 198.040 185.960 ;
        RECT 198.120 185.640 198.440 185.960 ;
        RECT 198.520 185.640 198.840 185.960 ;
        RECT 198.920 185.640 199.240 185.960 ;
        RECT 199.320 185.640 199.640 185.960 ;
        RECT 199.720 185.640 200.040 185.960 ;
        RECT 200.120 185.640 200.440 185.960 ;
        RECT 200.520 185.640 200.840 185.960 ;
        RECT 200.920 185.640 201.240 185.960 ;
        RECT 201.320 185.640 201.640 185.960 ;
        RECT 201.720 185.640 202.040 185.960 ;
        RECT 202.120 185.640 202.440 185.960 ;
        RECT 202.520 185.640 202.840 185.960 ;
        RECT 202.920 185.640 203.240 185.960 ;
        RECT 203.320 185.640 203.640 185.960 ;
        RECT 203.720 185.640 204.040 185.960 ;
        RECT 204.120 185.640 204.440 185.960 ;
        RECT 204.520 185.640 204.840 185.960 ;
        RECT 204.920 185.640 205.240 185.960 ;
        RECT 205.320 185.640 205.640 185.960 ;
        RECT 0.040 185.240 0.360 185.560 ;
        RECT 0.440 185.240 0.760 185.560 ;
        RECT 0.840 185.240 1.160 185.560 ;
        RECT 1.240 185.240 1.560 185.560 ;
        RECT 1.640 185.240 1.960 185.560 ;
        RECT 2.040 185.240 2.360 185.560 ;
        RECT 2.440 185.240 2.760 185.560 ;
        RECT 2.840 185.240 3.160 185.560 ;
        RECT 3.240 185.240 3.560 185.560 ;
        RECT 3.640 185.240 3.960 185.560 ;
        RECT 4.040 185.240 4.360 185.560 ;
        RECT 4.440 185.240 4.760 185.560 ;
        RECT 4.840 185.240 5.160 185.560 ;
        RECT 5.240 185.240 5.560 185.560 ;
        RECT 5.640 185.240 5.960 185.560 ;
        RECT 6.040 185.240 6.360 185.560 ;
        RECT 6.440 185.240 6.760 185.560 ;
        RECT 6.840 185.240 7.160 185.560 ;
        RECT 7.240 185.240 7.560 185.560 ;
        RECT 7.640 185.240 7.960 185.560 ;
        RECT 8.040 185.240 8.360 185.560 ;
        RECT 8.440 185.240 8.760 185.560 ;
        RECT 8.840 185.240 9.160 185.560 ;
        RECT 9.240 185.240 9.560 185.560 ;
        RECT 9.640 185.240 9.960 185.560 ;
        RECT 10.040 185.240 10.360 185.560 ;
        RECT 10.440 185.240 10.760 185.560 ;
        RECT 10.840 185.240 11.160 185.560 ;
        RECT 11.240 185.240 11.560 185.560 ;
        RECT 11.640 185.240 11.960 185.560 ;
        RECT 12.040 185.240 12.360 185.560 ;
        RECT 12.440 185.240 12.760 185.560 ;
        RECT 12.840 185.240 13.160 185.560 ;
        RECT 13.240 185.240 13.560 185.560 ;
        RECT 13.640 185.240 13.960 185.560 ;
        RECT 14.040 185.240 14.360 185.560 ;
        RECT 14.440 185.240 14.760 185.560 ;
        RECT 14.840 185.240 15.160 185.560 ;
        RECT 15.240 185.240 15.560 185.560 ;
        RECT 15.640 185.240 15.960 185.560 ;
        RECT 16.040 185.240 16.360 185.560 ;
        RECT 16.440 185.240 16.760 185.560 ;
        RECT 16.840 185.240 17.160 185.560 ;
        RECT 17.240 185.240 17.560 185.560 ;
        RECT 17.640 185.240 17.960 185.560 ;
        RECT 18.040 185.240 18.360 185.560 ;
        RECT 18.440 185.240 18.760 185.560 ;
        RECT 18.840 185.240 19.160 185.560 ;
        RECT 19.240 185.240 19.560 185.560 ;
        RECT 19.640 185.240 19.960 185.560 ;
        RECT 95.560 185.240 95.880 185.560 ;
        RECT 95.960 185.240 96.280 185.560 ;
        RECT 96.360 185.240 96.680 185.560 ;
        RECT 96.760 185.240 97.080 185.560 ;
        RECT 145.560 185.240 145.880 185.560 ;
        RECT 145.960 185.240 146.280 185.560 ;
        RECT 146.360 185.240 146.680 185.560 ;
        RECT 146.760 185.240 147.080 185.560 ;
        RECT 185.720 185.240 186.040 185.560 ;
        RECT 186.120 185.240 186.440 185.560 ;
        RECT 186.520 185.240 186.840 185.560 ;
        RECT 186.920 185.240 187.240 185.560 ;
        RECT 187.320 185.240 187.640 185.560 ;
        RECT 187.720 185.240 188.040 185.560 ;
        RECT 188.120 185.240 188.440 185.560 ;
        RECT 188.520 185.240 188.840 185.560 ;
        RECT 188.920 185.240 189.240 185.560 ;
        RECT 189.320 185.240 189.640 185.560 ;
        RECT 189.720 185.240 190.040 185.560 ;
        RECT 190.120 185.240 190.440 185.560 ;
        RECT 190.520 185.240 190.840 185.560 ;
        RECT 190.920 185.240 191.240 185.560 ;
        RECT 191.320 185.240 191.640 185.560 ;
        RECT 191.720 185.240 192.040 185.560 ;
        RECT 192.120 185.240 192.440 185.560 ;
        RECT 192.520 185.240 192.840 185.560 ;
        RECT 192.920 185.240 193.240 185.560 ;
        RECT 193.320 185.240 193.640 185.560 ;
        RECT 193.720 185.240 194.040 185.560 ;
        RECT 194.120 185.240 194.440 185.560 ;
        RECT 194.520 185.240 194.840 185.560 ;
        RECT 194.920 185.240 195.240 185.560 ;
        RECT 195.320 185.240 195.640 185.560 ;
        RECT 195.720 185.240 196.040 185.560 ;
        RECT 196.120 185.240 196.440 185.560 ;
        RECT 196.520 185.240 196.840 185.560 ;
        RECT 196.920 185.240 197.240 185.560 ;
        RECT 197.320 185.240 197.640 185.560 ;
        RECT 197.720 185.240 198.040 185.560 ;
        RECT 198.120 185.240 198.440 185.560 ;
        RECT 198.520 185.240 198.840 185.560 ;
        RECT 198.920 185.240 199.240 185.560 ;
        RECT 199.320 185.240 199.640 185.560 ;
        RECT 199.720 185.240 200.040 185.560 ;
        RECT 200.120 185.240 200.440 185.560 ;
        RECT 200.520 185.240 200.840 185.560 ;
        RECT 200.920 185.240 201.240 185.560 ;
        RECT 201.320 185.240 201.640 185.560 ;
        RECT 201.720 185.240 202.040 185.560 ;
        RECT 202.120 185.240 202.440 185.560 ;
        RECT 202.520 185.240 202.840 185.560 ;
        RECT 202.920 185.240 203.240 185.560 ;
        RECT 203.320 185.240 203.640 185.560 ;
        RECT 203.720 185.240 204.040 185.560 ;
        RECT 204.120 185.240 204.440 185.560 ;
        RECT 204.520 185.240 204.840 185.560 ;
        RECT 204.920 185.240 205.240 185.560 ;
        RECT 205.320 185.240 205.640 185.560 ;
        RECT 0.040 19.640 0.360 19.960 ;
        RECT 0.440 19.640 0.760 19.960 ;
        RECT 0.840 19.640 1.160 19.960 ;
        RECT 1.240 19.640 1.560 19.960 ;
        RECT 1.640 19.640 1.960 19.960 ;
        RECT 2.040 19.640 2.360 19.960 ;
        RECT 2.440 19.640 2.760 19.960 ;
        RECT 2.840 19.640 3.160 19.960 ;
        RECT 3.240 19.640 3.560 19.960 ;
        RECT 3.640 19.640 3.960 19.960 ;
        RECT 4.040 19.640 4.360 19.960 ;
        RECT 4.440 19.640 4.760 19.960 ;
        RECT 4.840 19.640 5.160 19.960 ;
        RECT 5.240 19.640 5.560 19.960 ;
        RECT 5.640 19.640 5.960 19.960 ;
        RECT 6.040 19.640 6.360 19.960 ;
        RECT 6.440 19.640 6.760 19.960 ;
        RECT 6.840 19.640 7.160 19.960 ;
        RECT 7.240 19.640 7.560 19.960 ;
        RECT 7.640 19.640 7.960 19.960 ;
        RECT 8.040 19.640 8.360 19.960 ;
        RECT 8.440 19.640 8.760 19.960 ;
        RECT 8.840 19.640 9.160 19.960 ;
        RECT 9.240 19.640 9.560 19.960 ;
        RECT 9.640 19.640 9.960 19.960 ;
        RECT 10.040 19.640 10.360 19.960 ;
        RECT 10.440 19.640 10.760 19.960 ;
        RECT 10.840 19.640 11.160 19.960 ;
        RECT 11.240 19.640 11.560 19.960 ;
        RECT 11.640 19.640 11.960 19.960 ;
        RECT 12.040 19.640 12.360 19.960 ;
        RECT 12.440 19.640 12.760 19.960 ;
        RECT 12.840 19.640 13.160 19.960 ;
        RECT 13.240 19.640 13.560 19.960 ;
        RECT 13.640 19.640 13.960 19.960 ;
        RECT 14.040 19.640 14.360 19.960 ;
        RECT 14.440 19.640 14.760 19.960 ;
        RECT 14.840 19.640 15.160 19.960 ;
        RECT 15.240 19.640 15.560 19.960 ;
        RECT 15.640 19.640 15.960 19.960 ;
        RECT 16.040 19.640 16.360 19.960 ;
        RECT 16.440 19.640 16.760 19.960 ;
        RECT 16.840 19.640 17.160 19.960 ;
        RECT 17.240 19.640 17.560 19.960 ;
        RECT 17.640 19.640 17.960 19.960 ;
        RECT 18.040 19.640 18.360 19.960 ;
        RECT 18.440 19.640 18.760 19.960 ;
        RECT 18.840 19.640 19.160 19.960 ;
        RECT 19.240 19.640 19.560 19.960 ;
        RECT 19.640 19.640 19.960 19.960 ;
        RECT 95.560 19.640 95.880 19.960 ;
        RECT 95.960 19.640 96.280 19.960 ;
        RECT 96.360 19.640 96.680 19.960 ;
        RECT 96.760 19.640 97.080 19.960 ;
        RECT 145.560 19.640 145.880 19.960 ;
        RECT 145.960 19.640 146.280 19.960 ;
        RECT 146.360 19.640 146.680 19.960 ;
        RECT 146.760 19.640 147.080 19.960 ;
        RECT 185.720 19.640 186.040 19.960 ;
        RECT 186.120 19.640 186.440 19.960 ;
        RECT 186.520 19.640 186.840 19.960 ;
        RECT 186.920 19.640 187.240 19.960 ;
        RECT 187.320 19.640 187.640 19.960 ;
        RECT 187.720 19.640 188.040 19.960 ;
        RECT 188.120 19.640 188.440 19.960 ;
        RECT 188.520 19.640 188.840 19.960 ;
        RECT 188.920 19.640 189.240 19.960 ;
        RECT 189.320 19.640 189.640 19.960 ;
        RECT 189.720 19.640 190.040 19.960 ;
        RECT 190.120 19.640 190.440 19.960 ;
        RECT 190.520 19.640 190.840 19.960 ;
        RECT 190.920 19.640 191.240 19.960 ;
        RECT 191.320 19.640 191.640 19.960 ;
        RECT 191.720 19.640 192.040 19.960 ;
        RECT 192.120 19.640 192.440 19.960 ;
        RECT 192.520 19.640 192.840 19.960 ;
        RECT 192.920 19.640 193.240 19.960 ;
        RECT 193.320 19.640 193.640 19.960 ;
        RECT 193.720 19.640 194.040 19.960 ;
        RECT 194.120 19.640 194.440 19.960 ;
        RECT 194.520 19.640 194.840 19.960 ;
        RECT 194.920 19.640 195.240 19.960 ;
        RECT 195.320 19.640 195.640 19.960 ;
        RECT 195.720 19.640 196.040 19.960 ;
        RECT 196.120 19.640 196.440 19.960 ;
        RECT 196.520 19.640 196.840 19.960 ;
        RECT 196.920 19.640 197.240 19.960 ;
        RECT 197.320 19.640 197.640 19.960 ;
        RECT 197.720 19.640 198.040 19.960 ;
        RECT 198.120 19.640 198.440 19.960 ;
        RECT 198.520 19.640 198.840 19.960 ;
        RECT 198.920 19.640 199.240 19.960 ;
        RECT 199.320 19.640 199.640 19.960 ;
        RECT 199.720 19.640 200.040 19.960 ;
        RECT 200.120 19.640 200.440 19.960 ;
        RECT 200.520 19.640 200.840 19.960 ;
        RECT 200.920 19.640 201.240 19.960 ;
        RECT 201.320 19.640 201.640 19.960 ;
        RECT 201.720 19.640 202.040 19.960 ;
        RECT 202.120 19.640 202.440 19.960 ;
        RECT 202.520 19.640 202.840 19.960 ;
        RECT 202.920 19.640 203.240 19.960 ;
        RECT 203.320 19.640 203.640 19.960 ;
        RECT 203.720 19.640 204.040 19.960 ;
        RECT 204.120 19.640 204.440 19.960 ;
        RECT 204.520 19.640 204.840 19.960 ;
        RECT 204.920 19.640 205.240 19.960 ;
        RECT 205.320 19.640 205.640 19.960 ;
        RECT 0.040 19.240 0.360 19.560 ;
        RECT 0.440 19.240 0.760 19.560 ;
        RECT 0.840 19.240 1.160 19.560 ;
        RECT 1.240 19.240 1.560 19.560 ;
        RECT 1.640 19.240 1.960 19.560 ;
        RECT 2.040 19.240 2.360 19.560 ;
        RECT 2.440 19.240 2.760 19.560 ;
        RECT 2.840 19.240 3.160 19.560 ;
        RECT 3.240 19.240 3.560 19.560 ;
        RECT 3.640 19.240 3.960 19.560 ;
        RECT 4.040 19.240 4.360 19.560 ;
        RECT 4.440 19.240 4.760 19.560 ;
        RECT 4.840 19.240 5.160 19.560 ;
        RECT 5.240 19.240 5.560 19.560 ;
        RECT 5.640 19.240 5.960 19.560 ;
        RECT 6.040 19.240 6.360 19.560 ;
        RECT 6.440 19.240 6.760 19.560 ;
        RECT 6.840 19.240 7.160 19.560 ;
        RECT 7.240 19.240 7.560 19.560 ;
        RECT 7.640 19.240 7.960 19.560 ;
        RECT 8.040 19.240 8.360 19.560 ;
        RECT 8.440 19.240 8.760 19.560 ;
        RECT 8.840 19.240 9.160 19.560 ;
        RECT 9.240 19.240 9.560 19.560 ;
        RECT 9.640 19.240 9.960 19.560 ;
        RECT 10.040 19.240 10.360 19.560 ;
        RECT 10.440 19.240 10.760 19.560 ;
        RECT 10.840 19.240 11.160 19.560 ;
        RECT 11.240 19.240 11.560 19.560 ;
        RECT 11.640 19.240 11.960 19.560 ;
        RECT 12.040 19.240 12.360 19.560 ;
        RECT 12.440 19.240 12.760 19.560 ;
        RECT 12.840 19.240 13.160 19.560 ;
        RECT 13.240 19.240 13.560 19.560 ;
        RECT 13.640 19.240 13.960 19.560 ;
        RECT 14.040 19.240 14.360 19.560 ;
        RECT 14.440 19.240 14.760 19.560 ;
        RECT 14.840 19.240 15.160 19.560 ;
        RECT 15.240 19.240 15.560 19.560 ;
        RECT 15.640 19.240 15.960 19.560 ;
        RECT 16.040 19.240 16.360 19.560 ;
        RECT 16.440 19.240 16.760 19.560 ;
        RECT 16.840 19.240 17.160 19.560 ;
        RECT 17.240 19.240 17.560 19.560 ;
        RECT 17.640 19.240 17.960 19.560 ;
        RECT 18.040 19.240 18.360 19.560 ;
        RECT 18.440 19.240 18.760 19.560 ;
        RECT 18.840 19.240 19.160 19.560 ;
        RECT 19.240 19.240 19.560 19.560 ;
        RECT 19.640 19.240 19.960 19.560 ;
        RECT 95.560 19.240 95.880 19.560 ;
        RECT 95.960 19.240 96.280 19.560 ;
        RECT 96.360 19.240 96.680 19.560 ;
        RECT 96.760 19.240 97.080 19.560 ;
        RECT 145.560 19.240 145.880 19.560 ;
        RECT 145.960 19.240 146.280 19.560 ;
        RECT 146.360 19.240 146.680 19.560 ;
        RECT 146.760 19.240 147.080 19.560 ;
        RECT 185.720 19.240 186.040 19.560 ;
        RECT 186.120 19.240 186.440 19.560 ;
        RECT 186.520 19.240 186.840 19.560 ;
        RECT 186.920 19.240 187.240 19.560 ;
        RECT 187.320 19.240 187.640 19.560 ;
        RECT 187.720 19.240 188.040 19.560 ;
        RECT 188.120 19.240 188.440 19.560 ;
        RECT 188.520 19.240 188.840 19.560 ;
        RECT 188.920 19.240 189.240 19.560 ;
        RECT 189.320 19.240 189.640 19.560 ;
        RECT 189.720 19.240 190.040 19.560 ;
        RECT 190.120 19.240 190.440 19.560 ;
        RECT 190.520 19.240 190.840 19.560 ;
        RECT 190.920 19.240 191.240 19.560 ;
        RECT 191.320 19.240 191.640 19.560 ;
        RECT 191.720 19.240 192.040 19.560 ;
        RECT 192.120 19.240 192.440 19.560 ;
        RECT 192.520 19.240 192.840 19.560 ;
        RECT 192.920 19.240 193.240 19.560 ;
        RECT 193.320 19.240 193.640 19.560 ;
        RECT 193.720 19.240 194.040 19.560 ;
        RECT 194.120 19.240 194.440 19.560 ;
        RECT 194.520 19.240 194.840 19.560 ;
        RECT 194.920 19.240 195.240 19.560 ;
        RECT 195.320 19.240 195.640 19.560 ;
        RECT 195.720 19.240 196.040 19.560 ;
        RECT 196.120 19.240 196.440 19.560 ;
        RECT 196.520 19.240 196.840 19.560 ;
        RECT 196.920 19.240 197.240 19.560 ;
        RECT 197.320 19.240 197.640 19.560 ;
        RECT 197.720 19.240 198.040 19.560 ;
        RECT 198.120 19.240 198.440 19.560 ;
        RECT 198.520 19.240 198.840 19.560 ;
        RECT 198.920 19.240 199.240 19.560 ;
        RECT 199.320 19.240 199.640 19.560 ;
        RECT 199.720 19.240 200.040 19.560 ;
        RECT 200.120 19.240 200.440 19.560 ;
        RECT 200.520 19.240 200.840 19.560 ;
        RECT 200.920 19.240 201.240 19.560 ;
        RECT 201.320 19.240 201.640 19.560 ;
        RECT 201.720 19.240 202.040 19.560 ;
        RECT 202.120 19.240 202.440 19.560 ;
        RECT 202.520 19.240 202.840 19.560 ;
        RECT 202.920 19.240 203.240 19.560 ;
        RECT 203.320 19.240 203.640 19.560 ;
        RECT 203.720 19.240 204.040 19.560 ;
        RECT 204.120 19.240 204.440 19.560 ;
        RECT 204.520 19.240 204.840 19.560 ;
        RECT 204.920 19.240 205.240 19.560 ;
        RECT 205.320 19.240 205.640 19.560 ;
        RECT 0.040 18.840 0.360 19.160 ;
        RECT 0.440 18.840 0.760 19.160 ;
        RECT 0.840 18.840 1.160 19.160 ;
        RECT 1.240 18.840 1.560 19.160 ;
        RECT 1.640 18.840 1.960 19.160 ;
        RECT 2.040 18.840 2.360 19.160 ;
        RECT 2.440 18.840 2.760 19.160 ;
        RECT 2.840 18.840 3.160 19.160 ;
        RECT 3.240 18.840 3.560 19.160 ;
        RECT 3.640 18.840 3.960 19.160 ;
        RECT 4.040 18.840 4.360 19.160 ;
        RECT 4.440 18.840 4.760 19.160 ;
        RECT 4.840 18.840 5.160 19.160 ;
        RECT 5.240 18.840 5.560 19.160 ;
        RECT 5.640 18.840 5.960 19.160 ;
        RECT 6.040 18.840 6.360 19.160 ;
        RECT 6.440 18.840 6.760 19.160 ;
        RECT 6.840 18.840 7.160 19.160 ;
        RECT 7.240 18.840 7.560 19.160 ;
        RECT 7.640 18.840 7.960 19.160 ;
        RECT 8.040 18.840 8.360 19.160 ;
        RECT 8.440 18.840 8.760 19.160 ;
        RECT 8.840 18.840 9.160 19.160 ;
        RECT 9.240 18.840 9.560 19.160 ;
        RECT 9.640 18.840 9.960 19.160 ;
        RECT 10.040 18.840 10.360 19.160 ;
        RECT 10.440 18.840 10.760 19.160 ;
        RECT 10.840 18.840 11.160 19.160 ;
        RECT 11.240 18.840 11.560 19.160 ;
        RECT 11.640 18.840 11.960 19.160 ;
        RECT 12.040 18.840 12.360 19.160 ;
        RECT 12.440 18.840 12.760 19.160 ;
        RECT 12.840 18.840 13.160 19.160 ;
        RECT 13.240 18.840 13.560 19.160 ;
        RECT 13.640 18.840 13.960 19.160 ;
        RECT 14.040 18.840 14.360 19.160 ;
        RECT 14.440 18.840 14.760 19.160 ;
        RECT 14.840 18.840 15.160 19.160 ;
        RECT 15.240 18.840 15.560 19.160 ;
        RECT 15.640 18.840 15.960 19.160 ;
        RECT 16.040 18.840 16.360 19.160 ;
        RECT 16.440 18.840 16.760 19.160 ;
        RECT 16.840 18.840 17.160 19.160 ;
        RECT 17.240 18.840 17.560 19.160 ;
        RECT 17.640 18.840 17.960 19.160 ;
        RECT 18.040 18.840 18.360 19.160 ;
        RECT 18.440 18.840 18.760 19.160 ;
        RECT 18.840 18.840 19.160 19.160 ;
        RECT 19.240 18.840 19.560 19.160 ;
        RECT 19.640 18.840 19.960 19.160 ;
        RECT 95.560 18.840 95.880 19.160 ;
        RECT 95.960 18.840 96.280 19.160 ;
        RECT 96.360 18.840 96.680 19.160 ;
        RECT 96.760 18.840 97.080 19.160 ;
        RECT 145.560 18.840 145.880 19.160 ;
        RECT 145.960 18.840 146.280 19.160 ;
        RECT 146.360 18.840 146.680 19.160 ;
        RECT 146.760 18.840 147.080 19.160 ;
        RECT 185.720 18.840 186.040 19.160 ;
        RECT 186.120 18.840 186.440 19.160 ;
        RECT 186.520 18.840 186.840 19.160 ;
        RECT 186.920 18.840 187.240 19.160 ;
        RECT 187.320 18.840 187.640 19.160 ;
        RECT 187.720 18.840 188.040 19.160 ;
        RECT 188.120 18.840 188.440 19.160 ;
        RECT 188.520 18.840 188.840 19.160 ;
        RECT 188.920 18.840 189.240 19.160 ;
        RECT 189.320 18.840 189.640 19.160 ;
        RECT 189.720 18.840 190.040 19.160 ;
        RECT 190.120 18.840 190.440 19.160 ;
        RECT 190.520 18.840 190.840 19.160 ;
        RECT 190.920 18.840 191.240 19.160 ;
        RECT 191.320 18.840 191.640 19.160 ;
        RECT 191.720 18.840 192.040 19.160 ;
        RECT 192.120 18.840 192.440 19.160 ;
        RECT 192.520 18.840 192.840 19.160 ;
        RECT 192.920 18.840 193.240 19.160 ;
        RECT 193.320 18.840 193.640 19.160 ;
        RECT 193.720 18.840 194.040 19.160 ;
        RECT 194.120 18.840 194.440 19.160 ;
        RECT 194.520 18.840 194.840 19.160 ;
        RECT 194.920 18.840 195.240 19.160 ;
        RECT 195.320 18.840 195.640 19.160 ;
        RECT 195.720 18.840 196.040 19.160 ;
        RECT 196.120 18.840 196.440 19.160 ;
        RECT 196.520 18.840 196.840 19.160 ;
        RECT 196.920 18.840 197.240 19.160 ;
        RECT 197.320 18.840 197.640 19.160 ;
        RECT 197.720 18.840 198.040 19.160 ;
        RECT 198.120 18.840 198.440 19.160 ;
        RECT 198.520 18.840 198.840 19.160 ;
        RECT 198.920 18.840 199.240 19.160 ;
        RECT 199.320 18.840 199.640 19.160 ;
        RECT 199.720 18.840 200.040 19.160 ;
        RECT 200.120 18.840 200.440 19.160 ;
        RECT 200.520 18.840 200.840 19.160 ;
        RECT 200.920 18.840 201.240 19.160 ;
        RECT 201.320 18.840 201.640 19.160 ;
        RECT 201.720 18.840 202.040 19.160 ;
        RECT 202.120 18.840 202.440 19.160 ;
        RECT 202.520 18.840 202.840 19.160 ;
        RECT 202.920 18.840 203.240 19.160 ;
        RECT 203.320 18.840 203.640 19.160 ;
        RECT 203.720 18.840 204.040 19.160 ;
        RECT 204.120 18.840 204.440 19.160 ;
        RECT 204.520 18.840 204.840 19.160 ;
        RECT 204.920 18.840 205.240 19.160 ;
        RECT 205.320 18.840 205.640 19.160 ;
        RECT 0.040 18.440 0.360 18.760 ;
        RECT 0.440 18.440 0.760 18.760 ;
        RECT 0.840 18.440 1.160 18.760 ;
        RECT 1.240 18.440 1.560 18.760 ;
        RECT 1.640 18.440 1.960 18.760 ;
        RECT 2.040 18.440 2.360 18.760 ;
        RECT 2.440 18.440 2.760 18.760 ;
        RECT 2.840 18.440 3.160 18.760 ;
        RECT 3.240 18.440 3.560 18.760 ;
        RECT 3.640 18.440 3.960 18.760 ;
        RECT 4.040 18.440 4.360 18.760 ;
        RECT 4.440 18.440 4.760 18.760 ;
        RECT 4.840 18.440 5.160 18.760 ;
        RECT 5.240 18.440 5.560 18.760 ;
        RECT 5.640 18.440 5.960 18.760 ;
        RECT 6.040 18.440 6.360 18.760 ;
        RECT 6.440 18.440 6.760 18.760 ;
        RECT 6.840 18.440 7.160 18.760 ;
        RECT 7.240 18.440 7.560 18.760 ;
        RECT 7.640 18.440 7.960 18.760 ;
        RECT 8.040 18.440 8.360 18.760 ;
        RECT 8.440 18.440 8.760 18.760 ;
        RECT 8.840 18.440 9.160 18.760 ;
        RECT 9.240 18.440 9.560 18.760 ;
        RECT 9.640 18.440 9.960 18.760 ;
        RECT 10.040 18.440 10.360 18.760 ;
        RECT 10.440 18.440 10.760 18.760 ;
        RECT 10.840 18.440 11.160 18.760 ;
        RECT 11.240 18.440 11.560 18.760 ;
        RECT 11.640 18.440 11.960 18.760 ;
        RECT 12.040 18.440 12.360 18.760 ;
        RECT 12.440 18.440 12.760 18.760 ;
        RECT 12.840 18.440 13.160 18.760 ;
        RECT 13.240 18.440 13.560 18.760 ;
        RECT 13.640 18.440 13.960 18.760 ;
        RECT 14.040 18.440 14.360 18.760 ;
        RECT 14.440 18.440 14.760 18.760 ;
        RECT 14.840 18.440 15.160 18.760 ;
        RECT 15.240 18.440 15.560 18.760 ;
        RECT 15.640 18.440 15.960 18.760 ;
        RECT 16.040 18.440 16.360 18.760 ;
        RECT 16.440 18.440 16.760 18.760 ;
        RECT 16.840 18.440 17.160 18.760 ;
        RECT 17.240 18.440 17.560 18.760 ;
        RECT 17.640 18.440 17.960 18.760 ;
        RECT 18.040 18.440 18.360 18.760 ;
        RECT 18.440 18.440 18.760 18.760 ;
        RECT 18.840 18.440 19.160 18.760 ;
        RECT 19.240 18.440 19.560 18.760 ;
        RECT 19.640 18.440 19.960 18.760 ;
        RECT 95.560 18.440 95.880 18.760 ;
        RECT 95.960 18.440 96.280 18.760 ;
        RECT 96.360 18.440 96.680 18.760 ;
        RECT 96.760 18.440 97.080 18.760 ;
        RECT 145.560 18.440 145.880 18.760 ;
        RECT 145.960 18.440 146.280 18.760 ;
        RECT 146.360 18.440 146.680 18.760 ;
        RECT 146.760 18.440 147.080 18.760 ;
        RECT 185.720 18.440 186.040 18.760 ;
        RECT 186.120 18.440 186.440 18.760 ;
        RECT 186.520 18.440 186.840 18.760 ;
        RECT 186.920 18.440 187.240 18.760 ;
        RECT 187.320 18.440 187.640 18.760 ;
        RECT 187.720 18.440 188.040 18.760 ;
        RECT 188.120 18.440 188.440 18.760 ;
        RECT 188.520 18.440 188.840 18.760 ;
        RECT 188.920 18.440 189.240 18.760 ;
        RECT 189.320 18.440 189.640 18.760 ;
        RECT 189.720 18.440 190.040 18.760 ;
        RECT 190.120 18.440 190.440 18.760 ;
        RECT 190.520 18.440 190.840 18.760 ;
        RECT 190.920 18.440 191.240 18.760 ;
        RECT 191.320 18.440 191.640 18.760 ;
        RECT 191.720 18.440 192.040 18.760 ;
        RECT 192.120 18.440 192.440 18.760 ;
        RECT 192.520 18.440 192.840 18.760 ;
        RECT 192.920 18.440 193.240 18.760 ;
        RECT 193.320 18.440 193.640 18.760 ;
        RECT 193.720 18.440 194.040 18.760 ;
        RECT 194.120 18.440 194.440 18.760 ;
        RECT 194.520 18.440 194.840 18.760 ;
        RECT 194.920 18.440 195.240 18.760 ;
        RECT 195.320 18.440 195.640 18.760 ;
        RECT 195.720 18.440 196.040 18.760 ;
        RECT 196.120 18.440 196.440 18.760 ;
        RECT 196.520 18.440 196.840 18.760 ;
        RECT 196.920 18.440 197.240 18.760 ;
        RECT 197.320 18.440 197.640 18.760 ;
        RECT 197.720 18.440 198.040 18.760 ;
        RECT 198.120 18.440 198.440 18.760 ;
        RECT 198.520 18.440 198.840 18.760 ;
        RECT 198.920 18.440 199.240 18.760 ;
        RECT 199.320 18.440 199.640 18.760 ;
        RECT 199.720 18.440 200.040 18.760 ;
        RECT 200.120 18.440 200.440 18.760 ;
        RECT 200.520 18.440 200.840 18.760 ;
        RECT 200.920 18.440 201.240 18.760 ;
        RECT 201.320 18.440 201.640 18.760 ;
        RECT 201.720 18.440 202.040 18.760 ;
        RECT 202.120 18.440 202.440 18.760 ;
        RECT 202.520 18.440 202.840 18.760 ;
        RECT 202.920 18.440 203.240 18.760 ;
        RECT 203.320 18.440 203.640 18.760 ;
        RECT 203.720 18.440 204.040 18.760 ;
        RECT 204.120 18.440 204.440 18.760 ;
        RECT 204.520 18.440 204.840 18.760 ;
        RECT 204.920 18.440 205.240 18.760 ;
        RECT 205.320 18.440 205.640 18.760 ;
        RECT 0.040 18.040 0.360 18.360 ;
        RECT 0.440 18.040 0.760 18.360 ;
        RECT 0.840 18.040 1.160 18.360 ;
        RECT 1.240 18.040 1.560 18.360 ;
        RECT 1.640 18.040 1.960 18.360 ;
        RECT 2.040 18.040 2.360 18.360 ;
        RECT 2.440 18.040 2.760 18.360 ;
        RECT 2.840 18.040 3.160 18.360 ;
        RECT 3.240 18.040 3.560 18.360 ;
        RECT 3.640 18.040 3.960 18.360 ;
        RECT 4.040 18.040 4.360 18.360 ;
        RECT 4.440 18.040 4.760 18.360 ;
        RECT 4.840 18.040 5.160 18.360 ;
        RECT 5.240 18.040 5.560 18.360 ;
        RECT 5.640 18.040 5.960 18.360 ;
        RECT 6.040 18.040 6.360 18.360 ;
        RECT 6.440 18.040 6.760 18.360 ;
        RECT 6.840 18.040 7.160 18.360 ;
        RECT 7.240 18.040 7.560 18.360 ;
        RECT 7.640 18.040 7.960 18.360 ;
        RECT 8.040 18.040 8.360 18.360 ;
        RECT 8.440 18.040 8.760 18.360 ;
        RECT 8.840 18.040 9.160 18.360 ;
        RECT 9.240 18.040 9.560 18.360 ;
        RECT 9.640 18.040 9.960 18.360 ;
        RECT 10.040 18.040 10.360 18.360 ;
        RECT 10.440 18.040 10.760 18.360 ;
        RECT 10.840 18.040 11.160 18.360 ;
        RECT 11.240 18.040 11.560 18.360 ;
        RECT 11.640 18.040 11.960 18.360 ;
        RECT 12.040 18.040 12.360 18.360 ;
        RECT 12.440 18.040 12.760 18.360 ;
        RECT 12.840 18.040 13.160 18.360 ;
        RECT 13.240 18.040 13.560 18.360 ;
        RECT 13.640 18.040 13.960 18.360 ;
        RECT 14.040 18.040 14.360 18.360 ;
        RECT 14.440 18.040 14.760 18.360 ;
        RECT 14.840 18.040 15.160 18.360 ;
        RECT 15.240 18.040 15.560 18.360 ;
        RECT 15.640 18.040 15.960 18.360 ;
        RECT 16.040 18.040 16.360 18.360 ;
        RECT 16.440 18.040 16.760 18.360 ;
        RECT 16.840 18.040 17.160 18.360 ;
        RECT 17.240 18.040 17.560 18.360 ;
        RECT 17.640 18.040 17.960 18.360 ;
        RECT 18.040 18.040 18.360 18.360 ;
        RECT 18.440 18.040 18.760 18.360 ;
        RECT 18.840 18.040 19.160 18.360 ;
        RECT 19.240 18.040 19.560 18.360 ;
        RECT 19.640 18.040 19.960 18.360 ;
        RECT 95.560 18.040 95.880 18.360 ;
        RECT 95.960 18.040 96.280 18.360 ;
        RECT 96.360 18.040 96.680 18.360 ;
        RECT 96.760 18.040 97.080 18.360 ;
        RECT 145.560 18.040 145.880 18.360 ;
        RECT 145.960 18.040 146.280 18.360 ;
        RECT 146.360 18.040 146.680 18.360 ;
        RECT 146.760 18.040 147.080 18.360 ;
        RECT 185.720 18.040 186.040 18.360 ;
        RECT 186.120 18.040 186.440 18.360 ;
        RECT 186.520 18.040 186.840 18.360 ;
        RECT 186.920 18.040 187.240 18.360 ;
        RECT 187.320 18.040 187.640 18.360 ;
        RECT 187.720 18.040 188.040 18.360 ;
        RECT 188.120 18.040 188.440 18.360 ;
        RECT 188.520 18.040 188.840 18.360 ;
        RECT 188.920 18.040 189.240 18.360 ;
        RECT 189.320 18.040 189.640 18.360 ;
        RECT 189.720 18.040 190.040 18.360 ;
        RECT 190.120 18.040 190.440 18.360 ;
        RECT 190.520 18.040 190.840 18.360 ;
        RECT 190.920 18.040 191.240 18.360 ;
        RECT 191.320 18.040 191.640 18.360 ;
        RECT 191.720 18.040 192.040 18.360 ;
        RECT 192.120 18.040 192.440 18.360 ;
        RECT 192.520 18.040 192.840 18.360 ;
        RECT 192.920 18.040 193.240 18.360 ;
        RECT 193.320 18.040 193.640 18.360 ;
        RECT 193.720 18.040 194.040 18.360 ;
        RECT 194.120 18.040 194.440 18.360 ;
        RECT 194.520 18.040 194.840 18.360 ;
        RECT 194.920 18.040 195.240 18.360 ;
        RECT 195.320 18.040 195.640 18.360 ;
        RECT 195.720 18.040 196.040 18.360 ;
        RECT 196.120 18.040 196.440 18.360 ;
        RECT 196.520 18.040 196.840 18.360 ;
        RECT 196.920 18.040 197.240 18.360 ;
        RECT 197.320 18.040 197.640 18.360 ;
        RECT 197.720 18.040 198.040 18.360 ;
        RECT 198.120 18.040 198.440 18.360 ;
        RECT 198.520 18.040 198.840 18.360 ;
        RECT 198.920 18.040 199.240 18.360 ;
        RECT 199.320 18.040 199.640 18.360 ;
        RECT 199.720 18.040 200.040 18.360 ;
        RECT 200.120 18.040 200.440 18.360 ;
        RECT 200.520 18.040 200.840 18.360 ;
        RECT 200.920 18.040 201.240 18.360 ;
        RECT 201.320 18.040 201.640 18.360 ;
        RECT 201.720 18.040 202.040 18.360 ;
        RECT 202.120 18.040 202.440 18.360 ;
        RECT 202.520 18.040 202.840 18.360 ;
        RECT 202.920 18.040 203.240 18.360 ;
        RECT 203.320 18.040 203.640 18.360 ;
        RECT 203.720 18.040 204.040 18.360 ;
        RECT 204.120 18.040 204.440 18.360 ;
        RECT 204.520 18.040 204.840 18.360 ;
        RECT 204.920 18.040 205.240 18.360 ;
        RECT 205.320 18.040 205.640 18.360 ;
        RECT 0.040 17.640 0.360 17.960 ;
        RECT 0.440 17.640 0.760 17.960 ;
        RECT 0.840 17.640 1.160 17.960 ;
        RECT 1.240 17.640 1.560 17.960 ;
        RECT 1.640 17.640 1.960 17.960 ;
        RECT 2.040 17.640 2.360 17.960 ;
        RECT 2.440 17.640 2.760 17.960 ;
        RECT 2.840 17.640 3.160 17.960 ;
        RECT 3.240 17.640 3.560 17.960 ;
        RECT 3.640 17.640 3.960 17.960 ;
        RECT 4.040 17.640 4.360 17.960 ;
        RECT 4.440 17.640 4.760 17.960 ;
        RECT 4.840 17.640 5.160 17.960 ;
        RECT 5.240 17.640 5.560 17.960 ;
        RECT 5.640 17.640 5.960 17.960 ;
        RECT 6.040 17.640 6.360 17.960 ;
        RECT 6.440 17.640 6.760 17.960 ;
        RECT 6.840 17.640 7.160 17.960 ;
        RECT 7.240 17.640 7.560 17.960 ;
        RECT 7.640 17.640 7.960 17.960 ;
        RECT 8.040 17.640 8.360 17.960 ;
        RECT 8.440 17.640 8.760 17.960 ;
        RECT 8.840 17.640 9.160 17.960 ;
        RECT 9.240 17.640 9.560 17.960 ;
        RECT 9.640 17.640 9.960 17.960 ;
        RECT 10.040 17.640 10.360 17.960 ;
        RECT 10.440 17.640 10.760 17.960 ;
        RECT 10.840 17.640 11.160 17.960 ;
        RECT 11.240 17.640 11.560 17.960 ;
        RECT 11.640 17.640 11.960 17.960 ;
        RECT 12.040 17.640 12.360 17.960 ;
        RECT 12.440 17.640 12.760 17.960 ;
        RECT 12.840 17.640 13.160 17.960 ;
        RECT 13.240 17.640 13.560 17.960 ;
        RECT 13.640 17.640 13.960 17.960 ;
        RECT 14.040 17.640 14.360 17.960 ;
        RECT 14.440 17.640 14.760 17.960 ;
        RECT 14.840 17.640 15.160 17.960 ;
        RECT 15.240 17.640 15.560 17.960 ;
        RECT 15.640 17.640 15.960 17.960 ;
        RECT 16.040 17.640 16.360 17.960 ;
        RECT 16.440 17.640 16.760 17.960 ;
        RECT 16.840 17.640 17.160 17.960 ;
        RECT 17.240 17.640 17.560 17.960 ;
        RECT 17.640 17.640 17.960 17.960 ;
        RECT 18.040 17.640 18.360 17.960 ;
        RECT 18.440 17.640 18.760 17.960 ;
        RECT 18.840 17.640 19.160 17.960 ;
        RECT 19.240 17.640 19.560 17.960 ;
        RECT 19.640 17.640 19.960 17.960 ;
        RECT 95.560 17.640 95.880 17.960 ;
        RECT 95.960 17.640 96.280 17.960 ;
        RECT 96.360 17.640 96.680 17.960 ;
        RECT 96.760 17.640 97.080 17.960 ;
        RECT 145.560 17.640 145.880 17.960 ;
        RECT 145.960 17.640 146.280 17.960 ;
        RECT 146.360 17.640 146.680 17.960 ;
        RECT 146.760 17.640 147.080 17.960 ;
        RECT 185.720 17.640 186.040 17.960 ;
        RECT 186.120 17.640 186.440 17.960 ;
        RECT 186.520 17.640 186.840 17.960 ;
        RECT 186.920 17.640 187.240 17.960 ;
        RECT 187.320 17.640 187.640 17.960 ;
        RECT 187.720 17.640 188.040 17.960 ;
        RECT 188.120 17.640 188.440 17.960 ;
        RECT 188.520 17.640 188.840 17.960 ;
        RECT 188.920 17.640 189.240 17.960 ;
        RECT 189.320 17.640 189.640 17.960 ;
        RECT 189.720 17.640 190.040 17.960 ;
        RECT 190.120 17.640 190.440 17.960 ;
        RECT 190.520 17.640 190.840 17.960 ;
        RECT 190.920 17.640 191.240 17.960 ;
        RECT 191.320 17.640 191.640 17.960 ;
        RECT 191.720 17.640 192.040 17.960 ;
        RECT 192.120 17.640 192.440 17.960 ;
        RECT 192.520 17.640 192.840 17.960 ;
        RECT 192.920 17.640 193.240 17.960 ;
        RECT 193.320 17.640 193.640 17.960 ;
        RECT 193.720 17.640 194.040 17.960 ;
        RECT 194.120 17.640 194.440 17.960 ;
        RECT 194.520 17.640 194.840 17.960 ;
        RECT 194.920 17.640 195.240 17.960 ;
        RECT 195.320 17.640 195.640 17.960 ;
        RECT 195.720 17.640 196.040 17.960 ;
        RECT 196.120 17.640 196.440 17.960 ;
        RECT 196.520 17.640 196.840 17.960 ;
        RECT 196.920 17.640 197.240 17.960 ;
        RECT 197.320 17.640 197.640 17.960 ;
        RECT 197.720 17.640 198.040 17.960 ;
        RECT 198.120 17.640 198.440 17.960 ;
        RECT 198.520 17.640 198.840 17.960 ;
        RECT 198.920 17.640 199.240 17.960 ;
        RECT 199.320 17.640 199.640 17.960 ;
        RECT 199.720 17.640 200.040 17.960 ;
        RECT 200.120 17.640 200.440 17.960 ;
        RECT 200.520 17.640 200.840 17.960 ;
        RECT 200.920 17.640 201.240 17.960 ;
        RECT 201.320 17.640 201.640 17.960 ;
        RECT 201.720 17.640 202.040 17.960 ;
        RECT 202.120 17.640 202.440 17.960 ;
        RECT 202.520 17.640 202.840 17.960 ;
        RECT 202.920 17.640 203.240 17.960 ;
        RECT 203.320 17.640 203.640 17.960 ;
        RECT 203.720 17.640 204.040 17.960 ;
        RECT 204.120 17.640 204.440 17.960 ;
        RECT 204.520 17.640 204.840 17.960 ;
        RECT 204.920 17.640 205.240 17.960 ;
        RECT 205.320 17.640 205.640 17.960 ;
        RECT 0.040 17.240 0.360 17.560 ;
        RECT 0.440 17.240 0.760 17.560 ;
        RECT 0.840 17.240 1.160 17.560 ;
        RECT 1.240 17.240 1.560 17.560 ;
        RECT 1.640 17.240 1.960 17.560 ;
        RECT 2.040 17.240 2.360 17.560 ;
        RECT 2.440 17.240 2.760 17.560 ;
        RECT 2.840 17.240 3.160 17.560 ;
        RECT 3.240 17.240 3.560 17.560 ;
        RECT 3.640 17.240 3.960 17.560 ;
        RECT 4.040 17.240 4.360 17.560 ;
        RECT 4.440 17.240 4.760 17.560 ;
        RECT 4.840 17.240 5.160 17.560 ;
        RECT 5.240 17.240 5.560 17.560 ;
        RECT 5.640 17.240 5.960 17.560 ;
        RECT 6.040 17.240 6.360 17.560 ;
        RECT 6.440 17.240 6.760 17.560 ;
        RECT 6.840 17.240 7.160 17.560 ;
        RECT 7.240 17.240 7.560 17.560 ;
        RECT 7.640 17.240 7.960 17.560 ;
        RECT 8.040 17.240 8.360 17.560 ;
        RECT 8.440 17.240 8.760 17.560 ;
        RECT 8.840 17.240 9.160 17.560 ;
        RECT 9.240 17.240 9.560 17.560 ;
        RECT 9.640 17.240 9.960 17.560 ;
        RECT 10.040 17.240 10.360 17.560 ;
        RECT 10.440 17.240 10.760 17.560 ;
        RECT 10.840 17.240 11.160 17.560 ;
        RECT 11.240 17.240 11.560 17.560 ;
        RECT 11.640 17.240 11.960 17.560 ;
        RECT 12.040 17.240 12.360 17.560 ;
        RECT 12.440 17.240 12.760 17.560 ;
        RECT 12.840 17.240 13.160 17.560 ;
        RECT 13.240 17.240 13.560 17.560 ;
        RECT 13.640 17.240 13.960 17.560 ;
        RECT 14.040 17.240 14.360 17.560 ;
        RECT 14.440 17.240 14.760 17.560 ;
        RECT 14.840 17.240 15.160 17.560 ;
        RECT 15.240 17.240 15.560 17.560 ;
        RECT 15.640 17.240 15.960 17.560 ;
        RECT 16.040 17.240 16.360 17.560 ;
        RECT 16.440 17.240 16.760 17.560 ;
        RECT 16.840 17.240 17.160 17.560 ;
        RECT 17.240 17.240 17.560 17.560 ;
        RECT 17.640 17.240 17.960 17.560 ;
        RECT 18.040 17.240 18.360 17.560 ;
        RECT 18.440 17.240 18.760 17.560 ;
        RECT 18.840 17.240 19.160 17.560 ;
        RECT 19.240 17.240 19.560 17.560 ;
        RECT 19.640 17.240 19.960 17.560 ;
        RECT 95.560 17.240 95.880 17.560 ;
        RECT 95.960 17.240 96.280 17.560 ;
        RECT 96.360 17.240 96.680 17.560 ;
        RECT 96.760 17.240 97.080 17.560 ;
        RECT 145.560 17.240 145.880 17.560 ;
        RECT 145.960 17.240 146.280 17.560 ;
        RECT 146.360 17.240 146.680 17.560 ;
        RECT 146.760 17.240 147.080 17.560 ;
        RECT 185.720 17.240 186.040 17.560 ;
        RECT 186.120 17.240 186.440 17.560 ;
        RECT 186.520 17.240 186.840 17.560 ;
        RECT 186.920 17.240 187.240 17.560 ;
        RECT 187.320 17.240 187.640 17.560 ;
        RECT 187.720 17.240 188.040 17.560 ;
        RECT 188.120 17.240 188.440 17.560 ;
        RECT 188.520 17.240 188.840 17.560 ;
        RECT 188.920 17.240 189.240 17.560 ;
        RECT 189.320 17.240 189.640 17.560 ;
        RECT 189.720 17.240 190.040 17.560 ;
        RECT 190.120 17.240 190.440 17.560 ;
        RECT 190.520 17.240 190.840 17.560 ;
        RECT 190.920 17.240 191.240 17.560 ;
        RECT 191.320 17.240 191.640 17.560 ;
        RECT 191.720 17.240 192.040 17.560 ;
        RECT 192.120 17.240 192.440 17.560 ;
        RECT 192.520 17.240 192.840 17.560 ;
        RECT 192.920 17.240 193.240 17.560 ;
        RECT 193.320 17.240 193.640 17.560 ;
        RECT 193.720 17.240 194.040 17.560 ;
        RECT 194.120 17.240 194.440 17.560 ;
        RECT 194.520 17.240 194.840 17.560 ;
        RECT 194.920 17.240 195.240 17.560 ;
        RECT 195.320 17.240 195.640 17.560 ;
        RECT 195.720 17.240 196.040 17.560 ;
        RECT 196.120 17.240 196.440 17.560 ;
        RECT 196.520 17.240 196.840 17.560 ;
        RECT 196.920 17.240 197.240 17.560 ;
        RECT 197.320 17.240 197.640 17.560 ;
        RECT 197.720 17.240 198.040 17.560 ;
        RECT 198.120 17.240 198.440 17.560 ;
        RECT 198.520 17.240 198.840 17.560 ;
        RECT 198.920 17.240 199.240 17.560 ;
        RECT 199.320 17.240 199.640 17.560 ;
        RECT 199.720 17.240 200.040 17.560 ;
        RECT 200.120 17.240 200.440 17.560 ;
        RECT 200.520 17.240 200.840 17.560 ;
        RECT 200.920 17.240 201.240 17.560 ;
        RECT 201.320 17.240 201.640 17.560 ;
        RECT 201.720 17.240 202.040 17.560 ;
        RECT 202.120 17.240 202.440 17.560 ;
        RECT 202.520 17.240 202.840 17.560 ;
        RECT 202.920 17.240 203.240 17.560 ;
        RECT 203.320 17.240 203.640 17.560 ;
        RECT 203.720 17.240 204.040 17.560 ;
        RECT 204.120 17.240 204.440 17.560 ;
        RECT 204.520 17.240 204.840 17.560 ;
        RECT 204.920 17.240 205.240 17.560 ;
        RECT 205.320 17.240 205.640 17.560 ;
        RECT 0.040 16.840 0.360 17.160 ;
        RECT 0.440 16.840 0.760 17.160 ;
        RECT 0.840 16.840 1.160 17.160 ;
        RECT 1.240 16.840 1.560 17.160 ;
        RECT 1.640 16.840 1.960 17.160 ;
        RECT 2.040 16.840 2.360 17.160 ;
        RECT 2.440 16.840 2.760 17.160 ;
        RECT 2.840 16.840 3.160 17.160 ;
        RECT 3.240 16.840 3.560 17.160 ;
        RECT 3.640 16.840 3.960 17.160 ;
        RECT 4.040 16.840 4.360 17.160 ;
        RECT 4.440 16.840 4.760 17.160 ;
        RECT 4.840 16.840 5.160 17.160 ;
        RECT 5.240 16.840 5.560 17.160 ;
        RECT 5.640 16.840 5.960 17.160 ;
        RECT 6.040 16.840 6.360 17.160 ;
        RECT 6.440 16.840 6.760 17.160 ;
        RECT 6.840 16.840 7.160 17.160 ;
        RECT 7.240 16.840 7.560 17.160 ;
        RECT 7.640 16.840 7.960 17.160 ;
        RECT 8.040 16.840 8.360 17.160 ;
        RECT 8.440 16.840 8.760 17.160 ;
        RECT 8.840 16.840 9.160 17.160 ;
        RECT 9.240 16.840 9.560 17.160 ;
        RECT 9.640 16.840 9.960 17.160 ;
        RECT 10.040 16.840 10.360 17.160 ;
        RECT 10.440 16.840 10.760 17.160 ;
        RECT 10.840 16.840 11.160 17.160 ;
        RECT 11.240 16.840 11.560 17.160 ;
        RECT 11.640 16.840 11.960 17.160 ;
        RECT 12.040 16.840 12.360 17.160 ;
        RECT 12.440 16.840 12.760 17.160 ;
        RECT 12.840 16.840 13.160 17.160 ;
        RECT 13.240 16.840 13.560 17.160 ;
        RECT 13.640 16.840 13.960 17.160 ;
        RECT 14.040 16.840 14.360 17.160 ;
        RECT 14.440 16.840 14.760 17.160 ;
        RECT 14.840 16.840 15.160 17.160 ;
        RECT 15.240 16.840 15.560 17.160 ;
        RECT 15.640 16.840 15.960 17.160 ;
        RECT 16.040 16.840 16.360 17.160 ;
        RECT 16.440 16.840 16.760 17.160 ;
        RECT 16.840 16.840 17.160 17.160 ;
        RECT 17.240 16.840 17.560 17.160 ;
        RECT 17.640 16.840 17.960 17.160 ;
        RECT 18.040 16.840 18.360 17.160 ;
        RECT 18.440 16.840 18.760 17.160 ;
        RECT 18.840 16.840 19.160 17.160 ;
        RECT 19.240 16.840 19.560 17.160 ;
        RECT 19.640 16.840 19.960 17.160 ;
        RECT 95.560 16.840 95.880 17.160 ;
        RECT 95.960 16.840 96.280 17.160 ;
        RECT 96.360 16.840 96.680 17.160 ;
        RECT 96.760 16.840 97.080 17.160 ;
        RECT 145.560 16.840 145.880 17.160 ;
        RECT 145.960 16.840 146.280 17.160 ;
        RECT 146.360 16.840 146.680 17.160 ;
        RECT 146.760 16.840 147.080 17.160 ;
        RECT 185.720 16.840 186.040 17.160 ;
        RECT 186.120 16.840 186.440 17.160 ;
        RECT 186.520 16.840 186.840 17.160 ;
        RECT 186.920 16.840 187.240 17.160 ;
        RECT 187.320 16.840 187.640 17.160 ;
        RECT 187.720 16.840 188.040 17.160 ;
        RECT 188.120 16.840 188.440 17.160 ;
        RECT 188.520 16.840 188.840 17.160 ;
        RECT 188.920 16.840 189.240 17.160 ;
        RECT 189.320 16.840 189.640 17.160 ;
        RECT 189.720 16.840 190.040 17.160 ;
        RECT 190.120 16.840 190.440 17.160 ;
        RECT 190.520 16.840 190.840 17.160 ;
        RECT 190.920 16.840 191.240 17.160 ;
        RECT 191.320 16.840 191.640 17.160 ;
        RECT 191.720 16.840 192.040 17.160 ;
        RECT 192.120 16.840 192.440 17.160 ;
        RECT 192.520 16.840 192.840 17.160 ;
        RECT 192.920 16.840 193.240 17.160 ;
        RECT 193.320 16.840 193.640 17.160 ;
        RECT 193.720 16.840 194.040 17.160 ;
        RECT 194.120 16.840 194.440 17.160 ;
        RECT 194.520 16.840 194.840 17.160 ;
        RECT 194.920 16.840 195.240 17.160 ;
        RECT 195.320 16.840 195.640 17.160 ;
        RECT 195.720 16.840 196.040 17.160 ;
        RECT 196.120 16.840 196.440 17.160 ;
        RECT 196.520 16.840 196.840 17.160 ;
        RECT 196.920 16.840 197.240 17.160 ;
        RECT 197.320 16.840 197.640 17.160 ;
        RECT 197.720 16.840 198.040 17.160 ;
        RECT 198.120 16.840 198.440 17.160 ;
        RECT 198.520 16.840 198.840 17.160 ;
        RECT 198.920 16.840 199.240 17.160 ;
        RECT 199.320 16.840 199.640 17.160 ;
        RECT 199.720 16.840 200.040 17.160 ;
        RECT 200.120 16.840 200.440 17.160 ;
        RECT 200.520 16.840 200.840 17.160 ;
        RECT 200.920 16.840 201.240 17.160 ;
        RECT 201.320 16.840 201.640 17.160 ;
        RECT 201.720 16.840 202.040 17.160 ;
        RECT 202.120 16.840 202.440 17.160 ;
        RECT 202.520 16.840 202.840 17.160 ;
        RECT 202.920 16.840 203.240 17.160 ;
        RECT 203.320 16.840 203.640 17.160 ;
        RECT 203.720 16.840 204.040 17.160 ;
        RECT 204.120 16.840 204.440 17.160 ;
        RECT 204.520 16.840 204.840 17.160 ;
        RECT 204.920 16.840 205.240 17.160 ;
        RECT 205.320 16.840 205.640 17.160 ;
        RECT 0.040 16.440 0.360 16.760 ;
        RECT 0.440 16.440 0.760 16.760 ;
        RECT 0.840 16.440 1.160 16.760 ;
        RECT 1.240 16.440 1.560 16.760 ;
        RECT 1.640 16.440 1.960 16.760 ;
        RECT 2.040 16.440 2.360 16.760 ;
        RECT 2.440 16.440 2.760 16.760 ;
        RECT 2.840 16.440 3.160 16.760 ;
        RECT 3.240 16.440 3.560 16.760 ;
        RECT 3.640 16.440 3.960 16.760 ;
        RECT 4.040 16.440 4.360 16.760 ;
        RECT 4.440 16.440 4.760 16.760 ;
        RECT 4.840 16.440 5.160 16.760 ;
        RECT 5.240 16.440 5.560 16.760 ;
        RECT 5.640 16.440 5.960 16.760 ;
        RECT 6.040 16.440 6.360 16.760 ;
        RECT 6.440 16.440 6.760 16.760 ;
        RECT 6.840 16.440 7.160 16.760 ;
        RECT 7.240 16.440 7.560 16.760 ;
        RECT 7.640 16.440 7.960 16.760 ;
        RECT 8.040 16.440 8.360 16.760 ;
        RECT 8.440 16.440 8.760 16.760 ;
        RECT 8.840 16.440 9.160 16.760 ;
        RECT 9.240 16.440 9.560 16.760 ;
        RECT 9.640 16.440 9.960 16.760 ;
        RECT 10.040 16.440 10.360 16.760 ;
        RECT 10.440 16.440 10.760 16.760 ;
        RECT 10.840 16.440 11.160 16.760 ;
        RECT 11.240 16.440 11.560 16.760 ;
        RECT 11.640 16.440 11.960 16.760 ;
        RECT 12.040 16.440 12.360 16.760 ;
        RECT 12.440 16.440 12.760 16.760 ;
        RECT 12.840 16.440 13.160 16.760 ;
        RECT 13.240 16.440 13.560 16.760 ;
        RECT 13.640 16.440 13.960 16.760 ;
        RECT 14.040 16.440 14.360 16.760 ;
        RECT 14.440 16.440 14.760 16.760 ;
        RECT 14.840 16.440 15.160 16.760 ;
        RECT 15.240 16.440 15.560 16.760 ;
        RECT 15.640 16.440 15.960 16.760 ;
        RECT 16.040 16.440 16.360 16.760 ;
        RECT 16.440 16.440 16.760 16.760 ;
        RECT 16.840 16.440 17.160 16.760 ;
        RECT 17.240 16.440 17.560 16.760 ;
        RECT 17.640 16.440 17.960 16.760 ;
        RECT 18.040 16.440 18.360 16.760 ;
        RECT 18.440 16.440 18.760 16.760 ;
        RECT 18.840 16.440 19.160 16.760 ;
        RECT 19.240 16.440 19.560 16.760 ;
        RECT 19.640 16.440 19.960 16.760 ;
        RECT 95.560 16.440 95.880 16.760 ;
        RECT 95.960 16.440 96.280 16.760 ;
        RECT 96.360 16.440 96.680 16.760 ;
        RECT 96.760 16.440 97.080 16.760 ;
        RECT 145.560 16.440 145.880 16.760 ;
        RECT 145.960 16.440 146.280 16.760 ;
        RECT 146.360 16.440 146.680 16.760 ;
        RECT 146.760 16.440 147.080 16.760 ;
        RECT 185.720 16.440 186.040 16.760 ;
        RECT 186.120 16.440 186.440 16.760 ;
        RECT 186.520 16.440 186.840 16.760 ;
        RECT 186.920 16.440 187.240 16.760 ;
        RECT 187.320 16.440 187.640 16.760 ;
        RECT 187.720 16.440 188.040 16.760 ;
        RECT 188.120 16.440 188.440 16.760 ;
        RECT 188.520 16.440 188.840 16.760 ;
        RECT 188.920 16.440 189.240 16.760 ;
        RECT 189.320 16.440 189.640 16.760 ;
        RECT 189.720 16.440 190.040 16.760 ;
        RECT 190.120 16.440 190.440 16.760 ;
        RECT 190.520 16.440 190.840 16.760 ;
        RECT 190.920 16.440 191.240 16.760 ;
        RECT 191.320 16.440 191.640 16.760 ;
        RECT 191.720 16.440 192.040 16.760 ;
        RECT 192.120 16.440 192.440 16.760 ;
        RECT 192.520 16.440 192.840 16.760 ;
        RECT 192.920 16.440 193.240 16.760 ;
        RECT 193.320 16.440 193.640 16.760 ;
        RECT 193.720 16.440 194.040 16.760 ;
        RECT 194.120 16.440 194.440 16.760 ;
        RECT 194.520 16.440 194.840 16.760 ;
        RECT 194.920 16.440 195.240 16.760 ;
        RECT 195.320 16.440 195.640 16.760 ;
        RECT 195.720 16.440 196.040 16.760 ;
        RECT 196.120 16.440 196.440 16.760 ;
        RECT 196.520 16.440 196.840 16.760 ;
        RECT 196.920 16.440 197.240 16.760 ;
        RECT 197.320 16.440 197.640 16.760 ;
        RECT 197.720 16.440 198.040 16.760 ;
        RECT 198.120 16.440 198.440 16.760 ;
        RECT 198.520 16.440 198.840 16.760 ;
        RECT 198.920 16.440 199.240 16.760 ;
        RECT 199.320 16.440 199.640 16.760 ;
        RECT 199.720 16.440 200.040 16.760 ;
        RECT 200.120 16.440 200.440 16.760 ;
        RECT 200.520 16.440 200.840 16.760 ;
        RECT 200.920 16.440 201.240 16.760 ;
        RECT 201.320 16.440 201.640 16.760 ;
        RECT 201.720 16.440 202.040 16.760 ;
        RECT 202.120 16.440 202.440 16.760 ;
        RECT 202.520 16.440 202.840 16.760 ;
        RECT 202.920 16.440 203.240 16.760 ;
        RECT 203.320 16.440 203.640 16.760 ;
        RECT 203.720 16.440 204.040 16.760 ;
        RECT 204.120 16.440 204.440 16.760 ;
        RECT 204.520 16.440 204.840 16.760 ;
        RECT 204.920 16.440 205.240 16.760 ;
        RECT 205.320 16.440 205.640 16.760 ;
        RECT 0.040 16.040 0.360 16.360 ;
        RECT 0.440 16.040 0.760 16.360 ;
        RECT 0.840 16.040 1.160 16.360 ;
        RECT 1.240 16.040 1.560 16.360 ;
        RECT 1.640 16.040 1.960 16.360 ;
        RECT 2.040 16.040 2.360 16.360 ;
        RECT 2.440 16.040 2.760 16.360 ;
        RECT 2.840 16.040 3.160 16.360 ;
        RECT 3.240 16.040 3.560 16.360 ;
        RECT 3.640 16.040 3.960 16.360 ;
        RECT 4.040 16.040 4.360 16.360 ;
        RECT 4.440 16.040 4.760 16.360 ;
        RECT 4.840 16.040 5.160 16.360 ;
        RECT 5.240 16.040 5.560 16.360 ;
        RECT 5.640 16.040 5.960 16.360 ;
        RECT 6.040 16.040 6.360 16.360 ;
        RECT 6.440 16.040 6.760 16.360 ;
        RECT 6.840 16.040 7.160 16.360 ;
        RECT 7.240 16.040 7.560 16.360 ;
        RECT 7.640 16.040 7.960 16.360 ;
        RECT 8.040 16.040 8.360 16.360 ;
        RECT 8.440 16.040 8.760 16.360 ;
        RECT 8.840 16.040 9.160 16.360 ;
        RECT 9.240 16.040 9.560 16.360 ;
        RECT 9.640 16.040 9.960 16.360 ;
        RECT 10.040 16.040 10.360 16.360 ;
        RECT 10.440 16.040 10.760 16.360 ;
        RECT 10.840 16.040 11.160 16.360 ;
        RECT 11.240 16.040 11.560 16.360 ;
        RECT 11.640 16.040 11.960 16.360 ;
        RECT 12.040 16.040 12.360 16.360 ;
        RECT 12.440 16.040 12.760 16.360 ;
        RECT 12.840 16.040 13.160 16.360 ;
        RECT 13.240 16.040 13.560 16.360 ;
        RECT 13.640 16.040 13.960 16.360 ;
        RECT 14.040 16.040 14.360 16.360 ;
        RECT 14.440 16.040 14.760 16.360 ;
        RECT 14.840 16.040 15.160 16.360 ;
        RECT 15.240 16.040 15.560 16.360 ;
        RECT 15.640 16.040 15.960 16.360 ;
        RECT 16.040 16.040 16.360 16.360 ;
        RECT 16.440 16.040 16.760 16.360 ;
        RECT 16.840 16.040 17.160 16.360 ;
        RECT 17.240 16.040 17.560 16.360 ;
        RECT 17.640 16.040 17.960 16.360 ;
        RECT 18.040 16.040 18.360 16.360 ;
        RECT 18.440 16.040 18.760 16.360 ;
        RECT 18.840 16.040 19.160 16.360 ;
        RECT 19.240 16.040 19.560 16.360 ;
        RECT 19.640 16.040 19.960 16.360 ;
        RECT 95.560 16.040 95.880 16.360 ;
        RECT 95.960 16.040 96.280 16.360 ;
        RECT 96.360 16.040 96.680 16.360 ;
        RECT 96.760 16.040 97.080 16.360 ;
        RECT 145.560 16.040 145.880 16.360 ;
        RECT 145.960 16.040 146.280 16.360 ;
        RECT 146.360 16.040 146.680 16.360 ;
        RECT 146.760 16.040 147.080 16.360 ;
        RECT 185.720 16.040 186.040 16.360 ;
        RECT 186.120 16.040 186.440 16.360 ;
        RECT 186.520 16.040 186.840 16.360 ;
        RECT 186.920 16.040 187.240 16.360 ;
        RECT 187.320 16.040 187.640 16.360 ;
        RECT 187.720 16.040 188.040 16.360 ;
        RECT 188.120 16.040 188.440 16.360 ;
        RECT 188.520 16.040 188.840 16.360 ;
        RECT 188.920 16.040 189.240 16.360 ;
        RECT 189.320 16.040 189.640 16.360 ;
        RECT 189.720 16.040 190.040 16.360 ;
        RECT 190.120 16.040 190.440 16.360 ;
        RECT 190.520 16.040 190.840 16.360 ;
        RECT 190.920 16.040 191.240 16.360 ;
        RECT 191.320 16.040 191.640 16.360 ;
        RECT 191.720 16.040 192.040 16.360 ;
        RECT 192.120 16.040 192.440 16.360 ;
        RECT 192.520 16.040 192.840 16.360 ;
        RECT 192.920 16.040 193.240 16.360 ;
        RECT 193.320 16.040 193.640 16.360 ;
        RECT 193.720 16.040 194.040 16.360 ;
        RECT 194.120 16.040 194.440 16.360 ;
        RECT 194.520 16.040 194.840 16.360 ;
        RECT 194.920 16.040 195.240 16.360 ;
        RECT 195.320 16.040 195.640 16.360 ;
        RECT 195.720 16.040 196.040 16.360 ;
        RECT 196.120 16.040 196.440 16.360 ;
        RECT 196.520 16.040 196.840 16.360 ;
        RECT 196.920 16.040 197.240 16.360 ;
        RECT 197.320 16.040 197.640 16.360 ;
        RECT 197.720 16.040 198.040 16.360 ;
        RECT 198.120 16.040 198.440 16.360 ;
        RECT 198.520 16.040 198.840 16.360 ;
        RECT 198.920 16.040 199.240 16.360 ;
        RECT 199.320 16.040 199.640 16.360 ;
        RECT 199.720 16.040 200.040 16.360 ;
        RECT 200.120 16.040 200.440 16.360 ;
        RECT 200.520 16.040 200.840 16.360 ;
        RECT 200.920 16.040 201.240 16.360 ;
        RECT 201.320 16.040 201.640 16.360 ;
        RECT 201.720 16.040 202.040 16.360 ;
        RECT 202.120 16.040 202.440 16.360 ;
        RECT 202.520 16.040 202.840 16.360 ;
        RECT 202.920 16.040 203.240 16.360 ;
        RECT 203.320 16.040 203.640 16.360 ;
        RECT 203.720 16.040 204.040 16.360 ;
        RECT 204.120 16.040 204.440 16.360 ;
        RECT 204.520 16.040 204.840 16.360 ;
        RECT 204.920 16.040 205.240 16.360 ;
        RECT 205.320 16.040 205.640 16.360 ;
        RECT 0.040 15.640 0.360 15.960 ;
        RECT 0.440 15.640 0.760 15.960 ;
        RECT 0.840 15.640 1.160 15.960 ;
        RECT 1.240 15.640 1.560 15.960 ;
        RECT 1.640 15.640 1.960 15.960 ;
        RECT 2.040 15.640 2.360 15.960 ;
        RECT 2.440 15.640 2.760 15.960 ;
        RECT 2.840 15.640 3.160 15.960 ;
        RECT 3.240 15.640 3.560 15.960 ;
        RECT 3.640 15.640 3.960 15.960 ;
        RECT 4.040 15.640 4.360 15.960 ;
        RECT 4.440 15.640 4.760 15.960 ;
        RECT 4.840 15.640 5.160 15.960 ;
        RECT 5.240 15.640 5.560 15.960 ;
        RECT 5.640 15.640 5.960 15.960 ;
        RECT 6.040 15.640 6.360 15.960 ;
        RECT 6.440 15.640 6.760 15.960 ;
        RECT 6.840 15.640 7.160 15.960 ;
        RECT 7.240 15.640 7.560 15.960 ;
        RECT 7.640 15.640 7.960 15.960 ;
        RECT 8.040 15.640 8.360 15.960 ;
        RECT 8.440 15.640 8.760 15.960 ;
        RECT 8.840 15.640 9.160 15.960 ;
        RECT 9.240 15.640 9.560 15.960 ;
        RECT 9.640 15.640 9.960 15.960 ;
        RECT 10.040 15.640 10.360 15.960 ;
        RECT 10.440 15.640 10.760 15.960 ;
        RECT 10.840 15.640 11.160 15.960 ;
        RECT 11.240 15.640 11.560 15.960 ;
        RECT 11.640 15.640 11.960 15.960 ;
        RECT 12.040 15.640 12.360 15.960 ;
        RECT 12.440 15.640 12.760 15.960 ;
        RECT 12.840 15.640 13.160 15.960 ;
        RECT 13.240 15.640 13.560 15.960 ;
        RECT 13.640 15.640 13.960 15.960 ;
        RECT 14.040 15.640 14.360 15.960 ;
        RECT 14.440 15.640 14.760 15.960 ;
        RECT 14.840 15.640 15.160 15.960 ;
        RECT 15.240 15.640 15.560 15.960 ;
        RECT 15.640 15.640 15.960 15.960 ;
        RECT 16.040 15.640 16.360 15.960 ;
        RECT 16.440 15.640 16.760 15.960 ;
        RECT 16.840 15.640 17.160 15.960 ;
        RECT 17.240 15.640 17.560 15.960 ;
        RECT 17.640 15.640 17.960 15.960 ;
        RECT 18.040 15.640 18.360 15.960 ;
        RECT 18.440 15.640 18.760 15.960 ;
        RECT 18.840 15.640 19.160 15.960 ;
        RECT 19.240 15.640 19.560 15.960 ;
        RECT 19.640 15.640 19.960 15.960 ;
        RECT 95.560 15.640 95.880 15.960 ;
        RECT 95.960 15.640 96.280 15.960 ;
        RECT 96.360 15.640 96.680 15.960 ;
        RECT 96.760 15.640 97.080 15.960 ;
        RECT 145.560 15.640 145.880 15.960 ;
        RECT 145.960 15.640 146.280 15.960 ;
        RECT 146.360 15.640 146.680 15.960 ;
        RECT 146.760 15.640 147.080 15.960 ;
        RECT 185.720 15.640 186.040 15.960 ;
        RECT 186.120 15.640 186.440 15.960 ;
        RECT 186.520 15.640 186.840 15.960 ;
        RECT 186.920 15.640 187.240 15.960 ;
        RECT 187.320 15.640 187.640 15.960 ;
        RECT 187.720 15.640 188.040 15.960 ;
        RECT 188.120 15.640 188.440 15.960 ;
        RECT 188.520 15.640 188.840 15.960 ;
        RECT 188.920 15.640 189.240 15.960 ;
        RECT 189.320 15.640 189.640 15.960 ;
        RECT 189.720 15.640 190.040 15.960 ;
        RECT 190.120 15.640 190.440 15.960 ;
        RECT 190.520 15.640 190.840 15.960 ;
        RECT 190.920 15.640 191.240 15.960 ;
        RECT 191.320 15.640 191.640 15.960 ;
        RECT 191.720 15.640 192.040 15.960 ;
        RECT 192.120 15.640 192.440 15.960 ;
        RECT 192.520 15.640 192.840 15.960 ;
        RECT 192.920 15.640 193.240 15.960 ;
        RECT 193.320 15.640 193.640 15.960 ;
        RECT 193.720 15.640 194.040 15.960 ;
        RECT 194.120 15.640 194.440 15.960 ;
        RECT 194.520 15.640 194.840 15.960 ;
        RECT 194.920 15.640 195.240 15.960 ;
        RECT 195.320 15.640 195.640 15.960 ;
        RECT 195.720 15.640 196.040 15.960 ;
        RECT 196.120 15.640 196.440 15.960 ;
        RECT 196.520 15.640 196.840 15.960 ;
        RECT 196.920 15.640 197.240 15.960 ;
        RECT 197.320 15.640 197.640 15.960 ;
        RECT 197.720 15.640 198.040 15.960 ;
        RECT 198.120 15.640 198.440 15.960 ;
        RECT 198.520 15.640 198.840 15.960 ;
        RECT 198.920 15.640 199.240 15.960 ;
        RECT 199.320 15.640 199.640 15.960 ;
        RECT 199.720 15.640 200.040 15.960 ;
        RECT 200.120 15.640 200.440 15.960 ;
        RECT 200.520 15.640 200.840 15.960 ;
        RECT 200.920 15.640 201.240 15.960 ;
        RECT 201.320 15.640 201.640 15.960 ;
        RECT 201.720 15.640 202.040 15.960 ;
        RECT 202.120 15.640 202.440 15.960 ;
        RECT 202.520 15.640 202.840 15.960 ;
        RECT 202.920 15.640 203.240 15.960 ;
        RECT 203.320 15.640 203.640 15.960 ;
        RECT 203.720 15.640 204.040 15.960 ;
        RECT 204.120 15.640 204.440 15.960 ;
        RECT 204.520 15.640 204.840 15.960 ;
        RECT 204.920 15.640 205.240 15.960 ;
        RECT 205.320 15.640 205.640 15.960 ;
        RECT 0.040 15.240 0.360 15.560 ;
        RECT 0.440 15.240 0.760 15.560 ;
        RECT 0.840 15.240 1.160 15.560 ;
        RECT 1.240 15.240 1.560 15.560 ;
        RECT 1.640 15.240 1.960 15.560 ;
        RECT 2.040 15.240 2.360 15.560 ;
        RECT 2.440 15.240 2.760 15.560 ;
        RECT 2.840 15.240 3.160 15.560 ;
        RECT 3.240 15.240 3.560 15.560 ;
        RECT 3.640 15.240 3.960 15.560 ;
        RECT 4.040 15.240 4.360 15.560 ;
        RECT 4.440 15.240 4.760 15.560 ;
        RECT 4.840 15.240 5.160 15.560 ;
        RECT 5.240 15.240 5.560 15.560 ;
        RECT 5.640 15.240 5.960 15.560 ;
        RECT 6.040 15.240 6.360 15.560 ;
        RECT 6.440 15.240 6.760 15.560 ;
        RECT 6.840 15.240 7.160 15.560 ;
        RECT 7.240 15.240 7.560 15.560 ;
        RECT 7.640 15.240 7.960 15.560 ;
        RECT 8.040 15.240 8.360 15.560 ;
        RECT 8.440 15.240 8.760 15.560 ;
        RECT 8.840 15.240 9.160 15.560 ;
        RECT 9.240 15.240 9.560 15.560 ;
        RECT 9.640 15.240 9.960 15.560 ;
        RECT 10.040 15.240 10.360 15.560 ;
        RECT 10.440 15.240 10.760 15.560 ;
        RECT 10.840 15.240 11.160 15.560 ;
        RECT 11.240 15.240 11.560 15.560 ;
        RECT 11.640 15.240 11.960 15.560 ;
        RECT 12.040 15.240 12.360 15.560 ;
        RECT 12.440 15.240 12.760 15.560 ;
        RECT 12.840 15.240 13.160 15.560 ;
        RECT 13.240 15.240 13.560 15.560 ;
        RECT 13.640 15.240 13.960 15.560 ;
        RECT 14.040 15.240 14.360 15.560 ;
        RECT 14.440 15.240 14.760 15.560 ;
        RECT 14.840 15.240 15.160 15.560 ;
        RECT 15.240 15.240 15.560 15.560 ;
        RECT 15.640 15.240 15.960 15.560 ;
        RECT 16.040 15.240 16.360 15.560 ;
        RECT 16.440 15.240 16.760 15.560 ;
        RECT 16.840 15.240 17.160 15.560 ;
        RECT 17.240 15.240 17.560 15.560 ;
        RECT 17.640 15.240 17.960 15.560 ;
        RECT 18.040 15.240 18.360 15.560 ;
        RECT 18.440 15.240 18.760 15.560 ;
        RECT 18.840 15.240 19.160 15.560 ;
        RECT 19.240 15.240 19.560 15.560 ;
        RECT 19.640 15.240 19.960 15.560 ;
        RECT 95.560 15.240 95.880 15.560 ;
        RECT 95.960 15.240 96.280 15.560 ;
        RECT 96.360 15.240 96.680 15.560 ;
        RECT 96.760 15.240 97.080 15.560 ;
        RECT 145.560 15.240 145.880 15.560 ;
        RECT 145.960 15.240 146.280 15.560 ;
        RECT 146.360 15.240 146.680 15.560 ;
        RECT 146.760 15.240 147.080 15.560 ;
        RECT 185.720 15.240 186.040 15.560 ;
        RECT 186.120 15.240 186.440 15.560 ;
        RECT 186.520 15.240 186.840 15.560 ;
        RECT 186.920 15.240 187.240 15.560 ;
        RECT 187.320 15.240 187.640 15.560 ;
        RECT 187.720 15.240 188.040 15.560 ;
        RECT 188.120 15.240 188.440 15.560 ;
        RECT 188.520 15.240 188.840 15.560 ;
        RECT 188.920 15.240 189.240 15.560 ;
        RECT 189.320 15.240 189.640 15.560 ;
        RECT 189.720 15.240 190.040 15.560 ;
        RECT 190.120 15.240 190.440 15.560 ;
        RECT 190.520 15.240 190.840 15.560 ;
        RECT 190.920 15.240 191.240 15.560 ;
        RECT 191.320 15.240 191.640 15.560 ;
        RECT 191.720 15.240 192.040 15.560 ;
        RECT 192.120 15.240 192.440 15.560 ;
        RECT 192.520 15.240 192.840 15.560 ;
        RECT 192.920 15.240 193.240 15.560 ;
        RECT 193.320 15.240 193.640 15.560 ;
        RECT 193.720 15.240 194.040 15.560 ;
        RECT 194.120 15.240 194.440 15.560 ;
        RECT 194.520 15.240 194.840 15.560 ;
        RECT 194.920 15.240 195.240 15.560 ;
        RECT 195.320 15.240 195.640 15.560 ;
        RECT 195.720 15.240 196.040 15.560 ;
        RECT 196.120 15.240 196.440 15.560 ;
        RECT 196.520 15.240 196.840 15.560 ;
        RECT 196.920 15.240 197.240 15.560 ;
        RECT 197.320 15.240 197.640 15.560 ;
        RECT 197.720 15.240 198.040 15.560 ;
        RECT 198.120 15.240 198.440 15.560 ;
        RECT 198.520 15.240 198.840 15.560 ;
        RECT 198.920 15.240 199.240 15.560 ;
        RECT 199.320 15.240 199.640 15.560 ;
        RECT 199.720 15.240 200.040 15.560 ;
        RECT 200.120 15.240 200.440 15.560 ;
        RECT 200.520 15.240 200.840 15.560 ;
        RECT 200.920 15.240 201.240 15.560 ;
        RECT 201.320 15.240 201.640 15.560 ;
        RECT 201.720 15.240 202.040 15.560 ;
        RECT 202.120 15.240 202.440 15.560 ;
        RECT 202.520 15.240 202.840 15.560 ;
        RECT 202.920 15.240 203.240 15.560 ;
        RECT 203.320 15.240 203.640 15.560 ;
        RECT 203.720 15.240 204.040 15.560 ;
        RECT 204.120 15.240 204.440 15.560 ;
        RECT 204.520 15.240 204.840 15.560 ;
        RECT 204.920 15.240 205.240 15.560 ;
        RECT 205.320 15.240 205.640 15.560 ;
        RECT 0.040 14.840 0.360 15.160 ;
        RECT 0.440 14.840 0.760 15.160 ;
        RECT 0.840 14.840 1.160 15.160 ;
        RECT 1.240 14.840 1.560 15.160 ;
        RECT 1.640 14.840 1.960 15.160 ;
        RECT 2.040 14.840 2.360 15.160 ;
        RECT 2.440 14.840 2.760 15.160 ;
        RECT 2.840 14.840 3.160 15.160 ;
        RECT 3.240 14.840 3.560 15.160 ;
        RECT 3.640 14.840 3.960 15.160 ;
        RECT 4.040 14.840 4.360 15.160 ;
        RECT 4.440 14.840 4.760 15.160 ;
        RECT 4.840 14.840 5.160 15.160 ;
        RECT 5.240 14.840 5.560 15.160 ;
        RECT 5.640 14.840 5.960 15.160 ;
        RECT 6.040 14.840 6.360 15.160 ;
        RECT 6.440 14.840 6.760 15.160 ;
        RECT 6.840 14.840 7.160 15.160 ;
        RECT 7.240 14.840 7.560 15.160 ;
        RECT 7.640 14.840 7.960 15.160 ;
        RECT 8.040 14.840 8.360 15.160 ;
        RECT 8.440 14.840 8.760 15.160 ;
        RECT 8.840 14.840 9.160 15.160 ;
        RECT 9.240 14.840 9.560 15.160 ;
        RECT 9.640 14.840 9.960 15.160 ;
        RECT 10.040 14.840 10.360 15.160 ;
        RECT 10.440 14.840 10.760 15.160 ;
        RECT 10.840 14.840 11.160 15.160 ;
        RECT 11.240 14.840 11.560 15.160 ;
        RECT 11.640 14.840 11.960 15.160 ;
        RECT 12.040 14.840 12.360 15.160 ;
        RECT 12.440 14.840 12.760 15.160 ;
        RECT 12.840 14.840 13.160 15.160 ;
        RECT 13.240 14.840 13.560 15.160 ;
        RECT 13.640 14.840 13.960 15.160 ;
        RECT 14.040 14.840 14.360 15.160 ;
        RECT 14.440 14.840 14.760 15.160 ;
        RECT 14.840 14.840 15.160 15.160 ;
        RECT 15.240 14.840 15.560 15.160 ;
        RECT 15.640 14.840 15.960 15.160 ;
        RECT 16.040 14.840 16.360 15.160 ;
        RECT 16.440 14.840 16.760 15.160 ;
        RECT 16.840 14.840 17.160 15.160 ;
        RECT 17.240 14.840 17.560 15.160 ;
        RECT 17.640 14.840 17.960 15.160 ;
        RECT 18.040 14.840 18.360 15.160 ;
        RECT 18.440 14.840 18.760 15.160 ;
        RECT 18.840 14.840 19.160 15.160 ;
        RECT 19.240 14.840 19.560 15.160 ;
        RECT 19.640 14.840 19.960 15.160 ;
        RECT 95.560 14.840 95.880 15.160 ;
        RECT 95.960 14.840 96.280 15.160 ;
        RECT 96.360 14.840 96.680 15.160 ;
        RECT 96.760 14.840 97.080 15.160 ;
        RECT 145.560 14.840 145.880 15.160 ;
        RECT 145.960 14.840 146.280 15.160 ;
        RECT 146.360 14.840 146.680 15.160 ;
        RECT 146.760 14.840 147.080 15.160 ;
        RECT 185.720 14.840 186.040 15.160 ;
        RECT 186.120 14.840 186.440 15.160 ;
        RECT 186.520 14.840 186.840 15.160 ;
        RECT 186.920 14.840 187.240 15.160 ;
        RECT 187.320 14.840 187.640 15.160 ;
        RECT 187.720 14.840 188.040 15.160 ;
        RECT 188.120 14.840 188.440 15.160 ;
        RECT 188.520 14.840 188.840 15.160 ;
        RECT 188.920 14.840 189.240 15.160 ;
        RECT 189.320 14.840 189.640 15.160 ;
        RECT 189.720 14.840 190.040 15.160 ;
        RECT 190.120 14.840 190.440 15.160 ;
        RECT 190.520 14.840 190.840 15.160 ;
        RECT 190.920 14.840 191.240 15.160 ;
        RECT 191.320 14.840 191.640 15.160 ;
        RECT 191.720 14.840 192.040 15.160 ;
        RECT 192.120 14.840 192.440 15.160 ;
        RECT 192.520 14.840 192.840 15.160 ;
        RECT 192.920 14.840 193.240 15.160 ;
        RECT 193.320 14.840 193.640 15.160 ;
        RECT 193.720 14.840 194.040 15.160 ;
        RECT 194.120 14.840 194.440 15.160 ;
        RECT 194.520 14.840 194.840 15.160 ;
        RECT 194.920 14.840 195.240 15.160 ;
        RECT 195.320 14.840 195.640 15.160 ;
        RECT 195.720 14.840 196.040 15.160 ;
        RECT 196.120 14.840 196.440 15.160 ;
        RECT 196.520 14.840 196.840 15.160 ;
        RECT 196.920 14.840 197.240 15.160 ;
        RECT 197.320 14.840 197.640 15.160 ;
        RECT 197.720 14.840 198.040 15.160 ;
        RECT 198.120 14.840 198.440 15.160 ;
        RECT 198.520 14.840 198.840 15.160 ;
        RECT 198.920 14.840 199.240 15.160 ;
        RECT 199.320 14.840 199.640 15.160 ;
        RECT 199.720 14.840 200.040 15.160 ;
        RECT 200.120 14.840 200.440 15.160 ;
        RECT 200.520 14.840 200.840 15.160 ;
        RECT 200.920 14.840 201.240 15.160 ;
        RECT 201.320 14.840 201.640 15.160 ;
        RECT 201.720 14.840 202.040 15.160 ;
        RECT 202.120 14.840 202.440 15.160 ;
        RECT 202.520 14.840 202.840 15.160 ;
        RECT 202.920 14.840 203.240 15.160 ;
        RECT 203.320 14.840 203.640 15.160 ;
        RECT 203.720 14.840 204.040 15.160 ;
        RECT 204.120 14.840 204.440 15.160 ;
        RECT 204.520 14.840 204.840 15.160 ;
        RECT 204.920 14.840 205.240 15.160 ;
        RECT 205.320 14.840 205.640 15.160 ;
        RECT 0.040 14.440 0.360 14.760 ;
        RECT 0.440 14.440 0.760 14.760 ;
        RECT 0.840 14.440 1.160 14.760 ;
        RECT 1.240 14.440 1.560 14.760 ;
        RECT 1.640 14.440 1.960 14.760 ;
        RECT 2.040 14.440 2.360 14.760 ;
        RECT 2.440 14.440 2.760 14.760 ;
        RECT 2.840 14.440 3.160 14.760 ;
        RECT 3.240 14.440 3.560 14.760 ;
        RECT 3.640 14.440 3.960 14.760 ;
        RECT 4.040 14.440 4.360 14.760 ;
        RECT 4.440 14.440 4.760 14.760 ;
        RECT 4.840 14.440 5.160 14.760 ;
        RECT 5.240 14.440 5.560 14.760 ;
        RECT 5.640 14.440 5.960 14.760 ;
        RECT 6.040 14.440 6.360 14.760 ;
        RECT 6.440 14.440 6.760 14.760 ;
        RECT 6.840 14.440 7.160 14.760 ;
        RECT 7.240 14.440 7.560 14.760 ;
        RECT 7.640 14.440 7.960 14.760 ;
        RECT 8.040 14.440 8.360 14.760 ;
        RECT 8.440 14.440 8.760 14.760 ;
        RECT 8.840 14.440 9.160 14.760 ;
        RECT 9.240 14.440 9.560 14.760 ;
        RECT 9.640 14.440 9.960 14.760 ;
        RECT 10.040 14.440 10.360 14.760 ;
        RECT 10.440 14.440 10.760 14.760 ;
        RECT 10.840 14.440 11.160 14.760 ;
        RECT 11.240 14.440 11.560 14.760 ;
        RECT 11.640 14.440 11.960 14.760 ;
        RECT 12.040 14.440 12.360 14.760 ;
        RECT 12.440 14.440 12.760 14.760 ;
        RECT 12.840 14.440 13.160 14.760 ;
        RECT 13.240 14.440 13.560 14.760 ;
        RECT 13.640 14.440 13.960 14.760 ;
        RECT 14.040 14.440 14.360 14.760 ;
        RECT 14.440 14.440 14.760 14.760 ;
        RECT 14.840 14.440 15.160 14.760 ;
        RECT 15.240 14.440 15.560 14.760 ;
        RECT 15.640 14.440 15.960 14.760 ;
        RECT 16.040 14.440 16.360 14.760 ;
        RECT 16.440 14.440 16.760 14.760 ;
        RECT 16.840 14.440 17.160 14.760 ;
        RECT 17.240 14.440 17.560 14.760 ;
        RECT 17.640 14.440 17.960 14.760 ;
        RECT 18.040 14.440 18.360 14.760 ;
        RECT 18.440 14.440 18.760 14.760 ;
        RECT 18.840 14.440 19.160 14.760 ;
        RECT 19.240 14.440 19.560 14.760 ;
        RECT 19.640 14.440 19.960 14.760 ;
        RECT 95.560 14.440 95.880 14.760 ;
        RECT 95.960 14.440 96.280 14.760 ;
        RECT 96.360 14.440 96.680 14.760 ;
        RECT 96.760 14.440 97.080 14.760 ;
        RECT 145.560 14.440 145.880 14.760 ;
        RECT 145.960 14.440 146.280 14.760 ;
        RECT 146.360 14.440 146.680 14.760 ;
        RECT 146.760 14.440 147.080 14.760 ;
        RECT 185.720 14.440 186.040 14.760 ;
        RECT 186.120 14.440 186.440 14.760 ;
        RECT 186.520 14.440 186.840 14.760 ;
        RECT 186.920 14.440 187.240 14.760 ;
        RECT 187.320 14.440 187.640 14.760 ;
        RECT 187.720 14.440 188.040 14.760 ;
        RECT 188.120 14.440 188.440 14.760 ;
        RECT 188.520 14.440 188.840 14.760 ;
        RECT 188.920 14.440 189.240 14.760 ;
        RECT 189.320 14.440 189.640 14.760 ;
        RECT 189.720 14.440 190.040 14.760 ;
        RECT 190.120 14.440 190.440 14.760 ;
        RECT 190.520 14.440 190.840 14.760 ;
        RECT 190.920 14.440 191.240 14.760 ;
        RECT 191.320 14.440 191.640 14.760 ;
        RECT 191.720 14.440 192.040 14.760 ;
        RECT 192.120 14.440 192.440 14.760 ;
        RECT 192.520 14.440 192.840 14.760 ;
        RECT 192.920 14.440 193.240 14.760 ;
        RECT 193.320 14.440 193.640 14.760 ;
        RECT 193.720 14.440 194.040 14.760 ;
        RECT 194.120 14.440 194.440 14.760 ;
        RECT 194.520 14.440 194.840 14.760 ;
        RECT 194.920 14.440 195.240 14.760 ;
        RECT 195.320 14.440 195.640 14.760 ;
        RECT 195.720 14.440 196.040 14.760 ;
        RECT 196.120 14.440 196.440 14.760 ;
        RECT 196.520 14.440 196.840 14.760 ;
        RECT 196.920 14.440 197.240 14.760 ;
        RECT 197.320 14.440 197.640 14.760 ;
        RECT 197.720 14.440 198.040 14.760 ;
        RECT 198.120 14.440 198.440 14.760 ;
        RECT 198.520 14.440 198.840 14.760 ;
        RECT 198.920 14.440 199.240 14.760 ;
        RECT 199.320 14.440 199.640 14.760 ;
        RECT 199.720 14.440 200.040 14.760 ;
        RECT 200.120 14.440 200.440 14.760 ;
        RECT 200.520 14.440 200.840 14.760 ;
        RECT 200.920 14.440 201.240 14.760 ;
        RECT 201.320 14.440 201.640 14.760 ;
        RECT 201.720 14.440 202.040 14.760 ;
        RECT 202.120 14.440 202.440 14.760 ;
        RECT 202.520 14.440 202.840 14.760 ;
        RECT 202.920 14.440 203.240 14.760 ;
        RECT 203.320 14.440 203.640 14.760 ;
        RECT 203.720 14.440 204.040 14.760 ;
        RECT 204.120 14.440 204.440 14.760 ;
        RECT 204.520 14.440 204.840 14.760 ;
        RECT 204.920 14.440 205.240 14.760 ;
        RECT 205.320 14.440 205.640 14.760 ;
        RECT 0.040 14.040 0.360 14.360 ;
        RECT 0.440 14.040 0.760 14.360 ;
        RECT 0.840 14.040 1.160 14.360 ;
        RECT 1.240 14.040 1.560 14.360 ;
        RECT 1.640 14.040 1.960 14.360 ;
        RECT 2.040 14.040 2.360 14.360 ;
        RECT 2.440 14.040 2.760 14.360 ;
        RECT 2.840 14.040 3.160 14.360 ;
        RECT 3.240 14.040 3.560 14.360 ;
        RECT 3.640 14.040 3.960 14.360 ;
        RECT 4.040 14.040 4.360 14.360 ;
        RECT 4.440 14.040 4.760 14.360 ;
        RECT 4.840 14.040 5.160 14.360 ;
        RECT 5.240 14.040 5.560 14.360 ;
        RECT 5.640 14.040 5.960 14.360 ;
        RECT 6.040 14.040 6.360 14.360 ;
        RECT 6.440 14.040 6.760 14.360 ;
        RECT 6.840 14.040 7.160 14.360 ;
        RECT 7.240 14.040 7.560 14.360 ;
        RECT 7.640 14.040 7.960 14.360 ;
        RECT 8.040 14.040 8.360 14.360 ;
        RECT 8.440 14.040 8.760 14.360 ;
        RECT 8.840 14.040 9.160 14.360 ;
        RECT 9.240 14.040 9.560 14.360 ;
        RECT 9.640 14.040 9.960 14.360 ;
        RECT 10.040 14.040 10.360 14.360 ;
        RECT 10.440 14.040 10.760 14.360 ;
        RECT 10.840 14.040 11.160 14.360 ;
        RECT 11.240 14.040 11.560 14.360 ;
        RECT 11.640 14.040 11.960 14.360 ;
        RECT 12.040 14.040 12.360 14.360 ;
        RECT 12.440 14.040 12.760 14.360 ;
        RECT 12.840 14.040 13.160 14.360 ;
        RECT 13.240 14.040 13.560 14.360 ;
        RECT 13.640 14.040 13.960 14.360 ;
        RECT 14.040 14.040 14.360 14.360 ;
        RECT 14.440 14.040 14.760 14.360 ;
        RECT 14.840 14.040 15.160 14.360 ;
        RECT 15.240 14.040 15.560 14.360 ;
        RECT 15.640 14.040 15.960 14.360 ;
        RECT 16.040 14.040 16.360 14.360 ;
        RECT 16.440 14.040 16.760 14.360 ;
        RECT 16.840 14.040 17.160 14.360 ;
        RECT 17.240 14.040 17.560 14.360 ;
        RECT 17.640 14.040 17.960 14.360 ;
        RECT 18.040 14.040 18.360 14.360 ;
        RECT 18.440 14.040 18.760 14.360 ;
        RECT 18.840 14.040 19.160 14.360 ;
        RECT 19.240 14.040 19.560 14.360 ;
        RECT 19.640 14.040 19.960 14.360 ;
        RECT 95.560 14.040 95.880 14.360 ;
        RECT 95.960 14.040 96.280 14.360 ;
        RECT 96.360 14.040 96.680 14.360 ;
        RECT 96.760 14.040 97.080 14.360 ;
        RECT 145.560 14.040 145.880 14.360 ;
        RECT 145.960 14.040 146.280 14.360 ;
        RECT 146.360 14.040 146.680 14.360 ;
        RECT 146.760 14.040 147.080 14.360 ;
        RECT 185.720 14.040 186.040 14.360 ;
        RECT 186.120 14.040 186.440 14.360 ;
        RECT 186.520 14.040 186.840 14.360 ;
        RECT 186.920 14.040 187.240 14.360 ;
        RECT 187.320 14.040 187.640 14.360 ;
        RECT 187.720 14.040 188.040 14.360 ;
        RECT 188.120 14.040 188.440 14.360 ;
        RECT 188.520 14.040 188.840 14.360 ;
        RECT 188.920 14.040 189.240 14.360 ;
        RECT 189.320 14.040 189.640 14.360 ;
        RECT 189.720 14.040 190.040 14.360 ;
        RECT 190.120 14.040 190.440 14.360 ;
        RECT 190.520 14.040 190.840 14.360 ;
        RECT 190.920 14.040 191.240 14.360 ;
        RECT 191.320 14.040 191.640 14.360 ;
        RECT 191.720 14.040 192.040 14.360 ;
        RECT 192.120 14.040 192.440 14.360 ;
        RECT 192.520 14.040 192.840 14.360 ;
        RECT 192.920 14.040 193.240 14.360 ;
        RECT 193.320 14.040 193.640 14.360 ;
        RECT 193.720 14.040 194.040 14.360 ;
        RECT 194.120 14.040 194.440 14.360 ;
        RECT 194.520 14.040 194.840 14.360 ;
        RECT 194.920 14.040 195.240 14.360 ;
        RECT 195.320 14.040 195.640 14.360 ;
        RECT 195.720 14.040 196.040 14.360 ;
        RECT 196.120 14.040 196.440 14.360 ;
        RECT 196.520 14.040 196.840 14.360 ;
        RECT 196.920 14.040 197.240 14.360 ;
        RECT 197.320 14.040 197.640 14.360 ;
        RECT 197.720 14.040 198.040 14.360 ;
        RECT 198.120 14.040 198.440 14.360 ;
        RECT 198.520 14.040 198.840 14.360 ;
        RECT 198.920 14.040 199.240 14.360 ;
        RECT 199.320 14.040 199.640 14.360 ;
        RECT 199.720 14.040 200.040 14.360 ;
        RECT 200.120 14.040 200.440 14.360 ;
        RECT 200.520 14.040 200.840 14.360 ;
        RECT 200.920 14.040 201.240 14.360 ;
        RECT 201.320 14.040 201.640 14.360 ;
        RECT 201.720 14.040 202.040 14.360 ;
        RECT 202.120 14.040 202.440 14.360 ;
        RECT 202.520 14.040 202.840 14.360 ;
        RECT 202.920 14.040 203.240 14.360 ;
        RECT 203.320 14.040 203.640 14.360 ;
        RECT 203.720 14.040 204.040 14.360 ;
        RECT 204.120 14.040 204.440 14.360 ;
        RECT 204.520 14.040 204.840 14.360 ;
        RECT 204.920 14.040 205.240 14.360 ;
        RECT 205.320 14.040 205.640 14.360 ;
        RECT 0.040 13.640 0.360 13.960 ;
        RECT 0.440 13.640 0.760 13.960 ;
        RECT 0.840 13.640 1.160 13.960 ;
        RECT 1.240 13.640 1.560 13.960 ;
        RECT 1.640 13.640 1.960 13.960 ;
        RECT 2.040 13.640 2.360 13.960 ;
        RECT 2.440 13.640 2.760 13.960 ;
        RECT 2.840 13.640 3.160 13.960 ;
        RECT 3.240 13.640 3.560 13.960 ;
        RECT 3.640 13.640 3.960 13.960 ;
        RECT 4.040 13.640 4.360 13.960 ;
        RECT 4.440 13.640 4.760 13.960 ;
        RECT 4.840 13.640 5.160 13.960 ;
        RECT 5.240 13.640 5.560 13.960 ;
        RECT 5.640 13.640 5.960 13.960 ;
        RECT 6.040 13.640 6.360 13.960 ;
        RECT 6.440 13.640 6.760 13.960 ;
        RECT 6.840 13.640 7.160 13.960 ;
        RECT 7.240 13.640 7.560 13.960 ;
        RECT 7.640 13.640 7.960 13.960 ;
        RECT 8.040 13.640 8.360 13.960 ;
        RECT 8.440 13.640 8.760 13.960 ;
        RECT 8.840 13.640 9.160 13.960 ;
        RECT 9.240 13.640 9.560 13.960 ;
        RECT 9.640 13.640 9.960 13.960 ;
        RECT 10.040 13.640 10.360 13.960 ;
        RECT 10.440 13.640 10.760 13.960 ;
        RECT 10.840 13.640 11.160 13.960 ;
        RECT 11.240 13.640 11.560 13.960 ;
        RECT 11.640 13.640 11.960 13.960 ;
        RECT 12.040 13.640 12.360 13.960 ;
        RECT 12.440 13.640 12.760 13.960 ;
        RECT 12.840 13.640 13.160 13.960 ;
        RECT 13.240 13.640 13.560 13.960 ;
        RECT 13.640 13.640 13.960 13.960 ;
        RECT 14.040 13.640 14.360 13.960 ;
        RECT 14.440 13.640 14.760 13.960 ;
        RECT 14.840 13.640 15.160 13.960 ;
        RECT 15.240 13.640 15.560 13.960 ;
        RECT 15.640 13.640 15.960 13.960 ;
        RECT 16.040 13.640 16.360 13.960 ;
        RECT 16.440 13.640 16.760 13.960 ;
        RECT 16.840 13.640 17.160 13.960 ;
        RECT 17.240 13.640 17.560 13.960 ;
        RECT 17.640 13.640 17.960 13.960 ;
        RECT 18.040 13.640 18.360 13.960 ;
        RECT 18.440 13.640 18.760 13.960 ;
        RECT 18.840 13.640 19.160 13.960 ;
        RECT 19.240 13.640 19.560 13.960 ;
        RECT 19.640 13.640 19.960 13.960 ;
        RECT 95.560 13.640 95.880 13.960 ;
        RECT 95.960 13.640 96.280 13.960 ;
        RECT 96.360 13.640 96.680 13.960 ;
        RECT 96.760 13.640 97.080 13.960 ;
        RECT 145.560 13.640 145.880 13.960 ;
        RECT 145.960 13.640 146.280 13.960 ;
        RECT 146.360 13.640 146.680 13.960 ;
        RECT 146.760 13.640 147.080 13.960 ;
        RECT 185.720 13.640 186.040 13.960 ;
        RECT 186.120 13.640 186.440 13.960 ;
        RECT 186.520 13.640 186.840 13.960 ;
        RECT 186.920 13.640 187.240 13.960 ;
        RECT 187.320 13.640 187.640 13.960 ;
        RECT 187.720 13.640 188.040 13.960 ;
        RECT 188.120 13.640 188.440 13.960 ;
        RECT 188.520 13.640 188.840 13.960 ;
        RECT 188.920 13.640 189.240 13.960 ;
        RECT 189.320 13.640 189.640 13.960 ;
        RECT 189.720 13.640 190.040 13.960 ;
        RECT 190.120 13.640 190.440 13.960 ;
        RECT 190.520 13.640 190.840 13.960 ;
        RECT 190.920 13.640 191.240 13.960 ;
        RECT 191.320 13.640 191.640 13.960 ;
        RECT 191.720 13.640 192.040 13.960 ;
        RECT 192.120 13.640 192.440 13.960 ;
        RECT 192.520 13.640 192.840 13.960 ;
        RECT 192.920 13.640 193.240 13.960 ;
        RECT 193.320 13.640 193.640 13.960 ;
        RECT 193.720 13.640 194.040 13.960 ;
        RECT 194.120 13.640 194.440 13.960 ;
        RECT 194.520 13.640 194.840 13.960 ;
        RECT 194.920 13.640 195.240 13.960 ;
        RECT 195.320 13.640 195.640 13.960 ;
        RECT 195.720 13.640 196.040 13.960 ;
        RECT 196.120 13.640 196.440 13.960 ;
        RECT 196.520 13.640 196.840 13.960 ;
        RECT 196.920 13.640 197.240 13.960 ;
        RECT 197.320 13.640 197.640 13.960 ;
        RECT 197.720 13.640 198.040 13.960 ;
        RECT 198.120 13.640 198.440 13.960 ;
        RECT 198.520 13.640 198.840 13.960 ;
        RECT 198.920 13.640 199.240 13.960 ;
        RECT 199.320 13.640 199.640 13.960 ;
        RECT 199.720 13.640 200.040 13.960 ;
        RECT 200.120 13.640 200.440 13.960 ;
        RECT 200.520 13.640 200.840 13.960 ;
        RECT 200.920 13.640 201.240 13.960 ;
        RECT 201.320 13.640 201.640 13.960 ;
        RECT 201.720 13.640 202.040 13.960 ;
        RECT 202.120 13.640 202.440 13.960 ;
        RECT 202.520 13.640 202.840 13.960 ;
        RECT 202.920 13.640 203.240 13.960 ;
        RECT 203.320 13.640 203.640 13.960 ;
        RECT 203.720 13.640 204.040 13.960 ;
        RECT 204.120 13.640 204.440 13.960 ;
        RECT 204.520 13.640 204.840 13.960 ;
        RECT 204.920 13.640 205.240 13.960 ;
        RECT 205.320 13.640 205.640 13.960 ;
        RECT 0.040 13.240 0.360 13.560 ;
        RECT 0.440 13.240 0.760 13.560 ;
        RECT 0.840 13.240 1.160 13.560 ;
        RECT 1.240 13.240 1.560 13.560 ;
        RECT 1.640 13.240 1.960 13.560 ;
        RECT 2.040 13.240 2.360 13.560 ;
        RECT 2.440 13.240 2.760 13.560 ;
        RECT 2.840 13.240 3.160 13.560 ;
        RECT 3.240 13.240 3.560 13.560 ;
        RECT 3.640 13.240 3.960 13.560 ;
        RECT 4.040 13.240 4.360 13.560 ;
        RECT 4.440 13.240 4.760 13.560 ;
        RECT 4.840 13.240 5.160 13.560 ;
        RECT 5.240 13.240 5.560 13.560 ;
        RECT 5.640 13.240 5.960 13.560 ;
        RECT 6.040 13.240 6.360 13.560 ;
        RECT 6.440 13.240 6.760 13.560 ;
        RECT 6.840 13.240 7.160 13.560 ;
        RECT 7.240 13.240 7.560 13.560 ;
        RECT 7.640 13.240 7.960 13.560 ;
        RECT 8.040 13.240 8.360 13.560 ;
        RECT 8.440 13.240 8.760 13.560 ;
        RECT 8.840 13.240 9.160 13.560 ;
        RECT 9.240 13.240 9.560 13.560 ;
        RECT 9.640 13.240 9.960 13.560 ;
        RECT 10.040 13.240 10.360 13.560 ;
        RECT 10.440 13.240 10.760 13.560 ;
        RECT 10.840 13.240 11.160 13.560 ;
        RECT 11.240 13.240 11.560 13.560 ;
        RECT 11.640 13.240 11.960 13.560 ;
        RECT 12.040 13.240 12.360 13.560 ;
        RECT 12.440 13.240 12.760 13.560 ;
        RECT 12.840 13.240 13.160 13.560 ;
        RECT 13.240 13.240 13.560 13.560 ;
        RECT 13.640 13.240 13.960 13.560 ;
        RECT 14.040 13.240 14.360 13.560 ;
        RECT 14.440 13.240 14.760 13.560 ;
        RECT 14.840 13.240 15.160 13.560 ;
        RECT 15.240 13.240 15.560 13.560 ;
        RECT 15.640 13.240 15.960 13.560 ;
        RECT 16.040 13.240 16.360 13.560 ;
        RECT 16.440 13.240 16.760 13.560 ;
        RECT 16.840 13.240 17.160 13.560 ;
        RECT 17.240 13.240 17.560 13.560 ;
        RECT 17.640 13.240 17.960 13.560 ;
        RECT 18.040 13.240 18.360 13.560 ;
        RECT 18.440 13.240 18.760 13.560 ;
        RECT 18.840 13.240 19.160 13.560 ;
        RECT 19.240 13.240 19.560 13.560 ;
        RECT 19.640 13.240 19.960 13.560 ;
        RECT 95.560 13.240 95.880 13.560 ;
        RECT 95.960 13.240 96.280 13.560 ;
        RECT 96.360 13.240 96.680 13.560 ;
        RECT 96.760 13.240 97.080 13.560 ;
        RECT 145.560 13.240 145.880 13.560 ;
        RECT 145.960 13.240 146.280 13.560 ;
        RECT 146.360 13.240 146.680 13.560 ;
        RECT 146.760 13.240 147.080 13.560 ;
        RECT 185.720 13.240 186.040 13.560 ;
        RECT 186.120 13.240 186.440 13.560 ;
        RECT 186.520 13.240 186.840 13.560 ;
        RECT 186.920 13.240 187.240 13.560 ;
        RECT 187.320 13.240 187.640 13.560 ;
        RECT 187.720 13.240 188.040 13.560 ;
        RECT 188.120 13.240 188.440 13.560 ;
        RECT 188.520 13.240 188.840 13.560 ;
        RECT 188.920 13.240 189.240 13.560 ;
        RECT 189.320 13.240 189.640 13.560 ;
        RECT 189.720 13.240 190.040 13.560 ;
        RECT 190.120 13.240 190.440 13.560 ;
        RECT 190.520 13.240 190.840 13.560 ;
        RECT 190.920 13.240 191.240 13.560 ;
        RECT 191.320 13.240 191.640 13.560 ;
        RECT 191.720 13.240 192.040 13.560 ;
        RECT 192.120 13.240 192.440 13.560 ;
        RECT 192.520 13.240 192.840 13.560 ;
        RECT 192.920 13.240 193.240 13.560 ;
        RECT 193.320 13.240 193.640 13.560 ;
        RECT 193.720 13.240 194.040 13.560 ;
        RECT 194.120 13.240 194.440 13.560 ;
        RECT 194.520 13.240 194.840 13.560 ;
        RECT 194.920 13.240 195.240 13.560 ;
        RECT 195.320 13.240 195.640 13.560 ;
        RECT 195.720 13.240 196.040 13.560 ;
        RECT 196.120 13.240 196.440 13.560 ;
        RECT 196.520 13.240 196.840 13.560 ;
        RECT 196.920 13.240 197.240 13.560 ;
        RECT 197.320 13.240 197.640 13.560 ;
        RECT 197.720 13.240 198.040 13.560 ;
        RECT 198.120 13.240 198.440 13.560 ;
        RECT 198.520 13.240 198.840 13.560 ;
        RECT 198.920 13.240 199.240 13.560 ;
        RECT 199.320 13.240 199.640 13.560 ;
        RECT 199.720 13.240 200.040 13.560 ;
        RECT 200.120 13.240 200.440 13.560 ;
        RECT 200.520 13.240 200.840 13.560 ;
        RECT 200.920 13.240 201.240 13.560 ;
        RECT 201.320 13.240 201.640 13.560 ;
        RECT 201.720 13.240 202.040 13.560 ;
        RECT 202.120 13.240 202.440 13.560 ;
        RECT 202.520 13.240 202.840 13.560 ;
        RECT 202.920 13.240 203.240 13.560 ;
        RECT 203.320 13.240 203.640 13.560 ;
        RECT 203.720 13.240 204.040 13.560 ;
        RECT 204.120 13.240 204.440 13.560 ;
        RECT 204.520 13.240 204.840 13.560 ;
        RECT 204.920 13.240 205.240 13.560 ;
        RECT 205.320 13.240 205.640 13.560 ;
        RECT 0.040 12.840 0.360 13.160 ;
        RECT 0.440 12.840 0.760 13.160 ;
        RECT 0.840 12.840 1.160 13.160 ;
        RECT 1.240 12.840 1.560 13.160 ;
        RECT 1.640 12.840 1.960 13.160 ;
        RECT 2.040 12.840 2.360 13.160 ;
        RECT 2.440 12.840 2.760 13.160 ;
        RECT 2.840 12.840 3.160 13.160 ;
        RECT 3.240 12.840 3.560 13.160 ;
        RECT 3.640 12.840 3.960 13.160 ;
        RECT 4.040 12.840 4.360 13.160 ;
        RECT 4.440 12.840 4.760 13.160 ;
        RECT 4.840 12.840 5.160 13.160 ;
        RECT 5.240 12.840 5.560 13.160 ;
        RECT 5.640 12.840 5.960 13.160 ;
        RECT 6.040 12.840 6.360 13.160 ;
        RECT 6.440 12.840 6.760 13.160 ;
        RECT 6.840 12.840 7.160 13.160 ;
        RECT 7.240 12.840 7.560 13.160 ;
        RECT 7.640 12.840 7.960 13.160 ;
        RECT 8.040 12.840 8.360 13.160 ;
        RECT 8.440 12.840 8.760 13.160 ;
        RECT 8.840 12.840 9.160 13.160 ;
        RECT 9.240 12.840 9.560 13.160 ;
        RECT 9.640 12.840 9.960 13.160 ;
        RECT 10.040 12.840 10.360 13.160 ;
        RECT 10.440 12.840 10.760 13.160 ;
        RECT 10.840 12.840 11.160 13.160 ;
        RECT 11.240 12.840 11.560 13.160 ;
        RECT 11.640 12.840 11.960 13.160 ;
        RECT 12.040 12.840 12.360 13.160 ;
        RECT 12.440 12.840 12.760 13.160 ;
        RECT 12.840 12.840 13.160 13.160 ;
        RECT 13.240 12.840 13.560 13.160 ;
        RECT 13.640 12.840 13.960 13.160 ;
        RECT 14.040 12.840 14.360 13.160 ;
        RECT 14.440 12.840 14.760 13.160 ;
        RECT 14.840 12.840 15.160 13.160 ;
        RECT 15.240 12.840 15.560 13.160 ;
        RECT 15.640 12.840 15.960 13.160 ;
        RECT 16.040 12.840 16.360 13.160 ;
        RECT 16.440 12.840 16.760 13.160 ;
        RECT 16.840 12.840 17.160 13.160 ;
        RECT 17.240 12.840 17.560 13.160 ;
        RECT 17.640 12.840 17.960 13.160 ;
        RECT 18.040 12.840 18.360 13.160 ;
        RECT 18.440 12.840 18.760 13.160 ;
        RECT 18.840 12.840 19.160 13.160 ;
        RECT 19.240 12.840 19.560 13.160 ;
        RECT 19.640 12.840 19.960 13.160 ;
        RECT 95.560 12.840 95.880 13.160 ;
        RECT 95.960 12.840 96.280 13.160 ;
        RECT 96.360 12.840 96.680 13.160 ;
        RECT 96.760 12.840 97.080 13.160 ;
        RECT 145.560 12.840 145.880 13.160 ;
        RECT 145.960 12.840 146.280 13.160 ;
        RECT 146.360 12.840 146.680 13.160 ;
        RECT 146.760 12.840 147.080 13.160 ;
        RECT 185.720 12.840 186.040 13.160 ;
        RECT 186.120 12.840 186.440 13.160 ;
        RECT 186.520 12.840 186.840 13.160 ;
        RECT 186.920 12.840 187.240 13.160 ;
        RECT 187.320 12.840 187.640 13.160 ;
        RECT 187.720 12.840 188.040 13.160 ;
        RECT 188.120 12.840 188.440 13.160 ;
        RECT 188.520 12.840 188.840 13.160 ;
        RECT 188.920 12.840 189.240 13.160 ;
        RECT 189.320 12.840 189.640 13.160 ;
        RECT 189.720 12.840 190.040 13.160 ;
        RECT 190.120 12.840 190.440 13.160 ;
        RECT 190.520 12.840 190.840 13.160 ;
        RECT 190.920 12.840 191.240 13.160 ;
        RECT 191.320 12.840 191.640 13.160 ;
        RECT 191.720 12.840 192.040 13.160 ;
        RECT 192.120 12.840 192.440 13.160 ;
        RECT 192.520 12.840 192.840 13.160 ;
        RECT 192.920 12.840 193.240 13.160 ;
        RECT 193.320 12.840 193.640 13.160 ;
        RECT 193.720 12.840 194.040 13.160 ;
        RECT 194.120 12.840 194.440 13.160 ;
        RECT 194.520 12.840 194.840 13.160 ;
        RECT 194.920 12.840 195.240 13.160 ;
        RECT 195.320 12.840 195.640 13.160 ;
        RECT 195.720 12.840 196.040 13.160 ;
        RECT 196.120 12.840 196.440 13.160 ;
        RECT 196.520 12.840 196.840 13.160 ;
        RECT 196.920 12.840 197.240 13.160 ;
        RECT 197.320 12.840 197.640 13.160 ;
        RECT 197.720 12.840 198.040 13.160 ;
        RECT 198.120 12.840 198.440 13.160 ;
        RECT 198.520 12.840 198.840 13.160 ;
        RECT 198.920 12.840 199.240 13.160 ;
        RECT 199.320 12.840 199.640 13.160 ;
        RECT 199.720 12.840 200.040 13.160 ;
        RECT 200.120 12.840 200.440 13.160 ;
        RECT 200.520 12.840 200.840 13.160 ;
        RECT 200.920 12.840 201.240 13.160 ;
        RECT 201.320 12.840 201.640 13.160 ;
        RECT 201.720 12.840 202.040 13.160 ;
        RECT 202.120 12.840 202.440 13.160 ;
        RECT 202.520 12.840 202.840 13.160 ;
        RECT 202.920 12.840 203.240 13.160 ;
        RECT 203.320 12.840 203.640 13.160 ;
        RECT 203.720 12.840 204.040 13.160 ;
        RECT 204.120 12.840 204.440 13.160 ;
        RECT 204.520 12.840 204.840 13.160 ;
        RECT 204.920 12.840 205.240 13.160 ;
        RECT 205.320 12.840 205.640 13.160 ;
        RECT 0.040 12.440 0.360 12.760 ;
        RECT 0.440 12.440 0.760 12.760 ;
        RECT 0.840 12.440 1.160 12.760 ;
        RECT 1.240 12.440 1.560 12.760 ;
        RECT 1.640 12.440 1.960 12.760 ;
        RECT 2.040 12.440 2.360 12.760 ;
        RECT 2.440 12.440 2.760 12.760 ;
        RECT 2.840 12.440 3.160 12.760 ;
        RECT 3.240 12.440 3.560 12.760 ;
        RECT 3.640 12.440 3.960 12.760 ;
        RECT 4.040 12.440 4.360 12.760 ;
        RECT 4.440 12.440 4.760 12.760 ;
        RECT 4.840 12.440 5.160 12.760 ;
        RECT 5.240 12.440 5.560 12.760 ;
        RECT 5.640 12.440 5.960 12.760 ;
        RECT 6.040 12.440 6.360 12.760 ;
        RECT 6.440 12.440 6.760 12.760 ;
        RECT 6.840 12.440 7.160 12.760 ;
        RECT 7.240 12.440 7.560 12.760 ;
        RECT 7.640 12.440 7.960 12.760 ;
        RECT 8.040 12.440 8.360 12.760 ;
        RECT 8.440 12.440 8.760 12.760 ;
        RECT 8.840 12.440 9.160 12.760 ;
        RECT 9.240 12.440 9.560 12.760 ;
        RECT 9.640 12.440 9.960 12.760 ;
        RECT 10.040 12.440 10.360 12.760 ;
        RECT 10.440 12.440 10.760 12.760 ;
        RECT 10.840 12.440 11.160 12.760 ;
        RECT 11.240 12.440 11.560 12.760 ;
        RECT 11.640 12.440 11.960 12.760 ;
        RECT 12.040 12.440 12.360 12.760 ;
        RECT 12.440 12.440 12.760 12.760 ;
        RECT 12.840 12.440 13.160 12.760 ;
        RECT 13.240 12.440 13.560 12.760 ;
        RECT 13.640 12.440 13.960 12.760 ;
        RECT 14.040 12.440 14.360 12.760 ;
        RECT 14.440 12.440 14.760 12.760 ;
        RECT 14.840 12.440 15.160 12.760 ;
        RECT 15.240 12.440 15.560 12.760 ;
        RECT 15.640 12.440 15.960 12.760 ;
        RECT 16.040 12.440 16.360 12.760 ;
        RECT 16.440 12.440 16.760 12.760 ;
        RECT 16.840 12.440 17.160 12.760 ;
        RECT 17.240 12.440 17.560 12.760 ;
        RECT 17.640 12.440 17.960 12.760 ;
        RECT 18.040 12.440 18.360 12.760 ;
        RECT 18.440 12.440 18.760 12.760 ;
        RECT 18.840 12.440 19.160 12.760 ;
        RECT 19.240 12.440 19.560 12.760 ;
        RECT 19.640 12.440 19.960 12.760 ;
        RECT 95.560 12.440 95.880 12.760 ;
        RECT 95.960 12.440 96.280 12.760 ;
        RECT 96.360 12.440 96.680 12.760 ;
        RECT 96.760 12.440 97.080 12.760 ;
        RECT 145.560 12.440 145.880 12.760 ;
        RECT 145.960 12.440 146.280 12.760 ;
        RECT 146.360 12.440 146.680 12.760 ;
        RECT 146.760 12.440 147.080 12.760 ;
        RECT 185.720 12.440 186.040 12.760 ;
        RECT 186.120 12.440 186.440 12.760 ;
        RECT 186.520 12.440 186.840 12.760 ;
        RECT 186.920 12.440 187.240 12.760 ;
        RECT 187.320 12.440 187.640 12.760 ;
        RECT 187.720 12.440 188.040 12.760 ;
        RECT 188.120 12.440 188.440 12.760 ;
        RECT 188.520 12.440 188.840 12.760 ;
        RECT 188.920 12.440 189.240 12.760 ;
        RECT 189.320 12.440 189.640 12.760 ;
        RECT 189.720 12.440 190.040 12.760 ;
        RECT 190.120 12.440 190.440 12.760 ;
        RECT 190.520 12.440 190.840 12.760 ;
        RECT 190.920 12.440 191.240 12.760 ;
        RECT 191.320 12.440 191.640 12.760 ;
        RECT 191.720 12.440 192.040 12.760 ;
        RECT 192.120 12.440 192.440 12.760 ;
        RECT 192.520 12.440 192.840 12.760 ;
        RECT 192.920 12.440 193.240 12.760 ;
        RECT 193.320 12.440 193.640 12.760 ;
        RECT 193.720 12.440 194.040 12.760 ;
        RECT 194.120 12.440 194.440 12.760 ;
        RECT 194.520 12.440 194.840 12.760 ;
        RECT 194.920 12.440 195.240 12.760 ;
        RECT 195.320 12.440 195.640 12.760 ;
        RECT 195.720 12.440 196.040 12.760 ;
        RECT 196.120 12.440 196.440 12.760 ;
        RECT 196.520 12.440 196.840 12.760 ;
        RECT 196.920 12.440 197.240 12.760 ;
        RECT 197.320 12.440 197.640 12.760 ;
        RECT 197.720 12.440 198.040 12.760 ;
        RECT 198.120 12.440 198.440 12.760 ;
        RECT 198.520 12.440 198.840 12.760 ;
        RECT 198.920 12.440 199.240 12.760 ;
        RECT 199.320 12.440 199.640 12.760 ;
        RECT 199.720 12.440 200.040 12.760 ;
        RECT 200.120 12.440 200.440 12.760 ;
        RECT 200.520 12.440 200.840 12.760 ;
        RECT 200.920 12.440 201.240 12.760 ;
        RECT 201.320 12.440 201.640 12.760 ;
        RECT 201.720 12.440 202.040 12.760 ;
        RECT 202.120 12.440 202.440 12.760 ;
        RECT 202.520 12.440 202.840 12.760 ;
        RECT 202.920 12.440 203.240 12.760 ;
        RECT 203.320 12.440 203.640 12.760 ;
        RECT 203.720 12.440 204.040 12.760 ;
        RECT 204.120 12.440 204.440 12.760 ;
        RECT 204.520 12.440 204.840 12.760 ;
        RECT 204.920 12.440 205.240 12.760 ;
        RECT 205.320 12.440 205.640 12.760 ;
        RECT 0.040 12.040 0.360 12.360 ;
        RECT 0.440 12.040 0.760 12.360 ;
        RECT 0.840 12.040 1.160 12.360 ;
        RECT 1.240 12.040 1.560 12.360 ;
        RECT 1.640 12.040 1.960 12.360 ;
        RECT 2.040 12.040 2.360 12.360 ;
        RECT 2.440 12.040 2.760 12.360 ;
        RECT 2.840 12.040 3.160 12.360 ;
        RECT 3.240 12.040 3.560 12.360 ;
        RECT 3.640 12.040 3.960 12.360 ;
        RECT 4.040 12.040 4.360 12.360 ;
        RECT 4.440 12.040 4.760 12.360 ;
        RECT 4.840 12.040 5.160 12.360 ;
        RECT 5.240 12.040 5.560 12.360 ;
        RECT 5.640 12.040 5.960 12.360 ;
        RECT 6.040 12.040 6.360 12.360 ;
        RECT 6.440 12.040 6.760 12.360 ;
        RECT 6.840 12.040 7.160 12.360 ;
        RECT 7.240 12.040 7.560 12.360 ;
        RECT 7.640 12.040 7.960 12.360 ;
        RECT 8.040 12.040 8.360 12.360 ;
        RECT 8.440 12.040 8.760 12.360 ;
        RECT 8.840 12.040 9.160 12.360 ;
        RECT 9.240 12.040 9.560 12.360 ;
        RECT 9.640 12.040 9.960 12.360 ;
        RECT 10.040 12.040 10.360 12.360 ;
        RECT 10.440 12.040 10.760 12.360 ;
        RECT 10.840 12.040 11.160 12.360 ;
        RECT 11.240 12.040 11.560 12.360 ;
        RECT 11.640 12.040 11.960 12.360 ;
        RECT 12.040 12.040 12.360 12.360 ;
        RECT 12.440 12.040 12.760 12.360 ;
        RECT 12.840 12.040 13.160 12.360 ;
        RECT 13.240 12.040 13.560 12.360 ;
        RECT 13.640 12.040 13.960 12.360 ;
        RECT 14.040 12.040 14.360 12.360 ;
        RECT 14.440 12.040 14.760 12.360 ;
        RECT 14.840 12.040 15.160 12.360 ;
        RECT 15.240 12.040 15.560 12.360 ;
        RECT 15.640 12.040 15.960 12.360 ;
        RECT 16.040 12.040 16.360 12.360 ;
        RECT 16.440 12.040 16.760 12.360 ;
        RECT 16.840 12.040 17.160 12.360 ;
        RECT 17.240 12.040 17.560 12.360 ;
        RECT 17.640 12.040 17.960 12.360 ;
        RECT 18.040 12.040 18.360 12.360 ;
        RECT 18.440 12.040 18.760 12.360 ;
        RECT 18.840 12.040 19.160 12.360 ;
        RECT 19.240 12.040 19.560 12.360 ;
        RECT 19.640 12.040 19.960 12.360 ;
        RECT 95.560 12.040 95.880 12.360 ;
        RECT 95.960 12.040 96.280 12.360 ;
        RECT 96.360 12.040 96.680 12.360 ;
        RECT 96.760 12.040 97.080 12.360 ;
        RECT 145.560 12.040 145.880 12.360 ;
        RECT 145.960 12.040 146.280 12.360 ;
        RECT 146.360 12.040 146.680 12.360 ;
        RECT 146.760 12.040 147.080 12.360 ;
        RECT 185.720 12.040 186.040 12.360 ;
        RECT 186.120 12.040 186.440 12.360 ;
        RECT 186.520 12.040 186.840 12.360 ;
        RECT 186.920 12.040 187.240 12.360 ;
        RECT 187.320 12.040 187.640 12.360 ;
        RECT 187.720 12.040 188.040 12.360 ;
        RECT 188.120 12.040 188.440 12.360 ;
        RECT 188.520 12.040 188.840 12.360 ;
        RECT 188.920 12.040 189.240 12.360 ;
        RECT 189.320 12.040 189.640 12.360 ;
        RECT 189.720 12.040 190.040 12.360 ;
        RECT 190.120 12.040 190.440 12.360 ;
        RECT 190.520 12.040 190.840 12.360 ;
        RECT 190.920 12.040 191.240 12.360 ;
        RECT 191.320 12.040 191.640 12.360 ;
        RECT 191.720 12.040 192.040 12.360 ;
        RECT 192.120 12.040 192.440 12.360 ;
        RECT 192.520 12.040 192.840 12.360 ;
        RECT 192.920 12.040 193.240 12.360 ;
        RECT 193.320 12.040 193.640 12.360 ;
        RECT 193.720 12.040 194.040 12.360 ;
        RECT 194.120 12.040 194.440 12.360 ;
        RECT 194.520 12.040 194.840 12.360 ;
        RECT 194.920 12.040 195.240 12.360 ;
        RECT 195.320 12.040 195.640 12.360 ;
        RECT 195.720 12.040 196.040 12.360 ;
        RECT 196.120 12.040 196.440 12.360 ;
        RECT 196.520 12.040 196.840 12.360 ;
        RECT 196.920 12.040 197.240 12.360 ;
        RECT 197.320 12.040 197.640 12.360 ;
        RECT 197.720 12.040 198.040 12.360 ;
        RECT 198.120 12.040 198.440 12.360 ;
        RECT 198.520 12.040 198.840 12.360 ;
        RECT 198.920 12.040 199.240 12.360 ;
        RECT 199.320 12.040 199.640 12.360 ;
        RECT 199.720 12.040 200.040 12.360 ;
        RECT 200.120 12.040 200.440 12.360 ;
        RECT 200.520 12.040 200.840 12.360 ;
        RECT 200.920 12.040 201.240 12.360 ;
        RECT 201.320 12.040 201.640 12.360 ;
        RECT 201.720 12.040 202.040 12.360 ;
        RECT 202.120 12.040 202.440 12.360 ;
        RECT 202.520 12.040 202.840 12.360 ;
        RECT 202.920 12.040 203.240 12.360 ;
        RECT 203.320 12.040 203.640 12.360 ;
        RECT 203.720 12.040 204.040 12.360 ;
        RECT 204.120 12.040 204.440 12.360 ;
        RECT 204.520 12.040 204.840 12.360 ;
        RECT 204.920 12.040 205.240 12.360 ;
        RECT 205.320 12.040 205.640 12.360 ;
        RECT 0.040 11.640 0.360 11.960 ;
        RECT 0.440 11.640 0.760 11.960 ;
        RECT 0.840 11.640 1.160 11.960 ;
        RECT 1.240 11.640 1.560 11.960 ;
        RECT 1.640 11.640 1.960 11.960 ;
        RECT 2.040 11.640 2.360 11.960 ;
        RECT 2.440 11.640 2.760 11.960 ;
        RECT 2.840 11.640 3.160 11.960 ;
        RECT 3.240 11.640 3.560 11.960 ;
        RECT 3.640 11.640 3.960 11.960 ;
        RECT 4.040 11.640 4.360 11.960 ;
        RECT 4.440 11.640 4.760 11.960 ;
        RECT 4.840 11.640 5.160 11.960 ;
        RECT 5.240 11.640 5.560 11.960 ;
        RECT 5.640 11.640 5.960 11.960 ;
        RECT 6.040 11.640 6.360 11.960 ;
        RECT 6.440 11.640 6.760 11.960 ;
        RECT 6.840 11.640 7.160 11.960 ;
        RECT 7.240 11.640 7.560 11.960 ;
        RECT 7.640 11.640 7.960 11.960 ;
        RECT 8.040 11.640 8.360 11.960 ;
        RECT 8.440 11.640 8.760 11.960 ;
        RECT 8.840 11.640 9.160 11.960 ;
        RECT 9.240 11.640 9.560 11.960 ;
        RECT 9.640 11.640 9.960 11.960 ;
        RECT 10.040 11.640 10.360 11.960 ;
        RECT 10.440 11.640 10.760 11.960 ;
        RECT 10.840 11.640 11.160 11.960 ;
        RECT 11.240 11.640 11.560 11.960 ;
        RECT 11.640 11.640 11.960 11.960 ;
        RECT 12.040 11.640 12.360 11.960 ;
        RECT 12.440 11.640 12.760 11.960 ;
        RECT 12.840 11.640 13.160 11.960 ;
        RECT 13.240 11.640 13.560 11.960 ;
        RECT 13.640 11.640 13.960 11.960 ;
        RECT 14.040 11.640 14.360 11.960 ;
        RECT 14.440 11.640 14.760 11.960 ;
        RECT 14.840 11.640 15.160 11.960 ;
        RECT 15.240 11.640 15.560 11.960 ;
        RECT 15.640 11.640 15.960 11.960 ;
        RECT 16.040 11.640 16.360 11.960 ;
        RECT 16.440 11.640 16.760 11.960 ;
        RECT 16.840 11.640 17.160 11.960 ;
        RECT 17.240 11.640 17.560 11.960 ;
        RECT 17.640 11.640 17.960 11.960 ;
        RECT 18.040 11.640 18.360 11.960 ;
        RECT 18.440 11.640 18.760 11.960 ;
        RECT 18.840 11.640 19.160 11.960 ;
        RECT 19.240 11.640 19.560 11.960 ;
        RECT 19.640 11.640 19.960 11.960 ;
        RECT 95.560 11.640 95.880 11.960 ;
        RECT 95.960 11.640 96.280 11.960 ;
        RECT 96.360 11.640 96.680 11.960 ;
        RECT 96.760 11.640 97.080 11.960 ;
        RECT 145.560 11.640 145.880 11.960 ;
        RECT 145.960 11.640 146.280 11.960 ;
        RECT 146.360 11.640 146.680 11.960 ;
        RECT 146.760 11.640 147.080 11.960 ;
        RECT 185.720 11.640 186.040 11.960 ;
        RECT 186.120 11.640 186.440 11.960 ;
        RECT 186.520 11.640 186.840 11.960 ;
        RECT 186.920 11.640 187.240 11.960 ;
        RECT 187.320 11.640 187.640 11.960 ;
        RECT 187.720 11.640 188.040 11.960 ;
        RECT 188.120 11.640 188.440 11.960 ;
        RECT 188.520 11.640 188.840 11.960 ;
        RECT 188.920 11.640 189.240 11.960 ;
        RECT 189.320 11.640 189.640 11.960 ;
        RECT 189.720 11.640 190.040 11.960 ;
        RECT 190.120 11.640 190.440 11.960 ;
        RECT 190.520 11.640 190.840 11.960 ;
        RECT 190.920 11.640 191.240 11.960 ;
        RECT 191.320 11.640 191.640 11.960 ;
        RECT 191.720 11.640 192.040 11.960 ;
        RECT 192.120 11.640 192.440 11.960 ;
        RECT 192.520 11.640 192.840 11.960 ;
        RECT 192.920 11.640 193.240 11.960 ;
        RECT 193.320 11.640 193.640 11.960 ;
        RECT 193.720 11.640 194.040 11.960 ;
        RECT 194.120 11.640 194.440 11.960 ;
        RECT 194.520 11.640 194.840 11.960 ;
        RECT 194.920 11.640 195.240 11.960 ;
        RECT 195.320 11.640 195.640 11.960 ;
        RECT 195.720 11.640 196.040 11.960 ;
        RECT 196.120 11.640 196.440 11.960 ;
        RECT 196.520 11.640 196.840 11.960 ;
        RECT 196.920 11.640 197.240 11.960 ;
        RECT 197.320 11.640 197.640 11.960 ;
        RECT 197.720 11.640 198.040 11.960 ;
        RECT 198.120 11.640 198.440 11.960 ;
        RECT 198.520 11.640 198.840 11.960 ;
        RECT 198.920 11.640 199.240 11.960 ;
        RECT 199.320 11.640 199.640 11.960 ;
        RECT 199.720 11.640 200.040 11.960 ;
        RECT 200.120 11.640 200.440 11.960 ;
        RECT 200.520 11.640 200.840 11.960 ;
        RECT 200.920 11.640 201.240 11.960 ;
        RECT 201.320 11.640 201.640 11.960 ;
        RECT 201.720 11.640 202.040 11.960 ;
        RECT 202.120 11.640 202.440 11.960 ;
        RECT 202.520 11.640 202.840 11.960 ;
        RECT 202.920 11.640 203.240 11.960 ;
        RECT 203.320 11.640 203.640 11.960 ;
        RECT 203.720 11.640 204.040 11.960 ;
        RECT 204.120 11.640 204.440 11.960 ;
        RECT 204.520 11.640 204.840 11.960 ;
        RECT 204.920 11.640 205.240 11.960 ;
        RECT 205.320 11.640 205.640 11.960 ;
        RECT 0.040 11.240 0.360 11.560 ;
        RECT 0.440 11.240 0.760 11.560 ;
        RECT 0.840 11.240 1.160 11.560 ;
        RECT 1.240 11.240 1.560 11.560 ;
        RECT 1.640 11.240 1.960 11.560 ;
        RECT 2.040 11.240 2.360 11.560 ;
        RECT 2.440 11.240 2.760 11.560 ;
        RECT 2.840 11.240 3.160 11.560 ;
        RECT 3.240 11.240 3.560 11.560 ;
        RECT 3.640 11.240 3.960 11.560 ;
        RECT 4.040 11.240 4.360 11.560 ;
        RECT 4.440 11.240 4.760 11.560 ;
        RECT 4.840 11.240 5.160 11.560 ;
        RECT 5.240 11.240 5.560 11.560 ;
        RECT 5.640 11.240 5.960 11.560 ;
        RECT 6.040 11.240 6.360 11.560 ;
        RECT 6.440 11.240 6.760 11.560 ;
        RECT 6.840 11.240 7.160 11.560 ;
        RECT 7.240 11.240 7.560 11.560 ;
        RECT 7.640 11.240 7.960 11.560 ;
        RECT 8.040 11.240 8.360 11.560 ;
        RECT 8.440 11.240 8.760 11.560 ;
        RECT 8.840 11.240 9.160 11.560 ;
        RECT 9.240 11.240 9.560 11.560 ;
        RECT 9.640 11.240 9.960 11.560 ;
        RECT 10.040 11.240 10.360 11.560 ;
        RECT 10.440 11.240 10.760 11.560 ;
        RECT 10.840 11.240 11.160 11.560 ;
        RECT 11.240 11.240 11.560 11.560 ;
        RECT 11.640 11.240 11.960 11.560 ;
        RECT 12.040 11.240 12.360 11.560 ;
        RECT 12.440 11.240 12.760 11.560 ;
        RECT 12.840 11.240 13.160 11.560 ;
        RECT 13.240 11.240 13.560 11.560 ;
        RECT 13.640 11.240 13.960 11.560 ;
        RECT 14.040 11.240 14.360 11.560 ;
        RECT 14.440 11.240 14.760 11.560 ;
        RECT 14.840 11.240 15.160 11.560 ;
        RECT 15.240 11.240 15.560 11.560 ;
        RECT 15.640 11.240 15.960 11.560 ;
        RECT 16.040 11.240 16.360 11.560 ;
        RECT 16.440 11.240 16.760 11.560 ;
        RECT 16.840 11.240 17.160 11.560 ;
        RECT 17.240 11.240 17.560 11.560 ;
        RECT 17.640 11.240 17.960 11.560 ;
        RECT 18.040 11.240 18.360 11.560 ;
        RECT 18.440 11.240 18.760 11.560 ;
        RECT 18.840 11.240 19.160 11.560 ;
        RECT 19.240 11.240 19.560 11.560 ;
        RECT 19.640 11.240 19.960 11.560 ;
        RECT 95.560 11.240 95.880 11.560 ;
        RECT 95.960 11.240 96.280 11.560 ;
        RECT 96.360 11.240 96.680 11.560 ;
        RECT 96.760 11.240 97.080 11.560 ;
        RECT 145.560 11.240 145.880 11.560 ;
        RECT 145.960 11.240 146.280 11.560 ;
        RECT 146.360 11.240 146.680 11.560 ;
        RECT 146.760 11.240 147.080 11.560 ;
        RECT 185.720 11.240 186.040 11.560 ;
        RECT 186.120 11.240 186.440 11.560 ;
        RECT 186.520 11.240 186.840 11.560 ;
        RECT 186.920 11.240 187.240 11.560 ;
        RECT 187.320 11.240 187.640 11.560 ;
        RECT 187.720 11.240 188.040 11.560 ;
        RECT 188.120 11.240 188.440 11.560 ;
        RECT 188.520 11.240 188.840 11.560 ;
        RECT 188.920 11.240 189.240 11.560 ;
        RECT 189.320 11.240 189.640 11.560 ;
        RECT 189.720 11.240 190.040 11.560 ;
        RECT 190.120 11.240 190.440 11.560 ;
        RECT 190.520 11.240 190.840 11.560 ;
        RECT 190.920 11.240 191.240 11.560 ;
        RECT 191.320 11.240 191.640 11.560 ;
        RECT 191.720 11.240 192.040 11.560 ;
        RECT 192.120 11.240 192.440 11.560 ;
        RECT 192.520 11.240 192.840 11.560 ;
        RECT 192.920 11.240 193.240 11.560 ;
        RECT 193.320 11.240 193.640 11.560 ;
        RECT 193.720 11.240 194.040 11.560 ;
        RECT 194.120 11.240 194.440 11.560 ;
        RECT 194.520 11.240 194.840 11.560 ;
        RECT 194.920 11.240 195.240 11.560 ;
        RECT 195.320 11.240 195.640 11.560 ;
        RECT 195.720 11.240 196.040 11.560 ;
        RECT 196.120 11.240 196.440 11.560 ;
        RECT 196.520 11.240 196.840 11.560 ;
        RECT 196.920 11.240 197.240 11.560 ;
        RECT 197.320 11.240 197.640 11.560 ;
        RECT 197.720 11.240 198.040 11.560 ;
        RECT 198.120 11.240 198.440 11.560 ;
        RECT 198.520 11.240 198.840 11.560 ;
        RECT 198.920 11.240 199.240 11.560 ;
        RECT 199.320 11.240 199.640 11.560 ;
        RECT 199.720 11.240 200.040 11.560 ;
        RECT 200.120 11.240 200.440 11.560 ;
        RECT 200.520 11.240 200.840 11.560 ;
        RECT 200.920 11.240 201.240 11.560 ;
        RECT 201.320 11.240 201.640 11.560 ;
        RECT 201.720 11.240 202.040 11.560 ;
        RECT 202.120 11.240 202.440 11.560 ;
        RECT 202.520 11.240 202.840 11.560 ;
        RECT 202.920 11.240 203.240 11.560 ;
        RECT 203.320 11.240 203.640 11.560 ;
        RECT 203.720 11.240 204.040 11.560 ;
        RECT 204.120 11.240 204.440 11.560 ;
        RECT 204.520 11.240 204.840 11.560 ;
        RECT 204.920 11.240 205.240 11.560 ;
        RECT 205.320 11.240 205.640 11.560 ;
        RECT 0.040 10.840 0.360 11.160 ;
        RECT 0.440 10.840 0.760 11.160 ;
        RECT 0.840 10.840 1.160 11.160 ;
        RECT 1.240 10.840 1.560 11.160 ;
        RECT 1.640 10.840 1.960 11.160 ;
        RECT 2.040 10.840 2.360 11.160 ;
        RECT 2.440 10.840 2.760 11.160 ;
        RECT 2.840 10.840 3.160 11.160 ;
        RECT 3.240 10.840 3.560 11.160 ;
        RECT 3.640 10.840 3.960 11.160 ;
        RECT 4.040 10.840 4.360 11.160 ;
        RECT 4.440 10.840 4.760 11.160 ;
        RECT 4.840 10.840 5.160 11.160 ;
        RECT 5.240 10.840 5.560 11.160 ;
        RECT 5.640 10.840 5.960 11.160 ;
        RECT 6.040 10.840 6.360 11.160 ;
        RECT 6.440 10.840 6.760 11.160 ;
        RECT 6.840 10.840 7.160 11.160 ;
        RECT 7.240 10.840 7.560 11.160 ;
        RECT 7.640 10.840 7.960 11.160 ;
        RECT 8.040 10.840 8.360 11.160 ;
        RECT 8.440 10.840 8.760 11.160 ;
        RECT 8.840 10.840 9.160 11.160 ;
        RECT 9.240 10.840 9.560 11.160 ;
        RECT 9.640 10.840 9.960 11.160 ;
        RECT 10.040 10.840 10.360 11.160 ;
        RECT 10.440 10.840 10.760 11.160 ;
        RECT 10.840 10.840 11.160 11.160 ;
        RECT 11.240 10.840 11.560 11.160 ;
        RECT 11.640 10.840 11.960 11.160 ;
        RECT 12.040 10.840 12.360 11.160 ;
        RECT 12.440 10.840 12.760 11.160 ;
        RECT 12.840 10.840 13.160 11.160 ;
        RECT 13.240 10.840 13.560 11.160 ;
        RECT 13.640 10.840 13.960 11.160 ;
        RECT 14.040 10.840 14.360 11.160 ;
        RECT 14.440 10.840 14.760 11.160 ;
        RECT 14.840 10.840 15.160 11.160 ;
        RECT 15.240 10.840 15.560 11.160 ;
        RECT 15.640 10.840 15.960 11.160 ;
        RECT 16.040 10.840 16.360 11.160 ;
        RECT 16.440 10.840 16.760 11.160 ;
        RECT 16.840 10.840 17.160 11.160 ;
        RECT 17.240 10.840 17.560 11.160 ;
        RECT 17.640 10.840 17.960 11.160 ;
        RECT 18.040 10.840 18.360 11.160 ;
        RECT 18.440 10.840 18.760 11.160 ;
        RECT 18.840 10.840 19.160 11.160 ;
        RECT 19.240 10.840 19.560 11.160 ;
        RECT 19.640 10.840 19.960 11.160 ;
        RECT 95.560 10.840 95.880 11.160 ;
        RECT 95.960 10.840 96.280 11.160 ;
        RECT 96.360 10.840 96.680 11.160 ;
        RECT 96.760 10.840 97.080 11.160 ;
        RECT 145.560 10.840 145.880 11.160 ;
        RECT 145.960 10.840 146.280 11.160 ;
        RECT 146.360 10.840 146.680 11.160 ;
        RECT 146.760 10.840 147.080 11.160 ;
        RECT 185.720 10.840 186.040 11.160 ;
        RECT 186.120 10.840 186.440 11.160 ;
        RECT 186.520 10.840 186.840 11.160 ;
        RECT 186.920 10.840 187.240 11.160 ;
        RECT 187.320 10.840 187.640 11.160 ;
        RECT 187.720 10.840 188.040 11.160 ;
        RECT 188.120 10.840 188.440 11.160 ;
        RECT 188.520 10.840 188.840 11.160 ;
        RECT 188.920 10.840 189.240 11.160 ;
        RECT 189.320 10.840 189.640 11.160 ;
        RECT 189.720 10.840 190.040 11.160 ;
        RECT 190.120 10.840 190.440 11.160 ;
        RECT 190.520 10.840 190.840 11.160 ;
        RECT 190.920 10.840 191.240 11.160 ;
        RECT 191.320 10.840 191.640 11.160 ;
        RECT 191.720 10.840 192.040 11.160 ;
        RECT 192.120 10.840 192.440 11.160 ;
        RECT 192.520 10.840 192.840 11.160 ;
        RECT 192.920 10.840 193.240 11.160 ;
        RECT 193.320 10.840 193.640 11.160 ;
        RECT 193.720 10.840 194.040 11.160 ;
        RECT 194.120 10.840 194.440 11.160 ;
        RECT 194.520 10.840 194.840 11.160 ;
        RECT 194.920 10.840 195.240 11.160 ;
        RECT 195.320 10.840 195.640 11.160 ;
        RECT 195.720 10.840 196.040 11.160 ;
        RECT 196.120 10.840 196.440 11.160 ;
        RECT 196.520 10.840 196.840 11.160 ;
        RECT 196.920 10.840 197.240 11.160 ;
        RECT 197.320 10.840 197.640 11.160 ;
        RECT 197.720 10.840 198.040 11.160 ;
        RECT 198.120 10.840 198.440 11.160 ;
        RECT 198.520 10.840 198.840 11.160 ;
        RECT 198.920 10.840 199.240 11.160 ;
        RECT 199.320 10.840 199.640 11.160 ;
        RECT 199.720 10.840 200.040 11.160 ;
        RECT 200.120 10.840 200.440 11.160 ;
        RECT 200.520 10.840 200.840 11.160 ;
        RECT 200.920 10.840 201.240 11.160 ;
        RECT 201.320 10.840 201.640 11.160 ;
        RECT 201.720 10.840 202.040 11.160 ;
        RECT 202.120 10.840 202.440 11.160 ;
        RECT 202.520 10.840 202.840 11.160 ;
        RECT 202.920 10.840 203.240 11.160 ;
        RECT 203.320 10.840 203.640 11.160 ;
        RECT 203.720 10.840 204.040 11.160 ;
        RECT 204.120 10.840 204.440 11.160 ;
        RECT 204.520 10.840 204.840 11.160 ;
        RECT 204.920 10.840 205.240 11.160 ;
        RECT 205.320 10.840 205.640 11.160 ;
        RECT 0.040 10.440 0.360 10.760 ;
        RECT 0.440 10.440 0.760 10.760 ;
        RECT 0.840 10.440 1.160 10.760 ;
        RECT 1.240 10.440 1.560 10.760 ;
        RECT 1.640 10.440 1.960 10.760 ;
        RECT 2.040 10.440 2.360 10.760 ;
        RECT 2.440 10.440 2.760 10.760 ;
        RECT 2.840 10.440 3.160 10.760 ;
        RECT 3.240 10.440 3.560 10.760 ;
        RECT 3.640 10.440 3.960 10.760 ;
        RECT 4.040 10.440 4.360 10.760 ;
        RECT 4.440 10.440 4.760 10.760 ;
        RECT 4.840 10.440 5.160 10.760 ;
        RECT 5.240 10.440 5.560 10.760 ;
        RECT 5.640 10.440 5.960 10.760 ;
        RECT 6.040 10.440 6.360 10.760 ;
        RECT 6.440 10.440 6.760 10.760 ;
        RECT 6.840 10.440 7.160 10.760 ;
        RECT 7.240 10.440 7.560 10.760 ;
        RECT 7.640 10.440 7.960 10.760 ;
        RECT 8.040 10.440 8.360 10.760 ;
        RECT 8.440 10.440 8.760 10.760 ;
        RECT 8.840 10.440 9.160 10.760 ;
        RECT 9.240 10.440 9.560 10.760 ;
        RECT 9.640 10.440 9.960 10.760 ;
        RECT 10.040 10.440 10.360 10.760 ;
        RECT 10.440 10.440 10.760 10.760 ;
        RECT 10.840 10.440 11.160 10.760 ;
        RECT 11.240 10.440 11.560 10.760 ;
        RECT 11.640 10.440 11.960 10.760 ;
        RECT 12.040 10.440 12.360 10.760 ;
        RECT 12.440 10.440 12.760 10.760 ;
        RECT 12.840 10.440 13.160 10.760 ;
        RECT 13.240 10.440 13.560 10.760 ;
        RECT 13.640 10.440 13.960 10.760 ;
        RECT 14.040 10.440 14.360 10.760 ;
        RECT 14.440 10.440 14.760 10.760 ;
        RECT 14.840 10.440 15.160 10.760 ;
        RECT 15.240 10.440 15.560 10.760 ;
        RECT 15.640 10.440 15.960 10.760 ;
        RECT 16.040 10.440 16.360 10.760 ;
        RECT 16.440 10.440 16.760 10.760 ;
        RECT 16.840 10.440 17.160 10.760 ;
        RECT 17.240 10.440 17.560 10.760 ;
        RECT 17.640 10.440 17.960 10.760 ;
        RECT 18.040 10.440 18.360 10.760 ;
        RECT 18.440 10.440 18.760 10.760 ;
        RECT 18.840 10.440 19.160 10.760 ;
        RECT 19.240 10.440 19.560 10.760 ;
        RECT 19.640 10.440 19.960 10.760 ;
        RECT 95.560 10.440 95.880 10.760 ;
        RECT 95.960 10.440 96.280 10.760 ;
        RECT 96.360 10.440 96.680 10.760 ;
        RECT 96.760 10.440 97.080 10.760 ;
        RECT 145.560 10.440 145.880 10.760 ;
        RECT 145.960 10.440 146.280 10.760 ;
        RECT 146.360 10.440 146.680 10.760 ;
        RECT 146.760 10.440 147.080 10.760 ;
        RECT 185.720 10.440 186.040 10.760 ;
        RECT 186.120 10.440 186.440 10.760 ;
        RECT 186.520 10.440 186.840 10.760 ;
        RECT 186.920 10.440 187.240 10.760 ;
        RECT 187.320 10.440 187.640 10.760 ;
        RECT 187.720 10.440 188.040 10.760 ;
        RECT 188.120 10.440 188.440 10.760 ;
        RECT 188.520 10.440 188.840 10.760 ;
        RECT 188.920 10.440 189.240 10.760 ;
        RECT 189.320 10.440 189.640 10.760 ;
        RECT 189.720 10.440 190.040 10.760 ;
        RECT 190.120 10.440 190.440 10.760 ;
        RECT 190.520 10.440 190.840 10.760 ;
        RECT 190.920 10.440 191.240 10.760 ;
        RECT 191.320 10.440 191.640 10.760 ;
        RECT 191.720 10.440 192.040 10.760 ;
        RECT 192.120 10.440 192.440 10.760 ;
        RECT 192.520 10.440 192.840 10.760 ;
        RECT 192.920 10.440 193.240 10.760 ;
        RECT 193.320 10.440 193.640 10.760 ;
        RECT 193.720 10.440 194.040 10.760 ;
        RECT 194.120 10.440 194.440 10.760 ;
        RECT 194.520 10.440 194.840 10.760 ;
        RECT 194.920 10.440 195.240 10.760 ;
        RECT 195.320 10.440 195.640 10.760 ;
        RECT 195.720 10.440 196.040 10.760 ;
        RECT 196.120 10.440 196.440 10.760 ;
        RECT 196.520 10.440 196.840 10.760 ;
        RECT 196.920 10.440 197.240 10.760 ;
        RECT 197.320 10.440 197.640 10.760 ;
        RECT 197.720 10.440 198.040 10.760 ;
        RECT 198.120 10.440 198.440 10.760 ;
        RECT 198.520 10.440 198.840 10.760 ;
        RECT 198.920 10.440 199.240 10.760 ;
        RECT 199.320 10.440 199.640 10.760 ;
        RECT 199.720 10.440 200.040 10.760 ;
        RECT 200.120 10.440 200.440 10.760 ;
        RECT 200.520 10.440 200.840 10.760 ;
        RECT 200.920 10.440 201.240 10.760 ;
        RECT 201.320 10.440 201.640 10.760 ;
        RECT 201.720 10.440 202.040 10.760 ;
        RECT 202.120 10.440 202.440 10.760 ;
        RECT 202.520 10.440 202.840 10.760 ;
        RECT 202.920 10.440 203.240 10.760 ;
        RECT 203.320 10.440 203.640 10.760 ;
        RECT 203.720 10.440 204.040 10.760 ;
        RECT 204.120 10.440 204.440 10.760 ;
        RECT 204.520 10.440 204.840 10.760 ;
        RECT 204.920 10.440 205.240 10.760 ;
        RECT 205.320 10.440 205.640 10.760 ;
        RECT 0.040 10.040 0.360 10.360 ;
        RECT 0.440 10.040 0.760 10.360 ;
        RECT 0.840 10.040 1.160 10.360 ;
        RECT 1.240 10.040 1.560 10.360 ;
        RECT 1.640 10.040 1.960 10.360 ;
        RECT 2.040 10.040 2.360 10.360 ;
        RECT 2.440 10.040 2.760 10.360 ;
        RECT 2.840 10.040 3.160 10.360 ;
        RECT 3.240 10.040 3.560 10.360 ;
        RECT 3.640 10.040 3.960 10.360 ;
        RECT 4.040 10.040 4.360 10.360 ;
        RECT 4.440 10.040 4.760 10.360 ;
        RECT 4.840 10.040 5.160 10.360 ;
        RECT 5.240 10.040 5.560 10.360 ;
        RECT 5.640 10.040 5.960 10.360 ;
        RECT 6.040 10.040 6.360 10.360 ;
        RECT 6.440 10.040 6.760 10.360 ;
        RECT 6.840 10.040 7.160 10.360 ;
        RECT 7.240 10.040 7.560 10.360 ;
        RECT 7.640 10.040 7.960 10.360 ;
        RECT 8.040 10.040 8.360 10.360 ;
        RECT 8.440 10.040 8.760 10.360 ;
        RECT 8.840 10.040 9.160 10.360 ;
        RECT 9.240 10.040 9.560 10.360 ;
        RECT 9.640 10.040 9.960 10.360 ;
        RECT 10.040 10.040 10.360 10.360 ;
        RECT 10.440 10.040 10.760 10.360 ;
        RECT 10.840 10.040 11.160 10.360 ;
        RECT 11.240 10.040 11.560 10.360 ;
        RECT 11.640 10.040 11.960 10.360 ;
        RECT 12.040 10.040 12.360 10.360 ;
        RECT 12.440 10.040 12.760 10.360 ;
        RECT 12.840 10.040 13.160 10.360 ;
        RECT 13.240 10.040 13.560 10.360 ;
        RECT 13.640 10.040 13.960 10.360 ;
        RECT 14.040 10.040 14.360 10.360 ;
        RECT 14.440 10.040 14.760 10.360 ;
        RECT 14.840 10.040 15.160 10.360 ;
        RECT 15.240 10.040 15.560 10.360 ;
        RECT 15.640 10.040 15.960 10.360 ;
        RECT 16.040 10.040 16.360 10.360 ;
        RECT 16.440 10.040 16.760 10.360 ;
        RECT 16.840 10.040 17.160 10.360 ;
        RECT 17.240 10.040 17.560 10.360 ;
        RECT 17.640 10.040 17.960 10.360 ;
        RECT 18.040 10.040 18.360 10.360 ;
        RECT 18.440 10.040 18.760 10.360 ;
        RECT 18.840 10.040 19.160 10.360 ;
        RECT 19.240 10.040 19.560 10.360 ;
        RECT 19.640 10.040 19.960 10.360 ;
        RECT 95.560 10.040 95.880 10.360 ;
        RECT 95.960 10.040 96.280 10.360 ;
        RECT 96.360 10.040 96.680 10.360 ;
        RECT 96.760 10.040 97.080 10.360 ;
        RECT 145.560 10.040 145.880 10.360 ;
        RECT 145.960 10.040 146.280 10.360 ;
        RECT 146.360 10.040 146.680 10.360 ;
        RECT 146.760 10.040 147.080 10.360 ;
        RECT 185.720 10.040 186.040 10.360 ;
        RECT 186.120 10.040 186.440 10.360 ;
        RECT 186.520 10.040 186.840 10.360 ;
        RECT 186.920 10.040 187.240 10.360 ;
        RECT 187.320 10.040 187.640 10.360 ;
        RECT 187.720 10.040 188.040 10.360 ;
        RECT 188.120 10.040 188.440 10.360 ;
        RECT 188.520 10.040 188.840 10.360 ;
        RECT 188.920 10.040 189.240 10.360 ;
        RECT 189.320 10.040 189.640 10.360 ;
        RECT 189.720 10.040 190.040 10.360 ;
        RECT 190.120 10.040 190.440 10.360 ;
        RECT 190.520 10.040 190.840 10.360 ;
        RECT 190.920 10.040 191.240 10.360 ;
        RECT 191.320 10.040 191.640 10.360 ;
        RECT 191.720 10.040 192.040 10.360 ;
        RECT 192.120 10.040 192.440 10.360 ;
        RECT 192.520 10.040 192.840 10.360 ;
        RECT 192.920 10.040 193.240 10.360 ;
        RECT 193.320 10.040 193.640 10.360 ;
        RECT 193.720 10.040 194.040 10.360 ;
        RECT 194.120 10.040 194.440 10.360 ;
        RECT 194.520 10.040 194.840 10.360 ;
        RECT 194.920 10.040 195.240 10.360 ;
        RECT 195.320 10.040 195.640 10.360 ;
        RECT 195.720 10.040 196.040 10.360 ;
        RECT 196.120 10.040 196.440 10.360 ;
        RECT 196.520 10.040 196.840 10.360 ;
        RECT 196.920 10.040 197.240 10.360 ;
        RECT 197.320 10.040 197.640 10.360 ;
        RECT 197.720 10.040 198.040 10.360 ;
        RECT 198.120 10.040 198.440 10.360 ;
        RECT 198.520 10.040 198.840 10.360 ;
        RECT 198.920 10.040 199.240 10.360 ;
        RECT 199.320 10.040 199.640 10.360 ;
        RECT 199.720 10.040 200.040 10.360 ;
        RECT 200.120 10.040 200.440 10.360 ;
        RECT 200.520 10.040 200.840 10.360 ;
        RECT 200.920 10.040 201.240 10.360 ;
        RECT 201.320 10.040 201.640 10.360 ;
        RECT 201.720 10.040 202.040 10.360 ;
        RECT 202.120 10.040 202.440 10.360 ;
        RECT 202.520 10.040 202.840 10.360 ;
        RECT 202.920 10.040 203.240 10.360 ;
        RECT 203.320 10.040 203.640 10.360 ;
        RECT 203.720 10.040 204.040 10.360 ;
        RECT 204.120 10.040 204.440 10.360 ;
        RECT 204.520 10.040 204.840 10.360 ;
        RECT 204.920 10.040 205.240 10.360 ;
        RECT 205.320 10.040 205.640 10.360 ;
        RECT 0.040 9.640 0.360 9.960 ;
        RECT 0.440 9.640 0.760 9.960 ;
        RECT 0.840 9.640 1.160 9.960 ;
        RECT 1.240 9.640 1.560 9.960 ;
        RECT 1.640 9.640 1.960 9.960 ;
        RECT 2.040 9.640 2.360 9.960 ;
        RECT 2.440 9.640 2.760 9.960 ;
        RECT 2.840 9.640 3.160 9.960 ;
        RECT 3.240 9.640 3.560 9.960 ;
        RECT 3.640 9.640 3.960 9.960 ;
        RECT 4.040 9.640 4.360 9.960 ;
        RECT 4.440 9.640 4.760 9.960 ;
        RECT 4.840 9.640 5.160 9.960 ;
        RECT 5.240 9.640 5.560 9.960 ;
        RECT 5.640 9.640 5.960 9.960 ;
        RECT 6.040 9.640 6.360 9.960 ;
        RECT 6.440 9.640 6.760 9.960 ;
        RECT 6.840 9.640 7.160 9.960 ;
        RECT 7.240 9.640 7.560 9.960 ;
        RECT 7.640 9.640 7.960 9.960 ;
        RECT 8.040 9.640 8.360 9.960 ;
        RECT 8.440 9.640 8.760 9.960 ;
        RECT 8.840 9.640 9.160 9.960 ;
        RECT 9.240 9.640 9.560 9.960 ;
        RECT 9.640 9.640 9.960 9.960 ;
        RECT 10.040 9.640 10.360 9.960 ;
        RECT 10.440 9.640 10.760 9.960 ;
        RECT 10.840 9.640 11.160 9.960 ;
        RECT 11.240 9.640 11.560 9.960 ;
        RECT 11.640 9.640 11.960 9.960 ;
        RECT 12.040 9.640 12.360 9.960 ;
        RECT 12.440 9.640 12.760 9.960 ;
        RECT 12.840 9.640 13.160 9.960 ;
        RECT 13.240 9.640 13.560 9.960 ;
        RECT 13.640 9.640 13.960 9.960 ;
        RECT 14.040 9.640 14.360 9.960 ;
        RECT 14.440 9.640 14.760 9.960 ;
        RECT 14.840 9.640 15.160 9.960 ;
        RECT 15.240 9.640 15.560 9.960 ;
        RECT 15.640 9.640 15.960 9.960 ;
        RECT 16.040 9.640 16.360 9.960 ;
        RECT 16.440 9.640 16.760 9.960 ;
        RECT 16.840 9.640 17.160 9.960 ;
        RECT 17.240 9.640 17.560 9.960 ;
        RECT 17.640 9.640 17.960 9.960 ;
        RECT 18.040 9.640 18.360 9.960 ;
        RECT 18.440 9.640 18.760 9.960 ;
        RECT 18.840 9.640 19.160 9.960 ;
        RECT 19.240 9.640 19.560 9.960 ;
        RECT 19.640 9.640 19.960 9.960 ;
        RECT 95.560 9.640 95.880 9.960 ;
        RECT 95.960 9.640 96.280 9.960 ;
        RECT 96.360 9.640 96.680 9.960 ;
        RECT 96.760 9.640 97.080 9.960 ;
        RECT 145.560 9.640 145.880 9.960 ;
        RECT 145.960 9.640 146.280 9.960 ;
        RECT 146.360 9.640 146.680 9.960 ;
        RECT 146.760 9.640 147.080 9.960 ;
        RECT 185.720 9.640 186.040 9.960 ;
        RECT 186.120 9.640 186.440 9.960 ;
        RECT 186.520 9.640 186.840 9.960 ;
        RECT 186.920 9.640 187.240 9.960 ;
        RECT 187.320 9.640 187.640 9.960 ;
        RECT 187.720 9.640 188.040 9.960 ;
        RECT 188.120 9.640 188.440 9.960 ;
        RECT 188.520 9.640 188.840 9.960 ;
        RECT 188.920 9.640 189.240 9.960 ;
        RECT 189.320 9.640 189.640 9.960 ;
        RECT 189.720 9.640 190.040 9.960 ;
        RECT 190.120 9.640 190.440 9.960 ;
        RECT 190.520 9.640 190.840 9.960 ;
        RECT 190.920 9.640 191.240 9.960 ;
        RECT 191.320 9.640 191.640 9.960 ;
        RECT 191.720 9.640 192.040 9.960 ;
        RECT 192.120 9.640 192.440 9.960 ;
        RECT 192.520 9.640 192.840 9.960 ;
        RECT 192.920 9.640 193.240 9.960 ;
        RECT 193.320 9.640 193.640 9.960 ;
        RECT 193.720 9.640 194.040 9.960 ;
        RECT 194.120 9.640 194.440 9.960 ;
        RECT 194.520 9.640 194.840 9.960 ;
        RECT 194.920 9.640 195.240 9.960 ;
        RECT 195.320 9.640 195.640 9.960 ;
        RECT 195.720 9.640 196.040 9.960 ;
        RECT 196.120 9.640 196.440 9.960 ;
        RECT 196.520 9.640 196.840 9.960 ;
        RECT 196.920 9.640 197.240 9.960 ;
        RECT 197.320 9.640 197.640 9.960 ;
        RECT 197.720 9.640 198.040 9.960 ;
        RECT 198.120 9.640 198.440 9.960 ;
        RECT 198.520 9.640 198.840 9.960 ;
        RECT 198.920 9.640 199.240 9.960 ;
        RECT 199.320 9.640 199.640 9.960 ;
        RECT 199.720 9.640 200.040 9.960 ;
        RECT 200.120 9.640 200.440 9.960 ;
        RECT 200.520 9.640 200.840 9.960 ;
        RECT 200.920 9.640 201.240 9.960 ;
        RECT 201.320 9.640 201.640 9.960 ;
        RECT 201.720 9.640 202.040 9.960 ;
        RECT 202.120 9.640 202.440 9.960 ;
        RECT 202.520 9.640 202.840 9.960 ;
        RECT 202.920 9.640 203.240 9.960 ;
        RECT 203.320 9.640 203.640 9.960 ;
        RECT 203.720 9.640 204.040 9.960 ;
        RECT 204.120 9.640 204.440 9.960 ;
        RECT 204.520 9.640 204.840 9.960 ;
        RECT 204.920 9.640 205.240 9.960 ;
        RECT 205.320 9.640 205.640 9.960 ;
        RECT 0.040 9.240 0.360 9.560 ;
        RECT 0.440 9.240 0.760 9.560 ;
        RECT 0.840 9.240 1.160 9.560 ;
        RECT 1.240 9.240 1.560 9.560 ;
        RECT 1.640 9.240 1.960 9.560 ;
        RECT 2.040 9.240 2.360 9.560 ;
        RECT 2.440 9.240 2.760 9.560 ;
        RECT 2.840 9.240 3.160 9.560 ;
        RECT 3.240 9.240 3.560 9.560 ;
        RECT 3.640 9.240 3.960 9.560 ;
        RECT 4.040 9.240 4.360 9.560 ;
        RECT 4.440 9.240 4.760 9.560 ;
        RECT 4.840 9.240 5.160 9.560 ;
        RECT 5.240 9.240 5.560 9.560 ;
        RECT 5.640 9.240 5.960 9.560 ;
        RECT 6.040 9.240 6.360 9.560 ;
        RECT 6.440 9.240 6.760 9.560 ;
        RECT 6.840 9.240 7.160 9.560 ;
        RECT 7.240 9.240 7.560 9.560 ;
        RECT 7.640 9.240 7.960 9.560 ;
        RECT 8.040 9.240 8.360 9.560 ;
        RECT 8.440 9.240 8.760 9.560 ;
        RECT 8.840 9.240 9.160 9.560 ;
        RECT 9.240 9.240 9.560 9.560 ;
        RECT 9.640 9.240 9.960 9.560 ;
        RECT 10.040 9.240 10.360 9.560 ;
        RECT 10.440 9.240 10.760 9.560 ;
        RECT 10.840 9.240 11.160 9.560 ;
        RECT 11.240 9.240 11.560 9.560 ;
        RECT 11.640 9.240 11.960 9.560 ;
        RECT 12.040 9.240 12.360 9.560 ;
        RECT 12.440 9.240 12.760 9.560 ;
        RECT 12.840 9.240 13.160 9.560 ;
        RECT 13.240 9.240 13.560 9.560 ;
        RECT 13.640 9.240 13.960 9.560 ;
        RECT 14.040 9.240 14.360 9.560 ;
        RECT 14.440 9.240 14.760 9.560 ;
        RECT 14.840 9.240 15.160 9.560 ;
        RECT 15.240 9.240 15.560 9.560 ;
        RECT 15.640 9.240 15.960 9.560 ;
        RECT 16.040 9.240 16.360 9.560 ;
        RECT 16.440 9.240 16.760 9.560 ;
        RECT 16.840 9.240 17.160 9.560 ;
        RECT 17.240 9.240 17.560 9.560 ;
        RECT 17.640 9.240 17.960 9.560 ;
        RECT 18.040 9.240 18.360 9.560 ;
        RECT 18.440 9.240 18.760 9.560 ;
        RECT 18.840 9.240 19.160 9.560 ;
        RECT 19.240 9.240 19.560 9.560 ;
        RECT 19.640 9.240 19.960 9.560 ;
        RECT 95.560 9.240 95.880 9.560 ;
        RECT 95.960 9.240 96.280 9.560 ;
        RECT 96.360 9.240 96.680 9.560 ;
        RECT 96.760 9.240 97.080 9.560 ;
        RECT 145.560 9.240 145.880 9.560 ;
        RECT 145.960 9.240 146.280 9.560 ;
        RECT 146.360 9.240 146.680 9.560 ;
        RECT 146.760 9.240 147.080 9.560 ;
        RECT 185.720 9.240 186.040 9.560 ;
        RECT 186.120 9.240 186.440 9.560 ;
        RECT 186.520 9.240 186.840 9.560 ;
        RECT 186.920 9.240 187.240 9.560 ;
        RECT 187.320 9.240 187.640 9.560 ;
        RECT 187.720 9.240 188.040 9.560 ;
        RECT 188.120 9.240 188.440 9.560 ;
        RECT 188.520 9.240 188.840 9.560 ;
        RECT 188.920 9.240 189.240 9.560 ;
        RECT 189.320 9.240 189.640 9.560 ;
        RECT 189.720 9.240 190.040 9.560 ;
        RECT 190.120 9.240 190.440 9.560 ;
        RECT 190.520 9.240 190.840 9.560 ;
        RECT 190.920 9.240 191.240 9.560 ;
        RECT 191.320 9.240 191.640 9.560 ;
        RECT 191.720 9.240 192.040 9.560 ;
        RECT 192.120 9.240 192.440 9.560 ;
        RECT 192.520 9.240 192.840 9.560 ;
        RECT 192.920 9.240 193.240 9.560 ;
        RECT 193.320 9.240 193.640 9.560 ;
        RECT 193.720 9.240 194.040 9.560 ;
        RECT 194.120 9.240 194.440 9.560 ;
        RECT 194.520 9.240 194.840 9.560 ;
        RECT 194.920 9.240 195.240 9.560 ;
        RECT 195.320 9.240 195.640 9.560 ;
        RECT 195.720 9.240 196.040 9.560 ;
        RECT 196.120 9.240 196.440 9.560 ;
        RECT 196.520 9.240 196.840 9.560 ;
        RECT 196.920 9.240 197.240 9.560 ;
        RECT 197.320 9.240 197.640 9.560 ;
        RECT 197.720 9.240 198.040 9.560 ;
        RECT 198.120 9.240 198.440 9.560 ;
        RECT 198.520 9.240 198.840 9.560 ;
        RECT 198.920 9.240 199.240 9.560 ;
        RECT 199.320 9.240 199.640 9.560 ;
        RECT 199.720 9.240 200.040 9.560 ;
        RECT 200.120 9.240 200.440 9.560 ;
        RECT 200.520 9.240 200.840 9.560 ;
        RECT 200.920 9.240 201.240 9.560 ;
        RECT 201.320 9.240 201.640 9.560 ;
        RECT 201.720 9.240 202.040 9.560 ;
        RECT 202.120 9.240 202.440 9.560 ;
        RECT 202.520 9.240 202.840 9.560 ;
        RECT 202.920 9.240 203.240 9.560 ;
        RECT 203.320 9.240 203.640 9.560 ;
        RECT 203.720 9.240 204.040 9.560 ;
        RECT 204.120 9.240 204.440 9.560 ;
        RECT 204.520 9.240 204.840 9.560 ;
        RECT 204.920 9.240 205.240 9.560 ;
        RECT 205.320 9.240 205.640 9.560 ;
        RECT 0.040 8.840 0.360 9.160 ;
        RECT 0.440 8.840 0.760 9.160 ;
        RECT 0.840 8.840 1.160 9.160 ;
        RECT 1.240 8.840 1.560 9.160 ;
        RECT 1.640 8.840 1.960 9.160 ;
        RECT 2.040 8.840 2.360 9.160 ;
        RECT 2.440 8.840 2.760 9.160 ;
        RECT 2.840 8.840 3.160 9.160 ;
        RECT 3.240 8.840 3.560 9.160 ;
        RECT 3.640 8.840 3.960 9.160 ;
        RECT 4.040 8.840 4.360 9.160 ;
        RECT 4.440 8.840 4.760 9.160 ;
        RECT 4.840 8.840 5.160 9.160 ;
        RECT 5.240 8.840 5.560 9.160 ;
        RECT 5.640 8.840 5.960 9.160 ;
        RECT 6.040 8.840 6.360 9.160 ;
        RECT 6.440 8.840 6.760 9.160 ;
        RECT 6.840 8.840 7.160 9.160 ;
        RECT 7.240 8.840 7.560 9.160 ;
        RECT 7.640 8.840 7.960 9.160 ;
        RECT 8.040 8.840 8.360 9.160 ;
        RECT 8.440 8.840 8.760 9.160 ;
        RECT 8.840 8.840 9.160 9.160 ;
        RECT 9.240 8.840 9.560 9.160 ;
        RECT 9.640 8.840 9.960 9.160 ;
        RECT 10.040 8.840 10.360 9.160 ;
        RECT 10.440 8.840 10.760 9.160 ;
        RECT 10.840 8.840 11.160 9.160 ;
        RECT 11.240 8.840 11.560 9.160 ;
        RECT 11.640 8.840 11.960 9.160 ;
        RECT 12.040 8.840 12.360 9.160 ;
        RECT 12.440 8.840 12.760 9.160 ;
        RECT 12.840 8.840 13.160 9.160 ;
        RECT 13.240 8.840 13.560 9.160 ;
        RECT 13.640 8.840 13.960 9.160 ;
        RECT 14.040 8.840 14.360 9.160 ;
        RECT 14.440 8.840 14.760 9.160 ;
        RECT 14.840 8.840 15.160 9.160 ;
        RECT 15.240 8.840 15.560 9.160 ;
        RECT 15.640 8.840 15.960 9.160 ;
        RECT 16.040 8.840 16.360 9.160 ;
        RECT 16.440 8.840 16.760 9.160 ;
        RECT 16.840 8.840 17.160 9.160 ;
        RECT 17.240 8.840 17.560 9.160 ;
        RECT 17.640 8.840 17.960 9.160 ;
        RECT 18.040 8.840 18.360 9.160 ;
        RECT 18.440 8.840 18.760 9.160 ;
        RECT 18.840 8.840 19.160 9.160 ;
        RECT 19.240 8.840 19.560 9.160 ;
        RECT 19.640 8.840 19.960 9.160 ;
        RECT 95.560 8.840 95.880 9.160 ;
        RECT 95.960 8.840 96.280 9.160 ;
        RECT 96.360 8.840 96.680 9.160 ;
        RECT 96.760 8.840 97.080 9.160 ;
        RECT 145.560 8.840 145.880 9.160 ;
        RECT 145.960 8.840 146.280 9.160 ;
        RECT 146.360 8.840 146.680 9.160 ;
        RECT 146.760 8.840 147.080 9.160 ;
        RECT 185.720 8.840 186.040 9.160 ;
        RECT 186.120 8.840 186.440 9.160 ;
        RECT 186.520 8.840 186.840 9.160 ;
        RECT 186.920 8.840 187.240 9.160 ;
        RECT 187.320 8.840 187.640 9.160 ;
        RECT 187.720 8.840 188.040 9.160 ;
        RECT 188.120 8.840 188.440 9.160 ;
        RECT 188.520 8.840 188.840 9.160 ;
        RECT 188.920 8.840 189.240 9.160 ;
        RECT 189.320 8.840 189.640 9.160 ;
        RECT 189.720 8.840 190.040 9.160 ;
        RECT 190.120 8.840 190.440 9.160 ;
        RECT 190.520 8.840 190.840 9.160 ;
        RECT 190.920 8.840 191.240 9.160 ;
        RECT 191.320 8.840 191.640 9.160 ;
        RECT 191.720 8.840 192.040 9.160 ;
        RECT 192.120 8.840 192.440 9.160 ;
        RECT 192.520 8.840 192.840 9.160 ;
        RECT 192.920 8.840 193.240 9.160 ;
        RECT 193.320 8.840 193.640 9.160 ;
        RECT 193.720 8.840 194.040 9.160 ;
        RECT 194.120 8.840 194.440 9.160 ;
        RECT 194.520 8.840 194.840 9.160 ;
        RECT 194.920 8.840 195.240 9.160 ;
        RECT 195.320 8.840 195.640 9.160 ;
        RECT 195.720 8.840 196.040 9.160 ;
        RECT 196.120 8.840 196.440 9.160 ;
        RECT 196.520 8.840 196.840 9.160 ;
        RECT 196.920 8.840 197.240 9.160 ;
        RECT 197.320 8.840 197.640 9.160 ;
        RECT 197.720 8.840 198.040 9.160 ;
        RECT 198.120 8.840 198.440 9.160 ;
        RECT 198.520 8.840 198.840 9.160 ;
        RECT 198.920 8.840 199.240 9.160 ;
        RECT 199.320 8.840 199.640 9.160 ;
        RECT 199.720 8.840 200.040 9.160 ;
        RECT 200.120 8.840 200.440 9.160 ;
        RECT 200.520 8.840 200.840 9.160 ;
        RECT 200.920 8.840 201.240 9.160 ;
        RECT 201.320 8.840 201.640 9.160 ;
        RECT 201.720 8.840 202.040 9.160 ;
        RECT 202.120 8.840 202.440 9.160 ;
        RECT 202.520 8.840 202.840 9.160 ;
        RECT 202.920 8.840 203.240 9.160 ;
        RECT 203.320 8.840 203.640 9.160 ;
        RECT 203.720 8.840 204.040 9.160 ;
        RECT 204.120 8.840 204.440 9.160 ;
        RECT 204.520 8.840 204.840 9.160 ;
        RECT 204.920 8.840 205.240 9.160 ;
        RECT 205.320 8.840 205.640 9.160 ;
        RECT 0.040 8.440 0.360 8.760 ;
        RECT 0.440 8.440 0.760 8.760 ;
        RECT 0.840 8.440 1.160 8.760 ;
        RECT 1.240 8.440 1.560 8.760 ;
        RECT 1.640 8.440 1.960 8.760 ;
        RECT 2.040 8.440 2.360 8.760 ;
        RECT 2.440 8.440 2.760 8.760 ;
        RECT 2.840 8.440 3.160 8.760 ;
        RECT 3.240 8.440 3.560 8.760 ;
        RECT 3.640 8.440 3.960 8.760 ;
        RECT 4.040 8.440 4.360 8.760 ;
        RECT 4.440 8.440 4.760 8.760 ;
        RECT 4.840 8.440 5.160 8.760 ;
        RECT 5.240 8.440 5.560 8.760 ;
        RECT 5.640 8.440 5.960 8.760 ;
        RECT 6.040 8.440 6.360 8.760 ;
        RECT 6.440 8.440 6.760 8.760 ;
        RECT 6.840 8.440 7.160 8.760 ;
        RECT 7.240 8.440 7.560 8.760 ;
        RECT 7.640 8.440 7.960 8.760 ;
        RECT 8.040 8.440 8.360 8.760 ;
        RECT 8.440 8.440 8.760 8.760 ;
        RECT 8.840 8.440 9.160 8.760 ;
        RECT 9.240 8.440 9.560 8.760 ;
        RECT 9.640 8.440 9.960 8.760 ;
        RECT 10.040 8.440 10.360 8.760 ;
        RECT 10.440 8.440 10.760 8.760 ;
        RECT 10.840 8.440 11.160 8.760 ;
        RECT 11.240 8.440 11.560 8.760 ;
        RECT 11.640 8.440 11.960 8.760 ;
        RECT 12.040 8.440 12.360 8.760 ;
        RECT 12.440 8.440 12.760 8.760 ;
        RECT 12.840 8.440 13.160 8.760 ;
        RECT 13.240 8.440 13.560 8.760 ;
        RECT 13.640 8.440 13.960 8.760 ;
        RECT 14.040 8.440 14.360 8.760 ;
        RECT 14.440 8.440 14.760 8.760 ;
        RECT 14.840 8.440 15.160 8.760 ;
        RECT 15.240 8.440 15.560 8.760 ;
        RECT 15.640 8.440 15.960 8.760 ;
        RECT 16.040 8.440 16.360 8.760 ;
        RECT 16.440 8.440 16.760 8.760 ;
        RECT 16.840 8.440 17.160 8.760 ;
        RECT 17.240 8.440 17.560 8.760 ;
        RECT 17.640 8.440 17.960 8.760 ;
        RECT 18.040 8.440 18.360 8.760 ;
        RECT 18.440 8.440 18.760 8.760 ;
        RECT 18.840 8.440 19.160 8.760 ;
        RECT 19.240 8.440 19.560 8.760 ;
        RECT 19.640 8.440 19.960 8.760 ;
        RECT 95.560 8.440 95.880 8.760 ;
        RECT 95.960 8.440 96.280 8.760 ;
        RECT 96.360 8.440 96.680 8.760 ;
        RECT 96.760 8.440 97.080 8.760 ;
        RECT 145.560 8.440 145.880 8.760 ;
        RECT 145.960 8.440 146.280 8.760 ;
        RECT 146.360 8.440 146.680 8.760 ;
        RECT 146.760 8.440 147.080 8.760 ;
        RECT 185.720 8.440 186.040 8.760 ;
        RECT 186.120 8.440 186.440 8.760 ;
        RECT 186.520 8.440 186.840 8.760 ;
        RECT 186.920 8.440 187.240 8.760 ;
        RECT 187.320 8.440 187.640 8.760 ;
        RECT 187.720 8.440 188.040 8.760 ;
        RECT 188.120 8.440 188.440 8.760 ;
        RECT 188.520 8.440 188.840 8.760 ;
        RECT 188.920 8.440 189.240 8.760 ;
        RECT 189.320 8.440 189.640 8.760 ;
        RECT 189.720 8.440 190.040 8.760 ;
        RECT 190.120 8.440 190.440 8.760 ;
        RECT 190.520 8.440 190.840 8.760 ;
        RECT 190.920 8.440 191.240 8.760 ;
        RECT 191.320 8.440 191.640 8.760 ;
        RECT 191.720 8.440 192.040 8.760 ;
        RECT 192.120 8.440 192.440 8.760 ;
        RECT 192.520 8.440 192.840 8.760 ;
        RECT 192.920 8.440 193.240 8.760 ;
        RECT 193.320 8.440 193.640 8.760 ;
        RECT 193.720 8.440 194.040 8.760 ;
        RECT 194.120 8.440 194.440 8.760 ;
        RECT 194.520 8.440 194.840 8.760 ;
        RECT 194.920 8.440 195.240 8.760 ;
        RECT 195.320 8.440 195.640 8.760 ;
        RECT 195.720 8.440 196.040 8.760 ;
        RECT 196.120 8.440 196.440 8.760 ;
        RECT 196.520 8.440 196.840 8.760 ;
        RECT 196.920 8.440 197.240 8.760 ;
        RECT 197.320 8.440 197.640 8.760 ;
        RECT 197.720 8.440 198.040 8.760 ;
        RECT 198.120 8.440 198.440 8.760 ;
        RECT 198.520 8.440 198.840 8.760 ;
        RECT 198.920 8.440 199.240 8.760 ;
        RECT 199.320 8.440 199.640 8.760 ;
        RECT 199.720 8.440 200.040 8.760 ;
        RECT 200.120 8.440 200.440 8.760 ;
        RECT 200.520 8.440 200.840 8.760 ;
        RECT 200.920 8.440 201.240 8.760 ;
        RECT 201.320 8.440 201.640 8.760 ;
        RECT 201.720 8.440 202.040 8.760 ;
        RECT 202.120 8.440 202.440 8.760 ;
        RECT 202.520 8.440 202.840 8.760 ;
        RECT 202.920 8.440 203.240 8.760 ;
        RECT 203.320 8.440 203.640 8.760 ;
        RECT 203.720 8.440 204.040 8.760 ;
        RECT 204.120 8.440 204.440 8.760 ;
        RECT 204.520 8.440 204.840 8.760 ;
        RECT 204.920 8.440 205.240 8.760 ;
        RECT 205.320 8.440 205.640 8.760 ;
        RECT 0.040 8.040 0.360 8.360 ;
        RECT 0.440 8.040 0.760 8.360 ;
        RECT 0.840 8.040 1.160 8.360 ;
        RECT 1.240 8.040 1.560 8.360 ;
        RECT 1.640 8.040 1.960 8.360 ;
        RECT 2.040 8.040 2.360 8.360 ;
        RECT 2.440 8.040 2.760 8.360 ;
        RECT 2.840 8.040 3.160 8.360 ;
        RECT 3.240 8.040 3.560 8.360 ;
        RECT 3.640 8.040 3.960 8.360 ;
        RECT 4.040 8.040 4.360 8.360 ;
        RECT 4.440 8.040 4.760 8.360 ;
        RECT 4.840 8.040 5.160 8.360 ;
        RECT 5.240 8.040 5.560 8.360 ;
        RECT 5.640 8.040 5.960 8.360 ;
        RECT 6.040 8.040 6.360 8.360 ;
        RECT 6.440 8.040 6.760 8.360 ;
        RECT 6.840 8.040 7.160 8.360 ;
        RECT 7.240 8.040 7.560 8.360 ;
        RECT 7.640 8.040 7.960 8.360 ;
        RECT 8.040 8.040 8.360 8.360 ;
        RECT 8.440 8.040 8.760 8.360 ;
        RECT 8.840 8.040 9.160 8.360 ;
        RECT 9.240 8.040 9.560 8.360 ;
        RECT 9.640 8.040 9.960 8.360 ;
        RECT 10.040 8.040 10.360 8.360 ;
        RECT 10.440 8.040 10.760 8.360 ;
        RECT 10.840 8.040 11.160 8.360 ;
        RECT 11.240 8.040 11.560 8.360 ;
        RECT 11.640 8.040 11.960 8.360 ;
        RECT 12.040 8.040 12.360 8.360 ;
        RECT 12.440 8.040 12.760 8.360 ;
        RECT 12.840 8.040 13.160 8.360 ;
        RECT 13.240 8.040 13.560 8.360 ;
        RECT 13.640 8.040 13.960 8.360 ;
        RECT 14.040 8.040 14.360 8.360 ;
        RECT 14.440 8.040 14.760 8.360 ;
        RECT 14.840 8.040 15.160 8.360 ;
        RECT 15.240 8.040 15.560 8.360 ;
        RECT 15.640 8.040 15.960 8.360 ;
        RECT 16.040 8.040 16.360 8.360 ;
        RECT 16.440 8.040 16.760 8.360 ;
        RECT 16.840 8.040 17.160 8.360 ;
        RECT 17.240 8.040 17.560 8.360 ;
        RECT 17.640 8.040 17.960 8.360 ;
        RECT 18.040 8.040 18.360 8.360 ;
        RECT 18.440 8.040 18.760 8.360 ;
        RECT 18.840 8.040 19.160 8.360 ;
        RECT 19.240 8.040 19.560 8.360 ;
        RECT 19.640 8.040 19.960 8.360 ;
        RECT 95.560 8.040 95.880 8.360 ;
        RECT 95.960 8.040 96.280 8.360 ;
        RECT 96.360 8.040 96.680 8.360 ;
        RECT 96.760 8.040 97.080 8.360 ;
        RECT 145.560 8.040 145.880 8.360 ;
        RECT 145.960 8.040 146.280 8.360 ;
        RECT 146.360 8.040 146.680 8.360 ;
        RECT 146.760 8.040 147.080 8.360 ;
        RECT 185.720 8.040 186.040 8.360 ;
        RECT 186.120 8.040 186.440 8.360 ;
        RECT 186.520 8.040 186.840 8.360 ;
        RECT 186.920 8.040 187.240 8.360 ;
        RECT 187.320 8.040 187.640 8.360 ;
        RECT 187.720 8.040 188.040 8.360 ;
        RECT 188.120 8.040 188.440 8.360 ;
        RECT 188.520 8.040 188.840 8.360 ;
        RECT 188.920 8.040 189.240 8.360 ;
        RECT 189.320 8.040 189.640 8.360 ;
        RECT 189.720 8.040 190.040 8.360 ;
        RECT 190.120 8.040 190.440 8.360 ;
        RECT 190.520 8.040 190.840 8.360 ;
        RECT 190.920 8.040 191.240 8.360 ;
        RECT 191.320 8.040 191.640 8.360 ;
        RECT 191.720 8.040 192.040 8.360 ;
        RECT 192.120 8.040 192.440 8.360 ;
        RECT 192.520 8.040 192.840 8.360 ;
        RECT 192.920 8.040 193.240 8.360 ;
        RECT 193.320 8.040 193.640 8.360 ;
        RECT 193.720 8.040 194.040 8.360 ;
        RECT 194.120 8.040 194.440 8.360 ;
        RECT 194.520 8.040 194.840 8.360 ;
        RECT 194.920 8.040 195.240 8.360 ;
        RECT 195.320 8.040 195.640 8.360 ;
        RECT 195.720 8.040 196.040 8.360 ;
        RECT 196.120 8.040 196.440 8.360 ;
        RECT 196.520 8.040 196.840 8.360 ;
        RECT 196.920 8.040 197.240 8.360 ;
        RECT 197.320 8.040 197.640 8.360 ;
        RECT 197.720 8.040 198.040 8.360 ;
        RECT 198.120 8.040 198.440 8.360 ;
        RECT 198.520 8.040 198.840 8.360 ;
        RECT 198.920 8.040 199.240 8.360 ;
        RECT 199.320 8.040 199.640 8.360 ;
        RECT 199.720 8.040 200.040 8.360 ;
        RECT 200.120 8.040 200.440 8.360 ;
        RECT 200.520 8.040 200.840 8.360 ;
        RECT 200.920 8.040 201.240 8.360 ;
        RECT 201.320 8.040 201.640 8.360 ;
        RECT 201.720 8.040 202.040 8.360 ;
        RECT 202.120 8.040 202.440 8.360 ;
        RECT 202.520 8.040 202.840 8.360 ;
        RECT 202.920 8.040 203.240 8.360 ;
        RECT 203.320 8.040 203.640 8.360 ;
        RECT 203.720 8.040 204.040 8.360 ;
        RECT 204.120 8.040 204.440 8.360 ;
        RECT 204.520 8.040 204.840 8.360 ;
        RECT 204.920 8.040 205.240 8.360 ;
        RECT 205.320 8.040 205.640 8.360 ;
        RECT 0.040 7.640 0.360 7.960 ;
        RECT 0.440 7.640 0.760 7.960 ;
        RECT 0.840 7.640 1.160 7.960 ;
        RECT 1.240 7.640 1.560 7.960 ;
        RECT 1.640 7.640 1.960 7.960 ;
        RECT 2.040 7.640 2.360 7.960 ;
        RECT 2.440 7.640 2.760 7.960 ;
        RECT 2.840 7.640 3.160 7.960 ;
        RECT 3.240 7.640 3.560 7.960 ;
        RECT 3.640 7.640 3.960 7.960 ;
        RECT 4.040 7.640 4.360 7.960 ;
        RECT 4.440 7.640 4.760 7.960 ;
        RECT 4.840 7.640 5.160 7.960 ;
        RECT 5.240 7.640 5.560 7.960 ;
        RECT 5.640 7.640 5.960 7.960 ;
        RECT 6.040 7.640 6.360 7.960 ;
        RECT 6.440 7.640 6.760 7.960 ;
        RECT 6.840 7.640 7.160 7.960 ;
        RECT 7.240 7.640 7.560 7.960 ;
        RECT 7.640 7.640 7.960 7.960 ;
        RECT 8.040 7.640 8.360 7.960 ;
        RECT 8.440 7.640 8.760 7.960 ;
        RECT 8.840 7.640 9.160 7.960 ;
        RECT 9.240 7.640 9.560 7.960 ;
        RECT 9.640 7.640 9.960 7.960 ;
        RECT 10.040 7.640 10.360 7.960 ;
        RECT 10.440 7.640 10.760 7.960 ;
        RECT 10.840 7.640 11.160 7.960 ;
        RECT 11.240 7.640 11.560 7.960 ;
        RECT 11.640 7.640 11.960 7.960 ;
        RECT 12.040 7.640 12.360 7.960 ;
        RECT 12.440 7.640 12.760 7.960 ;
        RECT 12.840 7.640 13.160 7.960 ;
        RECT 13.240 7.640 13.560 7.960 ;
        RECT 13.640 7.640 13.960 7.960 ;
        RECT 14.040 7.640 14.360 7.960 ;
        RECT 14.440 7.640 14.760 7.960 ;
        RECT 14.840 7.640 15.160 7.960 ;
        RECT 15.240 7.640 15.560 7.960 ;
        RECT 15.640 7.640 15.960 7.960 ;
        RECT 16.040 7.640 16.360 7.960 ;
        RECT 16.440 7.640 16.760 7.960 ;
        RECT 16.840 7.640 17.160 7.960 ;
        RECT 17.240 7.640 17.560 7.960 ;
        RECT 17.640 7.640 17.960 7.960 ;
        RECT 18.040 7.640 18.360 7.960 ;
        RECT 18.440 7.640 18.760 7.960 ;
        RECT 18.840 7.640 19.160 7.960 ;
        RECT 19.240 7.640 19.560 7.960 ;
        RECT 19.640 7.640 19.960 7.960 ;
        RECT 95.560 7.640 95.880 7.960 ;
        RECT 95.960 7.640 96.280 7.960 ;
        RECT 96.360 7.640 96.680 7.960 ;
        RECT 96.760 7.640 97.080 7.960 ;
        RECT 145.560 7.640 145.880 7.960 ;
        RECT 145.960 7.640 146.280 7.960 ;
        RECT 146.360 7.640 146.680 7.960 ;
        RECT 146.760 7.640 147.080 7.960 ;
        RECT 185.720 7.640 186.040 7.960 ;
        RECT 186.120 7.640 186.440 7.960 ;
        RECT 186.520 7.640 186.840 7.960 ;
        RECT 186.920 7.640 187.240 7.960 ;
        RECT 187.320 7.640 187.640 7.960 ;
        RECT 187.720 7.640 188.040 7.960 ;
        RECT 188.120 7.640 188.440 7.960 ;
        RECT 188.520 7.640 188.840 7.960 ;
        RECT 188.920 7.640 189.240 7.960 ;
        RECT 189.320 7.640 189.640 7.960 ;
        RECT 189.720 7.640 190.040 7.960 ;
        RECT 190.120 7.640 190.440 7.960 ;
        RECT 190.520 7.640 190.840 7.960 ;
        RECT 190.920 7.640 191.240 7.960 ;
        RECT 191.320 7.640 191.640 7.960 ;
        RECT 191.720 7.640 192.040 7.960 ;
        RECT 192.120 7.640 192.440 7.960 ;
        RECT 192.520 7.640 192.840 7.960 ;
        RECT 192.920 7.640 193.240 7.960 ;
        RECT 193.320 7.640 193.640 7.960 ;
        RECT 193.720 7.640 194.040 7.960 ;
        RECT 194.120 7.640 194.440 7.960 ;
        RECT 194.520 7.640 194.840 7.960 ;
        RECT 194.920 7.640 195.240 7.960 ;
        RECT 195.320 7.640 195.640 7.960 ;
        RECT 195.720 7.640 196.040 7.960 ;
        RECT 196.120 7.640 196.440 7.960 ;
        RECT 196.520 7.640 196.840 7.960 ;
        RECT 196.920 7.640 197.240 7.960 ;
        RECT 197.320 7.640 197.640 7.960 ;
        RECT 197.720 7.640 198.040 7.960 ;
        RECT 198.120 7.640 198.440 7.960 ;
        RECT 198.520 7.640 198.840 7.960 ;
        RECT 198.920 7.640 199.240 7.960 ;
        RECT 199.320 7.640 199.640 7.960 ;
        RECT 199.720 7.640 200.040 7.960 ;
        RECT 200.120 7.640 200.440 7.960 ;
        RECT 200.520 7.640 200.840 7.960 ;
        RECT 200.920 7.640 201.240 7.960 ;
        RECT 201.320 7.640 201.640 7.960 ;
        RECT 201.720 7.640 202.040 7.960 ;
        RECT 202.120 7.640 202.440 7.960 ;
        RECT 202.520 7.640 202.840 7.960 ;
        RECT 202.920 7.640 203.240 7.960 ;
        RECT 203.320 7.640 203.640 7.960 ;
        RECT 203.720 7.640 204.040 7.960 ;
        RECT 204.120 7.640 204.440 7.960 ;
        RECT 204.520 7.640 204.840 7.960 ;
        RECT 204.920 7.640 205.240 7.960 ;
        RECT 205.320 7.640 205.640 7.960 ;
        RECT 0.040 7.240 0.360 7.560 ;
        RECT 0.440 7.240 0.760 7.560 ;
        RECT 0.840 7.240 1.160 7.560 ;
        RECT 1.240 7.240 1.560 7.560 ;
        RECT 1.640 7.240 1.960 7.560 ;
        RECT 2.040 7.240 2.360 7.560 ;
        RECT 2.440 7.240 2.760 7.560 ;
        RECT 2.840 7.240 3.160 7.560 ;
        RECT 3.240 7.240 3.560 7.560 ;
        RECT 3.640 7.240 3.960 7.560 ;
        RECT 4.040 7.240 4.360 7.560 ;
        RECT 4.440 7.240 4.760 7.560 ;
        RECT 4.840 7.240 5.160 7.560 ;
        RECT 5.240 7.240 5.560 7.560 ;
        RECT 5.640 7.240 5.960 7.560 ;
        RECT 6.040 7.240 6.360 7.560 ;
        RECT 6.440 7.240 6.760 7.560 ;
        RECT 6.840 7.240 7.160 7.560 ;
        RECT 7.240 7.240 7.560 7.560 ;
        RECT 7.640 7.240 7.960 7.560 ;
        RECT 8.040 7.240 8.360 7.560 ;
        RECT 8.440 7.240 8.760 7.560 ;
        RECT 8.840 7.240 9.160 7.560 ;
        RECT 9.240 7.240 9.560 7.560 ;
        RECT 9.640 7.240 9.960 7.560 ;
        RECT 10.040 7.240 10.360 7.560 ;
        RECT 10.440 7.240 10.760 7.560 ;
        RECT 10.840 7.240 11.160 7.560 ;
        RECT 11.240 7.240 11.560 7.560 ;
        RECT 11.640 7.240 11.960 7.560 ;
        RECT 12.040 7.240 12.360 7.560 ;
        RECT 12.440 7.240 12.760 7.560 ;
        RECT 12.840 7.240 13.160 7.560 ;
        RECT 13.240 7.240 13.560 7.560 ;
        RECT 13.640 7.240 13.960 7.560 ;
        RECT 14.040 7.240 14.360 7.560 ;
        RECT 14.440 7.240 14.760 7.560 ;
        RECT 14.840 7.240 15.160 7.560 ;
        RECT 15.240 7.240 15.560 7.560 ;
        RECT 15.640 7.240 15.960 7.560 ;
        RECT 16.040 7.240 16.360 7.560 ;
        RECT 16.440 7.240 16.760 7.560 ;
        RECT 16.840 7.240 17.160 7.560 ;
        RECT 17.240 7.240 17.560 7.560 ;
        RECT 17.640 7.240 17.960 7.560 ;
        RECT 18.040 7.240 18.360 7.560 ;
        RECT 18.440 7.240 18.760 7.560 ;
        RECT 18.840 7.240 19.160 7.560 ;
        RECT 19.240 7.240 19.560 7.560 ;
        RECT 19.640 7.240 19.960 7.560 ;
        RECT 95.560 7.240 95.880 7.560 ;
        RECT 95.960 7.240 96.280 7.560 ;
        RECT 96.360 7.240 96.680 7.560 ;
        RECT 96.760 7.240 97.080 7.560 ;
        RECT 145.560 7.240 145.880 7.560 ;
        RECT 145.960 7.240 146.280 7.560 ;
        RECT 146.360 7.240 146.680 7.560 ;
        RECT 146.760 7.240 147.080 7.560 ;
        RECT 185.720 7.240 186.040 7.560 ;
        RECT 186.120 7.240 186.440 7.560 ;
        RECT 186.520 7.240 186.840 7.560 ;
        RECT 186.920 7.240 187.240 7.560 ;
        RECT 187.320 7.240 187.640 7.560 ;
        RECT 187.720 7.240 188.040 7.560 ;
        RECT 188.120 7.240 188.440 7.560 ;
        RECT 188.520 7.240 188.840 7.560 ;
        RECT 188.920 7.240 189.240 7.560 ;
        RECT 189.320 7.240 189.640 7.560 ;
        RECT 189.720 7.240 190.040 7.560 ;
        RECT 190.120 7.240 190.440 7.560 ;
        RECT 190.520 7.240 190.840 7.560 ;
        RECT 190.920 7.240 191.240 7.560 ;
        RECT 191.320 7.240 191.640 7.560 ;
        RECT 191.720 7.240 192.040 7.560 ;
        RECT 192.120 7.240 192.440 7.560 ;
        RECT 192.520 7.240 192.840 7.560 ;
        RECT 192.920 7.240 193.240 7.560 ;
        RECT 193.320 7.240 193.640 7.560 ;
        RECT 193.720 7.240 194.040 7.560 ;
        RECT 194.120 7.240 194.440 7.560 ;
        RECT 194.520 7.240 194.840 7.560 ;
        RECT 194.920 7.240 195.240 7.560 ;
        RECT 195.320 7.240 195.640 7.560 ;
        RECT 195.720 7.240 196.040 7.560 ;
        RECT 196.120 7.240 196.440 7.560 ;
        RECT 196.520 7.240 196.840 7.560 ;
        RECT 196.920 7.240 197.240 7.560 ;
        RECT 197.320 7.240 197.640 7.560 ;
        RECT 197.720 7.240 198.040 7.560 ;
        RECT 198.120 7.240 198.440 7.560 ;
        RECT 198.520 7.240 198.840 7.560 ;
        RECT 198.920 7.240 199.240 7.560 ;
        RECT 199.320 7.240 199.640 7.560 ;
        RECT 199.720 7.240 200.040 7.560 ;
        RECT 200.120 7.240 200.440 7.560 ;
        RECT 200.520 7.240 200.840 7.560 ;
        RECT 200.920 7.240 201.240 7.560 ;
        RECT 201.320 7.240 201.640 7.560 ;
        RECT 201.720 7.240 202.040 7.560 ;
        RECT 202.120 7.240 202.440 7.560 ;
        RECT 202.520 7.240 202.840 7.560 ;
        RECT 202.920 7.240 203.240 7.560 ;
        RECT 203.320 7.240 203.640 7.560 ;
        RECT 203.720 7.240 204.040 7.560 ;
        RECT 204.120 7.240 204.440 7.560 ;
        RECT 204.520 7.240 204.840 7.560 ;
        RECT 204.920 7.240 205.240 7.560 ;
        RECT 205.320 7.240 205.640 7.560 ;
        RECT 0.040 6.840 0.360 7.160 ;
        RECT 0.440 6.840 0.760 7.160 ;
        RECT 0.840 6.840 1.160 7.160 ;
        RECT 1.240 6.840 1.560 7.160 ;
        RECT 1.640 6.840 1.960 7.160 ;
        RECT 2.040 6.840 2.360 7.160 ;
        RECT 2.440 6.840 2.760 7.160 ;
        RECT 2.840 6.840 3.160 7.160 ;
        RECT 3.240 6.840 3.560 7.160 ;
        RECT 3.640 6.840 3.960 7.160 ;
        RECT 4.040 6.840 4.360 7.160 ;
        RECT 4.440 6.840 4.760 7.160 ;
        RECT 4.840 6.840 5.160 7.160 ;
        RECT 5.240 6.840 5.560 7.160 ;
        RECT 5.640 6.840 5.960 7.160 ;
        RECT 6.040 6.840 6.360 7.160 ;
        RECT 6.440 6.840 6.760 7.160 ;
        RECT 6.840 6.840 7.160 7.160 ;
        RECT 7.240 6.840 7.560 7.160 ;
        RECT 7.640 6.840 7.960 7.160 ;
        RECT 8.040 6.840 8.360 7.160 ;
        RECT 8.440 6.840 8.760 7.160 ;
        RECT 8.840 6.840 9.160 7.160 ;
        RECT 9.240 6.840 9.560 7.160 ;
        RECT 9.640 6.840 9.960 7.160 ;
        RECT 10.040 6.840 10.360 7.160 ;
        RECT 10.440 6.840 10.760 7.160 ;
        RECT 10.840 6.840 11.160 7.160 ;
        RECT 11.240 6.840 11.560 7.160 ;
        RECT 11.640 6.840 11.960 7.160 ;
        RECT 12.040 6.840 12.360 7.160 ;
        RECT 12.440 6.840 12.760 7.160 ;
        RECT 12.840 6.840 13.160 7.160 ;
        RECT 13.240 6.840 13.560 7.160 ;
        RECT 13.640 6.840 13.960 7.160 ;
        RECT 14.040 6.840 14.360 7.160 ;
        RECT 14.440 6.840 14.760 7.160 ;
        RECT 14.840 6.840 15.160 7.160 ;
        RECT 15.240 6.840 15.560 7.160 ;
        RECT 15.640 6.840 15.960 7.160 ;
        RECT 16.040 6.840 16.360 7.160 ;
        RECT 16.440 6.840 16.760 7.160 ;
        RECT 16.840 6.840 17.160 7.160 ;
        RECT 17.240 6.840 17.560 7.160 ;
        RECT 17.640 6.840 17.960 7.160 ;
        RECT 18.040 6.840 18.360 7.160 ;
        RECT 18.440 6.840 18.760 7.160 ;
        RECT 18.840 6.840 19.160 7.160 ;
        RECT 19.240 6.840 19.560 7.160 ;
        RECT 19.640 6.840 19.960 7.160 ;
        RECT 95.560 6.840 95.880 7.160 ;
        RECT 95.960 6.840 96.280 7.160 ;
        RECT 96.360 6.840 96.680 7.160 ;
        RECT 96.760 6.840 97.080 7.160 ;
        RECT 145.560 6.840 145.880 7.160 ;
        RECT 145.960 6.840 146.280 7.160 ;
        RECT 146.360 6.840 146.680 7.160 ;
        RECT 146.760 6.840 147.080 7.160 ;
        RECT 185.720 6.840 186.040 7.160 ;
        RECT 186.120 6.840 186.440 7.160 ;
        RECT 186.520 6.840 186.840 7.160 ;
        RECT 186.920 6.840 187.240 7.160 ;
        RECT 187.320 6.840 187.640 7.160 ;
        RECT 187.720 6.840 188.040 7.160 ;
        RECT 188.120 6.840 188.440 7.160 ;
        RECT 188.520 6.840 188.840 7.160 ;
        RECT 188.920 6.840 189.240 7.160 ;
        RECT 189.320 6.840 189.640 7.160 ;
        RECT 189.720 6.840 190.040 7.160 ;
        RECT 190.120 6.840 190.440 7.160 ;
        RECT 190.520 6.840 190.840 7.160 ;
        RECT 190.920 6.840 191.240 7.160 ;
        RECT 191.320 6.840 191.640 7.160 ;
        RECT 191.720 6.840 192.040 7.160 ;
        RECT 192.120 6.840 192.440 7.160 ;
        RECT 192.520 6.840 192.840 7.160 ;
        RECT 192.920 6.840 193.240 7.160 ;
        RECT 193.320 6.840 193.640 7.160 ;
        RECT 193.720 6.840 194.040 7.160 ;
        RECT 194.120 6.840 194.440 7.160 ;
        RECT 194.520 6.840 194.840 7.160 ;
        RECT 194.920 6.840 195.240 7.160 ;
        RECT 195.320 6.840 195.640 7.160 ;
        RECT 195.720 6.840 196.040 7.160 ;
        RECT 196.120 6.840 196.440 7.160 ;
        RECT 196.520 6.840 196.840 7.160 ;
        RECT 196.920 6.840 197.240 7.160 ;
        RECT 197.320 6.840 197.640 7.160 ;
        RECT 197.720 6.840 198.040 7.160 ;
        RECT 198.120 6.840 198.440 7.160 ;
        RECT 198.520 6.840 198.840 7.160 ;
        RECT 198.920 6.840 199.240 7.160 ;
        RECT 199.320 6.840 199.640 7.160 ;
        RECT 199.720 6.840 200.040 7.160 ;
        RECT 200.120 6.840 200.440 7.160 ;
        RECT 200.520 6.840 200.840 7.160 ;
        RECT 200.920 6.840 201.240 7.160 ;
        RECT 201.320 6.840 201.640 7.160 ;
        RECT 201.720 6.840 202.040 7.160 ;
        RECT 202.120 6.840 202.440 7.160 ;
        RECT 202.520 6.840 202.840 7.160 ;
        RECT 202.920 6.840 203.240 7.160 ;
        RECT 203.320 6.840 203.640 7.160 ;
        RECT 203.720 6.840 204.040 7.160 ;
        RECT 204.120 6.840 204.440 7.160 ;
        RECT 204.520 6.840 204.840 7.160 ;
        RECT 204.920 6.840 205.240 7.160 ;
        RECT 205.320 6.840 205.640 7.160 ;
        RECT 0.040 6.440 0.360 6.760 ;
        RECT 0.440 6.440 0.760 6.760 ;
        RECT 0.840 6.440 1.160 6.760 ;
        RECT 1.240 6.440 1.560 6.760 ;
        RECT 1.640 6.440 1.960 6.760 ;
        RECT 2.040 6.440 2.360 6.760 ;
        RECT 2.440 6.440 2.760 6.760 ;
        RECT 2.840 6.440 3.160 6.760 ;
        RECT 3.240 6.440 3.560 6.760 ;
        RECT 3.640 6.440 3.960 6.760 ;
        RECT 4.040 6.440 4.360 6.760 ;
        RECT 4.440 6.440 4.760 6.760 ;
        RECT 4.840 6.440 5.160 6.760 ;
        RECT 5.240 6.440 5.560 6.760 ;
        RECT 5.640 6.440 5.960 6.760 ;
        RECT 6.040 6.440 6.360 6.760 ;
        RECT 6.440 6.440 6.760 6.760 ;
        RECT 6.840 6.440 7.160 6.760 ;
        RECT 7.240 6.440 7.560 6.760 ;
        RECT 7.640 6.440 7.960 6.760 ;
        RECT 8.040 6.440 8.360 6.760 ;
        RECT 8.440 6.440 8.760 6.760 ;
        RECT 8.840 6.440 9.160 6.760 ;
        RECT 9.240 6.440 9.560 6.760 ;
        RECT 9.640 6.440 9.960 6.760 ;
        RECT 10.040 6.440 10.360 6.760 ;
        RECT 10.440 6.440 10.760 6.760 ;
        RECT 10.840 6.440 11.160 6.760 ;
        RECT 11.240 6.440 11.560 6.760 ;
        RECT 11.640 6.440 11.960 6.760 ;
        RECT 12.040 6.440 12.360 6.760 ;
        RECT 12.440 6.440 12.760 6.760 ;
        RECT 12.840 6.440 13.160 6.760 ;
        RECT 13.240 6.440 13.560 6.760 ;
        RECT 13.640 6.440 13.960 6.760 ;
        RECT 14.040 6.440 14.360 6.760 ;
        RECT 14.440 6.440 14.760 6.760 ;
        RECT 14.840 6.440 15.160 6.760 ;
        RECT 15.240 6.440 15.560 6.760 ;
        RECT 15.640 6.440 15.960 6.760 ;
        RECT 16.040 6.440 16.360 6.760 ;
        RECT 16.440 6.440 16.760 6.760 ;
        RECT 16.840 6.440 17.160 6.760 ;
        RECT 17.240 6.440 17.560 6.760 ;
        RECT 17.640 6.440 17.960 6.760 ;
        RECT 18.040 6.440 18.360 6.760 ;
        RECT 18.440 6.440 18.760 6.760 ;
        RECT 18.840 6.440 19.160 6.760 ;
        RECT 19.240 6.440 19.560 6.760 ;
        RECT 19.640 6.440 19.960 6.760 ;
        RECT 95.560 6.440 95.880 6.760 ;
        RECT 95.960 6.440 96.280 6.760 ;
        RECT 96.360 6.440 96.680 6.760 ;
        RECT 96.760 6.440 97.080 6.760 ;
        RECT 145.560 6.440 145.880 6.760 ;
        RECT 145.960 6.440 146.280 6.760 ;
        RECT 146.360 6.440 146.680 6.760 ;
        RECT 146.760 6.440 147.080 6.760 ;
        RECT 185.720 6.440 186.040 6.760 ;
        RECT 186.120 6.440 186.440 6.760 ;
        RECT 186.520 6.440 186.840 6.760 ;
        RECT 186.920 6.440 187.240 6.760 ;
        RECT 187.320 6.440 187.640 6.760 ;
        RECT 187.720 6.440 188.040 6.760 ;
        RECT 188.120 6.440 188.440 6.760 ;
        RECT 188.520 6.440 188.840 6.760 ;
        RECT 188.920 6.440 189.240 6.760 ;
        RECT 189.320 6.440 189.640 6.760 ;
        RECT 189.720 6.440 190.040 6.760 ;
        RECT 190.120 6.440 190.440 6.760 ;
        RECT 190.520 6.440 190.840 6.760 ;
        RECT 190.920 6.440 191.240 6.760 ;
        RECT 191.320 6.440 191.640 6.760 ;
        RECT 191.720 6.440 192.040 6.760 ;
        RECT 192.120 6.440 192.440 6.760 ;
        RECT 192.520 6.440 192.840 6.760 ;
        RECT 192.920 6.440 193.240 6.760 ;
        RECT 193.320 6.440 193.640 6.760 ;
        RECT 193.720 6.440 194.040 6.760 ;
        RECT 194.120 6.440 194.440 6.760 ;
        RECT 194.520 6.440 194.840 6.760 ;
        RECT 194.920 6.440 195.240 6.760 ;
        RECT 195.320 6.440 195.640 6.760 ;
        RECT 195.720 6.440 196.040 6.760 ;
        RECT 196.120 6.440 196.440 6.760 ;
        RECT 196.520 6.440 196.840 6.760 ;
        RECT 196.920 6.440 197.240 6.760 ;
        RECT 197.320 6.440 197.640 6.760 ;
        RECT 197.720 6.440 198.040 6.760 ;
        RECT 198.120 6.440 198.440 6.760 ;
        RECT 198.520 6.440 198.840 6.760 ;
        RECT 198.920 6.440 199.240 6.760 ;
        RECT 199.320 6.440 199.640 6.760 ;
        RECT 199.720 6.440 200.040 6.760 ;
        RECT 200.120 6.440 200.440 6.760 ;
        RECT 200.520 6.440 200.840 6.760 ;
        RECT 200.920 6.440 201.240 6.760 ;
        RECT 201.320 6.440 201.640 6.760 ;
        RECT 201.720 6.440 202.040 6.760 ;
        RECT 202.120 6.440 202.440 6.760 ;
        RECT 202.520 6.440 202.840 6.760 ;
        RECT 202.920 6.440 203.240 6.760 ;
        RECT 203.320 6.440 203.640 6.760 ;
        RECT 203.720 6.440 204.040 6.760 ;
        RECT 204.120 6.440 204.440 6.760 ;
        RECT 204.520 6.440 204.840 6.760 ;
        RECT 204.920 6.440 205.240 6.760 ;
        RECT 205.320 6.440 205.640 6.760 ;
        RECT 0.040 6.040 0.360 6.360 ;
        RECT 0.440 6.040 0.760 6.360 ;
        RECT 0.840 6.040 1.160 6.360 ;
        RECT 1.240 6.040 1.560 6.360 ;
        RECT 1.640 6.040 1.960 6.360 ;
        RECT 2.040 6.040 2.360 6.360 ;
        RECT 2.440 6.040 2.760 6.360 ;
        RECT 2.840 6.040 3.160 6.360 ;
        RECT 3.240 6.040 3.560 6.360 ;
        RECT 3.640 6.040 3.960 6.360 ;
        RECT 4.040 6.040 4.360 6.360 ;
        RECT 4.440 6.040 4.760 6.360 ;
        RECT 4.840 6.040 5.160 6.360 ;
        RECT 5.240 6.040 5.560 6.360 ;
        RECT 5.640 6.040 5.960 6.360 ;
        RECT 6.040 6.040 6.360 6.360 ;
        RECT 6.440 6.040 6.760 6.360 ;
        RECT 6.840 6.040 7.160 6.360 ;
        RECT 7.240 6.040 7.560 6.360 ;
        RECT 7.640 6.040 7.960 6.360 ;
        RECT 8.040 6.040 8.360 6.360 ;
        RECT 8.440 6.040 8.760 6.360 ;
        RECT 8.840 6.040 9.160 6.360 ;
        RECT 9.240 6.040 9.560 6.360 ;
        RECT 9.640 6.040 9.960 6.360 ;
        RECT 10.040 6.040 10.360 6.360 ;
        RECT 10.440 6.040 10.760 6.360 ;
        RECT 10.840 6.040 11.160 6.360 ;
        RECT 11.240 6.040 11.560 6.360 ;
        RECT 11.640 6.040 11.960 6.360 ;
        RECT 12.040 6.040 12.360 6.360 ;
        RECT 12.440 6.040 12.760 6.360 ;
        RECT 12.840 6.040 13.160 6.360 ;
        RECT 13.240 6.040 13.560 6.360 ;
        RECT 13.640 6.040 13.960 6.360 ;
        RECT 14.040 6.040 14.360 6.360 ;
        RECT 14.440 6.040 14.760 6.360 ;
        RECT 14.840 6.040 15.160 6.360 ;
        RECT 15.240 6.040 15.560 6.360 ;
        RECT 15.640 6.040 15.960 6.360 ;
        RECT 16.040 6.040 16.360 6.360 ;
        RECT 16.440 6.040 16.760 6.360 ;
        RECT 16.840 6.040 17.160 6.360 ;
        RECT 17.240 6.040 17.560 6.360 ;
        RECT 17.640 6.040 17.960 6.360 ;
        RECT 18.040 6.040 18.360 6.360 ;
        RECT 18.440 6.040 18.760 6.360 ;
        RECT 18.840 6.040 19.160 6.360 ;
        RECT 19.240 6.040 19.560 6.360 ;
        RECT 19.640 6.040 19.960 6.360 ;
        RECT 95.560 6.040 95.880 6.360 ;
        RECT 95.960 6.040 96.280 6.360 ;
        RECT 96.360 6.040 96.680 6.360 ;
        RECT 96.760 6.040 97.080 6.360 ;
        RECT 145.560 6.040 145.880 6.360 ;
        RECT 145.960 6.040 146.280 6.360 ;
        RECT 146.360 6.040 146.680 6.360 ;
        RECT 146.760 6.040 147.080 6.360 ;
        RECT 185.720 6.040 186.040 6.360 ;
        RECT 186.120 6.040 186.440 6.360 ;
        RECT 186.520 6.040 186.840 6.360 ;
        RECT 186.920 6.040 187.240 6.360 ;
        RECT 187.320 6.040 187.640 6.360 ;
        RECT 187.720 6.040 188.040 6.360 ;
        RECT 188.120 6.040 188.440 6.360 ;
        RECT 188.520 6.040 188.840 6.360 ;
        RECT 188.920 6.040 189.240 6.360 ;
        RECT 189.320 6.040 189.640 6.360 ;
        RECT 189.720 6.040 190.040 6.360 ;
        RECT 190.120 6.040 190.440 6.360 ;
        RECT 190.520 6.040 190.840 6.360 ;
        RECT 190.920 6.040 191.240 6.360 ;
        RECT 191.320 6.040 191.640 6.360 ;
        RECT 191.720 6.040 192.040 6.360 ;
        RECT 192.120 6.040 192.440 6.360 ;
        RECT 192.520 6.040 192.840 6.360 ;
        RECT 192.920 6.040 193.240 6.360 ;
        RECT 193.320 6.040 193.640 6.360 ;
        RECT 193.720 6.040 194.040 6.360 ;
        RECT 194.120 6.040 194.440 6.360 ;
        RECT 194.520 6.040 194.840 6.360 ;
        RECT 194.920 6.040 195.240 6.360 ;
        RECT 195.320 6.040 195.640 6.360 ;
        RECT 195.720 6.040 196.040 6.360 ;
        RECT 196.120 6.040 196.440 6.360 ;
        RECT 196.520 6.040 196.840 6.360 ;
        RECT 196.920 6.040 197.240 6.360 ;
        RECT 197.320 6.040 197.640 6.360 ;
        RECT 197.720 6.040 198.040 6.360 ;
        RECT 198.120 6.040 198.440 6.360 ;
        RECT 198.520 6.040 198.840 6.360 ;
        RECT 198.920 6.040 199.240 6.360 ;
        RECT 199.320 6.040 199.640 6.360 ;
        RECT 199.720 6.040 200.040 6.360 ;
        RECT 200.120 6.040 200.440 6.360 ;
        RECT 200.520 6.040 200.840 6.360 ;
        RECT 200.920 6.040 201.240 6.360 ;
        RECT 201.320 6.040 201.640 6.360 ;
        RECT 201.720 6.040 202.040 6.360 ;
        RECT 202.120 6.040 202.440 6.360 ;
        RECT 202.520 6.040 202.840 6.360 ;
        RECT 202.920 6.040 203.240 6.360 ;
        RECT 203.320 6.040 203.640 6.360 ;
        RECT 203.720 6.040 204.040 6.360 ;
        RECT 204.120 6.040 204.440 6.360 ;
        RECT 204.520 6.040 204.840 6.360 ;
        RECT 204.920 6.040 205.240 6.360 ;
        RECT 205.320 6.040 205.640 6.360 ;
        RECT 0.040 5.640 0.360 5.960 ;
        RECT 0.440 5.640 0.760 5.960 ;
        RECT 0.840 5.640 1.160 5.960 ;
        RECT 1.240 5.640 1.560 5.960 ;
        RECT 1.640 5.640 1.960 5.960 ;
        RECT 2.040 5.640 2.360 5.960 ;
        RECT 2.440 5.640 2.760 5.960 ;
        RECT 2.840 5.640 3.160 5.960 ;
        RECT 3.240 5.640 3.560 5.960 ;
        RECT 3.640 5.640 3.960 5.960 ;
        RECT 4.040 5.640 4.360 5.960 ;
        RECT 4.440 5.640 4.760 5.960 ;
        RECT 4.840 5.640 5.160 5.960 ;
        RECT 5.240 5.640 5.560 5.960 ;
        RECT 5.640 5.640 5.960 5.960 ;
        RECT 6.040 5.640 6.360 5.960 ;
        RECT 6.440 5.640 6.760 5.960 ;
        RECT 6.840 5.640 7.160 5.960 ;
        RECT 7.240 5.640 7.560 5.960 ;
        RECT 7.640 5.640 7.960 5.960 ;
        RECT 8.040 5.640 8.360 5.960 ;
        RECT 8.440 5.640 8.760 5.960 ;
        RECT 8.840 5.640 9.160 5.960 ;
        RECT 9.240 5.640 9.560 5.960 ;
        RECT 9.640 5.640 9.960 5.960 ;
        RECT 10.040 5.640 10.360 5.960 ;
        RECT 10.440 5.640 10.760 5.960 ;
        RECT 10.840 5.640 11.160 5.960 ;
        RECT 11.240 5.640 11.560 5.960 ;
        RECT 11.640 5.640 11.960 5.960 ;
        RECT 12.040 5.640 12.360 5.960 ;
        RECT 12.440 5.640 12.760 5.960 ;
        RECT 12.840 5.640 13.160 5.960 ;
        RECT 13.240 5.640 13.560 5.960 ;
        RECT 13.640 5.640 13.960 5.960 ;
        RECT 14.040 5.640 14.360 5.960 ;
        RECT 14.440 5.640 14.760 5.960 ;
        RECT 14.840 5.640 15.160 5.960 ;
        RECT 15.240 5.640 15.560 5.960 ;
        RECT 15.640 5.640 15.960 5.960 ;
        RECT 16.040 5.640 16.360 5.960 ;
        RECT 16.440 5.640 16.760 5.960 ;
        RECT 16.840 5.640 17.160 5.960 ;
        RECT 17.240 5.640 17.560 5.960 ;
        RECT 17.640 5.640 17.960 5.960 ;
        RECT 18.040 5.640 18.360 5.960 ;
        RECT 18.440 5.640 18.760 5.960 ;
        RECT 18.840 5.640 19.160 5.960 ;
        RECT 19.240 5.640 19.560 5.960 ;
        RECT 19.640 5.640 19.960 5.960 ;
        RECT 95.560 5.640 95.880 5.960 ;
        RECT 95.960 5.640 96.280 5.960 ;
        RECT 96.360 5.640 96.680 5.960 ;
        RECT 96.760 5.640 97.080 5.960 ;
        RECT 145.560 5.640 145.880 5.960 ;
        RECT 145.960 5.640 146.280 5.960 ;
        RECT 146.360 5.640 146.680 5.960 ;
        RECT 146.760 5.640 147.080 5.960 ;
        RECT 185.720 5.640 186.040 5.960 ;
        RECT 186.120 5.640 186.440 5.960 ;
        RECT 186.520 5.640 186.840 5.960 ;
        RECT 186.920 5.640 187.240 5.960 ;
        RECT 187.320 5.640 187.640 5.960 ;
        RECT 187.720 5.640 188.040 5.960 ;
        RECT 188.120 5.640 188.440 5.960 ;
        RECT 188.520 5.640 188.840 5.960 ;
        RECT 188.920 5.640 189.240 5.960 ;
        RECT 189.320 5.640 189.640 5.960 ;
        RECT 189.720 5.640 190.040 5.960 ;
        RECT 190.120 5.640 190.440 5.960 ;
        RECT 190.520 5.640 190.840 5.960 ;
        RECT 190.920 5.640 191.240 5.960 ;
        RECT 191.320 5.640 191.640 5.960 ;
        RECT 191.720 5.640 192.040 5.960 ;
        RECT 192.120 5.640 192.440 5.960 ;
        RECT 192.520 5.640 192.840 5.960 ;
        RECT 192.920 5.640 193.240 5.960 ;
        RECT 193.320 5.640 193.640 5.960 ;
        RECT 193.720 5.640 194.040 5.960 ;
        RECT 194.120 5.640 194.440 5.960 ;
        RECT 194.520 5.640 194.840 5.960 ;
        RECT 194.920 5.640 195.240 5.960 ;
        RECT 195.320 5.640 195.640 5.960 ;
        RECT 195.720 5.640 196.040 5.960 ;
        RECT 196.120 5.640 196.440 5.960 ;
        RECT 196.520 5.640 196.840 5.960 ;
        RECT 196.920 5.640 197.240 5.960 ;
        RECT 197.320 5.640 197.640 5.960 ;
        RECT 197.720 5.640 198.040 5.960 ;
        RECT 198.120 5.640 198.440 5.960 ;
        RECT 198.520 5.640 198.840 5.960 ;
        RECT 198.920 5.640 199.240 5.960 ;
        RECT 199.320 5.640 199.640 5.960 ;
        RECT 199.720 5.640 200.040 5.960 ;
        RECT 200.120 5.640 200.440 5.960 ;
        RECT 200.520 5.640 200.840 5.960 ;
        RECT 200.920 5.640 201.240 5.960 ;
        RECT 201.320 5.640 201.640 5.960 ;
        RECT 201.720 5.640 202.040 5.960 ;
        RECT 202.120 5.640 202.440 5.960 ;
        RECT 202.520 5.640 202.840 5.960 ;
        RECT 202.920 5.640 203.240 5.960 ;
        RECT 203.320 5.640 203.640 5.960 ;
        RECT 203.720 5.640 204.040 5.960 ;
        RECT 204.120 5.640 204.440 5.960 ;
        RECT 204.520 5.640 204.840 5.960 ;
        RECT 204.920 5.640 205.240 5.960 ;
        RECT 205.320 5.640 205.640 5.960 ;
        RECT 0.040 5.240 0.360 5.560 ;
        RECT 0.440 5.240 0.760 5.560 ;
        RECT 0.840 5.240 1.160 5.560 ;
        RECT 1.240 5.240 1.560 5.560 ;
        RECT 1.640 5.240 1.960 5.560 ;
        RECT 2.040 5.240 2.360 5.560 ;
        RECT 2.440 5.240 2.760 5.560 ;
        RECT 2.840 5.240 3.160 5.560 ;
        RECT 3.240 5.240 3.560 5.560 ;
        RECT 3.640 5.240 3.960 5.560 ;
        RECT 4.040 5.240 4.360 5.560 ;
        RECT 4.440 5.240 4.760 5.560 ;
        RECT 4.840 5.240 5.160 5.560 ;
        RECT 5.240 5.240 5.560 5.560 ;
        RECT 5.640 5.240 5.960 5.560 ;
        RECT 6.040 5.240 6.360 5.560 ;
        RECT 6.440 5.240 6.760 5.560 ;
        RECT 6.840 5.240 7.160 5.560 ;
        RECT 7.240 5.240 7.560 5.560 ;
        RECT 7.640 5.240 7.960 5.560 ;
        RECT 8.040 5.240 8.360 5.560 ;
        RECT 8.440 5.240 8.760 5.560 ;
        RECT 8.840 5.240 9.160 5.560 ;
        RECT 9.240 5.240 9.560 5.560 ;
        RECT 9.640 5.240 9.960 5.560 ;
        RECT 10.040 5.240 10.360 5.560 ;
        RECT 10.440 5.240 10.760 5.560 ;
        RECT 10.840 5.240 11.160 5.560 ;
        RECT 11.240 5.240 11.560 5.560 ;
        RECT 11.640 5.240 11.960 5.560 ;
        RECT 12.040 5.240 12.360 5.560 ;
        RECT 12.440 5.240 12.760 5.560 ;
        RECT 12.840 5.240 13.160 5.560 ;
        RECT 13.240 5.240 13.560 5.560 ;
        RECT 13.640 5.240 13.960 5.560 ;
        RECT 14.040 5.240 14.360 5.560 ;
        RECT 14.440 5.240 14.760 5.560 ;
        RECT 14.840 5.240 15.160 5.560 ;
        RECT 15.240 5.240 15.560 5.560 ;
        RECT 15.640 5.240 15.960 5.560 ;
        RECT 16.040 5.240 16.360 5.560 ;
        RECT 16.440 5.240 16.760 5.560 ;
        RECT 16.840 5.240 17.160 5.560 ;
        RECT 17.240 5.240 17.560 5.560 ;
        RECT 17.640 5.240 17.960 5.560 ;
        RECT 18.040 5.240 18.360 5.560 ;
        RECT 18.440 5.240 18.760 5.560 ;
        RECT 18.840 5.240 19.160 5.560 ;
        RECT 19.240 5.240 19.560 5.560 ;
        RECT 19.640 5.240 19.960 5.560 ;
        RECT 95.560 5.240 95.880 5.560 ;
        RECT 95.960 5.240 96.280 5.560 ;
        RECT 96.360 5.240 96.680 5.560 ;
        RECT 96.760 5.240 97.080 5.560 ;
        RECT 145.560 5.240 145.880 5.560 ;
        RECT 145.960 5.240 146.280 5.560 ;
        RECT 146.360 5.240 146.680 5.560 ;
        RECT 146.760 5.240 147.080 5.560 ;
        RECT 185.720 5.240 186.040 5.560 ;
        RECT 186.120 5.240 186.440 5.560 ;
        RECT 186.520 5.240 186.840 5.560 ;
        RECT 186.920 5.240 187.240 5.560 ;
        RECT 187.320 5.240 187.640 5.560 ;
        RECT 187.720 5.240 188.040 5.560 ;
        RECT 188.120 5.240 188.440 5.560 ;
        RECT 188.520 5.240 188.840 5.560 ;
        RECT 188.920 5.240 189.240 5.560 ;
        RECT 189.320 5.240 189.640 5.560 ;
        RECT 189.720 5.240 190.040 5.560 ;
        RECT 190.120 5.240 190.440 5.560 ;
        RECT 190.520 5.240 190.840 5.560 ;
        RECT 190.920 5.240 191.240 5.560 ;
        RECT 191.320 5.240 191.640 5.560 ;
        RECT 191.720 5.240 192.040 5.560 ;
        RECT 192.120 5.240 192.440 5.560 ;
        RECT 192.520 5.240 192.840 5.560 ;
        RECT 192.920 5.240 193.240 5.560 ;
        RECT 193.320 5.240 193.640 5.560 ;
        RECT 193.720 5.240 194.040 5.560 ;
        RECT 194.120 5.240 194.440 5.560 ;
        RECT 194.520 5.240 194.840 5.560 ;
        RECT 194.920 5.240 195.240 5.560 ;
        RECT 195.320 5.240 195.640 5.560 ;
        RECT 195.720 5.240 196.040 5.560 ;
        RECT 196.120 5.240 196.440 5.560 ;
        RECT 196.520 5.240 196.840 5.560 ;
        RECT 196.920 5.240 197.240 5.560 ;
        RECT 197.320 5.240 197.640 5.560 ;
        RECT 197.720 5.240 198.040 5.560 ;
        RECT 198.120 5.240 198.440 5.560 ;
        RECT 198.520 5.240 198.840 5.560 ;
        RECT 198.920 5.240 199.240 5.560 ;
        RECT 199.320 5.240 199.640 5.560 ;
        RECT 199.720 5.240 200.040 5.560 ;
        RECT 200.120 5.240 200.440 5.560 ;
        RECT 200.520 5.240 200.840 5.560 ;
        RECT 200.920 5.240 201.240 5.560 ;
        RECT 201.320 5.240 201.640 5.560 ;
        RECT 201.720 5.240 202.040 5.560 ;
        RECT 202.120 5.240 202.440 5.560 ;
        RECT 202.520 5.240 202.840 5.560 ;
        RECT 202.920 5.240 203.240 5.560 ;
        RECT 203.320 5.240 203.640 5.560 ;
        RECT 203.720 5.240 204.040 5.560 ;
        RECT 204.120 5.240 204.440 5.560 ;
        RECT 204.520 5.240 204.840 5.560 ;
        RECT 204.920 5.240 205.240 5.560 ;
        RECT 205.320 5.240 205.640 5.560 ;
        RECT 0.040 4.840 0.360 5.160 ;
        RECT 0.440 4.840 0.760 5.160 ;
        RECT 0.840 4.840 1.160 5.160 ;
        RECT 1.240 4.840 1.560 5.160 ;
        RECT 1.640 4.840 1.960 5.160 ;
        RECT 2.040 4.840 2.360 5.160 ;
        RECT 2.440 4.840 2.760 5.160 ;
        RECT 2.840 4.840 3.160 5.160 ;
        RECT 3.240 4.840 3.560 5.160 ;
        RECT 3.640 4.840 3.960 5.160 ;
        RECT 4.040 4.840 4.360 5.160 ;
        RECT 4.440 4.840 4.760 5.160 ;
        RECT 4.840 4.840 5.160 5.160 ;
        RECT 5.240 4.840 5.560 5.160 ;
        RECT 5.640 4.840 5.960 5.160 ;
        RECT 6.040 4.840 6.360 5.160 ;
        RECT 6.440 4.840 6.760 5.160 ;
        RECT 6.840 4.840 7.160 5.160 ;
        RECT 7.240 4.840 7.560 5.160 ;
        RECT 7.640 4.840 7.960 5.160 ;
        RECT 8.040 4.840 8.360 5.160 ;
        RECT 8.440 4.840 8.760 5.160 ;
        RECT 8.840 4.840 9.160 5.160 ;
        RECT 9.240 4.840 9.560 5.160 ;
        RECT 9.640 4.840 9.960 5.160 ;
        RECT 10.040 4.840 10.360 5.160 ;
        RECT 10.440 4.840 10.760 5.160 ;
        RECT 10.840 4.840 11.160 5.160 ;
        RECT 11.240 4.840 11.560 5.160 ;
        RECT 11.640 4.840 11.960 5.160 ;
        RECT 12.040 4.840 12.360 5.160 ;
        RECT 12.440 4.840 12.760 5.160 ;
        RECT 12.840 4.840 13.160 5.160 ;
        RECT 13.240 4.840 13.560 5.160 ;
        RECT 13.640 4.840 13.960 5.160 ;
        RECT 14.040 4.840 14.360 5.160 ;
        RECT 14.440 4.840 14.760 5.160 ;
        RECT 14.840 4.840 15.160 5.160 ;
        RECT 15.240 4.840 15.560 5.160 ;
        RECT 15.640 4.840 15.960 5.160 ;
        RECT 16.040 4.840 16.360 5.160 ;
        RECT 16.440 4.840 16.760 5.160 ;
        RECT 16.840 4.840 17.160 5.160 ;
        RECT 17.240 4.840 17.560 5.160 ;
        RECT 17.640 4.840 17.960 5.160 ;
        RECT 18.040 4.840 18.360 5.160 ;
        RECT 18.440 4.840 18.760 5.160 ;
        RECT 18.840 4.840 19.160 5.160 ;
        RECT 19.240 4.840 19.560 5.160 ;
        RECT 19.640 4.840 19.960 5.160 ;
        RECT 95.560 4.840 95.880 5.160 ;
        RECT 95.960 4.840 96.280 5.160 ;
        RECT 96.360 4.840 96.680 5.160 ;
        RECT 96.760 4.840 97.080 5.160 ;
        RECT 145.560 4.840 145.880 5.160 ;
        RECT 145.960 4.840 146.280 5.160 ;
        RECT 146.360 4.840 146.680 5.160 ;
        RECT 146.760 4.840 147.080 5.160 ;
        RECT 185.720 4.840 186.040 5.160 ;
        RECT 186.120 4.840 186.440 5.160 ;
        RECT 186.520 4.840 186.840 5.160 ;
        RECT 186.920 4.840 187.240 5.160 ;
        RECT 187.320 4.840 187.640 5.160 ;
        RECT 187.720 4.840 188.040 5.160 ;
        RECT 188.120 4.840 188.440 5.160 ;
        RECT 188.520 4.840 188.840 5.160 ;
        RECT 188.920 4.840 189.240 5.160 ;
        RECT 189.320 4.840 189.640 5.160 ;
        RECT 189.720 4.840 190.040 5.160 ;
        RECT 190.120 4.840 190.440 5.160 ;
        RECT 190.520 4.840 190.840 5.160 ;
        RECT 190.920 4.840 191.240 5.160 ;
        RECT 191.320 4.840 191.640 5.160 ;
        RECT 191.720 4.840 192.040 5.160 ;
        RECT 192.120 4.840 192.440 5.160 ;
        RECT 192.520 4.840 192.840 5.160 ;
        RECT 192.920 4.840 193.240 5.160 ;
        RECT 193.320 4.840 193.640 5.160 ;
        RECT 193.720 4.840 194.040 5.160 ;
        RECT 194.120 4.840 194.440 5.160 ;
        RECT 194.520 4.840 194.840 5.160 ;
        RECT 194.920 4.840 195.240 5.160 ;
        RECT 195.320 4.840 195.640 5.160 ;
        RECT 195.720 4.840 196.040 5.160 ;
        RECT 196.120 4.840 196.440 5.160 ;
        RECT 196.520 4.840 196.840 5.160 ;
        RECT 196.920 4.840 197.240 5.160 ;
        RECT 197.320 4.840 197.640 5.160 ;
        RECT 197.720 4.840 198.040 5.160 ;
        RECT 198.120 4.840 198.440 5.160 ;
        RECT 198.520 4.840 198.840 5.160 ;
        RECT 198.920 4.840 199.240 5.160 ;
        RECT 199.320 4.840 199.640 5.160 ;
        RECT 199.720 4.840 200.040 5.160 ;
        RECT 200.120 4.840 200.440 5.160 ;
        RECT 200.520 4.840 200.840 5.160 ;
        RECT 200.920 4.840 201.240 5.160 ;
        RECT 201.320 4.840 201.640 5.160 ;
        RECT 201.720 4.840 202.040 5.160 ;
        RECT 202.120 4.840 202.440 5.160 ;
        RECT 202.520 4.840 202.840 5.160 ;
        RECT 202.920 4.840 203.240 5.160 ;
        RECT 203.320 4.840 203.640 5.160 ;
        RECT 203.720 4.840 204.040 5.160 ;
        RECT 204.120 4.840 204.440 5.160 ;
        RECT 204.520 4.840 204.840 5.160 ;
        RECT 204.920 4.840 205.240 5.160 ;
        RECT 205.320 4.840 205.640 5.160 ;
        RECT 0.040 4.440 0.360 4.760 ;
        RECT 0.440 4.440 0.760 4.760 ;
        RECT 0.840 4.440 1.160 4.760 ;
        RECT 1.240 4.440 1.560 4.760 ;
        RECT 1.640 4.440 1.960 4.760 ;
        RECT 2.040 4.440 2.360 4.760 ;
        RECT 2.440 4.440 2.760 4.760 ;
        RECT 2.840 4.440 3.160 4.760 ;
        RECT 3.240 4.440 3.560 4.760 ;
        RECT 3.640 4.440 3.960 4.760 ;
        RECT 4.040 4.440 4.360 4.760 ;
        RECT 4.440 4.440 4.760 4.760 ;
        RECT 4.840 4.440 5.160 4.760 ;
        RECT 5.240 4.440 5.560 4.760 ;
        RECT 5.640 4.440 5.960 4.760 ;
        RECT 6.040 4.440 6.360 4.760 ;
        RECT 6.440 4.440 6.760 4.760 ;
        RECT 6.840 4.440 7.160 4.760 ;
        RECT 7.240 4.440 7.560 4.760 ;
        RECT 7.640 4.440 7.960 4.760 ;
        RECT 8.040 4.440 8.360 4.760 ;
        RECT 8.440 4.440 8.760 4.760 ;
        RECT 8.840 4.440 9.160 4.760 ;
        RECT 9.240 4.440 9.560 4.760 ;
        RECT 9.640 4.440 9.960 4.760 ;
        RECT 10.040 4.440 10.360 4.760 ;
        RECT 10.440 4.440 10.760 4.760 ;
        RECT 10.840 4.440 11.160 4.760 ;
        RECT 11.240 4.440 11.560 4.760 ;
        RECT 11.640 4.440 11.960 4.760 ;
        RECT 12.040 4.440 12.360 4.760 ;
        RECT 12.440 4.440 12.760 4.760 ;
        RECT 12.840 4.440 13.160 4.760 ;
        RECT 13.240 4.440 13.560 4.760 ;
        RECT 13.640 4.440 13.960 4.760 ;
        RECT 14.040 4.440 14.360 4.760 ;
        RECT 14.440 4.440 14.760 4.760 ;
        RECT 14.840 4.440 15.160 4.760 ;
        RECT 15.240 4.440 15.560 4.760 ;
        RECT 15.640 4.440 15.960 4.760 ;
        RECT 16.040 4.440 16.360 4.760 ;
        RECT 16.440 4.440 16.760 4.760 ;
        RECT 16.840 4.440 17.160 4.760 ;
        RECT 17.240 4.440 17.560 4.760 ;
        RECT 17.640 4.440 17.960 4.760 ;
        RECT 18.040 4.440 18.360 4.760 ;
        RECT 18.440 4.440 18.760 4.760 ;
        RECT 18.840 4.440 19.160 4.760 ;
        RECT 19.240 4.440 19.560 4.760 ;
        RECT 19.640 4.440 19.960 4.760 ;
        RECT 95.560 4.440 95.880 4.760 ;
        RECT 95.960 4.440 96.280 4.760 ;
        RECT 96.360 4.440 96.680 4.760 ;
        RECT 96.760 4.440 97.080 4.760 ;
        RECT 145.560 4.440 145.880 4.760 ;
        RECT 145.960 4.440 146.280 4.760 ;
        RECT 146.360 4.440 146.680 4.760 ;
        RECT 146.760 4.440 147.080 4.760 ;
        RECT 185.720 4.440 186.040 4.760 ;
        RECT 186.120 4.440 186.440 4.760 ;
        RECT 186.520 4.440 186.840 4.760 ;
        RECT 186.920 4.440 187.240 4.760 ;
        RECT 187.320 4.440 187.640 4.760 ;
        RECT 187.720 4.440 188.040 4.760 ;
        RECT 188.120 4.440 188.440 4.760 ;
        RECT 188.520 4.440 188.840 4.760 ;
        RECT 188.920 4.440 189.240 4.760 ;
        RECT 189.320 4.440 189.640 4.760 ;
        RECT 189.720 4.440 190.040 4.760 ;
        RECT 190.120 4.440 190.440 4.760 ;
        RECT 190.520 4.440 190.840 4.760 ;
        RECT 190.920 4.440 191.240 4.760 ;
        RECT 191.320 4.440 191.640 4.760 ;
        RECT 191.720 4.440 192.040 4.760 ;
        RECT 192.120 4.440 192.440 4.760 ;
        RECT 192.520 4.440 192.840 4.760 ;
        RECT 192.920 4.440 193.240 4.760 ;
        RECT 193.320 4.440 193.640 4.760 ;
        RECT 193.720 4.440 194.040 4.760 ;
        RECT 194.120 4.440 194.440 4.760 ;
        RECT 194.520 4.440 194.840 4.760 ;
        RECT 194.920 4.440 195.240 4.760 ;
        RECT 195.320 4.440 195.640 4.760 ;
        RECT 195.720 4.440 196.040 4.760 ;
        RECT 196.120 4.440 196.440 4.760 ;
        RECT 196.520 4.440 196.840 4.760 ;
        RECT 196.920 4.440 197.240 4.760 ;
        RECT 197.320 4.440 197.640 4.760 ;
        RECT 197.720 4.440 198.040 4.760 ;
        RECT 198.120 4.440 198.440 4.760 ;
        RECT 198.520 4.440 198.840 4.760 ;
        RECT 198.920 4.440 199.240 4.760 ;
        RECT 199.320 4.440 199.640 4.760 ;
        RECT 199.720 4.440 200.040 4.760 ;
        RECT 200.120 4.440 200.440 4.760 ;
        RECT 200.520 4.440 200.840 4.760 ;
        RECT 200.920 4.440 201.240 4.760 ;
        RECT 201.320 4.440 201.640 4.760 ;
        RECT 201.720 4.440 202.040 4.760 ;
        RECT 202.120 4.440 202.440 4.760 ;
        RECT 202.520 4.440 202.840 4.760 ;
        RECT 202.920 4.440 203.240 4.760 ;
        RECT 203.320 4.440 203.640 4.760 ;
        RECT 203.720 4.440 204.040 4.760 ;
        RECT 204.120 4.440 204.440 4.760 ;
        RECT 204.520 4.440 204.840 4.760 ;
        RECT 204.920 4.440 205.240 4.760 ;
        RECT 205.320 4.440 205.640 4.760 ;
        RECT 0.040 4.040 0.360 4.360 ;
        RECT 0.440 4.040 0.760 4.360 ;
        RECT 0.840 4.040 1.160 4.360 ;
        RECT 1.240 4.040 1.560 4.360 ;
        RECT 1.640 4.040 1.960 4.360 ;
        RECT 2.040 4.040 2.360 4.360 ;
        RECT 2.440 4.040 2.760 4.360 ;
        RECT 2.840 4.040 3.160 4.360 ;
        RECT 3.240 4.040 3.560 4.360 ;
        RECT 3.640 4.040 3.960 4.360 ;
        RECT 4.040 4.040 4.360 4.360 ;
        RECT 4.440 4.040 4.760 4.360 ;
        RECT 4.840 4.040 5.160 4.360 ;
        RECT 5.240 4.040 5.560 4.360 ;
        RECT 5.640 4.040 5.960 4.360 ;
        RECT 6.040 4.040 6.360 4.360 ;
        RECT 6.440 4.040 6.760 4.360 ;
        RECT 6.840 4.040 7.160 4.360 ;
        RECT 7.240 4.040 7.560 4.360 ;
        RECT 7.640 4.040 7.960 4.360 ;
        RECT 8.040 4.040 8.360 4.360 ;
        RECT 8.440 4.040 8.760 4.360 ;
        RECT 8.840 4.040 9.160 4.360 ;
        RECT 9.240 4.040 9.560 4.360 ;
        RECT 9.640 4.040 9.960 4.360 ;
        RECT 10.040 4.040 10.360 4.360 ;
        RECT 10.440 4.040 10.760 4.360 ;
        RECT 10.840 4.040 11.160 4.360 ;
        RECT 11.240 4.040 11.560 4.360 ;
        RECT 11.640 4.040 11.960 4.360 ;
        RECT 12.040 4.040 12.360 4.360 ;
        RECT 12.440 4.040 12.760 4.360 ;
        RECT 12.840 4.040 13.160 4.360 ;
        RECT 13.240 4.040 13.560 4.360 ;
        RECT 13.640 4.040 13.960 4.360 ;
        RECT 14.040 4.040 14.360 4.360 ;
        RECT 14.440 4.040 14.760 4.360 ;
        RECT 14.840 4.040 15.160 4.360 ;
        RECT 15.240 4.040 15.560 4.360 ;
        RECT 15.640 4.040 15.960 4.360 ;
        RECT 16.040 4.040 16.360 4.360 ;
        RECT 16.440 4.040 16.760 4.360 ;
        RECT 16.840 4.040 17.160 4.360 ;
        RECT 17.240 4.040 17.560 4.360 ;
        RECT 17.640 4.040 17.960 4.360 ;
        RECT 18.040 4.040 18.360 4.360 ;
        RECT 18.440 4.040 18.760 4.360 ;
        RECT 18.840 4.040 19.160 4.360 ;
        RECT 19.240 4.040 19.560 4.360 ;
        RECT 19.640 4.040 19.960 4.360 ;
        RECT 95.560 4.040 95.880 4.360 ;
        RECT 95.960 4.040 96.280 4.360 ;
        RECT 96.360 4.040 96.680 4.360 ;
        RECT 96.760 4.040 97.080 4.360 ;
        RECT 145.560 4.040 145.880 4.360 ;
        RECT 145.960 4.040 146.280 4.360 ;
        RECT 146.360 4.040 146.680 4.360 ;
        RECT 146.760 4.040 147.080 4.360 ;
        RECT 185.720 4.040 186.040 4.360 ;
        RECT 186.120 4.040 186.440 4.360 ;
        RECT 186.520 4.040 186.840 4.360 ;
        RECT 186.920 4.040 187.240 4.360 ;
        RECT 187.320 4.040 187.640 4.360 ;
        RECT 187.720 4.040 188.040 4.360 ;
        RECT 188.120 4.040 188.440 4.360 ;
        RECT 188.520 4.040 188.840 4.360 ;
        RECT 188.920 4.040 189.240 4.360 ;
        RECT 189.320 4.040 189.640 4.360 ;
        RECT 189.720 4.040 190.040 4.360 ;
        RECT 190.120 4.040 190.440 4.360 ;
        RECT 190.520 4.040 190.840 4.360 ;
        RECT 190.920 4.040 191.240 4.360 ;
        RECT 191.320 4.040 191.640 4.360 ;
        RECT 191.720 4.040 192.040 4.360 ;
        RECT 192.120 4.040 192.440 4.360 ;
        RECT 192.520 4.040 192.840 4.360 ;
        RECT 192.920 4.040 193.240 4.360 ;
        RECT 193.320 4.040 193.640 4.360 ;
        RECT 193.720 4.040 194.040 4.360 ;
        RECT 194.120 4.040 194.440 4.360 ;
        RECT 194.520 4.040 194.840 4.360 ;
        RECT 194.920 4.040 195.240 4.360 ;
        RECT 195.320 4.040 195.640 4.360 ;
        RECT 195.720 4.040 196.040 4.360 ;
        RECT 196.120 4.040 196.440 4.360 ;
        RECT 196.520 4.040 196.840 4.360 ;
        RECT 196.920 4.040 197.240 4.360 ;
        RECT 197.320 4.040 197.640 4.360 ;
        RECT 197.720 4.040 198.040 4.360 ;
        RECT 198.120 4.040 198.440 4.360 ;
        RECT 198.520 4.040 198.840 4.360 ;
        RECT 198.920 4.040 199.240 4.360 ;
        RECT 199.320 4.040 199.640 4.360 ;
        RECT 199.720 4.040 200.040 4.360 ;
        RECT 200.120 4.040 200.440 4.360 ;
        RECT 200.520 4.040 200.840 4.360 ;
        RECT 200.920 4.040 201.240 4.360 ;
        RECT 201.320 4.040 201.640 4.360 ;
        RECT 201.720 4.040 202.040 4.360 ;
        RECT 202.120 4.040 202.440 4.360 ;
        RECT 202.520 4.040 202.840 4.360 ;
        RECT 202.920 4.040 203.240 4.360 ;
        RECT 203.320 4.040 203.640 4.360 ;
        RECT 203.720 4.040 204.040 4.360 ;
        RECT 204.120 4.040 204.440 4.360 ;
        RECT 204.520 4.040 204.840 4.360 ;
        RECT 204.920 4.040 205.240 4.360 ;
        RECT 205.320 4.040 205.640 4.360 ;
        RECT 0.040 3.640 0.360 3.960 ;
        RECT 0.440 3.640 0.760 3.960 ;
        RECT 0.840 3.640 1.160 3.960 ;
        RECT 1.240 3.640 1.560 3.960 ;
        RECT 1.640 3.640 1.960 3.960 ;
        RECT 2.040 3.640 2.360 3.960 ;
        RECT 2.440 3.640 2.760 3.960 ;
        RECT 2.840 3.640 3.160 3.960 ;
        RECT 3.240 3.640 3.560 3.960 ;
        RECT 3.640 3.640 3.960 3.960 ;
        RECT 4.040 3.640 4.360 3.960 ;
        RECT 4.440 3.640 4.760 3.960 ;
        RECT 4.840 3.640 5.160 3.960 ;
        RECT 5.240 3.640 5.560 3.960 ;
        RECT 5.640 3.640 5.960 3.960 ;
        RECT 6.040 3.640 6.360 3.960 ;
        RECT 6.440 3.640 6.760 3.960 ;
        RECT 6.840 3.640 7.160 3.960 ;
        RECT 7.240 3.640 7.560 3.960 ;
        RECT 7.640 3.640 7.960 3.960 ;
        RECT 8.040 3.640 8.360 3.960 ;
        RECT 8.440 3.640 8.760 3.960 ;
        RECT 8.840 3.640 9.160 3.960 ;
        RECT 9.240 3.640 9.560 3.960 ;
        RECT 9.640 3.640 9.960 3.960 ;
        RECT 10.040 3.640 10.360 3.960 ;
        RECT 10.440 3.640 10.760 3.960 ;
        RECT 10.840 3.640 11.160 3.960 ;
        RECT 11.240 3.640 11.560 3.960 ;
        RECT 11.640 3.640 11.960 3.960 ;
        RECT 12.040 3.640 12.360 3.960 ;
        RECT 12.440 3.640 12.760 3.960 ;
        RECT 12.840 3.640 13.160 3.960 ;
        RECT 13.240 3.640 13.560 3.960 ;
        RECT 13.640 3.640 13.960 3.960 ;
        RECT 14.040 3.640 14.360 3.960 ;
        RECT 14.440 3.640 14.760 3.960 ;
        RECT 14.840 3.640 15.160 3.960 ;
        RECT 15.240 3.640 15.560 3.960 ;
        RECT 15.640 3.640 15.960 3.960 ;
        RECT 16.040 3.640 16.360 3.960 ;
        RECT 16.440 3.640 16.760 3.960 ;
        RECT 16.840 3.640 17.160 3.960 ;
        RECT 17.240 3.640 17.560 3.960 ;
        RECT 17.640 3.640 17.960 3.960 ;
        RECT 18.040 3.640 18.360 3.960 ;
        RECT 18.440 3.640 18.760 3.960 ;
        RECT 18.840 3.640 19.160 3.960 ;
        RECT 19.240 3.640 19.560 3.960 ;
        RECT 19.640 3.640 19.960 3.960 ;
        RECT 95.560 3.640 95.880 3.960 ;
        RECT 95.960 3.640 96.280 3.960 ;
        RECT 96.360 3.640 96.680 3.960 ;
        RECT 96.760 3.640 97.080 3.960 ;
        RECT 145.560 3.640 145.880 3.960 ;
        RECT 145.960 3.640 146.280 3.960 ;
        RECT 146.360 3.640 146.680 3.960 ;
        RECT 146.760 3.640 147.080 3.960 ;
        RECT 185.720 3.640 186.040 3.960 ;
        RECT 186.120 3.640 186.440 3.960 ;
        RECT 186.520 3.640 186.840 3.960 ;
        RECT 186.920 3.640 187.240 3.960 ;
        RECT 187.320 3.640 187.640 3.960 ;
        RECT 187.720 3.640 188.040 3.960 ;
        RECT 188.120 3.640 188.440 3.960 ;
        RECT 188.520 3.640 188.840 3.960 ;
        RECT 188.920 3.640 189.240 3.960 ;
        RECT 189.320 3.640 189.640 3.960 ;
        RECT 189.720 3.640 190.040 3.960 ;
        RECT 190.120 3.640 190.440 3.960 ;
        RECT 190.520 3.640 190.840 3.960 ;
        RECT 190.920 3.640 191.240 3.960 ;
        RECT 191.320 3.640 191.640 3.960 ;
        RECT 191.720 3.640 192.040 3.960 ;
        RECT 192.120 3.640 192.440 3.960 ;
        RECT 192.520 3.640 192.840 3.960 ;
        RECT 192.920 3.640 193.240 3.960 ;
        RECT 193.320 3.640 193.640 3.960 ;
        RECT 193.720 3.640 194.040 3.960 ;
        RECT 194.120 3.640 194.440 3.960 ;
        RECT 194.520 3.640 194.840 3.960 ;
        RECT 194.920 3.640 195.240 3.960 ;
        RECT 195.320 3.640 195.640 3.960 ;
        RECT 195.720 3.640 196.040 3.960 ;
        RECT 196.120 3.640 196.440 3.960 ;
        RECT 196.520 3.640 196.840 3.960 ;
        RECT 196.920 3.640 197.240 3.960 ;
        RECT 197.320 3.640 197.640 3.960 ;
        RECT 197.720 3.640 198.040 3.960 ;
        RECT 198.120 3.640 198.440 3.960 ;
        RECT 198.520 3.640 198.840 3.960 ;
        RECT 198.920 3.640 199.240 3.960 ;
        RECT 199.320 3.640 199.640 3.960 ;
        RECT 199.720 3.640 200.040 3.960 ;
        RECT 200.120 3.640 200.440 3.960 ;
        RECT 200.520 3.640 200.840 3.960 ;
        RECT 200.920 3.640 201.240 3.960 ;
        RECT 201.320 3.640 201.640 3.960 ;
        RECT 201.720 3.640 202.040 3.960 ;
        RECT 202.120 3.640 202.440 3.960 ;
        RECT 202.520 3.640 202.840 3.960 ;
        RECT 202.920 3.640 203.240 3.960 ;
        RECT 203.320 3.640 203.640 3.960 ;
        RECT 203.720 3.640 204.040 3.960 ;
        RECT 204.120 3.640 204.440 3.960 ;
        RECT 204.520 3.640 204.840 3.960 ;
        RECT 204.920 3.640 205.240 3.960 ;
        RECT 205.320 3.640 205.640 3.960 ;
        RECT 0.040 3.240 0.360 3.560 ;
        RECT 0.440 3.240 0.760 3.560 ;
        RECT 0.840 3.240 1.160 3.560 ;
        RECT 1.240 3.240 1.560 3.560 ;
        RECT 1.640 3.240 1.960 3.560 ;
        RECT 2.040 3.240 2.360 3.560 ;
        RECT 2.440 3.240 2.760 3.560 ;
        RECT 2.840 3.240 3.160 3.560 ;
        RECT 3.240 3.240 3.560 3.560 ;
        RECT 3.640 3.240 3.960 3.560 ;
        RECT 4.040 3.240 4.360 3.560 ;
        RECT 4.440 3.240 4.760 3.560 ;
        RECT 4.840 3.240 5.160 3.560 ;
        RECT 5.240 3.240 5.560 3.560 ;
        RECT 5.640 3.240 5.960 3.560 ;
        RECT 6.040 3.240 6.360 3.560 ;
        RECT 6.440 3.240 6.760 3.560 ;
        RECT 6.840 3.240 7.160 3.560 ;
        RECT 7.240 3.240 7.560 3.560 ;
        RECT 7.640 3.240 7.960 3.560 ;
        RECT 8.040 3.240 8.360 3.560 ;
        RECT 8.440 3.240 8.760 3.560 ;
        RECT 8.840 3.240 9.160 3.560 ;
        RECT 9.240 3.240 9.560 3.560 ;
        RECT 9.640 3.240 9.960 3.560 ;
        RECT 10.040 3.240 10.360 3.560 ;
        RECT 10.440 3.240 10.760 3.560 ;
        RECT 10.840 3.240 11.160 3.560 ;
        RECT 11.240 3.240 11.560 3.560 ;
        RECT 11.640 3.240 11.960 3.560 ;
        RECT 12.040 3.240 12.360 3.560 ;
        RECT 12.440 3.240 12.760 3.560 ;
        RECT 12.840 3.240 13.160 3.560 ;
        RECT 13.240 3.240 13.560 3.560 ;
        RECT 13.640 3.240 13.960 3.560 ;
        RECT 14.040 3.240 14.360 3.560 ;
        RECT 14.440 3.240 14.760 3.560 ;
        RECT 14.840 3.240 15.160 3.560 ;
        RECT 15.240 3.240 15.560 3.560 ;
        RECT 15.640 3.240 15.960 3.560 ;
        RECT 16.040 3.240 16.360 3.560 ;
        RECT 16.440 3.240 16.760 3.560 ;
        RECT 16.840 3.240 17.160 3.560 ;
        RECT 17.240 3.240 17.560 3.560 ;
        RECT 17.640 3.240 17.960 3.560 ;
        RECT 18.040 3.240 18.360 3.560 ;
        RECT 18.440 3.240 18.760 3.560 ;
        RECT 18.840 3.240 19.160 3.560 ;
        RECT 19.240 3.240 19.560 3.560 ;
        RECT 19.640 3.240 19.960 3.560 ;
        RECT 95.560 3.240 95.880 3.560 ;
        RECT 95.960 3.240 96.280 3.560 ;
        RECT 96.360 3.240 96.680 3.560 ;
        RECT 96.760 3.240 97.080 3.560 ;
        RECT 145.560 3.240 145.880 3.560 ;
        RECT 145.960 3.240 146.280 3.560 ;
        RECT 146.360 3.240 146.680 3.560 ;
        RECT 146.760 3.240 147.080 3.560 ;
        RECT 185.720 3.240 186.040 3.560 ;
        RECT 186.120 3.240 186.440 3.560 ;
        RECT 186.520 3.240 186.840 3.560 ;
        RECT 186.920 3.240 187.240 3.560 ;
        RECT 187.320 3.240 187.640 3.560 ;
        RECT 187.720 3.240 188.040 3.560 ;
        RECT 188.120 3.240 188.440 3.560 ;
        RECT 188.520 3.240 188.840 3.560 ;
        RECT 188.920 3.240 189.240 3.560 ;
        RECT 189.320 3.240 189.640 3.560 ;
        RECT 189.720 3.240 190.040 3.560 ;
        RECT 190.120 3.240 190.440 3.560 ;
        RECT 190.520 3.240 190.840 3.560 ;
        RECT 190.920 3.240 191.240 3.560 ;
        RECT 191.320 3.240 191.640 3.560 ;
        RECT 191.720 3.240 192.040 3.560 ;
        RECT 192.120 3.240 192.440 3.560 ;
        RECT 192.520 3.240 192.840 3.560 ;
        RECT 192.920 3.240 193.240 3.560 ;
        RECT 193.320 3.240 193.640 3.560 ;
        RECT 193.720 3.240 194.040 3.560 ;
        RECT 194.120 3.240 194.440 3.560 ;
        RECT 194.520 3.240 194.840 3.560 ;
        RECT 194.920 3.240 195.240 3.560 ;
        RECT 195.320 3.240 195.640 3.560 ;
        RECT 195.720 3.240 196.040 3.560 ;
        RECT 196.120 3.240 196.440 3.560 ;
        RECT 196.520 3.240 196.840 3.560 ;
        RECT 196.920 3.240 197.240 3.560 ;
        RECT 197.320 3.240 197.640 3.560 ;
        RECT 197.720 3.240 198.040 3.560 ;
        RECT 198.120 3.240 198.440 3.560 ;
        RECT 198.520 3.240 198.840 3.560 ;
        RECT 198.920 3.240 199.240 3.560 ;
        RECT 199.320 3.240 199.640 3.560 ;
        RECT 199.720 3.240 200.040 3.560 ;
        RECT 200.120 3.240 200.440 3.560 ;
        RECT 200.520 3.240 200.840 3.560 ;
        RECT 200.920 3.240 201.240 3.560 ;
        RECT 201.320 3.240 201.640 3.560 ;
        RECT 201.720 3.240 202.040 3.560 ;
        RECT 202.120 3.240 202.440 3.560 ;
        RECT 202.520 3.240 202.840 3.560 ;
        RECT 202.920 3.240 203.240 3.560 ;
        RECT 203.320 3.240 203.640 3.560 ;
        RECT 203.720 3.240 204.040 3.560 ;
        RECT 204.120 3.240 204.440 3.560 ;
        RECT 204.520 3.240 204.840 3.560 ;
        RECT 204.920 3.240 205.240 3.560 ;
        RECT 205.320 3.240 205.640 3.560 ;
        RECT 0.040 2.840 0.360 3.160 ;
        RECT 0.440 2.840 0.760 3.160 ;
        RECT 0.840 2.840 1.160 3.160 ;
        RECT 1.240 2.840 1.560 3.160 ;
        RECT 1.640 2.840 1.960 3.160 ;
        RECT 2.040 2.840 2.360 3.160 ;
        RECT 2.440 2.840 2.760 3.160 ;
        RECT 2.840 2.840 3.160 3.160 ;
        RECT 3.240 2.840 3.560 3.160 ;
        RECT 3.640 2.840 3.960 3.160 ;
        RECT 4.040 2.840 4.360 3.160 ;
        RECT 4.440 2.840 4.760 3.160 ;
        RECT 4.840 2.840 5.160 3.160 ;
        RECT 5.240 2.840 5.560 3.160 ;
        RECT 5.640 2.840 5.960 3.160 ;
        RECT 6.040 2.840 6.360 3.160 ;
        RECT 6.440 2.840 6.760 3.160 ;
        RECT 6.840 2.840 7.160 3.160 ;
        RECT 7.240 2.840 7.560 3.160 ;
        RECT 7.640 2.840 7.960 3.160 ;
        RECT 8.040 2.840 8.360 3.160 ;
        RECT 8.440 2.840 8.760 3.160 ;
        RECT 8.840 2.840 9.160 3.160 ;
        RECT 9.240 2.840 9.560 3.160 ;
        RECT 9.640 2.840 9.960 3.160 ;
        RECT 10.040 2.840 10.360 3.160 ;
        RECT 10.440 2.840 10.760 3.160 ;
        RECT 10.840 2.840 11.160 3.160 ;
        RECT 11.240 2.840 11.560 3.160 ;
        RECT 11.640 2.840 11.960 3.160 ;
        RECT 12.040 2.840 12.360 3.160 ;
        RECT 12.440 2.840 12.760 3.160 ;
        RECT 12.840 2.840 13.160 3.160 ;
        RECT 13.240 2.840 13.560 3.160 ;
        RECT 13.640 2.840 13.960 3.160 ;
        RECT 14.040 2.840 14.360 3.160 ;
        RECT 14.440 2.840 14.760 3.160 ;
        RECT 14.840 2.840 15.160 3.160 ;
        RECT 15.240 2.840 15.560 3.160 ;
        RECT 15.640 2.840 15.960 3.160 ;
        RECT 16.040 2.840 16.360 3.160 ;
        RECT 16.440 2.840 16.760 3.160 ;
        RECT 16.840 2.840 17.160 3.160 ;
        RECT 17.240 2.840 17.560 3.160 ;
        RECT 17.640 2.840 17.960 3.160 ;
        RECT 18.040 2.840 18.360 3.160 ;
        RECT 18.440 2.840 18.760 3.160 ;
        RECT 18.840 2.840 19.160 3.160 ;
        RECT 19.240 2.840 19.560 3.160 ;
        RECT 19.640 2.840 19.960 3.160 ;
        RECT 95.560 2.840 95.880 3.160 ;
        RECT 95.960 2.840 96.280 3.160 ;
        RECT 96.360 2.840 96.680 3.160 ;
        RECT 96.760 2.840 97.080 3.160 ;
        RECT 145.560 2.840 145.880 3.160 ;
        RECT 145.960 2.840 146.280 3.160 ;
        RECT 146.360 2.840 146.680 3.160 ;
        RECT 146.760 2.840 147.080 3.160 ;
        RECT 185.720 2.840 186.040 3.160 ;
        RECT 186.120 2.840 186.440 3.160 ;
        RECT 186.520 2.840 186.840 3.160 ;
        RECT 186.920 2.840 187.240 3.160 ;
        RECT 187.320 2.840 187.640 3.160 ;
        RECT 187.720 2.840 188.040 3.160 ;
        RECT 188.120 2.840 188.440 3.160 ;
        RECT 188.520 2.840 188.840 3.160 ;
        RECT 188.920 2.840 189.240 3.160 ;
        RECT 189.320 2.840 189.640 3.160 ;
        RECT 189.720 2.840 190.040 3.160 ;
        RECT 190.120 2.840 190.440 3.160 ;
        RECT 190.520 2.840 190.840 3.160 ;
        RECT 190.920 2.840 191.240 3.160 ;
        RECT 191.320 2.840 191.640 3.160 ;
        RECT 191.720 2.840 192.040 3.160 ;
        RECT 192.120 2.840 192.440 3.160 ;
        RECT 192.520 2.840 192.840 3.160 ;
        RECT 192.920 2.840 193.240 3.160 ;
        RECT 193.320 2.840 193.640 3.160 ;
        RECT 193.720 2.840 194.040 3.160 ;
        RECT 194.120 2.840 194.440 3.160 ;
        RECT 194.520 2.840 194.840 3.160 ;
        RECT 194.920 2.840 195.240 3.160 ;
        RECT 195.320 2.840 195.640 3.160 ;
        RECT 195.720 2.840 196.040 3.160 ;
        RECT 196.120 2.840 196.440 3.160 ;
        RECT 196.520 2.840 196.840 3.160 ;
        RECT 196.920 2.840 197.240 3.160 ;
        RECT 197.320 2.840 197.640 3.160 ;
        RECT 197.720 2.840 198.040 3.160 ;
        RECT 198.120 2.840 198.440 3.160 ;
        RECT 198.520 2.840 198.840 3.160 ;
        RECT 198.920 2.840 199.240 3.160 ;
        RECT 199.320 2.840 199.640 3.160 ;
        RECT 199.720 2.840 200.040 3.160 ;
        RECT 200.120 2.840 200.440 3.160 ;
        RECT 200.520 2.840 200.840 3.160 ;
        RECT 200.920 2.840 201.240 3.160 ;
        RECT 201.320 2.840 201.640 3.160 ;
        RECT 201.720 2.840 202.040 3.160 ;
        RECT 202.120 2.840 202.440 3.160 ;
        RECT 202.520 2.840 202.840 3.160 ;
        RECT 202.920 2.840 203.240 3.160 ;
        RECT 203.320 2.840 203.640 3.160 ;
        RECT 203.720 2.840 204.040 3.160 ;
        RECT 204.120 2.840 204.440 3.160 ;
        RECT 204.520 2.840 204.840 3.160 ;
        RECT 204.920 2.840 205.240 3.160 ;
        RECT 205.320 2.840 205.640 3.160 ;
        RECT 0.040 2.440 0.360 2.760 ;
        RECT 0.440 2.440 0.760 2.760 ;
        RECT 0.840 2.440 1.160 2.760 ;
        RECT 1.240 2.440 1.560 2.760 ;
        RECT 1.640 2.440 1.960 2.760 ;
        RECT 2.040 2.440 2.360 2.760 ;
        RECT 2.440 2.440 2.760 2.760 ;
        RECT 2.840 2.440 3.160 2.760 ;
        RECT 3.240 2.440 3.560 2.760 ;
        RECT 3.640 2.440 3.960 2.760 ;
        RECT 4.040 2.440 4.360 2.760 ;
        RECT 4.440 2.440 4.760 2.760 ;
        RECT 4.840 2.440 5.160 2.760 ;
        RECT 5.240 2.440 5.560 2.760 ;
        RECT 5.640 2.440 5.960 2.760 ;
        RECT 6.040 2.440 6.360 2.760 ;
        RECT 6.440 2.440 6.760 2.760 ;
        RECT 6.840 2.440 7.160 2.760 ;
        RECT 7.240 2.440 7.560 2.760 ;
        RECT 7.640 2.440 7.960 2.760 ;
        RECT 8.040 2.440 8.360 2.760 ;
        RECT 8.440 2.440 8.760 2.760 ;
        RECT 8.840 2.440 9.160 2.760 ;
        RECT 9.240 2.440 9.560 2.760 ;
        RECT 9.640 2.440 9.960 2.760 ;
        RECT 10.040 2.440 10.360 2.760 ;
        RECT 10.440 2.440 10.760 2.760 ;
        RECT 10.840 2.440 11.160 2.760 ;
        RECT 11.240 2.440 11.560 2.760 ;
        RECT 11.640 2.440 11.960 2.760 ;
        RECT 12.040 2.440 12.360 2.760 ;
        RECT 12.440 2.440 12.760 2.760 ;
        RECT 12.840 2.440 13.160 2.760 ;
        RECT 13.240 2.440 13.560 2.760 ;
        RECT 13.640 2.440 13.960 2.760 ;
        RECT 14.040 2.440 14.360 2.760 ;
        RECT 14.440 2.440 14.760 2.760 ;
        RECT 14.840 2.440 15.160 2.760 ;
        RECT 15.240 2.440 15.560 2.760 ;
        RECT 15.640 2.440 15.960 2.760 ;
        RECT 16.040 2.440 16.360 2.760 ;
        RECT 16.440 2.440 16.760 2.760 ;
        RECT 16.840 2.440 17.160 2.760 ;
        RECT 17.240 2.440 17.560 2.760 ;
        RECT 17.640 2.440 17.960 2.760 ;
        RECT 18.040 2.440 18.360 2.760 ;
        RECT 18.440 2.440 18.760 2.760 ;
        RECT 18.840 2.440 19.160 2.760 ;
        RECT 19.240 2.440 19.560 2.760 ;
        RECT 19.640 2.440 19.960 2.760 ;
        RECT 95.560 2.440 95.880 2.760 ;
        RECT 95.960 2.440 96.280 2.760 ;
        RECT 96.360 2.440 96.680 2.760 ;
        RECT 96.760 2.440 97.080 2.760 ;
        RECT 145.560 2.440 145.880 2.760 ;
        RECT 145.960 2.440 146.280 2.760 ;
        RECT 146.360 2.440 146.680 2.760 ;
        RECT 146.760 2.440 147.080 2.760 ;
        RECT 185.720 2.440 186.040 2.760 ;
        RECT 186.120 2.440 186.440 2.760 ;
        RECT 186.520 2.440 186.840 2.760 ;
        RECT 186.920 2.440 187.240 2.760 ;
        RECT 187.320 2.440 187.640 2.760 ;
        RECT 187.720 2.440 188.040 2.760 ;
        RECT 188.120 2.440 188.440 2.760 ;
        RECT 188.520 2.440 188.840 2.760 ;
        RECT 188.920 2.440 189.240 2.760 ;
        RECT 189.320 2.440 189.640 2.760 ;
        RECT 189.720 2.440 190.040 2.760 ;
        RECT 190.120 2.440 190.440 2.760 ;
        RECT 190.520 2.440 190.840 2.760 ;
        RECT 190.920 2.440 191.240 2.760 ;
        RECT 191.320 2.440 191.640 2.760 ;
        RECT 191.720 2.440 192.040 2.760 ;
        RECT 192.120 2.440 192.440 2.760 ;
        RECT 192.520 2.440 192.840 2.760 ;
        RECT 192.920 2.440 193.240 2.760 ;
        RECT 193.320 2.440 193.640 2.760 ;
        RECT 193.720 2.440 194.040 2.760 ;
        RECT 194.120 2.440 194.440 2.760 ;
        RECT 194.520 2.440 194.840 2.760 ;
        RECT 194.920 2.440 195.240 2.760 ;
        RECT 195.320 2.440 195.640 2.760 ;
        RECT 195.720 2.440 196.040 2.760 ;
        RECT 196.120 2.440 196.440 2.760 ;
        RECT 196.520 2.440 196.840 2.760 ;
        RECT 196.920 2.440 197.240 2.760 ;
        RECT 197.320 2.440 197.640 2.760 ;
        RECT 197.720 2.440 198.040 2.760 ;
        RECT 198.120 2.440 198.440 2.760 ;
        RECT 198.520 2.440 198.840 2.760 ;
        RECT 198.920 2.440 199.240 2.760 ;
        RECT 199.320 2.440 199.640 2.760 ;
        RECT 199.720 2.440 200.040 2.760 ;
        RECT 200.120 2.440 200.440 2.760 ;
        RECT 200.520 2.440 200.840 2.760 ;
        RECT 200.920 2.440 201.240 2.760 ;
        RECT 201.320 2.440 201.640 2.760 ;
        RECT 201.720 2.440 202.040 2.760 ;
        RECT 202.120 2.440 202.440 2.760 ;
        RECT 202.520 2.440 202.840 2.760 ;
        RECT 202.920 2.440 203.240 2.760 ;
        RECT 203.320 2.440 203.640 2.760 ;
        RECT 203.720 2.440 204.040 2.760 ;
        RECT 204.120 2.440 204.440 2.760 ;
        RECT 204.520 2.440 204.840 2.760 ;
        RECT 204.920 2.440 205.240 2.760 ;
        RECT 205.320 2.440 205.640 2.760 ;
        RECT 0.040 2.040 0.360 2.360 ;
        RECT 0.440 2.040 0.760 2.360 ;
        RECT 0.840 2.040 1.160 2.360 ;
        RECT 1.240 2.040 1.560 2.360 ;
        RECT 1.640 2.040 1.960 2.360 ;
        RECT 2.040 2.040 2.360 2.360 ;
        RECT 2.440 2.040 2.760 2.360 ;
        RECT 2.840 2.040 3.160 2.360 ;
        RECT 3.240 2.040 3.560 2.360 ;
        RECT 3.640 2.040 3.960 2.360 ;
        RECT 4.040 2.040 4.360 2.360 ;
        RECT 4.440 2.040 4.760 2.360 ;
        RECT 4.840 2.040 5.160 2.360 ;
        RECT 5.240 2.040 5.560 2.360 ;
        RECT 5.640 2.040 5.960 2.360 ;
        RECT 6.040 2.040 6.360 2.360 ;
        RECT 6.440 2.040 6.760 2.360 ;
        RECT 6.840 2.040 7.160 2.360 ;
        RECT 7.240 2.040 7.560 2.360 ;
        RECT 7.640 2.040 7.960 2.360 ;
        RECT 8.040 2.040 8.360 2.360 ;
        RECT 8.440 2.040 8.760 2.360 ;
        RECT 8.840 2.040 9.160 2.360 ;
        RECT 9.240 2.040 9.560 2.360 ;
        RECT 9.640 2.040 9.960 2.360 ;
        RECT 10.040 2.040 10.360 2.360 ;
        RECT 10.440 2.040 10.760 2.360 ;
        RECT 10.840 2.040 11.160 2.360 ;
        RECT 11.240 2.040 11.560 2.360 ;
        RECT 11.640 2.040 11.960 2.360 ;
        RECT 12.040 2.040 12.360 2.360 ;
        RECT 12.440 2.040 12.760 2.360 ;
        RECT 12.840 2.040 13.160 2.360 ;
        RECT 13.240 2.040 13.560 2.360 ;
        RECT 13.640 2.040 13.960 2.360 ;
        RECT 14.040 2.040 14.360 2.360 ;
        RECT 14.440 2.040 14.760 2.360 ;
        RECT 14.840 2.040 15.160 2.360 ;
        RECT 15.240 2.040 15.560 2.360 ;
        RECT 15.640 2.040 15.960 2.360 ;
        RECT 16.040 2.040 16.360 2.360 ;
        RECT 16.440 2.040 16.760 2.360 ;
        RECT 16.840 2.040 17.160 2.360 ;
        RECT 17.240 2.040 17.560 2.360 ;
        RECT 17.640 2.040 17.960 2.360 ;
        RECT 18.040 2.040 18.360 2.360 ;
        RECT 18.440 2.040 18.760 2.360 ;
        RECT 18.840 2.040 19.160 2.360 ;
        RECT 19.240 2.040 19.560 2.360 ;
        RECT 19.640 2.040 19.960 2.360 ;
        RECT 95.560 2.040 95.880 2.360 ;
        RECT 95.960 2.040 96.280 2.360 ;
        RECT 96.360 2.040 96.680 2.360 ;
        RECT 96.760 2.040 97.080 2.360 ;
        RECT 145.560 2.040 145.880 2.360 ;
        RECT 145.960 2.040 146.280 2.360 ;
        RECT 146.360 2.040 146.680 2.360 ;
        RECT 146.760 2.040 147.080 2.360 ;
        RECT 185.720 2.040 186.040 2.360 ;
        RECT 186.120 2.040 186.440 2.360 ;
        RECT 186.520 2.040 186.840 2.360 ;
        RECT 186.920 2.040 187.240 2.360 ;
        RECT 187.320 2.040 187.640 2.360 ;
        RECT 187.720 2.040 188.040 2.360 ;
        RECT 188.120 2.040 188.440 2.360 ;
        RECT 188.520 2.040 188.840 2.360 ;
        RECT 188.920 2.040 189.240 2.360 ;
        RECT 189.320 2.040 189.640 2.360 ;
        RECT 189.720 2.040 190.040 2.360 ;
        RECT 190.120 2.040 190.440 2.360 ;
        RECT 190.520 2.040 190.840 2.360 ;
        RECT 190.920 2.040 191.240 2.360 ;
        RECT 191.320 2.040 191.640 2.360 ;
        RECT 191.720 2.040 192.040 2.360 ;
        RECT 192.120 2.040 192.440 2.360 ;
        RECT 192.520 2.040 192.840 2.360 ;
        RECT 192.920 2.040 193.240 2.360 ;
        RECT 193.320 2.040 193.640 2.360 ;
        RECT 193.720 2.040 194.040 2.360 ;
        RECT 194.120 2.040 194.440 2.360 ;
        RECT 194.520 2.040 194.840 2.360 ;
        RECT 194.920 2.040 195.240 2.360 ;
        RECT 195.320 2.040 195.640 2.360 ;
        RECT 195.720 2.040 196.040 2.360 ;
        RECT 196.120 2.040 196.440 2.360 ;
        RECT 196.520 2.040 196.840 2.360 ;
        RECT 196.920 2.040 197.240 2.360 ;
        RECT 197.320 2.040 197.640 2.360 ;
        RECT 197.720 2.040 198.040 2.360 ;
        RECT 198.120 2.040 198.440 2.360 ;
        RECT 198.520 2.040 198.840 2.360 ;
        RECT 198.920 2.040 199.240 2.360 ;
        RECT 199.320 2.040 199.640 2.360 ;
        RECT 199.720 2.040 200.040 2.360 ;
        RECT 200.120 2.040 200.440 2.360 ;
        RECT 200.520 2.040 200.840 2.360 ;
        RECT 200.920 2.040 201.240 2.360 ;
        RECT 201.320 2.040 201.640 2.360 ;
        RECT 201.720 2.040 202.040 2.360 ;
        RECT 202.120 2.040 202.440 2.360 ;
        RECT 202.520 2.040 202.840 2.360 ;
        RECT 202.920 2.040 203.240 2.360 ;
        RECT 203.320 2.040 203.640 2.360 ;
        RECT 203.720 2.040 204.040 2.360 ;
        RECT 204.120 2.040 204.440 2.360 ;
        RECT 204.520 2.040 204.840 2.360 ;
        RECT 204.920 2.040 205.240 2.360 ;
        RECT 205.320 2.040 205.640 2.360 ;
        RECT 0.040 1.640 0.360 1.960 ;
        RECT 0.440 1.640 0.760 1.960 ;
        RECT 0.840 1.640 1.160 1.960 ;
        RECT 1.240 1.640 1.560 1.960 ;
        RECT 1.640 1.640 1.960 1.960 ;
        RECT 2.040 1.640 2.360 1.960 ;
        RECT 2.440 1.640 2.760 1.960 ;
        RECT 2.840 1.640 3.160 1.960 ;
        RECT 3.240 1.640 3.560 1.960 ;
        RECT 3.640 1.640 3.960 1.960 ;
        RECT 4.040 1.640 4.360 1.960 ;
        RECT 4.440 1.640 4.760 1.960 ;
        RECT 4.840 1.640 5.160 1.960 ;
        RECT 5.240 1.640 5.560 1.960 ;
        RECT 5.640 1.640 5.960 1.960 ;
        RECT 6.040 1.640 6.360 1.960 ;
        RECT 6.440 1.640 6.760 1.960 ;
        RECT 6.840 1.640 7.160 1.960 ;
        RECT 7.240 1.640 7.560 1.960 ;
        RECT 7.640 1.640 7.960 1.960 ;
        RECT 8.040 1.640 8.360 1.960 ;
        RECT 8.440 1.640 8.760 1.960 ;
        RECT 8.840 1.640 9.160 1.960 ;
        RECT 9.240 1.640 9.560 1.960 ;
        RECT 9.640 1.640 9.960 1.960 ;
        RECT 10.040 1.640 10.360 1.960 ;
        RECT 10.440 1.640 10.760 1.960 ;
        RECT 10.840 1.640 11.160 1.960 ;
        RECT 11.240 1.640 11.560 1.960 ;
        RECT 11.640 1.640 11.960 1.960 ;
        RECT 12.040 1.640 12.360 1.960 ;
        RECT 12.440 1.640 12.760 1.960 ;
        RECT 12.840 1.640 13.160 1.960 ;
        RECT 13.240 1.640 13.560 1.960 ;
        RECT 13.640 1.640 13.960 1.960 ;
        RECT 14.040 1.640 14.360 1.960 ;
        RECT 14.440 1.640 14.760 1.960 ;
        RECT 14.840 1.640 15.160 1.960 ;
        RECT 15.240 1.640 15.560 1.960 ;
        RECT 15.640 1.640 15.960 1.960 ;
        RECT 16.040 1.640 16.360 1.960 ;
        RECT 16.440 1.640 16.760 1.960 ;
        RECT 16.840 1.640 17.160 1.960 ;
        RECT 17.240 1.640 17.560 1.960 ;
        RECT 17.640 1.640 17.960 1.960 ;
        RECT 18.040 1.640 18.360 1.960 ;
        RECT 18.440 1.640 18.760 1.960 ;
        RECT 18.840 1.640 19.160 1.960 ;
        RECT 19.240 1.640 19.560 1.960 ;
        RECT 19.640 1.640 19.960 1.960 ;
        RECT 95.560 1.640 95.880 1.960 ;
        RECT 95.960 1.640 96.280 1.960 ;
        RECT 96.360 1.640 96.680 1.960 ;
        RECT 96.760 1.640 97.080 1.960 ;
        RECT 145.560 1.640 145.880 1.960 ;
        RECT 145.960 1.640 146.280 1.960 ;
        RECT 146.360 1.640 146.680 1.960 ;
        RECT 146.760 1.640 147.080 1.960 ;
        RECT 185.720 1.640 186.040 1.960 ;
        RECT 186.120 1.640 186.440 1.960 ;
        RECT 186.520 1.640 186.840 1.960 ;
        RECT 186.920 1.640 187.240 1.960 ;
        RECT 187.320 1.640 187.640 1.960 ;
        RECT 187.720 1.640 188.040 1.960 ;
        RECT 188.120 1.640 188.440 1.960 ;
        RECT 188.520 1.640 188.840 1.960 ;
        RECT 188.920 1.640 189.240 1.960 ;
        RECT 189.320 1.640 189.640 1.960 ;
        RECT 189.720 1.640 190.040 1.960 ;
        RECT 190.120 1.640 190.440 1.960 ;
        RECT 190.520 1.640 190.840 1.960 ;
        RECT 190.920 1.640 191.240 1.960 ;
        RECT 191.320 1.640 191.640 1.960 ;
        RECT 191.720 1.640 192.040 1.960 ;
        RECT 192.120 1.640 192.440 1.960 ;
        RECT 192.520 1.640 192.840 1.960 ;
        RECT 192.920 1.640 193.240 1.960 ;
        RECT 193.320 1.640 193.640 1.960 ;
        RECT 193.720 1.640 194.040 1.960 ;
        RECT 194.120 1.640 194.440 1.960 ;
        RECT 194.520 1.640 194.840 1.960 ;
        RECT 194.920 1.640 195.240 1.960 ;
        RECT 195.320 1.640 195.640 1.960 ;
        RECT 195.720 1.640 196.040 1.960 ;
        RECT 196.120 1.640 196.440 1.960 ;
        RECT 196.520 1.640 196.840 1.960 ;
        RECT 196.920 1.640 197.240 1.960 ;
        RECT 197.320 1.640 197.640 1.960 ;
        RECT 197.720 1.640 198.040 1.960 ;
        RECT 198.120 1.640 198.440 1.960 ;
        RECT 198.520 1.640 198.840 1.960 ;
        RECT 198.920 1.640 199.240 1.960 ;
        RECT 199.320 1.640 199.640 1.960 ;
        RECT 199.720 1.640 200.040 1.960 ;
        RECT 200.120 1.640 200.440 1.960 ;
        RECT 200.520 1.640 200.840 1.960 ;
        RECT 200.920 1.640 201.240 1.960 ;
        RECT 201.320 1.640 201.640 1.960 ;
        RECT 201.720 1.640 202.040 1.960 ;
        RECT 202.120 1.640 202.440 1.960 ;
        RECT 202.520 1.640 202.840 1.960 ;
        RECT 202.920 1.640 203.240 1.960 ;
        RECT 203.320 1.640 203.640 1.960 ;
        RECT 203.720 1.640 204.040 1.960 ;
        RECT 204.120 1.640 204.440 1.960 ;
        RECT 204.520 1.640 204.840 1.960 ;
        RECT 204.920 1.640 205.240 1.960 ;
        RECT 205.320 1.640 205.640 1.960 ;
        RECT 0.040 1.240 0.360 1.560 ;
        RECT 0.440 1.240 0.760 1.560 ;
        RECT 0.840 1.240 1.160 1.560 ;
        RECT 1.240 1.240 1.560 1.560 ;
        RECT 1.640 1.240 1.960 1.560 ;
        RECT 2.040 1.240 2.360 1.560 ;
        RECT 2.440 1.240 2.760 1.560 ;
        RECT 2.840 1.240 3.160 1.560 ;
        RECT 3.240 1.240 3.560 1.560 ;
        RECT 3.640 1.240 3.960 1.560 ;
        RECT 4.040 1.240 4.360 1.560 ;
        RECT 4.440 1.240 4.760 1.560 ;
        RECT 4.840 1.240 5.160 1.560 ;
        RECT 5.240 1.240 5.560 1.560 ;
        RECT 5.640 1.240 5.960 1.560 ;
        RECT 6.040 1.240 6.360 1.560 ;
        RECT 6.440 1.240 6.760 1.560 ;
        RECT 6.840 1.240 7.160 1.560 ;
        RECT 7.240 1.240 7.560 1.560 ;
        RECT 7.640 1.240 7.960 1.560 ;
        RECT 8.040 1.240 8.360 1.560 ;
        RECT 8.440 1.240 8.760 1.560 ;
        RECT 8.840 1.240 9.160 1.560 ;
        RECT 9.240 1.240 9.560 1.560 ;
        RECT 9.640 1.240 9.960 1.560 ;
        RECT 10.040 1.240 10.360 1.560 ;
        RECT 10.440 1.240 10.760 1.560 ;
        RECT 10.840 1.240 11.160 1.560 ;
        RECT 11.240 1.240 11.560 1.560 ;
        RECT 11.640 1.240 11.960 1.560 ;
        RECT 12.040 1.240 12.360 1.560 ;
        RECT 12.440 1.240 12.760 1.560 ;
        RECT 12.840 1.240 13.160 1.560 ;
        RECT 13.240 1.240 13.560 1.560 ;
        RECT 13.640 1.240 13.960 1.560 ;
        RECT 14.040 1.240 14.360 1.560 ;
        RECT 14.440 1.240 14.760 1.560 ;
        RECT 14.840 1.240 15.160 1.560 ;
        RECT 15.240 1.240 15.560 1.560 ;
        RECT 15.640 1.240 15.960 1.560 ;
        RECT 16.040 1.240 16.360 1.560 ;
        RECT 16.440 1.240 16.760 1.560 ;
        RECT 16.840 1.240 17.160 1.560 ;
        RECT 17.240 1.240 17.560 1.560 ;
        RECT 17.640 1.240 17.960 1.560 ;
        RECT 18.040 1.240 18.360 1.560 ;
        RECT 18.440 1.240 18.760 1.560 ;
        RECT 18.840 1.240 19.160 1.560 ;
        RECT 19.240 1.240 19.560 1.560 ;
        RECT 19.640 1.240 19.960 1.560 ;
        RECT 95.560 1.240 95.880 1.560 ;
        RECT 95.960 1.240 96.280 1.560 ;
        RECT 96.360 1.240 96.680 1.560 ;
        RECT 96.760 1.240 97.080 1.560 ;
        RECT 145.560 1.240 145.880 1.560 ;
        RECT 145.960 1.240 146.280 1.560 ;
        RECT 146.360 1.240 146.680 1.560 ;
        RECT 146.760 1.240 147.080 1.560 ;
        RECT 185.720 1.240 186.040 1.560 ;
        RECT 186.120 1.240 186.440 1.560 ;
        RECT 186.520 1.240 186.840 1.560 ;
        RECT 186.920 1.240 187.240 1.560 ;
        RECT 187.320 1.240 187.640 1.560 ;
        RECT 187.720 1.240 188.040 1.560 ;
        RECT 188.120 1.240 188.440 1.560 ;
        RECT 188.520 1.240 188.840 1.560 ;
        RECT 188.920 1.240 189.240 1.560 ;
        RECT 189.320 1.240 189.640 1.560 ;
        RECT 189.720 1.240 190.040 1.560 ;
        RECT 190.120 1.240 190.440 1.560 ;
        RECT 190.520 1.240 190.840 1.560 ;
        RECT 190.920 1.240 191.240 1.560 ;
        RECT 191.320 1.240 191.640 1.560 ;
        RECT 191.720 1.240 192.040 1.560 ;
        RECT 192.120 1.240 192.440 1.560 ;
        RECT 192.520 1.240 192.840 1.560 ;
        RECT 192.920 1.240 193.240 1.560 ;
        RECT 193.320 1.240 193.640 1.560 ;
        RECT 193.720 1.240 194.040 1.560 ;
        RECT 194.120 1.240 194.440 1.560 ;
        RECT 194.520 1.240 194.840 1.560 ;
        RECT 194.920 1.240 195.240 1.560 ;
        RECT 195.320 1.240 195.640 1.560 ;
        RECT 195.720 1.240 196.040 1.560 ;
        RECT 196.120 1.240 196.440 1.560 ;
        RECT 196.520 1.240 196.840 1.560 ;
        RECT 196.920 1.240 197.240 1.560 ;
        RECT 197.320 1.240 197.640 1.560 ;
        RECT 197.720 1.240 198.040 1.560 ;
        RECT 198.120 1.240 198.440 1.560 ;
        RECT 198.520 1.240 198.840 1.560 ;
        RECT 198.920 1.240 199.240 1.560 ;
        RECT 199.320 1.240 199.640 1.560 ;
        RECT 199.720 1.240 200.040 1.560 ;
        RECT 200.120 1.240 200.440 1.560 ;
        RECT 200.520 1.240 200.840 1.560 ;
        RECT 200.920 1.240 201.240 1.560 ;
        RECT 201.320 1.240 201.640 1.560 ;
        RECT 201.720 1.240 202.040 1.560 ;
        RECT 202.120 1.240 202.440 1.560 ;
        RECT 202.520 1.240 202.840 1.560 ;
        RECT 202.920 1.240 203.240 1.560 ;
        RECT 203.320 1.240 203.640 1.560 ;
        RECT 203.720 1.240 204.040 1.560 ;
        RECT 204.120 1.240 204.440 1.560 ;
        RECT 204.520 1.240 204.840 1.560 ;
        RECT 204.920 1.240 205.240 1.560 ;
        RECT 205.320 1.240 205.640 1.560 ;
        RECT 0.040 0.840 0.360 1.160 ;
        RECT 0.440 0.840 0.760 1.160 ;
        RECT 0.840 0.840 1.160 1.160 ;
        RECT 1.240 0.840 1.560 1.160 ;
        RECT 1.640 0.840 1.960 1.160 ;
        RECT 2.040 0.840 2.360 1.160 ;
        RECT 2.440 0.840 2.760 1.160 ;
        RECT 2.840 0.840 3.160 1.160 ;
        RECT 3.240 0.840 3.560 1.160 ;
        RECT 3.640 0.840 3.960 1.160 ;
        RECT 4.040 0.840 4.360 1.160 ;
        RECT 4.440 0.840 4.760 1.160 ;
        RECT 4.840 0.840 5.160 1.160 ;
        RECT 5.240 0.840 5.560 1.160 ;
        RECT 5.640 0.840 5.960 1.160 ;
        RECT 6.040 0.840 6.360 1.160 ;
        RECT 6.440 0.840 6.760 1.160 ;
        RECT 6.840 0.840 7.160 1.160 ;
        RECT 7.240 0.840 7.560 1.160 ;
        RECT 7.640 0.840 7.960 1.160 ;
        RECT 8.040 0.840 8.360 1.160 ;
        RECT 8.440 0.840 8.760 1.160 ;
        RECT 8.840 0.840 9.160 1.160 ;
        RECT 9.240 0.840 9.560 1.160 ;
        RECT 9.640 0.840 9.960 1.160 ;
        RECT 10.040 0.840 10.360 1.160 ;
        RECT 10.440 0.840 10.760 1.160 ;
        RECT 10.840 0.840 11.160 1.160 ;
        RECT 11.240 0.840 11.560 1.160 ;
        RECT 11.640 0.840 11.960 1.160 ;
        RECT 12.040 0.840 12.360 1.160 ;
        RECT 12.440 0.840 12.760 1.160 ;
        RECT 12.840 0.840 13.160 1.160 ;
        RECT 13.240 0.840 13.560 1.160 ;
        RECT 13.640 0.840 13.960 1.160 ;
        RECT 14.040 0.840 14.360 1.160 ;
        RECT 14.440 0.840 14.760 1.160 ;
        RECT 14.840 0.840 15.160 1.160 ;
        RECT 15.240 0.840 15.560 1.160 ;
        RECT 15.640 0.840 15.960 1.160 ;
        RECT 16.040 0.840 16.360 1.160 ;
        RECT 16.440 0.840 16.760 1.160 ;
        RECT 16.840 0.840 17.160 1.160 ;
        RECT 17.240 0.840 17.560 1.160 ;
        RECT 17.640 0.840 17.960 1.160 ;
        RECT 18.040 0.840 18.360 1.160 ;
        RECT 18.440 0.840 18.760 1.160 ;
        RECT 18.840 0.840 19.160 1.160 ;
        RECT 19.240 0.840 19.560 1.160 ;
        RECT 19.640 0.840 19.960 1.160 ;
        RECT 95.560 0.840 95.880 1.160 ;
        RECT 95.960 0.840 96.280 1.160 ;
        RECT 96.360 0.840 96.680 1.160 ;
        RECT 96.760 0.840 97.080 1.160 ;
        RECT 145.560 0.840 145.880 1.160 ;
        RECT 145.960 0.840 146.280 1.160 ;
        RECT 146.360 0.840 146.680 1.160 ;
        RECT 146.760 0.840 147.080 1.160 ;
        RECT 185.720 0.840 186.040 1.160 ;
        RECT 186.120 0.840 186.440 1.160 ;
        RECT 186.520 0.840 186.840 1.160 ;
        RECT 186.920 0.840 187.240 1.160 ;
        RECT 187.320 0.840 187.640 1.160 ;
        RECT 187.720 0.840 188.040 1.160 ;
        RECT 188.120 0.840 188.440 1.160 ;
        RECT 188.520 0.840 188.840 1.160 ;
        RECT 188.920 0.840 189.240 1.160 ;
        RECT 189.320 0.840 189.640 1.160 ;
        RECT 189.720 0.840 190.040 1.160 ;
        RECT 190.120 0.840 190.440 1.160 ;
        RECT 190.520 0.840 190.840 1.160 ;
        RECT 190.920 0.840 191.240 1.160 ;
        RECT 191.320 0.840 191.640 1.160 ;
        RECT 191.720 0.840 192.040 1.160 ;
        RECT 192.120 0.840 192.440 1.160 ;
        RECT 192.520 0.840 192.840 1.160 ;
        RECT 192.920 0.840 193.240 1.160 ;
        RECT 193.320 0.840 193.640 1.160 ;
        RECT 193.720 0.840 194.040 1.160 ;
        RECT 194.120 0.840 194.440 1.160 ;
        RECT 194.520 0.840 194.840 1.160 ;
        RECT 194.920 0.840 195.240 1.160 ;
        RECT 195.320 0.840 195.640 1.160 ;
        RECT 195.720 0.840 196.040 1.160 ;
        RECT 196.120 0.840 196.440 1.160 ;
        RECT 196.520 0.840 196.840 1.160 ;
        RECT 196.920 0.840 197.240 1.160 ;
        RECT 197.320 0.840 197.640 1.160 ;
        RECT 197.720 0.840 198.040 1.160 ;
        RECT 198.120 0.840 198.440 1.160 ;
        RECT 198.520 0.840 198.840 1.160 ;
        RECT 198.920 0.840 199.240 1.160 ;
        RECT 199.320 0.840 199.640 1.160 ;
        RECT 199.720 0.840 200.040 1.160 ;
        RECT 200.120 0.840 200.440 1.160 ;
        RECT 200.520 0.840 200.840 1.160 ;
        RECT 200.920 0.840 201.240 1.160 ;
        RECT 201.320 0.840 201.640 1.160 ;
        RECT 201.720 0.840 202.040 1.160 ;
        RECT 202.120 0.840 202.440 1.160 ;
        RECT 202.520 0.840 202.840 1.160 ;
        RECT 202.920 0.840 203.240 1.160 ;
        RECT 203.320 0.840 203.640 1.160 ;
        RECT 203.720 0.840 204.040 1.160 ;
        RECT 204.120 0.840 204.440 1.160 ;
        RECT 204.520 0.840 204.840 1.160 ;
        RECT 204.920 0.840 205.240 1.160 ;
        RECT 205.320 0.840 205.640 1.160 ;
        RECT 0.040 0.440 0.360 0.760 ;
        RECT 0.440 0.440 0.760 0.760 ;
        RECT 0.840 0.440 1.160 0.760 ;
        RECT 1.240 0.440 1.560 0.760 ;
        RECT 1.640 0.440 1.960 0.760 ;
        RECT 2.040 0.440 2.360 0.760 ;
        RECT 2.440 0.440 2.760 0.760 ;
        RECT 2.840 0.440 3.160 0.760 ;
        RECT 3.240 0.440 3.560 0.760 ;
        RECT 3.640 0.440 3.960 0.760 ;
        RECT 4.040 0.440 4.360 0.760 ;
        RECT 4.440 0.440 4.760 0.760 ;
        RECT 4.840 0.440 5.160 0.760 ;
        RECT 5.240 0.440 5.560 0.760 ;
        RECT 5.640 0.440 5.960 0.760 ;
        RECT 6.040 0.440 6.360 0.760 ;
        RECT 6.440 0.440 6.760 0.760 ;
        RECT 6.840 0.440 7.160 0.760 ;
        RECT 7.240 0.440 7.560 0.760 ;
        RECT 7.640 0.440 7.960 0.760 ;
        RECT 8.040 0.440 8.360 0.760 ;
        RECT 8.440 0.440 8.760 0.760 ;
        RECT 8.840 0.440 9.160 0.760 ;
        RECT 9.240 0.440 9.560 0.760 ;
        RECT 9.640 0.440 9.960 0.760 ;
        RECT 10.040 0.440 10.360 0.760 ;
        RECT 10.440 0.440 10.760 0.760 ;
        RECT 10.840 0.440 11.160 0.760 ;
        RECT 11.240 0.440 11.560 0.760 ;
        RECT 11.640 0.440 11.960 0.760 ;
        RECT 12.040 0.440 12.360 0.760 ;
        RECT 12.440 0.440 12.760 0.760 ;
        RECT 12.840 0.440 13.160 0.760 ;
        RECT 13.240 0.440 13.560 0.760 ;
        RECT 13.640 0.440 13.960 0.760 ;
        RECT 14.040 0.440 14.360 0.760 ;
        RECT 14.440 0.440 14.760 0.760 ;
        RECT 14.840 0.440 15.160 0.760 ;
        RECT 15.240 0.440 15.560 0.760 ;
        RECT 15.640 0.440 15.960 0.760 ;
        RECT 16.040 0.440 16.360 0.760 ;
        RECT 16.440 0.440 16.760 0.760 ;
        RECT 16.840 0.440 17.160 0.760 ;
        RECT 17.240 0.440 17.560 0.760 ;
        RECT 17.640 0.440 17.960 0.760 ;
        RECT 18.040 0.440 18.360 0.760 ;
        RECT 18.440 0.440 18.760 0.760 ;
        RECT 18.840 0.440 19.160 0.760 ;
        RECT 19.240 0.440 19.560 0.760 ;
        RECT 19.640 0.440 19.960 0.760 ;
        RECT 95.560 0.440 95.880 0.760 ;
        RECT 95.960 0.440 96.280 0.760 ;
        RECT 96.360 0.440 96.680 0.760 ;
        RECT 96.760 0.440 97.080 0.760 ;
        RECT 145.560 0.440 145.880 0.760 ;
        RECT 145.960 0.440 146.280 0.760 ;
        RECT 146.360 0.440 146.680 0.760 ;
        RECT 146.760 0.440 147.080 0.760 ;
        RECT 185.720 0.440 186.040 0.760 ;
        RECT 186.120 0.440 186.440 0.760 ;
        RECT 186.520 0.440 186.840 0.760 ;
        RECT 186.920 0.440 187.240 0.760 ;
        RECT 187.320 0.440 187.640 0.760 ;
        RECT 187.720 0.440 188.040 0.760 ;
        RECT 188.120 0.440 188.440 0.760 ;
        RECT 188.520 0.440 188.840 0.760 ;
        RECT 188.920 0.440 189.240 0.760 ;
        RECT 189.320 0.440 189.640 0.760 ;
        RECT 189.720 0.440 190.040 0.760 ;
        RECT 190.120 0.440 190.440 0.760 ;
        RECT 190.520 0.440 190.840 0.760 ;
        RECT 190.920 0.440 191.240 0.760 ;
        RECT 191.320 0.440 191.640 0.760 ;
        RECT 191.720 0.440 192.040 0.760 ;
        RECT 192.120 0.440 192.440 0.760 ;
        RECT 192.520 0.440 192.840 0.760 ;
        RECT 192.920 0.440 193.240 0.760 ;
        RECT 193.320 0.440 193.640 0.760 ;
        RECT 193.720 0.440 194.040 0.760 ;
        RECT 194.120 0.440 194.440 0.760 ;
        RECT 194.520 0.440 194.840 0.760 ;
        RECT 194.920 0.440 195.240 0.760 ;
        RECT 195.320 0.440 195.640 0.760 ;
        RECT 195.720 0.440 196.040 0.760 ;
        RECT 196.120 0.440 196.440 0.760 ;
        RECT 196.520 0.440 196.840 0.760 ;
        RECT 196.920 0.440 197.240 0.760 ;
        RECT 197.320 0.440 197.640 0.760 ;
        RECT 197.720 0.440 198.040 0.760 ;
        RECT 198.120 0.440 198.440 0.760 ;
        RECT 198.520 0.440 198.840 0.760 ;
        RECT 198.920 0.440 199.240 0.760 ;
        RECT 199.320 0.440 199.640 0.760 ;
        RECT 199.720 0.440 200.040 0.760 ;
        RECT 200.120 0.440 200.440 0.760 ;
        RECT 200.520 0.440 200.840 0.760 ;
        RECT 200.920 0.440 201.240 0.760 ;
        RECT 201.320 0.440 201.640 0.760 ;
        RECT 201.720 0.440 202.040 0.760 ;
        RECT 202.120 0.440 202.440 0.760 ;
        RECT 202.520 0.440 202.840 0.760 ;
        RECT 202.920 0.440 203.240 0.760 ;
        RECT 203.320 0.440 203.640 0.760 ;
        RECT 203.720 0.440 204.040 0.760 ;
        RECT 204.120 0.440 204.440 0.760 ;
        RECT 204.520 0.440 204.840 0.760 ;
        RECT 204.920 0.440 205.240 0.760 ;
        RECT 205.320 0.440 205.640 0.760 ;
        RECT 0.040 0.040 0.360 0.360 ;
        RECT 0.440 0.040 0.760 0.360 ;
        RECT 0.840 0.040 1.160 0.360 ;
        RECT 1.240 0.040 1.560 0.360 ;
        RECT 1.640 0.040 1.960 0.360 ;
        RECT 2.040 0.040 2.360 0.360 ;
        RECT 2.440 0.040 2.760 0.360 ;
        RECT 2.840 0.040 3.160 0.360 ;
        RECT 3.240 0.040 3.560 0.360 ;
        RECT 3.640 0.040 3.960 0.360 ;
        RECT 4.040 0.040 4.360 0.360 ;
        RECT 4.440 0.040 4.760 0.360 ;
        RECT 4.840 0.040 5.160 0.360 ;
        RECT 5.240 0.040 5.560 0.360 ;
        RECT 5.640 0.040 5.960 0.360 ;
        RECT 6.040 0.040 6.360 0.360 ;
        RECT 6.440 0.040 6.760 0.360 ;
        RECT 6.840 0.040 7.160 0.360 ;
        RECT 7.240 0.040 7.560 0.360 ;
        RECT 7.640 0.040 7.960 0.360 ;
        RECT 8.040 0.040 8.360 0.360 ;
        RECT 8.440 0.040 8.760 0.360 ;
        RECT 8.840 0.040 9.160 0.360 ;
        RECT 9.240 0.040 9.560 0.360 ;
        RECT 9.640 0.040 9.960 0.360 ;
        RECT 10.040 0.040 10.360 0.360 ;
        RECT 10.440 0.040 10.760 0.360 ;
        RECT 10.840 0.040 11.160 0.360 ;
        RECT 11.240 0.040 11.560 0.360 ;
        RECT 11.640 0.040 11.960 0.360 ;
        RECT 12.040 0.040 12.360 0.360 ;
        RECT 12.440 0.040 12.760 0.360 ;
        RECT 12.840 0.040 13.160 0.360 ;
        RECT 13.240 0.040 13.560 0.360 ;
        RECT 13.640 0.040 13.960 0.360 ;
        RECT 14.040 0.040 14.360 0.360 ;
        RECT 14.440 0.040 14.760 0.360 ;
        RECT 14.840 0.040 15.160 0.360 ;
        RECT 15.240 0.040 15.560 0.360 ;
        RECT 15.640 0.040 15.960 0.360 ;
        RECT 16.040 0.040 16.360 0.360 ;
        RECT 16.440 0.040 16.760 0.360 ;
        RECT 16.840 0.040 17.160 0.360 ;
        RECT 17.240 0.040 17.560 0.360 ;
        RECT 17.640 0.040 17.960 0.360 ;
        RECT 18.040 0.040 18.360 0.360 ;
        RECT 18.440 0.040 18.760 0.360 ;
        RECT 18.840 0.040 19.160 0.360 ;
        RECT 19.240 0.040 19.560 0.360 ;
        RECT 19.640 0.040 19.960 0.360 ;
        RECT 95.560 0.040 95.880 0.360 ;
        RECT 95.960 0.040 96.280 0.360 ;
        RECT 96.360 0.040 96.680 0.360 ;
        RECT 96.760 0.040 97.080 0.360 ;
        RECT 145.560 0.040 145.880 0.360 ;
        RECT 145.960 0.040 146.280 0.360 ;
        RECT 146.360 0.040 146.680 0.360 ;
        RECT 146.760 0.040 147.080 0.360 ;
        RECT 185.720 0.040 186.040 0.360 ;
        RECT 186.120 0.040 186.440 0.360 ;
        RECT 186.520 0.040 186.840 0.360 ;
        RECT 186.920 0.040 187.240 0.360 ;
        RECT 187.320 0.040 187.640 0.360 ;
        RECT 187.720 0.040 188.040 0.360 ;
        RECT 188.120 0.040 188.440 0.360 ;
        RECT 188.520 0.040 188.840 0.360 ;
        RECT 188.920 0.040 189.240 0.360 ;
        RECT 189.320 0.040 189.640 0.360 ;
        RECT 189.720 0.040 190.040 0.360 ;
        RECT 190.120 0.040 190.440 0.360 ;
        RECT 190.520 0.040 190.840 0.360 ;
        RECT 190.920 0.040 191.240 0.360 ;
        RECT 191.320 0.040 191.640 0.360 ;
        RECT 191.720 0.040 192.040 0.360 ;
        RECT 192.120 0.040 192.440 0.360 ;
        RECT 192.520 0.040 192.840 0.360 ;
        RECT 192.920 0.040 193.240 0.360 ;
        RECT 193.320 0.040 193.640 0.360 ;
        RECT 193.720 0.040 194.040 0.360 ;
        RECT 194.120 0.040 194.440 0.360 ;
        RECT 194.520 0.040 194.840 0.360 ;
        RECT 194.920 0.040 195.240 0.360 ;
        RECT 195.320 0.040 195.640 0.360 ;
        RECT 195.720 0.040 196.040 0.360 ;
        RECT 196.120 0.040 196.440 0.360 ;
        RECT 196.520 0.040 196.840 0.360 ;
        RECT 196.920 0.040 197.240 0.360 ;
        RECT 197.320 0.040 197.640 0.360 ;
        RECT 197.720 0.040 198.040 0.360 ;
        RECT 198.120 0.040 198.440 0.360 ;
        RECT 198.520 0.040 198.840 0.360 ;
        RECT 198.920 0.040 199.240 0.360 ;
        RECT 199.320 0.040 199.640 0.360 ;
        RECT 199.720 0.040 200.040 0.360 ;
        RECT 200.120 0.040 200.440 0.360 ;
        RECT 200.520 0.040 200.840 0.360 ;
        RECT 200.920 0.040 201.240 0.360 ;
        RECT 201.320 0.040 201.640 0.360 ;
        RECT 201.720 0.040 202.040 0.360 ;
        RECT 202.120 0.040 202.440 0.360 ;
        RECT 202.520 0.040 202.840 0.360 ;
        RECT 202.920 0.040 203.240 0.360 ;
        RECT 203.320 0.040 203.640 0.360 ;
        RECT 203.720 0.040 204.040 0.360 ;
        RECT 204.120 0.040 204.440 0.360 ;
        RECT 204.520 0.040 204.840 0.360 ;
        RECT 204.920 0.040 205.240 0.360 ;
        RECT 205.320 0.040 205.640 0.360 ;
      LAYER met4 ;
        RECT 0.000 0.000 20.000 205.200 ;
        RECT 95.520 151.200 97.120 205.200 ;
        RECT 145.520 151.200 147.120 205.200 ;
        RECT 95.520 0.000 97.120 54.000 ;
        RECT 145.520 0.000 147.120 54.000 ;
        RECT 185.680 0.000 205.680 205.200 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 55.000 54.915 150.680 150.285 ;
      LAYER met1 ;
        RECT 54.000 54.760 150.680 150.440 ;
      LAYER met2 ;
        RECT 56.480 54.000 150.120 151.200 ;
      LAYER met3 ;
        RECT 54.000 54.835 151.680 150.690 ;
      LAYER met4 ;
        RECT 70.520 54.000 147.120 151.200 ;
  END
END digital_pll
END LIBRARY

