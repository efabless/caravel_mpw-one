.subckt decred_hash_macro CLK DATA_AVAILABLE DATA_FROM_HASH[0] DATA_FROM_HASH[1] DATA_FROM_HASH[2]
+ DATA_FROM_HASH[3] DATA_FROM_HASH[4] DATA_FROM_HASH[5] DATA_FROM_HASH[6] DATA_FROM_HASH[7]
+ DATA_TO_HASH[0] DATA_TO_HASH[1] DATA_TO_HASH[2] DATA_TO_HASH[3] DATA_TO_HASH[4]
+ DATA_TO_HASH[5] DATA_TO_HASH[6] DATA_TO_HASH[7] HASH_ADDR[0] HASH_ADDR[1] HASH_ADDR[2]
+ HASH_ADDR[3] HASH_ADDR[4] HASH_ADDR[5] HASH_EN MACRO_RD_SELECT MACRO_WR_SELECT THREAD_COUNT[0]
+ THREAD_COUNT[1] THREAD_COUNT[2] THREAD_COUNT[3] VPWR VGND
X_48709_ _46423_/X _82338_/Q _48708_/X _48874_/B sky130_fd_sc_hd__o21ai_4
X_67543_ _67522_/X _67532_/Y _67507_/X _67542_/Y _67543_/X sky130_fd_sc_hd__a211o_4
X_79529_ _79528_/Y _79529_/B _79529_/Y sky130_fd_sc_hd__nand2_4
X_64755_ _64883_/A _64755_/B _64755_/X sky130_fd_sc_hd__and2_4
X_61967_ _61510_/X _61933_/X _61967_/C _61952_/D _61967_/Y sky130_fd_sc_hd__nand4_4
X_49689_ _49688_/X _49699_/A sky130_fd_sc_hd__buf_2
X_51720_ _52688_/A _52605_/A sky130_fd_sc_hd__buf_2
X_63706_ _63697_/A _64544_/C _63458_/A _63706_/X sky130_fd_sc_hd__and3_4
X_82540_ _82553_/CLK _82540_/D _82540_/Q sky130_fd_sc_hd__dfxtp_4
X_60918_ _64172_/C _60918_/X sky130_fd_sc_hd__buf_2
X_67474_ _67497_/A _87661_/Q _67474_/X sky130_fd_sc_hd__and2_4
X_64686_ _64682_/X _64937_/B _64685_/X _64686_/Y sky130_fd_sc_hd__nand3_4
X_61898_ _61820_/A _61960_/B sky130_fd_sc_hd__buf_2
X_69213_ _68507_/X _68511_/X _69212_/X _69213_/Y sky130_fd_sc_hd__a21oi_4
X_66425_ _84126_/Q _65296_/X _66424_/Y _66425_/X sky130_fd_sc_hd__a21o_4
X_51651_ _51629_/X _51651_/B _51651_/C _53177_/D _51651_/X sky130_fd_sc_hd__and4_4
X_63637_ _63634_/Y _63635_/X _63636_/Y _63637_/Y sky130_fd_sc_hd__a21oi_4
X_82471_ _82589_/CLK _82471_/D _78296_/B sky130_fd_sc_hd__dfxtp_4
X_60849_ _60844_/X _60857_/D _60909_/A sky130_fd_sc_hd__and2_4
X_84210_ _84210_/CLK _84210_/D _84210_/Q sky130_fd_sc_hd__dfxtp_4
X_50602_ _50598_/Y _50577_/X _50601_/Y _86170_/D sky130_fd_sc_hd__a21boi_4
X_81422_ _81333_/CLK _81454_/Q _76013_/B sky130_fd_sc_hd__dfxtp_4
X_69144_ _68929_/X _68357_/Y _69095_/X _69143_/Y _69144_/X sky130_fd_sc_hd__a211o_4
X_54370_ _85454_/Q _54349_/X _54369_/Y _54370_/Y sky130_fd_sc_hd__o21ai_4
X_66356_ _66104_/A _66367_/B sky130_fd_sc_hd__buf_2
X_85190_ _85190_/CLK _56447_/Y _85190_/Q sky130_fd_sc_hd__dfxtp_4
X_51582_ _51590_/A _53109_/B _51582_/Y sky130_fd_sc_hd__nand2_4
X_63568_ _63566_/Y _63516_/X _63567_/Y _84313_/D sky130_fd_sc_hd__a21oi_4
X_53321_ _53347_/A _53330_/B sky130_fd_sc_hd__buf_2
X_65307_ _65307_/A _65833_/B sky130_fd_sc_hd__buf_2
X_84141_ _84175_/CLK _84141_/D _66319_/C sky130_fd_sc_hd__dfxtp_4
X_50533_ _50506_/A _50533_/X sky130_fd_sc_hd__buf_2
X_62519_ _59951_/B _62198_/Y _62520_/A sky130_fd_sc_hd__and2_4
X_81353_ _81351_/CLK _76707_/X _81353_/Q sky130_fd_sc_hd__dfxtp_4
X_69075_ _69071_/X _69074_/X _60014_/X _69075_/Y sky130_fd_sc_hd__a21oi_4
X_66287_ _66284_/X _66286_/X _65937_/X _66287_/X sky130_fd_sc_hd__a21o_4
X_63499_ _58546_/Y _63497_/X _61468_/A _63498_/X _63499_/X sky130_fd_sc_hd__a2bb2o_4
X_56040_ _56039_/Y _56040_/X sky130_fd_sc_hd__buf_2
X_80304_ _80304_/A _80304_/B _82244_/D sky130_fd_sc_hd__xnor2_4
X_68026_ _87138_/Q _68023_/X _68024_/X _68025_/X _68027_/B sky130_fd_sc_hd__a211o_4
X_53252_ _85668_/Q _51929_/X _53251_/Y _53252_/Y sky130_fd_sc_hd__o21ai_4
X_65238_ _65235_/X _65237_/X _65161_/X _65238_/X sky130_fd_sc_hd__a21o_4
X_84072_ _81322_/CLK _84072_/D _81504_/D sky130_fd_sc_hd__dfxtp_4
X_50464_ _50464_/A _50464_/X sky130_fd_sc_hd__buf_2
X_81284_ _81284_/CLK _76972_/X _81284_/Q sky130_fd_sc_hd__dfxtp_4
X_52203_ _52203_/A _52203_/X sky130_fd_sc_hd__buf_2
X_83023_ _83022_/CLK _74593_/Y _45181_/A sky130_fd_sc_hd__dfxtp_4
X_87900_ _87195_/CLK _87900_/D _87900_/Q sky130_fd_sc_hd__dfxtp_4
X_80235_ _80213_/X _80216_/Y _80235_/X sky130_fd_sc_hd__or2_4
X_53183_ _53187_/A _53183_/B _53183_/Y sky130_fd_sc_hd__nand2_4
X_65169_ _84212_/Q _65170_/C sky130_fd_sc_hd__inv_2
X_50395_ _50491_/A _50395_/X sky130_fd_sc_hd__buf_2
X_52134_ _51956_/X _52156_/C sky130_fd_sc_hd__buf_2
X_87831_ _88326_/CLK _87831_/D _69052_/A sky130_fd_sc_hd__dfxtp_4
X_80166_ _60032_/C _84289_/Q _80166_/X sky130_fd_sc_hd__xor2_4
X_57991_ _57991_/A _57991_/B _57991_/Y sky130_fd_sc_hd__nor2_4
X_69977_ _83882_/Q _69955_/X _69976_/X _83882_/D sky130_fd_sc_hd__a21bo_4
X_59730_ _59730_/A _59754_/A sky130_fd_sc_hd__buf_2
X_52065_ _66283_/B _52041_/X _52064_/Y _52065_/Y sky130_fd_sc_hd__o21ai_4
X_56942_ _56561_/X _56930_/X _56931_/X _85121_/Q _57084_/A _56942_/X
+ sky130_fd_sc_hd__a32o_4
X_68928_ _83955_/Q _68838_/X _68927_/X _68928_/X sky130_fd_sc_hd__a21bo_4
X_87762_ _87260_/CLK _42703_/X _68403_/B sky130_fd_sc_hd__dfxtp_4
X_84974_ _86541_/CLK _84974_/D _84974_/Q sky130_fd_sc_hd__dfxtp_4
X_80097_ _80094_/Y _80077_/Y _80096_/X _80098_/B sky130_fd_sc_hd__o21ai_4
X_51016_ _51003_/A _51016_/B _51016_/Y sky130_fd_sc_hd__nand2_4
X_86713_ _86713_/CLK _86713_/D _58672_/A sky130_fd_sc_hd__dfxtp_4
X_83925_ _81473_/CLK _83925_/D _83925_/Q sky130_fd_sc_hd__dfxtp_4
X_59661_ _59661_/A _59662_/C _59805_/A _59661_/D _59679_/A sky130_fd_sc_hd__and4_4
X_56873_ _56872_/Y _56873_/X sky130_fd_sc_hd__buf_2
X_68859_ _68669_/A _68859_/B _68859_/Y sky130_fd_sc_hd__nor2_4
X_87693_ _87126_/CLK _87693_/D _66710_/B sky130_fd_sc_hd__dfxtp_4
X_58612_ _84814_/Q _58599_/X _58604_/X _58611_/X _84814_/D sky130_fd_sc_hd__a2bb2oi_4
X_55824_ _56424_/C _55454_/X _55457_/X _55823_/X _55824_/X sky130_fd_sc_hd__a211o_4
X_86644_ _86005_/CLK _86644_/D _57919_/A sky130_fd_sc_hd__dfxtp_4
X_71870_ _71870_/A _71870_/Y sky130_fd_sc_hd__inv_2
X_59592_ _59539_/A _59598_/A _44003_/X _59564_/A _59579_/A _60392_/B
+ sky130_fd_sc_hd__a41oi_4
X_83856_ _82596_/CLK _83856_/D _82536_/D sky130_fd_sc_hd__dfxtp_4
X_70821_ _47195_/X _70802_/A _70820_/Y _83692_/D sky130_fd_sc_hd__o21ai_4
X_58543_ _58543_/A _58543_/Y sky130_fd_sc_hd__inv_2
X_82807_ _82740_/CLK _82839_/Q _78617_/B sky130_fd_sc_hd__dfxtp_4
X_55755_ _55752_/Y _44095_/X _55754_/X _56117_/B sky130_fd_sc_hd__a21boi_4
X_86575_ _86576_/CLK _48029_/Y _66168_/B sky130_fd_sc_hd__dfxtp_4
X_40981_ _40931_/X _81720_/Q _40980_/X _40982_/A sky130_fd_sc_hd__o21ai_4
X_52967_ _52947_/X _52982_/B _52977_/C _52967_/D _52967_/X sky130_fd_sc_hd__and4_4
X_83787_ _83787_/CLK _70349_/X _74745_/A sky130_fd_sc_hd__dfxtp_4
X_80999_ _80776_/CLK _65294_/C _75617_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_593_0_CLK clkbuf_9_296_0_CLK/X _82084_/CLK sky130_fd_sc_hd__clkbuf_1
X_88314_ _88085_/CLK _40900_/X _88314_/Q sky130_fd_sc_hd__dfxtp_4
X_42720_ _42465_/A _42720_/X sky130_fd_sc_hd__buf_2
X_54706_ _85393_/Q _54703_/X _54705_/Y _54706_/Y sky130_fd_sc_hd__o21ai_4
X_85526_ _85815_/CLK _53999_/Y _85526_/Q sky130_fd_sc_hd__dfxtp_4
X_73540_ _73476_/A _86498_/Q _73540_/X sky130_fd_sc_hd__and2_4
X_51918_ _52626_/A _51919_/C sky130_fd_sc_hd__buf_2
X_70752_ _53127_/B _70740_/A _70751_/Y _83708_/D sky130_fd_sc_hd__o21ai_4
X_82738_ _82152_/CLK _84122_/Q _82738_/Q sky130_fd_sc_hd__dfxtp_4
X_58474_ _58474_/A _58474_/B _58474_/Y sky130_fd_sc_hd__nor2_4
X_55686_ _73024_/B _56171_/A _55686_/C _56171_/C _55686_/Y sky130_fd_sc_hd__nand4_4
X_52898_ _85734_/Q _52874_/X _52897_/Y _52898_/Y sky130_fd_sc_hd__o21ai_4
X_57425_ _55317_/B _57413_/X _57425_/X sky130_fd_sc_hd__or2_4
X_88245_ _88245_/CLK _41279_/Y _69104_/B sky130_fd_sc_hd__dfxtp_4
X_42651_ _52754_/A _42651_/X sky130_fd_sc_hd__buf_2
X_54637_ _85405_/Q _54621_/X _54636_/Y _54637_/Y sky130_fd_sc_hd__o21ai_4
X_73471_ _72721_/X _86181_/Q _73351_/X _73470_/X _73471_/X sky130_fd_sc_hd__a211o_4
X_85457_ _85459_/CLK _85457_/D _85457_/Q sky130_fd_sc_hd__dfxtp_4
X_51849_ _85935_/Q _51846_/X _51848_/Y _51849_/Y sky130_fd_sc_hd__o21ai_4
X_70683_ _70664_/X _47489_/A _70682_/Y _83725_/D sky130_fd_sc_hd__a21o_4
X_82669_ _82675_/CLK _82669_/D _82669_/Q sky130_fd_sc_hd__dfxtp_4
X_75210_ _75217_/B _75210_/B _81035_/D sky130_fd_sc_hd__xor2_4
X_41602_ _41601_/X _41581_/X _67231_/B _41582_/X _88184_/D sky130_fd_sc_hd__a2bb2o_4
X_72422_ _58126_/A _72422_/X sky130_fd_sc_hd__buf_2
X_84408_ _84408_/CLK _62469_/Y _76984_/B sky130_fd_sc_hd__dfxtp_4
X_45370_ _45452_/A _45370_/X sky130_fd_sc_hd__buf_2
X_57356_ _57238_/X _57354_/Y _57355_/Y _85030_/D sky130_fd_sc_hd__o21ai_4
X_88176_ _87473_/CLK _88176_/D _67421_/B sky130_fd_sc_hd__dfxtp_4
X_76190_ _76176_/Y _76171_/Y _76175_/A _76190_/X sky130_fd_sc_hd__o21a_4
X_42582_ _42581_/Y _87813_/D sky130_fd_sc_hd__inv_2
X_54568_ _54486_/A _54578_/A sky130_fd_sc_hd__buf_2
X_85388_ _85484_/CLK _54735_/Y _85388_/Q sky130_fd_sc_hd__dfxtp_4
X_44321_ _41839_/X _40488_/X _41631_/X _87167_/Q _40492_/X _44321_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56307_ _56040_/X _56305_/X _56306_/Y _85242_/D sky130_fd_sc_hd__o21ai_4
X_87127_ _87126_/CLK _87127_/D _87127_/Q sky130_fd_sc_hd__dfxtp_4
X_75141_ _75142_/A _75140_/Y _81063_/Q _75141_/X sky130_fd_sc_hd__a21o_4
X_41533_ _40380_/A _41533_/X sky130_fd_sc_hd__buf_2
X_53519_ _85621_/Q _53506_/X _53518_/Y _53519_/Y sky130_fd_sc_hd__o21ai_4
X_72353_ _72258_/X _85678_/Q _72308_/X _72353_/X sky130_fd_sc_hd__o21a_4
X_84339_ _84263_/CLK _84339_/D _84339_/Q sky130_fd_sc_hd__dfxtp_4
X_57287_ _57286_/X _85040_/D sky130_fd_sc_hd__inv_2
X_54499_ _54497_/Y _54475_/X _54498_/X _54499_/Y sky130_fd_sc_hd__a21oi_4
X_47040_ _47034_/Y _47035_/X _47039_/X _86677_/D sky130_fd_sc_hd__a21oi_4
X_59026_ _84775_/Q _58956_/X _59020_/X _59025_/X _84775_/D sky130_fd_sc_hd__a2bb2oi_4
X_71304_ _50328_/B _71290_/X _71303_/Y _83542_/D sky130_fd_sc_hd__o21ai_4
X_44252_ _58020_/A _44252_/X sky130_fd_sc_hd__buf_2
X_56238_ _56099_/X _56225_/X _56237_/Y _85264_/D sky130_fd_sc_hd__o21ai_4
X_75072_ _75069_/Y _75071_/Y _75072_/Y sky130_fd_sc_hd__nand2_4
X_87058_ _88060_/CLK _87058_/D _73104_/A sky130_fd_sc_hd__dfxtp_4
X_41464_ _41449_/X _82336_/Q _41463_/X _41464_/Y sky130_fd_sc_hd__o21ai_4
X_72284_ _72281_/Y _72283_/Y _72201_/X _72284_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_10_531_0_CLK clkbuf_9_265_0_CLK/X _81346_/CLK sky130_fd_sc_hd__clkbuf_1
X_43203_ _87540_/Q _43203_/Y sky130_fd_sc_hd__inv_2
X_74023_ _74022_/X _86542_/Q _74023_/X sky130_fd_sc_hd__and2_4
X_78900_ _78900_/A _78899_/Y _78901_/B sky130_fd_sc_hd__xor2_4
Xclkbuf_6_22_0_CLK clkbuf_6_23_0_CLK/A clkbuf_6_22_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_86009_ _86008_/CLK _86009_/D _86009_/Q sky130_fd_sc_hd__dfxtp_4
X_40415_ _40414_/X _40416_/A sky130_fd_sc_hd__buf_2
X_71235_ _71235_/A _71091_/B _71232_/C _71235_/Y sky130_fd_sc_hd__nand3_4
X_44183_ _44036_/Y _44184_/A sky130_fd_sc_hd__buf_2
X_56169_ _56169_/A _56150_/B _85283_/Q _56169_/Y sky130_fd_sc_hd__nand3_4
X_79880_ _79878_/Y _79874_/X _79882_/A sky130_fd_sc_hd__nand2_4
X_41395_ _81740_/Q _41325_/X _41395_/X sky130_fd_sc_hd__or2_4
X_43134_ _43046_/X _43125_/X _40802_/X _43133_/Y _43127_/X _87564_/D
+ sky130_fd_sc_hd__o32ai_4
X_78831_ _78831_/A _78831_/B _78831_/X sky130_fd_sc_hd__xor2_4
X_40346_ _40326_/A _86757_/Q _43175_/B _40361_/A sky130_fd_sc_hd__o21a_4
X_71166_ _71170_/A _74531_/B sky130_fd_sc_hd__buf_2
X_48991_ _83614_/Q _72012_/B sky130_fd_sc_hd__inv_2
X_70117_ _70117_/A _70114_/Y _70117_/C _70117_/D _70118_/D sky130_fd_sc_hd__nand4_4
X_47942_ _66055_/B _47897_/X _47941_/Y _47942_/Y sky130_fd_sc_hd__o21ai_4
X_59928_ _59927_/Y _59985_/A sky130_fd_sc_hd__buf_2
X_43065_ _43065_/A _43065_/Y sky130_fd_sc_hd__inv_2
X_78762_ _78762_/A _78761_/X _78762_/X sky130_fd_sc_hd__xor2_4
X_71097_ _71088_/A _71073_/B _71099_/C _71097_/Y sky130_fd_sc_hd__nand3_4
X_75974_ _75948_/Y _75974_/B _75980_/A sky130_fd_sc_hd__nand2_4
Xclkbuf_10_546_0_CLK clkbuf_9_273_0_CLK/X _82642_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_37_0_CLK clkbuf_6_37_0_CLK/A clkbuf_7_74_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_42016_ _42013_/X _42006_/X _40831_/X _73106_/A _42007_/X _42017_/A
+ sky130_fd_sc_hd__o32ai_4
X_77713_ _77698_/Y _77711_/Y _77712_/Y _77713_/Y sky130_fd_sc_hd__o21ai_4
X_74925_ _74930_/A _74912_/X _74924_/Y _74925_/Y sky130_fd_sc_hd__a21boi_4
X_70048_ _70048_/A _70048_/X sky130_fd_sc_hd__buf_2
X_47873_ _52139_/A _52309_/A sky130_fd_sc_hd__buf_2
X_59859_ _59689_/A _59859_/Y sky130_fd_sc_hd__inv_2
X_78693_ _78689_/Y _78690_/Y _78693_/C _78693_/X sky130_fd_sc_hd__or3_4
X_49612_ _49607_/X _52829_/B _49612_/Y sky130_fd_sc_hd__nand2_4
X_46824_ _46824_/A _52696_/B sky130_fd_sc_hd__inv_2
X_77644_ _77643_/B _77644_/Y sky130_fd_sc_hd__inv_2
X_62870_ _61549_/X _62858_/X _62859_/X _62889_/D _62870_/Y sky130_fd_sc_hd__nand4_4
X_74856_ _74855_/Y _74856_/Y sky130_fd_sc_hd__inv_2
X_61821_ _61865_/A _61865_/B _78075_/B _61821_/Y sky130_fd_sc_hd__nor3_4
X_49543_ _49571_/A _49561_/A sky130_fd_sc_hd__buf_2
X_73807_ _73711_/A _66055_/B _73807_/X sky130_fd_sc_hd__and2_4
X_46755_ _46737_/A _46784_/B _46717_/C _52654_/D _46755_/X sky130_fd_sc_hd__and4_4
X_77575_ _77575_/A _77575_/B _77571_/Y _77576_/B sky130_fd_sc_hd__nand3_4
X_43967_ _43957_/A _87186_/Q _43967_/X sky130_fd_sc_hd__and2_4
X_74787_ _70317_/Y _71012_/B _74786_/Y _74787_/Y sky130_fd_sc_hd__o21ai_4
X_71999_ _71997_/Y _71969_/X _71998_/Y _83305_/D sky130_fd_sc_hd__a21boi_4
X_79314_ _79286_/X _79304_/B _79303_/A _79302_/Y _79314_/X sky130_fd_sc_hd__o22a_4
X_45706_ _57430_/A _45705_/X _45691_/X _45706_/X sky130_fd_sc_hd__o21a_4
X_64540_ _64533_/Y _64539_/X _60074_/X _64540_/Y sky130_fd_sc_hd__o21ai_4
X_76526_ _76524_/X _76525_/Y _76526_/X sky130_fd_sc_hd__and2_4
X_42918_ _42916_/X _42917_/X _41710_/X _67691_/B _42905_/X _42919_/A
+ sky130_fd_sc_hd__o32ai_4
X_49474_ _49467_/A _49456_/B _49467_/C _46810_/X _49474_/X sky130_fd_sc_hd__and4_4
X_61752_ _61752_/A _61723_/X _78079_/B _61752_/Y sky130_fd_sc_hd__nor3_4
X_73738_ _73262_/A _73738_/X sky130_fd_sc_hd__buf_2
X_46686_ _46712_/A _46685_/X _46686_/Y sky130_fd_sc_hd__nand2_4
X_43898_ _43895_/X _43876_/X _41332_/X _87210_/Q _43897_/X _43898_/Y
+ sky130_fd_sc_hd__o32ai_4
X_48425_ _65525_/B _48419_/X _48424_/Y _48425_/Y sky130_fd_sc_hd__o21ai_4
X_60703_ _60724_/B _60702_/Y _60703_/Y sky130_fd_sc_hd__nor2_4
X_79245_ _79245_/A _79245_/B _79246_/B sky130_fd_sc_hd__xor2_4
X_45637_ _82994_/Q _45638_/A sky130_fd_sc_hd__inv_2
X_64471_ _64464_/Y _64470_/X _64442_/X _64471_/X sky130_fd_sc_hd__o21a_4
X_76457_ _76456_/Y _76457_/Y sky130_fd_sc_hd__inv_2
X_42849_ _42945_/A _42849_/X sky130_fd_sc_hd__buf_2
X_61683_ _59443_/A _61683_/X sky130_fd_sc_hd__buf_2
X_73669_ _47880_/Y _73668_/Y _73669_/X sky130_fd_sc_hd__xor2_4
X_66210_ _64598_/X _86220_/Q _65761_/X _66209_/X _66210_/X sky130_fd_sc_hd__a211o_4
X_63422_ _60731_/A _63484_/A sky130_fd_sc_hd__buf_2
X_75408_ _75408_/A _75407_/X _80760_/D sky130_fd_sc_hd__xor2_4
X_48356_ _48353_/Y _48302_/X _48355_/X _86530_/D sky130_fd_sc_hd__a21oi_4
X_60634_ _60659_/A _60725_/A sky130_fd_sc_hd__buf_2
X_67190_ _67241_/A _86780_/Q _67190_/X sky130_fd_sc_hd__and2_4
X_79176_ _79176_/A _79175_/Y _79176_/Y sky130_fd_sc_hd__nand2_4
X_45568_ _55514_/B _45516_/X _45396_/X _45567_/Y _45568_/X sky130_fd_sc_hd__a211o_4
X_76388_ _81362_/Q _81618_/D _76388_/X sky130_fd_sc_hd__xor2_4
X_47307_ _47287_/X _52973_/B _47307_/Y sky130_fd_sc_hd__nand2_4
X_66141_ _65932_/A _66141_/B _66141_/X sky130_fd_sc_hd__and2_4
X_78127_ _78130_/D _78126_/Y _78128_/B sky130_fd_sc_hd__xor2_4
X_44519_ _44512_/X _44513_/X _40770_/Y _44518_/Y _44516_/X _87070_/D
+ sky130_fd_sc_hd__o32ai_4
X_63353_ _63351_/Y _63284_/X _63352_/Y _63353_/Y sky130_fd_sc_hd__a21oi_4
X_75339_ _75334_/X _75337_/Y _75339_/C _75339_/Y sky130_fd_sc_hd__nand3_4
X_48287_ _48287_/A _48286_/X _48287_/C _48287_/X sky130_fd_sc_hd__and3_4
X_60565_ _60564_/X _84599_/D sky130_fd_sc_hd__inv_2
X_45499_ _45492_/X _45496_/Y _45498_/Y _45499_/Y sky130_fd_sc_hd__a21oi_4
X_62304_ _62304_/A _58241_/X _62244_/C _62286_/X _62304_/X sky130_fd_sc_hd__and4_4
X_47238_ _47233_/Y _47224_/X _47237_/X _47238_/Y sky130_fd_sc_hd__a21oi_4
X_66072_ _65300_/X _85622_/Q _65301_/X _66071_/X _66072_/X sky130_fd_sc_hd__a211o_4
X_78058_ _84563_/Q _78058_/B _78058_/X sky130_fd_sc_hd__xor2_4
X_63284_ _63516_/A _63284_/X sky130_fd_sc_hd__buf_2
X_60496_ _60105_/X _60526_/A sky130_fd_sc_hd__buf_2
X_69900_ _69900_/A _88314_/Q _69900_/X sky130_fd_sc_hd__and2_4
X_65023_ _64946_/A _85809_/Q _65023_/X sky130_fd_sc_hd__and2_4
X_77009_ _77009_/A _82276_/D _77010_/A sky130_fd_sc_hd__nand2_4
X_62235_ _62193_/A _62628_/C sky130_fd_sc_hd__buf_2
X_47169_ _82375_/Q _47169_/Y sky130_fd_sc_hd__inv_2
X_80020_ _80016_/Y _80019_/Y _80023_/A sky130_fd_sc_hd__xor2_4
X_69831_ _69988_/A _69831_/X sky130_fd_sc_hd__buf_2
X_50180_ _50178_/Y _50166_/X _50179_/X _50180_/Y sky130_fd_sc_hd__a21oi_4
X_62166_ _62033_/A _62166_/X sky130_fd_sc_hd__buf_2
X_61117_ _64546_/A _61117_/X sky130_fd_sc_hd__buf_2
X_69762_ _70009_/A _69988_/A sky130_fd_sc_hd__buf_2
X_66974_ _87874_/Q _66875_/X _66926_/X _66973_/X _66974_/X sky130_fd_sc_hd__a211o_4
X_62097_ _58279_/A _62097_/X sky130_fd_sc_hd__buf_2
X_68713_ _68586_/A _68713_/X sky130_fd_sc_hd__buf_2
X_65925_ _65896_/A _73588_/B _65925_/X sky130_fd_sc_hd__and2_4
Xclkbuf_8_5_0_CLK clkbuf_8_5_0_CLK/A clkbuf_8_5_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_61048_ _60953_/X _61044_/X _61016_/Y _60952_/X _61047_/X _84529_/D
+ sky130_fd_sc_hd__o41a_4
X_81971_ _82116_/CLK _81971_/D _77737_/B sky130_fd_sc_hd__dfxtp_4
X_69693_ _69689_/X _69692_/X _69655_/X _69693_/Y sky130_fd_sc_hd__a21oi_4
X_83710_ _83711_/CLK _70748_/Y _83710_/Q sky130_fd_sc_hd__dfxtp_4
X_80922_ _80928_/CLK _84098_/Q _75787_/A sky130_fd_sc_hd__dfxtp_4
X_68644_ _68644_/A _69092_/A sky130_fd_sc_hd__buf_2
X_53870_ _53661_/A _54295_/A sky130_fd_sc_hd__buf_2
X_65856_ _65854_/Y _65830_/X _65855_/X _84173_/D sky130_fd_sc_hd__a21o_4
X_84690_ _84358_/CLK _59844_/Y _80379_/A sky130_fd_sc_hd__dfxtp_4
X_52821_ _52821_/A _52821_/X sky130_fd_sc_hd__buf_2
X_64807_ _64807_/A _64807_/X sky130_fd_sc_hd__buf_2
X_83641_ _86422_/CLK _70988_/Y _83641_/Q sky130_fd_sc_hd__dfxtp_4
X_80853_ _80854_/CLK _80885_/Q _74980_/B sky130_fd_sc_hd__dfxtp_4
X_68575_ _68553_/A _87755_/Q _68575_/X sky130_fd_sc_hd__and2_4
X_65787_ _65855_/A _65775_/B _84178_/Q _65787_/X sky130_fd_sc_hd__and3_4
X_62999_ _63060_/A _62999_/X sky130_fd_sc_hd__buf_2
X_55540_ _85048_/Q _55510_/X _55512_/X _55539_/Y _55540_/X sky130_fd_sc_hd__a211o_4
X_67526_ _87979_/Q _67473_/X _67524_/X _67525_/X _67526_/X sky130_fd_sc_hd__a211o_4
X_86360_ _86361_/CLK _86360_/D _86360_/Q sky130_fd_sc_hd__dfxtp_4
X_52752_ _52744_/A _52752_/B _52752_/Y sky130_fd_sc_hd__nand2_4
X_64738_ _64738_/A _64739_/A sky130_fd_sc_hd__buf_2
X_83572_ _83572_/CLK _71208_/Y _83572_/Q sky130_fd_sc_hd__dfxtp_4
X_80784_ _80784_/CLK _75719_/Y _80784_/Q sky130_fd_sc_hd__dfxtp_4
X_85311_ _85311_/CLK _56018_/Y _85311_/Q sky130_fd_sc_hd__dfxtp_4
X_51703_ _51717_/A _53227_/B _51703_/Y sky130_fd_sc_hd__nand2_4
X_82523_ _82491_/CLK _79119_/Y _82523_/Q sky130_fd_sc_hd__dfxtp_4
X_55471_ _85107_/Q _55468_/X _55469_/X _55470_/Y _55471_/X sky130_fd_sc_hd__a211o_4
X_67457_ _86970_/Q _67432_/X _67433_/X _67456_/X _67457_/X sky130_fd_sc_hd__a211o_4
X_86291_ _86611_/CLK _86291_/D _72294_/B sky130_fd_sc_hd__dfxtp_4
X_52683_ _52515_/A _52684_/A sky130_fd_sc_hd__buf_2
X_64669_ _64666_/X _86142_/Q _64566_/X _64668_/X _64669_/X sky130_fd_sc_hd__a211o_4
X_57210_ _57049_/A _57210_/B _57086_/X _57210_/Y sky130_fd_sc_hd__nor3_4
X_88030_ _88036_/CLK _42112_/Y _88030_/Q sky130_fd_sc_hd__dfxtp_4
X_54422_ _54475_/A _54422_/X sky130_fd_sc_hd__buf_2
X_66408_ _66405_/Y _66377_/X _66407_/Y _84129_/D sky130_fd_sc_hd__a21o_4
X_85242_ _85241_/CLK _85242_/D _56306_/C sky130_fd_sc_hd__dfxtp_4
X_51634_ _51608_/A _51651_/C sky130_fd_sc_hd__buf_2
X_58190_ _44282_/X _58341_/A sky130_fd_sc_hd__buf_2
X_82454_ _82248_/CLK _79146_/X _82454_/Q sky130_fd_sc_hd__dfxtp_4
X_67388_ _57754_/X _67388_/X sky130_fd_sc_hd__buf_2
X_57141_ _57141_/A _57141_/X sky130_fd_sc_hd__buf_2
X_81405_ _83940_/CLK _81405_/D _76747_/B sky130_fd_sc_hd__dfxtp_4
X_69127_ _69123_/X _69126_/X _69035_/X _69127_/X sky130_fd_sc_hd__a21o_4
X_54353_ _54362_/A _54353_/B _54362_/C _54353_/D _54353_/X sky130_fd_sc_hd__and4_4
X_66339_ _64710_/A _86531_/Q _66339_/X sky130_fd_sc_hd__and2_4
X_85173_ _86900_/CLK _85173_/D _55876_/B sky130_fd_sc_hd__dfxtp_4
X_51565_ _50991_/A _51621_/A sky130_fd_sc_hd__buf_2
X_82385_ _84757_/CLK _82193_/Q _82385_/Q sky130_fd_sc_hd__dfxtp_4
X_53304_ _53299_/Y _53301_/X _53303_/X _53304_/Y sky130_fd_sc_hd__a21oi_4
X_84124_ _84161_/CLK _84124_/D _66433_/C sky130_fd_sc_hd__dfxtp_4
X_50516_ _50514_/Y _50491_/X _50515_/X _50516_/Y sky130_fd_sc_hd__a21oi_4
X_81336_ _81333_/CLK _81336_/D _81712_/D sky130_fd_sc_hd__dfxtp_4
X_57072_ _57070_/X _57071_/Y _56953_/X _57072_/Y sky130_fd_sc_hd__a21oi_4
X_69058_ _69485_/A _69058_/X sky130_fd_sc_hd__buf_2
X_54284_ _54284_/A _54366_/A sky130_fd_sc_hd__buf_2
X_51496_ _51491_/A _53021_/B _51496_/Y sky130_fd_sc_hd__nand2_4
X_56023_ _56023_/A _56017_/B _55963_/B _56023_/Y sky130_fd_sc_hd__nand3_4
X_68009_ _67914_/X _86915_/Q _68009_/X sky130_fd_sc_hd__and2_4
X_53235_ _53233_/Y _53215_/X _53234_/X _53235_/Y sky130_fd_sc_hd__a21oi_4
X_84055_ _81492_/CLK _84055_/D _84055_/Q sky130_fd_sc_hd__dfxtp_4
X_50447_ _50447_/A _50456_/B _50462_/C _50447_/X sky130_fd_sc_hd__and3_4
X_81267_ _81631_/CLK _81267_/D _76393_/A sky130_fd_sc_hd__dfxtp_4
X_71020_ _70768_/A _71171_/A sky130_fd_sc_hd__buf_2
X_83006_ _83008_/CLK _83006_/D _45448_/A sky130_fd_sc_hd__dfxtp_4
X_80218_ _80244_/A _80228_/A sky130_fd_sc_hd__inv_2
X_53166_ _53162_/Y _53163_/X _53165_/X _53166_/Y sky130_fd_sc_hd__a21oi_4
X_41180_ _40717_/X _41181_/A sky130_fd_sc_hd__buf_2
X_50378_ _50383_/A _50378_/B _50378_/Y sky130_fd_sc_hd__nand2_4
X_81198_ _81198_/CLK _81198_/D _49077_/A sky130_fd_sc_hd__dfxtp_4
X_52117_ _52462_/A _52117_/X sky130_fd_sc_hd__buf_2
X_87814_ _87814_/CLK _87814_/D _69734_/A sky130_fd_sc_hd__dfxtp_4
X_80149_ _80157_/A _80149_/B _81687_/D sky130_fd_sc_hd__xnor2_4
X_53097_ _53097_/A _53097_/X sky130_fd_sc_hd__buf_2
X_57974_ _57903_/X _85487_/Q _57962_/X _57974_/X sky130_fd_sc_hd__o21a_4
X_59713_ _59713_/A _59713_/Y sky130_fd_sc_hd__inv_2
X_52048_ _85899_/Q _52013_/X _52047_/Y _52048_/Y sky130_fd_sc_hd__o21ai_4
X_56925_ _55218_/Y _56924_/X _56649_/X _56927_/A sky130_fd_sc_hd__a21o_4
X_87745_ _87748_/CLK _87745_/D _87745_/Q sky130_fd_sc_hd__dfxtp_4
X_72971_ _72968_/X _72969_/Y _72970_/X _72971_/Y sky130_fd_sc_hd__a21oi_4
X_84957_ _84869_/CLK _57671_/Y _84957_/Q sky130_fd_sc_hd__dfxtp_4
X_74710_ _74711_/A _74710_/Y sky130_fd_sc_hd__inv_2
X_71922_ _71920_/Y _57270_/X _71921_/Y _83328_/D sky130_fd_sc_hd__a21o_4
X_59644_ _59797_/B _59651_/B sky130_fd_sc_hd__inv_2
X_83908_ _83905_/CLK _83908_/D _81980_/D sky130_fd_sc_hd__dfxtp_4
X_44870_ _45612_/A _45297_/A sky130_fd_sc_hd__buf_2
X_56856_ _83335_/Q _56856_/Y sky130_fd_sc_hd__inv_2
X_75690_ _75678_/A _75677_/Y _75690_/Y sky130_fd_sc_hd__nor2_4
X_87676_ _87675_/CLK _42871_/X _67118_/B sky130_fd_sc_hd__dfxtp_4
X_84888_ _84888_/CLK _84888_/D _84888_/Q sky130_fd_sc_hd__dfxtp_4
X_43821_ _43821_/A _43821_/Y sky130_fd_sc_hd__inv_2
X_55807_ _55804_/X _55806_/X _44111_/X _55807_/X sky130_fd_sc_hd__a21o_4
X_86627_ _86627_/CLK _86627_/D _58132_/A sky130_fd_sc_hd__dfxtp_4
X_74641_ _74685_/C _74641_/X sky130_fd_sc_hd__buf_2
X_71853_ _70534_/Y _71857_/B _71851_/X _71857_/D _71853_/Y sky130_fd_sc_hd__nor4_4
X_59575_ _60639_/A _60620_/B _60620_/C _59575_/Y sky130_fd_sc_hd__nand3_4
X_83839_ _83835_/CLK _70201_/X _74789_/C sky130_fd_sc_hd__dfxtp_4
X_56787_ _56755_/X _56787_/X sky130_fd_sc_hd__buf_2
X_53999_ _53996_/Y _53982_/X _53998_/Y _53999_/Y sky130_fd_sc_hd__a21boi_4
X_46540_ _46531_/A _50854_/B _46540_/Y sky130_fd_sc_hd__nand2_4
X_70804_ _70804_/A _70810_/A sky130_fd_sc_hd__buf_2
X_58526_ _58526_/A _58526_/Y sky130_fd_sc_hd__inv_2
X_77360_ _77360_/A _77354_/X _77360_/C _77361_/A sky130_fd_sc_hd__nand3_4
X_43752_ _43752_/A _43752_/X sky130_fd_sc_hd__buf_2
X_55738_ _55235_/A _55738_/B _55738_/X sky130_fd_sc_hd__and2_4
X_74572_ _45067_/A _74568_/X _74571_/X _83031_/D sky130_fd_sc_hd__o21ai_4
X_86558_ _86558_/CLK _48197_/Y _86558_/Q sky130_fd_sc_hd__dfxtp_4
X_40964_ _40964_/A _40964_/X sky130_fd_sc_hd__buf_2
X_71784_ _71783_/Y _71784_/X sky130_fd_sc_hd__buf_2
X_76311_ _76311_/A _76310_/Y _76312_/B sky130_fd_sc_hd__xnor2_4
X_42703_ _41121_/X _42695_/X _68403_/B _42696_/X _42703_/X sky130_fd_sc_hd__a2bb2o_4
X_73523_ _73524_/B _73524_/C _73522_/X _73523_/X sky130_fd_sc_hd__a21o_4
X_85509_ _86733_/CLK _54080_/Y _85509_/Q sky130_fd_sc_hd__dfxtp_4
X_46471_ _46471_/A _51330_/A sky130_fd_sc_hd__buf_2
X_70735_ _71263_/D _70735_/X sky130_fd_sc_hd__buf_2
X_58457_ _58457_/A _58474_/B _58457_/Y sky130_fd_sc_hd__nor2_4
X_77291_ _81926_/Q _82182_/D _77291_/X sky130_fd_sc_hd__xor2_4
X_43683_ _40787_/A _43659_/X _69622_/B _43661_/X _43683_/X sky130_fd_sc_hd__a2bb2o_4
X_55669_ _55669_/A _55289_/X _55670_/B sky130_fd_sc_hd__and2_4
X_86489_ _85879_/CLK _48753_/Y _65551_/B sky130_fd_sc_hd__dfxtp_4
X_40895_ _40870_/X _40871_/X _40894_/X _69888_/B _40867_/X _40895_/Y
+ sky130_fd_sc_hd__o32ai_4
X_48210_ _48204_/X _50264_/B _48210_/Y sky130_fd_sc_hd__nand2_4
X_79030_ _82827_/Q _82539_/Q _79031_/B sky130_fd_sc_hd__xnor2_4
X_45422_ _45422_/A _45422_/Y sky130_fd_sc_hd__inv_2
X_57408_ _57470_/B _57408_/X sky130_fd_sc_hd__buf_2
X_88228_ _88232_/CLK _88228_/D _67707_/B sky130_fd_sc_hd__dfxtp_4
X_76242_ _76240_/Y _76211_/Y _76241_/X _76242_/Y sky130_fd_sc_hd__o21ai_4
X_42634_ _42634_/A _42634_/X sky130_fd_sc_hd__buf_2
X_49190_ _49190_/A _49161_/B _49190_/Y sky130_fd_sc_hd__nor2_4
X_73454_ _73448_/X _73453_/X _73383_/X _73457_/A sky130_fd_sc_hd__a21o_4
X_70666_ _70410_/Y _70667_/A sky130_fd_sc_hd__buf_2
X_58388_ _58328_/A _58388_/X sky130_fd_sc_hd__buf_2
X_48141_ _48141_/A _50383_/B sky130_fd_sc_hd__buf_2
X_72405_ _72405_/A _72428_/B _72405_/Y sky130_fd_sc_hd__nor2_4
X_45353_ _45342_/X _45349_/Y _45352_/Y _45353_/Y sky130_fd_sc_hd__a21oi_4
X_57339_ _57338_/Y _57290_/A _44039_/X _57339_/X sky130_fd_sc_hd__o21a_4
X_76173_ _76171_/A _76171_/B _76175_/A sky130_fd_sc_hd__nand2_4
X_88159_ _88164_/CLK _88159_/D _67826_/B sky130_fd_sc_hd__dfxtp_4
X_42565_ _42554_/X _42547_/X _40810_/X _42564_/Y _42556_/X _42565_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73385_ _72880_/A _73385_/X sky130_fd_sc_hd__buf_2
X_70597_ DATA_TO_HASH[6] _70768_/A sky130_fd_sc_hd__buf_2
X_44304_ _44313_/A _43987_/A _46228_/A _44304_/Y sky130_fd_sc_hd__nand3_4
X_75124_ _80678_/Q _75124_/B _75124_/X sky130_fd_sc_hd__or2_4
Xclkbuf_10_470_0_CLK clkbuf_9_235_0_CLK/X _85447_/CLK sky130_fd_sc_hd__clkbuf_1
X_41516_ _41489_/X _41490_/X _41515_/X _88200_/Q _41474_/X _41517_/A
+ sky130_fd_sc_hd__o32ai_4
X_72336_ _72336_/A _72348_/B _72336_/Y sky130_fd_sc_hd__nor2_4
X_48072_ _57605_/B _48073_/B sky130_fd_sc_hd__buf_2
X_60350_ _60350_/A _60350_/Y sky130_fd_sc_hd__inv_2
X_45284_ _45284_/A _45284_/X sky130_fd_sc_hd__buf_2
X_42496_ _42574_/A _42496_/X sky130_fd_sc_hd__buf_2
X_47023_ _83046_/Q _47023_/Y sky130_fd_sc_hd__inv_2
X_59009_ _58918_/X _59006_/Y _59008_/Y _58959_/X _58923_/X _59009_/X
+ sky130_fd_sc_hd__o32a_4
X_44235_ _72881_/A _44235_/X sky130_fd_sc_hd__buf_2
X_75055_ _75062_/A _75062_/B _75055_/Y sky130_fd_sc_hd__xnor2_4
X_79932_ _79932_/A _79932_/B _79932_/Y sky130_fd_sc_hd__xnor2_4
X_41447_ _41446_/Y _41447_/X sky130_fd_sc_hd__buf_2
X_60281_ _60281_/A _60284_/A sky130_fd_sc_hd__inv_2
X_72267_ _72240_/X _85685_/Q _72241_/X _72267_/X sky130_fd_sc_hd__o21a_4
X_62020_ _61787_/X _62020_/X sky130_fd_sc_hd__buf_2
X_74006_ _41947_/Y _56182_/X _73962_/X _74005_/Y _74006_/X sky130_fd_sc_hd__a211o_4
X_71218_ _48628_/B _71216_/X _71217_/Y _71218_/Y sky130_fd_sc_hd__o21ai_4
X_44166_ _64619_/A _57736_/A _58834_/A _44265_/D _44166_/Y sky130_fd_sc_hd__nor4_4
X_79863_ _79863_/A _79863_/B _79864_/B sky130_fd_sc_hd__xor2_4
X_41378_ _41378_/A _41378_/Y sky130_fd_sc_hd__inv_2
X_72198_ _72143_/X _85371_/Q _72197_/X _72198_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_485_0_CLK clkbuf_9_242_0_CLK/X _84797_/CLK sky130_fd_sc_hd__clkbuf_1
X_43117_ _87569_/Q _43117_/Y sky130_fd_sc_hd__inv_2
X_78814_ _78814_/A _82547_/Q _79122_/B sky130_fd_sc_hd__nand2_4
X_40329_ _40402_/A _81184_/Q _40329_/X sky130_fd_sc_hd__or2_4
X_71149_ _70611_/X _71160_/D sky130_fd_sc_hd__buf_2
X_48974_ _48964_/A _52307_/B _48974_/Y sky130_fd_sc_hd__nand2_4
X_44097_ _44096_/X _44097_/X sky130_fd_sc_hd__buf_2
X_79794_ _79794_/A _79794_/B _79794_/Y sky130_fd_sc_hd__nand2_4
X_47925_ _66024_/B _47897_/X _47924_/Y _47925_/Y sky130_fd_sc_hd__o21ai_4
X_43048_ _87595_/Q _43048_/Y sky130_fd_sc_hd__inv_2
X_78745_ _78745_/A _78745_/Y sky130_fd_sc_hd__inv_2
X_63971_ _61954_/X _63955_/X _63905_/C _64033_/D _63971_/Y sky130_fd_sc_hd__nand4_4
X_75957_ _75957_/A _75957_/B _75957_/Y sky130_fd_sc_hd__nand2_4
X_65710_ _65710_/A _65710_/B _65710_/Y sky130_fd_sc_hd__nand2_4
X_62922_ _62920_/X _62893_/X _62921_/Y _84370_/D sky130_fd_sc_hd__a21oi_4
X_74908_ _81130_/D _80842_/Q _74908_/Y sky130_fd_sc_hd__nand2_4
X_47856_ _65935_/B _47840_/X _47855_/Y _47856_/Y sky130_fd_sc_hd__o21ai_4
X_66690_ _87950_/Q _66639_/X _66688_/X _66689_/X _66690_/X sky130_fd_sc_hd__a211o_4
X_78676_ _82522_/Q _82778_/D _78676_/X sky130_fd_sc_hd__xor2_4
X_75888_ _75888_/A _75580_/Y _75888_/Y sky130_fd_sc_hd__nand2_4
X_46807_ _86701_/Q _46767_/X _46806_/Y _46807_/Y sky130_fd_sc_hd__o21ai_4
X_65641_ _65638_/X _85587_/Q _65470_/X _65640_/X _65641_/X sky130_fd_sc_hd__a211o_4
X_77627_ _77627_/A _77626_/Y _82204_/D sky130_fd_sc_hd__xor2_4
X_62853_ _62894_/A _62852_/X _75907_/B _62853_/Y sky130_fd_sc_hd__nor3_4
X_74839_ _74844_/A _46121_/A _74839_/Y sky130_fd_sc_hd__nand2_4
X_47787_ _47787_/A _47788_/A sky130_fd_sc_hd__inv_2
X_44999_ _56303_/C _44979_/X _44926_/X _44999_/X sky130_fd_sc_hd__o21a_4
X_49526_ _49546_/A _46899_/X _49526_/Y sky130_fd_sc_hd__nand2_4
X_61804_ _59721_/X _61823_/A sky130_fd_sc_hd__buf_2
X_68360_ _65117_/A _68360_/X sky130_fd_sc_hd__buf_2
X_46738_ _46734_/Y _46704_/X _46737_/X _86709_/D sky130_fd_sc_hd__a21oi_4
X_65572_ _65516_/X _64855_/Y _65571_/Y _65572_/Y sky130_fd_sc_hd__o21ai_4
X_77558_ _77553_/X _77556_/Y _77558_/C _77559_/B sky130_fd_sc_hd__nand3_4
X_62784_ _57664_/X _62749_/X _62768_/X _62759_/X _62783_/X _62784_/Y
+ sky130_fd_sc_hd__a41oi_4
X_67311_ _66953_/X _67311_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_423_0_CLK clkbuf_9_211_0_CLK/X _82462_/CLK sky130_fd_sc_hd__clkbuf_1
X_64523_ _64234_/A _64523_/B _58201_/A _64523_/D _64523_/X sky130_fd_sc_hd__and4_4
X_76509_ _76510_/A _76510_/C _76510_/B _76509_/X sky130_fd_sc_hd__a21o_4
X_49457_ _49455_/Y _49434_/X _49456_/X _86384_/D sky130_fd_sc_hd__a21oi_4
X_61735_ _61704_/Y _61736_/A sky130_fd_sc_hd__buf_2
X_68291_ _67800_/X _67802_/X _68283_/X _68291_/Y sky130_fd_sc_hd__a21oi_4
X_46669_ _54298_/D _51777_/D sky130_fd_sc_hd__buf_2
X_77489_ _77488_/Y _77489_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_4_15_1_CLK clkbuf_4_15_0_CLK/X clkbuf_5_30_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_48408_ _48557_/A _52119_/B _48408_/Y sky130_fd_sc_hd__nand2_4
X_67242_ _87351_/Q _67239_/X _67240_/X _67241_/X _67242_/X sky130_fd_sc_hd__a211o_4
X_79228_ _84791_/Q _84111_/Q _79230_/A sky130_fd_sc_hd__or2_4
X_64454_ _64454_/A _64454_/B _64454_/Y sky130_fd_sc_hd__nor2_4
X_49388_ _49415_/A _49388_/X sky130_fd_sc_hd__buf_2
X_61666_ _61666_/A _61653_/X _61654_/X _61639_/X _61666_/Y sky130_fd_sc_hd__nand4_4
X_63405_ _62851_/A _63468_/A sky130_fd_sc_hd__buf_2
X_60617_ _61078_/B _61075_/B sky130_fd_sc_hd__buf_2
X_48339_ _48336_/Y _48322_/X _48338_/Y _48339_/Y sky130_fd_sc_hd__a21boi_4
X_67173_ _67149_/A _88186_/Q _67173_/X sky130_fd_sc_hd__and2_4
X_79159_ _79158_/B _79159_/Y sky130_fd_sc_hd__inv_2
X_64385_ _64376_/X _64378_/X _64379_/X _64383_/Y _64384_/X _64385_/X
+ sky130_fd_sc_hd__o41a_4
X_61597_ _61597_/A _61611_/B _61611_/C _61572_/D _61597_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_10_438_0_CLK clkbuf_9_219_0_CLK/X _81227_/CLK sky130_fd_sc_hd__clkbuf_1
X_66124_ _66122_/Y _66065_/X _66123_/X _84155_/D sky130_fd_sc_hd__a21o_4
X_51350_ _51350_/A _51350_/B _51350_/Y sky130_fd_sc_hd__nand2_4
X_63336_ _63334_/Y _63335_/X _63317_/X _63336_/X sky130_fd_sc_hd__a21o_4
X_82170_ _84166_/CLK _84162_/Q _82170_/Q sky130_fd_sc_hd__dfxtp_4
X_60548_ _60413_/X _60455_/Y _60571_/B _60546_/Y _60547_/Y _60548_/Y
+ sky130_fd_sc_hd__a41oi_4
X_50301_ _50298_/Y _50299_/X _50300_/Y _50301_/Y sky130_fd_sc_hd__a21boi_4
X_81121_ _81121_/CLK _79892_/Y _81121_/Q sky130_fd_sc_hd__dfxtp_4
X_66055_ _66054_/X _66055_/B _66055_/X sky130_fd_sc_hd__and2_4
X_51281_ _64860_/B _51259_/X _51280_/Y _51281_/Y sky130_fd_sc_hd__o21ai_4
X_63267_ _58459_/Y _63316_/B _63295_/C _63267_/D _63267_/X sky130_fd_sc_hd__or4_4
X_60479_ _60572_/A _60572_/B _60572_/C _60479_/Y sky130_fd_sc_hd__nand3_4
X_53020_ _53018_/Y _53001_/X _53019_/X _53020_/Y sky130_fd_sc_hd__a21oi_4
X_65006_ _65005_/X _86418_/Q _65006_/X sky130_fd_sc_hd__and2_4
X_50232_ _51737_/A _50232_/B _50232_/Y sky130_fd_sc_hd__nand2_4
X_62218_ _62218_/A _62618_/C sky130_fd_sc_hd__buf_2
X_81052_ _84276_/CLK _81052_/D _81052_/Q sky130_fd_sc_hd__dfxtp_4
X_63198_ _63198_/A _63170_/X _63161_/C _63149_/X _63198_/X sky130_fd_sc_hd__or4_4
X_80003_ _79997_/X _80003_/B _80003_/Y sky130_fd_sc_hd__nand2_4
X_69814_ _69814_/A _70012_/A sky130_fd_sc_hd__buf_2
X_50163_ _50064_/A _50169_/A sky130_fd_sc_hd__buf_2
X_62149_ _61665_/B _62149_/B _62149_/C _61749_/B _62153_/B sky130_fd_sc_hd__nand4_4
X_85860_ _85859_/CLK _85860_/D _85860_/Q sky130_fd_sc_hd__dfxtp_4
X_84811_ _85955_/CLK _84811_/D _84811_/Q sky130_fd_sc_hd__dfxtp_4
X_69745_ _83900_/Q _69696_/X _69744_/X _83900_/D sky130_fd_sc_hd__a21bo_4
X_50094_ _50091_/Y _50092_/X _50093_/X _50094_/Y sky130_fd_sc_hd__a21oi_4
X_54971_ _54253_/A _54971_/X sky130_fd_sc_hd__buf_2
X_66957_ _88387_/Q _66954_/X _66955_/X _66956_/X _66957_/X sky130_fd_sc_hd__a211o_4
X_85791_ _83685_/CLK _52589_/Y _85791_/Q sky130_fd_sc_hd__dfxtp_4
X_56710_ _56661_/C _56721_/D sky130_fd_sc_hd__buf_2
X_87530_ _87533_/CLK _43224_/X _87530_/Q sky130_fd_sc_hd__dfxtp_4
X_53922_ _53956_/A _53951_/A sky130_fd_sc_hd__buf_2
X_65908_ _65807_/A _65908_/B _65908_/X sky130_fd_sc_hd__and2_4
X_84742_ _83766_/CLK _84742_/D _84742_/Q sky130_fd_sc_hd__dfxtp_4
X_57690_ _58094_/A _57896_/A sky130_fd_sc_hd__buf_2
X_81954_ _81954_/CLK _83882_/Q _77872_/B sky130_fd_sc_hd__dfxtp_4
X_69676_ _69687_/A _69676_/B _69676_/Y sky130_fd_sc_hd__nor2_4
X_66888_ _87878_/Q _66816_/X _66794_/X _66887_/X _66888_/X sky130_fd_sc_hd__a211o_4
X_56641_ _56636_/X _56639_/X _85140_/Q _56753_/A _56641_/X sky130_fd_sc_hd__a2bb2o_4
X_80905_ _83932_/CLK _84081_/Q _75630_/A sky130_fd_sc_hd__dfxtp_4
X_68627_ _68604_/A _68627_/B _68627_/X sky130_fd_sc_hd__and2_4
X_87461_ _87149_/CLK _87461_/D _87461_/Q sky130_fd_sc_hd__dfxtp_4
X_53853_ _85555_/Q _53846_/X _53852_/Y _53853_/Y sky130_fd_sc_hd__o21ai_4
X_65839_ _65319_/A _86502_/Q _65839_/X sky130_fd_sc_hd__and2_4
X_84673_ _84671_/CLK _84673_/D _60032_/C sky130_fd_sc_hd__dfxtp_4
X_81885_ _81839_/CLK _78076_/X _81885_/Q sky130_fd_sc_hd__dfxtp_4
X_86412_ _86414_/CLK _49313_/Y _65152_/B sky130_fd_sc_hd__dfxtp_4
X_52804_ _85751_/Q _52792_/X _52803_/Y _52804_/Y sky130_fd_sc_hd__o21ai_4
X_59360_ _59238_/X _59360_/B _59360_/Y sky130_fd_sc_hd__nor2_4
X_83624_ _83310_/CLK _71053_/Y _83624_/Q sky130_fd_sc_hd__dfxtp_4
X_56572_ _56552_/Y _56572_/X sky130_fd_sc_hd__buf_2
X_80836_ _81125_/CLK _80868_/Q _74854_/B sky130_fd_sc_hd__dfxtp_4
X_68558_ _68429_/A _68558_/X sky130_fd_sc_hd__buf_2
X_87392_ _87646_/CLK _87392_/D _87392_/Q sky130_fd_sc_hd__dfxtp_4
X_53784_ _53729_/A _53784_/X sky130_fd_sc_hd__buf_2
X_50996_ _50973_/X _50985_/B _50985_/C _46810_/X _50996_/X sky130_fd_sc_hd__and4_4
X_58311_ _84881_/Q _58314_/A sky130_fd_sc_hd__inv_2
Xclkbuf_8_50_0_CLK clkbuf_8_51_0_CLK/A clkbuf_8_50_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_55523_ _55458_/X _55523_/X sky130_fd_sc_hd__buf_2
X_86343_ _82381_/CLK _86343_/D _86343_/Q sky130_fd_sc_hd__dfxtp_4
X_67509_ _67460_/A _87724_/Q _67509_/X sky130_fd_sc_hd__and2_4
X_52735_ _52729_/X _52724_/B _52746_/C _52735_/D _52735_/X sky130_fd_sc_hd__and4_4
X_59291_ _84753_/Q _59291_/Y sky130_fd_sc_hd__inv_2
X_83555_ _83556_/CLK _83555_/D _47899_/A sky130_fd_sc_hd__dfxtp_4
X_80767_ _80740_/CLK _75535_/Y _81143_/D sky130_fd_sc_hd__dfxtp_4
X_68489_ _83973_/Q _68462_/X _68488_/X _83973_/D sky130_fd_sc_hd__a21bo_4
X_70520_ _70504_/A _70526_/A sky130_fd_sc_hd__buf_2
X_58242_ _44184_/X _58510_/A sky130_fd_sc_hd__buf_2
X_82506_ _82498_/CLK _82506_/D _82506_/Q sky130_fd_sc_hd__dfxtp_4
X_55454_ _55342_/X _55454_/X sky130_fd_sc_hd__buf_2
X_86274_ _85955_/CLK _86274_/D _72475_/B sky130_fd_sc_hd__dfxtp_4
X_52666_ _52664_/Y _52647_/X _52665_/X _52666_/Y sky130_fd_sc_hd__a21oi_4
X_40680_ _40829_/A _82864_/Q _40680_/X sky130_fd_sc_hd__or2_4
X_83486_ _83482_/CLK _83486_/D _83486_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_702 sky130_fd_sc_hd__decap_3
X_80698_ _81048_/CLK _80730_/Q _75424_/A sky130_fd_sc_hd__dfxtp_4
XPHY_713 sky130_fd_sc_hd__decap_3
X_88013_ _87766_/CLK _42145_/X _88013_/Q sky130_fd_sc_hd__dfxtp_4
X_54405_ _54322_/A _54425_/A sky130_fd_sc_hd__buf_2
X_85225_ _85192_/CLK _56353_/Y _55764_/B sky130_fd_sc_hd__dfxtp_4
X_51617_ _51617_/A _53141_/B _51617_/Y sky130_fd_sc_hd__nand2_4
X_70451_ _50306_/B _70421_/Y _70450_/Y _70451_/Y sky130_fd_sc_hd__o21ai_4
X_58173_ _63081_/A _64282_/A sky130_fd_sc_hd__buf_2
X_82437_ _82443_/CLK _82437_/D _82437_/Q sky130_fd_sc_hd__dfxtp_4
X_55385_ _55384_/Y _55375_/Y _55382_/A _56719_/B sky130_fd_sc_hd__o21ai_4
X_52597_ _85789_/Q _52575_/X _52596_/Y _52597_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_8_65_0_CLK clkbuf_8_65_0_CLK/A clkbuf_8_65_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_57124_ _56972_/Y _56664_/Y _57221_/A _57123_/Y _57124_/X sky130_fd_sc_hd__a211o_4
X_42350_ _42417_/A _42350_/X sky130_fd_sc_hd__buf_2
X_54336_ _54332_/A _52645_/B _54336_/Y sky130_fd_sc_hd__nand2_4
X_73170_ _73156_/Y _73169_/X _73170_/Y sky130_fd_sc_hd__xnor2_4
X_85156_ _85156_/CLK _56541_/Y _55724_/B sky130_fd_sc_hd__dfxtp_4
X_51548_ _51553_/A _51553_/B _51533_/C _53074_/D _51548_/X sky130_fd_sc_hd__and4_4
X_70382_ _70382_/A _70994_/A sky130_fd_sc_hd__buf_2
X_82368_ _82368_/CLK _82368_/D _82368_/Q sky130_fd_sc_hd__dfxtp_4
X_41301_ _41290_/X _82910_/Q _41300_/X _41301_/Y sky130_fd_sc_hd__o21ai_4
X_72121_ _59346_/X _85345_/Q _72120_/X _72121_/X sky130_fd_sc_hd__o21a_4
X_84107_ _82425_/CLK _84107_/D _82723_/D sky130_fd_sc_hd__dfxtp_4
X_57055_ _57055_/A _56849_/X _56985_/D _57055_/Y sky130_fd_sc_hd__nor3_4
X_81319_ _84079_/CLK _76226_/X _81727_/D sky130_fd_sc_hd__dfxtp_4
X_54267_ _54295_/A _54288_/A sky130_fd_sc_hd__buf_2
X_42281_ _42281_/A _42281_/Y sky130_fd_sc_hd__inv_2
X_85087_ _85152_/CLK _57101_/X _45422_/A sky130_fd_sc_hd__dfxtp_4
X_51479_ _51473_/A _51494_/B _51494_/C _53003_/D _51479_/X sky130_fd_sc_hd__and4_4
X_82299_ _82299_/CLK _82299_/D _82299_/Q sky130_fd_sc_hd__dfxtp_4
X_44020_ _44020_/A _64717_/A sky130_fd_sc_hd__buf_2
X_56006_ _45765_/A _56017_/B sky130_fd_sc_hd__buf_2
X_41232_ _41062_/B _41223_/B _41232_/X sky130_fd_sc_hd__or2_4
X_53218_ _53214_/Y _53215_/X _53217_/X _53218_/Y sky130_fd_sc_hd__a21oi_4
X_72052_ _72052_/A _72053_/A sky130_fd_sc_hd__buf_2
X_84038_ _81160_/CLK _84038_/D _82078_/D sky130_fd_sc_hd__dfxtp_4
X_54198_ _54254_/A _54209_/C sky130_fd_sc_hd__buf_2
X_71003_ _71003_/A _71071_/A sky130_fd_sc_hd__buf_2
X_41163_ _40984_/B _41145_/B _41163_/X sky130_fd_sc_hd__or2_4
X_53149_ _85688_/Q _53146_/X _53148_/Y _53149_/Y sky130_fd_sc_hd__o21ai_4
X_76860_ _76854_/A _76854_/B _76860_/Y sky130_fd_sc_hd__nor2_4
X_75811_ _75811_/A _75810_/Y _75811_/X sky130_fd_sc_hd__and2_4
X_45971_ _44857_/X _44865_/X _40394_/X _66700_/B _44858_/X _45971_/Y
+ sky130_fd_sc_hd__o32ai_4
X_41094_ _41093_/X _41065_/X _69526_/B _41066_/X _41094_/X sky130_fd_sc_hd__a2bb2o_4
X_57957_ _57944_/Y _57758_/X _57951_/X _57956_/X _84937_/D sky130_fd_sc_hd__a22oi_4
X_76791_ _81490_/Q _76806_/A sky130_fd_sc_hd__inv_2
X_85989_ _85990_/CLK _85989_/D _85989_/Q sky130_fd_sc_hd__dfxtp_4
X_47710_ _47710_/A _53203_/D sky130_fd_sc_hd__buf_2
X_78530_ _78519_/A _78519_/B _78510_/Y _78530_/X sky130_fd_sc_hd__o21a_4
X_44922_ _64223_/B _61329_/B sky130_fd_sc_hd__buf_2
X_56908_ _56908_/A _56907_/X _56908_/X sky130_fd_sc_hd__xor2_4
X_87728_ _87472_/CLK _87728_/D _67406_/B sky130_fd_sc_hd__dfxtp_4
X_75742_ _80917_/Q _75742_/Y sky130_fd_sc_hd__inv_2
X_48690_ _48635_/A _48894_/B sky130_fd_sc_hd__buf_2
X_72954_ _44535_/Y _72775_/X _72953_/Y _72969_/C sky130_fd_sc_hd__a21o_4
X_57888_ _72476_/B _86006_/Q _57887_/X _57888_/Y sky130_fd_sc_hd__o21ai_4
X_47641_ _47649_/A _53161_/B _47641_/Y sky130_fd_sc_hd__nand2_4
X_71905_ _74527_/A _71893_/X _71902_/X _71898_/D _71905_/Y sky130_fd_sc_hd__nand4_4
X_59627_ _61755_/A _59628_/A sky130_fd_sc_hd__buf_2
X_78461_ _78461_/A _78458_/Y _78460_/Y _78463_/A sky130_fd_sc_hd__or3_4
X_44853_ _44852_/Y _86919_/D sky130_fd_sc_hd__inv_2
X_56839_ _56838_/Y _56839_/Y sky130_fd_sc_hd__inv_2
X_75673_ _75656_/A _80780_/D _75672_/Y _75673_/Y sky130_fd_sc_hd__a21oi_4
X_87659_ _87653_/CLK _87659_/D _87659_/Q sky130_fd_sc_hd__dfxtp_4
X_72885_ _72869_/Y _72884_/X _72885_/Y sky130_fd_sc_hd__xnor2_4
X_77412_ _77412_/A _77412_/B _77412_/C _77412_/X sky130_fd_sc_hd__or3_4
X_43804_ _41070_/X _43801_/X _69469_/B _43802_/X _87259_/D sky130_fd_sc_hd__a2bb2o_4
X_74624_ _45365_/A _74612_/X _74623_/X _74624_/Y sky130_fd_sc_hd__o21ai_4
X_47572_ _83708_/Q _47572_/Y sky130_fd_sc_hd__inv_2
X_71836_ _71825_/X _58548_/B _71835_/X _83358_/D sky130_fd_sc_hd__a21o_4
X_59558_ _43959_/A _44008_/A _43959_/B _59558_/Y sky130_fd_sc_hd__nand3_4
X_78392_ _78391_/Y _78371_/Y _78375_/C _78394_/C sky130_fd_sc_hd__o21ai_4
X_44784_ _44766_/X _44767_/X _41387_/A _86956_/Q _44768_/X _44784_/Y
+ sky130_fd_sc_hd__o32ai_4
X_41996_ _41996_/A _41996_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_18_0_CLK clkbuf_7_9_0_CLK/X clkbuf_9_37_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_49311_ _65152_/B _49300_/X _49310_/Y _49311_/Y sky130_fd_sc_hd__o21ai_4
X_46523_ _46399_/A _46523_/X sky130_fd_sc_hd__buf_2
X_58509_ _64335_/C _58511_/A sky130_fd_sc_hd__buf_2
X_77343_ _77339_/X _77340_/Y _77342_/Y _77345_/A sky130_fd_sc_hd__a21o_4
X_43735_ _40899_/X _43695_/X _87290_/Q _43696_/X _43735_/X sky130_fd_sc_hd__a2bb2o_4
X_74555_ _46155_/X _74553_/X _56025_/X _74554_/X _74555_/X sky130_fd_sc_hd__a211o_4
X_40947_ _40947_/A _40970_/B sky130_fd_sc_hd__buf_2
X_71767_ _71762_/X _83384_/Q _71766_/X _71767_/X sky130_fd_sc_hd__a21o_4
X_59489_ _64248_/C _63396_/B sky130_fd_sc_hd__buf_2
X_49242_ _64798_/B _49222_/X _49241_/Y _49242_/Y sky130_fd_sc_hd__o21ai_4
X_61520_ _72561_/C _61538_/C sky130_fd_sc_hd__buf_2
X_73506_ _83148_/Q _73437_/X _73505_/Y _73506_/X sky130_fd_sc_hd__a21o_4
X_70718_ _52768_/B _70699_/X _70717_/Y _70718_/Y sky130_fd_sc_hd__o21ai_4
X_46454_ _46444_/Y _46445_/X _46453_/X _46454_/Y sky130_fd_sc_hd__a21oi_4
X_77274_ _77272_/Y _77274_/B _77270_/X _77274_/Y sky130_fd_sc_hd__nand3_4
X_43666_ _40739_/X _43656_/X _74186_/A _43657_/X _87320_/D sky130_fd_sc_hd__a2bb2o_4
X_74486_ _83056_/Q _74474_/X _74485_/Y _74486_/Y sky130_fd_sc_hd__o21ai_4
X_40878_ _40878_/A _46469_/B sky130_fd_sc_hd__buf_2
X_71698_ _71698_/A _71690_/A _71874_/D _71698_/Y sky130_fd_sc_hd__nor3_4
X_79013_ _82825_/Q _82537_/Q _79014_/B sky130_fd_sc_hd__xnor2_4
X_45405_ _61714_/A _61315_/A sky130_fd_sc_hd__buf_2
X_76225_ _76223_/Y _76225_/B _81607_/D sky130_fd_sc_hd__xor2_4
X_42617_ _42616_/Y _87800_/D sky130_fd_sc_hd__inv_2
X_49173_ _49173_/A _50710_/B _49173_/X sky130_fd_sc_hd__and2_4
X_61451_ _61451_/A _61404_/X _61406_/C _61451_/D _61451_/Y sky130_fd_sc_hd__nand4_4
X_73437_ _73193_/A _73437_/X sky130_fd_sc_hd__buf_2
X_46385_ _46385_/A _52480_/B sky130_fd_sc_hd__inv_2
X_70649_ _70719_/A _70639_/B _70642_/X _70638_/X _70649_/Y sky130_fd_sc_hd__nand4_4
X_43597_ _40573_/A _43586_/X _68387_/B _43593_/X _43598_/A sky130_fd_sc_hd__a2bb2o_4
X_48124_ _48142_/A _48335_/B _48124_/Y sky130_fd_sc_hd__nand2_4
X_60402_ _60402_/A _60403_/B sky130_fd_sc_hd__buf_2
X_45336_ _45329_/X _45333_/Y _45335_/Y _45336_/Y sky130_fd_sc_hd__a21oi_4
X_64170_ _64166_/Y _64167_/Y _64168_/Y _64169_/Y _64170_/X sky130_fd_sc_hd__and4_4
X_76156_ _81634_/Q _76155_/X _81602_/D sky130_fd_sc_hd__xor2_4
X_42548_ _42548_/A _42548_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_3_4_1_CLK clkbuf_3_4_0_CLK/X clkbuf_4_9_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_61382_ _61381_/Y _61382_/Y sky130_fd_sc_hd__inv_2
X_73368_ _73364_/X _73365_/Y _73367_/X _73368_/Y sky130_fd_sc_hd__a21oi_4
X_63121_ _63097_/A _64334_/B _63108_/C _63121_/D _63121_/X sky130_fd_sc_hd__and4_4
X_75107_ _75107_/A _75107_/B _75107_/Y sky130_fd_sc_hd__xnor2_4
X_60333_ _60256_/X _60285_/A _60330_/Y _60331_/Y _60332_/Y _60333_/Y
+ sky130_fd_sc_hd__a41oi_4
X_72319_ _72366_/A _86289_/Q _72319_/Y sky130_fd_sc_hd__nor2_4
X_48055_ _48734_/A _48055_/X sky130_fd_sc_hd__buf_2
X_45267_ _85193_/Q _45252_/X _45266_/X _45267_/Y sky130_fd_sc_hd__o21ai_4
X_76087_ _76077_/Y _76080_/X _76082_/A _76087_/Y sky130_fd_sc_hd__a21boi_4
X_42479_ _42460_/X _40632_/Y _42477_/X _68567_/B _42463_/X _42479_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73299_ _73299_/A _73003_/B _73299_/Y sky130_fd_sc_hd__nor2_4
X_47006_ _83048_/Q _47006_/Y sky130_fd_sc_hd__inv_2
X_44218_ _44216_/X _44217_/X _44153_/X _44218_/X sky130_fd_sc_hd__a21o_4
X_79915_ _79915_/A _79915_/B _80262_/B sky130_fd_sc_hd__nand2_4
X_63052_ _63047_/Y _63049_/X _63050_/X _63051_/X _63020_/X _63052_/Y
+ sky130_fd_sc_hd__o41ai_4
X_75038_ _81149_/D _75040_/B _75038_/X sky130_fd_sc_hd__or2_4
X_60264_ _60207_/Y _60264_/Y sky130_fd_sc_hd__inv_2
X_45198_ _45272_/A _45199_/B sky130_fd_sc_hd__buf_2
X_62003_ _62001_/Y _61959_/X _62002_/Y _84440_/D sky130_fd_sc_hd__a21oi_4
X_44149_ _44149_/A _44149_/X sky130_fd_sc_hd__buf_2
X_67860_ _67909_/A _67860_/B _67860_/X sky130_fd_sc_hd__and2_4
X_79846_ _79846_/A _79846_/B _79860_/B sky130_fd_sc_hd__xor2_4
X_60195_ _60179_/A _62737_/A sky130_fd_sc_hd__buf_2
X_66811_ _87369_/Q _66762_/X _66764_/X _66810_/X _66811_/X sky130_fd_sc_hd__a211o_4
X_48957_ _86458_/Q _48952_/X _48956_/Y _48957_/Y sky130_fd_sc_hd__o21ai_4
X_67791_ _87148_/Q _67788_/X _67789_/X _67790_/X _67791_/X sky130_fd_sc_hd__a211o_4
X_79777_ _79790_/B _79776_/Y _79777_/X sky130_fd_sc_hd__xor2_4
X_76989_ _76989_/A _62397_/C _76989_/X sky130_fd_sc_hd__xor2_4
X_69530_ _81381_/D _69504_/X _69529_/X _83917_/D sky130_fd_sc_hd__a21bo_4
X_47908_ _47887_/A _48212_/A _47908_/X sky130_fd_sc_hd__and2_4
X_66742_ _88396_/Q _66715_/X _66717_/X _66741_/X _66742_/X sky130_fd_sc_hd__a211o_4
X_78728_ _78728_/A _78732_/A sky130_fd_sc_hd__inv_2
X_63954_ _63947_/Y _63949_/Y _63951_/Y _63954_/D _63954_/X sky130_fd_sc_hd__and4_4
X_48888_ _48887_/Y _48889_/B sky130_fd_sc_hd__buf_2
X_62905_ _58495_/A _62658_/A _60197_/C _60202_/A _62905_/Y sky130_fd_sc_hd__nand4_4
X_69461_ _69461_/A _69461_/B _69461_/Y sky130_fd_sc_hd__nand2_4
X_47839_ _47838_/X _47840_/A sky130_fd_sc_hd__buf_2
X_66673_ _45920_/A _66673_/X sky130_fd_sc_hd__buf_2
X_78659_ _82810_/Q _78663_/A sky130_fd_sc_hd__inv_2
X_63885_ _61437_/B _63920_/B _63840_/C _63920_/D _63885_/Y sky130_fd_sc_hd__nand4_4
X_68412_ _68376_/X _66524_/B _68401_/Y _68411_/Y _68412_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_362_0_CLK clkbuf_9_181_0_CLK/X _84926_/CLK sky130_fd_sc_hd__clkbuf_1
X_65624_ _65777_/A _85876_/Q _65624_/X sky130_fd_sc_hd__and2_4
X_50850_ _50845_/A _50850_/B _50850_/Y sky130_fd_sc_hd__nand2_4
X_62836_ _62789_/A _59419_/A _62848_/C _62880_/D _62836_/X sky130_fd_sc_hd__and4_4
X_69392_ _81391_/D _69367_/X _69391_/X _83927_/D sky130_fd_sc_hd__a21bo_4
X_81670_ _81582_/CLK _79967_/Y _81670_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_992_0_CLK clkbuf_9_496_0_CLK/X _86210_/CLK sky130_fd_sc_hd__clkbuf_1
X_49509_ _86374_/Q _49496_/X _49508_/Y _49509_/Y sky130_fd_sc_hd__o21ai_4
X_80621_ _80622_/B _80622_/A _82272_/D sky130_fd_sc_hd__xor2_4
X_68343_ _64898_/A _68343_/B _68343_/X sky130_fd_sc_hd__and2_4
X_65555_ _65524_/X _83073_/Q _65391_/X _65554_/X _65556_/C sky130_fd_sc_hd__a211o_4
X_50781_ _50777_/A _50781_/B _50781_/Y sky130_fd_sc_hd__nand2_4
X_62767_ _62765_/X _62721_/X _62766_/Y _62767_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_483_0_CLK clkbuf_9_483_0_CLK/A clkbuf_9_483_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_52520_ _51330_/A _52509_/B _52498_/C _52520_/X sky130_fd_sc_hd__and3_4
X_64506_ _58976_/A _61085_/X _64505_/Y _64506_/Y sky130_fd_sc_hd__o21ai_4
X_83340_ _83362_/CLK _71886_/X _83340_/Q sky130_fd_sc_hd__dfxtp_4
X_61718_ _61704_/Y _61719_/A sky130_fd_sc_hd__buf_2
X_80552_ _80542_/A _80527_/Y _80537_/X _80541_/B _80552_/X sky130_fd_sc_hd__o22a_4
X_68274_ _68272_/X _67674_/Y _68268_/X _68273_/Y _68274_/X sky130_fd_sc_hd__a211o_4
X_65486_ _65486_/A _65667_/A sky130_fd_sc_hd__buf_2
X_62698_ _62696_/X _62652_/X _62697_/Y _62698_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_377_0_CLK clkbuf_9_188_0_CLK/X _83716_/CLK sky130_fd_sc_hd__clkbuf_1
X_67225_ _66572_/X _67226_/A sky130_fd_sc_hd__buf_2
X_52451_ _52449_/Y _52415_/X _52450_/X _52451_/Y sky130_fd_sc_hd__a21oi_4
X_64437_ _61101_/A _64515_/C sky130_fd_sc_hd__buf_2
X_83271_ _83627_/CLK _72249_/Y _72236_/A sky130_fd_sc_hd__dfxtp_4
X_61649_ _61636_/A _61649_/B _61682_/C _61649_/Y sky130_fd_sc_hd__nand3_4
X_80483_ _59159_/A _84156_/Q _80494_/A sky130_fd_sc_hd__xor2_4
X_85010_ _85041_/CLK _57407_/X _55483_/A sky130_fd_sc_hd__dfxtp_4
X_51402_ _51128_/A _51402_/X sky130_fd_sc_hd__buf_2
X_82222_ _81883_/CLK _82254_/Q _77392_/A sky130_fd_sc_hd__dfxtp_4
X_55170_ _85036_/Q _55157_/X _55168_/X _55169_/X _55170_/X sky130_fd_sc_hd__a211o_4
X_67156_ _66915_/A _67156_/X sky130_fd_sc_hd__buf_2
X_52382_ _52380_/Y _52364_/X _52381_/X _85834_/D sky130_fd_sc_hd__a21oi_4
X_64368_ _64336_/A _84820_/Q _64323_/X _64368_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_9_498_0_CLK clkbuf_9_499_0_CLK/A clkbuf_9_498_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_54121_ _54134_/A _54121_/B _54121_/Y sky130_fd_sc_hd__nand2_4
X_66107_ _65045_/A _66164_/B sky130_fd_sc_hd__buf_2
X_51333_ _50063_/A _51790_/A sky130_fd_sc_hd__buf_2
X_63319_ _79212_/A _63310_/X _63318_/X _63319_/Y sky130_fd_sc_hd__o21ai_4
X_82153_ _84175_/CLK _84145_/Q _82153_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_300_0_CLK clkbuf_9_150_0_CLK/X _84308_/CLK sky130_fd_sc_hd__clkbuf_1
X_67087_ _67087_/A _67087_/B _67087_/X sky130_fd_sc_hd__and2_4
X_64299_ _64292_/Y _64298_/X _64269_/X _64299_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_10_930_0_CLK clkbuf_9_465_0_CLK/X _87288_/CLK sky130_fd_sc_hd__clkbuf_1
X_81104_ _81104_/CLK _79709_/X _81104_/Q sky130_fd_sc_hd__dfxtp_4
X_54052_ _46507_/A _54043_/B _51749_/X _54052_/X sky130_fd_sc_hd__and3_4
X_66038_ _65876_/X _85624_/Q _65976_/X _66037_/X _66038_/X sky130_fd_sc_hd__a211o_4
X_51264_ _52139_/A _51265_/A sky130_fd_sc_hd__buf_2
X_86961_ _88232_/CLK _44777_/X _86961_/Q sky130_fd_sc_hd__dfxtp_4
X_82084_ _82084_/CLK _82084_/D _77017_/A sky130_fd_sc_hd__dfxtp_4
X_53003_ _53019_/A _52997_/B _52997_/C _53003_/D _53003_/X sky130_fd_sc_hd__and4_4
Xclkbuf_9_421_0_CLK clkbuf_8_210_0_CLK/X clkbuf_9_421_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_50215_ _42373_/X _57491_/C _50214_/Y _50215_/X sky130_fd_sc_hd__o21a_4
X_85912_ _86587_/CLK _51984_/Y _73780_/B sky130_fd_sc_hd__dfxtp_4
X_81035_ _81061_/CLK _81035_/D _81035_/Q sky130_fd_sc_hd__dfxtp_4
X_58860_ _58858_/X _85450_/Q _58859_/X _58860_/Y sky130_fd_sc_hd__o21ai_4
X_51195_ _86056_/Q _51183_/X _51194_/Y _51195_/Y sky130_fd_sc_hd__o21ai_4
X_86892_ _86861_/CLK _45205_/Y _64434_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_315_0_CLK clkbuf_9_157_0_CLK/X _83476_/CLK sky130_fd_sc_hd__clkbuf_1
X_57811_ _57811_/A _57811_/X sky130_fd_sc_hd__buf_2
X_50146_ _48853_/A _50147_/C sky130_fd_sc_hd__buf_2
X_85843_ _85555_/CLK _52337_/Y _85843_/Q sky130_fd_sc_hd__dfxtp_4
X_58791_ _84800_/Q _58725_/X _58781_/X _58790_/X _84800_/D sky130_fd_sc_hd__a2bb2oi_4
X_67989_ _87384_/Q _67987_/X _67938_/X _67988_/X _67989_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_945_0_CLK clkbuf_9_472_0_CLK/X _87063_/CLK sky130_fd_sc_hd__clkbuf_1
X_57742_ _57738_/Y _57741_/Y _57718_/X _57742_/X sky130_fd_sc_hd__a21o_4
X_69728_ _69575_/A _69728_/X sky130_fd_sc_hd__buf_2
X_50077_ _48833_/A _50082_/B sky130_fd_sc_hd__buf_2
X_54954_ _85346_/Q _53449_/X _54953_/Y _54954_/Y sky130_fd_sc_hd__o21ai_4
X_85774_ _85778_/CLK _52682_/Y _85774_/Q sky130_fd_sc_hd__dfxtp_4
X_82986_ _82987_/CLK _74684_/Y _82986_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_436_0_CLK clkbuf_8_218_0_CLK/X clkbuf_9_436_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_87513_ _87520_/CLK _87513_/D _87513_/Q sky130_fd_sc_hd__dfxtp_4
X_53905_ _85545_/Q _53896_/X _53904_/Y _53905_/Y sky130_fd_sc_hd__o21ai_4
X_84725_ _83464_/CLK _84725_/D _59463_/A sky130_fd_sc_hd__dfxtp_4
X_81937_ _81989_/CLK _77876_/Y _77453_/A sky130_fd_sc_hd__dfxtp_4
X_57673_ _57673_/A _58230_/A sky130_fd_sc_hd__buf_2
X_69659_ _69086_/A _72947_/A _69659_/X sky130_fd_sc_hd__and2_4
X_54885_ _54885_/A _54885_/B _54885_/Y sky130_fd_sc_hd__nand2_4
X_59412_ _59394_/X _83484_/Q _59411_/Y _84740_/D sky130_fd_sc_hd__o21a_4
X_56624_ _56629_/B _72664_/C _72662_/C _56624_/Y sky130_fd_sc_hd__a21oi_4
X_87444_ _88201_/CLK _87444_/D _87444_/Q sky130_fd_sc_hd__dfxtp_4
X_41850_ _41839_/X _41841_/X _40515_/X _88123_/Q _41835_/X _41851_/A
+ sky130_fd_sc_hd__o32ai_4
X_53836_ _53819_/A _72012_/B _53836_/Y sky130_fd_sc_hd__nand2_4
X_72670_ _72668_/A _72668_/B _55646_/X _72670_/Y sky130_fd_sc_hd__nand3_4
X_84656_ _84672_/CLK _84656_/D _84656_/Q sky130_fd_sc_hd__dfxtp_4
X_81868_ _84441_/CLK _78059_/X _81868_/Q sky130_fd_sc_hd__dfxtp_4
X_40801_ _40628_/X _82874_/Q _40800_/X _40802_/A sky130_fd_sc_hd__o21ai_4
X_59343_ _59325_/X _59340_/Y _59341_/Y _59342_/X _59329_/X _59343_/X
+ sky130_fd_sc_hd__o32a_4
X_71621_ _71603_/Y _83435_/Q _71620_/Y _83435_/D sky130_fd_sc_hd__a21o_4
X_83607_ _85837_/CLK _83607_/D _83607_/Q sky130_fd_sc_hd__dfxtp_4
X_56555_ _55504_/Y _56580_/B _55552_/X _56556_/A sky130_fd_sc_hd__nand3_4
X_80819_ _80991_/CLK _83963_/Q _80819_/Q sky130_fd_sc_hd__dfxtp_4
X_87375_ _86834_/CLK _87375_/D _87375_/Q sky130_fd_sc_hd__dfxtp_4
X_53767_ _85572_/Q _53754_/X _53766_/Y _53767_/Y sky130_fd_sc_hd__o21ai_4
X_41781_ _40621_/X _41440_/A _41780_/X _41781_/Y sky130_fd_sc_hd__o21ai_4
X_84587_ _84333_/CLK _60611_/X _79127_/A sky130_fd_sc_hd__dfxtp_4
X_50979_ _50973_/X _50963_/B _50985_/C _46783_/X _50979_/X sky130_fd_sc_hd__and4_4
X_81799_ _81801_/CLK _81607_/Q _47473_/A sky130_fd_sc_hd__dfxtp_4
X_43520_ _43519_/Y _43520_/Y sky130_fd_sc_hd__inv_2
X_55506_ _55469_/X _55506_/X sky130_fd_sc_hd__buf_2
X_74340_ _72943_/A _74340_/X sky130_fd_sc_hd__buf_2
X_86326_ _86322_/CLK _49773_/Y _57891_/B sky130_fd_sc_hd__dfxtp_4
X_40732_ _40732_/A _40710_/B _40732_/X sky130_fd_sc_hd__or2_4
X_52718_ _52718_/A _52718_/B _52718_/Y sky130_fd_sc_hd__nand2_4
X_59274_ _59273_/X _85643_/Q _59196_/X _59274_/X sky130_fd_sc_hd__o21a_4
X_71552_ _71585_/A _71553_/B sky130_fd_sc_hd__buf_2
X_83538_ _86570_/CLK _83538_/D _83538_/Q sky130_fd_sc_hd__dfxtp_4
X_56486_ _56040_/X _56483_/X _56485_/Y _56486_/Y sky130_fd_sc_hd__o21ai_4
X_53698_ _53695_/Y _53696_/X _53697_/Y _53698_/Y sky130_fd_sc_hd__a21boi_4
XPHY_510 sky130_fd_sc_hd__decap_3
X_70503_ _70502_/Y _70504_/A sky130_fd_sc_hd__buf_2
X_58225_ _58225_/A _58225_/X sky130_fd_sc_hd__buf_2
X_43451_ _43450_/Y _87415_/D sky130_fd_sc_hd__inv_2
X_55437_ _55436_/Y _55438_/B sky130_fd_sc_hd__inv_2
X_74271_ _74038_/A _85890_/Q _74271_/X sky130_fd_sc_hd__and2_4
X_86257_ _85557_/CLK _86257_/D _65037_/B sky130_fd_sc_hd__dfxtp_4
XPHY_521 sky130_fd_sc_hd__decap_3
X_40663_ _40663_/A _40663_/Y sky130_fd_sc_hd__inv_2
X_52649_ _52648_/X _52654_/B _52643_/C _46744_/X _52649_/X sky130_fd_sc_hd__and4_4
X_71483_ _71827_/A _71483_/B _71439_/C _71716_/D _71483_/X sky130_fd_sc_hd__and4_4
X_83469_ _85959_/CLK _83469_/D _47787_/A sky130_fd_sc_hd__dfxtp_4
XPHY_532 sky130_fd_sc_hd__decap_3
XPHY_543 sky130_fd_sc_hd__decap_3
X_76010_ _76010_/A _76009_/Y _81742_/D sky130_fd_sc_hd__xor2_4
X_42402_ _42401_/X _42397_/X _40432_/X _87880_/Q _42398_/X _42403_/A
+ sky130_fd_sc_hd__o32ai_4
XPHY_554 sky130_fd_sc_hd__decap_3
X_73222_ _73219_/X _73220_/Y _73221_/X _73222_/Y sky130_fd_sc_hd__a21oi_4
X_85208_ _85269_/CLK _85208_/D _85208_/Q sky130_fd_sc_hd__dfxtp_4
X_70434_ _47932_/B _70422_/X _70433_/Y _83776_/D sky130_fd_sc_hd__o21ai_4
X_46170_ _46166_/A _45898_/X _46170_/C _46170_/Y sky130_fd_sc_hd__nand3_4
X_58156_ _63389_/A _58160_/B _58156_/Y sky130_fd_sc_hd__nand2_4
XPHY_565 sky130_fd_sc_hd__decap_3
X_43382_ _43367_/X _43375_/X _41424_/X _87450_/Q _43378_/X _43382_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55368_ _55360_/X _55368_/Y sky130_fd_sc_hd__inv_2
X_86188_ _83307_/CLK _86188_/D _86188_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_576 sky130_fd_sc_hd__decap_3
X_40594_ _48192_/A _49569_/A sky130_fd_sc_hd__buf_2
XPHY_587 sky130_fd_sc_hd__decap_3
XPHY_598 sky130_fd_sc_hd__decap_3
X_45121_ _56080_/C _45120_/X _45079_/X _45121_/X sky130_fd_sc_hd__o21a_4
X_57107_ _56960_/X _85083_/Q _57087_/X _57107_/Y sky130_fd_sc_hd__nor3_4
X_42333_ _41663_/X _42325_/X _87917_/Q _42326_/X _87917_/D sky130_fd_sc_hd__a2bb2o_4
X_54319_ _54315_/Y _54311_/X _54318_/X _85464_/D sky130_fd_sc_hd__a21oi_4
X_85139_ _85138_/CLK _85139_/D _85139_/Q sky130_fd_sc_hd__dfxtp_4
X_73153_ _73152_/X _73153_/X sky130_fd_sc_hd__buf_2
X_70365_ _71003_/A _71129_/A sky130_fd_sc_hd__buf_2
X_58087_ _58085_/X _85382_/Q _58086_/X _58087_/Y sky130_fd_sc_hd__o21ai_4
X_55299_ _55288_/Y _55292_/X _55298_/X _55299_/Y sky130_fd_sc_hd__a21boi_4
X_72104_ _72102_/Y _72083_/X _72103_/Y _72104_/Y sky130_fd_sc_hd__a21boi_4
X_45052_ _45350_/A _45052_/X sky130_fd_sc_hd__buf_2
X_57038_ _56732_/X _57038_/B _57038_/X sky130_fd_sc_hd__xor2_4
X_42264_ _41479_/X _42258_/X _87951_/Q _42259_/X _42264_/X sky130_fd_sc_hd__a2bb2o_4
X_77961_ _77960_/C _77961_/B _77944_/B _77961_/Y sky130_fd_sc_hd__nand3_4
X_73084_ _69722_/B _57377_/X _73055_/X _73083_/Y _73084_/X sky130_fd_sc_hd__a211o_4
X_70296_ _70246_/A _70296_/X sky130_fd_sc_hd__buf_2
Xclkbuf_5_15_0_CLK clkbuf_4_7_1_CLK/X clkbuf_6_31_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_44003_ _44003_/A _44003_/X sky130_fd_sc_hd__buf_2
X_79700_ _79700_/A _79700_/B _79710_/B sky130_fd_sc_hd__xor2_4
X_41215_ _41205_/X _41206_/X _41214_/X _88256_/Q _41194_/X _41216_/A
+ sky130_fd_sc_hd__o32ai_4
X_72035_ _72032_/Y _72033_/X _72034_/Y _72035_/Y sky130_fd_sc_hd__a21boi_4
X_76912_ _76899_/B _76899_/A _76888_/C _76888_/B _76911_/Y _76912_/X
+ sky130_fd_sc_hd__o41a_4
X_49860_ _58081_/B _49853_/X _49859_/Y _49860_/Y sky130_fd_sc_hd__o21ai_4
X_42195_ _41298_/X _42192_/X _87985_/Q _42193_/X _87985_/D sky130_fd_sc_hd__a2bb2o_4
X_77892_ _77892_/A _77902_/A sky130_fd_sc_hd__inv_2
X_48811_ _48831_/A _48811_/B _48811_/Y sky130_fd_sc_hd__nand2_4
X_79631_ _79627_/Y _79630_/X _79633_/A sky130_fd_sc_hd__xor2_4
X_41146_ _41143_/X _40615_/A _41145_/X _41147_/A sky130_fd_sc_hd__o21ai_4
X_76843_ _76837_/B _76837_/A _76842_/Y _76843_/Y sky130_fd_sc_hd__a21oi_4
X_49791_ _49769_/X _53005_/B _49791_/Y sky130_fd_sc_hd__nand2_4
X_58989_ _58982_/X _83436_/Q _58988_/Y _84780_/D sky130_fd_sc_hd__o21a_4
X_48742_ _65521_/B _48730_/X _48741_/Y _48742_/Y sky130_fd_sc_hd__o21ai_4
X_79562_ _79560_/Y _79561_/Y _79563_/B sky130_fd_sc_hd__nand2_4
X_45954_ _45883_/B _45954_/X sky130_fd_sc_hd__buf_2
X_41077_ _41040_/X _41041_/X _41076_/X _69486_/B _41037_/X _41078_/A
+ sky130_fd_sc_hd__o32ai_4
X_76774_ _76772_/Y _76773_/Y _76774_/X sky130_fd_sc_hd__xor2_4
X_73986_ _88353_/Q _56939_/X _72741_/X _73986_/Y sky130_fd_sc_hd__o21ai_4
X_78513_ _78499_/A _78482_/A _78513_/Y sky130_fd_sc_hd__nor2_4
X_44905_ _44975_/A _44905_/X sky130_fd_sc_hd__buf_2
X_75725_ _80915_/Q _75727_/A sky130_fd_sc_hd__inv_2
X_48673_ _48695_/A _48673_/B _48673_/Y sky130_fd_sc_hd__nand2_4
X_72937_ _72934_/X _72936_/X _72938_/B sky130_fd_sc_hd__nand2_4
X_60951_ _60905_/Y _60951_/Y sky130_fd_sc_hd__inv_2
X_79493_ _79493_/A _79493_/B _79494_/B sky130_fd_sc_hd__xor2_4
X_45885_ _73614_/A _45885_/X sky130_fd_sc_hd__buf_2
X_47624_ _47649_/A _53153_/B _47624_/Y sky130_fd_sc_hd__nand2_4
X_78444_ _82507_/Q _82763_/D _78444_/X sky130_fd_sc_hd__xor2_4
X_44836_ _44832_/X _44821_/X _41709_/X _67693_/B _44833_/X _44837_/A
+ sky130_fd_sc_hd__o32ai_4
X_63670_ _63670_/A _63670_/B _80347_/B _63670_/Y sky130_fd_sc_hd__nor3_4
X_75656_ _75656_/A _75658_/A sky130_fd_sc_hd__inv_2
X_60882_ _60997_/A _60882_/X sky130_fd_sc_hd__buf_2
X_72868_ _87067_/Q _73370_/B _72867_/X _72868_/Y sky130_fd_sc_hd__o21ai_4
X_62621_ _61683_/X _62515_/A _62534_/X _62621_/D _62621_/Y sky130_fd_sc_hd__nand4_4
X_74607_ _45257_/Y _74598_/X _74606_/X _83018_/D sky130_fd_sc_hd__o21ai_4
X_47555_ _47414_/A _47555_/X sky130_fd_sc_hd__buf_2
X_71819_ _71813_/A _71777_/B _71049_/A _71819_/X sky130_fd_sc_hd__and3_4
X_78375_ _78375_/A _78375_/B _78375_/C _78375_/Y sky130_fd_sc_hd__nand3_4
X_44767_ _41936_/A _44767_/X sky130_fd_sc_hd__buf_2
X_75587_ _80995_/Q _75587_/B _75587_/X sky130_fd_sc_hd__xor2_4
X_41979_ _41978_/Y _88084_/D sky130_fd_sc_hd__inv_2
X_72799_ _72798_/X _72799_/X sky130_fd_sc_hd__buf_2
X_46506_ _46493_/X _82923_/Q _46505_/Y _46507_/A sky130_fd_sc_hd__o21ai_4
X_65340_ _65984_/A _65340_/X sky130_fd_sc_hd__buf_2
X_77326_ _82217_/Q _77326_/Y sky130_fd_sc_hd__inv_2
X_43718_ _43606_/A _43718_/X sky130_fd_sc_hd__buf_2
X_62552_ _62851_/A _62672_/A sky130_fd_sc_hd__buf_2
X_74538_ _45909_/A _45933_/Y _74537_/Y _74538_/Y sky130_fd_sc_hd__o21ai_4
X_47486_ _47486_/A _53074_/D sky130_fd_sc_hd__buf_2
X_44698_ _44686_/X _44687_/X _40649_/Y _44697_/Y _44689_/X _44698_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49225_ _86430_/Q _49222_/X _49224_/Y _49225_/Y sky130_fd_sc_hd__o21ai_4
X_61503_ _61380_/A _61514_/D sky130_fd_sc_hd__buf_2
X_46437_ _46403_/X _49049_/A _46436_/X _46438_/A sky130_fd_sc_hd__o21ai_4
X_65271_ _65199_/X _86119_/Q _65224_/X _65270_/X _65271_/X sky130_fd_sc_hd__a211o_4
X_77257_ _77252_/Y _77255_/Y _77258_/A _77260_/A sky130_fd_sc_hd__a21oi_4
X_43649_ _40702_/A _43634_/X _68861_/B _43636_/X _43649_/X sky130_fd_sc_hd__a2bb2o_4
X_62483_ _62671_/A _62483_/X sky130_fd_sc_hd__buf_2
X_74469_ _74467_/Y _46300_/X _74468_/Y _83060_/D sky130_fd_sc_hd__a21boi_4
X_67010_ _67007_/X _67009_/X _66964_/X _67010_/X sky130_fd_sc_hd__a21o_4
X_64222_ _64234_/A _64234_/B _63376_/B _64221_/X _64222_/X sky130_fd_sc_hd__and4_4
X_76208_ _76207_/Y _76208_/Y sky130_fd_sc_hd__inv_2
X_61434_ _61434_/A _61434_/B _61434_/C _61434_/Y sky130_fd_sc_hd__nor3_4
X_49156_ _49205_/A _49156_/X sky130_fd_sc_hd__buf_2
X_46368_ _46367_/Y _50777_/B sky130_fd_sc_hd__buf_2
X_77188_ _77171_/A _77186_/Y _77187_/Y _77188_/X sky130_fd_sc_hd__a21o_4
X_48107_ _48142_/A _50365_/B _48107_/Y sky130_fd_sc_hd__nand2_4
X_45319_ _45319_/A _45272_/X _45319_/Y sky130_fd_sc_hd__nand2_4
X_64153_ _64187_/A _64187_/B _79950_/B _64153_/Y sky130_fd_sc_hd__nor3_4
X_76139_ _81727_/D _76139_/B _76139_/Y sky130_fd_sc_hd__nand2_4
X_49087_ _48976_/A _48586_/Y _49087_/Y sky130_fd_sc_hd__nand2_4
X_61365_ _84854_/Q _61365_/X sky130_fd_sc_hd__buf_2
X_46299_ _46653_/A _72083_/A sky130_fd_sc_hd__buf_2
X_63104_ _63101_/Y _63103_/X _63056_/X _63104_/Y sky130_fd_sc_hd__a21oi_4
X_48038_ _48033_/Y _48007_/X _48037_/X _86574_/D sky130_fd_sc_hd__a21oi_4
X_60316_ _60315_/X _60316_/Y sky130_fd_sc_hd__inv_2
X_64084_ _64077_/Y _64079_/Y _64083_/X _58457_/A _63736_/X _64084_/Y
+ sky130_fd_sc_hd__o32ai_4
X_68961_ _68957_/X _68960_/X _68748_/X _68961_/X sky130_fd_sc_hd__a21o_4
X_61296_ _61302_/A _72515_/D sky130_fd_sc_hd__buf_2
X_67912_ _67817_/X _67912_/B _67912_/X sky130_fd_sc_hd__and2_4
X_63035_ _79493_/A _63008_/X _63034_/Y _63035_/X sky130_fd_sc_hd__a21o_4
X_60247_ _60221_/A _60324_/B _60324_/C _60218_/A _60528_/A _60247_/Y
+ sky130_fd_sc_hd__a41oi_4
X_68892_ _68750_/A _68892_/B _68892_/X sky130_fd_sc_hd__and2_4
X_50000_ _49998_/Y _49977_/X _49999_/X _86284_/D sky130_fd_sc_hd__a21oi_4
X_67843_ _67817_/X _87710_/Q _67843_/X sky130_fd_sc_hd__and2_4
X_79829_ _79829_/A _79829_/B _79852_/B sky130_fd_sc_hd__and2_4
X_60178_ _60177_/X _60179_/A sky130_fd_sc_hd__buf_2
X_49989_ _72347_/B _49986_/X _49988_/Y _49989_/Y sky130_fd_sc_hd__o21ai_4
X_82840_ _82740_/CLK _82840_/D _82840_/Q sky130_fd_sc_hd__dfxtp_4
X_67774_ _87393_/Q _67751_/X _67702_/X _67773_/X _67774_/X sky130_fd_sc_hd__a211o_4
X_64986_ _64725_/A _65012_/A sky130_fd_sc_hd__buf_2
X_69513_ _69586_/A _69513_/B _69513_/X sky130_fd_sc_hd__and2_4
X_66725_ _87373_/Q _66678_/X _66629_/X _66724_/X _66725_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_7_113_0_CLK clkbuf_6_56_0_CLK/X clkbuf_8_227_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_51951_ _52486_/A _51951_/X sky130_fd_sc_hd__buf_2
X_63937_ _64353_/B _63920_/B _63951_/C _64015_/D _63937_/Y sky130_fd_sc_hd__nand4_4
X_82771_ _82774_/CLK _82771_/D _82771_/Q sky130_fd_sc_hd__dfxtp_4
X_84510_ _84503_/CLK _84510_/D _61192_/C sky130_fd_sc_hd__dfxtp_4
X_50902_ _50957_/A _50902_/X sky130_fd_sc_hd__buf_2
X_81722_ _84020_/CLK _81722_/D _41149_/A sky130_fd_sc_hd__dfxtp_4
X_69444_ _87517_/Q _69442_/X _69396_/X _69443_/X _69444_/X sky130_fd_sc_hd__a211o_4
X_54670_ _85399_/Q _54648_/X _54669_/Y _54670_/Y sky130_fd_sc_hd__o21ai_4
X_66656_ _66683_/A _66656_/B _66656_/X sky130_fd_sc_hd__and2_4
X_85490_ _83736_/CLK _54178_/Y _85490_/Q sky130_fd_sc_hd__dfxtp_4
X_51882_ _51870_/A _51870_/B _51870_/C _52709_/D _51882_/X sky130_fd_sc_hd__and4_4
X_63868_ _63751_/X _63900_/D sky130_fd_sc_hd__buf_2
Xclkbuf_10_83_0_CLK clkbuf_9_41_0_CLK/X _86757_/CLK sky130_fd_sc_hd__clkbuf_1
X_53621_ _53617_/Y _53619_/X _53620_/X _53621_/Y sky130_fd_sc_hd__a21oi_4
X_65607_ _65607_/A _65653_/B sky130_fd_sc_hd__buf_2
X_84441_ _84441_/CLK _61990_/Y _78064_/B sky130_fd_sc_hd__dfxtp_4
X_50833_ _86124_/Q _50820_/X _50832_/Y _50833_/Y sky130_fd_sc_hd__o21ai_4
X_62819_ _62819_/A _64379_/C _62819_/C _62782_/X _62819_/X sky130_fd_sc_hd__and4_4
X_81653_ _81682_/CLK _81685_/Q _76426_/A sky130_fd_sc_hd__dfxtp_4
X_69375_ _69651_/A _69612_/A sky130_fd_sc_hd__buf_2
X_66587_ _84105_/Q _59803_/X _66586_/X _84105_/D sky130_fd_sc_hd__a21bo_4
X_63799_ _63794_/X _63736_/X _63796_/Y _63797_/Y _63798_/X _63799_/X
+ sky130_fd_sc_hd__a41o_4
X_80604_ _84775_/Q _84167_/Q _80606_/A sky130_fd_sc_hd__xor2_4
X_56340_ _56109_/X _56337_/X _56339_/Y _85230_/D sky130_fd_sc_hd__o21ai_4
X_68326_ _68447_/A _68326_/X sky130_fd_sc_hd__buf_2
X_87160_ _86935_/CLK _87160_/D _87160_/Q sky130_fd_sc_hd__dfxtp_4
X_53552_ _53468_/A _53552_/B _53552_/Y sky130_fd_sc_hd__nand2_4
X_65538_ _65453_/X _85594_/Q _65470_/X _65537_/X _65538_/X sky130_fd_sc_hd__a211o_4
X_84372_ _84449_/CLK _84372_/D _84372_/Q sky130_fd_sc_hd__dfxtp_4
X_50764_ _50764_/A _53978_/B _50764_/Y sky130_fd_sc_hd__nand2_4
X_81584_ _83914_/CLK _65698_/C _81584_/Q sky130_fd_sc_hd__dfxtp_4
X_86111_ _83685_/CLK _50899_/Y _86111_/Q sky130_fd_sc_hd__dfxtp_4
X_52503_ _85809_/Q _52500_/X _52502_/Y _52503_/Y sky130_fd_sc_hd__o21ai_4
X_83323_ _83322_/CLK _83323_/D _56808_/A sky130_fd_sc_hd__dfxtp_4
X_56271_ _56168_/X _56188_/X _56270_/Y _56271_/Y sky130_fd_sc_hd__o21ai_4
X_80535_ _80529_/Y _80534_/Y _82264_/D sky130_fd_sc_hd__xor2_4
X_68257_ _83999_/Q _68238_/X _68256_/X _83999_/D sky130_fd_sc_hd__a21bo_4
X_87091_ _88263_/CLK _87091_/D _87091_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_98_0_CLK clkbuf_9_49_0_CLK/X _85067_/CLK sky130_fd_sc_hd__clkbuf_1
X_53483_ _85628_/Q _53476_/X _53482_/Y _53483_/Y sky130_fd_sc_hd__o21ai_4
X_65469_ _65350_/X _86206_/Q _65400_/X _65468_/X _65469_/X sky130_fd_sc_hd__a211o_4
X_50695_ _50695_/A _53910_/A _50695_/Y sky130_fd_sc_hd__nand2_4
X_58010_ _58696_/A _58010_/X sky130_fd_sc_hd__buf_2
X_67208_ _67205_/X _67207_/X _67113_/X _67208_/Y sky130_fd_sc_hd__a21oi_4
X_55222_ _85091_/Q _55152_/A _55133_/X _55221_/Y _55222_/X sky130_fd_sc_hd__a211o_4
X_86042_ _85818_/CLK _51275_/Y _64794_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_244_0_CLK clkbuf_8_245_0_CLK/A clkbuf_9_489_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_52434_ _52185_/X _53951_/B _52434_/Y sky130_fd_sc_hd__nand2_4
X_83254_ _85957_/CLK _72444_/Y _83254_/Q sky130_fd_sc_hd__dfxtp_4
X_80466_ _80478_/A _80478_/B _80471_/A sky130_fd_sc_hd__xor2_4
X_68188_ _68376_/A _68188_/X sky130_fd_sc_hd__buf_2
X_82205_ _82206_/CLK _77643_/X _82205_/Q sky130_fd_sc_hd__dfxtp_4
X_55153_ _80665_/Q _55168_/A sky130_fd_sc_hd__buf_2
X_67139_ _66899_/X _67130_/Y _67031_/X _67138_/Y _67139_/X sky130_fd_sc_hd__a211o_4
X_52365_ _52365_/A _52310_/B _52291_/C _52365_/X sky130_fd_sc_hd__and3_4
X_83185_ _81627_/CLK _83185_/D _70241_/C sky130_fd_sc_hd__dfxtp_4
X_80397_ _84755_/Q _80397_/B _80397_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_21_0_CLK clkbuf_9_10_0_CLK/X _85192_/CLK sky130_fd_sc_hd__clkbuf_1
X_54104_ _54123_/A _53428_/X _54111_/C _52938_/D _54104_/X sky130_fd_sc_hd__and4_4
X_51316_ _51310_/X _51316_/B _51316_/Y sky130_fd_sc_hd__nand2_4
X_70150_ _83524_/Q _83172_/Q _83519_/Q _83167_/Q _70150_/Y sky130_fd_sc_hd__a22oi_4
X_82136_ _81970_/CLK _82136_/D _77376_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_360_0_CLK clkbuf_8_180_0_CLK/X clkbuf_9_360_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_55084_ _55081_/Y _55076_/X _55083_/X _85322_/D sky130_fd_sc_hd__a21oi_4
X_59961_ _59961_/A _64386_/A sky130_fd_sc_hd__buf_2
X_52296_ _52294_/Y _52289_/X _52295_/X _52296_/Y sky130_fd_sc_hd__a21oi_4
X_87993_ _87993_/CLK _87993_/D _87993_/Q sky130_fd_sc_hd__dfxtp_4
X_58912_ _58877_/X _85926_/Q _58900_/X _58912_/X sky130_fd_sc_hd__o21a_4
X_54035_ _54320_/A _54035_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_254_0_CLK clkbuf_9_127_0_CLK/X _81094_/CLK sky130_fd_sc_hd__clkbuf_1
X_51247_ _51278_/A _46276_/A _51247_/X sky130_fd_sc_hd__and2_4
X_70081_ _70056_/A _70081_/X sky130_fd_sc_hd__buf_2
X_86944_ _88398_/CLK _86944_/D _86944_/Q sky130_fd_sc_hd__dfxtp_4
X_82067_ _82067_/CLK _82067_/D _82067_/Q sky130_fd_sc_hd__dfxtp_4
X_59892_ _60593_/B _61066_/B _59892_/Y sky130_fd_sc_hd__nor2_4
X_41000_ _40946_/A _41000_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_884_0_CLK clkbuf_9_442_0_CLK/X _86040_/CLK sky130_fd_sc_hd__clkbuf_1
X_81018_ _82152_/CLK _84226_/Q _81018_/Q sky130_fd_sc_hd__dfxtp_4
X_58843_ _84795_/Q _58843_/Y sky130_fd_sc_hd__inv_2
X_51178_ _51174_/Y _51175_/X _51177_/X _86060_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_36_0_CLK clkbuf_9_18_0_CLK/X _85144_/CLK sky130_fd_sc_hd__clkbuf_1
X_86875_ _86873_/CLK _86875_/D _63051_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_375_0_CLK clkbuf_9_375_0_CLK/A clkbuf_9_375_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_50129_ _65012_/B _50113_/X _50128_/Y _50129_/Y sky130_fd_sc_hd__o21ai_4
X_73840_ _73837_/X _73838_/Y _73839_/X _73840_/X sky130_fd_sc_hd__a21o_4
X_85826_ _85826_/CLK _85826_/D _85826_/Q sky130_fd_sc_hd__dfxtp_4
X_58774_ _58771_/Y _58773_/Y _58761_/X _58774_/X sky130_fd_sc_hd__a21o_4
X_55986_ _74284_/C _55985_/Y _55986_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_10_269_0_CLK clkbuf_9_134_0_CLK/X _83766_/CLK sky130_fd_sc_hd__clkbuf_1
X_57725_ _46224_/X _85408_/Q _57724_/X _57725_/Y sky130_fd_sc_hd__o21ai_4
X_42951_ _42951_/A _42951_/X sky130_fd_sc_hd__buf_2
X_54937_ _54932_/A _54942_/B _54932_/C _53244_/D _54937_/X sky130_fd_sc_hd__and4_4
X_73771_ _68588_/Y _73674_/X _73698_/X _73770_/Y _73771_/X sky130_fd_sc_hd__a211o_4
X_85757_ _85757_/CLK _52776_/Y _85757_/Q sky130_fd_sc_hd__dfxtp_4
X_70983_ _70983_/A _70983_/X sky130_fd_sc_hd__buf_2
X_82969_ _82206_/CLK _82777_/Q _46696_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_899_0_CLK clkbuf_9_449_0_CLK/X _86982_/CLK sky130_fd_sc_hd__clkbuf_1
X_75510_ _75510_/A _75482_/Y _75509_/Y _75510_/X sky130_fd_sc_hd__and3_4
X_41902_ _41902_/A _40591_/B _46616_/A _41902_/X sky130_fd_sc_hd__and3_4
X_72722_ _72721_/X _72722_/X sky130_fd_sc_hd__buf_2
X_84708_ _84355_/CLK _59719_/Y _80568_/A sky130_fd_sc_hd__dfxtp_4
X_57656_ _84960_/Q _57656_/X sky130_fd_sc_hd__buf_2
X_45670_ _45668_/X _61542_/A _45608_/X _45670_/Y sky130_fd_sc_hd__o21ai_4
X_76490_ _76489_/Y _76491_/C sky130_fd_sc_hd__inv_2
X_54868_ _85363_/Q _54865_/X _54867_/Y _54868_/Y sky130_fd_sc_hd__o21ai_4
X_42882_ _42874_/X _42875_/X _41616_/X _87670_/Q _42881_/X _42883_/A
+ sky130_fd_sc_hd__o32ai_4
X_85688_ _85688_/CLK _53152_/Y _85688_/Q sky130_fd_sc_hd__dfxtp_4
X_56607_ _56607_/A _56607_/X sky130_fd_sc_hd__buf_2
X_44621_ _40985_/Y _44618_/X _87029_/Q _44619_/X _87029_/D sky130_fd_sc_hd__a2bb2o_4
X_75441_ _75423_/Y _75427_/B _75426_/A _75441_/X sky130_fd_sc_hd__o21a_4
X_87427_ _87686_/CLK _43428_/Y _87427_/Q sky130_fd_sc_hd__dfxtp_4
X_41833_ _41824_/X _41825_/X _40474_/X _66978_/B _41821_/X _41834_/A
+ sky130_fd_sc_hd__o32ai_4
X_53819_ _53819_/A _53819_/B _53819_/Y sky130_fd_sc_hd__nand2_4
X_72653_ _70193_/A _72645_/X _72652_/Y _83202_/D sky130_fd_sc_hd__a21bo_4
X_84639_ _83216_/CLK _60301_/X _79775_/A sky130_fd_sc_hd__dfxtp_4
X_57587_ _71964_/A _71960_/C sky130_fd_sc_hd__buf_2
X_54799_ _54797_/Y _54774_/X _54798_/X _54799_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_822_0_CLK clkbuf_9_411_0_CLK/X _82931_/CLK sky130_fd_sc_hd__clkbuf_1
X_47340_ _54685_/D _52993_/D sky130_fd_sc_hd__buf_2
X_59326_ _59255_/A _59326_/X sky130_fd_sc_hd__buf_2
X_71604_ _71603_/Y _71604_/X sky130_fd_sc_hd__buf_2
X_78160_ _82669_/Q _78160_/B _78160_/X sky130_fd_sc_hd__xor2_4
X_44552_ _44547_/X _44548_/X _40839_/X _87057_/Q _44549_/X _44552_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56538_ _56538_/A _56535_/X _55732_/B _56538_/Y sky130_fd_sc_hd__nand3_4
X_75372_ _80694_/Q _80950_/D _75372_/Y sky130_fd_sc_hd__nor2_4
X_41764_ _41764_/A _41764_/Y sky130_fd_sc_hd__inv_2
X_87358_ _86784_/CLK _87358_/D _87358_/Q sky130_fd_sc_hd__dfxtp_4
X_72584_ _72584_/A _72530_/A _72584_/C _72585_/A sky130_fd_sc_hd__nand3_4
X_77111_ _77111_/A _82290_/D _77111_/X sky130_fd_sc_hd__xor2_4
X_43503_ _43425_/X _43503_/X sky130_fd_sc_hd__buf_2
X_74323_ _74325_/A _74325_/B _55854_/X _74323_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_9_313_0_CLK clkbuf_9_313_0_CLK/A clkbuf_9_313_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_86309_ _86627_/CLK _49867_/Y _58096_/B sky130_fd_sc_hd__dfxtp_4
X_40715_ _40621_/X _40888_/A _40714_/X _40716_/A sky130_fd_sc_hd__o21ai_4
X_59257_ _86668_/Q _59282_/B _59257_/Y sky130_fd_sc_hd__nor2_4
X_47271_ _47128_/A _47271_/X sky130_fd_sc_hd__buf_2
X_71535_ _71137_/B _71536_/A sky130_fd_sc_hd__buf_2
X_78091_ _82563_/Q _78091_/B _78091_/Y sky130_fd_sc_hd__nor2_4
X_44483_ _44624_/A _44549_/A sky130_fd_sc_hd__buf_2
X_56469_ _56545_/A _56454_/B _56469_/C _56469_/Y sky130_fd_sc_hd__nand3_4
X_87289_ _87824_/CLK _43738_/X _87289_/Q sky130_fd_sc_hd__dfxtp_4
X_41695_ _82901_/Q _41660_/X _41695_/X sky130_fd_sc_hd__or2_4
X_49010_ _48946_/X _48495_/Y _49009_/Y _52328_/B sky130_fd_sc_hd__a21o_4
X_46222_ _46222_/A _46222_/B _46221_/Y _46222_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_207_0_CLK clkbuf_9_103_0_CLK/X _80728_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_340 sky130_fd_sc_hd__decap_3
X_58208_ _58191_/X _58204_/Y _58207_/Y _84908_/D sky130_fd_sc_hd__a21oi_4
X_77042_ _77047_/A _77041_/Y _77042_/X sky130_fd_sc_hd__and2_4
X_43434_ _43329_/X _43434_/X sky130_fd_sc_hd__buf_2
X_74254_ _74016_/X _85603_/Q _56933_/X _74253_/X _74254_/X sky130_fd_sc_hd__a211o_4
XPHY_351 sky130_fd_sc_hd__decap_3
X_40646_ _40645_/Y _40646_/X sky130_fd_sc_hd__buf_2
X_59188_ _59154_/A _86354_/Q _59188_/Y sky130_fd_sc_hd__nor2_4
X_71466_ _70880_/B _71435_/B _70763_/A _71476_/D _71466_/X sky130_fd_sc_hd__and4_4
XPHY_362 sky130_fd_sc_hd__decap_3
Xclkbuf_10_837_0_CLK clkbuf_9_418_0_CLK/X _85955_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_373 sky130_fd_sc_hd__decap_3
XPHY_384 sky130_fd_sc_hd__decap_3
X_73205_ _73351_/A _73205_/X sky130_fd_sc_hd__buf_2
X_46153_ _46120_/A _46120_/B _46170_/C _46158_/A sky130_fd_sc_hd__a21o_4
X_58139_ _58085_/X _85378_/Q _58138_/X _58139_/Y sky130_fd_sc_hd__o21ai_4
X_70417_ _70416_/Y _71162_/B sky130_fd_sc_hd__buf_2
XPHY_395 sky130_fd_sc_hd__decap_3
X_43365_ _43347_/X _43350_/X _41382_/X _87457_/Q _43353_/X _43366_/A
+ sky130_fd_sc_hd__o32ai_4
X_74185_ _41969_/Y _73930_/X _73031_/X _74184_/Y _74185_/X sky130_fd_sc_hd__a211o_4
X_40577_ _49048_/A _40577_/X sky130_fd_sc_hd__buf_2
X_71397_ _71396_/Y _71397_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_328_0_CLK clkbuf_9_329_0_CLK/A clkbuf_9_328_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_45104_ _85204_/Q _45102_/X _45103_/X _45104_/Y sky130_fd_sc_hd__o21ai_4
X_42316_ _42316_/A _87925_/D sky130_fd_sc_hd__inv_2
X_61150_ _64523_/D _61176_/B sky130_fd_sc_hd__buf_2
X_73136_ _72959_/X _85587_/Q _73092_/X _73135_/X _73136_/X sky130_fd_sc_hd__a211o_4
X_70348_ _70348_/A _70348_/B _83083_/Q _70348_/D _70348_/X sky130_fd_sc_hd__and4_4
X_46084_ _46111_/B _46141_/A _46115_/A _46114_/A _46162_/A sky130_fd_sc_hd__nor4_4
X_43296_ _43296_/A _43296_/X sky130_fd_sc_hd__buf_2
X_78993_ _78993_/A _78993_/B _78994_/B sky130_fd_sc_hd__xor2_4
X_60101_ _60091_/B _60100_/Y _59951_/C _60102_/A sky130_fd_sc_hd__o21ai_4
X_49912_ _49928_/A _53127_/B _49912_/Y sky130_fd_sc_hd__nand2_4
X_45035_ _64305_/B _61427_/B sky130_fd_sc_hd__buf_2
X_42247_ _41429_/X _42222_/X _87961_/Q _42224_/X _87961_/D sky130_fd_sc_hd__a2bb2o_4
X_61081_ _61081_/A _61122_/A sky130_fd_sc_hd__buf_2
X_73067_ _73067_/A _73067_/X sky130_fd_sc_hd__buf_2
X_77944_ _77961_/B _77944_/B _77950_/A sky130_fd_sc_hd__xor2_4
X_70279_ _83812_/Q _74762_/A sky130_fd_sc_hd__inv_2
X_60032_ _60064_/A _59873_/B _60032_/C _60032_/Y sky130_fd_sc_hd__nor3_4
X_72018_ _72017_/X _53841_/B _72018_/Y sky130_fd_sc_hd__nand2_4
X_49843_ _49569_/A _49924_/A sky130_fd_sc_hd__buf_2
X_42178_ _42178_/A _42178_/Y sky130_fd_sc_hd__inv_2
X_77875_ _77875_/A _77874_/X _77879_/A sky130_fd_sc_hd__nand2_4
X_79614_ _65268_/C _83256_/Q _79614_/X sky130_fd_sc_hd__xor2_4
X_41129_ _41100_/X _40588_/A _41128_/X _41129_/Y sky130_fd_sc_hd__o21ai_4
X_64840_ _64508_/A _64870_/B sky130_fd_sc_hd__buf_2
X_76826_ _81589_/Q _76826_/B _76826_/X sky130_fd_sc_hd__xor2_4
X_49774_ _49769_/X _52991_/B _49774_/Y sky130_fd_sc_hd__nand2_4
X_46986_ _59090_/A _46955_/X _46985_/Y _46986_/Y sky130_fd_sc_hd__o21ai_4
X_48725_ _48725_/A _48391_/X _48725_/Y sky130_fd_sc_hd__nand2_4
X_79545_ _79543_/Y _79545_/B _79545_/Y sky130_fd_sc_hd__nand2_4
X_45937_ _44164_/X _44140_/X _44004_/Y _45918_/Y _45937_/Y sky130_fd_sc_hd__nand4_4
X_64771_ _64768_/X _64770_/X _64619_/X _64775_/A sky130_fd_sc_hd__a21o_4
X_76757_ _76744_/A _76757_/B _76758_/B sky130_fd_sc_hd__and2_4
X_61983_ _61522_/X _61933_/X _61967_/C _61952_/D _61983_/Y sky130_fd_sc_hd__nand4_4
X_73969_ _86990_/Q _73776_/X _73968_/X _73981_/C sky130_fd_sc_hd__o21ai_4
X_66510_ _66508_/Y _59756_/X _66509_/X _84109_/D sky130_fd_sc_hd__a21o_4
X_63722_ _61003_/A _64192_/B sky130_fd_sc_hd__buf_2
X_75708_ _75708_/A _75707_/Y _75711_/A sky130_fd_sc_hd__xor2_4
X_60934_ _60934_/A _60934_/X sky130_fd_sc_hd__buf_2
X_48656_ _48656_/A _48849_/A sky130_fd_sc_hd__buf_2
X_67490_ _67517_/A _88237_/Q _67490_/X sky130_fd_sc_hd__and2_4
X_79476_ _79476_/A _79476_/B _79476_/X sky130_fd_sc_hd__xor2_4
X_45868_ _55211_/B _45736_/B _45868_/Y sky130_fd_sc_hd__nor2_4
X_76688_ _76688_/A _76687_/Y _81446_/D sky130_fd_sc_hd__xor2_4
X_47607_ _47595_/A _47645_/B _47595_/C _53144_/D _47607_/X sky130_fd_sc_hd__and4_4
X_66441_ _65004_/X _66476_/B _65007_/X _66441_/Y sky130_fd_sc_hd__nand3_4
X_78427_ _78426_/B _78413_/A _78412_/A _78427_/X sky130_fd_sc_hd__o21a_4
X_44819_ _41662_/Y _44817_/X _86937_/Q _44818_/X _86937_/D sky130_fd_sc_hd__a2bb2o_4
X_63653_ _63670_/A _63670_/B _80371_/B _63653_/Y sky130_fd_sc_hd__nor3_4
X_75639_ _75632_/A _75639_/B _75641_/A sky130_fd_sc_hd__nor2_4
X_48587_ _48586_/Y _48565_/B _48587_/Y sky130_fd_sc_hd__nand2_4
X_60865_ _60997_/A _60865_/B _60865_/C _60864_/X _60866_/A sky130_fd_sc_hd__nand4_4
X_45799_ _55281_/A _45798_/X _45743_/X _45799_/X sky130_fd_sc_hd__o21a_4
X_62604_ _62671_/A _62653_/A sky130_fd_sc_hd__buf_2
X_69160_ _83944_/Q _69066_/X _69159_/X _83944_/D sky130_fd_sc_hd__a21bo_4
X_47538_ _72129_/A _47524_/X _47537_/Y _47538_/Y sky130_fd_sc_hd__o21ai_4
X_66372_ _66366_/X _64649_/Y _66371_/Y _66372_/Y sky130_fd_sc_hd__o21ai_4
X_78358_ _78358_/A _78358_/B _78376_/B sky130_fd_sc_hd__nand2_4
X_63584_ _63398_/A _63657_/A sky130_fd_sc_hd__buf_2
X_60796_ _60727_/A _60794_/Y _60795_/X _60796_/Y sky130_fd_sc_hd__nand3_4
X_68111_ _66702_/X _66705_/X _68106_/X _68111_/Y sky130_fd_sc_hd__a21oi_4
X_65323_ _84206_/Q _65296_/X _65322_/Y _84206_/D sky130_fd_sc_hd__a21o_4
X_77309_ _77310_/A _77307_/Y _77308_/Y _77315_/A sky130_fd_sc_hd__o21ai_4
X_62535_ _61593_/B _62504_/X _62534_/X _62475_/X _62536_/D sky130_fd_sc_hd__nand4_4
X_69091_ _69087_/X _69090_/X _68697_/X _69091_/X sky130_fd_sc_hd__a21o_4
X_47469_ _47469_/A _53067_/B sky130_fd_sc_hd__buf_2
X_78289_ _82590_/Q _78290_/B _78289_/X sky130_fd_sc_hd__or2_4
X_49208_ _64580_/B _49204_/X _49207_/Y _49208_/Y sky130_fd_sc_hd__o21ai_4
X_80320_ _80320_/A _80320_/B _80320_/Y sky130_fd_sc_hd__nand2_4
X_68042_ _68437_/A _87701_/Q _68042_/X sky130_fd_sc_hd__and2_4
X_65254_ _65252_/X _83288_/Q _65230_/X _65253_/X _65254_/X sky130_fd_sc_hd__a211o_4
X_50480_ _50478_/Y _50455_/X _50479_/X _86193_/D sky130_fd_sc_hd__a21oi_4
X_62466_ _62457_/X _62461_/Y _62465_/X _84848_/Q _62440_/X _62466_/Y
+ sky130_fd_sc_hd__o32ai_4
X_64205_ _64267_/A _64457_/C sky130_fd_sc_hd__buf_2
X_49139_ _49048_/A _49139_/B _50693_/A sky130_fd_sc_hd__nor2_4
X_61417_ _61375_/A _61417_/B _61398_/C _61417_/Y sky130_fd_sc_hd__nand3_4
X_80251_ _80251_/A _80250_/X _80259_/A sky130_fd_sc_hd__nand2_4
X_65185_ _65009_/X _86155_/Q _65182_/X _65184_/X _65185_/X sky130_fd_sc_hd__a211o_4
X_62397_ _62342_/A _62341_/X _62397_/C _62397_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_7_90_0_CLK clkbuf_7_91_0_CLK/A clkbuf_7_90_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_52150_ _50447_/A _52140_/X _52156_/C _52150_/X sky130_fd_sc_hd__and3_4
X_64136_ _84871_/Q _64136_/B _64136_/X sky130_fd_sc_hd__or2_4
X_61348_ _61348_/A _61394_/A sky130_fd_sc_hd__buf_2
X_80182_ _80198_/A _80189_/A _80182_/X sky130_fd_sc_hd__xor2_4
X_69993_ _68471_/X _68476_/X _69992_/X _69993_/X sky130_fd_sc_hd__a21o_4
X_51101_ _51101_/A _51101_/X sky130_fd_sc_hd__buf_2
X_52081_ _52121_/A _50378_/B _52081_/Y sky130_fd_sc_hd__nand2_4
X_68944_ _69011_/A _68944_/B _68944_/X sky130_fd_sc_hd__and2_4
X_64067_ _64067_/A _64161_/B sky130_fd_sc_hd__buf_2
X_61279_ _61312_/A _72502_/A sky130_fd_sc_hd__inv_2
X_84990_ _86558_/CLK _57508_/Y _84990_/Q sky130_fd_sc_hd__dfxtp_4
X_51032_ _86086_/Q _51020_/X _51031_/Y _51032_/Y sky130_fd_sc_hd__o21ai_4
X_63018_ _60472_/A _60443_/A _63001_/A _60404_/Y _63018_/X sky130_fd_sc_hd__a211o_4
X_83941_ _83940_/CLK _83941_/D _81405_/D sky130_fd_sc_hd__dfxtp_4
X_68875_ _68993_/A _68875_/X sky130_fd_sc_hd__buf_2
X_55840_ _55837_/X _55839_/X _55516_/X _55845_/B sky130_fd_sc_hd__a21o_4
X_67826_ _67873_/A _67826_/B _67826_/X sky130_fd_sc_hd__and2_4
X_86660_ _84746_/CLK _47203_/Y _59361_/A sky130_fd_sc_hd__dfxtp_4
X_83872_ _83133_/CLK _83872_/D _82552_/D sky130_fd_sc_hd__dfxtp_4
X_85611_ _85601_/CLK _85611_/D _85611_/Q sky130_fd_sc_hd__dfxtp_4
X_82823_ _82248_/CLK _82823_/D _82823_/Q sky130_fd_sc_hd__dfxtp_4
X_55771_ _55768_/X _55771_/B _55772_/A sky130_fd_sc_hd__and2_4
X_67757_ _86958_/Q _67706_/X _67755_/X _67756_/X _67757_/X sky130_fd_sc_hd__a211o_4
X_86591_ _86592_/CLK _47862_/Y _65935_/B sky130_fd_sc_hd__dfxtp_4
X_52983_ _52980_/Y _52975_/X _52982_/X _52983_/Y sky130_fd_sc_hd__a21oi_4
X_64969_ _65196_/A _64913_/B _84220_/Q _64969_/X sky130_fd_sc_hd__and3_4
X_57510_ _84989_/Q _57493_/X _57509_/Y _57510_/Y sky130_fd_sc_hd__o21ai_4
X_88330_ _84970_/CLK _40811_/X _88330_/Q sky130_fd_sc_hd__dfxtp_4
X_54722_ _54719_/Y _54720_/X _54721_/X _54722_/Y sky130_fd_sc_hd__a21oi_4
X_66708_ _66526_/X _66696_/Y _66672_/X _66707_/Y _66708_/X sky130_fd_sc_hd__a211o_4
X_85542_ _85542_/CLK _53920_/Y _85542_/Q sky130_fd_sc_hd__dfxtp_4
X_51934_ _51934_/A _51934_/X sky130_fd_sc_hd__buf_2
X_82754_ _82965_/CLK _82754_/D _82946_/D sky130_fd_sc_hd__dfxtp_4
X_58490_ _58490_/A _58498_/B _58490_/Y sky130_fd_sc_hd__nand2_4
X_67688_ _67806_/A _67688_/X sky130_fd_sc_hd__buf_2
X_81705_ _81703_/CLK _75976_/A _41068_/B sky130_fd_sc_hd__dfxtp_4
X_57441_ _58425_/A _57441_/X sky130_fd_sc_hd__buf_2
X_69427_ _69305_/A _69427_/B _69427_/X sky130_fd_sc_hd__and2_4
X_88261_ _87103_/CLK _88261_/D _68723_/B sky130_fd_sc_hd__dfxtp_4
X_54653_ _54651_/Y _54638_/X _54652_/X _54653_/Y sky130_fd_sc_hd__a21oi_4
X_66639_ _69315_/A _66639_/X sky130_fd_sc_hd__buf_2
X_85473_ _85471_/CLK _54271_/Y _85473_/Q sky130_fd_sc_hd__dfxtp_4
X_51865_ _51870_/A _51851_/B _51870_/C _52694_/D _51865_/X sky130_fd_sc_hd__and4_4
X_82685_ _82933_/CLK _82685_/D _78278_/A sky130_fd_sc_hd__dfxtp_4
X_87212_ _87446_/CLK _87212_/D _87212_/Q sky130_fd_sc_hd__dfxtp_4
X_53604_ _53604_/A _50381_/B _53604_/Y sky130_fd_sc_hd__nand2_4
X_84424_ _84424_/CLK _84424_/D _84424_/Q sky130_fd_sc_hd__dfxtp_4
X_50816_ _50787_/X _50816_/B _50816_/Y sky130_fd_sc_hd__nand2_4
X_57372_ _57440_/A _57372_/X sky130_fd_sc_hd__buf_2
X_81636_ _81684_/CLK _81668_/Q _76176_/A sky130_fd_sc_hd__dfxtp_4
X_69358_ _69383_/A _69358_/B _69358_/X sky130_fd_sc_hd__and2_4
X_88192_ _87116_/CLK _88192_/D _67041_/B sky130_fd_sc_hd__dfxtp_4
X_54584_ _54558_/A _54584_/X sky130_fd_sc_hd__buf_2
X_51796_ _51796_/A _46701_/X _51796_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_7_43_0_CLK clkbuf_7_42_0_CLK/A clkbuf_8_87_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_59111_ _58721_/A _59189_/B sky130_fd_sc_hd__buf_2
X_68309_ _67893_/X _67896_/X _68283_/X _68309_/Y sky130_fd_sc_hd__a21oi_4
X_56323_ _56332_/A _56312_/X _55865_/B _56323_/Y sky130_fd_sc_hd__nand3_4
X_87143_ _88220_/CLK _87143_/D _87143_/Q sky130_fd_sc_hd__dfxtp_4
X_53535_ _53468_/A _53535_/B _53535_/Y sky130_fd_sc_hd__nand2_4
X_84355_ _84355_/CLK _84355_/D _79447_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_183_0_CLK clkbuf_7_91_0_CLK/X clkbuf_9_367_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_50747_ _50745_/Y _50735_/X _50746_/Y _86142_/D sky130_fd_sc_hd__a21boi_4
X_81567_ _83926_/CLK _81567_/D _81567_/Q sky130_fd_sc_hd__dfxtp_4
X_69289_ _87528_/Q _69261_/X _69248_/X _69288_/X _69289_/X sky130_fd_sc_hd__a211o_4
X_40500_ _40456_/X _41572_/A _40499_/X _40500_/X sky130_fd_sc_hd__o21a_4
X_71320_ _71320_/A _71320_/X sky130_fd_sc_hd__buf_2
X_59042_ _58094_/A _59043_/A sky130_fd_sc_hd__buf_2
X_83306_ _83306_/CLK _71995_/Y _83306_/Q sky130_fd_sc_hd__dfxtp_4
X_56254_ _56134_/X _56242_/X _56253_/Y _56254_/Y sky130_fd_sc_hd__o21ai_4
X_80518_ _80518_/A _80518_/B _80531_/B sky130_fd_sc_hd__xnor2_4
X_41480_ _41479_/X _41455_/X _88207_/Q _41457_/X _41480_/X sky130_fd_sc_hd__a2bb2o_4
X_87074_ _87077_/CLK _87074_/D _87074_/Q sky130_fd_sc_hd__dfxtp_4
X_53466_ _53687_/A _53466_/X sky130_fd_sc_hd__buf_2
X_84286_ _84668_/CLK _84286_/D _80133_/B sky130_fd_sc_hd__dfxtp_4
X_50678_ _50675_/Y _50676_/X _50677_/X _86155_/D sky130_fd_sc_hd__a21oi_4
X_81498_ _81749_/CLK _81498_/D _81498_/Q sky130_fd_sc_hd__dfxtp_4
X_55205_ _85029_/Q _55157_/X _55168_/X _55204_/Y _55205_/X sky130_fd_sc_hd__a211o_4
X_86025_ _86122_/CLK _86025_/D _86025_/Q sky130_fd_sc_hd__dfxtp_4
X_52417_ _52414_/Y _52415_/X _52416_/X _85827_/D sky130_fd_sc_hd__a21oi_4
X_40431_ _40429_/X _82326_/Q _40430_/X _40431_/X sky130_fd_sc_hd__o21a_4
X_71251_ _51947_/B _71239_/X _71250_/Y _83558_/D sky130_fd_sc_hd__o21ai_4
X_83237_ _84350_/CLK _83237_/D _79467_/B sky130_fd_sc_hd__dfxtp_4
X_80449_ _80436_/X _80447_/X _80448_/X _80449_/Y sky130_fd_sc_hd__a21oi_4
X_56185_ _55684_/X _56460_/D sky130_fd_sc_hd__buf_2
Xclkbuf_7_58_0_CLK clkbuf_7_58_0_CLK/A clkbuf_7_58_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_53397_ _53397_/A _53388_/B _53388_/C _51192_/D _53397_/X sky130_fd_sc_hd__and4_4
X_70202_ _70231_/A _70214_/A sky130_fd_sc_hd__buf_2
X_43150_ _43146_/X _43149_/X _40839_/X _73126_/A _43121_/X _43151_/A
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_8_198_0_CLK clkbuf_7_99_0_CLK/X clkbuf_8_198_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_55136_ _57027_/A _55126_/X _55134_/X _55135_/X _55136_/X sky130_fd_sc_hd__a211o_4
X_40362_ _42081_/A _40362_/X sky130_fd_sc_hd__buf_2
X_52348_ _52271_/A _52349_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_193_0_CLK clkbuf_9_96_0_CLK/X _84280_/CLK sky130_fd_sc_hd__clkbuf_1
X_71182_ _52163_/B _71164_/Y _71181_/Y _71182_/Y sky130_fd_sc_hd__o21ai_4
X_83168_ _83167_/CLK _73023_/X _83168_/Q sky130_fd_sc_hd__dfxtp_4
X_42101_ _42101_/A _42101_/Y sky130_fd_sc_hd__inv_2
X_70133_ _70133_/A _70134_/C sky130_fd_sc_hd__inv_2
X_82119_ _82145_/CLK _82119_/D _82107_/D sky130_fd_sc_hd__dfxtp_4
X_43081_ _43072_/X _43075_/X _40702_/X _74033_/A _43080_/X _43081_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55067_ _55054_/A _54903_/B _55067_/Y sky130_fd_sc_hd__nand2_4
X_59944_ _59943_/X _62532_/A sky130_fd_sc_hd__buf_2
X_52279_ _52274_/A _52319_/A sky130_fd_sc_hd__buf_2
X_75990_ _75980_/Y _75990_/B _75990_/Y sky130_fd_sc_hd__nand2_4
X_87976_ _88158_/CLK _42217_/Y _87976_/Q sky130_fd_sc_hd__dfxtp_4
X_83099_ _83095_/CLK _83099_/D _70306_/C sky130_fd_sc_hd__dfxtp_4
X_54018_ _53921_/A _54018_/X sky130_fd_sc_hd__buf_2
X_42032_ _42031_/Y _88064_/D sky130_fd_sc_hd__inv_2
X_74941_ _81136_/D _74960_/C _74958_/A sky130_fd_sc_hd__xor2_4
X_70064_ _69864_/X _69866_/X _69994_/X _70064_/X sky130_fd_sc_hd__a21o_4
X_86927_ _87652_/CLK _44840_/X _67719_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_121_0_CLK clkbuf_7_60_0_CLK/X clkbuf_9_243_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_59875_ _59875_/A _59875_/X sky130_fd_sc_hd__buf_2
X_46840_ _46840_/A _52706_/B sky130_fd_sc_hd__inv_2
X_58826_ _84797_/Q _58725_/X _58820_/X _58825_/X _84797_/D sky130_fd_sc_hd__a2bb2oi_4
X_77660_ _77660_/A _77658_/Y _77656_/Y _77693_/C sky130_fd_sc_hd__nand3_4
X_74872_ _74870_/Y _74866_/Y _74871_/Y _74872_/Y sky130_fd_sc_hd__o21ai_4
X_86858_ _84534_/CLK _45732_/Y _62057_/D sky130_fd_sc_hd__dfxtp_4
X_76611_ _76611_/A _81375_/Q _76609_/Y _76611_/Y sky130_fd_sc_hd__nand3_4
X_73823_ _43057_/Y _72900_/X _73772_/X _73822_/Y _73823_/X sky130_fd_sc_hd__a211o_4
X_85809_ _86422_/CLK _85809_/D _85809_/Q sky130_fd_sc_hd__dfxtp_4
X_58757_ _58756_/X _85938_/Q _58664_/X _58757_/X sky130_fd_sc_hd__o21a_4
X_46771_ _46806_/A _50971_/B _46771_/Y sky130_fd_sc_hd__nand2_4
X_77591_ _77591_/A _77596_/A sky130_fd_sc_hd__buf_2
X_43983_ _43983_/A _44186_/A sky130_fd_sc_hd__inv_2
X_55969_ _55691_/A _85183_/Q _55969_/X sky130_fd_sc_hd__and2_4
X_86789_ _86814_/CLK _86789_/D _66985_/B sky130_fd_sc_hd__dfxtp_4
X_48510_ _74431_/A _52166_/A sky130_fd_sc_hd__buf_2
X_79330_ _79330_/A _79330_/B _79331_/B sky130_fd_sc_hd__xor2_4
X_45722_ _45719_/Y _45627_/X _45720_/X _45721_/Y _45722_/X sky130_fd_sc_hd__a211o_4
X_57708_ _57837_/A _57708_/X sky130_fd_sc_hd__buf_2
X_76542_ _76584_/C _76548_/A sky130_fd_sc_hd__inv_2
Xclkbuf_8_136_0_CLK clkbuf_7_68_0_CLK/X clkbuf_8_136_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_42934_ _42835_/X _42934_/X sky130_fd_sc_hd__buf_2
X_49490_ _49486_/Y _49487_/X _49489_/X _49490_/Y sky130_fd_sc_hd__a21oi_4
X_73754_ _73751_/X _73753_/X _73679_/X _73767_/B sky130_fd_sc_hd__a21o_4
Xclkbuf_10_131_0_CLK clkbuf_9_65_0_CLK/X _81808_/CLK sky130_fd_sc_hd__clkbuf_1
X_70966_ _70966_/A _70969_/C sky130_fd_sc_hd__buf_2
X_58688_ _58688_/A _58688_/B _58688_/Y sky130_fd_sc_hd__nor2_4
X_48441_ _46485_/X _48489_/B sky130_fd_sc_hd__buf_2
X_72705_ _72688_/A _72714_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_761_0_CLK clkbuf_9_380_0_CLK/X _88036_/CLK sky130_fd_sc_hd__clkbuf_1
X_79261_ _79257_/Y _79270_/B _79263_/A sky130_fd_sc_hd__xor2_4
X_45653_ _82993_/Q _45654_/A sky130_fd_sc_hd__inv_2
X_57639_ _71993_/A _71970_/A sky130_fd_sc_hd__buf_2
X_76473_ _76473_/A _76473_/Y sky130_fd_sc_hd__inv_2
X_42865_ _42865_/A _42865_/Y sky130_fd_sc_hd__inv_2
X_73685_ _73605_/X _86236_/Q _73683_/X _73684_/X _73685_/X sky130_fd_sc_hd__a211o_4
X_70897_ _70869_/A _70903_/B _70899_/C _70899_/D _70897_/Y sky130_fd_sc_hd__nand4_4
X_78212_ _78213_/A _78213_/B _78220_/B sky130_fd_sc_hd__or2_4
X_44604_ _40935_/A _44602_/X _87039_/Q _44603_/X _44604_/X sky130_fd_sc_hd__a2bb2o_4
X_75424_ _75424_/A _75424_/B _75427_/B sky130_fd_sc_hd__nor2_4
X_41816_ _40418_/X _41813_/X _66802_/B _41814_/X _88138_/D sky130_fd_sc_hd__a2bb2o_4
X_60650_ _60712_/B _60694_/B sky130_fd_sc_hd__buf_2
Xclkbuf_9_252_0_CLK clkbuf_9_253_0_CLK/A clkbuf_9_252_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_48372_ _48471_/A _48372_/X sky130_fd_sc_hd__buf_2
X_72636_ _70165_/A _72631_/X _72635_/Y _72636_/X sky130_fd_sc_hd__a21bo_4
X_79192_ _79190_/Y _79192_/B _79193_/B sky130_fd_sc_hd__nand2_4
X_45584_ _45584_/A _45584_/Y sky130_fd_sc_hd__inv_2
X_42796_ _42723_/A _42796_/X sky130_fd_sc_hd__buf_2
X_47323_ _47323_/A _47324_/A sky130_fd_sc_hd__inv_2
X_59309_ _59273_/X _85640_/Q _59308_/X _59309_/X sky130_fd_sc_hd__o21a_4
X_78143_ _78143_/A _78143_/B _78144_/B sky130_fd_sc_hd__xnor2_4
Xclkbuf_10_146_0_CLK clkbuf_9_73_0_CLK/X _83187_/CLK sky130_fd_sc_hd__clkbuf_1
X_44535_ _87064_/Q _44535_/Y sky130_fd_sc_hd__inv_2
X_75355_ _75347_/X _75354_/X _75355_/X sky130_fd_sc_hd__xor2_4
X_41747_ _41747_/A _41718_/X _41747_/X sky130_fd_sc_hd__or2_4
X_60581_ _60612_/A _60612_/B _79135_/A _60581_/Y sky130_fd_sc_hd__nor3_4
X_72567_ _72573_/A _72573_/B _79414_/B _72567_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_10_776_0_CLK clkbuf_9_388_0_CLK/X _82145_/CLK sky130_fd_sc_hd__clkbuf_1
X_62320_ _62471_/A _62334_/D sky130_fd_sc_hd__buf_2
X_74306_ _74302_/X _74310_/B _74306_/C _74306_/Y sky130_fd_sc_hd__nand3_4
X_47254_ _86654_/Q _47240_/X _47253_/Y _47254_/Y sky130_fd_sc_hd__o21ai_4
X_71518_ _53240_/B _71508_/X _71517_/Y _83470_/D sky130_fd_sc_hd__o21ai_4
X_78074_ _78074_/A _78074_/B _78074_/X sky130_fd_sc_hd__xor2_4
X_44466_ _44603_/A _44466_/X sky130_fd_sc_hd__buf_2
X_75286_ _75267_/Y _75268_/Y _75269_/Y _75294_/A sky130_fd_sc_hd__o21a_4
X_41678_ _41678_/A _41678_/Y sky130_fd_sc_hd__inv_2
X_72498_ _63630_/A _72498_/B _72498_/Y sky130_fd_sc_hd__nand2_4
X_46205_ _46120_/A _72527_/B _46204_/Y _46205_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_267_0_CLK clkbuf_9_267_0_CLK/A clkbuf_9_267_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_170 sky130_fd_sc_hd__decap_3
X_77025_ _77018_/A _82277_/D _77025_/Y sky130_fd_sc_hd__nand2_4
X_43417_ _43399_/X _43404_/X _41520_/X _87431_/Q _43407_/X _43418_/A
+ sky130_fd_sc_hd__o32ai_4
X_74237_ _74237_/A _66326_/B _74237_/X sky130_fd_sc_hd__and2_4
X_62251_ _62212_/A _62251_/B _62251_/C _62251_/D _62251_/Y sky130_fd_sc_hd__nand4_4
XPHY_181 sky130_fd_sc_hd__decap_3
X_40629_ _40629_/A _48631_/A sky130_fd_sc_hd__buf_2
X_47185_ _47150_/A _47184_/X _47185_/Y sky130_fd_sc_hd__nand2_4
X_71449_ _71445_/X _58151_/B _71448_/Y _83496_/D sky130_fd_sc_hd__a21o_4
X_44397_ _44381_/X _44382_/X _41493_/X _87129_/Q _44383_/X _44398_/A
+ sky130_fd_sc_hd__o32ai_4
XPHY_192 sky130_fd_sc_hd__decap_3
X_61202_ _61202_/A _61202_/B _61202_/Y sky130_fd_sc_hd__nor2_4
X_46136_ _44184_/X _57665_/A sky130_fd_sc_hd__buf_2
X_43348_ _43347_/X _43319_/X _41332_/X _87466_/Q _43330_/X _43349_/A
+ sky130_fd_sc_hd__o32ai_4
X_62182_ _62177_/Y _62166_/X _62181_/Y _84427_/D sky130_fd_sc_hd__a21oi_4
X_74168_ _74165_/X _74167_/X _73602_/X _74168_/X sky130_fd_sc_hd__a21o_4
X_61133_ _61110_/Y _61118_/X _61254_/B _61131_/Y _61132_/Y _84519_/D
+ sky130_fd_sc_hd__a41oi_4
X_73119_ _73116_/X _73118_/X _73120_/B sky130_fd_sc_hd__nand2_4
X_46067_ _40556_/A _46067_/X sky130_fd_sc_hd__buf_2
X_43279_ _41134_/X _43277_/X _87503_/Q _43278_/X _87503_/D sky130_fd_sc_hd__a2bb2o_4
X_66990_ _87118_/Q _66988_/X _66919_/X _66989_/X _66990_/X sky130_fd_sc_hd__a211o_4
X_78976_ _82645_/Q _78976_/Y sky130_fd_sc_hd__inv_2
X_74099_ _74096_/X _74098_/X _73489_/X _74102_/A sky130_fd_sc_hd__a21o_4
X_45018_ _56041_/C _44963_/X _45004_/X _45018_/X sky130_fd_sc_hd__o21a_4
X_65941_ _65938_/X _65868_/B _65940_/X _65941_/Y sky130_fd_sc_hd__nand3_4
X_61064_ _61055_/A _59771_/X _84522_/Q _61064_/X sky130_fd_sc_hd__or3_4
X_77927_ _77925_/Y _77927_/B _77928_/A sky130_fd_sc_hd__xor2_4
Xclkbuf_10_714_0_CLK clkbuf_9_357_0_CLK/X _86824_/CLK sky130_fd_sc_hd__clkbuf_1
X_60015_ _60011_/X _59995_/X _62548_/D _60014_/X _46199_/X _60015_/Y
+ sky130_fd_sc_hd__a32oi_4
X_49826_ _49416_/A _49854_/A sky130_fd_sc_hd__buf_2
X_68660_ _69654_/A _68660_/X sky130_fd_sc_hd__buf_2
X_65872_ _65888_/A _65888_/B _65872_/C _65872_/Y sky130_fd_sc_hd__nor3_4
X_77858_ _77844_/Y _77845_/Y _77832_/A _81934_/D _77858_/X sky130_fd_sc_hd__a2bb2o_4
X_67611_ _67522_/X _67602_/Y _67507_/X _67610_/Y _67611_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_9_205_0_CLK clkbuf_8_102_0_CLK/X clkbuf_9_205_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_64823_ _64810_/A _86425_/Q _64823_/X sky130_fd_sc_hd__and2_4
X_76809_ _76809_/A _76809_/B _76809_/X sky130_fd_sc_hd__xor2_4
X_49757_ _49757_/A _52973_/B _49757_/Y sky130_fd_sc_hd__nand2_4
X_68591_ _44148_/A _69661_/A sky130_fd_sc_hd__buf_2
X_46969_ _46959_/A _52777_/B _46969_/Y sky130_fd_sc_hd__nand2_4
X_77789_ _77788_/X _77789_/Y sky130_fd_sc_hd__inv_2
X_48708_ _81762_/Q _48959_/B _48708_/X sky130_fd_sc_hd__or2_4
X_67542_ _67538_/X _67541_/X _67423_/X _67542_/Y sky130_fd_sc_hd__a21oi_4
X_79528_ _60374_/C _79528_/Y sky130_fd_sc_hd__inv_2
X_64754_ _64752_/X _86172_/Q _64716_/X _64753_/X _64754_/X sky130_fd_sc_hd__a211o_4
X_49688_ _49416_/A _49688_/X sky130_fd_sc_hd__buf_2
X_61966_ _61966_/A _61967_/C sky130_fd_sc_hd__buf_2
Xclkbuf_10_729_0_CLK clkbuf_9_364_0_CLK/X _87026_/CLK sky130_fd_sc_hd__clkbuf_1
X_63705_ _63696_/A _62174_/X _63705_/X sky130_fd_sc_hd__and2_4
X_48639_ _48639_/A _48843_/B sky130_fd_sc_hd__buf_2
X_60917_ _64189_/C _64172_/C sky130_fd_sc_hd__buf_2
X_67473_ _67354_/X _67473_/X sky130_fd_sc_hd__buf_2
X_79459_ _79459_/A _79459_/B _79482_/B sky130_fd_sc_hd__and2_4
X_64685_ _64657_/X _83310_/Q _64600_/X _64684_/X _64685_/X sky130_fd_sc_hd__a211o_4
X_61897_ _61722_/A _61960_/A sky130_fd_sc_hd__buf_2
X_69212_ _68737_/A _69212_/X sky130_fd_sc_hd__buf_2
X_66424_ _66422_/Y _66423_/Y _65842_/X _66424_/Y sky130_fd_sc_hd__a21oi_4
X_51650_ _85971_/Q _51647_/X _51649_/Y _51650_/Y sky130_fd_sc_hd__o21ai_4
X_63636_ _63615_/A _63615_/B _63636_/C _63636_/Y sky130_fd_sc_hd__nor3_4
X_82470_ _82675_/CLK _82470_/D _78290_/B sky130_fd_sc_hd__dfxtp_4
X_60848_ _60848_/A _60857_/D sky130_fd_sc_hd__buf_2
X_50601_ _50580_/A _71994_/B _50601_/Y sky130_fd_sc_hd__nand2_4
X_81421_ _82648_/CLK _81453_/Q _81421_/Q sky130_fd_sc_hd__dfxtp_4
X_69143_ _69139_/X _69141_/X _69142_/X _69143_/Y sky130_fd_sc_hd__a21oi_4
X_66355_ _66352_/X _66354_/X _66355_/Y sky130_fd_sc_hd__nand2_4
X_51581_ _51578_/Y _51557_/X _51580_/X _51581_/Y sky130_fd_sc_hd__a21oi_4
X_63567_ _63554_/A _63554_/B _80455_/B _63567_/Y sky130_fd_sc_hd__nor3_4
X_60779_ _61075_/C _60629_/Y _60616_/Y _60644_/C _60667_/A _63371_/A
+ sky130_fd_sc_hd__a41oi_4
Xclkbuf_4_5_0_CLK clkbuf_4_5_0_CLK/A clkbuf_4_5_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_53320_ _51842_/A _53347_/A sky130_fd_sc_hd__buf_2
X_65306_ _64961_/A _65307_/A sky130_fd_sc_hd__buf_2
X_84140_ _84220_/CLK _84140_/D _84140_/Q sky130_fd_sc_hd__dfxtp_4
X_50532_ _50529_/Y _50525_/X _50531_/X _86183_/D sky130_fd_sc_hd__a21oi_4
X_62518_ _62517_/Y _64454_/A sky130_fd_sc_hd__buf_2
X_81352_ _81352_/CLK _76696_/X _81352_/Q sky130_fd_sc_hd__dfxtp_4
X_69074_ _44745_/A _68864_/X _68891_/X _69073_/X _69074_/X sky130_fd_sc_hd__a211o_4
X_66286_ _64722_/X _85607_/Q _64724_/X _66285_/X _66286_/X sky130_fd_sc_hd__a211o_4
X_63498_ _63372_/A _63498_/X sky130_fd_sc_hd__buf_2
X_80303_ _80301_/Y _80303_/B _80304_/B sky130_fd_sc_hd__nand2_4
X_68025_ _68025_/A _88150_/Q _68025_/X sky130_fd_sc_hd__and2_4
X_53251_ _53259_/A _51728_/B _53251_/Y sky130_fd_sc_hd__nand2_4
X_65237_ _65211_/X _85513_/Q _65212_/X _65236_/X _65237_/X sky130_fd_sc_hd__a211o_4
X_84071_ _81461_/CLK _67404_/X _84071_/Q sky130_fd_sc_hd__dfxtp_4
X_50463_ _50459_/Y _50455_/X _50462_/X _50463_/Y sky130_fd_sc_hd__a21oi_4
X_62449_ _62534_/A _62449_/X sky130_fd_sc_hd__buf_2
X_81283_ _81794_/CLK _76971_/X _81283_/Q sky130_fd_sc_hd__dfxtp_4
X_52202_ _85869_/Q _52178_/X _52201_/Y _52202_/Y sky130_fd_sc_hd__o21ai_4
X_83022_ _83022_/CLK _83022_/D _45196_/A sky130_fd_sc_hd__dfxtp_4
X_80234_ _80230_/Y _80233_/Y _80244_/B sky130_fd_sc_hd__xor2_4
X_53182_ _53180_/Y _53163_/X _53181_/X _85682_/D sky130_fd_sc_hd__a21oi_4
X_65168_ _64739_/A _65397_/A sky130_fd_sc_hd__buf_2
X_50394_ _86209_/Q _50333_/X _50393_/Y _50394_/Y sky130_fd_sc_hd__o21ai_4
X_52133_ _72957_/B _52125_/X _52132_/Y _52133_/Y sky130_fd_sc_hd__o21ai_4
X_64119_ _64012_/A _64178_/C sky130_fd_sc_hd__buf_2
X_87830_ _87834_/CLK _87830_/D _74224_/A sky130_fd_sc_hd__dfxtp_4
X_80165_ _84945_/Q _65559_/C _80167_/A sky130_fd_sc_hd__xor2_4
X_57990_ _58749_/A _57991_/A sky130_fd_sc_hd__buf_2
X_65099_ _64797_/A _65099_/X sky130_fd_sc_hd__buf_2
X_69976_ _69943_/X _69974_/Y _69938_/X _69975_/Y _69976_/X sky130_fd_sc_hd__a211o_4
X_52064_ _52070_/A _50365_/B _52064_/Y sky130_fd_sc_hd__nand2_4
X_56941_ _56940_/Y _57084_/A sky130_fd_sc_hd__buf_2
X_68927_ _68907_/X _68882_/X _68915_/Y _68926_/Y _68927_/X sky130_fd_sc_hd__a211o_4
X_87761_ _87758_/CLK _87761_/D _68425_/B sky130_fd_sc_hd__dfxtp_4
X_84973_ _86541_/CLK _57594_/Y _84973_/Q sky130_fd_sc_hd__dfxtp_4
X_80096_ _80080_/Y _80083_/Y _80095_/X _80096_/X sky130_fd_sc_hd__a21o_4
X_51015_ _51009_/Y _51011_/X _51014_/X _86090_/D sky130_fd_sc_hd__a21oi_4
X_86712_ _86393_/CLK _46709_/Y _58677_/A sky130_fd_sc_hd__dfxtp_4
X_59660_ _60414_/B _60353_/B _59660_/C _59660_/D _59805_/A sky130_fd_sc_hd__and4_4
X_83924_ _81322_/CLK _83924_/D _81388_/D sky130_fd_sc_hd__dfxtp_4
X_56872_ _56688_/X _56867_/X _56871_/Y _56872_/Y sky130_fd_sc_hd__o21ai_4
X_68858_ _87839_/Q _68859_/B sky130_fd_sc_hd__inv_2
X_87692_ _87126_/CLK _87692_/D _66745_/B sky130_fd_sc_hd__dfxtp_4
X_58611_ _58607_/Y _58609_/Y _58610_/X _58611_/X sky130_fd_sc_hd__a21o_4
X_55823_ _55817_/A _55823_/B _55823_/X sky130_fd_sc_hd__and2_4
X_67809_ _87967_/Q _67713_/X _67761_/X _67808_/X _67809_/X sky130_fd_sc_hd__a211o_4
X_86643_ _86005_/CLK _86643_/D _86643_/Q sky130_fd_sc_hd__dfxtp_4
X_83855_ _82536_/CLK _83855_/D _82535_/D sky130_fd_sc_hd__dfxtp_4
X_59591_ _59591_/A _59689_/A sky130_fd_sc_hd__buf_2
X_68789_ _83961_/Q _68713_/X _68788_/X _83961_/D sky130_fd_sc_hd__a21bo_4
X_70820_ _71219_/A _70952_/B _70703_/X _70820_/Y sky130_fd_sc_hd__nand3_4
X_58542_ _58538_/X _83360_/Q _58541_/Y _84824_/D sky130_fd_sc_hd__o21a_4
X_82806_ _82529_/CLK _82838_/Q _82806_/Q sky130_fd_sc_hd__dfxtp_4
X_55754_ _45290_/A _55190_/X _44095_/A _55753_/X _55754_/X sky130_fd_sc_hd__a211o_4
X_86574_ _86530_/CLK _86574_/D _66183_/B sky130_fd_sc_hd__dfxtp_4
X_40980_ _82296_/Q _40932_/X _40980_/X sky130_fd_sc_hd__or2_4
X_52966_ _85722_/Q _52957_/X _52965_/Y _52966_/Y sky130_fd_sc_hd__o21ai_4
X_83786_ _83787_/CLK _70351_/X _74727_/A sky130_fd_sc_hd__dfxtp_4
X_80998_ _82532_/CLK _84206_/Q _80998_/Q sky130_fd_sc_hd__dfxtp_4
X_88313_ _88324_/CLK _88313_/D _88313_/Q sky130_fd_sc_hd__dfxtp_4
X_54705_ _54718_/A _47372_/Y _54705_/Y sky130_fd_sc_hd__nand2_4
X_85525_ _85815_/CLK _85525_/D _85525_/Q sky130_fd_sc_hd__dfxtp_4
X_51917_ _85922_/Q _51900_/X _51916_/Y _51917_/Y sky130_fd_sc_hd__o21ai_4
X_70751_ _70753_/A _70722_/A _70751_/Y sky130_fd_sc_hd__nand2_4
X_58473_ _64412_/C _58474_/A sky130_fd_sc_hd__buf_2
X_82737_ _81019_/CLK _84121_/Q _82737_/Q sky130_fd_sc_hd__dfxtp_4
X_55685_ _55684_/X _56171_/C sky130_fd_sc_hd__buf_2
X_52897_ _52885_/A _47174_/X _52897_/Y sky130_fd_sc_hd__nand2_4
X_57424_ _57423_/Y _85007_/D sky130_fd_sc_hd__inv_2
X_88244_ _82629_/CLK _88244_/D _69129_/B sky130_fd_sc_hd__dfxtp_4
X_42650_ _42649_/Y _42650_/Y sky130_fd_sc_hd__inv_2
X_54636_ _54636_/A _47260_/A _54636_/Y sky130_fd_sc_hd__nand2_4
X_85456_ _85459_/CLK _85456_/D _85456_/Q sky130_fd_sc_hd__dfxtp_4
X_73470_ _73353_/A _85861_/Q _73470_/X sky130_fd_sc_hd__and2_4
X_51848_ _51853_/A _50981_/B _51848_/Y sky130_fd_sc_hd__nand2_4
X_70682_ _70682_/A _70676_/B _70676_/C _70682_/Y sky130_fd_sc_hd__nor3_4
X_82668_ _82803_/CLK _82668_/D _82668_/Q sky130_fd_sc_hd__dfxtp_4
X_41601_ _41600_/Y _41601_/X sky130_fd_sc_hd__buf_2
X_72421_ _72419_/X _85352_/Q _72420_/X _72421_/Y sky130_fd_sc_hd__o21ai_4
X_84407_ _84407_/CLK _84407_/D _62485_/C sky130_fd_sc_hd__dfxtp_4
X_57355_ _57236_/X _45811_/A _57355_/Y sky130_fd_sc_hd__nand2_4
X_81619_ _81259_/CLK _76407_/B _81619_/Q sky130_fd_sc_hd__dfxtp_4
X_88175_ _88175_/CLK _88175_/D _67434_/B sky130_fd_sc_hd__dfxtp_4
X_42581_ _42573_/X _42574_/X _40839_/X _87813_/Q _42580_/X _42581_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54567_ _54540_/A _54567_/X sky130_fd_sc_hd__buf_2
X_85387_ _85484_/CLK _85387_/D _85387_/Q sky130_fd_sc_hd__dfxtp_4
X_51779_ _51779_/A _51779_/B _51779_/Y sky130_fd_sc_hd__nand2_4
X_82599_ _82879_/CLK _78851_/B _82567_/D sky130_fd_sc_hd__dfxtp_4
X_44320_ _44320_/A _44318_/A _44320_/Y sky130_fd_sc_hd__nor2_4
X_56306_ _56296_/A _56298_/X _56306_/C _56306_/Y sky130_fd_sc_hd__nand3_4
X_75140_ _75138_/A _75138_/B _75140_/Y sky130_fd_sc_hd__nand2_4
X_87126_ _87126_/CLK _44402_/X _87126_/Q sky130_fd_sc_hd__dfxtp_4
X_53518_ _53509_/A _73864_/A _53518_/Y sky130_fd_sc_hd__nand2_4
X_41532_ _41529_/X _41530_/X _88197_/Q _41531_/X _88197_/D sky130_fd_sc_hd__a2bb2o_4
X_72352_ _59286_/A _72352_/X sky130_fd_sc_hd__buf_2
X_84338_ _83218_/CLK _84338_/D _79267_/A sky130_fd_sc_hd__dfxtp_4
X_57286_ _57280_/X _57282_/Y _57283_/Y _57285_/Y _57286_/X sky130_fd_sc_hd__a211o_4
X_54498_ _54483_/A _54503_/B _54483_/C _54498_/D _54498_/X sky130_fd_sc_hd__and4_4
X_71303_ _71303_/A _71303_/B _71302_/X _71303_/Y sky130_fd_sc_hd__nand3_4
X_59025_ _59022_/Y _59024_/Y _58966_/X _59025_/X sky130_fd_sc_hd__a21o_4
X_44251_ _59036_/A _58020_/A sky130_fd_sc_hd__buf_2
X_56237_ _56233_/A _56243_/B _85264_/Q _56237_/Y sky130_fd_sc_hd__nand3_4
X_75071_ _75070_/Y _75071_/Y sky130_fd_sc_hd__inv_2
X_41463_ _81184_/Q _41459_/B _41463_/X sky130_fd_sc_hd__or2_4
X_87057_ _88062_/CLK _44553_/Y _87057_/Q sky130_fd_sc_hd__dfxtp_4
X_53449_ _53448_/X _53449_/X sky130_fd_sc_hd__buf_2
X_72283_ _72209_/X _85972_/Q _72282_/X _72283_/Y sky130_fd_sc_hd__o21ai_4
X_84269_ _84269_/CLK _64165_/Y _79937_/B sky130_fd_sc_hd__dfxtp_4
X_43202_ _43047_/X _53944_/A _40925_/X _43201_/Y _43021_/X _87541_/D
+ sky130_fd_sc_hd__o32ai_4
X_74022_ _72874_/A _74022_/X sky130_fd_sc_hd__buf_2
X_86008_ _86008_/CLK _86008_/D _86008_/Q sky130_fd_sc_hd__dfxtp_4
X_40414_ _40413_/X _40414_/X sky130_fd_sc_hd__buf_2
X_71234_ _71221_/A _71235_/A sky130_fd_sc_hd__buf_2
X_44182_ _44181_/X _72461_/A sky130_fd_sc_hd__buf_2
X_56168_ _56168_/A _56168_/X sky130_fd_sc_hd__buf_2
X_41394_ _41393_/X _41362_/X _67813_/B _41363_/X _88223_/D sky130_fd_sc_hd__a2bb2o_4
X_55119_ _85314_/Q _55098_/X _55118_/Y _55119_/Y sky130_fd_sc_hd__o21ai_4
X_43133_ _43133_/A _43133_/Y sky130_fd_sc_hd__inv_2
X_78830_ _78830_/A _78829_/Y _78831_/B sky130_fd_sc_hd__xor2_4
X_40345_ _46610_/A _46725_/A sky130_fd_sc_hd__buf_2
X_71165_ _71164_/Y _71165_/X sky130_fd_sc_hd__buf_2
X_48990_ _48984_/Y _48985_/X _48989_/X _48990_/Y sky130_fd_sc_hd__a21oi_4
X_56099_ _56099_/A _56099_/X sky130_fd_sc_hd__buf_2
X_70116_ _83128_/Q _70117_/D sky130_fd_sc_hd__inv_2
X_47941_ _47912_/A _48231_/B _47941_/Y sky130_fd_sc_hd__nand2_4
X_43064_ _43038_/X _43050_/X _40661_/X _73873_/A _43061_/X _43065_/A
+ sky130_fd_sc_hd__o32ai_4
X_59927_ _59927_/A _59927_/Y sky130_fd_sc_hd__inv_2
X_78761_ _78747_/A _78746_/Y _78737_/Y _78761_/X sky130_fd_sc_hd__o21a_4
X_71096_ _70905_/D _71099_/C sky130_fd_sc_hd__buf_2
X_75973_ _75949_/A _75954_/A _75961_/A _75970_/A _75974_/B sky130_fd_sc_hd__and4_4
X_87959_ _87952_/CLK _87959_/D _87959_/Q sky130_fd_sc_hd__dfxtp_4
X_42015_ _42014_/Y _88071_/D sky130_fd_sc_hd__inv_2
X_77712_ _77712_/A _82124_/Q _77712_/Y sky130_fd_sc_hd__nand2_4
X_74924_ _81132_/D _74912_/B _74924_/Y sky130_fd_sc_hd__nand2_4
X_70047_ _82544_/D _70029_/X _70046_/X _70047_/X sky130_fd_sc_hd__a21bo_4
X_47872_ _47872_/A _52139_/A sky130_fd_sc_hd__buf_2
X_59858_ _59858_/A _59858_/Y sky130_fd_sc_hd__inv_2
X_78692_ _78691_/Y _78693_/C sky130_fd_sc_hd__inv_2
X_49611_ _49609_/Y _49596_/X _49610_/X _49611_/Y sky130_fd_sc_hd__a21oi_4
X_46823_ _46818_/Y _46798_/X _46822_/X _86700_/D sky130_fd_sc_hd__a21oi_4
X_58809_ _57848_/A _58810_/A sky130_fd_sc_hd__buf_2
X_77643_ _77643_/A _77643_/B _77643_/X sky130_fd_sc_hd__xor2_4
X_74855_ _81124_/D _74854_/B _74855_/Y sky130_fd_sc_hd__nand2_4
X_59789_ _59789_/A _59591_/A _59789_/Y sky130_fd_sc_hd__nor2_4
X_49542_ _49406_/A _49571_/A sky130_fd_sc_hd__buf_2
X_61820_ _61820_/A _61865_/B sky130_fd_sc_hd__buf_2
X_73806_ _73731_/X _86231_/Q _73804_/X _73805_/X _73806_/X sky130_fd_sc_hd__a211o_4
X_46754_ _46753_/Y _52654_/D sky130_fd_sc_hd__buf_2
X_77574_ _77575_/A _77571_/Y _77575_/B _77576_/A sky130_fd_sc_hd__a21o_4
X_43966_ _43963_/X _43965_/X _80669_/Q _43969_/A sky130_fd_sc_hd__a21o_4
X_74786_ _74786_/A _74720_/C _74804_/D _74780_/D _74786_/Y sky130_fd_sc_hd__nand4_4
X_71998_ _71993_/X _71998_/B _71998_/Y sky130_fd_sc_hd__nand2_4
X_79313_ _79291_/A _79303_/X _79313_/Y sky130_fd_sc_hd__nand2_4
X_45705_ _45705_/A _45705_/X sky130_fd_sc_hd__buf_2
X_76525_ _76521_/Y _76524_/C _76520_/Y _76525_/Y sky130_fd_sc_hd__o21ai_4
X_42917_ _42945_/A _42917_/X sky130_fd_sc_hd__buf_2
X_49473_ _86381_/Q _49470_/X _49472_/Y _49473_/Y sky130_fd_sc_hd__o21ai_4
X_73737_ _73735_/X _85626_/Q _73661_/X _73736_/X _73737_/X sky130_fd_sc_hd__a211o_4
X_61751_ _61726_/X _61734_/X _61750_/Y _58149_/A _61719_/X _61751_/Y
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_9_191_0_CLK clkbuf_8_95_0_CLK/X clkbuf_9_191_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_46685_ _46685_/A _46685_/X sky130_fd_sc_hd__buf_2
X_70949_ _70947_/A _70949_/B _70947_/C _70949_/Y sky130_fd_sc_hd__nand3_4
X_43897_ _43896_/X _43897_/X sky130_fd_sc_hd__buf_2
X_48424_ _48469_/A _52128_/B _48424_/Y sky130_fd_sc_hd__nand2_4
X_60702_ _60652_/A _60677_/A _60702_/C _60702_/Y sky130_fd_sc_hd__nand3_4
X_79244_ _84792_/Q _66495_/C _79244_/X sky130_fd_sc_hd__xor2_4
X_45636_ _85138_/Q _45556_/X _45378_/X _45636_/X sky130_fd_sc_hd__o21a_4
X_64470_ _64465_/Y _64466_/X _64467_/X _64469_/Y _64440_/X _64470_/X
+ sky130_fd_sc_hd__o41a_4
X_76456_ _76456_/A _76453_/A _76456_/Y sky130_fd_sc_hd__nand2_4
X_42848_ _42429_/A _42945_/A sky130_fd_sc_hd__buf_2
X_61682_ _61305_/A _61682_/B _61682_/C _61682_/Y sky130_fd_sc_hd__nand3_4
X_73668_ _73668_/A _73667_/X _73668_/Y sky130_fd_sc_hd__nand2_4
X_63421_ _63419_/Y _63391_/X _63420_/Y _63421_/Y sky130_fd_sc_hd__a21oi_4
X_75407_ _75403_/Y _75406_/Y _75407_/X sky130_fd_sc_hd__xor2_4
X_48355_ _50391_/A _48286_/X _48354_/X _48355_/X sky130_fd_sc_hd__and3_4
X_60633_ _60632_/X _60659_/A sky130_fd_sc_hd__buf_2
X_72619_ _72579_/A _72579_/B _65842_/X _72619_/Y sky130_fd_sc_hd__a21oi_4
X_79175_ _79171_/B _79171_/C _79175_/Y sky130_fd_sc_hd__nand2_4
X_45567_ _45567_/A _45597_/B _45567_/Y sky130_fd_sc_hd__nor2_4
X_76387_ _76387_/A _76387_/B _81618_/D sky130_fd_sc_hd__xor2_4
X_42779_ _42774_/X _42775_/X _41332_/X _87722_/Q _42750_/X _42779_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73599_ _73599_/A _73599_/B _73599_/Y sky130_fd_sc_hd__nor2_4
X_47306_ _47306_/A _52973_/B sky130_fd_sc_hd__buf_2
X_66140_ _66136_/Y _66137_/X _66139_/Y _84154_/D sky130_fd_sc_hd__a21o_4
X_78126_ _78119_/X _78125_/Y _78126_/Y sky130_fd_sc_hd__nand2_4
X_44518_ _44518_/A _44518_/Y sky130_fd_sc_hd__inv_2
X_75338_ _75334_/X _75339_/C _75337_/Y _75340_/A sky130_fd_sc_hd__a21o_4
X_63352_ _63305_/X _63392_/B _79158_/B _63352_/Y sky130_fd_sc_hd__nor3_4
X_48286_ _46485_/X _48286_/X sky130_fd_sc_hd__buf_2
X_60564_ _79139_/A _60132_/X _60562_/Y _60563_/X _60564_/X sky130_fd_sc_hd__a2bb2o_4
X_45498_ _45434_/X _61406_/A _45452_/X _45498_/Y sky130_fd_sc_hd__o21ai_4
X_62303_ _62301_/Y _62253_/X _62302_/Y _62303_/Y sky130_fd_sc_hd__a21oi_4
X_47237_ _47210_/A _47228_/B _47234_/X _52934_/D _47237_/X sky130_fd_sc_hd__and4_4
X_66071_ _64694_/A _73830_/B _66071_/X sky130_fd_sc_hd__and2_4
X_78057_ _84562_/Q _78057_/B _78057_/X sky130_fd_sc_hd__xor2_4
X_44449_ _44352_/X _44449_/X sky130_fd_sc_hd__buf_2
X_63283_ _63248_/X _63278_/Y _63279_/X _63280_/Y _63282_/Y _63283_/X
+ sky130_fd_sc_hd__a41o_4
X_75269_ _75269_/A _80944_/D _75269_/Y sky130_fd_sc_hd__nand2_4
X_60495_ _60476_/C _60570_/B _72590_/A _60495_/X sky130_fd_sc_hd__o21a_4
X_65022_ _64766_/A _65022_/X sky130_fd_sc_hd__buf_2
X_77008_ _77009_/A _82276_/D _77019_/A sky130_fd_sc_hd__nor2_4
X_62234_ _62362_/A _62234_/B _62229_/Y _62234_/D _62234_/Y sky130_fd_sc_hd__nand4_4
X_47168_ _86663_/Q _47145_/X _47167_/Y _47168_/Y sky130_fd_sc_hd__o21ai_4
X_46119_ _46119_/A _46120_/B sky130_fd_sc_hd__buf_2
X_69830_ _81966_/D _69763_/X _69829_/X _69830_/X sky130_fd_sc_hd__a21bo_4
X_62165_ _62157_/X _62159_/X _62164_/Y _84868_/Q _62117_/X _62165_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47099_ _53369_/B _52855_/B sky130_fd_sc_hd__buf_2
X_61116_ _64474_/A _64546_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_653_0_CLK clkbuf_9_326_0_CLK/X _87188_/CLK sky130_fd_sc_hd__clkbuf_1
X_69761_ _81971_/D _69696_/X _69760_/X _83899_/D sky130_fd_sc_hd__a21bo_4
X_66973_ _66972_/X _87618_/Q _66973_/X sky130_fd_sc_hd__and2_4
X_62096_ _84785_/Q _62128_/B _62128_/C _62060_/X _62096_/Y sky130_fd_sc_hd__nand4_4
X_78959_ _82643_/Q _78959_/Y sky130_fd_sc_hd__inv_2
X_68712_ _83964_/Q _68586_/X _68711_/X _68712_/X sky130_fd_sc_hd__a21bo_4
X_65924_ _65660_/A _65924_/X sky130_fd_sc_hd__buf_2
X_61047_ _61055_/A _61000_/X _76977_/A _61047_/X sky130_fd_sc_hd__or3_4
Xclkbuf_9_144_0_CLK clkbuf_8_72_0_CLK/X clkbuf_9_144_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_81970_ _81970_/CLK _83898_/Q _77732_/B sky130_fd_sc_hd__dfxtp_4
X_69692_ _44539_/A _69690_/X _69611_/X _69691_/X _69692_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_9_71_0_CLK clkbuf_9_71_0_CLK/A clkbuf_9_71_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_49809_ _49809_/A _53021_/B _49809_/Y sky130_fd_sc_hd__nand2_4
X_80921_ _84105_/CLK _80921_/D _75778_/A sky130_fd_sc_hd__dfxtp_4
X_68643_ _68639_/X _68642_/X _68442_/X _68647_/A sky130_fd_sc_hd__a21o_4
X_65855_ _65855_/A _65916_/B _65855_/C _65855_/X sky130_fd_sc_hd__and3_4
Xclkbuf_10_668_0_CLK clkbuf_9_334_0_CLK/X _88386_/CLK sky130_fd_sc_hd__clkbuf_1
X_52820_ _52515_/A _52821_/A sky130_fd_sc_hd__buf_2
X_64806_ _64806_/A _64807_/A sky130_fd_sc_hd__buf_2
X_83640_ _86424_/CLK _83640_/D _83640_/Q sky130_fd_sc_hd__dfxtp_4
X_80852_ _80854_/CLK _80852_/D _74989_/C sky130_fd_sc_hd__dfxtp_4
X_68574_ _68574_/A _68573_/X _68574_/Y sky130_fd_sc_hd__nand2_4
X_65786_ _65516_/X _65208_/Y _65785_/Y _65786_/Y sky130_fd_sc_hd__o21ai_4
X_62998_ _58403_/A _60493_/X _62998_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_9_159_0_CLK clkbuf_8_79_0_CLK/X clkbuf_9_159_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_67525_ _67497_/A _87723_/Q _67525_/X sky130_fd_sc_hd__and2_4
X_52751_ _52749_/Y _52728_/X _52750_/X _52751_/Y sky130_fd_sc_hd__a21oi_4
X_83571_ _86500_/CLK _71212_/Y _48602_/A sky130_fd_sc_hd__dfxtp_4
X_64737_ _64737_/A _64736_/Y _64737_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_2_2_2_CLK clkbuf_2_2_2_CLK/A clkbuf_2_2_2_CLK/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_9_86_0_CLK clkbuf_9_87_0_CLK/A clkbuf_9_86_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_61949_ _61949_/A _61949_/B _61949_/C _63168_/B _61949_/X sky130_fd_sc_hd__and4_4
X_80783_ _80849_/CLK _80783_/D _80783_/Q sky130_fd_sc_hd__dfxtp_4
X_85310_ _83001_/CLK _56024_/Y _55963_/B sky130_fd_sc_hd__dfxtp_4
X_51702_ _50222_/X _51717_/A sky130_fd_sc_hd__buf_2
X_82522_ _82711_/CLK _79021_/B _82522_/Q sky130_fd_sc_hd__dfxtp_4
X_55470_ _55470_/A _55470_/B _55470_/Y sky130_fd_sc_hd__nor2_4
X_67456_ _67364_/X _67456_/B _67456_/X sky130_fd_sc_hd__and2_4
X_86290_ _86610_/CLK _49970_/Y _72301_/B sky130_fd_sc_hd__dfxtp_4
X_52682_ _52678_/Y _52673_/X _52681_/X _52682_/Y sky130_fd_sc_hd__a21oi_4
X_64668_ _64767_/A _85822_/Q _64668_/X sky130_fd_sc_hd__and2_4
X_54421_ _54284_/A _54475_/A sky130_fd_sc_hd__buf_2
X_66407_ _66389_/A _66402_/B _66407_/C _66407_/Y sky130_fd_sc_hd__nor3_4
X_85241_ _85241_/CLK _56310_/Y _85241_/Q sky130_fd_sc_hd__dfxtp_4
X_51633_ _85974_/Q _51621_/X _51632_/Y _51633_/Y sky130_fd_sc_hd__o21ai_4
X_63619_ _58268_/A _60671_/C _62057_/D _63371_/A _63619_/X sky130_fd_sc_hd__a2bb2o_4
X_82453_ _82248_/CLK _79145_/X _82453_/Q sky130_fd_sc_hd__dfxtp_4
X_67387_ _67387_/A _67386_/X _67387_/Y sky130_fd_sc_hd__nand2_4
X_64599_ _64598_/X _64599_/X sky130_fd_sc_hd__buf_2
X_81404_ _81322_/CLK _81404_/D _76735_/B sky130_fd_sc_hd__dfxtp_4
X_57140_ _57140_/A _57140_/B _83322_/Q _57129_/Y _57141_/A sky130_fd_sc_hd__and4_4
X_69126_ _87476_/Q _69098_/X _69124_/X _69125_/X _69126_/X sky130_fd_sc_hd__a211o_4
X_54352_ _85458_/Q _54349_/X _54351_/Y _54352_/Y sky130_fd_sc_hd__o21ai_4
X_66338_ _66335_/X _66337_/X _64701_/X _66338_/X sky130_fd_sc_hd__a21o_4
X_85172_ _85168_/CLK _56502_/Y _56501_/C sky130_fd_sc_hd__dfxtp_4
X_51564_ _51562_/Y _51557_/X _51563_/X _51564_/Y sky130_fd_sc_hd__a21oi_4
X_82384_ _83703_/CLK _82192_/Q _47083_/A sky130_fd_sc_hd__dfxtp_4
X_53303_ _53293_/A _53293_/B _53302_/X _52785_/D _53303_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_606_0_CLK clkbuf_9_303_0_CLK/X _81954_/CLK sky130_fd_sc_hd__clkbuf_1
X_84123_ _84210_/CLK _84123_/D _66435_/A sky130_fd_sc_hd__dfxtp_4
X_50515_ _52218_/A _50526_/B _50526_/C _50515_/X sky130_fd_sc_hd__and3_4
X_57071_ _57179_/A _57071_/B _57071_/Y sky130_fd_sc_hd__nand2_4
X_81335_ _81352_/CLK _76469_/X _81711_/D sky130_fd_sc_hd__dfxtp_4
X_69057_ _69054_/X _69056_/X _69035_/X _69057_/X sky130_fd_sc_hd__a21o_4
X_54283_ _43177_/Y _54284_/A sky130_fd_sc_hd__buf_2
X_66269_ _66266_/X _86216_/Q _66180_/X _66268_/X _66269_/X sky130_fd_sc_hd__a211o_4
X_51495_ _51492_/Y _51477_/X _51494_/X _86000_/D sky130_fd_sc_hd__a21oi_4
X_56022_ _56142_/A _56023_/A sky130_fd_sc_hd__buf_2
X_68008_ _87895_/Q _68006_/X _67984_/X _68007_/X _68008_/X sky130_fd_sc_hd__a211o_4
X_53234_ _53217_/A _53244_/B _53222_/X _53234_/D _53234_/X sky130_fd_sc_hd__and4_4
X_84054_ _81492_/CLK _84054_/D _81486_/D sky130_fd_sc_hd__dfxtp_4
X_50446_ _86199_/Q _50437_/X _50445_/Y _50446_/Y sky130_fd_sc_hd__o21ai_4
X_81266_ _81362_/CLK _81298_/Q _81266_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_24_0_CLK clkbuf_9_25_0_CLK/A clkbuf_9_24_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_83005_ _85050_/CLK _83005_/D _83005_/Q sky130_fd_sc_hd__dfxtp_4
X_80217_ _80213_/X _80216_/Y _80244_/A sky130_fd_sc_hd__xor2_4
X_53165_ _53181_/A _53159_/B _53143_/X _53165_/D _53165_/X sky130_fd_sc_hd__and4_4
X_50377_ _50375_/Y _50351_/X _50376_/Y _50377_/Y sky130_fd_sc_hd__a21boi_4
X_81197_ _81197_/CLK _74978_/X _81197_/Q sky130_fd_sc_hd__dfxtp_4
X_52116_ _85885_/Q _52075_/X _52115_/Y _52116_/Y sky130_fd_sc_hd__o21ai_4
X_87813_ _87813_/CLK _87813_/D _87813_/Q sky130_fd_sc_hd__dfxtp_4
X_80148_ _80139_/Y _80135_/X _80147_/X _80149_/B sky130_fd_sc_hd__a21boi_4
X_57973_ _57868_/X _57971_/Y _57972_/Y _57899_/X _57872_/X _57973_/X
+ sky130_fd_sc_hd__o32a_4
X_53096_ _85698_/Q _53093_/X _53095_/Y _53096_/Y sky130_fd_sc_hd__o21ai_4
X_69959_ _88053_/Q _69468_/X _68745_/X _69958_/Y _69959_/X sky130_fd_sc_hd__a211o_4
X_59712_ _60403_/C _59790_/B _60414_/B _59710_/Y _59711_/Y _59712_/Y
+ sky130_fd_sc_hd__a41oi_4
X_52047_ _52014_/X _52047_/B _52047_/Y sky130_fd_sc_hd__nand2_4
X_56924_ _72718_/C _72718_/D _83314_/Q _56924_/X sky130_fd_sc_hd__a21o_4
X_87744_ _87748_/CLK _87744_/D _68848_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_39_0_CLK clkbuf_9_39_0_CLK/A clkbuf_9_39_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_72970_ _74140_/A _72970_/X sky130_fd_sc_hd__buf_2
X_84956_ _84892_/CLK _57676_/X _63524_/B sky130_fd_sc_hd__dfxtp_4
X_80079_ _84936_/Q _65698_/C _80079_/Y sky130_fd_sc_hd__nand2_4
X_71921_ _71586_/A _71930_/B _71574_/C _71921_/Y sky130_fd_sc_hd__nor3_4
X_59643_ _59635_/Y _59642_/X _59604_/X _59797_/B sky130_fd_sc_hd__and3_4
X_83907_ _83905_/CLK _83907_/D _83907_/Q sky130_fd_sc_hd__dfxtp_4
X_56855_ _56568_/X _57050_/A _56854_/X _56855_/Y sky130_fd_sc_hd__o21ai_4
X_87675_ _87675_/CLK _87675_/D _87675_/Q sky130_fd_sc_hd__dfxtp_4
X_84887_ _84921_/CLK _58289_/X _58287_/A sky130_fd_sc_hd__dfxtp_4
X_43820_ _43810_/X _43797_/X _41116_/X _87251_/Q _43811_/X _43821_/A
+ sky130_fd_sc_hd__o32ai_4
X_55806_ _85197_/Q _55342_/X _55457_/X _55805_/X _55806_/X sky130_fd_sc_hd__a211o_4
X_74640_ _74627_/Y _74685_/C sky130_fd_sc_hd__inv_2
X_86626_ _84922_/CLK _86626_/D _58136_/A sky130_fd_sc_hd__dfxtp_4
X_71852_ _71711_/A _71857_/D sky130_fd_sc_hd__buf_2
X_83838_ _83835_/CLK _70206_/X _83838_/Q sky130_fd_sc_hd__dfxtp_4
X_59574_ _59574_/A _60620_/C sky130_fd_sc_hd__buf_2
X_56786_ _56786_/A _56786_/Y sky130_fd_sc_hd__inv_2
X_53998_ _53998_/A _52478_/B _53998_/Y sky130_fd_sc_hd__nand2_4
X_70803_ _71221_/A _70804_/A sky130_fd_sc_hd__buf_2
X_58525_ _58517_/X _58522_/Y _58524_/Y _84828_/D sky130_fd_sc_hd__a21oi_4
X_43751_ _43602_/X _43752_/A sky130_fd_sc_hd__buf_2
X_55737_ _56280_/C _55278_/A _44043_/X _55736_/X _55737_/X sky130_fd_sc_hd__a211o_4
X_74571_ _74559_/X _74569_/X _56059_/Y _74570_/X _74571_/X sky130_fd_sc_hd__a211o_4
X_86557_ _86558_/CLK _48202_/Y _86557_/Q sky130_fd_sc_hd__dfxtp_4
X_40963_ _40931_/X _81724_/Q _40962_/X _40964_/A sky130_fd_sc_hd__o21ai_4
X_52949_ _52945_/Y _52946_/X _52948_/X _85725_/D sky130_fd_sc_hd__a21oi_4
X_71783_ _71783_/A _71507_/A _71783_/C _70361_/A _71783_/Y sky130_fd_sc_hd__nor4_4
X_83769_ _83476_/CLK _70465_/Y _58342_/A sky130_fd_sc_hd__dfxtp_4
X_76310_ _76296_/A _76295_/Y _76309_/X _76310_/Y sky130_fd_sc_hd__o21ai_4
X_42702_ _42701_/Y _42702_/Y sky130_fd_sc_hd__inv_2
X_73522_ _48694_/A _73521_/Y _73522_/X sky130_fd_sc_hd__xor2_4
X_85508_ _85507_/CLK _85508_/D _85508_/Q sky130_fd_sc_hd__dfxtp_4
X_46470_ _46423_/X _49077_/A _46469_/Y _46471_/A sky130_fd_sc_hd__o21ai_4
X_70734_ _70733_/Y _71263_/D sky130_fd_sc_hd__buf_2
X_58456_ _58510_/A _58474_/B sky130_fd_sc_hd__buf_2
X_77290_ _77318_/A _77290_/B _82182_/D sky130_fd_sc_hd__xnor2_4
X_55668_ _55288_/B _55288_/A _55287_/X _55669_/A sky130_fd_sc_hd__nand3_4
X_43682_ _87311_/Q _69622_/B sky130_fd_sc_hd__inv_2
X_86488_ _85879_/CLK _86488_/D _73012_/B sky130_fd_sc_hd__dfxtp_4
X_40894_ _40894_/A _40894_/X sky130_fd_sc_hd__buf_2
X_57407_ _55483_/Y _57391_/Y _44318_/A _56667_/Y _57407_/X sky130_fd_sc_hd__a2bb2o_4
X_45421_ _45415_/X _45418_/X _45420_/Y _86878_/D sky130_fd_sc_hd__a21oi_4
X_76241_ _76207_/Y _76221_/Y _76220_/Y _76241_/X sky130_fd_sc_hd__a21o_4
X_88227_ _88232_/CLK _88227_/D _67732_/B sky130_fd_sc_hd__dfxtp_4
X_54619_ _54625_/A _54607_/B _54618_/X _47227_/A _54619_/X sky130_fd_sc_hd__and4_4
X_42633_ _42680_/A _42634_/A sky130_fd_sc_hd__buf_2
X_73453_ _73449_/X _85574_/Q _73450_/X _73452_/X _73453_/X sky130_fd_sc_hd__a211o_4
X_85439_ _85439_/CLK _85439_/D _85439_/Q sky130_fd_sc_hd__dfxtp_4
X_70665_ _70534_/Y _70670_/A sky130_fd_sc_hd__buf_2
X_58387_ _58366_/X _83350_/Q _58386_/Y _84862_/D sky130_fd_sc_hd__o21a_4
X_55599_ _55908_/A _55599_/B _55599_/X sky130_fd_sc_hd__and2_4
X_48140_ _83531_/Q _48141_/A sky130_fd_sc_hd__inv_2
X_72404_ _72347_/A _86281_/Q _72404_/Y sky130_fd_sc_hd__nor2_4
X_45352_ _45350_/X _61673_/B _45294_/X _45352_/Y sky130_fd_sc_hd__o21ai_4
X_57338_ _57337_/Y _56659_/Y _56788_/X _57338_/Y sky130_fd_sc_hd__a21oi_4
X_76172_ _76171_/Y _76174_/A sky130_fd_sc_hd__inv_2
X_42564_ _87818_/Q _42564_/Y sky130_fd_sc_hd__inv_2
X_88158_ _88158_/CLK _88158_/D _67840_/B sky130_fd_sc_hd__dfxtp_4
X_73384_ _73380_/X _73382_/X _73383_/X _73384_/X sky130_fd_sc_hd__a21o_4
X_70596_ _52969_/B _70584_/X _70595_/Y _83745_/D sky130_fd_sc_hd__o21ai_4
X_44303_ _44231_/A _46228_/A sky130_fd_sc_hd__buf_2
X_75123_ _80773_/Q _75122_/A _80741_/D sky130_fd_sc_hd__xnor2_4
X_41515_ _41514_/X _41515_/X sky130_fd_sc_hd__buf_2
X_87109_ _87417_/CLK _44437_/Y _87109_/Q sky130_fd_sc_hd__dfxtp_4
X_48071_ _83538_/Q _57605_/B sky130_fd_sc_hd__inv_2
X_72335_ _72347_/A _86287_/Q _72335_/Y sky130_fd_sc_hd__nor2_4
X_45283_ _85256_/Q _45222_/X _45282_/X _45283_/Y sky130_fd_sc_hd__o21ai_4
X_57269_ _57268_/X _57149_/B _57149_/C _57149_/D _57271_/A sky130_fd_sc_hd__and4_4
X_88089_ _87588_/CLK _88089_/D _88089_/Q sky130_fd_sc_hd__dfxtp_4
X_42495_ _42610_/A _42495_/X sky130_fd_sc_hd__buf_2
X_59008_ _86688_/Q _59008_/B _59008_/Y sky130_fd_sc_hd__nor2_4
X_47022_ _47018_/Y _46987_/X _47021_/X _47022_/Y sky130_fd_sc_hd__a21oi_4
X_44234_ _73181_/A _72881_/A sky130_fd_sc_hd__buf_2
X_75054_ _80958_/Q _75053_/X _75054_/X sky130_fd_sc_hd__xor2_4
X_79931_ _79929_/Y _79931_/B _79932_/B sky130_fd_sc_hd__nand2_4
X_41446_ _41412_/X _82883_/Q _41445_/X _41446_/Y sky130_fd_sc_hd__o21ai_4
X_60280_ _60168_/A _60251_/A _60179_/A _60204_/A _60281_/A sky130_fd_sc_hd__and4_4
X_72266_ _72264_/X _85365_/Q _72265_/X _72266_/Y sky130_fd_sc_hd__o21ai_4
X_74005_ _74005_/A _74244_/B _74005_/Y sky130_fd_sc_hd__nor2_4
X_71217_ _71219_/A _71217_/B _71219_/C _71217_/Y sky130_fd_sc_hd__nand3_4
X_44165_ _64850_/A _64619_/A sky130_fd_sc_hd__buf_2
X_79862_ _64663_/C _83279_/Q _79862_/X sky130_fd_sc_hd__xor2_4
X_41377_ _41337_/X _41338_/X _41376_/X _67756_/B _41333_/X _41378_/A
+ sky130_fd_sc_hd__o32ai_4
X_72197_ _72196_/X _85339_/Q _72120_/X _72197_/X sky130_fd_sc_hd__o21a_4
X_43116_ _43105_/X _43106_/X _40771_/X _43115_/Y _43108_/X _87570_/D
+ sky130_fd_sc_hd__o32ai_4
X_78813_ _82835_/Q _78814_/A sky130_fd_sc_hd__inv_2
X_40328_ _40878_/A _40402_/A sky130_fd_sc_hd__buf_2
X_71148_ _48380_/X _71138_/X _71147_/Y _71148_/Y sky130_fd_sc_hd__o21ai_4
X_48973_ _48973_/A _52307_/B sky130_fd_sc_hd__buf_2
X_44096_ _44095_/X _44096_/X sky130_fd_sc_hd__buf_2
X_79793_ _79793_/A _79793_/B _79793_/X sky130_fd_sc_hd__xor2_4
X_47924_ _47912_/A _47924_/B _47924_/Y sky130_fd_sc_hd__nand2_4
X_43047_ _43047_/A _43047_/X sky130_fd_sc_hd__buf_2
X_78744_ _78742_/X _78718_/Y _78744_/C _78745_/A sky130_fd_sc_hd__and3_4
X_63970_ _60984_/A _64033_/D sky130_fd_sc_hd__buf_2
X_71079_ _48982_/X _71070_/X _71078_/Y _71079_/Y sky130_fd_sc_hd__o21ai_4
X_75956_ _75948_/Y _75949_/A _75954_/A _75956_/Y sky130_fd_sc_hd__nand3_4
X_62921_ _62930_/A _62930_/B _62921_/C _62921_/Y sky130_fd_sc_hd__nor3_4
X_74907_ _81131_/D _74916_/B _74910_/A sky130_fd_sc_hd__xor2_4
X_47855_ _47855_/A _50232_/B _47855_/Y sky130_fd_sc_hd__nand2_4
X_78675_ _78701_/B _78675_/B _82778_/D sky130_fd_sc_hd__xor2_4
X_75887_ _75887_/A _75887_/Y sky130_fd_sc_hd__inv_2
X_46806_ _46806_/A _46805_/X _46806_/Y sky130_fd_sc_hd__nand2_4
X_65640_ _65704_/A _86483_/Q _65640_/X sky130_fd_sc_hd__and2_4
X_77626_ _77596_/B _77622_/X _77625_/X _77626_/Y sky130_fd_sc_hd__a21boi_4
X_74838_ _46196_/A _74842_/B _46195_/Y _80670_/D sky130_fd_sc_hd__and3_4
X_62852_ _63306_/A _62852_/X sky130_fd_sc_hd__buf_2
X_47786_ _47782_/Y _47745_/X _47785_/X _86598_/D sky130_fd_sc_hd__a21oi_4
X_44998_ _45824_/B _44998_/X sky130_fd_sc_hd__buf_2
X_49525_ _49444_/A _49546_/A sky130_fd_sc_hd__buf_2
X_61803_ _61800_/Y _61801_/X _61802_/Y _61803_/Y sky130_fd_sc_hd__a21oi_4
X_46737_ _46737_/A _46717_/B _46717_/C _46736_/X _46737_/X sky130_fd_sc_hd__and4_4
X_65571_ _66044_/A _65631_/B _65570_/X _65571_/Y sky130_fd_sc_hd__nand3_4
X_77557_ _77553_/X _77558_/C _77556_/Y _77559_/A sky130_fd_sc_hd__a21o_4
X_43949_ _87180_/Q _43987_/B _43945_/Y _43948_/Y _43949_/X sky130_fd_sc_hd__a211o_4
X_62783_ _62819_/A _84830_/Q _62737_/X _62782_/X _62783_/X sky130_fd_sc_hd__and4_4
X_74769_ _74769_/A _74804_/C _74744_/X _74769_/D _74772_/B sky130_fd_sc_hd__nand4_4
X_67310_ _67307_/X _67309_/X _67264_/X _67316_/A sky130_fd_sc_hd__a21o_4
X_64522_ _58360_/A _64521_/X _64522_/Y sky130_fd_sc_hd__nor2_4
X_76508_ _76508_/A _76510_/B sky130_fd_sc_hd__inv_2
X_49456_ _49447_/A _49456_/B _49447_/C _46783_/X _49456_/X sky130_fd_sc_hd__and4_4
X_61734_ _58221_/X _61728_/X _62183_/D _59591_/A _61733_/X _61734_/X
+ sky130_fd_sc_hd__a41o_4
X_68290_ _82639_/D _68279_/X _68289_/X _83991_/D sky130_fd_sc_hd__a21bo_4
X_46668_ _82972_/Q _54298_/D sky130_fd_sc_hd__inv_2
X_77488_ _77488_/A _77488_/B _77488_/Y sky130_fd_sc_hd__nand2_4
X_48407_ _48407_/A _52119_/B sky130_fd_sc_hd__buf_2
X_67241_ _67241_/A _86810_/Q _67241_/X sky130_fd_sc_hd__and2_4
X_79227_ _79227_/A _82822_/D sky130_fd_sc_hd__inv_2
X_45619_ _45614_/X _45618_/X _45602_/X _45619_/X sky130_fd_sc_hd__a21o_4
X_76439_ _76459_/A _81526_/D _76439_/X sky130_fd_sc_hd__xor2_4
X_64453_ _84245_/Q _64429_/X _64452_/X _64453_/X sky130_fd_sc_hd__a21o_4
X_49387_ _49383_/Y _49378_/X _49386_/X _86397_/D sky130_fd_sc_hd__a21oi_4
X_61665_ _61292_/A _61665_/B _61675_/C _61665_/Y sky130_fd_sc_hd__nand3_4
X_46599_ _81186_/Q _46600_/B sky130_fd_sc_hd__inv_2
X_63404_ _63528_/A _63456_/A sky130_fd_sc_hd__buf_2
X_48338_ _48348_/A _52079_/B _48338_/Y sky130_fd_sc_hd__nand2_4
X_60616_ _60593_/B _60616_/B _60616_/Y sky130_fd_sc_hd__nor2_4
X_67172_ _67169_/X _67171_/X _67147_/X _67172_/X sky130_fd_sc_hd__a21o_4
X_79158_ _79158_/A _79158_/B _79158_/Y sky130_fd_sc_hd__nand2_4
X_64384_ _64267_/A _64384_/X sky130_fd_sc_hd__buf_2
X_61596_ _61340_/A _61611_/C sky130_fd_sc_hd__buf_2
X_66123_ _66123_/A _66004_/B _80481_/B _66123_/X sky130_fd_sc_hd__and3_4
X_78109_ _82566_/Q _78102_/B _78109_/Y sky130_fd_sc_hd__nand2_4
X_63335_ _63335_/A _63344_/B _60588_/X _63344_/D _63335_/X sky130_fd_sc_hd__or4_4
X_60547_ _60526_/A _60526_/B _79142_/A _60547_/Y sky130_fd_sc_hd__nor3_4
X_48269_ _50314_/A _48201_/B _48287_/C _48269_/X sky130_fd_sc_hd__and3_4
X_79089_ _79089_/A _82527_/D sky130_fd_sc_hd__inv_2
X_50300_ _50279_/X _50300_/B _50300_/Y sky130_fd_sc_hd__nand2_4
X_81120_ _81834_/CLK _79879_/X _81120_/Q sky130_fd_sc_hd__dfxtp_4
X_66054_ _65877_/A _66054_/X sky130_fd_sc_hd__buf_2
X_51280_ _51280_/A _46356_/X _51280_/Y sky130_fd_sc_hd__nand2_4
X_63266_ _63260_/Y _63261_/X _63263_/X _63265_/X _63242_/X _63266_/Y
+ sky130_fd_sc_hd__o41ai_4
X_60478_ _60465_/Y _60471_/X _60586_/A _60476_/Y _60477_/Y _60478_/Y
+ sky130_fd_sc_hd__a41oi_4
X_65005_ _64602_/A _65005_/X sky130_fd_sc_hd__buf_2
X_50231_ _50225_/Y _50227_/X _50230_/Y _50231_/Y sky130_fd_sc_hd__a21boi_4
X_62217_ _62215_/Y _62166_/X _62216_/Y _84425_/D sky130_fd_sc_hd__a21oi_4
X_81051_ _81082_/CLK _75451_/Y _81051_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_592_0_CLK clkbuf_9_296_0_CLK/X _81061_/CLK sky130_fd_sc_hd__clkbuf_1
X_63197_ _63191_/Y _63192_/X _63194_/X _63196_/X _63183_/X _63197_/Y
+ sky130_fd_sc_hd__o41ai_4
X_80002_ _80000_/X _80002_/B _80002_/X sky130_fd_sc_hd__xor2_4
X_69813_ _69810_/X _69813_/B _69813_/Y sky130_fd_sc_hd__nand2_4
X_50162_ _50113_/A _50162_/X sky130_fd_sc_hd__buf_2
X_62148_ _58201_/X _62105_/X _62065_/D _61948_/X _62147_/X _62148_/X
+ sky130_fd_sc_hd__a41o_4
X_84810_ _82973_/CLK _84810_/D _58653_/A sky130_fd_sc_hd__dfxtp_4
X_69744_ _69324_/Y _69732_/X _69733_/X _69743_/Y _69744_/X sky130_fd_sc_hd__a211o_4
X_50093_ _50599_/A _50599_/B _47848_/X _50093_/X sky130_fd_sc_hd__o21a_4
X_54970_ _85343_/Q _54967_/X _54969_/Y _54970_/Y sky130_fd_sc_hd__o21ai_4
X_66956_ _66956_/A _88131_/Q _66956_/X sky130_fd_sc_hd__and2_4
X_62079_ _62050_/X _62090_/B _78058_/B _62079_/Y sky130_fd_sc_hd__nor3_4
X_85790_ _84807_/CLK _85790_/D _85790_/Q sky130_fd_sc_hd__dfxtp_4
X_53921_ _53921_/A _53921_/X sky130_fd_sc_hd__buf_2
X_65907_ _65845_/X _86241_/Q _65904_/X _65906_/X _65907_/X sky130_fd_sc_hd__a211o_4
X_84741_ _83766_/CLK _84741_/D _84741_/Q sky130_fd_sc_hd__dfxtp_4
X_81953_ _82124_/CLK _78028_/X _77721_/A sky130_fd_sc_hd__dfxtp_4
X_69675_ _68386_/A _69687_/A sky130_fd_sc_hd__buf_2
X_66887_ _66912_/A _87622_/Q _66887_/X sky130_fd_sc_hd__and2_4
X_56640_ _56552_/Y _56753_/A sky130_fd_sc_hd__buf_2
X_80904_ _83933_/CLK _84080_/Q _75619_/A sky130_fd_sc_hd__dfxtp_4
X_68626_ _68757_/A _68626_/X sky130_fd_sc_hd__buf_2
X_87460_ _87149_/CLK _87460_/D _87460_/Q sky130_fd_sc_hd__dfxtp_4
X_53852_ _53848_/A _53852_/B _53852_/Y sky130_fd_sc_hd__nand2_4
X_65838_ _65835_/X _65837_/X _64574_/X _65838_/X sky130_fd_sc_hd__a21o_4
X_84672_ _84672_/CLK _60041_/Y _80153_/A sky130_fd_sc_hd__dfxtp_4
X_81884_ _81872_/CLK _78075_/X _81852_/D sky130_fd_sc_hd__dfxtp_4
X_86411_ _86733_/CLK _86411_/D _86411_/Q sky130_fd_sc_hd__dfxtp_4
X_52803_ _52803_/A _52803_/B _52803_/Y sky130_fd_sc_hd__nand2_4
X_83623_ _83623_/CLK _71056_/Y _83623_/Q sky130_fd_sc_hd__dfxtp_4
X_56571_ _56570_/Y _56571_/X sky130_fd_sc_hd__buf_2
X_80835_ _80835_/CLK _80835_/D _80835_/Q sky130_fd_sc_hd__dfxtp_4
X_68557_ _88108_/Q _68504_/X _68555_/X _68556_/Y _68557_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_530_0_CLK clkbuf_9_265_0_CLK/X _81352_/CLK sky130_fd_sc_hd__clkbuf_1
X_87391_ _87898_/CLK _43497_/Y _87391_/Q sky130_fd_sc_hd__dfxtp_4
X_53783_ _53781_/Y _53773_/X _53782_/X _53783_/Y sky130_fd_sc_hd__a21oi_4
X_65769_ _65769_/A _86507_/Q _65769_/X sky130_fd_sc_hd__and2_4
Xclkbuf_6_21_0_CLK clkbuf_6_21_0_CLK/A clkbuf_7_42_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_50995_ _86093_/Q _50992_/X _50994_/Y _50995_/Y sky130_fd_sc_hd__o21ai_4
X_58310_ _58328_/A _58310_/X sky130_fd_sc_hd__buf_2
X_55522_ _55489_/A _55522_/X sky130_fd_sc_hd__buf_2
X_67508_ _67270_/X _67508_/X sky130_fd_sc_hd__buf_2
X_86342_ _86342_/CLK _49686_/Y _59327_/B sky130_fd_sc_hd__dfxtp_4
X_52734_ _52708_/A _52746_/C sky130_fd_sc_hd__buf_2
X_59290_ _84754_/Q _59268_/X _59283_/X _59289_/X _84754_/D sky130_fd_sc_hd__a2bb2oi_4
X_83554_ _86554_/CLK _71262_/Y _47910_/A sky130_fd_sc_hd__dfxtp_4
X_80766_ _80991_/CLK _75514_/X _80766_/Q sky130_fd_sc_hd__dfxtp_4
X_68488_ _68376_/X _66524_/B _68478_/Y _68487_/Y _68488_/X sky130_fd_sc_hd__a211o_4
X_58241_ _64283_/C _58241_/X sky130_fd_sc_hd__buf_2
X_82505_ _82671_/CLK _78877_/A _78416_/A sky130_fd_sc_hd__dfxtp_4
X_55453_ _55311_/X _55453_/X sky130_fd_sc_hd__buf_2
X_67439_ _67082_/A _67513_/A sky130_fd_sc_hd__buf_2
X_86273_ _83623_/CLK _86273_/D _86273_/Q sky130_fd_sc_hd__dfxtp_4
X_52665_ _52648_/X _52661_/B _52654_/C _46775_/X _52665_/X sky130_fd_sc_hd__and4_4
X_83485_ _83482_/CLK _83485_/D _83485_/Q sky130_fd_sc_hd__dfxtp_4
X_80697_ _80697_/CLK _80729_/Q _75411_/A sky130_fd_sc_hd__dfxtp_4
XPHY_703 sky130_fd_sc_hd__decap_3
X_88012_ _88012_/CLK _42146_/X _88012_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_714 sky130_fd_sc_hd__decap_3
X_54404_ _54376_/A _54404_/X sky130_fd_sc_hd__buf_2
X_85224_ _85192_/CLK _56355_/Y _55748_/B sky130_fd_sc_hd__dfxtp_4
X_51616_ _51612_/Y _51613_/X _51615_/X _85978_/D sky130_fd_sc_hd__a21oi_4
X_70450_ _71650_/A _74533_/A _71194_/C _70450_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_545_0_CLK clkbuf_9_272_0_CLK/X _81755_/CLK sky130_fd_sc_hd__clkbuf_1
X_58172_ _84915_/Q _63081_/A sky130_fd_sc_hd__inv_2
X_82436_ _82436_/CLK _79128_/X _82436_/Q sky130_fd_sc_hd__dfxtp_4
X_55384_ _55384_/A _55384_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_6_36_0_CLK clkbuf_6_37_0_CLK/A clkbuf_6_36_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_52596_ _52590_/A _46650_/A _52596_/Y sky130_fd_sc_hd__nand2_4
X_57123_ _56893_/B _57193_/D _57086_/X _57123_/Y sky130_fd_sc_hd__a21oi_4
X_69109_ _60111_/X _69109_/X sky130_fd_sc_hd__buf_2
X_54335_ _54333_/Y _54311_/X _54334_/X _54335_/Y sky130_fd_sc_hd__a21oi_4
X_85155_ _85250_/CLK _85155_/D _55715_/B sky130_fd_sc_hd__dfxtp_4
X_51547_ _51629_/A _51553_/A sky130_fd_sc_hd__buf_2
X_70381_ DATA_TO_HASH[4] _70382_/A sky130_fd_sc_hd__buf_2
X_82367_ _84115_/CLK _77028_/X _82367_/Q sky130_fd_sc_hd__dfxtp_4
X_41300_ _81758_/Q _41292_/B _41300_/X sky130_fd_sc_hd__or2_4
X_72120_ _72255_/A _72120_/X sky130_fd_sc_hd__buf_2
X_84106_ _84111_/CLK _84106_/D _66524_/C sky130_fd_sc_hd__dfxtp_4
X_57054_ _57346_/C _57055_/A sky130_fd_sc_hd__inv_2
X_81318_ _84079_/CLK _76213_/X _81726_/D sky130_fd_sc_hd__dfxtp_4
X_42280_ _42279_/X _42275_/X _41520_/X _87943_/Q _42276_/X _42281_/A
+ sky130_fd_sc_hd__o32ai_4
X_54266_ _54320_/A _54266_/X sky130_fd_sc_hd__buf_2
X_85086_ _83008_/CLK _85086_/D _85086_/Q sky130_fd_sc_hd__dfxtp_4
X_51478_ _51504_/A _51494_/B sky130_fd_sc_hd__buf_2
X_82298_ _82343_/CLK _77170_/B _40800_/B sky130_fd_sc_hd__dfxtp_4
X_56005_ _56004_/X _56005_/X sky130_fd_sc_hd__buf_2
X_41231_ _41230_/X _41181_/X _68924_/B _41182_/X _88253_/D sky130_fd_sc_hd__a2bb2o_4
X_53217_ _53217_/A _53211_/B _53195_/X _53217_/D _53217_/X sky130_fd_sc_hd__and4_4
X_72051_ _71985_/A _72051_/X sky130_fd_sc_hd__buf_2
X_84037_ _81160_/CLK _68109_/X _84037_/Q sky130_fd_sc_hd__dfxtp_4
X_50429_ _50491_/A _50429_/X sky130_fd_sc_hd__buf_2
X_81249_ _85334_/CLK _81057_/Q _81249_/Q sky130_fd_sc_hd__dfxtp_4
X_54197_ _53436_/X _54197_/X sky130_fd_sc_hd__buf_2
X_71002_ _50832_/B _70983_/A _71001_/Y _83636_/D sky130_fd_sc_hd__o21ai_4
X_41162_ _41161_/X _41152_/X _68607_/B _41153_/X _88266_/D sky130_fd_sc_hd__a2bb2o_4
X_53148_ _53147_/X _53148_/B _53148_/Y sky130_fd_sc_hd__nand2_4
X_75810_ _75810_/A _75810_/B _75810_/C _75810_/Y sky130_fd_sc_hd__nand3_4
X_45970_ _40390_/Y _45963_/X _86834_/Q _45964_/X _86834_/D sky130_fd_sc_hd__a2bb2o_4
X_41093_ _41092_/Y _41093_/X sky130_fd_sc_hd__buf_2
X_53079_ _53077_/Y _53056_/X _53078_/X _53079_/Y sky130_fd_sc_hd__a21oi_4
X_57956_ _57781_/X _57952_/Y _57955_/Y _57893_/X _57795_/X _57956_/X
+ sky130_fd_sc_hd__o32a_4
X_76790_ _76790_/A _76790_/B _76790_/X sky130_fd_sc_hd__xor2_4
X_85988_ _85700_/CLK _85988_/D _85988_/Q sky130_fd_sc_hd__dfxtp_4
X_44921_ _44917_/Y _44920_/Y _44901_/X _44921_/X sky130_fd_sc_hd__o21a_4
X_56907_ _56906_/X _56907_/X sky130_fd_sc_hd__buf_2
X_75741_ _81012_/Q _75741_/B _80980_/D sky130_fd_sc_hd__xor2_4
X_87727_ _87472_/CLK _42770_/X _67437_/B sky130_fd_sc_hd__dfxtp_4
X_72953_ _88332_/Q _72803_/X _72776_/X _72953_/Y sky130_fd_sc_hd__o21ai_4
X_84939_ _84939_/CLK _57933_/Y _84939_/Q sky130_fd_sc_hd__dfxtp_4
X_57887_ _57773_/X _85718_/Q _44177_/X _57887_/X sky130_fd_sc_hd__o21a_4
X_47640_ _47639_/Y _53161_/B sky130_fd_sc_hd__buf_2
X_71904_ _57055_/A _71892_/X _71903_/Y _83334_/D sky130_fd_sc_hd__o21ai_4
X_59626_ _59664_/A _61755_/A sky130_fd_sc_hd__buf_2
X_78460_ _78460_/A _78460_/Y sky130_fd_sc_hd__inv_2
X_44852_ _44832_/X _44844_/X _41756_/X _67915_/B _44833_/X _44852_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56838_ _56838_/A _44135_/X _56837_/X _56838_/Y sky130_fd_sc_hd__nand3_4
X_75672_ _75665_/A _75665_/B _75666_/A _75672_/Y sky130_fd_sc_hd__a21boi_4
X_87658_ _86932_/CLK _42908_/X _67556_/B sky130_fd_sc_hd__dfxtp_4
X_72884_ _74383_/B _72884_/B _72884_/X sky130_fd_sc_hd__xor2_4
X_77411_ _77410_/Y _77412_/C sky130_fd_sc_hd__inv_2
X_43803_ _41064_/X _43801_/X _87260_/Q _43802_/X _87260_/D sky130_fd_sc_hd__a2bb2o_4
X_74623_ _58253_/A _74613_/X _56168_/A _74614_/X _74623_/X sky130_fd_sc_hd__a211o_4
X_86609_ _86611_/CLK _86609_/D _86609_/Q sky130_fd_sc_hd__dfxtp_4
X_47571_ _47525_/A _47574_/A sky130_fd_sc_hd__buf_2
X_71835_ _71829_/X _71839_/B _70778_/A _71826_/X _71835_/X sky130_fd_sc_hd__and4_4
X_59557_ _59557_/A _59557_/X sky130_fd_sc_hd__buf_2
X_78391_ _78375_/B _78391_/Y sky130_fd_sc_hd__inv_2
X_44783_ _44783_/A _44783_/Y sky130_fd_sc_hd__inv_2
X_56769_ _56768_/Y _57163_/C sky130_fd_sc_hd__buf_2
X_87589_ _88111_/CLK _87589_/D _73895_/A sky130_fd_sc_hd__dfxtp_4
X_41995_ _41982_/X _41993_/X _40792_/X _41994_/Y _41984_/X _88078_/D
+ sky130_fd_sc_hd__o32ai_4
X_49310_ _49302_/A _50832_/B _49310_/Y sky130_fd_sc_hd__nand2_4
X_46522_ _86729_/Q _46430_/X _46521_/Y _46522_/Y sky130_fd_sc_hd__o21ai_4
X_58508_ _58508_/A _58508_/Y sky130_fd_sc_hd__inv_2
X_77342_ _77341_/X _77342_/Y sky130_fd_sc_hd__inv_2
X_43734_ _43733_/X _87291_/D sky130_fd_sc_hd__inv_2
X_74554_ _74600_/A _74554_/X sky130_fd_sc_hd__buf_2
X_40946_ _40946_/A _40946_/X sky130_fd_sc_hd__buf_2
X_59488_ _83430_/Q _59488_/Y sky130_fd_sc_hd__inv_2
X_71766_ _71763_/X _71424_/C _70794_/X _71766_/X sky130_fd_sc_hd__and3_4
X_49241_ _49241_/A _49241_/B _49241_/Y sky130_fd_sc_hd__nand2_4
X_73505_ _73339_/A _73505_/B _73505_/Y sky130_fd_sc_hd__nor2_4
X_46453_ _50812_/A _46428_/B _46472_/C _46453_/X sky130_fd_sc_hd__and3_4
X_70717_ _70717_/A _70713_/X _70727_/C _70710_/D _70717_/Y sky130_fd_sc_hd__nand4_4
X_58439_ _58423_/X _83480_/Q _58438_/Y _58439_/X sky130_fd_sc_hd__o21a_4
X_77273_ _77270_/X _77274_/B _77272_/Y _77273_/X sky130_fd_sc_hd__a21o_4
X_43665_ _40734_/X _43656_/X _74166_/A _43657_/X _87321_/D sky130_fd_sc_hd__a2bb2o_4
X_74485_ _74490_/A _48639_/A _74485_/Y sky130_fd_sc_hd__nand2_4
X_40877_ _40365_/X _40877_/X sky130_fd_sc_hd__buf_2
X_71697_ _58283_/Y _71695_/X _71696_/Y _71697_/Y sky130_fd_sc_hd__o21ai_4
X_79012_ _79012_/A _79012_/Y sky130_fd_sc_hd__inv_2
X_45404_ _45403_/Y _45590_/B _45404_/X sky130_fd_sc_hd__and2_4
X_76224_ _76206_/Y _76211_/Y _76207_/Y _76225_/B sky130_fd_sc_hd__o21ai_4
X_42616_ _42614_/X _42615_/X _40909_/X _69917_/A _42597_/X _42616_/Y
+ sky130_fd_sc_hd__o32ai_4
X_61450_ _61342_/X _61451_/D sky130_fd_sc_hd__buf_2
X_49172_ _49172_/A _50710_/B sky130_fd_sc_hd__buf_2
X_73436_ _83151_/Q _73318_/X _73435_/Y _83151_/D sky130_fd_sc_hd__a21o_4
X_46384_ _46379_/Y _46346_/X _46383_/Y _46384_/Y sky130_fd_sc_hd__a21boi_4
X_70648_ _53025_/B _70632_/X _70647_/Y _83734_/D sky130_fd_sc_hd__o21ai_4
X_43596_ _43596_/A _68387_/B sky130_fd_sc_hd__inv_2
Xclkbuf_8_4_0_CLK clkbuf_8_5_0_CLK/A clkbuf_8_4_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_60401_ _60400_/Y _60472_/A sky130_fd_sc_hd__buf_2
X_48123_ _48122_/Y _48335_/B sky130_fd_sc_hd__buf_2
X_45335_ _45277_/X _61663_/B _45294_/X _45335_/Y sky130_fd_sc_hd__o21ai_4
X_76155_ _76155_/A _76155_/B _76155_/X sky130_fd_sc_hd__xor2_4
X_42547_ _42547_/A _42547_/X sky130_fd_sc_hd__buf_2
X_61381_ _64257_/A _61368_/B _61368_/C _61391_/D _61381_/Y sky130_fd_sc_hd__nand4_4
X_73367_ _73367_/A _73367_/X sky130_fd_sc_hd__buf_2
X_70579_ HASH_ADDR[3] _70356_/Y _70579_/Y sky130_fd_sc_hd__nor2_4
X_63120_ _60607_/A _63121_/D sky130_fd_sc_hd__buf_2
X_75106_ _75106_/A _75105_/Y _75107_/B sky130_fd_sc_hd__nor2_4
X_48054_ _66211_/B _48049_/X _48053_/Y _48054_/Y sky130_fd_sc_hd__o21ai_4
X_60332_ _60317_/A _60319_/X _79680_/A _60332_/Y sky130_fd_sc_hd__nor3_4
X_72318_ _72315_/Y _72317_/Y _72292_/X _72318_/X sky130_fd_sc_hd__a21o_4
X_45266_ _85161_/Q _45209_/X _45265_/X _45266_/X sky130_fd_sc_hd__o21a_4
X_76086_ _76096_/A _76097_/B _76086_/Y sky130_fd_sc_hd__nand2_4
X_42478_ _73750_/A _68567_/B sky130_fd_sc_hd__inv_2
X_73298_ _72829_/X _73298_/X sky130_fd_sc_hd__buf_2
X_47005_ _46909_/X _47008_/A sky130_fd_sc_hd__buf_2
X_44217_ _43959_/B _44217_/X sky130_fd_sc_hd__buf_2
X_63051_ _63041_/A _63051_/B _63030_/C _60541_/C _63051_/X sky130_fd_sc_hd__and4_4
X_75037_ _80956_/Q _75036_/X _75037_/X sky130_fd_sc_hd__xor2_4
X_79914_ _79912_/Y _79914_/B _79915_/B sky130_fd_sc_hd__nand2_4
X_41429_ _41428_/Y _41429_/X sky130_fd_sc_hd__buf_2
X_60263_ _60263_/A _60268_/A _60263_/C _60263_/Y sky130_fd_sc_hd__nor3_4
X_72249_ _72236_/Y _72237_/X _72244_/X _72248_/X _72249_/Y sky130_fd_sc_hd__a22oi_4
X_45197_ _45197_/A _45272_/A sky130_fd_sc_hd__buf_2
X_62002_ _62002_/A _62002_/B _78063_/B _62002_/Y sky130_fd_sc_hd__nor3_4
X_44148_ _44148_/A _44149_/A sky130_fd_sc_hd__buf_2
X_79845_ _84230_/Q _83278_/Q _79845_/X sky130_fd_sc_hd__xor2_4
X_60194_ _60239_/B _60253_/A sky130_fd_sc_hd__buf_2
X_66810_ _66785_/A _66810_/B _66810_/X sky130_fd_sc_hd__and2_4
X_48956_ _48964_/A _48955_/X _48956_/Y sky130_fd_sc_hd__nand2_4
X_44079_ _55817_/A _44079_/X sky130_fd_sc_hd__buf_2
X_67790_ _67790_/A _88160_/Q _67790_/X sky130_fd_sc_hd__and2_4
X_79776_ _79774_/X _79781_/B _79776_/Y sky130_fd_sc_hd__xnor2_4
X_76988_ _84540_/Q _84412_/Q _76988_/X sky130_fd_sc_hd__xor2_4
X_47907_ _47904_/X _82939_/Q _47906_/X _48212_/A sky130_fd_sc_hd__o21ai_4
X_66741_ _66669_/A _88140_/Q _66741_/X sky130_fd_sc_hd__and2_4
X_78727_ _78727_/A _78726_/Y _82493_/D sky130_fd_sc_hd__xnor2_4
X_75939_ _81508_/Q _75939_/B _75939_/Y sky130_fd_sc_hd__xnor2_4
X_63953_ _57672_/X _63902_/B _63902_/C _64016_/D _63954_/D sky130_fd_sc_hd__nand4_4
X_48887_ _83624_/Q _48887_/Y sky130_fd_sc_hd__inv_2
X_62904_ _62900_/X _62893_/X _62903_/Y _84372_/D sky130_fd_sc_hd__a21oi_4
X_69460_ _87016_/Q _69457_/X _69458_/X _69459_/X _69461_/B sky130_fd_sc_hd__a211o_4
X_47838_ _47832_/X _47838_/X sky130_fd_sc_hd__buf_2
X_66672_ _60781_/A _66672_/X sky130_fd_sc_hd__buf_2
X_78658_ _82521_/Q _82777_/D _82489_/D sky130_fd_sc_hd__xor2_4
X_63884_ _58506_/A _63900_/B _63900_/C _63900_/D _63884_/Y sky130_fd_sc_hd__nand4_4
X_68411_ _68407_/X _68410_/X _68331_/X _68411_/Y sky130_fd_sc_hd__a21oi_4
X_65623_ _64752_/A _65623_/X sky130_fd_sc_hd__buf_2
X_77609_ _77609_/A _82203_/D _81915_/D sky130_fd_sc_hd__xor2_4
X_62835_ _62717_/A _62880_/D sky130_fd_sc_hd__buf_2
X_69391_ _69329_/X _68822_/Y _69325_/X _69390_/Y _69391_/X sky130_fd_sc_hd__a211o_4
X_47769_ _47804_/A _47777_/B _47777_/C _53234_/D _47769_/X sky130_fd_sc_hd__and4_4
X_78589_ _78585_/Y _78587_/Y _78584_/Y _78589_/Y sky130_fd_sc_hd__o21ai_4
X_49508_ _49502_/A _51031_/B _49508_/Y sky130_fd_sc_hd__nand2_4
X_80620_ _80617_/Y _80600_/Y _80619_/X _80622_/A sky130_fd_sc_hd__o21ai_4
X_68342_ _68342_/A _69796_/A sky130_fd_sc_hd__buf_2
X_65554_ _65416_/X _72993_/B _65554_/X sky130_fd_sc_hd__and2_4
X_50780_ _50778_/Y _50768_/X _50779_/Y _50780_/Y sky130_fd_sc_hd__a21boi_4
X_62766_ _62766_/A _62766_/B _62766_/C _62766_/Y sky130_fd_sc_hd__nor3_4
X_64505_ _64455_/X _61637_/X _64211_/C _64505_/Y sky130_fd_sc_hd__nand3_4
X_49439_ _58750_/B _49415_/X _49438_/Y _49439_/Y sky130_fd_sc_hd__o21ai_4
X_61717_ _58403_/A _59858_/Y _61298_/B _61716_/X _61717_/X sky130_fd_sc_hd__a2bb2o_4
X_80551_ _80551_/A _80551_/B _80551_/Y sky130_fd_sc_hd__nand2_4
X_68273_ _67682_/X _67684_/X _68260_/X _68273_/Y sky130_fd_sc_hd__a21oi_4
X_65485_ _64567_/A _65486_/A sky130_fd_sc_hd__buf_2
X_62697_ _62673_/A _62673_/B _84390_/Q _62697_/Y sky130_fd_sc_hd__nor3_4
X_67224_ _87928_/Q _67176_/X _67153_/X _67223_/X _67224_/X sky130_fd_sc_hd__a211o_4
X_52450_ _50755_/A _52446_/B _52369_/X _52450_/X sky130_fd_sc_hd__and3_4
X_64436_ _61180_/A _64515_/A sky130_fd_sc_hd__buf_2
X_83270_ _83630_/CLK _83270_/D _83270_/Q sky130_fd_sc_hd__dfxtp_4
X_61648_ _72561_/C _61682_/C sky130_fd_sc_hd__buf_2
X_80482_ _80476_/A _80476_/B _80481_/Y _80482_/Y sky130_fd_sc_hd__a21boi_4
X_51401_ _51399_/Y _51229_/X _51400_/X _51401_/Y sky130_fd_sc_hd__a21oi_4
X_82221_ _82221_/CLK _82253_/Q _82221_/Q sky130_fd_sc_hd__dfxtp_4
X_67155_ _87931_/Q _67056_/X _67153_/X _67154_/X _67155_/X sky130_fd_sc_hd__a211o_4
X_52381_ _52385_/A _49121_/A _52381_/X sky130_fd_sc_hd__and2_4
X_64367_ _64367_/A _64367_/X sky130_fd_sc_hd__buf_2
X_61579_ _61329_/A _61579_/B _72549_/B _61579_/Y sky130_fd_sc_hd__nand3_4
X_54120_ _54116_/Y _54117_/X _54119_/X _85501_/D sky130_fd_sc_hd__a21oi_4
X_66106_ _66020_/X _66103_/Y _66105_/Y _66106_/Y sky130_fd_sc_hd__o21ai_4
X_51332_ _51259_/A _51332_/X sky130_fd_sc_hd__buf_2
X_63318_ _63315_/Y _63316_/X _63317_/X _63318_/X sky130_fd_sc_hd__a21o_4
X_82152_ _82152_/CLK _84144_/Q _82152_/Q sky130_fd_sc_hd__dfxtp_4
X_67086_ _67080_/X _67084_/X _67085_/X _67086_/X sky130_fd_sc_hd__a21o_4
X_64298_ _64293_/X _64294_/X _64295_/X _64297_/Y _64267_/X _64298_/X
+ sky130_fd_sc_hd__o41a_4
X_81103_ _80817_/CLK _79696_/Y _75839_/A sky130_fd_sc_hd__dfxtp_4
X_54051_ _53773_/A _54051_/X sky130_fd_sc_hd__buf_2
X_66037_ _65878_/A _66037_/B _66037_/X sky130_fd_sc_hd__and2_4
X_51263_ _51263_/A _51263_/X sky130_fd_sc_hd__buf_2
X_86960_ _88232_/CLK _86960_/D _86960_/Q sky130_fd_sc_hd__dfxtp_4
X_82083_ _81954_/CLK _82083_/D _82083_/Q sky130_fd_sc_hd__dfxtp_4
X_63249_ _60555_/A _61582_/A _60608_/X _61579_/B _63249_/Y sky130_fd_sc_hd__a22oi_4
X_53002_ _52893_/X _53019_/A sky130_fd_sc_hd__buf_2
X_50214_ _50473_/A _57489_/B _50213_/X _50214_/Y sky130_fd_sc_hd__nand3_4
X_85911_ _86554_/CLK _85911_/D _85911_/Q sky130_fd_sc_hd__dfxtp_4
X_81034_ _81065_/CLK _81034_/D _81034_/Q sky130_fd_sc_hd__dfxtp_4
X_51194_ _51184_/X _52885_/B _51194_/Y sky130_fd_sc_hd__nand2_4
X_86891_ _80672_/CLK _45221_/Y _63238_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_opt_22_CLK _86506_/CLK _86471_/CLK sky130_fd_sc_hd__clkbuf_16
X_57810_ _57801_/X _57807_/Y _57808_/Y _57700_/X _57809_/X _57810_/X
+ sky130_fd_sc_hd__o32a_4
X_50145_ _65084_/B _50137_/X _50144_/Y _50145_/Y sky130_fd_sc_hd__o21ai_4
X_85842_ _83303_/CLK _52342_/Y _85842_/Q sky130_fd_sc_hd__dfxtp_4
X_58790_ _58783_/Y _58789_/Y _58735_/X _58790_/X sky130_fd_sc_hd__a21o_4
X_67988_ _67914_/X _67988_/B _67988_/X sky130_fd_sc_hd__and2_4
X_57741_ _57726_/X _86015_/Q _57740_/X _57741_/Y sky130_fd_sc_hd__o21ai_4
X_69727_ _69727_/A _69727_/B _69727_/Y sky130_fd_sc_hd__nand2_4
X_50076_ _86269_/Q _50061_/X _50075_/Y _50076_/Y sky130_fd_sc_hd__o21ai_4
X_54953_ _53460_/A _47818_/A _54953_/Y sky130_fd_sc_hd__nand2_4
X_66939_ _87364_/Q _66915_/X _66863_/X _66938_/X _66939_/X sky130_fd_sc_hd__a211o_4
X_85773_ _85773_/CLK _52691_/Y _85773_/Q sky130_fd_sc_hd__dfxtp_4
X_82985_ _85096_/CLK _74687_/Y _82985_/Q sky130_fd_sc_hd__dfxtp_4
X_87512_ _87520_/CLK _43262_/Y _87512_/Q sky130_fd_sc_hd__dfxtp_4
X_53904_ _53898_/A _72077_/B _53904_/Y sky130_fd_sc_hd__nand2_4
X_84724_ _83464_/CLK _84724_/D _84724_/Q sky130_fd_sc_hd__dfxtp_4
X_57672_ _63524_/B _57672_/X sky130_fd_sc_hd__buf_2
X_81936_ _81985_/CLK _77866_/Y _77441_/A sky130_fd_sc_hd__dfxtp_4
X_69658_ _83907_/Q _69632_/X _69657_/X _83907_/D sky130_fd_sc_hd__a21bo_4
X_54884_ _54881_/Y _54882_/X _54883_/X _85360_/D sky130_fd_sc_hd__a21oi_4
X_59411_ _59411_/A _59399_/B _59411_/Y sky130_fd_sc_hd__nand2_4
X_56623_ _55526_/X _55536_/D _72662_/C sky130_fd_sc_hd__and2_4
X_68609_ _68606_/X _68608_/X _68512_/X _68609_/Y sky130_fd_sc_hd__a21oi_4
X_87443_ _87888_/CLK _87443_/D _87443_/Q sky130_fd_sc_hd__dfxtp_4
X_53835_ _53833_/Y _53799_/X _53834_/Y _53835_/Y sky130_fd_sc_hd__a21boi_4
X_84655_ _84672_/CLK _84655_/D _60136_/C sky130_fd_sc_hd__dfxtp_4
X_81867_ _82220_/CLK _78058_/X _81867_/Q sky130_fd_sc_hd__dfxtp_4
X_69589_ _69152_/X _69155_/X _69575_/X _69589_/Y sky130_fd_sc_hd__a21oi_4
X_40800_ _40817_/A _40800_/B _40800_/X sky130_fd_sc_hd__or2_4
X_83606_ _85554_/CLK _83606_/D _49072_/A sky130_fd_sc_hd__dfxtp_4
X_59342_ _59133_/A _59342_/X sky130_fd_sc_hd__buf_2
X_71620_ _71865_/A _70667_/A _71614_/C _71622_/D _71620_/Y sky130_fd_sc_hd__nor4_4
X_56554_ _55536_/X _56580_/B sky130_fd_sc_hd__buf_2
X_80818_ _80818_/CLK _80818_/D _80818_/Q sky130_fd_sc_hd__dfxtp_4
X_41780_ _82884_/Q _46240_/A _41780_/X sky130_fd_sc_hd__or2_4
X_87374_ _87373_/CLK _87374_/D _87374_/Q sky130_fd_sc_hd__dfxtp_4
X_53766_ _53766_/A _48683_/A _53766_/Y sky130_fd_sc_hd__nand2_4
X_84586_ _84590_/CLK _60613_/Y _60612_/C sky130_fd_sc_hd__dfxtp_4
X_50978_ _50952_/A _50985_/C sky130_fd_sc_hd__buf_2
X_81798_ _81671_/CLK _81606_/Q _47485_/A sky130_fd_sc_hd__dfxtp_4
X_55505_ _44063_/X _55505_/X sky130_fd_sc_hd__buf_2
X_86325_ _86322_/CLK _86325_/D _57897_/B sky130_fd_sc_hd__dfxtp_4
X_40731_ _40585_/A _40731_/X sky130_fd_sc_hd__buf_2
X_52717_ _52714_/Y _52702_/X _52716_/X _52717_/Y sky130_fd_sc_hd__a21oi_4
X_59273_ _58877_/A _59273_/X sky130_fd_sc_hd__buf_2
X_71551_ _71530_/Y _83459_/Q _71550_/Y _83459_/D sky130_fd_sc_hd__a21o_4
X_83537_ _86218_/CLK _83537_/D _83537_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_484_0_CLK clkbuf_9_242_0_CLK/X _85679_/CLK sky130_fd_sc_hd__clkbuf_1
X_56485_ _56474_/X _56484_/X _85178_/Q _56485_/Y sky130_fd_sc_hd__nand3_4
X_80749_ _81125_/CLK _80749_/D _81125_/D sky130_fd_sc_hd__dfxtp_4
X_53697_ _48533_/A _53697_/B _53697_/C _53697_/Y sky130_fd_sc_hd__nand3_4
X_58224_ _58224_/A _58224_/Y sky130_fd_sc_hd__inv_2
X_70502_ _70502_/A _70502_/Y sky130_fd_sc_hd__inv_2
XPHY_500 sky130_fd_sc_hd__decap_3
X_43450_ _43449_/X _43426_/X _41606_/X _87415_/Q _43434_/X _43450_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55436_ _55383_/A _55377_/Y _55379_/Y _55436_/Y sky130_fd_sc_hd__nand3_4
X_86256_ _86256_/CLK _86256_/D _65061_/B sky130_fd_sc_hd__dfxtp_4
X_74270_ _86976_/Q _73916_/B _74269_/X _74281_/C sky130_fd_sc_hd__o21ai_4
XPHY_511 sky130_fd_sc_hd__decap_3
X_40662_ _40635_/X _40638_/X _40661_/X _68699_/B _40612_/X _40663_/A
+ sky130_fd_sc_hd__o32ai_4
X_52648_ _52648_/A _52648_/X sky130_fd_sc_hd__buf_2
X_83468_ _85955_/CLK _83468_/D _47797_/A sky130_fd_sc_hd__dfxtp_4
X_71482_ _71463_/Y _83483_/Q _71481_/X _83483_/D sky130_fd_sc_hd__a21o_4
XPHY_522 sky130_fd_sc_hd__decap_3
XPHY_533 sky130_fd_sc_hd__decap_3
X_42401_ _42417_/A _42401_/X sky130_fd_sc_hd__buf_2
XPHY_544 sky130_fd_sc_hd__decap_3
X_73221_ _74140_/A _73221_/X sky130_fd_sc_hd__buf_2
X_85207_ _85269_/CLK _85207_/D _85207_/Q sky130_fd_sc_hd__dfxtp_4
X_70433_ _70442_/A _70374_/X _70431_/C _70433_/Y sky130_fd_sc_hd__nand3_4
X_58155_ _63033_/A _63389_/A sky130_fd_sc_hd__buf_2
XPHY_555 sky130_fd_sc_hd__decap_3
X_82419_ _82820_/CLK _82419_/D _78549_/A sky130_fd_sc_hd__dfxtp_4
X_43381_ _41416_/X _43371_/X _87451_/Q _43372_/X _43381_/X sky130_fd_sc_hd__a2bb2o_4
X_55367_ _55392_/B _55392_/A _55367_/Y sky130_fd_sc_hd__nand2_4
X_86187_ _86505_/CLK _86187_/D _86187_/Q sky130_fd_sc_hd__dfxtp_4
X_40593_ _48903_/A _48192_/A sky130_fd_sc_hd__inv_2
X_52579_ _52605_/A _52594_/B sky130_fd_sc_hd__buf_2
XPHY_566 sky130_fd_sc_hd__decap_3
X_83399_ _84939_/CLK _83399_/D _58224_/A sky130_fd_sc_hd__dfxtp_4
XPHY_577 sky130_fd_sc_hd__decap_3
X_45120_ _44895_/X _45120_/X sky130_fd_sc_hd__buf_2
XPHY_588 sky130_fd_sc_hd__decap_3
X_57106_ _57105_/Y _57106_/X sky130_fd_sc_hd__buf_2
X_42332_ _42331_/Y _87918_/D sky130_fd_sc_hd__inv_2
X_54318_ _54325_/A _54325_/B _54317_/X _46706_/Y _54318_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_499_0_CLK clkbuf_9_249_0_CLK/X _83676_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_599 sky130_fd_sc_hd__decap_3
X_73152_ _44270_/X _73152_/X sky130_fd_sc_hd__buf_2
X_85138_ _85138_/CLK _85138_/D _85138_/Q sky130_fd_sc_hd__dfxtp_4
X_70364_ _70364_/A _70364_/X sky130_fd_sc_hd__buf_2
X_58086_ _58030_/X _85478_/Q _58062_/X _58086_/X sky130_fd_sc_hd__o21a_4
X_55298_ _55298_/A _55417_/A _55297_/X _55400_/A _55298_/X sky130_fd_sc_hd__and4_4
X_72103_ _74391_/A _50714_/B _72103_/Y sky130_fd_sc_hd__nand2_4
X_45051_ _45819_/A _45350_/A sky130_fd_sc_hd__buf_2
X_57037_ _56787_/X _56788_/A _57024_/D _57038_/B sky130_fd_sc_hd__nand3_4
X_42263_ _42262_/Y _42263_/Y sky130_fd_sc_hd__inv_2
X_54249_ _54249_/A _54249_/X sky130_fd_sc_hd__buf_2
X_77960_ _77950_/B _77950_/A _77960_/C _77960_/Y sky130_fd_sc_hd__nand3_4
X_73083_ _73083_/A _73198_/B _73083_/Y sky130_fd_sc_hd__nor2_4
X_85069_ _85103_/CLK _85069_/D _85069_/Q sky130_fd_sc_hd__dfxtp_4
X_70295_ _70289_/X _83807_/Q _70294_/X _83807_/D sky130_fd_sc_hd__a21o_4
X_44002_ _62640_/C _62975_/D sky130_fd_sc_hd__buf_2
X_41214_ _41213_/X _41214_/X sky130_fd_sc_hd__buf_2
X_72034_ _72025_/A _53858_/B _72034_/Y sky130_fd_sc_hd__nand2_4
X_76911_ _76893_/A _76897_/Y _76899_/A _76911_/Y sky130_fd_sc_hd__a21oi_4
X_42194_ _41294_/X _42192_/X _87986_/Q _42193_/X _87986_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_10_422_0_CLK clkbuf_9_211_0_CLK/X _82828_/CLK sky130_fd_sc_hd__clkbuf_1
X_77891_ _77891_/A _77890_/Y _77892_/A sky130_fd_sc_hd__xor2_4
X_48810_ _48837_/A _48831_/A sky130_fd_sc_hd__buf_2
Xclkbuf_opt_13_CLK _84914_/CLK _84716_/CLK sky130_fd_sc_hd__clkbuf_16
X_79630_ _79630_/A _79629_/X _79630_/X sky130_fd_sc_hd__xor2_4
X_41145_ _81723_/Q _41145_/B _41145_/X sky130_fd_sc_hd__or2_4
X_76842_ _76829_/A _76828_/Y _76842_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_4_14_1_CLK clkbuf_4_14_1_CLK/A clkbuf_4_14_1_CLK/X sky130_fd_sc_hd__clkbuf_1
X_49790_ _49786_/Y _49787_/X _49789_/X _86323_/D sky130_fd_sc_hd__a21oi_4
X_58988_ _58987_/Y _58988_/B _58988_/Y sky130_fd_sc_hd__nand2_4
X_48741_ _48737_/A _52128_/B _48741_/Y sky130_fd_sc_hd__nand2_4
X_79561_ _79558_/Y _79548_/Y _79561_/Y sky130_fd_sc_hd__nand2_4
X_45953_ _45948_/Y _45950_/Y _45952_/X _86840_/D sky130_fd_sc_hd__o21a_4
X_41076_ _41076_/A _41076_/X sky130_fd_sc_hd__buf_2
X_57939_ _58618_/A _57939_/X sky130_fd_sc_hd__buf_2
X_76773_ _76773_/A _76773_/B _76773_/Y sky130_fd_sc_hd__xnor2_4
X_73985_ _73985_/A _73024_/B _73985_/Y sky130_fd_sc_hd__nor2_4
X_78512_ _78511_/X _78519_/A sky130_fd_sc_hd__inv_2
X_44904_ _44904_/A _44975_/A sky130_fd_sc_hd__buf_2
X_75724_ _81010_/Q _75724_/B _75724_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_10_437_0_CLK clkbuf_9_218_0_CLK/X _83550_/CLK sky130_fd_sc_hd__clkbuf_1
X_48672_ _48672_/A _48673_/B sky130_fd_sc_hd__buf_2
X_60950_ _64182_/D _60901_/A _60934_/X _60950_/Y sky130_fd_sc_hd__nor3_4
X_72936_ _72755_/X _83075_/Q _72785_/X _72935_/X _72936_/X sky130_fd_sc_hd__a211o_4
X_79492_ _84815_/Q _84135_/Q _79494_/A sky130_fd_sc_hd__xor2_4
X_45884_ _45884_/A _45884_/Y sky130_fd_sc_hd__inv_2
X_47623_ _47623_/A _53153_/B sky130_fd_sc_hd__buf_2
X_59609_ _59571_/B _59571_/C _59516_/A _59609_/D _59609_/X sky130_fd_sc_hd__and4_4
X_78443_ _78441_/X _78443_/B _82763_/D sky130_fd_sc_hd__xor2_4
X_44835_ _44835_/A _86929_/D sky130_fd_sc_hd__inv_2
X_75655_ _81003_/Q _75655_/B _75655_/X sky130_fd_sc_hd__xor2_4
X_60881_ _64102_/B _60881_/B _60880_/X _60881_/Y sky130_fd_sc_hd__nand3_4
X_72867_ _69627_/B _72865_/X _72866_/X _72867_/X sky130_fd_sc_hd__o21a_4
X_62620_ _62620_/A _63703_/B _62532_/X _62622_/C sky130_fd_sc_hd__nand3_4
X_74606_ _74605_/X _74599_/X _56134_/A _74600_/X _74606_/X sky130_fd_sc_hd__a211o_4
X_47554_ _72162_/A _47524_/X _47553_/Y _47554_/Y sky130_fd_sc_hd__o21ai_4
X_71818_ _71804_/Y _83364_/Q _71817_/X _83364_/D sky130_fd_sc_hd__a21o_4
X_78374_ _78375_/A _78375_/C _78375_/B _78374_/X sky130_fd_sc_hd__a21o_4
X_44766_ _44528_/A _44766_/X sky130_fd_sc_hd__buf_2
X_75586_ _75586_/A _75585_/Y _75587_/B sky130_fd_sc_hd__xnor2_4
X_41978_ _41960_/X _41951_/X _40762_/X _88084_/Q _41953_/X _41978_/Y
+ sky130_fd_sc_hd__o32ai_4
X_72798_ _44130_/X _72798_/X sky130_fd_sc_hd__buf_2
X_46505_ _46505_/A _49110_/A _46505_/Y sky130_fd_sc_hd__nand2_4
X_77325_ _77325_/A _77325_/Y sky130_fd_sc_hd__inv_2
X_43717_ _43717_/A _69808_/B sky130_fd_sc_hd__inv_2
X_62551_ _62671_/A _62551_/X sky130_fd_sc_hd__buf_2
X_74537_ _74600_/A _74537_/Y sky130_fd_sc_hd__inv_2
X_40929_ _40929_/A _40929_/X sky130_fd_sc_hd__buf_2
X_71749_ _71175_/A _71753_/B _71744_/C _71744_/D _71749_/Y sky130_fd_sc_hd__nand4_4
X_47485_ _47485_/A _47486_/A sky130_fd_sc_hd__inv_2
X_44697_ _44697_/A _44697_/Y sky130_fd_sc_hd__inv_2
X_61502_ _61502_/A _61468_/B _61467_/X _61451_/D _61502_/Y sky130_fd_sc_hd__nand4_4
X_49224_ _49241_/A _50744_/B _49224_/Y sky130_fd_sc_hd__nand2_4
X_46436_ _46436_/A _46459_/B _46436_/X sky130_fd_sc_hd__or2_4
X_65270_ _65225_/A _65270_/B _65270_/X sky130_fd_sc_hd__and2_4
X_77256_ _77245_/C _77239_/C _77258_/A sky130_fd_sc_hd__nand2_4
X_43648_ _87327_/Q _68861_/B sky130_fd_sc_hd__inv_2
X_62482_ _61412_/A _62671_/A sky130_fd_sc_hd__buf_2
X_74468_ _46347_/A _50503_/B _74468_/Y sky130_fd_sc_hd__nand2_4
X_64221_ _64221_/A _64221_/X sky130_fd_sc_hd__buf_2
X_76207_ _76205_/Y _76202_/X _76219_/A _76207_/Y sky130_fd_sc_hd__nand3_4
X_49155_ _49416_/A _49205_/A sky130_fd_sc_hd__buf_2
X_61433_ _61427_/Y _61429_/Y _61403_/X _61430_/Y _61432_/Y _61433_/X
+ sky130_fd_sc_hd__a41o_4
X_73419_ _73416_/X _73418_/X _73347_/X _73434_/B sky130_fd_sc_hd__a21o_4
X_46367_ _83647_/Q _46367_/Y sky130_fd_sc_hd__inv_2
X_77187_ _82011_/Q _82299_/D _77187_/Y sky130_fd_sc_hd__nor2_4
X_43579_ _40542_/X _53455_/A _87349_/Q _43185_/A _43579_/X sky130_fd_sc_hd__a2bb2o_4
X_74399_ _83074_/Q _74377_/X _74398_/Y _74399_/Y sky130_fd_sc_hd__o21ai_4
X_48106_ _53588_/B _50365_/B sky130_fd_sc_hd__buf_2
X_45318_ _83014_/Q _45319_/A sky130_fd_sc_hd__inv_2
X_64152_ _64147_/X _64048_/X _64149_/Y _64150_/Y _64151_/X _64152_/X
+ sky130_fd_sc_hd__a41o_4
X_76138_ _81727_/D _76139_/B _76138_/Y sky130_fd_sc_hd__nor2_4
X_49086_ _48985_/A _49086_/X sky130_fd_sc_hd__buf_2
X_61364_ _61329_/A _61364_/B _61375_/C _61364_/Y sky130_fd_sc_hd__nand3_4
X_46298_ _46298_/A _46653_/A sky130_fd_sc_hd__buf_2
X_63103_ _63103_/A _63081_/B _63103_/C _63092_/D _63103_/X sky130_fd_sc_hd__or4_4
X_48037_ _48287_/A _48069_/B _47919_/X _48037_/X sky130_fd_sc_hd__and3_4
X_60315_ _60198_/Y _60174_/X _60241_/A _60313_/Y _60314_/Y _60315_/X
+ sky130_fd_sc_hd__a41o_4
X_45249_ _45242_/X _45246_/Y _45248_/Y _45249_/Y sky130_fd_sc_hd__a21oi_4
X_64083_ _61582_/A _60967_/A _64082_/Y _64083_/X sky130_fd_sc_hd__a21o_4
X_68960_ _74123_/A _68958_/X _68494_/X _68959_/Y _68960_/X sky130_fd_sc_hd__a211o_4
X_76069_ _81526_/Q _76069_/B _76069_/X sky130_fd_sc_hd__xor2_4
X_61295_ _61295_/A _72540_/B _61302_/A sky130_fd_sc_hd__nor2_4
X_67911_ _67905_/X _67911_/B _67911_/Y sky130_fd_sc_hd__nand2_4
X_63034_ _63031_/Y _63033_/X _61194_/X _63034_/Y sky130_fd_sc_hd__a21oi_4
X_60246_ _59043_/A _60246_/X sky130_fd_sc_hd__buf_2
X_68891_ _44245_/A _68891_/X sky130_fd_sc_hd__buf_2
X_79828_ _79840_/A _79827_/Y _79828_/Y sky130_fd_sc_hd__xnor2_4
X_67842_ _67842_/A _67842_/B _67842_/Y sky130_fd_sc_hd__nand2_4
X_60177_ _60174_/X _61316_/A _60177_/X sky130_fd_sc_hd__and2_4
X_49988_ _50001_/A _53200_/B _49988_/Y sky130_fd_sc_hd__nand2_4
X_48939_ _48635_/A _48940_/B sky130_fd_sc_hd__buf_2
X_67773_ _67678_/X _67773_/B _67773_/X sky130_fd_sc_hd__and2_4
X_79759_ _79745_/Y _79750_/Y _79758_/X _79760_/B sky130_fd_sc_hd__o21ai_4
X_64985_ _64752_/X _86163_/Q _64902_/X _64984_/X _64985_/X sky130_fd_sc_hd__a211o_4
X_69512_ _69223_/A _69586_/A sky130_fd_sc_hd__buf_2
X_66724_ _66819_/A _86832_/Q _66724_/X sky130_fd_sc_hd__and2_4
X_51950_ _52618_/A _52486_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_64_0_CLK clkbuf_8_65_0_CLK/A clkbuf_8_64_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_63936_ _60926_/X _64015_/D sky130_fd_sc_hd__buf_2
X_82770_ _82961_/CLK _82770_/D _82770_/Q sky130_fd_sc_hd__dfxtp_4
X_50901_ _86110_/Q _50882_/X _50900_/Y _50901_/Y sky130_fd_sc_hd__o21ai_4
X_81721_ _81412_/CLK _81721_/D _81721_/Q sky130_fd_sc_hd__dfxtp_4
X_69443_ _69288_/A _69443_/B _69443_/X sky130_fd_sc_hd__and2_4
X_66655_ _66652_/X _66654_/X _66606_/X _66655_/X sky130_fd_sc_hd__a21o_4
X_51881_ _85929_/Q _51873_/X _51880_/Y _51881_/Y sky130_fd_sc_hd__o21ai_4
X_63867_ _61430_/A _63853_/B _63803_/C _63866_/X _63867_/Y sky130_fd_sc_hd__nand4_4
X_53620_ _53620_/A _53620_/B _53620_/C _53620_/X sky130_fd_sc_hd__and3_4
X_65606_ _65601_/Y _65602_/X _65605_/Y _65606_/X sky130_fd_sc_hd__a21o_4
X_84440_ _82221_/CLK _84440_/D _78063_/B sky130_fd_sc_hd__dfxtp_4
X_50832_ _50822_/A _50832_/B _50832_/Y sky130_fd_sc_hd__nand2_4
X_62818_ _60211_/A _62818_/X sky130_fd_sc_hd__buf_2
X_81652_ _81330_/CLK _81684_/Q _81652_/Q sky130_fd_sc_hd__dfxtp_4
X_69374_ _69370_/X _69373_/X _69138_/X _69374_/X sky130_fd_sc_hd__a21o_4
X_66586_ _66526_/X _66559_/Y _59782_/X _66585_/Y _66586_/X sky130_fd_sc_hd__a211o_4
X_63798_ _63765_/A _61368_/A _63765_/C _63798_/X sky130_fd_sc_hd__and3_4
X_80603_ _80587_/X _80589_/B _80602_/Y _80607_/A sky130_fd_sc_hd__a21boi_4
X_68325_ _83982_/Q _68318_/X _68324_/X _83982_/D sky130_fd_sc_hd__a21bo_4
Xclkbuf_8_79_0_CLK clkbuf_8_79_0_CLK/A clkbuf_8_79_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_65537_ _65592_/A _72960_/B _65537_/X sky130_fd_sc_hd__and2_4
X_53551_ _53549_/Y _53524_/X _53550_/Y _85615_/D sky130_fd_sc_hd__a21boi_4
X_84371_ _84449_/CLK _84371_/D _84371_/Q sky130_fd_sc_hd__dfxtp_4
X_50763_ _50718_/A _50764_/A sky130_fd_sc_hd__buf_2
X_81583_ _83918_/CLK _65713_/C _76771_/A sky130_fd_sc_hd__dfxtp_4
X_62749_ _60217_/A _62749_/X sky130_fd_sc_hd__buf_2
X_86110_ _84807_/CLK _50905_/Y _86110_/Q sky130_fd_sc_hd__dfxtp_4
X_52502_ _52501_/X _46433_/A _52502_/Y sky130_fd_sc_hd__nand2_4
X_83322_ _83322_/CLK _71937_/Y _83322_/Q sky130_fd_sc_hd__dfxtp_4
X_56270_ _56194_/X _56270_/B _56270_/C _56270_/Y sky130_fd_sc_hd__nand3_4
X_80534_ _80512_/Y _80530_/X _80533_/Y _80534_/Y sky130_fd_sc_hd__a21oi_4
X_68256_ _68254_/X _67577_/Y _68247_/X _68255_/Y _68256_/X sky130_fd_sc_hd__a211o_4
X_87090_ _88267_/CLK _44473_/X _87090_/Q sky130_fd_sc_hd__dfxtp_4
X_53482_ _53478_/A _73692_/A _53482_/Y sky130_fd_sc_hd__nand2_4
X_65468_ _65401_/A _72836_/B _65468_/X sky130_fd_sc_hd__and2_4
X_50694_ _50693_/X _53910_/A sky130_fd_sc_hd__buf_2
X_55221_ _55142_/A _55221_/B _55221_/Y sky130_fd_sc_hd__nor2_4
X_67207_ _88377_/Q _67110_/X _67160_/X _67206_/X _67207_/X sky130_fd_sc_hd__a211o_4
X_86041_ _85529_/CLK _51279_/Y _64820_/B sky130_fd_sc_hd__dfxtp_4
X_52433_ _52429_/Y _52430_/X _52432_/Y _52433_/Y sky130_fd_sc_hd__a21boi_4
X_64419_ _63586_/A _64419_/B _64419_/Y sky130_fd_sc_hd__nor2_4
X_83253_ _85317_/CLK _83253_/D _83253_/Q sky130_fd_sc_hd__dfxtp_4
X_80465_ _80472_/A _80472_/B _80478_/B sky130_fd_sc_hd__xnor2_4
X_68187_ _64636_/A _68376_/A sky130_fd_sc_hd__buf_2
X_65399_ _65198_/A _65399_/X sky130_fd_sc_hd__buf_2
X_82204_ _82961_/CLK _82204_/D _82204_/Q sky130_fd_sc_hd__dfxtp_4
X_55152_ _55152_/A _55152_/X sky130_fd_sc_hd__buf_2
X_67138_ _67135_/X _67137_/X _67113_/X _67138_/Y sky130_fd_sc_hd__a21oi_4
X_52364_ _52262_/A _52364_/X sky130_fd_sc_hd__buf_2
X_83184_ _83184_/CLK _72701_/X _83184_/Q sky130_fd_sc_hd__dfxtp_4
X_80396_ _80393_/X _80395_/Y _82251_/D sky130_fd_sc_hd__xnor2_4
X_54103_ _85503_/Q _53431_/X _54102_/Y _54103_/Y sky130_fd_sc_hd__o21ai_4
X_51315_ _51312_/Y _51313_/X _51314_/X _51315_/Y sky130_fd_sc_hd__a21oi_4
X_82135_ _82009_/CLK _82135_/D _82091_/D sky130_fd_sc_hd__dfxtp_4
X_55083_ _55083_/A _55104_/B _55083_/C _55083_/D _55083_/X sky130_fd_sc_hd__and4_4
X_59960_ _62515_/A _59913_/A _62621_/D _59962_/A sky130_fd_sc_hd__nand3_4
X_67069_ _66972_/X _87614_/Q _67069_/X sky130_fd_sc_hd__and2_4
X_52295_ _52295_/A _52295_/B _52295_/X sky130_fd_sc_hd__and2_4
X_87992_ _88002_/CLK _42185_/X _87992_/Q sky130_fd_sc_hd__dfxtp_4
X_54034_ _54034_/A _54320_/A sky130_fd_sc_hd__buf_2
X_58911_ _58828_/X _58909_/Y _58910_/Y _58874_/X _58832_/X _58911_/X
+ sky130_fd_sc_hd__o32a_4
X_51246_ _51282_/A _51278_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_17_0_CLK clkbuf_7_8_0_CLK/X clkbuf_9_35_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_70080_ _82535_/D _70067_/X _70079_/Y _83855_/D sky130_fd_sc_hd__a21bo_4
X_86943_ _83987_/CLK _86943_/D _86943_/Q sky130_fd_sc_hd__dfxtp_4
X_82066_ _86807_/CLK _82066_/D _82066_/Q sky130_fd_sc_hd__dfxtp_4
X_59891_ _59602_/C _60171_/B _60171_/A _61066_/B sky130_fd_sc_hd__nand3_4
X_81017_ _84150_/CLK _84225_/Q _81017_/Q sky130_fd_sc_hd__dfxtp_4
X_58842_ _84796_/Q _58725_/X _58833_/X _58841_/X _84796_/D sky130_fd_sc_hd__a2bb2oi_4
X_51177_ _51177_/A _51192_/B _51192_/C _52867_/D _51177_/X sky130_fd_sc_hd__and4_4
X_86874_ _86873_/CLK _45484_/Y _63066_/B sky130_fd_sc_hd__dfxtp_4
X_50128_ _50120_/A _52338_/B _50128_/Y sky130_fd_sc_hd__nand2_4
X_85825_ _86145_/CLK _85825_/D _85825_/Q sky130_fd_sc_hd__dfxtp_4
X_58773_ _58667_/X _86097_/Q _58772_/X _58773_/Y sky130_fd_sc_hd__o21ai_4
X_55985_ _56019_/B _55966_/X _55975_/X _74286_/C _55985_/Y sky130_fd_sc_hd__nand4_4
X_57724_ _57705_/X _85504_/Q _44031_/X _57724_/X sky130_fd_sc_hd__o21a_4
X_42950_ _42962_/A _42950_/X sky130_fd_sc_hd__buf_2
X_50059_ _48894_/A _48859_/B _50059_/C _50059_/X sky130_fd_sc_hd__and3_4
X_54936_ _54882_/A _54936_/X sky130_fd_sc_hd__buf_2
X_73770_ _88106_/Q _73649_/X _73770_/Y sky130_fd_sc_hd__nor2_4
X_85756_ _85757_/CLK _52780_/Y _85756_/Q sky130_fd_sc_hd__dfxtp_4
X_82968_ _82774_/CLK _82968_/D _82968_/Q sky130_fd_sc_hd__dfxtp_4
X_70982_ _70981_/X _70983_/A sky130_fd_sc_hd__buf_2
Xclkbuf_3_3_1_CLK clkbuf_3_3_0_CLK/X clkbuf_4_7_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_41901_ _43175_/B _46616_/A sky130_fd_sc_hd__buf_2
X_72721_ _73257_/A _72721_/X sky130_fd_sc_hd__buf_2
X_84707_ _84355_/CLK _84707_/D _80559_/A sky130_fd_sc_hd__dfxtp_4
X_57655_ _57655_/A _57655_/Y sky130_fd_sc_hd__inv_2
X_81919_ _82008_/CLK _77692_/Y _77157_/B sky130_fd_sc_hd__dfxtp_4
X_42881_ _42835_/X _42881_/X sky130_fd_sc_hd__buf_2
X_54867_ _54885_/A _54867_/B _54867_/Y sky130_fd_sc_hd__nand2_4
X_85687_ _84787_/CLK _85687_/D _85687_/Q sky130_fd_sc_hd__dfxtp_4
X_82899_ _82899_/CLK _78202_/B _82899_/Q sky130_fd_sc_hd__dfxtp_4
X_44620_ _40982_/A _44618_/X _87030_/Q _44619_/X _87030_/D sky130_fd_sc_hd__a2bb2o_4
X_56606_ _72652_/C _56556_/A _56607_/A sky130_fd_sc_hd__xor2_4
X_75440_ _80794_/Q _75440_/B _75440_/X sky130_fd_sc_hd__xor2_4
X_41832_ _40469_/X _41813_/X _88131_/Q _41814_/X _41832_/X sky130_fd_sc_hd__a2bb2o_4
X_87426_ _86784_/CLK _43429_/X _87426_/Q sky130_fd_sc_hd__dfxtp_4
X_53818_ _53956_/A _53819_/A sky130_fd_sc_hd__buf_2
X_72652_ _72656_/A _72656_/B _72652_/C _72652_/Y sky130_fd_sc_hd__nand3_4
X_84638_ _84620_/CLK _60307_/X _79764_/A sky130_fd_sc_hd__dfxtp_4
X_57586_ _50460_/A _71964_/A sky130_fd_sc_hd__buf_2
X_54798_ _54798_/A _54816_/B _54798_/C _53107_/D _54798_/X sky130_fd_sc_hd__and4_4
X_71603_ _71603_/A _71603_/Y sky130_fd_sc_hd__inv_2
X_59325_ _59325_/A _59325_/X sky130_fd_sc_hd__buf_2
X_44551_ _44551_/A _87058_/D sky130_fd_sc_hd__inv_2
X_56537_ _56153_/X _56528_/X _56536_/Y _85158_/D sky130_fd_sc_hd__o21ai_4
X_87357_ _86814_/CLK _43568_/Y _87357_/Q sky130_fd_sc_hd__dfxtp_4
X_75371_ _75371_/A _75370_/X _80758_/D sky130_fd_sc_hd__xor2_4
X_41763_ _41753_/X _41754_/X _41762_/X _67932_/B _41736_/X _41764_/A
+ sky130_fd_sc_hd__o32ai_4
X_53749_ _53746_/Y _53747_/X _53748_/X _53749_/Y sky130_fd_sc_hd__a21oi_4
X_72583_ _72525_/A _72597_/B _72583_/C _72583_/Y sky130_fd_sc_hd__nand3_4
X_84569_ _82436_/CLK _84569_/D _78064_/A sky130_fd_sc_hd__dfxtp_4
X_77110_ _77110_/A _77110_/B _82346_/D sky130_fd_sc_hd__xor2_4
X_43502_ _41749_/X _43498_/X _87388_/Q _43499_/X _43502_/X sky130_fd_sc_hd__a2bb2o_4
X_86308_ _86627_/CLK _86308_/D _58116_/B sky130_fd_sc_hd__dfxtp_4
X_74322_ _70306_/C _74314_/X _74321_/Y _83099_/D sky130_fd_sc_hd__a21bo_4
X_40714_ _40714_/A _40623_/X _40714_/X sky130_fd_sc_hd__or2_4
X_47270_ _86652_/Q _47240_/X _47269_/Y _47270_/Y sky130_fd_sc_hd__o21ai_4
X_59256_ _59256_/A _59256_/B _59256_/Y sky130_fd_sc_hd__nor2_4
X_71534_ _71585_/A _71622_/D sky130_fd_sc_hd__buf_2
X_78090_ _78087_/Y _78090_/B _78090_/Y sky130_fd_sc_hd__nor2_4
X_44482_ _44548_/A _44482_/X sky130_fd_sc_hd__buf_2
X_56468_ _56538_/A _56468_/X sky130_fd_sc_hd__buf_2
X_41694_ _41693_/X _41682_/X _67608_/B _41684_/X _41694_/X sky130_fd_sc_hd__a2bb2o_4
X_87288_ _87288_/CLK _87288_/D _87288_/Q sky130_fd_sc_hd__dfxtp_4
X_46221_ _46143_/B _46101_/A _46162_/C _46217_/B _46221_/Y sky130_fd_sc_hd__nand4_4
XPHY_330 sky130_fd_sc_hd__decap_3
X_58207_ _58207_/A _58238_/B _58207_/Y sky130_fd_sc_hd__nor2_4
X_77041_ _77041_/A _77041_/B _77041_/C _77041_/Y sky130_fd_sc_hd__nand3_4
X_43433_ _41560_/X _43431_/X _87424_/Q _43432_/X _87424_/D sky130_fd_sc_hd__a2bb2o_4
X_55419_ _55423_/B _55421_/B sky130_fd_sc_hd__inv_2
X_74253_ _73972_/X _86563_/Q _74253_/X sky130_fd_sc_hd__and2_4
X_86239_ _86436_/CLK _50235_/Y _86239_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_341 sky130_fd_sc_hd__decap_3
X_40645_ _40585_/X _82871_/Q _40644_/X _40645_/Y sky130_fd_sc_hd__o21ai_4
X_71465_ _71429_/A _71476_/D sky130_fd_sc_hd__buf_2
X_59187_ _59184_/Y _59186_/Y _59165_/X _59187_/X sky130_fd_sc_hd__a21o_4
XPHY_352 sky130_fd_sc_hd__decap_3
X_56399_ _56397_/X _56399_/B _85209_/Q _56399_/Y sky130_fd_sc_hd__nand3_4
XPHY_363 sky130_fd_sc_hd__decap_3
XPHY_374 sky130_fd_sc_hd__decap_3
X_73204_ _87054_/Q _73129_/X _73203_/X _73220_/C sky130_fd_sc_hd__o21ai_4
X_70416_ HASH_ADDR[1] _70416_/Y sky130_fd_sc_hd__inv_2
X_46152_ _46166_/C _46170_/C sky130_fd_sc_hd__buf_2
X_58138_ _58100_/X _85474_/Q _58062_/X _58138_/X sky130_fd_sc_hd__o21a_4
XPHY_385 sky130_fd_sc_hd__decap_3
X_43364_ _43364_/A _87458_/D sky130_fd_sc_hd__inv_2
X_74184_ _74184_/A _73152_/X _74184_/Y sky130_fd_sc_hd__nor2_4
X_40576_ _47825_/A _49048_/A sky130_fd_sc_hd__buf_2
XPHY_396 sky130_fd_sc_hd__decap_3
X_71396_ _71395_/Y _71396_/Y sky130_fd_sc_hd__inv_2
X_45103_ _56501_/C _45060_/X _45040_/X _45103_/X sky130_fd_sc_hd__o21a_4
X_42315_ _42307_/X _42297_/X _41621_/X _87925_/Q _42298_/X _42316_/A
+ sky130_fd_sc_hd__o32ai_4
X_73135_ _73260_/A _86483_/Q _73135_/X sky130_fd_sc_hd__and2_4
X_46083_ _41625_/Y _43586_/X _86775_/Q _43593_/X _86775_/D sky130_fd_sc_hd__a2bb2o_4
X_58069_ _84928_/Q _58025_/X _58061_/X _58068_/X _84928_/D sky130_fd_sc_hd__a2bb2oi_4
X_70347_ _70337_/X _74760_/A _70346_/X _83788_/D sky130_fd_sc_hd__a21o_4
X_43295_ _40362_/X _43296_/A sky130_fd_sc_hd__buf_2
X_78992_ _78987_/Y _78979_/B _78991_/Y _78993_/B sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_361_0_CLK clkbuf_9_180_0_CLK/X _86312_/CLK sky130_fd_sc_hd__clkbuf_1
X_60100_ _59913_/A _59881_/X _59884_/X _59973_/A _60100_/Y sky130_fd_sc_hd__nand4_4
X_49911_ _49909_/Y _49897_/X _49910_/X _49911_/Y sky130_fd_sc_hd__a21oi_4
X_45034_ _45031_/X _45033_/Y _44973_/X _45034_/Y sky130_fd_sc_hd__a21oi_4
X_42246_ _42245_/Y _87962_/D sky130_fd_sc_hd__inv_2
X_73066_ _72959_/X _85590_/Q _72839_/X _73065_/X _73066_/X sky130_fd_sc_hd__a211o_4
X_77943_ _82250_/Q _81962_/Q _77944_/B sky130_fd_sc_hd__xor2_4
X_61080_ _61205_/B _61079_/Y _59662_/C _61070_/C _61081_/A sky130_fd_sc_hd__and4_4
Xclkbuf_10_991_0_CLK clkbuf_9_495_0_CLK/X _85562_/CLK sky130_fd_sc_hd__clkbuf_1
X_70278_ _70269_/X _74775_/B _70277_/X _70278_/X sky130_fd_sc_hd__a21o_4
X_60031_ _59710_/Y _60620_/B _60620_/C _60031_/X sky130_fd_sc_hd__and3_4
X_72017_ _72017_/A _72017_/X sky130_fd_sc_hd__buf_2
X_49842_ _86313_/Q _49825_/X _49841_/Y _49842_/Y sky130_fd_sc_hd__o21ai_4
X_42177_ _42173_/X _42169_/X _41234_/X _87996_/Q _42170_/X _42178_/A
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_9_482_0_CLK clkbuf_9_483_0_CLK/A clkbuf_9_482_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_77874_ _77861_/A _77869_/A _77874_/X sky130_fd_sc_hd__and2_4
X_79613_ _79611_/Y _79612_/Y _79613_/X sky130_fd_sc_hd__xor2_4
X_41128_ _81726_/Q _41102_/B _41128_/X sky130_fd_sc_hd__or2_4
X_76825_ _76825_/A _76824_/Y _76826_/B sky130_fd_sc_hd__xor2_4
Xclkbuf_10_376_0_CLK clkbuf_9_188_0_CLK/X _86686_/CLK sky130_fd_sc_hd__clkbuf_1
X_49773_ _49771_/Y _49759_/X _49772_/X _49773_/Y sky130_fd_sc_hd__a21oi_4
X_46985_ _46959_/A _52787_/B _46985_/Y sky130_fd_sc_hd__nand2_4
X_48724_ _48722_/Y _48156_/X _48723_/X _86495_/D sky130_fd_sc_hd__a21oi_4
X_79544_ _79544_/A _79540_/C _79545_/B sky130_fd_sc_hd__nand2_4
X_45936_ _45919_/Y _45928_/X _45935_/X _86842_/D sky130_fd_sc_hd__a21oi_4
X_41059_ _41058_/Y _41059_/X sky130_fd_sc_hd__buf_2
X_64770_ _64615_/X _85563_/Q _64642_/X _64769_/X _64770_/X sky130_fd_sc_hd__a211o_4
X_76756_ _76768_/A _76755_/Y _76763_/A sky130_fd_sc_hd__xor2_4
X_61982_ _63562_/A _59841_/X _61528_/A _61981_/X _61982_/X sky130_fd_sc_hd__a2bb2o_4
X_73968_ _88354_/Q _73777_/X _73898_/X _73968_/X sky130_fd_sc_hd__o21a_4
X_63721_ _61714_/A _60870_/X _63721_/C _61012_/A _63721_/Y sky130_fd_sc_hd__nand4_4
X_75707_ _81121_/Q _75707_/B _75707_/Y sky130_fd_sc_hd__xnor2_4
Xclkbuf_9_497_0_CLK clkbuf_9_497_0_CLK/A clkbuf_9_497_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_48655_ _48652_/X _48110_/A _48654_/Y _48656_/A sky130_fd_sc_hd__o21ai_4
X_60933_ _60359_/A _60933_/X sky130_fd_sc_hd__buf_2
X_72919_ _73050_/A _72918_/Y _72919_/Y sky130_fd_sc_hd__nor2_4
X_79475_ _84814_/Q _84134_/Q _79475_/X sky130_fd_sc_hd__xor2_4
X_45867_ _85090_/Q _57084_/B sky130_fd_sc_hd__inv_2
X_76687_ _76680_/Y _76685_/Y _76686_/Y _76687_/Y sky130_fd_sc_hd__a21oi_4
X_73899_ _68735_/B _73777_/X _73898_/X _73899_/X sky130_fd_sc_hd__o21a_4
X_47606_ _55005_/D _53144_/D sky130_fd_sc_hd__buf_2
X_66440_ _66391_/A _66476_/B sky130_fd_sc_hd__buf_2
X_78426_ _78413_/Y _78426_/B _78426_/C _78426_/Y sky130_fd_sc_hd__nand3_4
X_44818_ _45964_/A _44818_/X sky130_fd_sc_hd__buf_2
X_63652_ _63648_/Y _63649_/X _63651_/X _58344_/A _63363_/X _63652_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75638_ _75638_/A _75637_/Y _75659_/A sky130_fd_sc_hd__xor2_4
X_48586_ _81773_/Q _48586_/Y sky130_fd_sc_hd__inv_2
X_60864_ _60863_/X _60864_/X sky130_fd_sc_hd__buf_2
X_45798_ _45734_/A _45798_/X sky130_fd_sc_hd__buf_2
X_62603_ _62596_/X _62600_/Y _62602_/X _84869_/Q _62572_/X _62603_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47537_ _47553_/A _53105_/B _47537_/Y sky130_fd_sc_hd__nand2_4
X_66371_ _65938_/X _66367_/B _65940_/X _66371_/Y sky130_fd_sc_hd__nand3_4
X_78357_ _78358_/A _78358_/B _78360_/A sky130_fd_sc_hd__or2_4
X_44749_ _44740_/X _44741_/X _40762_/X _86976_/Q _44742_/X _44749_/Y
+ sky130_fd_sc_hd__o32ai_4
X_63583_ _58383_/A _63558_/X _61551_/A _63559_/X _63583_/X sky130_fd_sc_hd__a2bb2o_4
X_75569_ _75574_/A _80818_/Q _75887_/A sky130_fd_sc_hd__xnor2_4
Xclkbuf_9_420_0_CLK clkbuf_8_210_0_CLK/X clkbuf_9_420_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_60795_ _60660_/X _60725_/B _60778_/Y _60795_/X sky130_fd_sc_hd__o21a_4
X_68110_ _68089_/A _68110_/X sky130_fd_sc_hd__buf_2
X_65322_ _65312_/Y _65321_/Y _63231_/X _65322_/Y sky130_fd_sc_hd__a21oi_4
X_77308_ _77308_/A _77308_/Y sky130_fd_sc_hd__inv_2
X_62534_ _62534_/A _62534_/X sky130_fd_sc_hd__buf_2
X_69090_ _88085_/Q _68640_/X _69088_/X _69089_/Y _69090_/X sky130_fd_sc_hd__a211o_4
X_47468_ _47468_/A _47469_/A sky130_fd_sc_hd__inv_2
Xclkbuf_10_314_0_CLK clkbuf_9_157_0_CLK/X _82251_/CLK sky130_fd_sc_hd__clkbuf_1
X_78288_ _78296_/A _78296_/B _78292_/A sky130_fd_sc_hd__xnor2_4
X_49207_ _49232_/A _51235_/B _49207_/Y sky130_fd_sc_hd__nand2_4
X_68041_ _68637_/A _68437_/A sky130_fd_sc_hd__buf_2
X_46419_ _46419_/A _52494_/B sky130_fd_sc_hd__inv_2
X_65253_ _65206_/A _65253_/B _65253_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_944_0_CLK clkbuf_9_472_0_CLK/X _88324_/CLK sky130_fd_sc_hd__clkbuf_1
X_77239_ _77239_/A _77239_/B _77239_/C _77245_/C sky130_fd_sc_hd__nand3_4
X_62465_ _61538_/B _62462_/X _62436_/X _62407_/X _62464_/X _62465_/X
+ sky130_fd_sc_hd__a41o_4
X_47399_ _47399_/A _53023_/D sky130_fd_sc_hd__buf_2
X_64204_ _64440_/A _64267_/A sky130_fd_sc_hd__buf_2
X_49138_ _48985_/A _49138_/X sky130_fd_sc_hd__buf_2
X_61416_ _61411_/X _61394_/X _61415_/Y _61416_/Y sky130_fd_sc_hd__a21oi_4
X_80250_ _80239_/Y _80242_/Y _80250_/X sky130_fd_sc_hd__or2_4
X_65184_ _65184_/A _85835_/Q _65184_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_435_0_CLK clkbuf_9_435_0_CLK/A clkbuf_9_435_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_62396_ _62395_/X _62396_/X sky130_fd_sc_hd__buf_2
X_64135_ _61640_/A _60967_/X _64134_/Y _64135_/X sky130_fd_sc_hd__a21bo_4
X_49069_ _49069_/A _52355_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_329_0_CLK clkbuf_9_164_0_CLK/X _86008_/CLK sky130_fd_sc_hd__clkbuf_1
X_61347_ _59961_/A _61348_/A sky130_fd_sc_hd__buf_2
X_80181_ _80178_/Y _80162_/B _80180_/X _80189_/A sky130_fd_sc_hd__o21ai_4
X_69992_ _59831_/X _69992_/X sky130_fd_sc_hd__buf_2
X_51100_ _51098_/Y _51093_/X _51099_/X _86074_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_959_0_CLK clkbuf_9_479_0_CLK/X _86213_/CLK sky130_fd_sc_hd__clkbuf_1
X_52080_ _52078_/Y _52066_/X _52079_/Y _52080_/Y sky130_fd_sc_hd__a21boi_4
X_68943_ _69357_/A _69011_/A sky130_fd_sc_hd__buf_2
X_64066_ _63610_/B _64095_/B _64095_/C _64095_/D _64066_/Y sky130_fd_sc_hd__nand4_4
X_61278_ _61278_/A _61278_/B _61281_/C _61312_/A sky130_fd_sc_hd__and3_4
X_51031_ _51022_/A _51031_/B _51031_/Y sky130_fd_sc_hd__nand2_4
X_63017_ _60476_/A _63017_/B _63030_/C _60541_/C _63017_/X sky130_fd_sc_hd__and4_4
X_60229_ _60224_/Y _60331_/B _60331_/D _60229_/Y sky130_fd_sc_hd__nand3_4
X_83940_ _83940_/CLK _83940_/D _81404_/D sky130_fd_sc_hd__dfxtp_4
X_68874_ _68869_/X _68873_/X _68806_/X _68874_/X sky130_fd_sc_hd__a21o_4
X_67825_ _67466_/X _67825_/X sky130_fd_sc_hd__buf_2
X_83871_ _82553_/CLK _70022_/X _83871_/Q sky130_fd_sc_hd__dfxtp_4
X_85610_ _84970_/CLK _85610_/D _85610_/Q sky130_fd_sc_hd__dfxtp_4
X_82822_ _82822_/CLK _82822_/D _82822_/Q sky130_fd_sc_hd__dfxtp_4
X_55770_ _83017_/Q _55157_/X _55172_/A _55769_/X _55771_/B sky130_fd_sc_hd__a211o_4
X_67756_ _67658_/X _67756_/B _67756_/X sky130_fd_sc_hd__and2_4
X_86590_ _86558_/CLK _86590_/D _73638_/B sky130_fd_sc_hd__dfxtp_4
X_52982_ _52997_/A _52982_/B _52997_/C _52982_/D _52982_/X sky130_fd_sc_hd__and4_4
X_64968_ _64967_/X _65196_/A sky130_fd_sc_hd__buf_2
X_54721_ _54699_/X _54734_/B _54721_/C _47407_/A _54721_/X sky130_fd_sc_hd__and4_4
X_66707_ _66702_/X _66705_/X _66706_/X _66707_/Y sky130_fd_sc_hd__a21oi_4
X_85541_ _86149_/CLK _85541_/D _85541_/Q sky130_fd_sc_hd__dfxtp_4
X_51933_ _73583_/B _51929_/X _51932_/Y _51933_/Y sky130_fd_sc_hd__o21ai_4
X_63919_ _60879_/B _63951_/C sky130_fd_sc_hd__buf_2
X_82753_ _82746_/CLK _66364_/C _82753_/Q sky130_fd_sc_hd__dfxtp_4
X_67687_ _84059_/Q _67568_/X _67686_/X _67687_/X sky130_fd_sc_hd__a21bo_4
X_64899_ _65319_/A _86422_/Q _64899_/X sky130_fd_sc_hd__and2_4
X_81704_ _81703_/CLK _81704_/D _81704_/Q sky130_fd_sc_hd__dfxtp_4
X_57440_ _57440_/A _57440_/X sky130_fd_sc_hd__buf_2
X_69426_ _88030_/Q _69424_/X _69202_/X _69425_/X _69426_/X sky130_fd_sc_hd__a211o_4
X_88260_ _88263_/CLK _88260_/D _68763_/B sky130_fd_sc_hd__dfxtp_4
X_54652_ _54667_/A _54645_/B _54644_/X _47283_/A _54652_/X sky130_fd_sc_hd__and4_4
X_66638_ _80927_/D _66614_/X _66637_/X _84103_/D sky130_fd_sc_hd__a21bo_4
X_85472_ _85471_/CLK _85472_/D _85472_/Q sky130_fd_sc_hd__dfxtp_4
X_51864_ _51781_/A _51870_/C sky130_fd_sc_hd__buf_2
X_82684_ _82933_/CLK _82684_/D _82684_/Q sky130_fd_sc_hd__dfxtp_4
X_87211_ _86934_/CLK _43894_/X _67527_/B sky130_fd_sc_hd__dfxtp_4
X_53603_ _53696_/A _53603_/X sky130_fd_sc_hd__buf_2
X_84423_ _84424_/CLK _62255_/Y _62254_/C sky130_fd_sc_hd__dfxtp_4
X_50815_ _86127_/Q _50804_/X _50814_/Y _50815_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_5_14_0_CLK clkbuf_4_7_1_CLK/X clkbuf_6_29_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_57371_ _44308_/X _57440_/A sky130_fd_sc_hd__buf_2
X_81635_ _81794_/CLK _81667_/Q _81635_/Q sky130_fd_sc_hd__dfxtp_4
X_69357_ _69357_/A _69383_/A sky130_fd_sc_hd__buf_2
X_88191_ _87686_/CLK _41567_/Y _67052_/B sky130_fd_sc_hd__dfxtp_4
X_54583_ _85415_/Q _54567_/X _54582_/Y _54583_/Y sky130_fd_sc_hd__o21ai_4
X_66569_ _44146_/A _68392_/A sky130_fd_sc_hd__buf_2
X_51795_ _51792_/Y _51793_/X _51794_/X _51795_/Y sky130_fd_sc_hd__a21oi_4
X_59110_ _58941_/A _86360_/Q _59110_/Y sky130_fd_sc_hd__nor2_4
X_56322_ _56347_/A _56332_/A sky130_fd_sc_hd__buf_2
X_68308_ _68447_/A _68308_/X sky130_fd_sc_hd__buf_2
X_87142_ _87141_/CLK _44372_/Y _87142_/Q sky130_fd_sc_hd__dfxtp_4
X_53534_ _53532_/Y _53472_/X _53533_/X _53534_/Y sky130_fd_sc_hd__a21oi_4
X_84354_ _84321_/CLK _84354_/D _79436_/A sky130_fd_sc_hd__dfxtp_4
X_50746_ _50740_/A _53959_/B _50746_/Y sky130_fd_sc_hd__nand2_4
X_81566_ _81482_/CLK _81566_/D _81522_/D sky130_fd_sc_hd__dfxtp_4
X_69288_ _69288_/A _69288_/B _69288_/X sky130_fd_sc_hd__and2_4
X_83305_ _83305_/CLK _83305_/D _83305_/Q sky130_fd_sc_hd__dfxtp_4
X_59041_ _84774_/Q _58956_/X _59032_/X _59040_/X _84774_/D sky130_fd_sc_hd__a2bb2oi_4
X_80517_ _80517_/A _63493_/C _80518_/B sky130_fd_sc_hd__xor2_4
X_56253_ _56263_/A _56253_/B _56253_/C _56253_/Y sky130_fd_sc_hd__nand3_4
X_68239_ _68208_/X _68239_/X sky130_fd_sc_hd__buf_2
X_87073_ _87073_/CLK _44509_/Y _87073_/Q sky130_fd_sc_hd__dfxtp_4
X_53465_ _53990_/A _53687_/A sky130_fd_sc_hd__buf_2
X_84285_ _84280_/CLK _84285_/D _63944_/C sky130_fd_sc_hd__dfxtp_4
X_50677_ _50677_/A _50651_/X _50668_/C _50677_/X sky130_fd_sc_hd__and3_4
X_81497_ _81749_/CLK _84065_/Q _81497_/Q sky130_fd_sc_hd__dfxtp_4
X_55204_ _55710_/B _45826_/Y _55204_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_5_29_0_CLK clkbuf_4_14_1_CLK/X clkbuf_6_59_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_86024_ _86121_/CLK _86024_/D _65260_/B sky130_fd_sc_hd__dfxtp_4
X_40430_ _40368_/X _40430_/B _40430_/X sky130_fd_sc_hd__or2_4
X_52416_ _52407_/A _49192_/A _52416_/X sky130_fd_sc_hd__and2_4
X_71250_ _71252_/A _71226_/B _71248_/C _71250_/Y sky130_fd_sc_hd__nand3_4
X_83236_ _83231_/CLK _72548_/Y _79456_/B sky130_fd_sc_hd__dfxtp_4
X_56184_ _74539_/A _56460_/B sky130_fd_sc_hd__buf_2
X_80448_ _80448_/A _80448_/B _80448_/X sky130_fd_sc_hd__and2_4
X_53396_ _85641_/Q _53378_/X _53395_/Y _53396_/Y sky130_fd_sc_hd__o21ai_4
X_70201_ _70195_/X _74789_/C _70200_/X _70201_/X sky130_fd_sc_hd__a21o_4
X_55135_ _55135_/A _57179_/B _55135_/X sky130_fd_sc_hd__and2_4
X_52347_ _52324_/A _52347_/X sky130_fd_sc_hd__buf_2
X_40361_ _40361_/A _42081_/A sky130_fd_sc_hd__inv_2
X_71181_ _71181_/A _71185_/B _71181_/C _74518_/D _71181_/Y sky130_fd_sc_hd__nand4_4
X_83167_ _83167_/CLK _83167_/D _83167_/Q sky130_fd_sc_hd__dfxtp_4
X_80379_ _80379_/A _80379_/B _80380_/B sky130_fd_sc_hd__xor2_4
X_42100_ _42099_/X _42094_/X _41021_/X _88036_/Q _42096_/X _42101_/A
+ sky130_fd_sc_hd__o32ai_4
X_70132_ _83115_/Q _70134_/B sky130_fd_sc_hd__inv_2
X_82118_ _82145_/CLK _77768_/X _82118_/Q sky130_fd_sc_hd__dfxtp_4
X_43080_ _43121_/A _43080_/X sky130_fd_sc_hd__buf_2
X_55066_ _55064_/Y _55050_/X _55065_/X _85325_/D sky130_fd_sc_hd__a21oi_4
X_59943_ _59943_/A _59943_/X sky130_fd_sc_hd__buf_2
X_52278_ _85854_/Q _52269_/X _52277_/Y _52278_/Y sky130_fd_sc_hd__o21ai_4
X_83098_ _83846_/CLK _83098_/D _83098_/Q sky130_fd_sc_hd__dfxtp_4
X_87975_ _87149_/CLK _87975_/D _87975_/Q sky130_fd_sc_hd__dfxtp_4
X_42031_ _42028_/X _42024_/X _40866_/X _73247_/A _42025_/X _42031_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54017_ _54014_/Y _54015_/X _54016_/X _85522_/D sky130_fd_sc_hd__a21oi_4
X_51229_ _51147_/A _51229_/X sky130_fd_sc_hd__buf_2
X_74940_ _74940_/A _74940_/B _74940_/X sky130_fd_sc_hd__xor2_4
X_70063_ _68912_/X _68914_/X _69992_/X _70063_/X sky130_fd_sc_hd__a21o_4
X_86926_ _87652_/CLK _44841_/X _86926_/Q sky130_fd_sc_hd__dfxtp_4
X_82049_ _82575_/CLK _78033_/Y _82017_/D sky130_fd_sc_hd__dfxtp_4
X_59874_ _59727_/X _59745_/X _59651_/C _59859_/Y _59873_/Y _59874_/Y
+ sky130_fd_sc_hd__a41oi_4
X_58825_ _58822_/Y _58824_/Y _58735_/X _58825_/X sky130_fd_sc_hd__a21o_4
X_74871_ _81125_/D _74870_/B _74871_/Y sky130_fd_sc_hd__nand2_4
X_86857_ _80664_/CLK _45751_/Y _63265_/B sky130_fd_sc_hd__dfxtp_4
X_76610_ _76611_/A _76609_/Y _81375_/Q _76613_/A sky130_fd_sc_hd__a21oi_4
X_85808_ _86030_/CLK _85808_/D _65049_/B sky130_fd_sc_hd__dfxtp_4
X_73822_ _73822_/A _74246_/B _73822_/Y sky130_fd_sc_hd__nor2_4
X_46770_ _52663_/B _50971_/B sky130_fd_sc_hd__buf_2
X_58756_ _58641_/A _58756_/X sky130_fd_sc_hd__buf_2
X_77590_ _77590_/A _77590_/B _77591_/A sky130_fd_sc_hd__and2_4
X_43982_ _59538_/C _60665_/C sky130_fd_sc_hd__buf_2
X_55968_ _56198_/C _55690_/A _44052_/X _55967_/X _55968_/X sky130_fd_sc_hd__a211o_4
X_86788_ _86814_/CLK _46060_/X _86788_/Q sky130_fd_sc_hd__dfxtp_4
X_45721_ _85068_/Q _45801_/A _45721_/Y sky130_fd_sc_hd__nor2_4
X_57707_ _46224_/X _85409_/Q _57706_/X _57707_/Y sky130_fd_sc_hd__o21ai_4
X_76541_ _76541_/A _76541_/B _76584_/C sky130_fd_sc_hd__and2_4
X_42933_ _41749_/X _42930_/X _87644_/Q _42931_/X _42933_/X sky130_fd_sc_hd__a2bb2o_4
X_54919_ _54919_/A _54919_/X sky130_fd_sc_hd__buf_2
X_73753_ _43048_/Y _73627_/X _73652_/X _73752_/Y _73753_/X sky130_fd_sc_hd__a211o_4
X_85739_ _85741_/CLK _52873_/Y _85739_/Q sky130_fd_sc_hd__dfxtp_4
X_70965_ _46356_/X _70961_/X _70964_/Y _70965_/Y sky130_fd_sc_hd__o21ai_4
X_58687_ _58687_/A _58687_/B _58687_/Y sky130_fd_sc_hd__nor2_4
X_55899_ _55908_/A _55949_/A sky130_fd_sc_hd__buf_2
X_48440_ _48440_/A _52135_/A sky130_fd_sc_hd__buf_2
X_72704_ _72704_/A _72714_/A sky130_fd_sc_hd__buf_2
X_79260_ _79258_/X _79260_/B _79270_/B sky130_fd_sc_hd__xor2_4
X_45652_ _85137_/Q _45556_/X _45651_/X _45652_/X sky130_fd_sc_hd__o21a_4
X_57638_ _84964_/Q _57635_/X _57637_/Y _57638_/Y sky130_fd_sc_hd__o21ai_4
X_76472_ _81272_/Q _81528_/D _76473_/A sky130_fd_sc_hd__nand2_4
X_42864_ _42847_/X _42849_/X _41565_/X _67047_/B _42858_/X _42865_/A
+ sky130_fd_sc_hd__o32ai_4
X_73684_ _73607_/A _65972_/B _73684_/X sky130_fd_sc_hd__and2_4
X_70896_ _70925_/A _70899_/C sky130_fd_sc_hd__buf_2
X_78211_ _82676_/Q _78211_/B _78211_/X sky130_fd_sc_hd__xor2_4
X_44603_ _44603_/A _44603_/X sky130_fd_sc_hd__buf_2
X_75423_ _81082_/Q _75423_/Y sky130_fd_sc_hd__inv_2
X_87409_ _87922_/CLK _87409_/D _87409_/Q sky130_fd_sc_hd__dfxtp_4
X_41815_ _40408_/X _41813_/X _88139_/Q _41814_/X _88139_/D sky130_fd_sc_hd__a2bb2o_4
X_48371_ _40420_/A _48471_/A sky130_fd_sc_hd__buf_2
X_72635_ _72633_/X _72643_/B _56564_/D _72635_/Y sky130_fd_sc_hd__nand3_4
X_79191_ _79189_/B _79189_/A _79192_/B sky130_fd_sc_hd__nand2_4
X_45583_ _45581_/Y _45516_/X _45548_/X _45582_/Y _45583_/X sky130_fd_sc_hd__a211o_4
X_57569_ _57564_/X _53535_/B _57569_/Y sky130_fd_sc_hd__nand2_4
X_88389_ _88133_/CLK _40454_/Y _88389_/Q sky130_fd_sc_hd__dfxtp_4
X_42795_ _42720_/X _42795_/X sky130_fd_sc_hd__buf_2
X_47322_ _47316_/Y _47317_/X _47321_/X _86647_/D sky130_fd_sc_hd__a21oi_4
X_59308_ _72255_/A _59308_/X sky130_fd_sc_hd__buf_2
X_78142_ _78137_/Y _78129_/X _78141_/Y _78143_/B sky130_fd_sc_hd__a21boi_4
X_44534_ _44529_/X _44530_/X _40798_/A _44531_/Y _44533_/X _87065_/D
+ sky130_fd_sc_hd__o32ai_4
X_75354_ _75354_/A _75353_/Y _75354_/X sky130_fd_sc_hd__and2_4
X_41746_ _41745_/X _41722_/X _67873_/B _41723_/X _88157_/D sky130_fd_sc_hd__a2bb2o_4
X_60580_ _60525_/A _60612_/B sky130_fd_sc_hd__buf_2
X_72566_ _60356_/Y _72522_/Y _72562_/Y _72570_/C _72565_/Y _72566_/Y
+ sky130_fd_sc_hd__a41oi_4
X_74305_ _83106_/Q _74301_/X _74304_/Y _83106_/D sky130_fd_sc_hd__a21bo_4
X_47253_ _47241_/X _52940_/B _47253_/Y sky130_fd_sc_hd__nand2_4
X_59239_ _59238_/X _86350_/Q _59239_/Y sky130_fd_sc_hd__nor2_4
X_71517_ _71521_/A _70717_/A _71517_/Y sky130_fd_sc_hd__nand2_4
X_78073_ _84578_/Q _78073_/B _81882_/D sky130_fd_sc_hd__xor2_4
X_44465_ _40353_/Y _44603_/A sky130_fd_sc_hd__buf_2
X_75285_ _80784_/Q _75284_/X _75285_/X sky130_fd_sc_hd__xor2_4
X_41677_ _41672_/X _41673_/X _41676_/X _88171_/Q _41668_/X _41678_/A
+ sky130_fd_sc_hd__o32ai_4
X_72497_ _46150_/B _83380_/Q _72496_/Y _72497_/X sky130_fd_sc_hd__o21a_4
X_46204_ _58160_/B _46204_/B _46204_/C _46204_/D _46204_/Y sky130_fd_sc_hd__nand4_4
XPHY_160 sky130_fd_sc_hd__decap_3
X_77024_ _77018_/A _82277_/D _77024_/Y sky130_fd_sc_hd__nor2_4
X_43416_ _43416_/A _43416_/Y sky130_fd_sc_hd__inv_2
X_62250_ _61356_/X _62560_/B _62560_/C _62211_/D _62251_/D sky130_fd_sc_hd__nand4_4
X_74236_ _74233_/X _74235_/X _56547_/X _74239_/A sky130_fd_sc_hd__a21o_4
XPHY_171 sky130_fd_sc_hd__decap_3
X_40628_ _40623_/X _40628_/X sky130_fd_sc_hd__buf_2
X_47184_ _47184_/A _47184_/X sky130_fd_sc_hd__buf_2
X_71448_ _70673_/A _71626_/C _71450_/C _71448_/Y sky130_fd_sc_hd__nor3_4
X_44396_ _41485_/X _44394_/X _87130_/Q _44395_/X _87130_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_182 sky130_fd_sc_hd__decap_3
XPHY_193 sky130_fd_sc_hd__decap_3
Xclkbuf_7_112_0_CLK clkbuf_6_56_0_CLK/X clkbuf_8_225_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_61201_ _61194_/X _61198_/X _61135_/X _61188_/Y _61200_/X _61201_/X
+ sky130_fd_sc_hd__o41a_4
X_46135_ _46135_/A _46204_/C _46135_/Y sky130_fd_sc_hd__nand2_4
X_43347_ _43296_/A _43347_/X sky130_fd_sc_hd__buf_2
X_62181_ _62181_/A _62181_/B _78050_/B _62181_/Y sky130_fd_sc_hd__nor3_4
X_74167_ _43096_/Y _56273_/X _73035_/X _74166_/Y _74167_/X sky130_fd_sc_hd__a211o_4
X_40559_ _40380_/X _82881_/Q _40558_/X _40559_/X sky130_fd_sc_hd__o21a_4
X_71379_ _70673_/A _71377_/B _71377_/C _71379_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_10_82_0_CLK clkbuf_9_41_0_CLK/X _86770_/CLK sky130_fd_sc_hd__clkbuf_1
X_61132_ _60946_/X _61138_/B _61132_/C _61132_/Y sky130_fd_sc_hd__nor3_4
X_73118_ _72978_/X _83068_/Q _72992_/X _73117_/X _73118_/X sky130_fd_sc_hd__a211o_4
X_46066_ _41569_/Y _46061_/X _86785_/Q _46062_/X _86785_/D sky130_fd_sc_hd__a2bb2o_4
X_43278_ _43218_/A _43278_/X sky130_fd_sc_hd__buf_2
X_74098_ _43089_/Y _72895_/X _73486_/X _74097_/Y _74098_/X sky130_fd_sc_hd__a211o_4
X_78975_ _78975_/A _78975_/B _78975_/X sky130_fd_sc_hd__xor2_4
X_45017_ _45014_/Y _45016_/Y _44986_/X _45017_/X sky130_fd_sc_hd__a21o_4
X_42229_ _42205_/X _42226_/X _41376_/X _87970_/Q _42228_/X _42230_/A
+ sky130_fd_sc_hd__o32ai_4
X_65940_ _65924_/X _84991_/Q _65865_/X _65939_/X _65940_/X sky130_fd_sc_hd__a211o_4
X_61063_ _60846_/Y _61063_/Y sky130_fd_sc_hd__inv_2
X_73049_ _73039_/Y _73048_/X _73049_/Y sky130_fd_sc_hd__xnor2_4
X_77926_ _82248_/Q _81960_/Q _77927_/B sky130_fd_sc_hd__xnor2_4
Xclkbuf_7_127_0_CLK clkbuf_6_63_0_CLK/X clkbuf_8_255_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_60014_ _60109_/A _60014_/X sky130_fd_sc_hd__buf_2
X_49825_ _49825_/A _49825_/X sky130_fd_sc_hd__buf_2
X_65871_ _84172_/Q _65872_/C sky130_fd_sc_hd__inv_2
X_77857_ _77833_/Y _81934_/D sky130_fd_sc_hd__inv_2
Xclkbuf_10_97_0_CLK clkbuf_9_48_0_CLK/X _82987_/CLK sky130_fd_sc_hd__clkbuf_1
X_67610_ _67607_/X _67609_/X _67423_/X _67610_/Y sky130_fd_sc_hd__a21oi_4
X_64822_ _64819_/X _64821_/X _64807_/X _64822_/X sky130_fd_sc_hd__a21o_4
X_76808_ _76808_/A _76807_/Y _76809_/B sky130_fd_sc_hd__xnor2_4
X_49756_ _49754_/Y _49732_/X _49755_/X _86329_/D sky130_fd_sc_hd__a21oi_4
X_68590_ _88106_/Q _68066_/X _67997_/X _68589_/Y _68590_/X sky130_fd_sc_hd__a211o_4
X_46968_ _54469_/B _52777_/B sky130_fd_sc_hd__buf_2
X_77788_ _81928_/D _77776_/A _77788_/X sky130_fd_sc_hd__and2_4
Xclkbuf_8_243_0_CLK clkbuf_8_243_0_CLK/A clkbuf_9_486_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_48707_ _86498_/Q _48548_/X _48706_/Y _48707_/Y sky130_fd_sc_hd__o21ai_4
X_67541_ _87159_/Q _67467_/X _67516_/X _67540_/X _67541_/X sky130_fd_sc_hd__a211o_4
X_79527_ _79526_/Y _60374_/C _79527_/Y sky130_fd_sc_hd__nand2_4
X_45919_ _44005_/X _44024_/A _45918_/Y _45919_/Y sky130_fd_sc_hd__nand3_4
X_64753_ _64826_/A _64753_/B _64753_/X sky130_fd_sc_hd__and2_4
X_76739_ _76728_/Y _81355_/D sky130_fd_sc_hd__inv_2
X_49687_ _49632_/A _49687_/X sky130_fd_sc_hd__buf_2
X_61965_ _57683_/X _61902_/X _61916_/X _61948_/X _61964_/X _61965_/X
+ sky130_fd_sc_hd__a41o_4
X_46899_ _52739_/B _46899_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_20_0_CLK clkbuf_9_10_0_CLK/X _85257_/CLK sky130_fd_sc_hd__clkbuf_1
X_63704_ _59445_/A _63370_/A _61685_/A _60780_/X _63704_/X sky130_fd_sc_hd__a2bb2o_4
X_48638_ _48638_/A _48639_/A sky130_fd_sc_hd__inv_2
X_60916_ _60915_/X _64189_/C sky130_fd_sc_hd__buf_2
X_67472_ _81500_/D _67449_/X _67471_/X _84068_/D sky130_fd_sc_hd__a21bo_4
X_79458_ _79470_/A _79470_/B _79481_/A sky130_fd_sc_hd__xnor2_4
X_64684_ _64684_/A _64684_/B _64684_/X sky130_fd_sc_hd__and2_4
X_61896_ _61885_/X _61887_/X _61894_/Y _84743_/Q _61895_/X _61896_/Y
+ sky130_fd_sc_hd__o32ai_4
X_69211_ _69208_/X _69210_/X _69171_/X _69211_/Y sky130_fd_sc_hd__a21oi_4
X_66423_ _64897_/X _66423_/B _64900_/X _66423_/Y sky130_fd_sc_hd__nand3_4
X_78409_ _78387_/Y _78384_/Y _78385_/Y _78409_/Y sky130_fd_sc_hd__o21ai_4
X_63635_ _63578_/A _63635_/X sky130_fd_sc_hd__buf_2
X_48569_ _52194_/A _48624_/B _48610_/C _48569_/X sky130_fd_sc_hd__and3_4
X_60847_ _60386_/A _60846_/Y _60848_/A sky130_fd_sc_hd__and2_4
X_79389_ _79375_/Y _79381_/B _79388_/X _79390_/B sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_253_0_CLK clkbuf_9_126_0_CLK/X _82436_/CLK sky130_fd_sc_hd__clkbuf_1
X_50600_ _50599_/X _71994_/B sky130_fd_sc_hd__buf_2
X_81420_ _84064_/CLK _81452_/Q _81420_/Q sky130_fd_sc_hd__dfxtp_4
X_69142_ _68660_/X _69142_/X sky130_fd_sc_hd__buf_2
X_66354_ _66117_/X _84962_/Q _66118_/X _66353_/X _66354_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_883_0_CLK clkbuf_9_441_0_CLK/X _85516_/CLK sky130_fd_sc_hd__clkbuf_1
X_51580_ _51580_/A _51580_/B _51603_/C _53107_/D _51580_/X sky130_fd_sc_hd__and4_4
X_63566_ _63556_/X _63557_/X _63560_/X _63563_/X _63565_/Y _63566_/Y
+ sky130_fd_sc_hd__o41ai_4
X_60778_ _60682_/A _63540_/A _60660_/A _60778_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_35_0_CLK clkbuf_9_17_0_CLK/X _85050_/CLK sky130_fd_sc_hd__clkbuf_1
X_65305_ _65299_/X _65303_/X _65304_/X _65305_/X sky130_fd_sc_hd__a21o_4
X_50531_ _48849_/A _50552_/B _50526_/C _50531_/X sky130_fd_sc_hd__and3_4
X_62517_ _62055_/B _62517_/Y sky130_fd_sc_hd__inv_2
X_81351_ _81351_/CLK _81351_/D _76226_/A sky130_fd_sc_hd__dfxtp_4
X_69073_ _69073_/A _88342_/Q _69073_/X sky130_fd_sc_hd__and2_4
X_66285_ _65934_/X _66285_/B _66285_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_374_0_CLK clkbuf_9_375_0_CLK/A clkbuf_9_374_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_63497_ _63436_/A _63497_/X sky130_fd_sc_hd__buf_2
X_80302_ _80299_/Y _80302_/B _80303_/B sky130_fd_sc_hd__nand2_4
X_68024_ _69797_/A _68024_/X sky130_fd_sc_hd__buf_2
X_53250_ _53247_/Y _53242_/X _53249_/X _85669_/D sky130_fd_sc_hd__a21oi_4
X_65236_ _65159_/A _86025_/Q _65236_/X sky130_fd_sc_hd__and2_4
X_84070_ _81461_/CLK _84070_/D _81502_/D sky130_fd_sc_hd__dfxtp_4
X_50462_ _52166_/A _50492_/B _50462_/C _50462_/X sky130_fd_sc_hd__and3_4
X_62448_ _62448_/A _63557_/B _62491_/C _62451_/C sky130_fd_sc_hd__nand3_4
X_81282_ _81282_/CLK _76970_/X _81250_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_268_0_CLK clkbuf_9_134_0_CLK/X _84823_/CLK sky130_fd_sc_hd__clkbuf_1
X_52201_ _52210_/A _48816_/B _52201_/Y sky130_fd_sc_hd__nand2_4
X_83021_ _85221_/CLK _83021_/D _45215_/A sky130_fd_sc_hd__dfxtp_4
X_80233_ _80233_/A _80232_/X _80233_/Y sky130_fd_sc_hd__xnor2_4
Xclkbuf_10_898_0_CLK clkbuf_9_449_0_CLK/X _86998_/CLK sky130_fd_sc_hd__clkbuf_1
X_53181_ _53181_/A _53181_/B _53169_/X _53181_/D _53181_/X sky130_fd_sc_hd__and4_4
X_65167_ _64915_/X _65154_/Y _65166_/Y _65167_/Y sky130_fd_sc_hd__o21ai_4
X_50393_ _50398_/A _48358_/X _50393_/Y sky130_fd_sc_hd__nand2_4
X_62379_ _62337_/A _61909_/X _62364_/X _62280_/D _62379_/X sky130_fd_sc_hd__and4_4
X_52132_ _52127_/X _48435_/B _52132_/Y sky130_fd_sc_hd__nand2_4
X_64118_ _61630_/A _64118_/B _64155_/C _64142_/D _64118_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_9_389_0_CLK clkbuf_9_389_0_CLK/A clkbuf_9_389_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_80164_ _80154_/A _80153_/X _80163_/Y _80164_/Y sky130_fd_sc_hd__a21boi_4
X_65098_ _65095_/X _65097_/X _64851_/X _65102_/A sky130_fd_sc_hd__a21o_4
X_69975_ _69557_/X _69559_/X _69939_/X _69975_/Y sky130_fd_sc_hd__a21oi_4
X_56940_ _45886_/X _45890_/X _56935_/X _56939_/X _44184_/A _56940_/Y
+ sky130_fd_sc_hd__a41oi_4
X_52063_ _52061_/Y _52049_/X _52062_/X _85896_/D sky130_fd_sc_hd__a21oi_4
X_68926_ _68923_/X _68925_/X _68878_/X _68926_/Y sky130_fd_sc_hd__a21oi_4
X_64049_ _60864_/X _64095_/D sky130_fd_sc_hd__buf_2
X_87760_ _87260_/CLK _42706_/X _87760_/Q sky130_fd_sc_hd__dfxtp_4
X_84972_ _83544_/CLK _84972_/D _84972_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_821_0_CLK clkbuf_9_410_0_CLK/X _82933_/CLK sky130_fd_sc_hd__clkbuf_1
X_80095_ _80071_/A _80070_/Y _80080_/Y _80083_/Y _80095_/X sky130_fd_sc_hd__o22a_4
X_51014_ _51018_/A _51029_/B _51029_/C _52704_/D _51014_/X sky130_fd_sc_hd__and4_4
X_86711_ _86711_/CLK _46718_/Y _58688_/A sky130_fd_sc_hd__dfxtp_4
X_83923_ _81507_/CLK _83923_/D _83923_/Q sky130_fd_sc_hd__dfxtp_4
X_56871_ _56869_/Y _55675_/X _56870_/Y _56871_/Y sky130_fd_sc_hd__o21ai_4
X_68857_ _83958_/Q _68838_/X _68856_/X _68857_/X sky130_fd_sc_hd__a21bo_4
X_87691_ _87950_/CLK _42841_/X _87691_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_312_0_CLK clkbuf_9_313_0_CLK/A clkbuf_9_312_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_58610_ _58610_/A _58610_/X sky130_fd_sc_hd__buf_2
X_55822_ _85263_/Q _55492_/X _44047_/X _55821_/X _55822_/X sky130_fd_sc_hd__a211o_4
X_67808_ _67901_/A _67808_/B _67808_/X sky130_fd_sc_hd__and2_4
X_86642_ _86640_/CLK _86642_/D _86642_/Q sky130_fd_sc_hd__dfxtp_4
X_59590_ _61948_/A _59591_/A sky130_fd_sc_hd__buf_2
X_83854_ _82536_/CLK _83854_/D _83854_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_206_0_CLK clkbuf_9_103_0_CLK/X _80697_/CLK sky130_fd_sc_hd__clkbuf_1
X_68788_ _68777_/Y _68358_/X _68649_/X _68787_/Y _68788_/X sky130_fd_sc_hd__a211o_4
X_58541_ _58541_/A _58557_/B _58541_/Y sky130_fd_sc_hd__nand2_4
X_82805_ _82529_/CLK _82837_/Q _82805_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_836_0_CLK clkbuf_9_418_0_CLK/X _85346_/CLK sky130_fd_sc_hd__clkbuf_1
X_67739_ _66554_/X _67739_/X sky130_fd_sc_hd__buf_2
X_55753_ _55192_/A _56145_/C _55753_/X sky130_fd_sc_hd__and2_4
X_86573_ _86530_/CLK _86573_/D _66198_/B sky130_fd_sc_hd__dfxtp_4
X_52965_ _52979_/A _52965_/B _52965_/Y sky130_fd_sc_hd__nand2_4
X_83785_ _85953_/CLK _70372_/Y _83785_/Q sky130_fd_sc_hd__dfxtp_4
X_80997_ _82610_/CLK _65348_/C _80997_/Q sky130_fd_sc_hd__dfxtp_4
X_88312_ _88326_/CLK _40911_/Y _69923_/B sky130_fd_sc_hd__dfxtp_4
X_54704_ _54594_/X _54718_/A sky130_fd_sc_hd__buf_2
X_85524_ _85815_/CLK _54008_/Y _85524_/Q sky130_fd_sc_hd__dfxtp_4
X_51916_ _51902_/A _46912_/X _51916_/Y sky130_fd_sc_hd__nand2_4
X_70750_ _53122_/B _70738_/X _70749_/Y _70750_/Y sky130_fd_sc_hd__o21ai_4
X_58472_ _83416_/Q _58472_/Y sky130_fd_sc_hd__inv_2
X_82736_ _82147_/CLK _84120_/Q _78939_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_327_0_CLK clkbuf_9_326_0_CLK/A clkbuf_9_327_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_55684_ _55683_/Y _55443_/Y _46234_/Y _55684_/X sky130_fd_sc_hd__o21a_4
X_52896_ _52890_/Y _52892_/X _52895_/X _52896_/Y sky130_fd_sc_hd__a21oi_4
X_57423_ _57408_/X _57420_/X _57422_/Y _57423_/Y sky130_fd_sc_hd__o21ai_4
X_69409_ _69302_/A _69409_/B _69409_/X sky130_fd_sc_hd__and2_4
X_88243_ _87416_/CLK _88243_/D _67338_/B sky130_fd_sc_hd__dfxtp_4
X_54635_ _54633_/Y _54611_/X _54634_/X _85406_/D sky130_fd_sc_hd__a21oi_4
X_85455_ _85778_/CLK _54368_/Y _85455_/Q sky130_fd_sc_hd__dfxtp_4
X_51847_ _53269_/A _51853_/A sky130_fd_sc_hd__buf_2
X_70681_ _71883_/A _70682_/A sky130_fd_sc_hd__buf_2
X_82667_ _82879_/CLK _82667_/D _82667_/Q sky130_fd_sc_hd__dfxtp_4
X_41600_ _41577_/X _81158_/Q _41599_/X _41600_/Y sky130_fd_sc_hd__o21ai_4
X_72420_ _72339_/X _85320_/Q _72386_/X _72420_/X sky130_fd_sc_hd__o21a_4
X_84406_ _84420_/CLK _84406_/D _62498_/C sky130_fd_sc_hd__dfxtp_4
X_57354_ _57261_/X _57352_/X _57353_/Y _57354_/Y sky130_fd_sc_hd__a21oi_4
X_81618_ _81631_/CLK _81618_/D _81618_/Q sky130_fd_sc_hd__dfxtp_4
X_88174_ _83987_/CLK _88174_/D _67468_/B sky130_fd_sc_hd__dfxtp_4
X_42580_ _42580_/A _42580_/X sky130_fd_sc_hd__buf_2
X_54566_ _54562_/Y _54558_/X _54565_/X _54566_/Y sky130_fd_sc_hd__a21oi_4
X_85386_ _85484_/CLK _54744_/Y _85386_/Q sky130_fd_sc_hd__dfxtp_4
X_51778_ _51775_/Y _51767_/X _51777_/X _85948_/D sky130_fd_sc_hd__a21oi_4
X_82598_ _82879_/CLK _78845_/B _82598_/Q sky130_fd_sc_hd__dfxtp_4
X_56305_ _56360_/A _56305_/X sky130_fd_sc_hd__buf_2
X_41531_ _41457_/A _41531_/X sky130_fd_sc_hd__buf_2
X_87125_ _88201_/CLK _44403_/X _87125_/Q sky130_fd_sc_hd__dfxtp_4
X_53517_ _53515_/Y _53498_/X _53516_/Y _53517_/Y sky130_fd_sc_hd__a21boi_4
X_72351_ _72305_/X _85358_/Q _72350_/X _72351_/Y sky130_fd_sc_hd__o21ai_4
X_84337_ _83218_/CLK _63286_/Y _79259_/A sky130_fd_sc_hd__dfxtp_4
X_50729_ _50799_/A _51235_/B _50729_/Y sky130_fd_sc_hd__nand2_4
X_57285_ _57284_/Y _57285_/Y sky130_fd_sc_hd__inv_2
X_81549_ _83940_/CLK _76753_/X _81537_/D sky130_fd_sc_hd__dfxtp_4
X_54497_ _85431_/Q _54485_/X _54496_/Y _54497_/Y sky130_fd_sc_hd__o21ai_4
X_59024_ _59001_/X _86079_/Q _59023_/X _59024_/Y sky130_fd_sc_hd__o21ai_4
X_71302_ _70382_/A _71302_/X sky130_fd_sc_hd__buf_2
X_56236_ _56280_/A _56094_/X _56235_/Y _56236_/Y sky130_fd_sc_hd__o21ai_4
X_44250_ _68385_/A _59036_/A sky130_fd_sc_hd__buf_2
X_75070_ _81153_/D _80865_/Q _75070_/Y sky130_fd_sc_hd__xnor2_4
X_87056_ _87045_/CLK _87056_/D _44556_/A sky130_fd_sc_hd__dfxtp_4
X_41462_ _41461_/X _41455_/X _88211_/Q _41457_/X _41462_/X sky130_fd_sc_hd__a2bb2o_4
X_72282_ _72258_/X _85684_/Q _72146_/X _72282_/X sky130_fd_sc_hd__o21a_4
X_53448_ _53661_/A _53448_/X sky130_fd_sc_hd__buf_2
X_84268_ _84269_/CLK _64176_/Y _79921_/A sky130_fd_sc_hd__dfxtp_4
X_43201_ _43201_/A _43201_/Y sky130_fd_sc_hd__inv_2
X_74021_ _72880_/A _74021_/X sky130_fd_sc_hd__buf_2
X_86007_ _86005_/CLK _51457_/Y _86007_/Q sky130_fd_sc_hd__dfxtp_4
X_40413_ _40629_/A _40413_/X sky130_fd_sc_hd__buf_2
X_71233_ _48695_/B _71233_/A2 _71232_/Y _71233_/Y sky130_fd_sc_hd__o21ai_4
X_83219_ _84350_/CLK _72605_/Y _79279_/B sky130_fd_sc_hd__dfxtp_4
X_44181_ _64817_/A _44181_/X sky130_fd_sc_hd__buf_2
X_56167_ _56167_/A _56167_/B _56168_/A sky130_fd_sc_hd__xnor2_4
X_41393_ _41392_/Y _41393_/X sky130_fd_sc_hd__buf_2
X_53379_ _53352_/A _53386_/A sky130_fd_sc_hd__buf_2
X_84199_ _84194_/CLK _84199_/D _65466_/C sky130_fd_sc_hd__dfxtp_4
X_43132_ _43129_/X _43130_/X _40798_/X _43131_/Y _43127_/X _43132_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55118_ _55118_/A _47818_/A _55118_/Y sky130_fd_sc_hd__nand2_4
X_40344_ _40344_/A _46610_/A sky130_fd_sc_hd__buf_2
X_71164_ _71137_/A _71164_/B _71164_/Y sky130_fd_sc_hd__nor2_4
X_56098_ _56098_/A _55830_/X _56099_/A sky130_fd_sc_hd__xnor2_4
X_70115_ _70115_/A _70117_/C sky130_fd_sc_hd__inv_2
X_47940_ _57537_/B _48231_/B sky130_fd_sc_hd__buf_2
X_43063_ _43062_/Y _87591_/D sky130_fd_sc_hd__inv_2
X_55049_ _85328_/Q _55046_/X _55048_/Y _55049_/Y sky130_fd_sc_hd__o21ai_4
X_78760_ _78759_/X _78762_/A sky130_fd_sc_hd__inv_2
X_59926_ _59926_/A _59929_/C sky130_fd_sc_hd__buf_2
X_71095_ _71095_/A _71095_/X sky130_fd_sc_hd__buf_2
X_87958_ _87221_/CLK _42254_/Y _87958_/Q sky130_fd_sc_hd__dfxtp_4
X_75972_ _81706_/D _75972_/B _75981_/A sky130_fd_sc_hd__xor2_4
X_42014_ _42013_/X _42006_/X _40826_/X _73081_/A _42007_/X _42014_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77711_ _77712_/A _82124_/Q _77711_/Y sky130_fd_sc_hd__nor2_4
X_74923_ _74923_/A _74923_/B _74926_/A sky130_fd_sc_hd__nand2_4
X_70046_ _70040_/X _69800_/Y _70033_/X _70045_/Y _70046_/X sky130_fd_sc_hd__a211o_4
X_86909_ _86878_/CLK _44942_/Y _64235_/B sky130_fd_sc_hd__dfxtp_4
X_47871_ _47871_/A _48196_/A sky130_fd_sc_hd__buf_2
X_59857_ _59823_/X _59637_/A _59648_/A _59858_/A sky130_fd_sc_hd__nor3_4
X_78691_ _78691_/A _82684_/D _78691_/Y sky130_fd_sc_hd__nand2_4
X_87889_ _87625_/CLK _87889_/D _87889_/Q sky130_fd_sc_hd__dfxtp_4
X_49610_ _49610_/A _49592_/B _49615_/C _52827_/D _49610_/X sky130_fd_sc_hd__and4_4
X_46822_ _46830_/A _46830_/B _46830_/C _52694_/D _46822_/X sky130_fd_sc_hd__and4_4
X_58808_ _58696_/X _58804_/Y _58807_/Y _58728_/X _58701_/X _58808_/X
+ sky130_fd_sc_hd__o32a_4
X_77642_ _77627_/A _77626_/Y _77666_/A _77643_/B sky130_fd_sc_hd__o21a_4
X_74854_ _81124_/D _74854_/B _74865_/A sky130_fd_sc_hd__nor2_4
X_59788_ _59512_/A _59789_/A sky130_fd_sc_hd__buf_2
X_49541_ _49434_/A _49541_/X sky130_fd_sc_hd__buf_2
X_73805_ _73733_/A _85911_/Q _73805_/X sky130_fd_sc_hd__and2_4
X_46753_ _82963_/Q _46753_/Y sky130_fd_sc_hd__inv_2
X_58739_ _58857_/A _58739_/X sky130_fd_sc_hd__buf_2
X_77573_ _77572_/X _77575_/B sky130_fd_sc_hd__inv_2
X_43965_ _87174_/Q _43944_/A _43945_/A _43964_/X _43965_/X sky130_fd_sc_hd__a211o_4
X_74785_ _83838_/Q _74731_/X _74778_/X _74779_/X _74784_/Y _74785_/X
+ sky130_fd_sc_hd__a2111o_4
X_71997_ _83305_/Q _71985_/X _71996_/Y _71997_/Y sky130_fd_sc_hd__o21ai_4
X_79312_ _79324_/A _79324_/B _79334_/B sky130_fd_sc_hd__xor2_4
X_45704_ _55186_/B _45596_/X _45644_/X _45703_/Y _45704_/X sky130_fd_sc_hd__a211o_4
X_76524_ _76520_/Y _76521_/Y _76524_/C _76524_/X sky130_fd_sc_hd__or3_4
X_42916_ _42846_/X _42916_/X sky130_fd_sc_hd__buf_2
X_49472_ _49481_/A _46805_/X _49472_/Y sky130_fd_sc_hd__nand2_4
X_61750_ _61782_/A _61750_/B _61743_/Y _61749_/Y _61750_/Y sky130_fd_sc_hd__nand4_4
X_73736_ _73711_/A _66008_/B _73736_/X sky130_fd_sc_hd__and2_4
X_46684_ _83682_/Q _46685_/A sky130_fd_sc_hd__inv_2
X_70948_ _50744_/B _70937_/X _70947_/Y _70948_/Y sky130_fd_sc_hd__o21ai_4
X_43896_ _43756_/A _43896_/X sky130_fd_sc_hd__buf_2
X_48423_ _53647_/B _52128_/B sky130_fd_sc_hd__buf_2
X_60701_ _60692_/X _60694_/Y _60696_/Y _60698_/X _60700_/Y _60701_/Y
+ sky130_fd_sc_hd__a41oi_4
X_79243_ _79251_/B _79242_/Y _82823_/D sky130_fd_sc_hd__xor2_4
X_45635_ _45630_/X _45634_/X _45602_/X _45635_/X sky130_fd_sc_hd__a21o_4
X_76455_ _76455_/A _76455_/B _76456_/A sky130_fd_sc_hd__nor2_4
X_42847_ _42846_/X _42847_/X sky130_fd_sc_hd__buf_2
X_73667_ _73665_/X _84989_/Q _73614_/X _73666_/X _73667_/X sky130_fd_sc_hd__a211o_4
X_61681_ _61679_/X _61645_/X _61680_/Y _84460_/D sky130_fd_sc_hd__a21oi_4
X_70879_ _70712_/A _70880_/C sky130_fd_sc_hd__buf_2
X_63420_ _63456_/A _63456_/B _80579_/B _63420_/Y sky130_fd_sc_hd__nor3_4
X_75406_ _75369_/Y _75404_/X _75405_/Y _75406_/Y sky130_fd_sc_hd__a21oi_4
X_48354_ _48545_/A _48354_/X sky130_fd_sc_hd__buf_2
X_60632_ _60632_/A _60632_/X sky130_fd_sc_hd__buf_2
X_72618_ _72576_/Y _72522_/Y _72535_/Y _72618_/X sky130_fd_sc_hd__a21bo_4
X_79174_ _79174_/A _79173_/Y _79176_/A sky130_fd_sc_hd__nor2_4
X_45566_ _85014_/Q _55514_/B sky130_fd_sc_hd__inv_2
X_76386_ _76382_/Y _76361_/Y _76385_/X _76387_/B sky130_fd_sc_hd__o21ai_4
X_42778_ _41328_/X _42767_/X _87723_/Q _42768_/X _42778_/X sky130_fd_sc_hd__a2bb2o_4
X_73598_ _72852_/X _73599_/B sky130_fd_sc_hd__buf_2
X_47305_ _47305_/A _47306_/A sky130_fd_sc_hd__inv_2
X_78125_ _82568_/Q _78125_/B _78125_/Y sky130_fd_sc_hd__nand2_4
X_44517_ _44512_/X _44513_/X _40767_/A _44514_/Y _44516_/X _87071_/D
+ sky130_fd_sc_hd__o32ai_4
X_63351_ _63003_/Y _63347_/X _63350_/X _58374_/A _63020_/X _63351_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75337_ _75336_/X _75337_/Y sky130_fd_sc_hd__inv_2
X_41729_ _41729_/A _41718_/X _41729_/X sky130_fd_sc_hd__or2_4
X_60563_ _60500_/Y _60501_/Y _60602_/B _60583_/A _60479_/Y _60563_/X
+ sky130_fd_sc_hd__o41a_4
X_48285_ _86542_/Q _48263_/X _48284_/Y _48285_/Y sky130_fd_sc_hd__o21ai_4
X_72549_ _72525_/A _72549_/B _72549_/Y sky130_fd_sc_hd__nand2_4
X_45497_ _63079_/B _61406_/A sky130_fd_sc_hd__buf_2
X_62302_ _62267_/A _62267_/B _62302_/C _62302_/Y sky130_fd_sc_hd__nor3_4
X_47236_ _47236_/A _52934_/D sky130_fd_sc_hd__buf_2
X_66070_ _64589_/X _86230_/Q _45922_/X _66069_/X _66070_/X sky130_fd_sc_hd__a211o_4
X_78056_ _60810_/C _78056_/B _78056_/X sky130_fd_sc_hd__xor2_4
X_44448_ _44548_/A _44448_/X sky130_fd_sc_hd__buf_2
X_63282_ _63281_/X _63282_/Y sky130_fd_sc_hd__inv_2
X_75268_ _75269_/A _80944_/D _75268_/Y sky130_fd_sc_hd__nor2_4
X_60494_ _59755_/A _72590_/A sky130_fd_sc_hd__buf_2
X_65021_ _65019_/Y _64939_/X _65020_/X _84218_/D sky130_fd_sc_hd__a21o_4
X_77007_ _82083_/Q _77006_/Y _77007_/X sky130_fd_sc_hd__xor2_4
X_62233_ _61330_/X _59898_/A _62233_/C _62597_/D _62234_/D sky130_fd_sc_hd__nand4_4
X_74219_ _74216_/X _74218_/X _74220_/B sky130_fd_sc_hd__nand2_4
X_47167_ _47150_/A _52889_/B _47167_/Y sky130_fd_sc_hd__nand2_4
X_44379_ _44454_/A _44379_/X sky130_fd_sc_hd__buf_2
X_75199_ _80683_/Q _80983_/Q _75201_/A sky130_fd_sc_hd__xor2_4
X_46118_ _46117_/X _46119_/A sky130_fd_sc_hd__buf_2
X_62164_ _61715_/A _62160_/Y _62161_/Y _62163_/Y _62164_/Y sky130_fd_sc_hd__nand4_4
X_47098_ _83702_/Q _53369_/B sky130_fd_sc_hd__inv_2
X_61115_ _64285_/A _64474_/A sky130_fd_sc_hd__buf_2
X_46049_ _46049_/A _86795_/D sky130_fd_sc_hd__inv_2
X_69760_ _69746_/X _69758_/Y _69733_/X _69759_/Y _69760_/X sky130_fd_sc_hd__a211o_4
X_66972_ _66534_/A _66972_/X sky130_fd_sc_hd__buf_2
X_62095_ _61716_/X _61617_/B _62094_/X _62095_/X sky130_fd_sc_hd__a21o_4
X_78958_ _82738_/Q _78958_/B _78958_/X sky130_fd_sc_hd__xor2_4
X_68711_ _68516_/X _68701_/Y _68649_/X _68710_/Y _68711_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_7_42_0_CLK clkbuf_7_42_0_CLK/A clkbuf_8_85_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_65923_ _65920_/X _65922_/X _65304_/X _65923_/X sky130_fd_sc_hd__a21o_4
X_61046_ _61412_/A _61055_/A sky130_fd_sc_hd__buf_2
X_77909_ _77892_/A _77904_/A _77909_/X sky130_fd_sc_hd__and2_4
X_69691_ _69680_/A _88330_/Q _69691_/X sky130_fd_sc_hd__and2_4
X_78889_ _78889_/A _78889_/B _82699_/D sky130_fd_sc_hd__xor2_4
Xclkbuf_8_182_0_CLK clkbuf_7_91_0_CLK/X clkbuf_9_365_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_49808_ _49805_/Y _49787_/X _49807_/X _49808_/Y sky130_fd_sc_hd__a21oi_4
X_80920_ _84105_/CLK _84096_/Q _80920_/Q sky130_fd_sc_hd__dfxtp_4
X_68642_ _41922_/A _68640_/X _68439_/X _68641_/Y _68642_/X sky130_fd_sc_hd__a211o_4
X_65854_ _65789_/X _65333_/Y _65853_/Y _65854_/Y sky130_fd_sc_hd__o21ai_4
X_64805_ _64678_/X _85562_/Q _64679_/X _64804_/X _64805_/X sky130_fd_sc_hd__a211o_4
X_49739_ _49751_/A _49724_/B _49761_/C _52954_/D _49739_/X sky130_fd_sc_hd__and4_4
X_80851_ _80792_/CLK _80851_/D _74965_/B sky130_fd_sc_hd__dfxtp_4
X_68573_ _44691_/A _68570_/X _68571_/X _68572_/X _68573_/X sky130_fd_sc_hd__a211o_4
X_65785_ _65781_/X _65725_/B _65784_/X _65785_/Y sky130_fd_sc_hd__nand3_4
X_62997_ _59478_/A _60571_/B _61298_/B _60608_/A _62997_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_57_0_CLK clkbuf_7_57_0_CLK/A clkbuf_7_57_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_67524_ _67997_/A _67524_/X sky130_fd_sc_hd__buf_2
X_52750_ _52729_/X _52746_/B _52746_/C _52750_/D _52750_/X sky130_fd_sc_hd__and4_4
X_64736_ _64730_/X _64761_/B _64735_/X _64736_/Y sky130_fd_sc_hd__nand3_4
X_83570_ _86505_/CLK _71214_/Y _48614_/A sky130_fd_sc_hd__dfxtp_4
X_61948_ _61948_/A _61948_/X sky130_fd_sc_hd__buf_2
X_80782_ _80784_/CLK _80782_/D _80782_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_197_0_CLK clkbuf_7_98_0_CLK/X clkbuf_9_395_0_CLK/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_192_0_CLK clkbuf_9_96_0_CLK/X _83753_/CLK sky130_fd_sc_hd__clkbuf_1
X_51701_ _50219_/X _51701_/X sky130_fd_sc_hd__buf_2
X_82521_ _82617_/CLK _79023_/Y _82521_/Q sky130_fd_sc_hd__dfxtp_4
X_67455_ _67452_/X _67454_/X _67383_/X _67455_/X sky130_fd_sc_hd__a21o_4
X_52681_ _52674_/X _52661_/B _52694_/C _52681_/D _52681_/X sky130_fd_sc_hd__and4_4
X_64667_ _64667_/A _64767_/A sky130_fd_sc_hd__buf_2
X_61879_ _61879_/A _61879_/B _61875_/Y _61879_/D _61879_/Y sky130_fd_sc_hd__nand4_4
X_54420_ _85445_/Q _54404_/X _54419_/Y _54420_/Y sky130_fd_sc_hd__o21ai_4
X_66406_ _84129_/Q _66407_/C sky130_fd_sc_hd__inv_2
X_85240_ _85269_/CLK _85240_/D _55908_/B sky130_fd_sc_hd__dfxtp_4
X_51632_ _51627_/A _53157_/B _51632_/Y sky130_fd_sc_hd__nand2_4
X_63618_ _64454_/A _60732_/C _60739_/X _58490_/A _60704_/Y _63618_/Y
+ sky130_fd_sc_hd__o32ai_4
X_82452_ _82452_/CLK _79144_/X _82452_/Q sky130_fd_sc_hd__dfxtp_4
X_67386_ _87165_/Q _67311_/X _67313_/X _67385_/X _67386_/X sky130_fd_sc_hd__a211o_4
X_64598_ _64678_/A _64598_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_120_0_CLK clkbuf_7_60_0_CLK/X clkbuf_8_120_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_81403_ _81352_/CLK _83939_/Q _76728_/B sky130_fd_sc_hd__dfxtp_4
X_69125_ _69236_/A _69125_/B _69125_/X sky130_fd_sc_hd__and2_4
X_54351_ _54355_/A _52658_/B _54351_/Y sky130_fd_sc_hd__nand2_4
X_66337_ _64971_/X _85603_/Q _44261_/X _66336_/X _66337_/X sky130_fd_sc_hd__a211o_4
X_85171_ _85297_/CLK _85171_/D _55857_/B sky130_fd_sc_hd__dfxtp_4
X_51563_ _51553_/A _51580_/B _51553_/C _53090_/D _51563_/X sky130_fd_sc_hd__and4_4
X_63549_ _63523_/A _61969_/X _63549_/X sky130_fd_sc_hd__and2_4
X_82383_ _83703_/CLK _82191_/Q _47092_/A sky130_fd_sc_hd__dfxtp_4
X_53302_ _53302_/A _53302_/X sky130_fd_sc_hd__buf_2
X_84122_ _84220_/CLK _66446_/X _84122_/Q sky130_fd_sc_hd__dfxtp_4
X_50514_ _86186_/Q _50506_/X _50513_/Y _50514_/Y sky130_fd_sc_hd__o21ai_4
X_81334_ _81352_/CLK _76449_/X _81710_/D sky130_fd_sc_hd__dfxtp_4
X_57070_ _56971_/C _56971_/B _56995_/X _57069_/Y _57070_/X sky130_fd_sc_hd__a211o_4
X_69056_ _74206_/A _68989_/X _69010_/X _69055_/Y _69056_/X sky130_fd_sc_hd__a211o_4
X_54282_ _85470_/Q _54266_/X _54281_/Y _54282_/Y sky130_fd_sc_hd__o21ai_4
X_66268_ _66267_/X _85896_/Q _66268_/X sky130_fd_sc_hd__and2_4
X_51494_ _51509_/A _51494_/B _51494_/C _53019_/D _51494_/X sky130_fd_sc_hd__and4_4
X_56021_ _55686_/Y _56142_/A sky130_fd_sc_hd__buf_2
X_68007_ _68028_/A _87639_/Q _68007_/X sky130_fd_sc_hd__and2_4
X_53233_ _85672_/Q _53225_/X _53232_/Y _53233_/Y sky130_fd_sc_hd__o21ai_4
X_65219_ _65198_/X _65208_/Y _65218_/Y _65219_/Y sky130_fd_sc_hd__o21ai_4
X_84053_ _81431_/CLK _84053_/D _81485_/D sky130_fd_sc_hd__dfxtp_4
X_50445_ _50439_/X _48763_/B _50445_/Y sky130_fd_sc_hd__nand2_4
X_81265_ _81265_/CLK _81265_/D _76366_/A sky130_fd_sc_hd__dfxtp_4
X_66199_ _57947_/A _85613_/Q _65301_/X _66198_/X _66199_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_8_135_0_CLK clkbuf_7_67_0_CLK/X clkbuf_9_271_0_CLK/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_130_0_CLK clkbuf_9_65_0_CLK/X _81615_/CLK sky130_fd_sc_hd__clkbuf_1
X_83004_ _85050_/CLK _83004_/D _45479_/A sky130_fd_sc_hd__dfxtp_4
X_80216_ _80216_/A _80215_/X _80216_/Y sky130_fd_sc_hd__xnor2_4
X_53164_ _53190_/A _53181_/A sky130_fd_sc_hd__buf_2
X_50376_ _50381_/A _52079_/B _50376_/Y sky130_fd_sc_hd__nand2_4
X_81196_ _83974_/CLK _74969_/X _81196_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_760_0_CLK clkbuf_9_380_0_CLK/X _87776_/CLK sky130_fd_sc_hd__clkbuf_1
X_52115_ _52121_/A _48401_/B _52115_/Y sky130_fd_sc_hd__nand2_4
X_87812_ _87820_/CLK _42584_/Y _42583_/A sky130_fd_sc_hd__dfxtp_4
X_80147_ _80131_/Y _80134_/Y _80147_/X sky130_fd_sc_hd__or2_4
X_53095_ _53115_/A _53095_/B _53095_/Y sky130_fd_sc_hd__nand2_4
X_57972_ _86639_/Q _58039_/B _57972_/Y sky130_fd_sc_hd__nor2_4
X_69958_ _69958_/A _69958_/B _69958_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_9_251_0_CLK clkbuf_9_251_0_CLK/A clkbuf_9_251_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_59711_ _59696_/A _59711_/B _80579_/A _59711_/Y sky130_fd_sc_hd__nor3_4
X_52046_ _52044_/Y _52022_/X _52045_/Y _85900_/D sky130_fd_sc_hd__a21boi_4
X_56923_ _44282_/X _56922_/X _56923_/Y sky130_fd_sc_hd__nand2_4
X_68909_ _87581_/Q _66538_/X _66540_/X _68908_/X _68909_/X sky130_fd_sc_hd__a211o_4
X_87743_ _87748_/CLK _87743_/D _68868_/B sky130_fd_sc_hd__dfxtp_4
X_80078_ _80072_/Y _80077_/Y _80078_/X sky130_fd_sc_hd__xor2_4
X_84955_ _84714_/CLK _84955_/D _84955_/Q sky130_fd_sc_hd__dfxtp_4
X_69889_ _73370_/A _69796_/X _69797_/X _69888_/X _69889_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_145_0_CLK clkbuf_9_72_0_CLK/X _83184_/CLK sky130_fd_sc_hd__clkbuf_1
X_71920_ _71916_/Y _71920_/Y sky130_fd_sc_hd__inv_2
X_83906_ _83906_/CLK _83906_/D _81978_/D sky130_fd_sc_hd__dfxtp_4
X_59642_ _59634_/B _59661_/A _59662_/B _59661_/D _59642_/X sky130_fd_sc_hd__and4_4
X_56854_ _56852_/X _56853_/Y _44137_/A _56854_/X sky130_fd_sc_hd__a21o_4
X_87674_ _87675_/CLK _42873_/X _87674_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_775_0_CLK clkbuf_9_387_0_CLK/X _82617_/CLK sky130_fd_sc_hd__clkbuf_1
X_84886_ _84886_/CLK _84886_/D _84886_/Q sky130_fd_sc_hd__dfxtp_4
X_55805_ _44077_/X _56518_/C _55805_/X sky130_fd_sc_hd__and2_4
X_86625_ _84922_/CLK _47534_/Y _86625_/Q sky130_fd_sc_hd__dfxtp_4
X_71851_ _70884_/B _71851_/X sky130_fd_sc_hd__buf_2
X_59573_ _59557_/A _59890_/B _59741_/C _59574_/A sky130_fd_sc_hd__nand3_4
X_83837_ _83835_/CLK _83837_/D _74773_/C sky130_fd_sc_hd__dfxtp_4
X_56785_ _56782_/X _56785_/B _56783_/X _56785_/D _56786_/A sky130_fd_sc_hd__and4_4
Xclkbuf_9_266_0_CLK clkbuf_9_267_0_CLK/A clkbuf_9_266_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_53997_ _53929_/A _53998_/A sky130_fd_sc_hd__buf_2
X_70802_ _70802_/A _70802_/X sky130_fd_sc_hd__buf_2
X_58524_ _63520_/B _58510_/X _58524_/Y sky130_fd_sc_hd__nor2_4
X_55736_ _55741_/A _55736_/B _55736_/X sky130_fd_sc_hd__and2_4
X_43750_ _40935_/X _43736_/X _87283_/Q _43737_/X _87283_/D sky130_fd_sc_hd__a2bb2o_4
X_74570_ _74600_/A _74570_/X sky130_fd_sc_hd__buf_2
X_86556_ _86560_/CLK _86556_/D _73689_/B sky130_fd_sc_hd__dfxtp_4
X_40962_ _40790_/B _40932_/X _40962_/X sky130_fd_sc_hd__or2_4
X_52948_ _52947_/X _52954_/B _52926_/X _52948_/D _52948_/X sky130_fd_sc_hd__and4_4
X_71782_ _71713_/Y _71783_/C sky130_fd_sc_hd__buf_2
X_83768_ _83482_/CLK _70471_/X _83768_/Q sky130_fd_sc_hd__dfxtp_4
X_42701_ _42687_/X _42688_/X _41116_/X _68343_/B _42700_/X _42701_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73521_ _73521_/A _73521_/B _73521_/Y sky130_fd_sc_hd__nand2_4
X_85507_ _85507_/CLK _54088_/Y _85507_/Q sky130_fd_sc_hd__dfxtp_4
X_70733_ HASH_ADDR[3] _70495_/A _70733_/Y sky130_fd_sc_hd__nor2_4
X_58455_ _84844_/Q _58457_/A sky130_fd_sc_hd__buf_2
X_82719_ _82715_/CLK _82719_/D _82675_/D sky130_fd_sc_hd__dfxtp_4
X_43681_ _40781_/X _43671_/X _72831_/A _43673_/X _43681_/X sky130_fd_sc_hd__a2bb2o_4
X_55667_ _55661_/X _55664_/Y _55665_/Y _55666_/Y _55676_/A sky130_fd_sc_hd__and4_4
X_86487_ _86196_/CLK _86487_/D _73042_/B sky130_fd_sc_hd__dfxtp_4
X_40893_ _40857_/X _82281_/Q _40892_/X _40894_/A sky130_fd_sc_hd__o21a_4
X_52879_ _52867_/A _52879_/B _52872_/C _52879_/D _52879_/X sky130_fd_sc_hd__and4_4
X_83699_ _83699_/CLK _70792_/Y _83699_/Q sky130_fd_sc_hd__dfxtp_4
X_45420_ _45350_/X _61338_/A _45370_/X _45420_/Y sky130_fd_sc_hd__o21ai_4
X_57406_ _57484_/A _56643_/X _85011_/Q _57380_/X _85011_/D sky130_fd_sc_hd__a2bb2o_4
X_76240_ _76209_/Y _76223_/Y _76240_/Y sky130_fd_sc_hd__nand2_4
X_88226_ _88224_/CLK _41378_/Y _67756_/B sky130_fd_sc_hd__dfxtp_4
X_42632_ _42449_/Y _42680_/A sky130_fd_sc_hd__buf_2
X_54618_ _54537_/A _54618_/X sky130_fd_sc_hd__buf_2
X_73452_ _73497_/A _86470_/Q _73452_/X sky130_fd_sc_hd__and2_4
X_85438_ _85439_/CLK _85438_/D _85438_/Q sky130_fd_sc_hd__dfxtp_4
X_70664_ _70664_/A _70664_/X sky130_fd_sc_hd__buf_2
X_58386_ _58385_/Y _58369_/X _58386_/Y sky130_fd_sc_hd__nand2_4
X_55598_ _55595_/X _55597_/X _55517_/X _55601_/A sky130_fd_sc_hd__a21o_4
X_72403_ _72394_/Y _72358_/X _72399_/X _72402_/X _83258_/D sky130_fd_sc_hd__a22oi_4
X_57337_ _57289_/B _56849_/X _57337_/Y sky130_fd_sc_hd__nor2_4
X_45351_ _64535_/B _61673_/B sky130_fd_sc_hd__buf_2
X_76171_ _76171_/A _76171_/B _76171_/Y sky130_fd_sc_hd__nor2_4
X_88157_ _87144_/CLK _88157_/D _67873_/B sky130_fd_sc_hd__dfxtp_4
X_42563_ _42554_/X _42547_/X _40806_/X _69676_/B _42556_/X _87819_/D
+ sky130_fd_sc_hd__o32ai_4
X_54549_ _54538_/A _54559_/B _54538_/C _47103_/Y _54549_/X sky130_fd_sc_hd__and4_4
X_73383_ _72877_/A _73383_/X sky130_fd_sc_hd__buf_2
X_85369_ _83275_/CLK _85369_/D _85369_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_713_0_CLK clkbuf_9_356_0_CLK/X _88247_/CLK sky130_fd_sc_hd__clkbuf_1
X_70595_ _70585_/X _70613_/B _74533_/D _70594_/X _70595_/Y sky130_fd_sc_hd__nand4_4
X_44302_ _44300_/Y _44313_/A sky130_fd_sc_hd__inv_2
X_87108_ _87110_/CLK _87108_/D _87108_/Q sky130_fd_sc_hd__dfxtp_4
X_75122_ _75122_/A _75122_/Y sky130_fd_sc_hd__inv_2
X_41514_ _41344_/X _40430_/B _41513_/X _41514_/X sky130_fd_sc_hd__o21a_4
X_48070_ _48063_/Y _48055_/X _48069_/X _48070_/Y sky130_fd_sc_hd__a21oi_4
X_72334_ _72323_/Y _72237_/X _72330_/X _72333_/X _83264_/D sky130_fd_sc_hd__a22oi_4
X_45282_ _55748_/B _45281_/X _45237_/X _45282_/X sky130_fd_sc_hd__o21a_4
X_57268_ _57267_/X _57268_/X sky130_fd_sc_hd__buf_2
X_42494_ _42494_/A _87846_/D sky130_fd_sc_hd__inv_2
X_88088_ _88086_/CLK _41970_/Y _88088_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_204_0_CLK clkbuf_8_102_0_CLK/X clkbuf_9_204_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_47021_ _47029_/A _47029_/B _47029_/C _52805_/D _47021_/X sky130_fd_sc_hd__and4_4
X_59007_ _58897_/A _59008_/B sky130_fd_sc_hd__buf_2
X_44233_ _72814_/A _73181_/A sky130_fd_sc_hd__buf_2
X_56219_ _56214_/A _56229_/B _56219_/C _56219_/Y sky130_fd_sc_hd__nand3_4
X_75053_ _75046_/X _75053_/B _75053_/X sky130_fd_sc_hd__xor2_4
X_79930_ _79928_/B _79928_/A _79931_/B sky130_fd_sc_hd__nand2_4
X_41445_ _41784_/B _41435_/B _41445_/X sky130_fd_sc_hd__or2_4
X_87039_ _86989_/CLK _44604_/X _87039_/Q sky130_fd_sc_hd__dfxtp_4
X_72265_ _72180_/X _85333_/Q _72225_/X _72265_/X sky130_fd_sc_hd__o21a_4
X_57199_ _57199_/A _44282_/X _57199_/Y sky130_fd_sc_hd__nor2_4
X_74004_ _70108_/Y _73939_/X _74003_/Y _74004_/Y sky130_fd_sc_hd__o21ai_4
X_71216_ _71216_/A _71216_/X sky130_fd_sc_hd__buf_2
X_44164_ _44024_/A _44164_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_728_0_CLK clkbuf_9_364_0_CLK/X _88288_/CLK sky130_fd_sc_hd__clkbuf_1
X_79861_ _64688_/Y _72151_/Y _79860_/Y _79861_/X sky130_fd_sc_hd__o21a_4
X_41376_ _41376_/A _41376_/X sky130_fd_sc_hd__buf_2
X_72196_ _59345_/X _72196_/X sky130_fd_sc_hd__buf_2
X_43115_ _43115_/A _43115_/Y sky130_fd_sc_hd__inv_2
X_78812_ _78812_/A _82835_/Q _79122_/A sky130_fd_sc_hd__nand2_4
X_40327_ _40629_/A _40878_/A sky130_fd_sc_hd__buf_2
X_71147_ _71173_/A _71155_/B _71152_/C _70875_/X _71147_/Y sky130_fd_sc_hd__nand4_4
X_48972_ _48972_/A _48973_/A sky130_fd_sc_hd__inv_2
X_44095_ _44095_/A _44095_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_219_0_CLK clkbuf_9_219_0_CLK/A clkbuf_9_219_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_79792_ _79770_/Y _79788_/X _79791_/Y _79793_/B sky130_fd_sc_hd__a21oi_4
X_47923_ _73765_/A _47924_/B sky130_fd_sc_hd__buf_2
X_59909_ _59909_/A _63632_/A _59909_/C _59909_/Y sky130_fd_sc_hd__nand3_4
X_43046_ _43046_/A _43046_/X sky130_fd_sc_hd__buf_2
X_78743_ _78717_/X _78722_/Y _78744_/C sky130_fd_sc_hd__nand2_4
X_71078_ _71078_/A _71055_/B _71078_/C _71078_/Y sky130_fd_sc_hd__nand3_4
X_75955_ _81511_/Q _75955_/B _75955_/X sky130_fd_sc_hd__xor2_4
X_74906_ _74906_/A _74906_/B _74906_/X sky130_fd_sc_hd__xor2_4
X_62920_ _62916_/Y _60337_/A _62660_/X _62918_/X _62919_/Y _62920_/X
+ sky130_fd_sc_hd__a41o_4
Xclkbuf_4_4_0_CLK clkbuf_4_5_0_CLK/A clkbuf_4_4_1_CLK/A sky130_fd_sc_hd__clkbuf_1
X_70029_ _70048_/A _70029_/X sky130_fd_sc_hd__buf_2
X_47854_ _47853_/Y _50232_/B sky130_fd_sc_hd__buf_2
X_78674_ _78672_/Y _78642_/Y _78673_/X _78675_/B sky130_fd_sc_hd__o21ai_4
X_75886_ _75817_/Y _75886_/Y sky130_fd_sc_hd__inv_2
X_46805_ _52686_/B _46805_/X sky130_fd_sc_hd__buf_2
X_77625_ _77606_/A _77623_/Y _77624_/Y _77625_/X sky130_fd_sc_hd__a21bo_4
X_62851_ _62851_/A _63306_/A sky130_fd_sc_hd__buf_2
X_74837_ _74836_/Y _80655_/D sky130_fd_sc_hd__inv_2
X_47785_ _47804_/A _47777_/B _47777_/C _53244_/D _47785_/X sky130_fd_sc_hd__and4_4
X_44997_ _44987_/X _44991_/Y _44996_/Y _44997_/Y sky130_fd_sc_hd__a21oi_4
X_61802_ _61752_/A _61723_/X _78076_/B _61802_/Y sky130_fd_sc_hd__nor3_4
X_49524_ _49496_/A _49524_/X sky130_fd_sc_hd__buf_2
X_46736_ _46735_/Y _46736_/X sky130_fd_sc_hd__buf_2
X_65570_ _65524_/X _83072_/Q _65568_/X _65569_/X _65570_/X sky130_fd_sc_hd__a211o_4
X_77556_ _77555_/X _77556_/Y sky130_fd_sc_hd__inv_2
X_43948_ _43979_/A _43948_/B _43948_/Y sky130_fd_sc_hd__nor2_4
X_62782_ _60199_/X _62782_/X sky130_fd_sc_hd__buf_2
X_74768_ _74723_/X _74768_/B _74780_/D _74768_/Y sky130_fd_sc_hd__nand3_4
X_76507_ _76487_/Y _76491_/B _76489_/Y _76508_/A sky130_fd_sc_hd__o21a_4
X_64521_ _64315_/A _64521_/X sky130_fd_sc_hd__buf_2
X_49455_ _86384_/Q _49443_/X _49454_/Y _49455_/Y sky130_fd_sc_hd__o21ai_4
X_61733_ _61730_/X _61791_/B _61732_/X _63017_/B _61733_/X sky130_fd_sc_hd__and4_4
X_73719_ _73717_/X _73719_/B _73719_/C _73719_/Y sky130_fd_sc_hd__nand3_4
X_46667_ _46667_/A _46682_/C sky130_fd_sc_hd__buf_2
X_77487_ _77488_/A _77488_/B _77487_/Y sky130_fd_sc_hd__nor2_4
X_43879_ _43842_/A _43879_/X sky130_fd_sc_hd__buf_2
X_74699_ _74698_/Y _82981_/D sky130_fd_sc_hd__inv_2
X_48406_ _48134_/X _82365_/Q _48405_/X _48407_/A sky130_fd_sc_hd__o21ai_4
X_67240_ _66879_/A _67240_/X sky130_fd_sc_hd__buf_2
X_79226_ _79251_/A _79225_/Y _79227_/A sky130_fd_sc_hd__xor2_4
X_45618_ _45615_/Y _45570_/X _45616_/X _45617_/Y _45618_/X sky130_fd_sc_hd__a211o_4
X_64452_ _64445_/Y _64451_/X _64442_/X _64452_/X sky130_fd_sc_hd__o21a_4
X_76438_ _76438_/A _76440_/A sky130_fd_sc_hd__inv_2
X_61664_ _64526_/B _61665_/B sky130_fd_sc_hd__buf_2
X_49386_ _49397_/A _49369_/X _49408_/C _51772_/D _49386_/X sky130_fd_sc_hd__and4_4
X_46598_ _72083_/A _46598_/X sky130_fd_sc_hd__buf_2
X_63403_ _63368_/X _63396_/X _63397_/X _63401_/X _63402_/Y _63403_/Y
+ sky130_fd_sc_hd__o41ai_4
X_60615_ _60615_/A _60312_/C _60312_/D _60616_/B sky130_fd_sc_hd__nand3_4
X_48337_ _48337_/A _52079_/B sky130_fd_sc_hd__buf_2
X_67171_ _87418_/Q _67121_/X _67122_/X _67170_/X _67171_/X sky130_fd_sc_hd__a211o_4
X_79157_ _79157_/A _84489_/Q _82465_/D sky130_fd_sc_hd__xor2_4
X_45549_ _45549_/A _45597_/B _45549_/Y sky130_fd_sc_hd__nor2_4
X_64383_ _58335_/Y _64367_/X _64382_/Y _64383_/Y sky130_fd_sc_hd__o21ai_4
X_76369_ _76369_/A _76369_/B _76368_/Y _76369_/X sky130_fd_sc_hd__or3_4
X_61595_ _72528_/A _61611_/B sky130_fd_sc_hd__buf_2
X_66122_ _66068_/X _65646_/Y _66121_/Y _66122_/Y sky130_fd_sc_hd__o21ai_4
X_78108_ _82567_/Q _78108_/B _78130_/B sky130_fd_sc_hd__xor2_4
X_63334_ _63330_/Y _63331_/X _63332_/X _63333_/X _63020_/A _63334_/Y
+ sky130_fd_sc_hd__o41ai_4
X_48268_ _48545_/A _48287_/C sky130_fd_sc_hd__buf_2
X_60546_ _60546_/A _60546_/Y sky130_fd_sc_hd__inv_2
X_79088_ _79088_/A _79088_/Y sky130_fd_sc_hd__inv_2
X_47219_ _47215_/Y _47177_/X _47218_/X _47219_/Y sky130_fd_sc_hd__a21oi_4
X_66053_ _66053_/A _66053_/X sky130_fd_sc_hd__buf_2
X_78039_ _77883_/Y _81939_/D sky130_fd_sc_hd__inv_2
X_63265_ _63216_/X _63265_/B _63333_/C _63240_/X _63265_/X sky130_fd_sc_hd__and4_4
X_48199_ _86557_/Q _48188_/X _48198_/Y _48199_/Y sky130_fd_sc_hd__o21ai_4
X_60477_ _60477_/A _60519_/B _79153_/A _60477_/Y sky130_fd_sc_hd__nor3_4
X_65004_ _65001_/X _65003_/X _64959_/X _65004_/X sky130_fd_sc_hd__a21o_4
X_50230_ _50230_/A _48178_/X _50230_/Y sky130_fd_sc_hd__nand2_4
X_81050_ _81048_/CLK _75440_/B _81050_/Q sky130_fd_sc_hd__dfxtp_4
X_62216_ _62181_/A _62181_/B _84425_/Q _62216_/Y sky130_fd_sc_hd__nor3_4
X_63196_ _63157_/X _63196_/B _63241_/C _63181_/X _63196_/X sky130_fd_sc_hd__and4_4
X_80001_ _79989_/Y _79992_/Y _79988_/A _80002_/B sky130_fd_sc_hd__o21ai_4
X_69812_ _87053_/Q _69796_/X _69797_/X _69811_/X _69813_/B sky130_fd_sc_hd__a211o_4
X_50161_ _50159_/Y _50141_/X _50160_/X _86252_/D sky130_fd_sc_hd__a21oi_4
X_62147_ _59730_/A _62170_/B _62158_/C _63324_/B _62147_/X sky130_fd_sc_hd__and4_4
X_69743_ _69739_/X _69741_/X _69742_/X _69743_/Y sky130_fd_sc_hd__a21oi_4
X_50092_ _50092_/A _50092_/X sky130_fd_sc_hd__buf_2
X_66955_ _66717_/A _66955_/X sky130_fd_sc_hd__buf_2
X_62078_ _62070_/X _62072_/X _62077_/Y _84843_/Q _62048_/X _62078_/Y
+ sky130_fd_sc_hd__o32ai_4
X_53920_ _53918_/Y _53914_/X _53919_/Y _53920_/Y sky130_fd_sc_hd__a21boi_4
X_65906_ _65932_/A _73561_/B _65906_/X sky130_fd_sc_hd__and2_4
X_61029_ _61028_/X _61030_/A sky130_fd_sc_hd__inv_2
X_84740_ _83766_/CLK _84740_/D _84740_/Q sky130_fd_sc_hd__dfxtp_4
X_69674_ _87563_/Q _69645_/X _68613_/X _69673_/X _69674_/X sky130_fd_sc_hd__a211o_4
X_81952_ _82145_/CLK _78024_/Y _81952_/Q sky130_fd_sc_hd__dfxtp_4
X_66886_ _66886_/A _66885_/X _66886_/Y sky130_fd_sc_hd__nand2_4
X_80903_ _83933_/CLK _80903_/D _75621_/A sky130_fd_sc_hd__dfxtp_4
X_68625_ _88009_/Q _68527_/X _68501_/X _68624_/X _68625_/X sky130_fd_sc_hd__a211o_4
X_53851_ _53849_/Y _53838_/X _53850_/Y _85556_/D sky130_fd_sc_hd__a21boi_4
X_65837_ _64696_/X _85574_/Q _64697_/X _65836_/X _65837_/X sky130_fd_sc_hd__a211o_4
X_84671_ _84671_/CLK _84671_/D _60047_/C sky130_fd_sc_hd__dfxtp_4
X_81883_ _81883_/CLK _78074_/X _81883_/Q sky130_fd_sc_hd__dfxtp_4
X_86410_ _86127_/CLK _86410_/D _86410_/Q sky130_fd_sc_hd__dfxtp_4
X_52802_ _52800_/Y _52783_/X _52801_/X _85752_/D sky130_fd_sc_hd__a21oi_4
X_83622_ _83310_/CLK _71059_/Y _83622_/Q sky130_fd_sc_hd__dfxtp_4
X_56570_ _56564_/C _56569_/X _56570_/Y sky130_fd_sc_hd__xnor2_4
X_80834_ _80835_/CLK _80834_/D _74848_/B sky130_fd_sc_hd__dfxtp_4
X_68556_ _68366_/X _42475_/Y _68556_/Y sky130_fd_sc_hd__nor2_4
X_87390_ _87644_/CLK _87390_/D _87390_/Q sky130_fd_sc_hd__dfxtp_4
X_53782_ _48885_/A _53774_/B _53774_/C _53782_/X sky130_fd_sc_hd__and3_4
X_65768_ _65768_/A _65768_/X sky130_fd_sc_hd__buf_2
X_50994_ _51003_/A _46805_/X _50994_/Y sky130_fd_sc_hd__nand2_4
X_55521_ _45549_/A _55511_/X _55506_/X _55520_/Y _55521_/X sky130_fd_sc_hd__a211o_4
X_67507_ _67863_/A _67507_/X sky130_fd_sc_hd__buf_2
X_86341_ _86342_/CLK _49693_/Y _86341_/Q sky130_fd_sc_hd__dfxtp_4
X_52733_ _85764_/Q _52711_/X _52732_/Y _52733_/Y sky130_fd_sc_hd__o21ai_4
X_64719_ _64826_/A _64719_/B _64719_/X sky130_fd_sc_hd__and2_4
X_83553_ _83550_/CLK _71270_/Y _83553_/Q sky130_fd_sc_hd__dfxtp_4
X_80765_ _80817_/CLK _75493_/Y _81141_/D sky130_fd_sc_hd__dfxtp_4
X_68487_ _68484_/X _68486_/X _68331_/X _68487_/Y sky130_fd_sc_hd__a21oi_4
X_65699_ _65696_/Y _65681_/X _65698_/X _84184_/D sky130_fd_sc_hd__a21o_4
X_58240_ _58240_/A _58240_/Y sky130_fd_sc_hd__inv_2
X_82504_ _81198_/CLK _78852_/X _82504_/Q sky130_fd_sc_hd__dfxtp_4
X_55452_ _55394_/Y _55444_/Y _55676_/B _55650_/A sky130_fd_sc_hd__o21ai_4
X_67438_ _87983_/Q _67414_/X _67391_/X _67437_/X _67438_/X sky130_fd_sc_hd__a211o_4
X_86272_ _83310_/CLK _50060_/Y _64627_/B sky130_fd_sc_hd__dfxtp_4
X_52664_ _85777_/Q _52656_/X _52663_/Y _52664_/Y sky130_fd_sc_hd__o21ai_4
X_83484_ _83414_/CLK _83484_/D _83484_/Q sky130_fd_sc_hd__dfxtp_4
X_80696_ _80696_/CLK _80696_/D _75393_/A sky130_fd_sc_hd__dfxtp_4
X_88011_ _87757_/CLK _88011_/D _88011_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_704 sky130_fd_sc_hd__decap_3
X_54403_ _54398_/Y _54394_/X _54402_/X _54403_/Y sky130_fd_sc_hd__a21oi_4
X_85223_ _85190_/CLK _85223_/D _55756_/B sky130_fd_sc_hd__dfxtp_4
X_51615_ _51619_/A _51619_/B _51608_/X _53139_/D _51615_/X sky130_fd_sc_hd__and4_4
X_58171_ _58253_/A _58171_/X sky130_fd_sc_hd__buf_2
X_82435_ _82443_/CLK _79127_/X _82435_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_715 sky130_fd_sc_hd__decap_3
X_55383_ _55383_/A _55384_/A _55383_/C _56719_/A sky130_fd_sc_hd__nand3_4
X_67369_ _87986_/Q _67293_/X _67271_/X _67368_/X _67369_/X sky130_fd_sc_hd__a211o_4
X_52595_ _52591_/Y _52592_/X _52594_/X _85790_/D sky130_fd_sc_hd__a21oi_4
X_57122_ _57121_/X _56643_/X _45611_/A _57192_/A _85075_/D sky130_fd_sc_hd__a2bb2o_4
X_69108_ _80803_/D _69066_/X _69107_/X _83947_/D sky130_fd_sc_hd__a21bo_4
X_54334_ _54325_/A _54353_/B _54317_/X _46735_/Y _54334_/X sky130_fd_sc_hd__and4_4
X_85154_ _82993_/CLK _85154_/D _55738_/B sky130_fd_sc_hd__dfxtp_4
X_51546_ _85990_/Q _51539_/X _51545_/Y _51546_/Y sky130_fd_sc_hd__o21ai_4
X_70380_ _50858_/B _70364_/X _70379_/Y _70380_/Y sky130_fd_sc_hd__o21ai_4
X_82366_ _83133_/CLK _82366_/D _82366_/Q sky130_fd_sc_hd__dfxtp_4
X_84105_ _84105_/CLK _84105_/D _84105_/Q sky130_fd_sc_hd__dfxtp_4
X_81317_ _84105_/CLK _76199_/Y _81725_/D sky130_fd_sc_hd__dfxtp_4
X_57053_ _57052_/X _85096_/D sky130_fd_sc_hd__inv_2
X_69039_ _69036_/X _69038_/X _69017_/X _69039_/Y sky130_fd_sc_hd__a21oi_4
X_54265_ _54262_/Y _54253_/X _54264_/X _54265_/Y sky130_fd_sc_hd__a21oi_4
X_85085_ _85152_/CLK _85085_/D _45455_/A sky130_fd_sc_hd__dfxtp_4
X_51477_ _51557_/A _51477_/X sky130_fd_sc_hd__buf_2
X_82297_ _82343_/CLK _81921_/Q _82297_/Q sky130_fd_sc_hd__dfxtp_4
X_56004_ _74286_/C _56003_/Y _56004_/X sky130_fd_sc_hd__xor2_4
X_41230_ _41230_/A _41230_/X sky130_fd_sc_hd__buf_2
X_53216_ _53190_/A _53217_/A sky130_fd_sc_hd__buf_2
X_72050_ _72047_/Y _71978_/X _72049_/X _72050_/Y sky130_fd_sc_hd__a21oi_4
X_84036_ _81160_/CLK _68113_/X _82076_/D sky130_fd_sc_hd__dfxtp_4
X_50428_ _86202_/Q _50403_/X _50427_/Y _50428_/Y sky130_fd_sc_hd__o21ai_4
X_81248_ _85375_/CLK _81056_/Q _47539_/A sky130_fd_sc_hd__dfxtp_4
X_54196_ _85486_/Q _54193_/X _54195_/Y _54196_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_190_0_CLK clkbuf_8_95_0_CLK/X clkbuf_9_190_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_71001_ _70990_/A _70952_/B _71001_/C _71001_/Y sky130_fd_sc_hd__nand3_4
X_53147_ _53147_/A _53147_/X sky130_fd_sc_hd__buf_2
X_41161_ _41161_/A _41161_/X sky130_fd_sc_hd__buf_2
X_50359_ _86216_/Q _50333_/X _50358_/Y _50359_/Y sky130_fd_sc_hd__o21ai_4
X_81179_ _81179_/CLK _75028_/B _81179_/Q sky130_fd_sc_hd__dfxtp_4
X_41092_ _41024_/X _41266_/A _41091_/X _41092_/Y sky130_fd_sc_hd__o21ai_4
X_53078_ _53074_/A _53069_/X _53074_/C _53078_/D _53078_/X sky130_fd_sc_hd__and4_4
X_57955_ _86641_/Q _57954_/X _57955_/Y sky130_fd_sc_hd__nor2_4
X_85987_ _85700_/CLK _51564_/Y _85987_/Q sky130_fd_sc_hd__dfxtp_4
X_44920_ _85312_/Q _45876_/B _44919_/X _44920_/Y sky130_fd_sc_hd__o21ai_4
X_52029_ _52058_/A _50326_/B _52029_/Y sky130_fd_sc_hd__nand2_4
X_56906_ _55227_/A _55225_/X _56906_/X sky130_fd_sc_hd__and2_4
X_75740_ _75735_/Y _75740_/B _75741_/B sky130_fd_sc_hd__xor2_4
X_87726_ _87472_/CLK _42771_/X _67451_/B sky130_fd_sc_hd__dfxtp_4
X_72952_ _72946_/X _72948_/X _72951_/X _72969_/B sky130_fd_sc_hd__a21o_4
X_84938_ _83736_/CLK _57943_/Y _84938_/Q sky130_fd_sc_hd__dfxtp_4
X_57886_ _57760_/X _85398_/Q _57885_/X _57886_/Y sky130_fd_sc_hd__o21ai_4
X_71903_ _70383_/X _71893_/X _71902_/X _71898_/D _71903_/Y sky130_fd_sc_hd__nand4_4
X_59625_ _59624_/X _59664_/A sky130_fd_sc_hd__buf_2
X_44851_ _41748_/Y _44848_/X _86920_/Q _44849_/X _86920_/D sky130_fd_sc_hd__a2bb2o_4
X_56837_ _56698_/Y _56836_/Y _56713_/A _56707_/X _56837_/X sky130_fd_sc_hd__a211o_4
X_75671_ _75657_/Y _80780_/D sky130_fd_sc_hd__inv_2
X_87657_ _87397_/CLK _42910_/Y _87657_/Q sky130_fd_sc_hd__dfxtp_4
X_72883_ _72883_/A _72883_/B _72884_/B sky130_fd_sc_hd__nand2_4
X_84869_ _84869_/CLK _84869_/D _84869_/Q sky130_fd_sc_hd__dfxtp_4
X_77410_ _77409_/A _82095_/D _77410_/Y sky130_fd_sc_hd__nand2_4
X_43802_ _43802_/A _43802_/X sky130_fd_sc_hd__buf_2
X_86608_ _86610_/CLK _86608_/D _72332_/A sky130_fd_sc_hd__dfxtp_4
X_74622_ _45347_/A _74612_/X _74621_/X _83012_/D sky130_fd_sc_hd__o21ai_4
X_47570_ _47619_/A _47570_/X sky130_fd_sc_hd__buf_2
X_71834_ _71825_/X _83359_/Q _71833_/X _83359_/D sky130_fd_sc_hd__a21o_4
X_59556_ _61276_/B _60599_/A sky130_fd_sc_hd__buf_2
X_78390_ _78390_/A _82792_/Q _78385_/Y _78394_/B sky130_fd_sc_hd__nand3_4
X_44782_ _44766_/X _44767_/X _41381_/X _86957_/Q _44768_/X _44783_/A
+ sky130_fd_sc_hd__o32ai_4
X_56768_ _56653_/Y _56768_/Y sky130_fd_sc_hd__inv_2
X_87588_ _87588_/CLK _43069_/Y _43068_/A sky130_fd_sc_hd__dfxtp_4
X_41994_ _88078_/Q _41994_/Y sky130_fd_sc_hd__inv_2
X_46521_ _46434_/A _51358_/B _46521_/Y sky130_fd_sc_hd__nand2_4
X_58507_ _58492_/X _58504_/Y _58506_/Y _84832_/D sky130_fd_sc_hd__a21oi_4
X_77341_ _77326_/Y _77323_/Y _77325_/A _77341_/X sky130_fd_sc_hd__o21a_4
X_43733_ _40894_/A _43716_/X _69885_/B _43718_/X _43733_/X sky130_fd_sc_hd__a2bb2o_4
X_55719_ _45345_/A _55710_/B _55719_/Y sky130_fd_sc_hd__nand2_4
X_74553_ _74552_/X _74553_/X sky130_fd_sc_hd__buf_2
X_86539_ _86210_/CLK _86539_/D _86539_/Q sky130_fd_sc_hd__dfxtp_4
X_40945_ _40637_/A _40946_/A sky130_fd_sc_hd__buf_2
X_71765_ _71762_/X _83385_/Q _71764_/X _83385_/D sky130_fd_sc_hd__a21o_4
X_59487_ _46159_/X _59484_/Y _59486_/Y _59487_/Y sky130_fd_sc_hd__a21oi_4
X_56699_ _83336_/Q _56842_/A sky130_fd_sc_hd__inv_2
X_49240_ _49238_/Y _49214_/X _49239_/Y _86427_/D sky130_fd_sc_hd__a21boi_4
X_73504_ _73494_/Y _73503_/X _73505_/B sky130_fd_sc_hd__xnor2_4
X_70716_ _70716_/A _70727_/C sky130_fd_sc_hd__buf_2
X_46452_ _53874_/A _46472_/C sky130_fd_sc_hd__buf_2
X_58438_ _58438_/A _58426_/X _58438_/Y sky130_fd_sc_hd__nand2_4
X_77272_ _77261_/A _77260_/A _77258_/Y _77272_/Y sky130_fd_sc_hd__o21ai_4
X_43664_ _40729_/X _43656_/X _74145_/A _43657_/X _87322_/D sky130_fd_sc_hd__a2bb2o_4
X_74484_ _74481_/Y _74463_/X _74483_/X _83057_/D sky130_fd_sc_hd__a21oi_4
X_40876_ _40875_/Y _88319_/D sky130_fd_sc_hd__inv_2
X_71696_ _71338_/A _71685_/X _71297_/X _71696_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_652_0_CLK clkbuf_9_326_0_CLK/X _87397_/CLK sky130_fd_sc_hd__clkbuf_1
X_79011_ _79011_/A _79011_/B _79011_/X sky130_fd_sc_hd__xor2_4
X_45403_ _83009_/Q _45401_/X _45402_/X _45403_/Y sky130_fd_sc_hd__o21ai_4
X_76223_ _76220_/Y _76222_/Y _76223_/Y sky130_fd_sc_hd__nor2_4
X_88209_ _87950_/CLK _41470_/X _66634_/B sky130_fd_sc_hd__dfxtp_4
X_42615_ _42592_/A _42615_/X sky130_fd_sc_hd__buf_2
X_49171_ _49128_/X _48676_/A _49170_/Y _49172_/A sky130_fd_sc_hd__a21o_4
X_73435_ _73433_/X _73434_/Y _73367_/X _73435_/Y sky130_fd_sc_hd__a21oi_4
X_46383_ _46362_/A _52478_/B _46383_/Y sky130_fd_sc_hd__nand2_4
X_70647_ _70717_/A _70639_/B _70642_/X _70638_/X _70647_/Y sky130_fd_sc_hd__nand4_4
X_58369_ _58408_/A _58369_/X sky130_fd_sc_hd__buf_2
X_43595_ _43595_/A _87347_/D sky130_fd_sc_hd__inv_2
Xclkbuf_9_143_0_CLK clkbuf_8_71_0_CLK/X clkbuf_9_143_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_48122_ _83533_/Q _48122_/Y sky130_fd_sc_hd__inv_2
X_60400_ _60395_/X _60400_/Y sky130_fd_sc_hd__inv_2
X_45334_ _64524_/B _61663_/B sky130_fd_sc_hd__buf_2
Xclkbuf_9_70_0_CLK clkbuf_9_71_0_CLK/A clkbuf_9_70_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_76154_ _76151_/Y _76153_/Y _76154_/Y sky130_fd_sc_hd__nor2_4
X_42546_ _42536_/X _42527_/X _40771_/X _69583_/B _42538_/X _87826_/D
+ sky130_fd_sc_hd__o32ai_4
X_61380_ _61380_/A _61391_/D sky130_fd_sc_hd__buf_2
X_73366_ _72765_/A _73367_/A sky130_fd_sc_hd__buf_2
X_70578_ _70578_/A _74515_/C sky130_fd_sc_hd__buf_2
X_75105_ _75105_/A _75105_/Y sky130_fd_sc_hd__inv_2
X_72317_ _72228_/X _85969_/Q _72316_/X _72317_/Y sky130_fd_sc_hd__o21ai_4
X_48053_ _48092_/A _50341_/B _48053_/Y sky130_fd_sc_hd__nand2_4
X_60331_ _60268_/C _60331_/B _60268_/A _60331_/D _60331_/Y sky130_fd_sc_hd__nand4_4
X_45265_ _45265_/A _45265_/X sky130_fd_sc_hd__buf_2
X_76085_ _81721_/D _76085_/B _76097_/B sky130_fd_sc_hd__nand2_4
Xclkbuf_10_667_0_CLK clkbuf_9_333_0_CLK/X _87137_/CLK sky130_fd_sc_hd__clkbuf_1
X_42477_ _42477_/A _42477_/X sky130_fd_sc_hd__buf_2
X_73297_ _42036_/Y _72921_/X _73194_/X _73296_/Y _73297_/X sky130_fd_sc_hd__a211o_4
X_47004_ _47004_/A _47004_/X sky130_fd_sc_hd__buf_2
X_44216_ _43959_/A _44216_/X sky130_fd_sc_hd__buf_2
X_63050_ _63039_/A _84717_/Q _63028_/X _63014_/D _63050_/X sky130_fd_sc_hd__and4_4
X_75036_ _75047_/A _75035_/Y _75036_/X sky130_fd_sc_hd__xor2_4
X_79913_ _79913_/A _79913_/B _79914_/B sky130_fd_sc_hd__nand2_4
X_41428_ _41412_/X _82887_/Q _41427_/X _41428_/Y sky130_fd_sc_hd__o21ai_4
X_60262_ _60211_/A _60263_/C sky130_fd_sc_hd__buf_2
X_72248_ _72172_/X _72245_/Y _72247_/Y _72189_/X _72176_/X _72248_/X
+ sky130_fd_sc_hd__o32a_4
X_45196_ _45196_/A _45199_/A sky130_fd_sc_hd__inv_2
Xclkbuf_9_158_0_CLK clkbuf_8_79_0_CLK/X clkbuf_9_158_0_CLK/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_1_2_CLK clkbuf_2_1_1_CLK/X clkbuf_3_3_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_62001_ _61991_/X _61993_/X _62000_/Y _84848_/Q _61973_/X _62001_/Y
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_9_85_0_CLK clkbuf_8_42_0_CLK/X clkbuf_9_85_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_44147_ _44147_/A _44148_/A sky130_fd_sc_hd__buf_2
X_79844_ _64741_/C _72165_/Y _79843_/Y _79844_/X sky130_fd_sc_hd__o21a_4
X_41359_ _41358_/X _82899_/Q _41359_/X sky130_fd_sc_hd__or2_4
X_72179_ _83276_/Q _72179_/Y sky130_fd_sc_hd__inv_2
X_60193_ _60193_/A _60239_/B sky130_fd_sc_hd__buf_2
X_48955_ _53819_/B _48955_/X sky130_fd_sc_hd__buf_2
X_44078_ _44077_/X _55817_/A sky130_fd_sc_hd__buf_2
X_79775_ _79775_/A _79775_/B _79781_/B sky130_fd_sc_hd__xor2_4
X_76987_ _76987_/A _62426_/C _76987_/X sky130_fd_sc_hd__xor2_4
X_47906_ _82363_/Q _47963_/B _47906_/X sky130_fd_sc_hd__or2_4
X_43029_ _43029_/A _43029_/Y sky130_fd_sc_hd__inv_2
X_66740_ _66737_/X _66739_/X _66667_/X _66743_/A sky130_fd_sc_hd__a21o_4
X_78726_ _78725_/A _78725_/B _78726_/Y sky130_fd_sc_hd__nand2_4
X_63952_ _64045_/A _64016_/D sky130_fd_sc_hd__buf_2
X_75938_ _75939_/B _75938_/Y sky130_fd_sc_hd__inv_2
X_48886_ _48879_/Y _48880_/X _48885_/X _86465_/D sky130_fd_sc_hd__a21oi_4
X_62903_ _62930_/A _62930_/B _84372_/Q _62903_/Y sky130_fd_sc_hd__nor3_4
X_47837_ _47836_/Y _86593_/D sky130_fd_sc_hd__inv_2
X_78657_ _78655_/X _78657_/B _82777_/D sky130_fd_sc_hd__xor2_4
X_66671_ _66668_/X _66670_/X _66671_/Y sky130_fd_sc_hd__nand2_4
X_63883_ _61440_/A _63853_/B _63947_/C _63866_/X _63883_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_10_605_0_CLK clkbuf_9_302_0_CLK/X _82116_/CLK sky130_fd_sc_hd__clkbuf_1
X_75869_ _75868_/X _75875_/B sky130_fd_sc_hd__inv_2
X_68410_ _87102_/Q _68059_/X _68370_/X _68409_/X _68410_/X sky130_fd_sc_hd__a211o_4
X_65622_ _65619_/Y _65602_/X _65621_/X _84189_/D sky130_fd_sc_hd__a21o_4
X_77608_ _77622_/A _77607_/Y _82203_/D sky130_fd_sc_hd__xnor2_4
X_62834_ _61510_/X _62834_/B _62801_/X _62834_/D _62834_/Y sky130_fd_sc_hd__nand4_4
X_69390_ _69386_/X _69388_/X _69389_/X _69390_/Y sky130_fd_sc_hd__a21oi_4
X_47768_ _47768_/A _53234_/D sky130_fd_sc_hd__buf_2
X_78588_ _78584_/Y _78585_/Y _78587_/Y _78588_/X sky130_fd_sc_hd__or3_4
X_49507_ _49503_/Y _49487_/X _49506_/X _86375_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_23_0_CLK clkbuf_9_23_0_CLK/A clkbuf_9_23_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_68341_ _82626_/D _68338_/X _68340_/X _68341_/X sky130_fd_sc_hd__a21bo_4
X_46719_ _46719_/A _46719_/X sky130_fd_sc_hd__buf_2
X_65553_ _65550_/X _65552_/X _65389_/X _65553_/X sky130_fd_sc_hd__a21o_4
X_77539_ _77539_/A _77540_/C sky130_fd_sc_hd__inv_2
X_62765_ _62761_/Y _62713_/X _62762_/Y _62763_/Y _62764_/X _62765_/X
+ sky130_fd_sc_hd__a41o_4
X_47699_ _47792_/A _47739_/B sky130_fd_sc_hd__buf_2
X_64504_ _64457_/B _64229_/X _64504_/C _64503_/Y _64504_/Y sky130_fd_sc_hd__nand4_4
X_49438_ _49418_/A _50961_/B _49438_/Y sky130_fd_sc_hd__nand2_4
X_80550_ _80550_/A _80549_/Y _80562_/B sky130_fd_sc_hd__xor2_4
X_61716_ _59638_/A _61716_/X sky130_fd_sc_hd__buf_2
X_68272_ _68376_/A _68272_/X sky130_fd_sc_hd__buf_2
X_65484_ _65484_/A _65484_/X sky130_fd_sc_hd__buf_2
X_62696_ _62691_/Y _62660_/X _62693_/Y _62694_/Y _62695_/X _62696_/X
+ sky130_fd_sc_hd__a41o_4
X_67223_ _67248_/A _67223_/B _67223_/X sky130_fd_sc_hd__and2_4
X_79209_ _79178_/Y _79192_/B _79189_/Y _79209_/Y sky130_fd_sc_hd__a21oi_4
X_64435_ _64402_/X _64421_/X _84838_/Q _64435_/X sky130_fd_sc_hd__and3_4
X_49369_ _49451_/A _49369_/X sky130_fd_sc_hd__buf_2
X_61647_ _61643_/X _61645_/X _61646_/Y _61647_/Y sky130_fd_sc_hd__a21oi_4
X_80481_ _84763_/Q _80481_/B _80481_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_38_0_CLK clkbuf_9_39_0_CLK/A clkbuf_9_38_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_51400_ _51220_/A _51230_/X _51225_/C _52927_/D _51400_/X sky130_fd_sc_hd__and4_4
X_82220_ _82220_/CLK _82252_/Q _82220_/Q sky130_fd_sc_hd__dfxtp_4
X_67154_ _67131_/A _87675_/Q _67154_/X sky130_fd_sc_hd__and2_4
X_52380_ _85834_/Q _52372_/X _52379_/Y _52380_/Y sky130_fd_sc_hd__o21ai_4
X_64366_ _64344_/X _64379_/B _84828_/Q _64366_/X sky130_fd_sc_hd__and3_4
X_61578_ _61575_/X _61576_/X _61577_/Y _61578_/Y sky130_fd_sc_hd__a21oi_4
X_66105_ _65628_/X _66135_/B _65630_/X _66105_/Y sky130_fd_sc_hd__nand3_4
X_51331_ _51329_/Y _51313_/X _51330_/X _86030_/D sky130_fd_sc_hd__a21oi_4
X_63317_ _63231_/A _63317_/X sky130_fd_sc_hd__buf_2
X_82151_ _82152_/CLK _84143_/Q _82151_/Q sky130_fd_sc_hd__dfxtp_4
X_60529_ _60529_/A _60529_/B _60529_/Y sky130_fd_sc_hd__nor2_4
X_67085_ _66606_/A _67085_/X sky130_fd_sc_hd__buf_2
X_64297_ _59474_/A _64249_/X _64296_/Y _64297_/Y sky130_fd_sc_hd__o21ai_4
X_81102_ _80817_/CLK _79687_/X _81102_/Q sky130_fd_sc_hd__dfxtp_4
X_54050_ _85515_/Q _54035_/X _54049_/Y _54050_/Y sky130_fd_sc_hd__o21ai_4
X_66036_ _65990_/X _86232_/Q _66021_/X _66035_/X _66036_/X sky130_fd_sc_hd__a211o_4
X_51262_ _64745_/B _51259_/X _51261_/Y _51262_/Y sky130_fd_sc_hd__o21ai_4
X_63248_ _63344_/B _60583_/A _60515_/B _63281_/D _60392_/A _63248_/X
+ sky130_fd_sc_hd__o41a_4
X_82082_ _82104_/CLK _82082_/D _82082_/Q sky130_fd_sc_hd__dfxtp_4
X_53001_ _52892_/A _53001_/X sky130_fd_sc_hd__buf_2
X_50213_ _50595_/A _50213_/X sky130_fd_sc_hd__buf_2
X_85910_ _86587_/CLK _85910_/D _73827_/B sky130_fd_sc_hd__dfxtp_4
X_81033_ _82084_/CLK _81033_/D _81033_/Q sky130_fd_sc_hd__dfxtp_4
X_51193_ _51190_/Y _51175_/X _51192_/X _51193_/Y sky130_fd_sc_hd__a21oi_4
X_63179_ _63154_/X _64392_/B _63165_/X _63192_/D _63179_/X sky130_fd_sc_hd__and4_4
X_86890_ _86861_/CLK _45236_/Y _64458_/B sky130_fd_sc_hd__dfxtp_4
X_50144_ _50153_/A _50144_/B _50144_/Y sky130_fd_sc_hd__nand2_4
X_85841_ _85555_/CLK _52346_/Y _65032_/B sky130_fd_sc_hd__dfxtp_4
X_67987_ _67987_/A _67987_/X sky130_fd_sc_hd__buf_2
X_57740_ _57739_/X _85727_/Q _44252_/X _57740_/X sky130_fd_sc_hd__o21a_4
X_69726_ _87059_/Q _69664_/X _69665_/X _69725_/X _69727_/B sky130_fd_sc_hd__a211o_4
X_54952_ _54949_/Y _54936_/X _54951_/X _85347_/D sky130_fd_sc_hd__a21oi_4
X_50075_ _50084_/A _48922_/B _50075_/Y sky130_fd_sc_hd__nand2_4
X_66938_ _66840_/X _66938_/B _66938_/X sky130_fd_sc_hd__and2_4
X_85772_ _85773_/CLK _52695_/Y _85772_/Q sky130_fd_sc_hd__dfxtp_4
X_82984_ _85134_/CLK _82984_/D _82984_/Q sky130_fd_sc_hd__dfxtp_4
X_87511_ _87767_/CLK _87511_/D _87511_/Q sky130_fd_sc_hd__dfxtp_4
X_53903_ _53899_/Y _53862_/X _53902_/Y _85546_/D sky130_fd_sc_hd__a21boi_4
X_84723_ _83464_/CLK _84723_/D _84723_/Q sky130_fd_sc_hd__dfxtp_4
X_57671_ _57650_/X _57668_/Y _57670_/Y _57671_/Y sky130_fd_sc_hd__a21oi_4
X_81935_ _81985_/CLK _77856_/Y _77421_/A sky130_fd_sc_hd__dfxtp_4
X_69657_ _69226_/Y _69644_/X _69604_/X _69656_/Y _69657_/X sky130_fd_sc_hd__a211o_4
X_54883_ _54883_/A _54883_/B _54883_/C _53191_/D _54883_/X sky130_fd_sc_hd__and4_4
X_66869_ _66823_/A _88135_/Q _66869_/X sky130_fd_sc_hd__and2_4
X_59410_ _63161_/A _59411_/A sky130_fd_sc_hd__buf_2
X_56622_ _56621_/X _72664_/C sky130_fd_sc_hd__buf_2
X_68608_ _87094_/Q _68580_/X _68509_/X _68607_/X _68608_/X sky130_fd_sc_hd__a211o_4
X_87442_ _87888_/CLK _87442_/D _87442_/Q sky130_fd_sc_hd__dfxtp_4
X_53834_ _53825_/A _53834_/B _53834_/Y sky130_fd_sc_hd__nand2_4
X_84654_ _84672_/CLK _60140_/Y _60139_/C sky130_fd_sc_hd__dfxtp_4
X_81866_ _84441_/CLK _78057_/X _81866_/Q sky130_fd_sc_hd__dfxtp_4
X_69588_ _69585_/X _69587_/X _69588_/Y sky130_fd_sc_hd__nand2_4
X_59341_ _86661_/Q _59306_/B _59341_/Y sky130_fd_sc_hd__nor2_4
X_83605_ _85837_/CLK _71107_/Y _49082_/A sky130_fd_sc_hd__dfxtp_4
X_56553_ _56552_/Y _56553_/Y sky130_fd_sc_hd__inv_2
X_80817_ _80817_/CLK _83961_/Q _80817_/Q sky130_fd_sc_hd__dfxtp_4
X_68539_ _80827_/D _68462_/X _68538_/X _83971_/D sky130_fd_sc_hd__a21bo_4
X_87373_ _87373_/CLK _87373_/D _87373_/Q sky130_fd_sc_hd__dfxtp_4
X_53765_ _53762_/Y _53747_/X _53764_/X _85573_/D sky130_fd_sc_hd__a21oi_4
X_84585_ _84458_/CLK _84585_/D _78080_/A sky130_fd_sc_hd__dfxtp_4
X_50977_ _86096_/Q _50965_/X _50976_/Y _50977_/Y sky130_fd_sc_hd__o21ai_4
X_81797_ _85381_/CLK _81605_/Q _47493_/A sky130_fd_sc_hd__dfxtp_4
X_55504_ _55447_/Y _55451_/B _55503_/Y _55504_/Y sky130_fd_sc_hd__a21oi_4
X_86324_ _86322_/CLK _49784_/Y _57918_/B sky130_fd_sc_hd__dfxtp_4
X_40730_ _40729_/X _40719_/X _88346_/Q _40720_/X _88346_/D sky130_fd_sc_hd__a2bb2o_4
X_52716_ _52704_/A _52724_/B _52708_/X _52716_/D _52716_/X sky130_fd_sc_hd__and4_4
X_59272_ _59253_/X _59269_/Y _59270_/Y _59271_/X _59258_/X _59272_/X
+ sky130_fd_sc_hd__o32a_4
X_71550_ _70689_/A _71546_/B _71536_/A _71550_/Y sky130_fd_sc_hd__nor3_4
X_83536_ _86210_/CLK _71324_/Y _83536_/Q sky130_fd_sc_hd__dfxtp_4
X_56484_ _56448_/X _56484_/X sky130_fd_sc_hd__buf_2
X_80748_ _81125_/CLK _80748_/D _81124_/D sky130_fd_sc_hd__dfxtp_4
X_53696_ _53696_/A _53696_/X sky130_fd_sc_hd__buf_2
X_70501_ _70500_/Y _70501_/X sky130_fd_sc_hd__buf_2
X_58223_ _58219_/X _58220_/Y _58222_/Y _58223_/Y sky130_fd_sc_hd__a21oi_4
X_55435_ _55431_/Y _55432_/Y _55434_/Y _55435_/X sky130_fd_sc_hd__o21a_4
X_86255_ _86256_/CLK _86255_/D _65084_/B sky130_fd_sc_hd__dfxtp_4
XPHY_501 sky130_fd_sc_hd__decap_3
X_40661_ _40660_/X _40661_/X sky130_fd_sc_hd__buf_2
X_52647_ _52619_/A _52647_/X sky130_fd_sc_hd__buf_2
X_71481_ _71827_/A _71479_/B _70790_/A _71716_/D _71481_/X sky130_fd_sc_hd__and4_4
X_83467_ _85955_/CLK _83467_/D _47808_/A sky130_fd_sc_hd__dfxtp_4
XPHY_512 sky130_fd_sc_hd__decap_3
X_80679_ _80679_/CLK _80679_/D _75138_/A sky130_fd_sc_hd__dfxtp_4
XPHY_523 sky130_fd_sc_hd__decap_3
X_42400_ _42400_/A _87881_/D sky130_fd_sc_hd__inv_2
XPHY_534 sky130_fd_sc_hd__decap_3
X_73220_ _73218_/X _73220_/B _73220_/C _73220_/Y sky130_fd_sc_hd__nand3_4
X_85206_ _85269_/CLK _56406_/Y _85206_/Q sky130_fd_sc_hd__dfxtp_4
X_70432_ _47924_/B _70422_/X _70431_/Y _70432_/Y sky130_fd_sc_hd__o21ai_4
X_58154_ _58154_/A _63033_/A sky130_fd_sc_hd__inv_2
X_82418_ _82820_/CLK _82450_/Q _78547_/A sky130_fd_sc_hd__dfxtp_4
XPHY_545 sky130_fd_sc_hd__decap_3
X_43380_ _43379_/Y _87452_/D sky130_fd_sc_hd__inv_2
X_55366_ _55366_/A _55392_/A sky130_fd_sc_hd__buf_2
X_86186_ _86186_/CLK _50516_/Y _86186_/Q sky130_fd_sc_hd__dfxtp_4
X_40592_ _40591_/X _48903_/A sky130_fd_sc_hd__buf_2
XPHY_556 sky130_fd_sc_hd__decap_3
X_52578_ _85793_/Q _52575_/X _52577_/Y _52578_/Y sky130_fd_sc_hd__o21ai_4
X_83398_ _83431_/CLK _71726_/Y _58229_/A sky130_fd_sc_hd__dfxtp_4
XPHY_567 sky130_fd_sc_hd__decap_3
XPHY_578 sky130_fd_sc_hd__decap_3
X_57105_ _57093_/Y _57105_/Y sky130_fd_sc_hd__inv_2
X_42331_ _42330_/X _42319_/X _41656_/X _87918_/Q _42320_/X _42331_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54317_ _54317_/A _54317_/X sky130_fd_sc_hd__buf_2
XPHY_589 sky130_fd_sc_hd__decap_3
X_73151_ _73148_/X _73150_/X _72862_/X _73156_/A sky130_fd_sc_hd__a21o_4
X_85137_ _85071_/CLK _56697_/X _85137_/Q sky130_fd_sc_hd__dfxtp_4
X_51529_ _51514_/A _53054_/B _51529_/Y sky130_fd_sc_hd__nand2_4
X_70363_ _70362_/X _70364_/A sky130_fd_sc_hd__buf_2
X_58085_ _58703_/A _58085_/X sky130_fd_sc_hd__buf_2
X_82349_ _82349_/CLK _77132_/X _82349_/Q sky130_fd_sc_hd__dfxtp_4
X_55297_ _55297_/A _55297_/X sky130_fd_sc_hd__buf_2
X_72102_ _83284_/Q _72090_/X _72101_/Y _72102_/Y sky130_fd_sc_hd__o21ai_4
X_45050_ _45045_/X _45048_/Y _45049_/X _45050_/Y sky130_fd_sc_hd__a21oi_4
X_57036_ _45752_/Y _56952_/X _57035_/X _85098_/D sky130_fd_sc_hd__o21ai_4
X_54248_ _54244_/Y _54226_/X _54247_/X _54248_/Y sky130_fd_sc_hd__a21oi_4
X_42262_ _42252_/X _42243_/X _41473_/X _87952_/Q _42244_/X _42262_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73082_ _69719_/B _73104_/B _72944_/X _73081_/Y _73082_/X sky130_fd_sc_hd__a211o_4
X_85068_ _84998_/CLK _85068_/D _85068_/Q sky130_fd_sc_hd__dfxtp_4
X_70294_ _70292_/A _70292_/B _83103_/Q _70292_/D _70294_/X sky130_fd_sc_hd__and4_4
X_44001_ _59544_/B _62640_/C sky130_fd_sc_hd__buf_2
X_41213_ _41042_/X _41043_/B _41212_/X _41213_/X sky130_fd_sc_hd__o21a_4
X_72033_ _72009_/A _72033_/X sky130_fd_sc_hd__buf_2
X_76910_ _76910_/A _76885_/X _76910_/C _76899_/Y _76910_/X sky130_fd_sc_hd__and4_4
X_84019_ _84020_/CLK _68179_/X _82059_/D sky130_fd_sc_hd__dfxtp_4
X_42193_ _42162_/A _42193_/X sky130_fd_sc_hd__buf_2
X_54179_ _54184_/A _47372_/Y _54179_/Y sky130_fd_sc_hd__nand2_4
X_77890_ _82244_/Q _77890_/B _77890_/Y sky130_fd_sc_hd__xnor2_4
X_41144_ _40932_/A _41145_/B sky130_fd_sc_hd__buf_2
X_76841_ _76841_/A _76840_/Y _76844_/A sky130_fd_sc_hd__xor2_4
X_58987_ _58987_/A _58987_/Y sky130_fd_sc_hd__inv_2
X_48740_ _48738_/Y _48734_/X _48739_/X _86492_/D sky130_fd_sc_hd__a21oi_4
X_79560_ _79559_/Y _79560_/Y sky130_fd_sc_hd__inv_2
X_57938_ _57875_/X _85394_/Q _57937_/X _57938_/Y sky130_fd_sc_hd__o21ai_4
X_45952_ _45951_/Y _45952_/X sky130_fd_sc_hd__buf_2
X_41075_ _41073_/X _81704_/Q _41074_/X _41076_/A sky130_fd_sc_hd__o21a_4
X_76772_ _81488_/Q _76772_/Y sky130_fd_sc_hd__inv_2
X_73984_ _70117_/D _73939_/X _73983_/X _83128_/D sky130_fd_sc_hd__o21ai_4
X_78511_ _78511_/A _78510_/Y _78511_/X sky130_fd_sc_hd__and2_4
X_44903_ _62195_/A _61298_/B sky130_fd_sc_hd__buf_2
X_87709_ _87708_/CLK _87709_/D _87709_/Q sky130_fd_sc_hd__dfxtp_4
X_75723_ _75723_/A _75723_/B _75724_/B sky130_fd_sc_hd__xor2_4
X_48671_ _48671_/A _48672_/A sky130_fd_sc_hd__inv_2
X_72935_ _72816_/X _65525_/B _72935_/X sky130_fd_sc_hd__and2_4
X_79491_ _79475_/X _79476_/X _79490_/Y _79491_/Y sky130_fd_sc_hd__a21boi_4
X_45883_ _45889_/A _45883_/B _45884_/A sky130_fd_sc_hd__nor2_4
X_57869_ _58080_/A _57971_/A sky130_fd_sc_hd__buf_2
X_47622_ _47622_/A _47623_/A sky130_fd_sc_hd__inv_2
X_59608_ _59608_/A _59689_/B sky130_fd_sc_hd__buf_2
X_78442_ _78429_/Y _78422_/X _78423_/Y _78443_/B sky130_fd_sc_hd__a21boi_4
X_44834_ _44832_/X _44821_/X _41704_/X _67679_/B _44833_/X _44835_/A
+ sky130_fd_sc_hd__o32ai_4
X_75654_ _75659_/B _75653_/Y _75655_/B sky130_fd_sc_hd__xnor2_4
X_60880_ _60879_/Y _60880_/X sky130_fd_sc_hd__buf_2
X_72866_ _72739_/X _72866_/X sky130_fd_sc_hd__buf_2
X_74605_ _46155_/A _74605_/X sky130_fd_sc_hd__buf_2
X_47553_ _47553_/A _53115_/B _47553_/Y sky130_fd_sc_hd__nand2_4
X_71817_ _71813_/A _71435_/C _71049_/A _71817_/X sky130_fd_sc_hd__and3_4
X_59539_ _59539_/A _61078_/B _60593_/A sky130_fd_sc_hd__nor2_4
X_78373_ _78373_/A _82663_/D _78375_/C sky130_fd_sc_hd__nand2_4
X_44765_ _44765_/A _86966_/D sky130_fd_sc_hd__inv_2
X_75585_ _75583_/Y _75584_/Y _75585_/Y sky130_fd_sc_hd__nand2_4
X_41977_ _41965_/X _41975_/X _40753_/X _41976_/Y _41967_/X _88085_/D
+ sky130_fd_sc_hd__o32ai_4
X_72797_ _41986_/Y _72723_/X _72725_/X _72796_/Y _72797_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_591_0_CLK clkbuf_9_295_0_CLK/X _80821_/CLK sky130_fd_sc_hd__clkbuf_1
X_46504_ _46504_/A _49110_/A sky130_fd_sc_hd__inv_2
X_77324_ _77324_/A _82089_/D _77325_/A sky130_fd_sc_hd__nand2_4
X_43716_ _47834_/A _43716_/X sky130_fd_sc_hd__buf_2
X_62550_ _62543_/X _62545_/X _62549_/Y _58465_/A _62511_/X _62550_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74536_ _74614_/A _74600_/A sky130_fd_sc_hd__buf_2
X_40928_ _40817_/X _82274_/Q _40927_/X _40929_/A sky130_fd_sc_hd__o21ai_4
X_47484_ _47530_/A _47513_/A sky130_fd_sc_hd__buf_2
X_71748_ _52936_/B _71737_/X _71747_/Y _83391_/D sky130_fd_sc_hd__o21ai_4
X_44696_ _44686_/X _44687_/X _40645_/Y _44695_/Y _44689_/X _44696_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49223_ _49223_/A _49241_/A sky130_fd_sc_hd__buf_2
X_61501_ _61482_/A _61500_/X _61482_/C _61501_/Y sky130_fd_sc_hd__nand3_4
X_46435_ _86737_/Q _46430_/X _46434_/Y _46435_/Y sky130_fd_sc_hd__o21ai_4
X_77255_ _77250_/A _77253_/Y _77254_/Y _77255_/Y sky130_fd_sc_hd__o21ai_4
X_62481_ _62470_/X _62477_/Y _62480_/X _84847_/Q _62440_/X _62481_/Y
+ sky130_fd_sc_hd__o32ai_4
X_43647_ _40696_/X _43624_/X _87328_/Q _43625_/X _87328_/D sky130_fd_sc_hd__a2bb2o_4
X_74467_ _83060_/Q _74387_/X _74466_/Y _74467_/Y sky130_fd_sc_hd__o21ai_4
X_40859_ _82863_/Q _40883_/B _40859_/X sky130_fd_sc_hd__or2_4
X_71679_ _58480_/Y _71669_/X _71678_/Y _83414_/D sky130_fd_sc_hd__o21ai_4
X_64220_ _64243_/A _64234_/A sky130_fd_sc_hd__buf_2
X_76206_ _76202_/X _76219_/A _76205_/Y _76206_/Y sky130_fd_sc_hd__a21oi_4
X_49154_ _48162_/A _49416_/A sky130_fd_sc_hd__buf_2
X_73418_ _43192_/Y _73298_/X _73251_/X _73417_/Y _73418_/X sky130_fd_sc_hd__a211o_4
X_61432_ _61431_/Y _61432_/Y sky130_fd_sc_hd__inv_2
X_46366_ _46366_/A _46387_/A sky130_fd_sc_hd__buf_2
X_77186_ _82011_/Q _82299_/D _77186_/Y sky130_fd_sc_hd__nand2_4
X_43578_ _40538_/X _53455_/A _87350_/Q _43185_/A _43578_/X sky130_fd_sc_hd__a2bb2o_4
X_74398_ _74408_/A _53651_/B _74398_/Y sky130_fd_sc_hd__nand2_4
X_48105_ _48105_/A _53588_/B sky130_fd_sc_hd__inv_2
X_45317_ _55707_/B _45269_/X _45303_/X _45317_/X sky130_fd_sc_hd__o21a_4
X_64151_ _64162_/A _61656_/A _64173_/C _64151_/X sky130_fd_sc_hd__and3_4
X_76137_ _81728_/D _76144_/B _76143_/B sky130_fd_sc_hd__xor2_4
X_42529_ _42517_/X _42527_/X _40734_/X _42528_/Y _42519_/X _87833_/D
+ sky130_fd_sc_hd__o32ai_4
X_49085_ _86445_/Q _49052_/X _49084_/Y _49085_/Y sky130_fd_sc_hd__o21ai_4
X_61363_ _61361_/X _61349_/X _61362_/Y _61363_/Y sky130_fd_sc_hd__a21oi_4
X_73349_ _88316_/Q _73059_/X _73007_/X _73349_/Y sky130_fd_sc_hd__o21ai_4
X_46297_ _86749_/Q _46292_/X _46296_/Y _46297_/Y sky130_fd_sc_hd__o21ai_4
X_63102_ _60489_/X _63103_/C sky130_fd_sc_hd__buf_2
X_48036_ _48036_/A _48287_/A sky130_fd_sc_hd__buf_2
X_60314_ _59772_/A _59837_/B _79742_/A _60314_/Y sky130_fd_sc_hd__nor3_4
X_45248_ _45202_/X _61590_/B _45219_/X _45248_/Y sky130_fd_sc_hd__o21ai_4
X_76068_ _76068_/A _76067_/Y _76069_/B sky130_fd_sc_hd__xor2_4
X_64082_ _62517_/Y _61030_/A _64081_/Y _64082_/Y sky130_fd_sc_hd__o21ai_4
X_61294_ _60353_/B _61287_/D _60403_/B _61294_/D _72540_/B sky130_fd_sc_hd__nand4_4
Xclkbuf_6_20_0_CLK clkbuf_6_21_0_CLK/A clkbuf_7_41_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_67910_ _86951_/Q _67906_/X _67908_/X _67909_/X _67911_/B sky130_fd_sc_hd__a211o_4
X_75019_ _74999_/X _75008_/X _75021_/B _75019_/X sky130_fd_sc_hd__and3_4
X_63033_ _63033_/A _63004_/B _63004_/C _63033_/D _63033_/X sky130_fd_sc_hd__or4_4
X_60245_ _60232_/Y _60238_/Y _59756_/X _60367_/B _60244_/Y _60245_/Y
+ sky130_fd_sc_hd__a41oi_4
X_45179_ _45175_/Y _45178_/Y _45137_/X _45179_/X sky130_fd_sc_hd__a21o_4
X_68890_ _68887_/X _68889_/X _68748_/X _68890_/X sky130_fd_sc_hd__a21o_4
X_67841_ _87146_/Q _67788_/X _67789_/X _67840_/X _67842_/B sky130_fd_sc_hd__a211o_4
X_79827_ _79825_/X _79834_/B _79827_/Y sky130_fd_sc_hd__xnor2_4
X_60176_ _61286_/B _61316_/A sky130_fd_sc_hd__inv_2
X_49987_ _48171_/X _50001_/A sky130_fd_sc_hd__buf_2
X_48938_ _48938_/A _52291_/A sky130_fd_sc_hd__buf_2
X_79758_ _79740_/X _79743_/Y _79758_/X sky130_fd_sc_hd__or2_4
X_67772_ _87905_/Q _67770_/X _67748_/X _67771_/X _67772_/X sky130_fd_sc_hd__a211o_4
X_64984_ _64904_/A _85843_/Q _64984_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_544_0_CLK clkbuf_9_272_0_CLK/X _81749_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_35_0_CLK clkbuf_6_35_0_CLK/A clkbuf_7_70_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_69511_ _69508_/X _69510_/X _69399_/X _69511_/X sky130_fd_sc_hd__a21o_4
X_66723_ _68721_/A _66819_/A sky130_fd_sc_hd__buf_2
X_78709_ _82813_/Q _78709_/Y sky130_fd_sc_hd__inv_2
X_63935_ _58520_/A _63934_/X _63949_/C _63900_/D _63935_/Y sky130_fd_sc_hd__nand4_4
X_48869_ _86467_/Q _48861_/X _48868_/Y _48869_/Y sky130_fd_sc_hd__o21ai_4
X_79689_ _79679_/X _79681_/B _79688_/Y _79689_/Y sky130_fd_sc_hd__a21boi_4
X_50900_ _50906_/A _51765_/B _50900_/Y sky130_fd_sc_hd__nand2_4
X_81720_ _81412_/CLK _81720_/D _81720_/Q sky130_fd_sc_hd__dfxtp_4
X_69442_ _69442_/A _69442_/X sky130_fd_sc_hd__buf_2
X_66654_ _87440_/Q _66571_/X _66629_/X _66653_/X _66654_/X sky130_fd_sc_hd__a211o_4
X_51880_ _51875_/A _51016_/B _51880_/Y sky130_fd_sc_hd__nand2_4
X_63866_ _64191_/D _63866_/X sky130_fd_sc_hd__buf_2
X_65605_ _65634_/A _65397_/B _65605_/C _65605_/Y sky130_fd_sc_hd__nor3_4
X_50831_ _50828_/Y _50801_/X _50830_/X _86125_/D sky130_fd_sc_hd__a21oi_4
X_62817_ _62815_/X _62779_/X _62816_/Y _62817_/Y sky130_fd_sc_hd__a21oi_4
X_81651_ _81330_/CLK _76656_/B _81651_/Q sky130_fd_sc_hd__dfxtp_4
X_69373_ _87522_/Q _69356_/X _69371_/X _69372_/X _69373_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_559_0_CLK clkbuf_9_279_0_CLK/X _82906_/CLK sky130_fd_sc_hd__clkbuf_1
X_66585_ _66580_/X _66584_/X _66411_/A _66585_/Y sky130_fd_sc_hd__a21oi_4
X_63797_ _61365_/X _63781_/B _63781_/C _63761_/X _63797_/Y sky130_fd_sc_hd__nand4_4
X_80602_ _84774_/Q _84166_/Q _80602_/Y sky130_fd_sc_hd__nand2_4
X_68324_ _68319_/X _67981_/Y _68308_/X _68323_/Y _68324_/X sky130_fd_sc_hd__a211o_4
X_53550_ _53565_/A _50326_/B _53550_/Y sky130_fd_sc_hd__nand2_4
X_65536_ _65484_/X _86202_/Q _65534_/X _65535_/X _65536_/X sky130_fd_sc_hd__a211o_4
X_84370_ _84449_/CLK _84370_/D _62921_/C sky130_fd_sc_hd__dfxtp_4
X_50762_ _86138_/Q _50742_/X _50761_/Y _50762_/Y sky130_fd_sc_hd__o21ai_4
X_62748_ _62746_/X _62721_/X _62747_/Y _84386_/D sky130_fd_sc_hd__a21oi_4
X_81582_ _81582_/CLK _84182_/Q _81582_/Q sky130_fd_sc_hd__dfxtp_4
X_52501_ _52177_/A _52501_/X sky130_fd_sc_hd__buf_2
X_83321_ _83316_/CLK _71941_/Y _83321_/Q sky130_fd_sc_hd__dfxtp_4
X_80533_ _80520_/X _80531_/X _80532_/X _80533_/Y sky130_fd_sc_hd__a21oi_4
X_68255_ _67584_/X _67587_/X _68239_/X _68255_/Y sky130_fd_sc_hd__a21oi_4
X_53481_ _53479_/Y _53455_/X _53480_/Y _85629_/D sky130_fd_sc_hd__a21boi_4
X_65467_ _65463_/Y _65448_/X _65466_/X _84199_/D sky130_fd_sc_hd__a21o_4
X_50693_ _50693_/A _50693_/B _50693_/X sky130_fd_sc_hd__or2_4
X_62679_ _60271_/X _62679_/X sky130_fd_sc_hd__buf_2
X_55220_ _85027_/Q _55152_/A _55128_/A _55219_/X _55220_/X sky130_fd_sc_hd__a211o_4
X_86040_ _86040_/CLK _86040_/D _64860_/B sky130_fd_sc_hd__dfxtp_4
X_67206_ _67183_/A _67206_/B _67206_/X sky130_fd_sc_hd__and2_4
X_52432_ _52436_/A _53949_/B _52432_/Y sky130_fd_sc_hd__nand2_4
X_64418_ _58442_/A _64418_/B _64418_/Y sky130_fd_sc_hd__nor2_4
X_83252_ _85317_/CLK _83252_/D _83252_/Q sky130_fd_sc_hd__dfxtp_4
X_80464_ _80464_/A _63554_/C _80472_/B sky130_fd_sc_hd__xor2_4
X_68186_ _82057_/D _68180_/X _68185_/X _84017_/D sky130_fd_sc_hd__a21bo_4
X_65398_ _65395_/Y _65347_/X _65397_/Y _84203_/D sky130_fd_sc_hd__a21o_4
X_82203_ _82965_/CLK _82203_/D _82395_/D sky130_fd_sc_hd__dfxtp_4
X_55151_ _85098_/Q _44058_/A _55134_/X _55150_/X _55151_/X sky130_fd_sc_hd__a211o_4
X_67137_ _88380_/Q _67110_/X _67040_/X _67136_/X _67137_/X sky130_fd_sc_hd__a211o_4
X_52363_ _65130_/B _52347_/X _52362_/Y _52363_/Y sky130_fd_sc_hd__o21ai_4
X_64349_ _64341_/Y _64348_/X _64328_/X _64349_/X sky130_fd_sc_hd__o21a_4
X_83183_ _83820_/CLK _72707_/X _70251_/C sky130_fd_sc_hd__dfxtp_4
X_80395_ _80386_/Y _80404_/B _80394_/X _80395_/Y sky130_fd_sc_hd__a21boi_4
X_54102_ _53434_/A _54102_/B _54102_/Y sky130_fd_sc_hd__nand2_4
X_51314_ _50802_/A _51266_/B _51330_/C _51314_/X sky130_fd_sc_hd__and3_4
X_82134_ _82009_/CLK _82134_/D _77338_/B sky130_fd_sc_hd__dfxtp_4
X_55082_ _47918_/A _55104_/B sky130_fd_sc_hd__buf_2
X_67068_ _84085_/Q _66971_/X _67067_/X _67068_/X sky130_fd_sc_hd__a21bo_4
X_52294_ _85851_/Q _52269_/X _52293_/Y _52294_/Y sky130_fd_sc_hd__o21ai_4
X_87991_ _87749_/CLK _87991_/D _87991_/Q sky130_fd_sc_hd__dfxtp_4
X_58910_ _86694_/Q _58898_/B _58910_/Y sky130_fd_sc_hd__nor2_4
X_54033_ _53817_/A _54034_/A sky130_fd_sc_hd__buf_2
X_66019_ _60150_/A _66366_/A sky130_fd_sc_hd__buf_2
X_51245_ _64643_/B _51233_/X _51244_/Y _51245_/Y sky130_fd_sc_hd__o21ai_4
X_86942_ _87416_/CLK _86942_/D _67361_/B sky130_fd_sc_hd__dfxtp_4
X_82065_ _80928_/CLK _82065_/D _82065_/Q sky130_fd_sc_hd__dfxtp_4
X_59890_ _59557_/X _59890_/B _59890_/C _60171_/A sky130_fd_sc_hd__nand3_4
X_81016_ _84150_/CLK _84224_/Q _81016_/Q sky130_fd_sc_hd__dfxtp_4
X_58841_ _58837_/Y _58840_/Y _58735_/X _58841_/X sky130_fd_sc_hd__a21o_4
X_51176_ _51149_/A _51192_/B sky130_fd_sc_hd__buf_2
X_86873_ _86873_/CLK _45499_/Y _63079_/B sky130_fd_sc_hd__dfxtp_4
X_50127_ _50125_/Y _50117_/X _50126_/X _50127_/Y sky130_fd_sc_hd__a21oi_4
X_85824_ _85535_/CLK _52433_/Y _85824_/Q sky130_fd_sc_hd__dfxtp_4
X_58772_ _58714_/X _85777_/Q _58716_/X _58772_/X sky130_fd_sc_hd__o21a_4
X_55984_ _55984_/A _74286_/C sky130_fd_sc_hd__buf_2
X_57723_ _46213_/X _57721_/Y _57722_/Y _57700_/X _57703_/X _57723_/X
+ sky130_fd_sc_hd__o32a_4
X_69709_ _43141_/A _69645_/X _68613_/X _69708_/X _69709_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_8_3_0_CLK clkbuf_8_3_0_CLK/A clkbuf_9_7_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_50058_ _48853_/A _50059_/C sky130_fd_sc_hd__buf_2
X_54935_ _85350_/Q _54918_/X _54934_/Y _54935_/Y sky130_fd_sc_hd__o21ai_4
X_85755_ _85754_/CLK _52786_/Y _85755_/Q sky130_fd_sc_hd__dfxtp_4
X_70981_ _70764_/A _70959_/B _70959_/C _71115_/B _70981_/X sky130_fd_sc_hd__and4_4
X_82967_ _82965_/CLK _82967_/D _46715_/A sky130_fd_sc_hd__dfxtp_4
X_41900_ _41887_/X _41888_/X _40617_/X _41899_/Y _41891_/X _41900_/Y
+ sky130_fd_sc_hd__o32ai_4
X_72720_ _72720_/A _73257_/A sky130_fd_sc_hd__buf_2
X_84706_ _84329_/CLK _59738_/Y _80548_/A sky130_fd_sc_hd__dfxtp_4
X_57654_ _57650_/X _57651_/Y _57653_/Y _84961_/D sky130_fd_sc_hd__a21oi_4
X_81918_ _82047_/CLK _77671_/X _81918_/Q sky130_fd_sc_hd__dfxtp_4
X_42880_ _42879_/Y _87671_/D sky130_fd_sc_hd__inv_2
X_54866_ _54919_/A _54885_/A sky130_fd_sc_hd__buf_2
X_85686_ _84787_/CLK _85686_/D _85686_/Q sky130_fd_sc_hd__dfxtp_4
X_82898_ _82327_/CLK _78197_/B _82898_/Q sky130_fd_sc_hd__dfxtp_4
X_56605_ _56600_/X _56553_/Y _56604_/Y _56605_/Y sky130_fd_sc_hd__a21oi_4
X_87425_ _86814_/CLK _87425_/D _87425_/Q sky130_fd_sc_hd__dfxtp_4
X_41831_ _41830_/Y _41831_/Y sky130_fd_sc_hd__inv_2
X_53817_ _53817_/A _53956_/A sky130_fd_sc_hd__buf_2
X_72651_ _83203_/Q _72645_/X _72650_/Y _83203_/D sky130_fd_sc_hd__a21bo_4
X_84637_ _83218_/CLK _84637_/D _79755_/A sky130_fd_sc_hd__dfxtp_4
X_57585_ _84974_/Q _57562_/X _57584_/Y _57585_/Y sky130_fd_sc_hd__o21ai_4
X_81849_ _82515_/CLK _81881_/Q _77568_/A sky130_fd_sc_hd__dfxtp_4
X_54797_ _85376_/Q _54784_/X _54796_/Y _54797_/Y sky130_fd_sc_hd__o21ai_4
X_59324_ _84751_/Q _59268_/X _59318_/X _59323_/X _59324_/Y sky130_fd_sc_hd__a2bb2oi_4
X_71602_ _70410_/Y _70361_/A _71602_/C _71603_/A sky130_fd_sc_hd__nor3_4
X_44550_ _44547_/X _44548_/X _40831_/X _73104_/A _44549_/X _44551_/A
+ sky130_fd_sc_hd__o32ai_4
X_56536_ _56533_/A _56535_/X _56536_/C _56536_/Y sky130_fd_sc_hd__nand3_4
X_75370_ _75370_/A _75369_/Y _75370_/X sky130_fd_sc_hd__xor2_4
X_87356_ _81182_/CLK _43569_/X _87356_/Q sky130_fd_sc_hd__dfxtp_4
X_53748_ _48845_/A _53748_/B _53748_/C _53748_/X sky130_fd_sc_hd__and3_4
X_41762_ _41761_/X _41762_/X sky130_fd_sc_hd__buf_2
X_72582_ _72510_/Y _72546_/Y _72584_/A _72579_/Y _72581_/Y _72582_/Y
+ sky130_fd_sc_hd__a41oi_4
X_84568_ _84583_/CLK _60787_/Y _84568_/Q sky130_fd_sc_hd__dfxtp_4
X_43501_ _41745_/X _43498_/X _87389_/Q _43499_/X _87389_/D sky130_fd_sc_hd__a2bb2o_4
X_74321_ _74325_/A _74325_/B _55863_/X _74321_/Y sky130_fd_sc_hd__nand3_4
X_86307_ _86627_/CLK _86307_/D _58130_/B sky130_fd_sc_hd__dfxtp_4
X_40713_ _40712_/X _40651_/X _88349_/Q _40652_/X _40713_/X sky130_fd_sc_hd__a2bb2o_4
X_71533_ _71602_/C _71585_/A sky130_fd_sc_hd__buf_2
X_59255_ _59255_/A _59256_/A sky130_fd_sc_hd__buf_2
X_83519_ _83521_/CLK _71382_/X _83519_/Q sky130_fd_sc_hd__dfxtp_4
X_44481_ _44547_/A _44481_/X sky130_fd_sc_hd__buf_2
X_56467_ _56463_/A _56538_/A sky130_fd_sc_hd__buf_2
X_41693_ _41692_/Y _41693_/X sky130_fd_sc_hd__buf_2
X_87287_ _87577_/CLK _87287_/D _43744_/A sky130_fd_sc_hd__dfxtp_4
X_53679_ _85589_/Q _53660_/X _53678_/Y _53679_/Y sky130_fd_sc_hd__o21ai_4
X_84499_ _84493_/CLK _84499_/D _75901_/A sky130_fd_sc_hd__dfxtp_4
X_46220_ _46220_/A _46220_/Y sky130_fd_sc_hd__inv_2
XPHY_320 sky130_fd_sc_hd__decap_3
X_58206_ _57665_/A _58238_/B sky130_fd_sc_hd__buf_2
X_77040_ _77041_/A _77041_/C _77041_/B _77047_/A sky130_fd_sc_hd__a21o_4
X_43432_ _43397_/A _43432_/X sky130_fd_sc_hd__buf_2
X_55418_ _55416_/Y _55296_/B _55417_/Y _56807_/A sky130_fd_sc_hd__a21o_4
X_74252_ _74012_/X _86211_/Q _45930_/X _74251_/X _74252_/X sky130_fd_sc_hd__a211o_4
X_86238_ _86238_/CLK _86238_/D _86238_/Q sky130_fd_sc_hd__dfxtp_4
X_40644_ _40644_/A _40588_/B _40644_/X sky130_fd_sc_hd__or2_4
XPHY_331 sky130_fd_sc_hd__decap_3
X_59186_ _59085_/X _86066_/Q _59185_/X _59186_/Y sky130_fd_sc_hd__o21ai_4
X_71464_ _71463_/Y _71464_/X sky130_fd_sc_hd__buf_2
X_56398_ _56436_/A _56399_/B sky130_fd_sc_hd__buf_2
XPHY_342 sky130_fd_sc_hd__decap_3
XPHY_353 sky130_fd_sc_hd__decap_3
XPHY_364 sky130_fd_sc_hd__decap_3
X_73203_ _88322_/Q _73086_/X _73202_/X _73203_/X sky130_fd_sc_hd__o21a_4
X_46151_ _46101_/A _46151_/B _46108_/D _46166_/C sky130_fd_sc_hd__and3_4
X_58137_ _58079_/X _58135_/Y _58136_/Y _58098_/X _58083_/X _58137_/X
+ sky130_fd_sc_hd__o32a_4
X_70415_ _70412_/X _70694_/A _70700_/B _70428_/A sky130_fd_sc_hd__nand3_4
XPHY_375 sky130_fd_sc_hd__decap_3
X_55349_ _55323_/A _85137_/Q _55349_/X sky130_fd_sc_hd__and2_4
X_43363_ _43347_/X _43350_/X _41376_/X _87458_/Q _43353_/X _43364_/A
+ sky130_fd_sc_hd__o32ai_4
X_74183_ _70129_/A _74139_/X _74182_/Y _74183_/X sky130_fd_sc_hd__a21o_4
X_86169_ _85562_/CLK _86169_/D _86169_/Q sky130_fd_sc_hd__dfxtp_4
X_40575_ _40574_/Y _40575_/Y sky130_fd_sc_hd__inv_2
XPHY_386 sky130_fd_sc_hd__decap_3
X_71395_ _71191_/A _71342_/B _71395_/Y sky130_fd_sc_hd__nor2_4
XPHY_397 sky130_fd_sc_hd__decap_3
X_45102_ _45827_/B _45102_/X sky130_fd_sc_hd__buf_2
X_42314_ _42314_/A _42314_/Y sky130_fd_sc_hd__inv_2
X_73134_ _73306_/A _73260_/A sky130_fd_sc_hd__buf_2
X_46082_ _46082_/A _46082_/Y sky130_fd_sc_hd__inv_2
X_58068_ _58064_/Y _58067_/Y _58035_/X _58068_/X sky130_fd_sc_hd__a21o_4
X_70346_ _70348_/A _70348_/B _70346_/C _70348_/D _70346_/X sky130_fd_sc_hd__and4_4
X_43294_ _41189_/X _43287_/X _87493_/Q _43288_/X _43294_/X sky130_fd_sc_hd__a2bb2o_4
X_78991_ _82645_/Q _82517_/D _78990_/X _78991_/Y sky130_fd_sc_hd__o21ai_4
X_49910_ _49904_/A _49893_/B _49904_/C _53125_/D _49910_/X sky130_fd_sc_hd__and4_4
X_45033_ _74564_/C _45033_/B _45033_/Y sky130_fd_sc_hd__nand2_4
X_57019_ _57019_/A _57011_/Y _57019_/C _57019_/X sky130_fd_sc_hd__and3_4
X_42245_ _42231_/X _42243_/X _41424_/X _87962_/Q _42244_/X _42245_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73065_ _73093_/A _86486_/Q _73065_/X sky130_fd_sc_hd__and2_4
X_77942_ _77942_/A _77942_/B _77942_/X sky130_fd_sc_hd__xor2_4
X_70277_ _70267_/A _70267_/B _70277_/C _70264_/X _70277_/X sky130_fd_sc_hd__and4_4
X_60030_ _60079_/B _59922_/C _60091_/A _60091_/C _60030_/Y sky130_fd_sc_hd__nand4_4
X_72016_ _71985_/A _72016_/X sky130_fd_sc_hd__buf_2
X_49841_ _49827_/X _53054_/B _49841_/Y sky130_fd_sc_hd__nand2_4
X_42176_ _41230_/X _42161_/X _87997_/Q _42162_/X _42176_/X sky130_fd_sc_hd__a2bb2o_4
X_77873_ _77885_/A _77872_/Y _77880_/A sky130_fd_sc_hd__xor2_4
X_79612_ _79596_/Y _79592_/Y _79594_/Y _79612_/Y sky130_fd_sc_hd__a21boi_4
X_41127_ _41127_/A _41127_/Y sky130_fd_sc_hd__inv_2
X_76824_ _76812_/A _76811_/Y _76823_/X _76824_/Y sky130_fd_sc_hd__o21ai_4
X_49772_ _49779_/A _49750_/X _49789_/C _52989_/D _49772_/X sky130_fd_sc_hd__and4_4
X_46984_ _54478_/B _52787_/B sky130_fd_sc_hd__buf_2
X_48723_ _48388_/A _48099_/X _48723_/C _48723_/X sky130_fd_sc_hd__and3_4
X_79543_ _79543_/A _79542_/Y _79543_/Y sky130_fd_sc_hd__nor2_4
X_45935_ _45935_/A _45935_/X sky130_fd_sc_hd__buf_2
X_41058_ _41024_/X _41228_/A _41057_/X _41058_/Y sky130_fd_sc_hd__o21ai_4
X_76755_ _76755_/A _76755_/B _76755_/Y sky130_fd_sc_hd__xnor2_4
X_61981_ _59807_/A _61981_/X sky130_fd_sc_hd__buf_2
X_73967_ _73964_/X _73966_/X _73944_/X _73967_/X sky130_fd_sc_hd__a21o_4
X_63720_ _60920_/A _63721_/C sky130_fd_sc_hd__buf_2
X_75706_ _80913_/Q _75708_/A sky130_fd_sc_hd__inv_2
X_72918_ _72904_/Y _72917_/X _72918_/Y sky130_fd_sc_hd__xnor2_4
X_48654_ _48654_/A _48632_/B _48654_/Y sky130_fd_sc_hd__nand2_4
X_60932_ _60707_/X _60913_/Y _60988_/A _60962_/A _60931_/Y _60932_/Y
+ sky130_fd_sc_hd__a41oi_4
X_79474_ _79466_/X _79468_/B _79473_/Y _79474_/Y sky130_fd_sc_hd__a21boi_4
X_45866_ _45859_/X _45863_/Y _45865_/Y _45866_/Y sky130_fd_sc_hd__a21oi_4
X_76686_ _76686_/A _76969_/A _76686_/Y sky130_fd_sc_hd__nor2_4
X_73898_ _72861_/X _73898_/X sky130_fd_sc_hd__buf_2
X_47605_ _81241_/Q _55005_/D sky130_fd_sc_hd__inv_2
X_78425_ _78369_/A _78397_/B _78400_/A _78413_/Y _78425_/Y sky130_fd_sc_hd__nand4_4
X_44817_ _43927_/X _44817_/X sky130_fd_sc_hd__buf_2
X_63651_ _62094_/D _60780_/X _63357_/X _60767_/X _63650_/Y _63651_/X
+ sky130_fd_sc_hd__a2111o_4
X_75637_ _75637_/A _80826_/Q _75637_/Y sky130_fd_sc_hd__xnor2_4
X_48585_ _48651_/A _48585_/X sky130_fd_sc_hd__buf_2
X_60863_ _60863_/A _60863_/X sky130_fd_sc_hd__buf_2
X_72849_ _72847_/X _72848_/Y _72766_/X _72849_/Y sky130_fd_sc_hd__a21oi_4
X_45797_ _45794_/X _45796_/Y _45757_/X _45797_/X sky130_fd_sc_hd__a21o_4
X_62602_ _61663_/B _62548_/C _62507_/X _62548_/B _62601_/X _62602_/X
+ sky130_fd_sc_hd__a41o_4
X_47536_ _47536_/A _53105_/B sky130_fd_sc_hd__buf_2
X_66370_ _66368_/Y _66343_/X _66369_/X _84136_/D sky130_fd_sc_hd__a21o_4
X_78356_ _78356_/A _78356_/B _82469_/D sky130_fd_sc_hd__xnor2_4
X_44748_ _49210_/A _50731_/B _40753_/A _44747_/Y _44736_/X _86977_/D
+ sky130_fd_sc_hd__o32ai_4
X_75568_ _75568_/A _75570_/A sky130_fd_sc_hd__inv_2
X_63582_ _63546_/A _58478_/A _63581_/X _63546_/D _63582_/X sky130_fd_sc_hd__and4_4
X_60794_ _60736_/X _60711_/X _60725_/A _60697_/B _60528_/A _60794_/Y
+ sky130_fd_sc_hd__a41oi_4
X_65321_ _65317_/X _66423_/B _65320_/X _65321_/Y sky130_fd_sc_hd__nand3_4
X_77307_ _77307_/A _77307_/Y sky130_fd_sc_hd__inv_2
X_74519_ _52794_/B _74517_/X _74518_/Y _74519_/Y sky130_fd_sc_hd__o21ai_4
X_62533_ _62533_/A _58495_/A _62532_/X _62536_/C sky130_fd_sc_hd__nand3_4
X_47467_ _47461_/Y _47462_/X _47466_/X _47467_/Y sky130_fd_sc_hd__a21oi_4
X_78287_ _82686_/Q _78287_/B _78287_/X sky130_fd_sc_hd__xor2_4
X_44679_ _44679_/A _44679_/X sky130_fd_sc_hd__buf_2
X_75499_ _75495_/Y _75497_/Y _75498_/A _75503_/C sky130_fd_sc_hd__o21ai_4
X_49206_ _46242_/Y _51235_/B sky130_fd_sc_hd__buf_2
X_68040_ _68120_/A _68040_/X sky130_fd_sc_hd__buf_2
X_46418_ _46413_/Y _46399_/X _46417_/Y _46418_/Y sky130_fd_sc_hd__a21boi_4
X_65252_ _64797_/A _65252_/X sky130_fd_sc_hd__buf_2
X_77238_ _77239_/A _77239_/C _77239_/B _77245_/A sky130_fd_sc_hd__a21o_4
X_62464_ _62479_/A _61997_/X _62479_/C _62463_/X _62464_/X sky130_fd_sc_hd__and4_4
X_47398_ _81807_/Q _47399_/A sky130_fd_sc_hd__inv_2
X_64203_ _59716_/A _64203_/B _72625_/A _64421_/A _64440_/A sky130_fd_sc_hd__nand4_4
X_61415_ _61434_/A _61434_/B _79151_/B _61415_/Y sky130_fd_sc_hd__nor3_4
X_49137_ _65253_/B _49104_/X _49136_/Y _49137_/Y sky130_fd_sc_hd__o21ai_4
X_46349_ _46349_/A _46380_/B sky130_fd_sc_hd__buf_2
X_65183_ _64903_/A _65184_/A sky130_fd_sc_hd__buf_2
X_77169_ _77170_/A _77170_/B _77172_/A sky130_fd_sc_hd__nor2_4
X_62395_ _61348_/A _62395_/X sky130_fd_sc_hd__buf_2
X_64134_ _62577_/Y _60879_/Y _62124_/B _61028_/X _64134_/Y sky130_fd_sc_hd__a2bb2oi_4
X_49068_ _48606_/X _81199_/Q _49067_/Y _49069_/A sky130_fd_sc_hd__o21ai_4
X_61346_ _61329_/Y _61332_/Y _61334_/X _61338_/Y _61345_/Y _61346_/X
+ sky130_fd_sc_hd__a41o_4
X_80180_ _80164_/Y _80167_/Y _80179_/X _80180_/X sky130_fd_sc_hd__a21o_4
X_69991_ _82558_/D _69988_/X _69990_/X _83878_/D sky130_fd_sc_hd__a21bo_4
X_48019_ _47971_/X _82928_/Q _48018_/X _48020_/B sky130_fd_sc_hd__o21ai_4
X_68942_ _87996_/Q _68895_/X _68916_/X _68941_/X _68942_/X sky130_fd_sc_hd__a211o_4
X_64065_ _60909_/X _64095_/C sky130_fd_sc_hd__buf_2
X_61277_ _59545_/A _61277_/B _61277_/C _61281_/C sky130_fd_sc_hd__nor3_4
X_51030_ _51027_/Y _51011_/X _51029_/X _51030_/Y sky130_fd_sc_hd__a21oi_4
X_63016_ _63342_/C _63030_/C sky130_fd_sc_hd__buf_2
X_60228_ _60228_/A _60331_/D sky130_fd_sc_hd__buf_2
X_68873_ _87487_/Q _68870_/X _68871_/X _68872_/X _68873_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_483_0_CLK clkbuf_9_241_0_CLK/X _85962_/CLK sky130_fd_sc_hd__clkbuf_1
X_67824_ _67819_/X _67823_/X _67799_/X _67824_/X sky130_fd_sc_hd__a21o_4
X_60159_ _60159_/A _60263_/A sky130_fd_sc_hd__buf_2
X_83870_ _82369_/CLK _83870_/D _82550_/D sky130_fd_sc_hd__dfxtp_4
X_82821_ _82822_/CLK _82821_/D _82821_/Q sky130_fd_sc_hd__dfxtp_4
X_67755_ _68370_/A _67755_/X sky130_fd_sc_hd__buf_2
X_52981_ _53062_/A _52997_/C sky130_fd_sc_hd__buf_2
X_64967_ _64961_/A _64967_/X sky130_fd_sc_hd__buf_2
X_54720_ _54693_/X _54720_/X sky130_fd_sc_hd__buf_2
X_66706_ _66410_/A _66706_/X sky130_fd_sc_hd__buf_2
X_85540_ _86149_/CLK _53931_/Y _85540_/Q sky130_fd_sc_hd__dfxtp_4
X_51932_ _53259_/A _50224_/B _51932_/Y sky130_fd_sc_hd__nand2_4
X_63918_ _63496_/B _63900_/B _63949_/C _63900_/D _63922_/B sky130_fd_sc_hd__nand4_4
X_82752_ _81019_/CLK _84136_/Q _82752_/Q sky130_fd_sc_hd__dfxtp_4
X_67686_ _67664_/X _67674_/Y _67624_/X _67685_/Y _67686_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_498_0_CLK clkbuf_9_249_0_CLK/X _86711_/CLK sky130_fd_sc_hd__clkbuf_1
X_64898_ _64898_/A _65319_/A sky130_fd_sc_hd__buf_2
X_81703_ _81703_/CLK _75957_/A _81703_/Q sky130_fd_sc_hd__dfxtp_4
X_69425_ _69302_/A _87774_/Q _69425_/X sky130_fd_sc_hd__and2_4
X_54651_ _85403_/Q _54648_/X _54650_/Y _54651_/Y sky130_fd_sc_hd__o21ai_4
X_66637_ _66499_/B _66623_/Y _59782_/X _66636_/Y _66637_/X sky130_fd_sc_hd__a211o_4
X_85471_ _85471_/CLK _54280_/Y _85471_/Q sky130_fd_sc_hd__dfxtp_4
X_51863_ _85932_/Q _51846_/X _51862_/Y _51863_/Y sky130_fd_sc_hd__o21ai_4
X_63849_ _63849_/A _63849_/X sky130_fd_sc_hd__buf_2
X_82683_ _82931_/CLK _78680_/B _82683_/Q sky130_fd_sc_hd__dfxtp_4
X_87210_ _87210_/CLK _87210_/D _87210_/Q sky130_fd_sc_hd__dfxtp_4
X_53602_ _85604_/Q _53586_/X _53601_/Y _53602_/Y sky130_fd_sc_hd__o21ai_4
X_84422_ _84538_/CLK _84422_/D _76998_/B sky130_fd_sc_hd__dfxtp_4
X_50814_ _50806_/A _51324_/B _50814_/Y sky130_fd_sc_hd__nand2_4
X_57370_ _57236_/X _57083_/X _57369_/Y _57370_/X sky130_fd_sc_hd__o21a_4
X_81634_ _83914_/CLK _81666_/Q _81634_/Q sky130_fd_sc_hd__dfxtp_4
X_69356_ _69607_/A _69356_/X sky130_fd_sc_hd__buf_2
X_88190_ _87116_/CLK _88190_/D _67087_/B sky130_fd_sc_hd__dfxtp_4
X_54582_ _54578_/A _47165_/Y _54582_/Y sky130_fd_sc_hd__nand2_4
X_66568_ _87891_/Q _66562_/X _66564_/X _66567_/X _66568_/X sky130_fd_sc_hd__a211o_4
X_51794_ _51794_/A _51794_/B _51794_/C _52622_/D _51794_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_421_0_CLK clkbuf_9_210_0_CLK/X _83507_/CLK sky130_fd_sc_hd__clkbuf_1
X_56321_ _56350_/A _56321_/X sky130_fd_sc_hd__buf_2
X_68307_ _82635_/D _68299_/X _68306_/X _68307_/X sky130_fd_sc_hd__a21bo_4
X_87141_ _87141_/CLK _87141_/D _87141_/Q sky130_fd_sc_hd__dfxtp_4
X_53533_ _50308_/A _53474_/B _53492_/X _53533_/X sky130_fd_sc_hd__and3_4
X_65519_ _65777_/A _65519_/B _65519_/X sky130_fd_sc_hd__and2_4
X_84353_ _83227_/CLK _63105_/X _79427_/A sky130_fd_sc_hd__dfxtp_4
X_50745_ _86142_/Q _50742_/X _50744_/Y _50745_/Y sky130_fd_sc_hd__o21ai_4
X_81565_ _84064_/CLK _76905_/Y _76366_/B sky130_fd_sc_hd__dfxtp_4
X_69287_ _88040_/Q _69217_/X _69245_/X _69286_/X _69287_/X sky130_fd_sc_hd__a211o_4
X_66499_ _66287_/X _66499_/B _66289_/X _66499_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_4_13_1_CLK clkbuf_4_13_0_CLK/X clkbuf_5_27_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_59040_ _59035_/Y _59039_/Y _58966_/X _59040_/X sky130_fd_sc_hd__a21o_4
X_83304_ _83304_/CLK _72006_/Y _83304_/Q sky130_fd_sc_hd__dfxtp_4
X_56252_ _56252_/A _56263_/A sky130_fd_sc_hd__buf_2
X_80516_ _84767_/Q _84159_/Q _80518_/A sky130_fd_sc_hd__xor2_4
X_68238_ _68160_/A _68238_/X sky130_fd_sc_hd__buf_2
X_87072_ _87077_/CLK _87072_/D _87072_/Q sky130_fd_sc_hd__dfxtp_4
X_53464_ _53817_/A _53990_/A sky130_fd_sc_hd__buf_2
X_84284_ _84668_/CLK _84284_/D _80111_/B sky130_fd_sc_hd__dfxtp_4
X_50676_ _50551_/A _50676_/X sky130_fd_sc_hd__buf_2
X_81496_ _82648_/CLK _84064_/Q _81496_/Q sky130_fd_sc_hd__dfxtp_4
X_55203_ _57071_/B _55157_/X _55165_/X _55202_/Y _55203_/X sky130_fd_sc_hd__a211o_4
X_86023_ _86118_/CLK _51373_/Y _65275_/B sky130_fd_sc_hd__dfxtp_4
X_52415_ _52496_/A _52415_/X sky130_fd_sc_hd__buf_2
X_83235_ _84487_/CLK _83235_/D _79447_/B sky130_fd_sc_hd__dfxtp_4
X_80447_ _80448_/B _80448_/A _80447_/X sky130_fd_sc_hd__or2_4
X_56183_ _56182_/X _56183_/X sky130_fd_sc_hd__buf_2
X_68169_ _68106_/A _68169_/X sky130_fd_sc_hd__buf_2
X_53395_ _53386_/A _53395_/B _53395_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_436_0_CLK clkbuf_9_218_0_CLK/X _81233_/CLK sky130_fd_sc_hd__clkbuf_1
X_70200_ _70200_/A _70200_/B _83199_/Q _70200_/D _70200_/X sky130_fd_sc_hd__and4_4
X_55134_ _55133_/X _55134_/X sky130_fd_sc_hd__buf_2
X_40360_ _44528_/A _57491_/A sky130_fd_sc_hd__buf_2
X_52346_ _52344_/Y _52340_/X _52345_/X _52346_/Y sky130_fd_sc_hd__a21oi_4
X_71180_ _70611_/X _74518_/D sky130_fd_sc_hd__buf_2
X_83166_ _83167_/CLK _73077_/X _83166_/Q sky130_fd_sc_hd__dfxtp_4
X_80378_ _84754_/Q _66247_/C _80378_/X sky130_fd_sc_hd__xor2_4
X_70131_ _70131_/A _70131_/B _70131_/C _70131_/X sky130_fd_sc_hd__and3_4
X_82117_ _82145_/CLK _77761_/X _82105_/D sky130_fd_sc_hd__dfxtp_4
X_59942_ _59923_/Y _62534_/A sky130_fd_sc_hd__buf_2
X_55065_ _55043_/X _55056_/X _55070_/C _47722_/A _55065_/X sky130_fd_sc_hd__and4_4
X_52277_ _52293_/A _48912_/B _52277_/Y sky130_fd_sc_hd__nand2_4
X_87974_ _87149_/CLK _87974_/D _87974_/Q sky130_fd_sc_hd__dfxtp_4
X_83097_ _83095_/CLK _83097_/D _70313_/C sky130_fd_sc_hd__dfxtp_4
X_42030_ _42029_/Y _88065_/D sky130_fd_sc_hd__inv_2
X_54016_ _46427_/A _53964_/B _53969_/C _54016_/X sky130_fd_sc_hd__and3_4
X_51228_ _86050_/Q _51209_/X _51227_/Y _51228_/Y sky130_fd_sc_hd__o21ai_4
X_86925_ _87652_/CLK _44842_/X _67773_/B sky130_fd_sc_hd__dfxtp_4
X_82048_ _82047_/CLK _78017_/X _82016_/D sky130_fd_sc_hd__dfxtp_4
X_70062_ _82540_/D _70048_/X _70061_/X _70062_/X sky130_fd_sc_hd__a21bo_4
X_59873_ _59873_/A _59873_/B _80266_/B _59873_/Y sky130_fd_sc_hd__nor3_4
X_58824_ _58787_/X _86093_/Q _58823_/X _58824_/Y sky130_fd_sc_hd__o21ai_4
X_51159_ _86063_/Q _51156_/X _51158_/Y _51159_/Y sky130_fd_sc_hd__o21ai_4
X_74870_ _81125_/D _74870_/B _74870_/Y sky130_fd_sc_hd__nor2_4
X_86856_ _86855_/CLK _45767_/Y _62083_/D sky130_fd_sc_hd__dfxtp_4
X_73821_ _41922_/Y _56182_/X _73819_/X _73820_/Y _73821_/X sky130_fd_sc_hd__a211o_4
X_85807_ _86127_/CLK _52514_/Y _65074_/B sky130_fd_sc_hd__dfxtp_4
X_58755_ _84802_/Q _58755_/Y sky130_fd_sc_hd__inv_2
X_43981_ _59899_/B _59899_/D _59538_/C sky130_fd_sc_hd__and2_4
X_55967_ _55695_/A _85247_/Q _55967_/X sky130_fd_sc_hd__and2_4
X_86787_ _86784_/CLK _46063_/X _86787_/Q sky130_fd_sc_hd__dfxtp_4
X_83999_ _81755_/CLK _83999_/D _83999_/Q sky130_fd_sc_hd__dfxtp_4
X_45720_ _45720_/A _45720_/X sky130_fd_sc_hd__buf_2
X_57706_ _57705_/X _85505_/Q _44031_/X _57706_/X sky130_fd_sc_hd__o21a_4
X_76540_ _76535_/X _76540_/B _76540_/C _76541_/B sky130_fd_sc_hd__nand3_4
X_42932_ _41745_/X _42930_/X _87645_/Q _42931_/X _42932_/X sky130_fd_sc_hd__a2bb2o_4
X_54918_ _53448_/X _54918_/X sky130_fd_sc_hd__buf_2
X_73752_ _73752_/A _73701_/B _73752_/Y sky130_fd_sc_hd__nor2_4
X_85738_ _85738_/CLK _52880_/Y _85738_/Q sky130_fd_sc_hd__dfxtp_4
X_70964_ _70969_/A _70942_/B _70962_/C _70964_/Y sky130_fd_sc_hd__nand3_4
X_58686_ _84808_/Q _58599_/X _58678_/X _58685_/X _84808_/D sky130_fd_sc_hd__a2bb2oi_4
X_55898_ _55895_/X _55897_/X _44118_/B _55902_/A sky130_fd_sc_hd__a21o_4
X_72703_ _45891_/X _72704_/A sky130_fd_sc_hd__buf_2
X_45651_ _45651_/A _45651_/X sky130_fd_sc_hd__buf_2
X_57637_ _71972_/A _57637_/B _57637_/Y sky130_fd_sc_hd__nand2_4
X_76471_ _81272_/Q _81528_/D _76471_/Y sky130_fd_sc_hd__nor2_4
X_54849_ _54846_/Y _54830_/X _54848_/X _54849_/Y sky130_fd_sc_hd__a21oi_4
X_42863_ _41560_/X _42852_/X _67033_/B _42853_/X _42863_/X sky130_fd_sc_hd__a2bb2o_4
X_73683_ _73948_/A _73683_/X sky130_fd_sc_hd__buf_2
X_85669_ _84815_/CLK _85669_/D _85669_/Q sky130_fd_sc_hd__dfxtp_4
X_70895_ _70866_/A _70903_/B sky130_fd_sc_hd__buf_2
X_78210_ _78220_/A _78210_/B _78211_/B sky130_fd_sc_hd__xor2_4
X_44602_ _44602_/A _44602_/X sky130_fd_sc_hd__buf_2
X_75422_ _80793_/Q _75421_/X _80761_/D sky130_fd_sc_hd__xor2_4
X_87408_ _87408_/CLK _87408_/D _87408_/Q sky130_fd_sc_hd__dfxtp_4
X_41814_ _41814_/A _41814_/X sky130_fd_sc_hd__buf_2
X_48370_ _65444_/B _48350_/X _48369_/Y _48370_/Y sky130_fd_sc_hd__o21ai_4
X_72634_ _44231_/A _72643_/B sky130_fd_sc_hd__buf_2
X_79190_ _79189_/Y _79190_/Y sky130_fd_sc_hd__inv_2
X_45582_ _45582_/A _45597_/B _45582_/Y sky130_fd_sc_hd__nor2_4
X_57568_ _57566_/Y _57506_/X _57567_/X _84978_/D sky130_fd_sc_hd__a21oi_4
X_42794_ _42794_/A _87714_/D sky130_fd_sc_hd__inv_2
X_88388_ _88394_/CLK _40461_/Y _88388_/Q sky130_fd_sc_hd__dfxtp_4
X_47321_ _47330_/A _47349_/B _47321_/C _52982_/D _47321_/X sky130_fd_sc_hd__and4_4
X_59307_ _59253_/X _59304_/Y _59306_/Y _59271_/X _59258_/X _59307_/X
+ sky130_fd_sc_hd__o32a_4
X_78141_ _82570_/Q _82858_/D _78141_/Y sky130_fd_sc_hd__nand2_4
X_44533_ _44533_/A _44533_/X sky130_fd_sc_hd__buf_2
X_56519_ _56114_/X _56515_/X _56518_/Y _85165_/D sky130_fd_sc_hd__o21ai_4
X_75353_ _75349_/Y _75351_/Y _75348_/Y _75353_/Y sky130_fd_sc_hd__o21ai_4
X_41745_ _41744_/Y _41745_/X sky130_fd_sc_hd__buf_2
X_87339_ _87070_/CLK _43619_/X _73752_/A sky130_fd_sc_hd__dfxtp_4
X_72565_ _72573_/A _72573_/B _79427_/B _72565_/Y sky130_fd_sc_hd__nor3_4
X_57499_ _57499_/A _47853_/Y _57499_/Y sky130_fd_sc_hd__nand2_4
X_74304_ _74302_/X _74310_/B _55927_/X _74304_/Y sky130_fd_sc_hd__nand3_4
X_59238_ _59238_/A _59238_/X sky130_fd_sc_hd__buf_2
X_71516_ _53236_/B _71508_/X _71515_/Y _83471_/D sky130_fd_sc_hd__o21ai_4
X_47252_ _54106_/B _52940_/B sky130_fd_sc_hd__buf_2
X_78072_ _60744_/C _78072_/B _78072_/X sky130_fd_sc_hd__xor2_4
X_44464_ _44602_/A _44464_/X sky130_fd_sc_hd__buf_2
X_75284_ _75284_/A _75283_/Y _75284_/X sky130_fd_sc_hd__xor2_4
X_41676_ _41675_/X _41676_/X sky130_fd_sc_hd__buf_2
X_72496_ _64454_/A _72498_/B _72496_/Y sky130_fd_sc_hd__nand2_4
X_46203_ _58273_/A _58160_/B sky130_fd_sc_hd__buf_2
XPHY_150 sky130_fd_sc_hd__decap_3
X_77023_ _77023_/A _77023_/B _77034_/B sky130_fd_sc_hd__xor2_4
X_43415_ _43399_/X _43404_/X _41515_/X _87432_/Q _43407_/X _43416_/A
+ sky130_fd_sc_hd__o32ai_4
X_74235_ _44270_/X _85604_/Q _44272_/X _74234_/X _74235_/X sky130_fd_sc_hd__a211o_4
XPHY_161 sky130_fd_sc_hd__decap_3
X_40627_ _40626_/X _40596_/X _88364_/Q _40599_/X _88364_/D sky130_fd_sc_hd__a2bb2o_4
X_47183_ _47183_/A _47184_/A sky130_fd_sc_hd__inv_2
X_59169_ _58766_/A _59169_/X sky130_fd_sc_hd__buf_2
X_71447_ _71446_/X _71626_/C sky130_fd_sc_hd__buf_2
X_44395_ _44454_/A _44395_/X sky130_fd_sc_hd__buf_2
XPHY_172 sky130_fd_sc_hd__decap_3
XPHY_183 sky130_fd_sc_hd__decap_3
Xclkbuf_8_63_0_CLK clkbuf_8_63_0_CLK/A clkbuf_8_63_0_CLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_194 sky130_fd_sc_hd__decap_3
X_61200_ _66518_/B _59771_/X _61200_/C _61200_/X sky130_fd_sc_hd__or3_4
X_46134_ _46134_/A _46135_/A sky130_fd_sc_hd__inv_2
X_43346_ _41328_/X _43336_/X _87467_/Q _43337_/X _87467_/D sky130_fd_sc_hd__a2bb2o_4
X_62180_ _62179_/X _62181_/B sky130_fd_sc_hd__buf_2
X_74166_ _74166_/A _74073_/X _74166_/Y sky130_fd_sc_hd__nor2_4
X_40558_ _40558_/A _48606_/A _40558_/X sky130_fd_sc_hd__or2_4
X_71378_ _71373_/X _83521_/Q _71377_/Y _83521_/D sky130_fd_sc_hd__a21o_4
X_61131_ _61153_/A _61202_/B _61131_/Y sky130_fd_sc_hd__nand2_4
X_73117_ _73186_/A _86516_/Q _73117_/X sky130_fd_sc_hd__and2_4
X_70329_ _70320_/X _74742_/B _70328_/X _70329_/X sky130_fd_sc_hd__a21o_4
X_46065_ _46065_/A _86786_/D sky130_fd_sc_hd__inv_2
X_43277_ _43180_/A _43277_/X sky130_fd_sc_hd__buf_2
X_74097_ _74097_/A _74073_/X _74097_/Y sky130_fd_sc_hd__nor2_4
X_78974_ _78979_/A _78979_/B _78975_/B sky130_fd_sc_hd__xor2_4
X_40489_ _40489_/A _40471_/X _40489_/X sky130_fd_sc_hd__or2_4
X_45016_ _56395_/C _44945_/X _45015_/X _45016_/Y sky130_fd_sc_hd__o21ai_4
X_42228_ _42276_/A _42228_/X sky130_fd_sc_hd__buf_2
X_61062_ _60880_/X _61037_/A _60891_/Y _61041_/Y _61061_/Y _61062_/Y
+ sky130_fd_sc_hd__a41oi_4
X_73048_ _74414_/B _73048_/B _73048_/X sky130_fd_sc_hd__xor2_4
X_77925_ _82072_/Q _77925_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_78_0_CLK clkbuf_8_79_0_CLK/A clkbuf_8_78_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_60013_ _45943_/A _60109_/A sky130_fd_sc_hd__buf_2
X_49824_ _49821_/Y _49815_/X _49823_/X _86317_/D sky130_fd_sc_hd__a21oi_4
X_65870_ _65045_/A _65888_/B sky130_fd_sc_hd__buf_2
X_42159_ _42154_/X _42141_/X _41193_/X _88004_/Q _42142_/X _42159_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77856_ _77845_/Y _77856_/Y sky130_fd_sc_hd__inv_2
X_64821_ _64678_/X _85529_/Q _64679_/X _64820_/X _64821_/X sky130_fd_sc_hd__a211o_4
X_76807_ _76801_/B _76801_/A _76806_/Y _76807_/Y sky130_fd_sc_hd__a21oi_4
X_49755_ _49751_/A _49750_/X _49761_/C _52971_/D _49755_/X sky130_fd_sc_hd__and4_4
X_46967_ _83716_/Q _54469_/B sky130_fd_sc_hd__inv_2
X_77787_ _77787_/A _77786_/X _77796_/B sky130_fd_sc_hd__xnor2_4
X_74999_ _80768_/Q _75020_/C _74999_/X sky130_fd_sc_hd__xor2_4
X_48706_ _49212_/A _48872_/B _48706_/Y sky130_fd_sc_hd__nand2_4
X_67540_ _67539_/X _88171_/Q _67540_/X sky130_fd_sc_hd__and2_4
X_79526_ _79529_/B _79526_/Y sky130_fd_sc_hd__inv_2
X_45918_ _65381_/A _44024_/A _44157_/Y _45918_/Y sky130_fd_sc_hd__a21oi_4
X_64752_ _64752_/A _64752_/X sky130_fd_sc_hd__buf_2
X_76738_ _76724_/Y _76737_/X _76738_/Y sky130_fd_sc_hd__nand2_4
X_49686_ _49683_/Y _49677_/X _49685_/X _49686_/Y sky130_fd_sc_hd__a21oi_4
X_61964_ _61949_/A _61949_/B _61949_/C _63182_/B _61964_/X sky130_fd_sc_hd__and4_4
X_46898_ _46898_/A _52739_/B sky130_fd_sc_hd__inv_2
X_63703_ _63484_/A _63703_/B _63672_/C _60682_/A _63703_/X sky130_fd_sc_hd__and4_4
X_60915_ _60915_/A _60915_/X sky130_fd_sc_hd__buf_2
X_48637_ _48629_/Y _48585_/X _48636_/X _86505_/D sky130_fd_sc_hd__a21oi_4
X_67471_ _67166_/X _67458_/Y _67390_/X _67470_/Y _67471_/X sky130_fd_sc_hd__a211o_4
X_79457_ _79455_/X _79457_/B _79470_/B sky130_fd_sc_hd__xnor2_4
X_45849_ _45846_/X _45848_/Y _45803_/X _45849_/Y sky130_fd_sc_hd__a21oi_4
X_64683_ _64683_/A _64937_/B sky130_fd_sc_hd__buf_2
X_76669_ _76667_/Y _81684_/Q _76669_/Y sky130_fd_sc_hd__nand2_4
X_61895_ _61719_/A _61895_/X sky130_fd_sc_hd__buf_2
X_69210_ _87034_/Q _69153_/X _69168_/X _69209_/X _69210_/X sky130_fd_sc_hd__a211o_4
X_66422_ _66073_/X _65833_/B _66075_/X _66422_/Y sky130_fd_sc_hd__nand3_4
X_78408_ _78407_/Y _78405_/A _78408_/C _78411_/B sky130_fd_sc_hd__nand3_4
X_63634_ _63624_/X _63625_/X _63628_/X _63631_/X _63633_/Y _63634_/Y
+ sky130_fd_sc_hd__o41ai_4
X_48568_ _48635_/A _48624_/B sky130_fd_sc_hd__buf_2
X_60846_ _60845_/Y _59579_/A _60846_/Y sky130_fd_sc_hd__nor2_4
X_79388_ _79374_/A _79373_/Y _79388_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_16_0_CLK clkbuf_7_8_0_CLK/X clkbuf_9_33_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_69141_ _87039_/Q _69058_/X _69103_/X _69140_/X _69141_/X sky130_fd_sc_hd__a211o_4
X_47519_ _47565_/A _47519_/X sky130_fd_sc_hd__buf_2
X_66353_ _64710_/A _86530_/Q _66353_/X sky130_fd_sc_hd__and2_4
X_78339_ _78339_/A _78339_/B _78340_/B sky130_fd_sc_hd__nor2_4
X_63565_ _58434_/A _63541_/B _63575_/C _63541_/D _63565_/Y sky130_fd_sc_hd__nand4_4
X_60777_ _78064_/A _59803_/X _60776_/Y _84569_/D sky130_fd_sc_hd__a21bo_4
X_48499_ _48499_/A _48635_/A sky130_fd_sc_hd__buf_2
X_65304_ _65614_/A _65304_/X sky130_fd_sc_hd__buf_2
X_50530_ _50496_/A _50552_/B sky130_fd_sc_hd__buf_2
X_62516_ _84836_/Q _60056_/A _62515_/X _62516_/X sky130_fd_sc_hd__a21o_4
X_81350_ _81346_/CLK _81350_/D _81350_/Q sky130_fd_sc_hd__dfxtp_4
X_69072_ _64777_/A _69073_/A sky130_fd_sc_hd__buf_2
X_66284_ _64714_/X _86215_/Q _64716_/X _66283_/X _66284_/X sky130_fd_sc_hd__a211o_4
X_63496_ _63496_/A _63496_/B _63458_/X _63496_/D _63496_/X sky130_fd_sc_hd__and4_4
X_80301_ _80300_/Y _80301_/Y sky130_fd_sc_hd__inv_2
X_68023_ _67550_/X _68023_/X sky130_fd_sc_hd__buf_2
X_65235_ _65172_/X _86121_/Q _65127_/X _65234_/X _65235_/X sky130_fd_sc_hd__a211o_4
X_50461_ _50496_/A _50492_/B sky130_fd_sc_hd__buf_2
X_62447_ _62532_/A _62491_/C sky130_fd_sc_hd__buf_2
X_81281_ _81697_/CLK _81313_/Q _76636_/A sky130_fd_sc_hd__dfxtp_4
X_52200_ _52197_/Y _52170_/X _52199_/X _85870_/D sky130_fd_sc_hd__a21oi_4
X_83020_ _80670_/CLK _74602_/Y _83020_/Q sky130_fd_sc_hd__dfxtp_4
X_80232_ _59982_/C _63784_/C _80232_/X sky130_fd_sc_hd__xor2_4
X_53180_ _85682_/Q _53172_/X _53179_/Y _53180_/Y sky130_fd_sc_hd__o21ai_4
X_65166_ _65162_/X _65631_/B _65165_/X _65166_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_3_2_1_CLK clkbuf_3_2_1_CLK/A clkbuf_4_5_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_50392_ _50390_/Y _50380_/X _50391_/Y _50392_/Y sky130_fd_sc_hd__a21boi_4
X_62378_ _62406_/A _62378_/B _62378_/C _62378_/D _62378_/Y sky130_fd_sc_hd__nand4_4
X_52131_ _52129_/Y _52108_/X _52130_/X _52131_/Y sky130_fd_sc_hd__a21oi_4
X_64117_ _64115_/Y _64073_/X _64116_/Y _84273_/D sky130_fd_sc_hd__a21oi_4
X_61329_ _61329_/A _61329_/B _61375_/C _61329_/Y sky130_fd_sc_hd__nand3_4
X_80163_ _84944_/Q _84192_/Q _80163_/Y sky130_fd_sc_hd__nand2_4
X_65097_ _64846_/X _85550_/Q _64919_/X _65096_/X _65097_/X sky130_fd_sc_hd__a211o_4
X_69974_ _69971_/X _69973_/X _69974_/Y sky130_fd_sc_hd__nand2_4
X_52062_ _50360_/A _52098_/B _52033_/X _52062_/X sky130_fd_sc_hd__and3_4
X_68925_ _87081_/Q _68832_/X _68875_/X _68924_/X _68925_/X sky130_fd_sc_hd__a211o_4
X_64048_ _63741_/A _64048_/X sky130_fd_sc_hd__buf_2
X_84971_ _86530_/CLK _84971_/D _84971_/Q sky130_fd_sc_hd__dfxtp_4
X_80094_ _80071_/X _80084_/X _80094_/Y sky130_fd_sc_hd__nand2_4
X_51013_ _51013_/A _51029_/B sky130_fd_sc_hd__buf_2
X_86710_ _86711_/CLK _86710_/D _58700_/A sky130_fd_sc_hd__dfxtp_4
X_83922_ _83932_/CLK _69464_/X _83922_/Q sky130_fd_sc_hd__dfxtp_4
X_56870_ _55675_/X _56869_/Y _56691_/A _56870_/Y sky130_fd_sc_hd__a21oi_4
X_68856_ _68666_/X _68612_/X _68847_/Y _68855_/Y _68856_/X sky130_fd_sc_hd__a211o_4
X_87690_ _87950_/CLK _42842_/X _87690_/Q sky130_fd_sc_hd__dfxtp_4
X_55821_ _55817_/A _55821_/B _55821_/X sky130_fd_sc_hd__and2_4
X_86641_ _86640_/CLK _47381_/Y _86641_/Q sky130_fd_sc_hd__dfxtp_4
X_67807_ _68637_/A _67901_/A sky130_fd_sc_hd__buf_2
X_83853_ _86988_/CLK _70088_/X _83853_/Q sky130_fd_sc_hd__dfxtp_4
X_68787_ _68783_/X _68786_/X _68737_/X _68787_/Y sky130_fd_sc_hd__a21oi_4
X_65999_ _65999_/A _65999_/B _65999_/Y sky130_fd_sc_hd__nand2_4
X_58540_ _58984_/A _58557_/B sky130_fd_sc_hd__buf_2
X_82804_ _82803_/CLK _82836_/Q _82804_/Q sky130_fd_sc_hd__dfxtp_4
X_55752_ _55749_/X _55752_/B _55752_/Y sky130_fd_sc_hd__nand2_4
X_67738_ _87906_/Q _67713_/X _67641_/X _67737_/X _67738_/X sky130_fd_sc_hd__a211o_4
X_86572_ _86570_/CLK _86572_/D _66211_/B sky130_fd_sc_hd__dfxtp_4
X_52964_ _52960_/Y _52946_/X _52963_/X _85723_/D sky130_fd_sc_hd__a21oi_4
X_83784_ _85953_/CLK _70376_/Y _83784_/Q sky130_fd_sc_hd__dfxtp_4
X_80996_ _85315_/CLK _84204_/Q _80996_/Q sky130_fd_sc_hd__dfxtp_4
X_88311_ _88056_/CLK _88311_/D _69935_/B sky130_fd_sc_hd__dfxtp_4
X_54703_ _54729_/A _54703_/X sky130_fd_sc_hd__buf_2
X_85523_ _85815_/CLK _54012_/Y _85523_/Q sky130_fd_sc_hd__dfxtp_4
X_51915_ _51912_/Y _51904_/X _51914_/X _51915_/Y sky130_fd_sc_hd__a21oi_4
X_82735_ _84177_/CLK _82735_/D _82735_/Q sky130_fd_sc_hd__dfxtp_4
X_58471_ _58467_/X _58468_/Y _58470_/Y _84841_/D sky130_fd_sc_hd__a21oi_4
X_55683_ _55683_/A _55683_/B _55429_/Y _55683_/D _55683_/Y sky130_fd_sc_hd__nand4_4
X_67669_ _67666_/X _67668_/X _67619_/X _67674_/A sky130_fd_sc_hd__a21o_4
X_52895_ _52895_/A _52879_/B _52872_/C _52895_/D _52895_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_360_0_CLK clkbuf_9_180_0_CLK/X _84930_/CLK sky130_fd_sc_hd__clkbuf_1
X_57422_ _56724_/A _57445_/B _56723_/Y _57422_/Y sky130_fd_sc_hd__nand3_4
X_69408_ _81390_/D _69367_/X _69407_/X _83926_/D sky130_fd_sc_hd__a21bo_4
X_88242_ _82906_/CLK _88242_/D _67373_/B sky130_fd_sc_hd__dfxtp_4
X_54634_ _54625_/A _54645_/B _54618_/X _54634_/D _54634_/X sky130_fd_sc_hd__and4_4
X_85454_ _85778_/CLK _85454_/D _85454_/Q sky130_fd_sc_hd__dfxtp_4
X_51846_ _51789_/A _51846_/X sky130_fd_sc_hd__buf_2
X_70680_ _70664_/X _47480_/A _70679_/Y _83726_/D sky130_fd_sc_hd__a21o_4
X_82666_ _82879_/CLK _82710_/Q _82666_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_990_0_CLK clkbuf_9_495_0_CLK/X _85561_/CLK sky130_fd_sc_hd__clkbuf_1
X_84405_ _84403_/CLK _84405_/D _76981_/B sky130_fd_sc_hd__dfxtp_4
X_57353_ _56885_/A _56884_/Y _44287_/X _57353_/Y sky130_fd_sc_hd__a21oi_4
X_81617_ _81260_/CLK _81617_/D _81809_/D sky130_fd_sc_hd__dfxtp_4
X_69339_ _83931_/Q _69299_/X _69338_/X _69339_/X sky130_fd_sc_hd__a21bo_4
X_88173_ _87472_/CLK _88173_/D _67482_/B sky130_fd_sc_hd__dfxtp_4
X_54565_ _54565_/A _54559_/B _54565_/C _54565_/D _54565_/X sky130_fd_sc_hd__and4_4
X_85385_ _85379_/CLK _54749_/Y _85385_/Q sky130_fd_sc_hd__dfxtp_4
X_51777_ _51794_/A _51782_/B _51755_/X _51777_/D _51777_/X sky130_fd_sc_hd__and4_4
X_82597_ _82879_/CLK _78838_/B _82565_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_481_0_CLK clkbuf_8_240_0_CLK/X clkbuf_9_481_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_56304_ _56035_/X _56290_/X _56303_/Y _85243_/D sky130_fd_sc_hd__o21ai_4
X_87124_ _87137_/CLK _87124_/D _87124_/Q sky130_fd_sc_hd__dfxtp_4
X_41530_ _41486_/A _41530_/X sky130_fd_sc_hd__buf_2
X_53516_ _53503_/X _53516_/B _53516_/Y sky130_fd_sc_hd__nand2_4
X_72350_ _72339_/X _85326_/Q _72255_/X _72350_/X sky130_fd_sc_hd__o21a_4
X_84336_ _84263_/CLK _84336_/D _79245_/A sky130_fd_sc_hd__dfxtp_4
X_50728_ _50728_/A _50799_/A sky130_fd_sc_hd__buf_2
X_81548_ _81352_/CLK _76745_/X _81548_/Q sky130_fd_sc_hd__dfxtp_4
X_57284_ _57284_/A _57340_/C _56715_/Y _57284_/Y sky130_fd_sc_hd__nand3_4
X_54496_ _54486_/X _47016_/A _54496_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_375_0_CLK clkbuf_9_187_0_CLK/X _85754_/CLK sky130_fd_sc_hd__clkbuf_1
X_59023_ _59013_/X _85759_/Q _58928_/X _59023_/X sky130_fd_sc_hd__o21a_4
X_71301_ _48024_/B _71290_/X _71300_/Y _83543_/D sky130_fd_sc_hd__o21ai_4
X_56235_ _56233_/A _56243_/B _85265_/Q _56235_/Y sky130_fd_sc_hd__nand3_4
X_41461_ _41460_/Y _41461_/X sky130_fd_sc_hd__buf_2
X_87055_ _88060_/CLK _87055_/D _87055_/Q sky130_fd_sc_hd__dfxtp_4
X_53447_ _53447_/A _53661_/A sky130_fd_sc_hd__buf_2
X_72281_ _72143_/X _85364_/Q _72280_/X _72281_/Y sky130_fd_sc_hd__o21ai_4
X_84267_ _84652_/CLK _64188_/Y _79908_/B sky130_fd_sc_hd__dfxtp_4
X_50659_ _50538_/A _50668_/C sky130_fd_sc_hd__buf_2
X_81479_ _81575_/CLK _81479_/D _76691_/A sky130_fd_sc_hd__dfxtp_4
X_43200_ _43031_/X _43125_/X _40921_/X _43199_/Y _43021_/X _87542_/D
+ sky130_fd_sc_hd__o32ai_4
X_74020_ _74015_/X _74018_/X _74019_/X _74025_/A sky130_fd_sc_hd__a21o_4
X_86006_ _86005_/CLK _86006_/D _86006_/Q sky130_fd_sc_hd__dfxtp_4
X_40412_ _40408_/X _40410_/X _88395_/Q _40411_/X _88395_/D sky130_fd_sc_hd__a2bb2o_4
X_71232_ _71232_/A _71232_/B _71232_/C _71232_/Y sky130_fd_sc_hd__nand3_4
X_83218_ _83218_/CLK _83218_/D _79267_/B sky130_fd_sc_hd__dfxtp_4
X_44180_ _64713_/A _64817_/A sky130_fd_sc_hd__buf_2
X_56166_ _56142_/X _56164_/X _56165_/Y _85284_/D sky130_fd_sc_hd__o21ai_4
X_41392_ _41324_/X _82893_/Q _41391_/X _41392_/Y sky130_fd_sc_hd__o21ai_4
X_53378_ _53351_/A _53378_/X sky130_fd_sc_hd__buf_2
X_84198_ _84194_/CLK _84198_/D _65481_/C sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_496_0_CLK clkbuf_9_497_0_CLK/A clkbuf_9_496_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_43131_ _87565_/Q _43131_/Y sky130_fd_sc_hd__inv_2
X_55117_ _55115_/Y _55102_/X _55116_/X _55117_/Y sky130_fd_sc_hd__a21oi_4
X_40343_ _40343_/A _40344_/A sky130_fd_sc_hd__buf_2
X_52329_ _52327_/Y _52314_/X _52328_/X _52329_/Y sky130_fd_sc_hd__a21oi_4
X_71163_ _71163_/A _71164_/B sky130_fd_sc_hd__buf_2
X_83149_ _86218_/CLK _73483_/X _83149_/Q sky130_fd_sc_hd__dfxtp_4
X_56097_ _56082_/X _56094_/X _56096_/Y _56097_/Y sky130_fd_sc_hd__o21ai_4
X_70114_ _83130_/Q _70114_/Y sky130_fd_sc_hd__inv_2
X_43062_ _43038_/X _43050_/X _40656_/X _73845_/A _43061_/X _43062_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55048_ _55054_/A _54880_/B _55048_/Y sky130_fd_sc_hd__nand2_4
X_59925_ _59880_/X _59883_/Y _59926_/A sky130_fd_sc_hd__and2_4
X_71094_ _71093_/X _71095_/A sky130_fd_sc_hd__buf_2
X_75971_ _75971_/A _81737_/D _81762_/D sky130_fd_sc_hd__xor2_4
X_87957_ _87952_/CLK _87957_/D _87957_/Q sky130_fd_sc_hd__dfxtp_4
X_42013_ _42013_/A _42013_/X sky130_fd_sc_hd__buf_2
X_77710_ _77710_/A _77709_/X _77718_/A sky130_fd_sc_hd__nand2_4
X_74922_ _80757_/Q _74921_/B _74923_/B sky130_fd_sc_hd__nand2_4
X_70045_ _68807_/X _68809_/X _70044_/X _70045_/Y sky130_fd_sc_hd__a21oi_4
X_86908_ _84538_/CLK _44955_/Y _64246_/B sky130_fd_sc_hd__dfxtp_4
X_47870_ _47867_/X _46285_/A _47869_/Y _47871_/A sky130_fd_sc_hd__o21ai_4
X_59856_ _59651_/A _59700_/Y _59717_/Y _59746_/Y _59855_/Y _84687_/D
+ sky130_fd_sc_hd__a41oi_4
X_78690_ _78691_/A _82684_/D _78690_/Y sky130_fd_sc_hd__nor2_4
X_87888_ _87888_/CLK _42387_/X _87888_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_313_0_CLK clkbuf_9_156_0_CLK/X _84760_/CLK sky130_fd_sc_hd__clkbuf_1
X_46821_ _46820_/Y _52694_/D sky130_fd_sc_hd__buf_2
X_58807_ _58807_/A _58873_/B _58807_/Y sky130_fd_sc_hd__nor2_4
X_77641_ _77645_/B _77643_/A sky130_fd_sc_hd__inv_2
X_74853_ _80931_/Q _74853_/B _74853_/X sky130_fd_sc_hd__xor2_4
X_86839_ _86841_/CLK _45961_/Y _44104_/A sky130_fd_sc_hd__dfxtp_4
X_59787_ _60132_/A _59787_/X sky130_fd_sc_hd__buf_2
X_56999_ _56996_/Y _56998_/Y _56982_/X _56999_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_943_0_CLK clkbuf_9_471_0_CLK/X _88062_/CLK sky130_fd_sc_hd__clkbuf_1
X_49540_ _86368_/Q _49524_/X _49539_/Y _49540_/Y sky130_fd_sc_hd__o21ai_4
X_73804_ _73948_/A _73804_/X sky130_fd_sc_hd__buf_2
X_46752_ _46845_/A _46784_/B sky130_fd_sc_hd__buf_2
X_58738_ _84803_/Q _58738_/Y sky130_fd_sc_hd__inv_2
X_77572_ _77553_/A _77553_/B _77552_/A _77572_/X sky130_fd_sc_hd__o21a_4
X_43964_ _43957_/A _44313_/B _43964_/X sky130_fd_sc_hd__and2_4
X_74784_ _74784_/A _74781_/Y _74782_/Y _74783_/Y _74784_/Y sky130_fd_sc_hd__nand4_4
X_71996_ _72007_/A _71996_/B _71996_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_434_0_CLK clkbuf_9_435_0_CLK/A clkbuf_9_434_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_79311_ _79309_/X _79311_/B _79324_/B sky130_fd_sc_hd__xnor2_4
X_45703_ _85101_/Q _45793_/B _45703_/Y sky130_fd_sc_hd__nor2_4
X_76523_ _76522_/Y _76524_/C sky130_fd_sc_hd__inv_2
X_42915_ _42914_/Y _87653_/D sky130_fd_sc_hd__inv_2
X_49471_ _49444_/A _49481_/A sky130_fd_sc_hd__buf_2
X_73735_ _74012_/A _73735_/X sky130_fd_sc_hd__buf_2
X_46683_ _46678_/Y _46654_/X _46682_/X _86715_/D sky130_fd_sc_hd__a21oi_4
X_58669_ _58667_/X _86105_/Q _58668_/X _58669_/Y sky130_fd_sc_hd__o21ai_4
X_70947_ _70947_/A _70947_/B _70947_/C _70947_/Y sky130_fd_sc_hd__nand3_4
X_43895_ _43810_/A _43895_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_328_0_CLK clkbuf_9_164_0_CLK/X _86647_/CLK sky130_fd_sc_hd__clkbuf_1
X_48422_ _83587_/Q _53647_/B sky130_fd_sc_hd__inv_2
X_60700_ _60700_/A _60612_/B _60700_/C _60700_/Y sky130_fd_sc_hd__nor3_4
X_79242_ _79225_/Y _79224_/A _79224_/B _79242_/Y sky130_fd_sc_hd__a21boi_4
X_45634_ _45631_/Y _45632_/X _45616_/X _45633_/Y _45634_/X sky130_fd_sc_hd__a211o_4
X_76454_ _76455_/A _76455_/B _76453_/Y _76454_/X sky130_fd_sc_hd__o21a_4
X_42846_ _40554_/X _42846_/X sky130_fd_sc_hd__buf_2
X_61680_ _61690_/A _61690_/B _79128_/B _61680_/Y sky130_fd_sc_hd__nor3_4
X_73666_ _73641_/A _86557_/Q _73666_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_958_0_CLK clkbuf_9_479_0_CLK/X _83158_/CLK sky130_fd_sc_hd__clkbuf_1
X_70878_ _71068_/B _70880_/B sky130_fd_sc_hd__buf_2
X_75405_ _75404_/A _75383_/X _75384_/X _75405_/Y sky130_fd_sc_hd__a21oi_4
X_60631_ _59619_/X _60299_/C _60629_/Y _60631_/D _60632_/A sky130_fd_sc_hd__nand4_4
X_48353_ _86530_/Q _48350_/X _48352_/Y _48353_/Y sky130_fd_sc_hd__o21ai_4
X_72617_ _72617_/A _79211_/A sky130_fd_sc_hd__inv_2
X_79173_ _79173_/A _79173_/Y sky130_fd_sc_hd__inv_2
X_45565_ _45555_/X _45562_/Y _45564_/Y _86869_/D sky130_fd_sc_hd__a21oi_4
X_76385_ _76383_/X _76353_/Y _76384_/Y _76385_/X sky130_fd_sc_hd__a21o_4
X_42777_ _42776_/Y _87724_/D sky130_fd_sc_hd__inv_2
X_73597_ _73250_/A _73597_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_449_0_CLK clkbuf_8_224_0_CLK/X clkbuf_9_449_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_47304_ _47300_/Y _47271_/X _47303_/X _86649_/D sky130_fd_sc_hd__a21oi_4
X_78124_ _82569_/Q _78124_/B _78130_/D sky130_fd_sc_hd__xor2_4
X_44516_ _44516_/A _44516_/X sky130_fd_sc_hd__buf_2
X_63350_ _62186_/X _60541_/Y _63348_/Y _63349_/X _63350_/X sky130_fd_sc_hd__a211o_4
X_75336_ _75317_/Y _75314_/Y _75315_/Y _75336_/X sky130_fd_sc_hd__o21a_4
X_41728_ _41727_/X _41722_/X _88161_/Q _41723_/X _88161_/D sky130_fd_sc_hd__a2bb2o_4
X_48284_ _48264_/X _50328_/B _48284_/Y sky130_fd_sc_hd__nand2_4
X_60562_ _65842_/A _60562_/B _60555_/A _60562_/Y sky130_fd_sc_hd__nor3_4
X_72548_ _72506_/Y _72546_/Y _72517_/A _72525_/Y _72547_/Y _72548_/Y
+ sky130_fd_sc_hd__a41oi_4
X_45496_ _45493_/X _45495_/Y _45348_/X _45496_/Y sky130_fd_sc_hd__a21oi_4
X_62301_ _62287_/X _62290_/X _62299_/Y _58166_/A _62300_/X _62301_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47235_ _81824_/Q _47236_/A sky130_fd_sc_hd__inv_2
X_78055_ _84560_/Q _62122_/C _78055_/X sky130_fd_sc_hd__xor2_4
X_44447_ _44547_/A _44447_/X sky130_fd_sc_hd__buf_2
X_63281_ _84873_/Q _63281_/B _63301_/C _63281_/D _63281_/X sky130_fd_sc_hd__or4_4
X_75267_ _75267_/A _75267_/Y sky130_fd_sc_hd__inv_2
X_41659_ _40421_/X _41659_/X sky130_fd_sc_hd__buf_2
X_60493_ _60493_/A _60493_/X sky130_fd_sc_hd__buf_2
X_72479_ _72419_/X _85346_/Q _72478_/X _72479_/Y sky130_fd_sc_hd__o21ai_4
X_65020_ _65196_/A _64913_/B _84218_/Q _65020_/X sky130_fd_sc_hd__and3_4
X_77006_ _77004_/Y _77006_/B _77006_/Y sky130_fd_sc_hd__xnor2_4
X_62232_ _62471_/A _62597_/D sky130_fd_sc_hd__buf_2
X_74218_ _74155_/X _84965_/Q _72992_/X _74217_/X _74218_/X sky130_fd_sc_hd__a211o_4
X_47166_ _47165_/Y _52889_/B sky130_fd_sc_hd__buf_2
X_44378_ _40353_/Y _44454_/A sky130_fd_sc_hd__buf_2
X_75198_ _80778_/Q _81034_/D _75198_/X sky130_fd_sc_hd__xor2_4
X_46117_ _46204_/B _46204_/C _46204_/D _46117_/X sky130_fd_sc_hd__and3_4
X_43329_ _43020_/A _43329_/X sky130_fd_sc_hd__buf_2
X_62163_ _62162_/X _62175_/B _61761_/C _62060_/X _62163_/Y sky130_fd_sc_hd__nand4_4
X_74149_ _72757_/A _74232_/A sky130_fd_sc_hd__buf_2
X_47097_ _46909_/X _47109_/A sky130_fd_sc_hd__buf_2
X_61114_ _61112_/X _61205_/A _61144_/A _64285_/A sky130_fd_sc_hd__a21boi_4
X_46048_ _46046_/X _46032_/X _41514_/X _66830_/B _46047_/X _46049_/A
+ sky130_fd_sc_hd__o32ai_4
X_66971_ _66971_/A _66971_/X sky130_fd_sc_hd__buf_2
X_62094_ _61730_/X _62094_/B _59722_/X _62094_/D _62094_/X sky130_fd_sc_hd__and4_4
X_78957_ _78957_/A _78957_/B _78958_/B sky130_fd_sc_hd__xor2_4
Xclkbuf_5_13_0_CLK clkbuf_4_6_1_CLK/X clkbuf_6_27_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_68710_ _68706_/X _68709_/X _68661_/X _68710_/Y sky130_fd_sc_hd__a21oi_4
X_65922_ _65733_/X _85632_/Q _65734_/X _65921_/X _65922_/X sky130_fd_sc_hd__a211o_4
X_77908_ _77908_/A _77907_/Y _77916_/A sky130_fd_sc_hd__xor2_4
X_61045_ _44315_/A _61412_/A sky130_fd_sc_hd__buf_2
X_69690_ _69485_/A _69690_/X sky130_fd_sc_hd__buf_2
X_78888_ _78888_/A _78888_/B _78889_/B sky130_fd_sc_hd__xnor2_4
X_49807_ _49807_/A _49830_/B _49795_/X _53019_/D _49807_/X sky130_fd_sc_hd__and4_4
X_68641_ _69661_/A _68641_/B _68641_/Y sky130_fd_sc_hd__nor2_4
X_65853_ _65850_/X _65725_/B _65852_/X _65853_/Y sky130_fd_sc_hd__nand3_4
X_77839_ _77827_/A _77826_/Y _77813_/A _77838_/Y _77839_/X sky130_fd_sc_hd__a2bb2o_4
X_47999_ _47832_/A _48755_/A sky130_fd_sc_hd__buf_2
X_64804_ _64804_/A _64804_/B _64804_/X sky130_fd_sc_hd__and2_4
X_49738_ _49657_/A _49761_/C sky130_fd_sc_hd__buf_2
X_80850_ _81130_/CLK _80882_/Q _74957_/B sky130_fd_sc_hd__dfxtp_4
X_68572_ _68444_/A _88363_/Q _68572_/X sky130_fd_sc_hd__and2_4
Xclkbuf_5_28_0_CLK clkbuf_4_14_1_CLK/X clkbuf_6_57_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_65784_ _65660_/X _83058_/Q _65768_/X _65783_/X _65784_/X sky130_fd_sc_hd__a211o_4
X_62996_ _62992_/Y _62987_/X _62995_/Y _84362_/D sky130_fd_sc_hd__a21oi_4
X_79509_ _79510_/B _79510_/A _82848_/D sky130_fd_sc_hd__xor2_4
X_67523_ _66563_/A _67997_/A sky130_fd_sc_hd__buf_2
X_64735_ _64657_/X _83309_/Q _64733_/X _64734_/X _64735_/X sky130_fd_sc_hd__a211o_4
X_49669_ _49651_/X _49669_/B _49669_/C _51192_/D _49669_/X sky130_fd_sc_hd__and4_4
X_61947_ _61915_/A _61945_/X _58528_/A _61947_/D _61947_/X sky130_fd_sc_hd__and4_4
X_80781_ _80849_/CLK _80781_/D _80781_/Q sky130_fd_sc_hd__dfxtp_4
X_51700_ _51698_/Y _51693_/X _51699_/X _85962_/D sky130_fd_sc_hd__a21oi_4
X_82520_ _82617_/CLK _82520_/D _78644_/A sky130_fd_sc_hd__dfxtp_4
X_67454_ _87470_/Q _67358_/X _67360_/X _67453_/X _67454_/X sky130_fd_sc_hd__a211o_4
X_52680_ _52708_/A _52694_/C sky130_fd_sc_hd__buf_2
X_64666_ _64666_/A _64666_/X sky130_fd_sc_hd__buf_2
X_61878_ _61876_/X _61846_/B _61878_/C _61846_/D _61879_/D sky130_fd_sc_hd__nand4_4
X_66405_ _66282_/X _66030_/Y _66404_/Y _66405_/Y sky130_fd_sc_hd__o21ai_4
X_51631_ _51628_/Y _51613_/X _51630_/X _51631_/Y sky130_fd_sc_hd__a21oi_4
X_63617_ _58393_/Y _63648_/B _63617_/Y sky130_fd_sc_hd__nor2_4
X_82451_ _82820_/CLK _79143_/X _82419_/D sky130_fd_sc_hd__dfxtp_4
X_60829_ _72592_/A _59837_/B _84556_/Q _60829_/Y sky130_fd_sc_hd__nor3_4
X_67385_ _67364_/X _67385_/B _67385_/X sky130_fd_sc_hd__and2_4
X_64597_ _64683_/A _64633_/B sky130_fd_sc_hd__buf_2
X_81402_ _81352_/CLK _83938_/Q _76715_/B sky130_fd_sc_hd__dfxtp_4
X_69124_ _69371_/A _69124_/X sky130_fd_sc_hd__buf_2
X_54350_ _54322_/A _54355_/A sky130_fd_sc_hd__buf_2
X_66336_ _65074_/A _86563_/Q _66336_/X sky130_fd_sc_hd__and2_4
X_85170_ _85297_/CLK _85170_/D _55848_/B sky130_fd_sc_hd__dfxtp_4
X_51562_ _85987_/Q _51539_/X _51561_/Y _51562_/Y sky130_fd_sc_hd__o21ai_4
X_63548_ _63487_/A _63548_/X sky130_fd_sc_hd__buf_2
X_82382_ _83703_/CLK _82190_/Q _82382_/Q sky130_fd_sc_hd__dfxtp_4
X_53301_ _53355_/A _53301_/X sky130_fd_sc_hd__buf_2
X_84121_ _82177_/CLK _84121_/D _84121_/Q sky130_fd_sc_hd__dfxtp_4
X_50513_ _50513_/A _52216_/B _50513_/Y sky130_fd_sc_hd__nand2_4
X_81333_ _81333_/CLK _81333_/D _81333_/Q sky130_fd_sc_hd__dfxtp_4
X_69055_ _69648_/A _69055_/B _69055_/Y sky130_fd_sc_hd__nor2_4
X_54281_ _54288_/A _52590_/B _54281_/Y sky130_fd_sc_hd__nand2_4
X_66267_ _65486_/A _66267_/X sky130_fd_sc_hd__buf_2
X_51493_ _51218_/X _51509_/A sky130_fd_sc_hd__buf_2
X_63479_ _63417_/A _63491_/D sky130_fd_sc_hd__buf_2
X_68006_ _68402_/A _68006_/X sky130_fd_sc_hd__buf_2
X_56020_ _56019_/Y _56020_/X sky130_fd_sc_hd__buf_2
X_53232_ _53246_/A _53232_/B _53232_/Y sky130_fd_sc_hd__nand2_4
X_65218_ _65215_/X _65111_/B _65217_/X _65218_/Y sky130_fd_sc_hd__nand3_4
X_84052_ _81431_/CLK _84052_/D _84052_/Q sky130_fd_sc_hd__dfxtp_4
X_50444_ _50441_/Y _50429_/X _50443_/X _86200_/D sky130_fd_sc_hd__a21oi_4
X_81264_ _81361_/CLK _81264_/D _76345_/A sky130_fd_sc_hd__dfxtp_4
X_66198_ _44263_/X _66198_/B _66198_/X sky130_fd_sc_hd__and2_4
X_83003_ _85144_/CLK _83003_/D _45494_/A sky130_fd_sc_hd__dfxtp_4
X_80215_ _80215_/A _63800_/C _80215_/X sky130_fd_sc_hd__xor2_4
X_53163_ _53189_/A _53163_/X sky130_fd_sc_hd__buf_2
X_65149_ _65145_/X _65148_/X _65122_/X _65154_/A sky130_fd_sc_hd__a21o_4
X_50375_ _86213_/Q _50363_/X _50374_/Y _50375_/Y sky130_fd_sc_hd__o21ai_4
X_81195_ _81195_/CLK _74964_/X _46504_/A sky130_fd_sc_hd__dfxtp_4
X_52114_ _52112_/Y _52108_/X _52113_/X _85886_/D sky130_fd_sc_hd__a21oi_4
X_87811_ _87553_/CLK _42586_/Y _87811_/Q sky130_fd_sc_hd__dfxtp_4
X_80146_ _80142_/X _80145_/Y _80157_/A sky130_fd_sc_hd__xor2_4
X_53094_ _53147_/A _53115_/A sky130_fd_sc_hd__buf_2
X_57971_ _57971_/A _57971_/B _57971_/Y sky130_fd_sc_hd__nor2_4
X_69957_ _43201_/A _66571_/X _68741_/X _69956_/X _69957_/X sky130_fd_sc_hd__a211o_4
X_59710_ _63344_/B _59741_/A _62975_/D _59890_/C _63055_/A _59710_/Y
+ sky130_fd_sc_hd__a41oi_4
X_52045_ _52058_/A _48297_/X _52045_/Y sky130_fd_sc_hd__nand2_4
X_56922_ _83330_/Q _56922_/X sky130_fd_sc_hd__buf_2
X_68908_ _69685_/A _87325_/Q _68908_/X sky130_fd_sc_hd__and2_4
X_87742_ _87487_/CLK _87742_/D _68896_/B sky130_fd_sc_hd__dfxtp_4
X_80077_ _80056_/B _80073_/X _80076_/Y _80077_/Y sky130_fd_sc_hd__a21oi_4
X_84954_ _84829_/CLK _84954_/D _84954_/Q sky130_fd_sc_hd__dfxtp_4
X_69888_ _69900_/A _69888_/B _69888_/X sky130_fd_sc_hd__and2_4
X_59641_ _61276_/B _60403_/A _60402_/A _59661_/A sky130_fd_sc_hd__and3_4
X_83905_ _83905_/CLK _83905_/D _83905_/Q sky130_fd_sc_hd__dfxtp_4
X_56853_ _56824_/X _85128_/Q _56853_/Y sky130_fd_sc_hd__nand2_4
X_68839_ _69685_/A _87328_/Q _68839_/X sky130_fd_sc_hd__and2_4
X_87673_ _87671_/CLK _87673_/D _67188_/B sky130_fd_sc_hd__dfxtp_4
X_84885_ _84885_/CLK _84885_/D _64525_/C sky130_fd_sc_hd__dfxtp_4
X_55804_ _56246_/C _55311_/X _44046_/X _55803_/X _55804_/X sky130_fd_sc_hd__a211o_4
X_86624_ _84922_/CLK _86624_/D _72129_/A sky130_fd_sc_hd__dfxtp_4
X_71850_ _71867_/B _71857_/B sky130_fd_sc_hd__buf_2
X_83836_ _83191_/CLK _83836_/D _74763_/C sky130_fd_sc_hd__dfxtp_4
X_59572_ _60160_/B _60620_/B sky130_fd_sc_hd__buf_2
X_56784_ _56768_/Y _56785_/D sky130_fd_sc_hd__buf_2
X_53996_ _85526_/Q _53989_/X _53995_/Y _53996_/Y sky130_fd_sc_hd__o21ai_4
X_70801_ _70800_/X _70802_/A sky130_fd_sc_hd__buf_2
X_58523_ _84828_/Q _63520_/B sky130_fd_sc_hd__buf_2
Xclkbuf_7_111_0_CLK clkbuf_6_55_0_CLK/X clkbuf_8_223_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_55735_ _55728_/Y _55729_/Y _55734_/Y _56158_/A sky130_fd_sc_hd__a21oi_4
X_86555_ _85915_/CLK _48214_/Y _65997_/B sky130_fd_sc_hd__dfxtp_4
X_40961_ _40960_/Y _88303_/D sky130_fd_sc_hd__inv_2
X_52947_ _52893_/X _52947_/X sky130_fd_sc_hd__buf_2
X_71781_ _71823_/A _71783_/A sky130_fd_sc_hd__buf_2
X_83767_ _82251_/CLK _70474_/Y _58350_/A sky130_fd_sc_hd__dfxtp_4
X_80979_ _81061_/CLK _75731_/X _75138_/B sky130_fd_sc_hd__dfxtp_4
X_42700_ _42700_/A _42700_/X sky130_fd_sc_hd__buf_2
X_73520_ _73359_/X _83051_/Q _73406_/X _73519_/X _73521_/B sky130_fd_sc_hd__a211o_4
X_85506_ _86733_/CLK _54092_/Y _85506_/Q sky130_fd_sc_hd__dfxtp_4
X_58454_ _83476_/Q _58454_/Y sky130_fd_sc_hd__inv_2
X_70732_ _71735_/D _70732_/X sky130_fd_sc_hd__buf_2
X_82718_ _81216_/CLK _79071_/X _82674_/D sky130_fd_sc_hd__dfxtp_4
X_43680_ _40776_/X _43671_/X _72800_/A _43673_/X _43680_/X sky130_fd_sc_hd__a2bb2o_4
X_55666_ _55657_/Y _55656_/X _55666_/Y sky130_fd_sc_hd__nand2_4
X_86486_ _85879_/CLK _86486_/D _86486_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_81_0_CLK clkbuf_9_40_0_CLK/X _86896_/CLK sky130_fd_sc_hd__clkbuf_1
X_40892_ _82857_/Q _40883_/B _40892_/X sky130_fd_sc_hd__or2_4
X_52878_ _52852_/A _52879_/B sky130_fd_sc_hd__buf_2
X_83698_ _83699_/CLK _70797_/Y _47135_/A sky130_fd_sc_hd__dfxtp_4
X_57405_ _57394_/X _56639_/X _45599_/A _57395_/X _85012_/D sky130_fd_sc_hd__a2bb2o_4
X_88225_ _88158_/CLK _88225_/D _67767_/B sky130_fd_sc_hd__dfxtp_4
X_42631_ _53189_/A _42631_/X sky130_fd_sc_hd__buf_2
X_54617_ _54616_/X _54625_/A sky130_fd_sc_hd__buf_2
X_85437_ _85757_/CLK _85437_/D _85437_/Q sky130_fd_sc_hd__dfxtp_4
X_73451_ _72910_/A _73497_/A sky130_fd_sc_hd__buf_2
X_51829_ _51827_/Y _51823_/X _51828_/X _85939_/D sky130_fd_sc_hd__a21oi_4
X_70663_ _70884_/A _70635_/A _70662_/X _70591_/A _70664_/A sky130_fd_sc_hd__nand4_4
X_58385_ _84862_/Q _58385_/Y sky130_fd_sc_hd__inv_2
X_82649_ _81755_/CLK _84001_/Q _79012_/A sky130_fd_sc_hd__dfxtp_4
X_55597_ _45444_/A _55571_/X _55610_/A _55596_/Y _55597_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_7_126_0_CLK clkbuf_6_63_0_CLK/X clkbuf_8_253_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_72402_ _57800_/X _72400_/Y _72401_/Y _64761_/B _59833_/X _72402_/X
+ sky130_fd_sc_hd__o32a_4
X_45350_ _45350_/A _45350_/X sky130_fd_sc_hd__buf_2
X_57336_ _57335_/Y _85033_/D sky130_fd_sc_hd__inv_2
X_76170_ _81347_/Q _81603_/D _76170_/X sky130_fd_sc_hd__xor2_4
X_88156_ _87141_/CLK _88156_/D _67885_/B sky130_fd_sc_hd__dfxtp_4
X_42562_ _87819_/Q _69676_/B sky130_fd_sc_hd__inv_2
X_54548_ _54521_/A _54559_/B sky130_fd_sc_hd__buf_2
X_73382_ _72908_/X _85577_/Q _72909_/X _73381_/X _73382_/X sky130_fd_sc_hd__a211o_4
X_85368_ _83275_/CLK _85368_/D _85368_/Q sky130_fd_sc_hd__dfxtp_4
X_70594_ _70620_/D _70594_/X sky130_fd_sc_hd__buf_2
X_44301_ _44006_/X _44164_/X _44300_/Y _44301_/Y sky130_fd_sc_hd__nand3_4
X_75121_ _75119_/X _75121_/B _75122_/A sky130_fd_sc_hd__nand2_4
X_87107_ _87417_/CLK _87107_/D _87107_/Q sky130_fd_sc_hd__dfxtp_4
X_41513_ _41513_/A _82326_/Q _41513_/X sky130_fd_sc_hd__or2_4
X_72333_ _72270_/X _72331_/Y _72332_/Y _72296_/X _72274_/X _72333_/X
+ sky130_fd_sc_hd__o32a_4
X_84319_ _84321_/CLK _84319_/D _63493_/C sky130_fd_sc_hd__dfxtp_4
X_45281_ _45281_/A _45281_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_96_0_CLK clkbuf_9_48_0_CLK/X _85134_/CLK sky130_fd_sc_hd__clkbuf_1
X_57267_ _56755_/X _57140_/B _56759_/X _57272_/D _57267_/X sky130_fd_sc_hd__and4_4
X_88087_ _88087_/CLK _41972_/Y _74204_/A sky130_fd_sc_hd__dfxtp_4
X_42493_ _42466_/X _42467_/X _40661_/X _68692_/A _42480_/X _42494_/A
+ sky130_fd_sc_hd__o32ai_4
X_54479_ _85434_/Q _54457_/X _54478_/Y _54479_/Y sky130_fd_sc_hd__o21ai_4
X_85299_ _85279_/CLK _85299_/D _56080_/C sky130_fd_sc_hd__dfxtp_4
X_47020_ _54498_/D _52805_/D sky130_fd_sc_hd__buf_2
X_59006_ _58920_/A _86368_/Q _59006_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_8_242_0_CLK clkbuf_8_243_0_CLK/A clkbuf_8_242_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_44232_ _44227_/Y _44232_/B _44242_/C _44232_/Y sky130_fd_sc_hd__nand3_4
X_56218_ _56123_/A _56229_/B sky130_fd_sc_hd__buf_2
X_75052_ _75047_/Y _75023_/B _75051_/X _75053_/B sky130_fd_sc_hd__o21ai_4
X_87038_ _86989_/CLK _44605_/X _87038_/Q sky130_fd_sc_hd__dfxtp_4
X_41444_ _41444_/A _41444_/Y sky130_fd_sc_hd__inv_2
X_72264_ _57708_/X _72264_/X sky130_fd_sc_hd__buf_2
X_57198_ _56842_/X _57198_/B _57198_/X sky130_fd_sc_hd__xor2_4
X_74003_ _74002_/X _74003_/B _74003_/Y sky130_fd_sc_hd__nand2_4
X_71215_ _71507_/A _70428_/A _71215_/C _71215_/Y sky130_fd_sc_hd__nor3_4
X_44163_ _44162_/Y _44163_/B _87184_/D sky130_fd_sc_hd__nor2_4
X_56149_ _56123_/A _56150_/B sky130_fd_sc_hd__buf_2
X_79860_ _79845_/X _79860_/B _79860_/Y sky130_fd_sc_hd__nand2_4
X_41375_ _41373_/X _41719_/A _41374_/X _41376_/A sky130_fd_sc_hd__o21a_4
X_72195_ _72137_/X _72192_/Y _72193_/Y _72194_/X _72141_/X _72195_/X
+ sky130_fd_sc_hd__o32a_4
X_43114_ _43105_/X _43106_/X _40767_/X _43113_/Y _43108_/X _43114_/Y
+ sky130_fd_sc_hd__o32ai_4
X_78811_ _82547_/Q _78812_/A sky130_fd_sc_hd__inv_2
X_40326_ _40326_/A _40629_/A sky130_fd_sc_hd__buf_2
X_71146_ _71225_/A _71155_/B sky130_fd_sc_hd__buf_2
X_48971_ _48965_/Y _48935_/X _48970_/X _86457_/D sky130_fd_sc_hd__a21oi_4
X_44094_ _55140_/A _44095_/A sky130_fd_sc_hd__buf_2
X_79791_ _79778_/X _79789_/X _79790_/X _79791_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_252_0_CLK clkbuf_9_126_0_CLK/X _81857_/CLK sky130_fd_sc_hd__clkbuf_1
X_47922_ _83777_/Q _73765_/A sky130_fd_sc_hd__inv_2
X_43045_ _43030_/A _43046_/A sky130_fd_sc_hd__buf_2
X_59908_ _61066_/B _61277_/C _59909_/C sky130_fd_sc_hd__nor2_4
X_78742_ _78742_/A _78742_/B _78742_/X sky130_fd_sc_hd__or2_4
X_71077_ _52307_/B _71070_/X _71076_/Y _83616_/D sky130_fd_sc_hd__o21ai_4
X_75954_ _75954_/A _75953_/Y _75955_/B sky130_fd_sc_hd__xnor2_4
Xclkbuf_10_882_0_CLK clkbuf_9_441_0_CLK/X _86414_/CLK sky130_fd_sc_hd__clkbuf_1
X_74905_ _74905_/A _74904_/Y _74906_/B sky130_fd_sc_hd__xor2_4
X_70028_ _82549_/D _70010_/X _70027_/X _70028_/X sky130_fd_sc_hd__a21bo_4
X_47853_ _83559_/Q _47853_/Y sky130_fd_sc_hd__inv_2
X_59839_ _59839_/A _59839_/Y sky130_fd_sc_hd__inv_2
X_78673_ _78638_/B _78655_/B _78653_/X _78673_/X sky130_fd_sc_hd__a21bo_4
Xclkbuf_10_34_0_CLK clkbuf_9_17_0_CLK/X _83008_/CLK sky130_fd_sc_hd__clkbuf_1
X_75885_ _75796_/Y _80795_/D sky130_fd_sc_hd__inv_2
Xclkbuf_9_373_0_CLK clkbuf_9_373_0_CLK/A clkbuf_9_373_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_46804_ _83669_/Q _52686_/B sky130_fd_sc_hd__inv_2
X_77624_ _77606_/A _77623_/Y _77590_/B _77624_/Y sky130_fd_sc_hd__o21ai_4
X_62850_ _62791_/X _62894_/A sky130_fd_sc_hd__buf_2
X_74836_ _74844_/A _46092_/X _74836_/Y sky130_fd_sc_hd__nand2_4
X_47784_ _47784_/A _53244_/D sky130_fd_sc_hd__buf_2
X_44996_ _44975_/X _61386_/B _44995_/X _44996_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_267_0_CLK clkbuf_9_133_0_CLK/X _84960_/CLK sky130_fd_sc_hd__clkbuf_1
X_49523_ _49519_/Y _49514_/X _49522_/X _86372_/D sky130_fd_sc_hd__a21oi_4
X_61801_ _61645_/A _61801_/X sky130_fd_sc_hd__buf_2
X_46735_ _46735_/A _46735_/Y sky130_fd_sc_hd__inv_2
X_77555_ _77535_/Y _77537_/A _77533_/Y _77555_/X sky130_fd_sc_hd__o21a_4
X_43947_ _87176_/Q _43948_/B sky130_fd_sc_hd__inv_2
X_62781_ _62778_/X _62779_/X _62780_/Y _84383_/D sky130_fd_sc_hd__a21oi_4
X_74767_ _83804_/Q _74738_/A _74761_/Y _74762_/Y _74766_/X _74767_/X
+ sky130_fd_sc_hd__a2111o_4
X_71979_ _48926_/A _71959_/X _71964_/X _71979_/X sky130_fd_sc_hd__and3_4
Xclkbuf_10_897_0_CLK clkbuf_9_448_0_CLK/X _86988_/CLK sky130_fd_sc_hd__clkbuf_1
X_64520_ _79568_/B _79566_/A sky130_fd_sc_hd__inv_2
X_76506_ _76502_/Y _76504_/Y _76501_/Y _76510_/C sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_49_0_CLK clkbuf_9_24_0_CLK/X _85041_/CLK sky130_fd_sc_hd__clkbuf_1
X_61732_ _59722_/A _61732_/X sky130_fd_sc_hd__buf_2
X_49454_ _49454_/A _50976_/B _49454_/Y sky130_fd_sc_hd__nand2_4
X_73718_ _73719_/B _73719_/C _73717_/X _73718_/X sky130_fd_sc_hd__a21o_4
X_46666_ _46902_/A _46667_/A sky130_fd_sc_hd__buf_2
X_77486_ _82228_/Q _77486_/Y sky130_fd_sc_hd__inv_2
X_43878_ _43877_/Y _87221_/D sky130_fd_sc_hd__inv_2
X_74698_ _74675_/X _57068_/X _74697_/Y _74698_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_388_0_CLK clkbuf_9_389_0_CLK/A clkbuf_9_388_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_48405_ _48405_/A _48136_/B _48405_/X sky130_fd_sc_hd__or2_4
X_79225_ _79208_/Y _79209_/Y _79205_/Y _79225_/Y sky130_fd_sc_hd__o21ai_4
X_45617_ _45617_/A _45617_/B _45617_/Y sky130_fd_sc_hd__nor2_4
X_64451_ _64446_/Y _64447_/X _64448_/X _64450_/Y _64440_/X _64451_/X
+ sky130_fd_sc_hd__o41a_4
X_76437_ _76430_/A _76430_/B _76429_/A _76437_/X sky130_fd_sc_hd__o21a_4
X_42829_ _42828_/Y _87696_/D sky130_fd_sc_hd__inv_2
X_49385_ _49493_/A _49408_/C sky130_fd_sc_hd__buf_2
X_61663_ _61636_/A _61663_/B _61682_/C _61663_/Y sky130_fd_sc_hd__nand3_4
X_73649_ _73227_/A _73649_/X sky130_fd_sc_hd__buf_2
X_46597_ _86722_/Q _46474_/X _46596_/Y _46597_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_820_0_CLK clkbuf_9_410_0_CLK/X _81190_/CLK sky130_fd_sc_hd__clkbuf_1
X_63402_ _61368_/A _63389_/B _63418_/C _63389_/D _63402_/Y sky130_fd_sc_hd__nand4_4
X_48336_ _86533_/Q _48333_/X _48335_/Y _48336_/Y sky130_fd_sc_hd__o21ai_4
X_60614_ _60182_/Y _59536_/A _61285_/C _60622_/A sky130_fd_sc_hd__and3_4
X_67170_ _67241_/A _86781_/Q _67170_/X sky130_fd_sc_hd__and2_4
X_79156_ _79156_/A _84488_/Q _79156_/X sky130_fd_sc_hd__xor2_4
X_45548_ _45389_/X _45548_/X sky130_fd_sc_hd__buf_2
X_64382_ _64380_/X _84819_/Q _64381_/X _64382_/Y sky130_fd_sc_hd__nand3_4
X_76368_ _76368_/A _76368_/Y sky130_fd_sc_hd__inv_2
X_61594_ _61323_/B _61594_/X sky130_fd_sc_hd__buf_2
X_66121_ _66116_/X _65967_/B _66120_/X _66121_/Y sky130_fd_sc_hd__nand3_4
X_78107_ _78107_/A _78107_/B _78107_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_9_311_0_CLK clkbuf_9_311_0_CLK/A clkbuf_9_311_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_63333_ _60433_/A _63333_/B _63333_/C _60484_/A _63333_/X sky130_fd_sc_hd__and4_4
X_75319_ _75314_/Y _75319_/B _75320_/A sky130_fd_sc_hd__nor2_4
X_48267_ _52139_/A _48545_/A sky130_fd_sc_hd__buf_2
X_60545_ _60515_/A _60488_/A _65842_/A _60546_/A sky130_fd_sc_hd__a21o_4
X_79087_ _79065_/A _79087_/B _79088_/A sky130_fd_sc_hd__and2_4
X_45479_ _45479_/A _45604_/B _45479_/Y sky130_fd_sc_hd__nor2_4
X_76299_ _76290_/B _81644_/Q _76298_/Y _76299_/Y sky130_fd_sc_hd__a21boi_4
Xclkbuf_10_205_0_CLK clkbuf_9_102_0_CLK/X _84652_/CLK sky130_fd_sc_hd__clkbuf_1
X_47218_ _47210_/A _47181_/B _47210_/C _47218_/D _47218_/X sky130_fd_sc_hd__and4_4
X_66052_ _65117_/A _66053_/A sky130_fd_sc_hd__buf_2
X_78038_ _77872_/Y _81938_/D sky130_fd_sc_hd__inv_2
X_63264_ _60410_/B _63333_/C sky130_fd_sc_hd__buf_2
X_48198_ _48190_/A _51954_/B _48198_/Y sky130_fd_sc_hd__nand2_4
X_60476_ _60476_/A _60488_/A _60476_/C _60476_/D _60476_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_10_835_0_CLK clkbuf_9_417_0_CLK/X _84175_/CLK sky130_fd_sc_hd__clkbuf_1
X_65003_ _64858_/X _85522_/Q _64859_/X _65002_/X _65003_/X sky130_fd_sc_hd__a211o_4
X_62215_ _62194_/X _62197_/X _62212_/Y _58147_/A _62214_/X _62215_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47149_ _53395_/B _52881_/B sky130_fd_sc_hd__buf_2
X_63195_ _63342_/C _63241_/C sky130_fd_sc_hd__buf_2
Xclkbuf_9_326_0_CLK clkbuf_9_326_0_CLK/A clkbuf_9_326_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_80000_ _80000_/A _79999_/X _80000_/X sky130_fd_sc_hd__xor2_4
X_69811_ _69770_/A _88321_/Q _69811_/X sky130_fd_sc_hd__and2_4
X_50160_ _52370_/A _51256_/B _50147_/C _50160_/X sky130_fd_sc_hd__and3_4
X_62146_ _62037_/X _62063_/X _58296_/A _62183_/D _62146_/X sky130_fd_sc_hd__and4_4
X_79989_ _79989_/A _79989_/Y sky130_fd_sc_hd__inv_2
X_69742_ _69655_/A _69742_/X sky130_fd_sc_hd__buf_2
X_50091_ _64804_/B _50088_/X _50090_/Y _50091_/Y sky130_fd_sc_hd__o21ai_4
X_66954_ _66953_/X _66954_/X sky130_fd_sc_hd__buf_2
X_62077_ _62142_/A _62077_/B _62077_/C _62077_/D _62077_/Y sky130_fd_sc_hd__nand4_4
X_65905_ _65791_/A _65932_/A sky130_fd_sc_hd__buf_2
X_61028_ _61027_/X _61028_/X sky130_fd_sc_hd__buf_2
X_81951_ _82124_/CLK _78012_/Y _77690_/B sky130_fd_sc_hd__dfxtp_4
X_69673_ _69605_/A _87307_/Q _69673_/X sky130_fd_sc_hd__and2_4
X_66885_ _87122_/Q _66833_/X _66834_/X _66884_/X _66885_/X sky130_fd_sc_hd__a211o_4
X_80902_ _84014_/CLK _84078_/Q _75606_/A sky130_fd_sc_hd__dfxtp_4
X_68624_ _68599_/A _68624_/B _68624_/X sky130_fd_sc_hd__and2_4
X_53850_ _53844_/A _72025_/B _53850_/Y sky130_fd_sc_hd__nand2_4
X_65836_ _65836_/A _86470_/Q _65836_/X sky130_fd_sc_hd__and2_4
X_84670_ _84668_/CLK _84670_/D _60051_/C sky130_fd_sc_hd__dfxtp_4
X_81882_ _81883_/CLK _81882_/D _81882_/Q sky130_fd_sc_hd__dfxtp_4
X_52801_ _52784_/X _52818_/B _52789_/X _52801_/D _52801_/X sky130_fd_sc_hd__and4_4
X_83621_ _85561_/CLK _83621_/D _48920_/A sky130_fd_sc_hd__dfxtp_4
X_80833_ _83944_/CLK _83977_/Q _75707_/B sky130_fd_sc_hd__dfxtp_4
X_68555_ _68617_/A _68555_/X sky130_fd_sc_hd__buf_2
X_53781_ _85569_/Q _53754_/X _53780_/Y _53781_/Y sky130_fd_sc_hd__o21ai_4
X_65767_ _65764_/X _65766_/X _65614_/X _65767_/X sky130_fd_sc_hd__a21o_4
X_50993_ _51021_/A _51003_/A sky130_fd_sc_hd__buf_2
X_62979_ _62979_/A _64546_/C _60302_/X _62979_/D _62979_/X sky130_fd_sc_hd__and4_4
X_55520_ _55524_/A _55520_/B _55520_/Y sky130_fd_sc_hd__nor2_4
X_67506_ _67506_/A _67506_/B _67506_/Y sky130_fd_sc_hd__nand2_4
X_86340_ _86340_/CLK _49698_/Y _59360_/B sky130_fd_sc_hd__dfxtp_4
X_52732_ _52718_/A _52732_/B _52732_/Y sky130_fd_sc_hd__nand2_4
X_64718_ _64903_/A _64826_/A sky130_fd_sc_hd__buf_2
X_83552_ _83550_/CLK _83552_/D _83552_/Q sky130_fd_sc_hd__dfxtp_4
X_80764_ _80740_/CLK _75472_/X _81140_/D sky130_fd_sc_hd__dfxtp_4
X_68486_ _87099_/Q _68455_/X _68370_/X _68485_/X _68486_/X sky130_fd_sc_hd__a211o_4
X_65698_ _65621_/A _65775_/B _65698_/C _65698_/X sky130_fd_sc_hd__and3_4
X_82503_ _82503_/CLK _78857_/A _78383_/A sky130_fd_sc_hd__dfxtp_4
X_55451_ _55447_/Y _55451_/B _55676_/B sky130_fd_sc_hd__and2_4
X_67437_ _67342_/A _67437_/B _67437_/X sky130_fd_sc_hd__and2_4
X_86271_ _83307_/CLK _50070_/Y _86271_/Q sky130_fd_sc_hd__dfxtp_4
X_52663_ _52657_/X _52663_/B _52663_/Y sky130_fd_sc_hd__nand2_4
X_64649_ _64649_/A _64648_/X _64649_/Y sky130_fd_sc_hd__nand2_4
X_83483_ _83414_/CLK _83483_/D _83483_/Q sky130_fd_sc_hd__dfxtp_4
X_80695_ _81111_/CLK _80695_/D _75376_/A sky130_fd_sc_hd__dfxtp_4
X_88010_ _87757_/CLK _42151_/X _88010_/Q sky130_fd_sc_hd__dfxtp_4
X_54402_ _54399_/X _54395_/B _54402_/C _46846_/Y _54402_/X sky130_fd_sc_hd__and4_4
X_85222_ _85190_/CLK _85222_/D _55702_/B sky130_fd_sc_hd__dfxtp_4
X_51614_ _51694_/A _51619_/B sky130_fd_sc_hd__buf_2
X_58170_ _46155_/A _58253_/A sky130_fd_sc_hd__buf_2
X_82434_ _82436_/CLK _79126_/X _82434_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_705 sky130_fd_sc_hd__decap_3
X_55382_ _55382_/A _55383_/C sky130_fd_sc_hd__inv_2
X_67368_ _67342_/A _67368_/B _67368_/X sky130_fd_sc_hd__and2_4
XPHY_716 sky130_fd_sc_hd__decap_3
X_52594_ _52614_/A _52594_/B _51919_/C _51768_/D _52594_/X sky130_fd_sc_hd__and4_4
X_57121_ _57096_/Y _57121_/X sky130_fd_sc_hd__buf_2
X_69107_ _68929_/X _69094_/Y _69095_/X _69106_/Y _69107_/X sky130_fd_sc_hd__a211o_4
X_54333_ _85461_/Q _54320_/X _54332_/Y _54333_/Y sky130_fd_sc_hd__o21ai_4
X_66319_ _66318_/X _66319_/B _66319_/C _66319_/X sky130_fd_sc_hd__and3_4
X_85153_ _85311_/CLK _85153_/D _55640_/A sky130_fd_sc_hd__dfxtp_4
X_51545_ _51545_/A _53072_/B _51545_/Y sky130_fd_sc_hd__nand2_4
X_82365_ _82369_/CLK _82365_/D _82365_/Q sky130_fd_sc_hd__dfxtp_4
X_67299_ _67062_/X _67324_/A sky130_fd_sc_hd__buf_2
X_84104_ _80928_/CLK _84104_/D _84104_/Q sky130_fd_sc_hd__dfxtp_4
X_57052_ _46159_/A _57047_/Y _57049_/Y _57051_/Y _57052_/X sky130_fd_sc_hd__a211o_4
X_81316_ _84105_/CLK _76184_/X _81724_/D sky130_fd_sc_hd__dfxtp_4
X_69038_ _87076_/Q _68948_/X _68993_/X _69037_/X _69038_/X sky130_fd_sc_hd__a211o_4
X_54264_ _54286_/A _54246_/X _54255_/C _53099_/D _54264_/X sky130_fd_sc_hd__and4_4
X_85084_ _83008_/CLK _57104_/X _45470_/A sky130_fd_sc_hd__dfxtp_4
X_51476_ _86003_/Q _51458_/X _51475_/Y _51476_/Y sky130_fd_sc_hd__o21ai_4
X_82296_ _82299_/CLK _81920_/Q _82296_/Q sky130_fd_sc_hd__dfxtp_4
X_56003_ _56002_/Y _56003_/B _55966_/X _55975_/X _56003_/Y sky130_fd_sc_hd__nand4_4
X_53215_ _53189_/A _53215_/X sky130_fd_sc_hd__buf_2
X_84035_ _81160_/CLK _68116_/X _84035_/Q sky130_fd_sc_hd__dfxtp_4
X_50427_ _50432_/A _48435_/B _50427_/Y sky130_fd_sc_hd__nand2_4
X_81247_ _85335_/CLK _81055_/Q _47547_/A sky130_fd_sc_hd__dfxtp_4
X_54195_ _54215_/A _47403_/A _54195_/Y sky130_fd_sc_hd__nand2_4
X_71000_ _70772_/A _71001_/C sky130_fd_sc_hd__buf_2
X_41160_ _41061_/X _81720_/Q _41159_/X _41161_/A sky130_fd_sc_hd__o21ai_4
X_53146_ _53172_/A _53146_/X sky130_fd_sc_hd__buf_2
X_50358_ _50398_/A _50358_/B _50358_/Y sky130_fd_sc_hd__nand2_4
X_81178_ _82335_/CLK _75024_/B _40402_/B sky130_fd_sc_hd__dfxtp_4
X_80129_ _80126_/X _80129_/B _81685_/D sky130_fd_sc_hd__xor2_4
X_53077_ _85701_/Q _53065_/X _53076_/Y _53077_/Y sky130_fd_sc_hd__o21ai_4
X_57954_ _58721_/A _57954_/X sky130_fd_sc_hd__buf_2
X_41091_ _40912_/B _41091_/B _41091_/X sky130_fd_sc_hd__or2_4
X_50289_ _50285_/A _48236_/B _50289_/Y sky130_fd_sc_hd__nand2_4
X_85986_ _85697_/CLK _51571_/Y _85986_/Q sky130_fd_sc_hd__dfxtp_4
X_56905_ _83315_/Q _56908_/A sky130_fd_sc_hd__inv_2
X_52028_ _66166_/B _51994_/X _52027_/Y _52028_/Y sky130_fd_sc_hd__o21ai_4
X_87725_ _87221_/CLK _42773_/Y _87725_/Q sky130_fd_sc_hd__dfxtp_4
X_84937_ _85485_/CLK _84937_/D _84937_/Q sky130_fd_sc_hd__dfxtp_4
X_72951_ _72951_/A _72951_/X sky130_fd_sc_hd__buf_2
X_57885_ _57884_/X _85494_/Q _57763_/X _57885_/X sky130_fd_sc_hd__o21a_4
X_71902_ _70591_/A _71902_/X sky130_fd_sc_hd__buf_2
X_59624_ _59619_/X _59621_/X _59753_/B _59624_/X sky130_fd_sc_hd__and3_4
X_44850_ _41744_/Y _44848_/X _86921_/Q _44849_/X _86921_/D sky130_fd_sc_hd__a2bb2o_4
X_56836_ _56759_/X _56866_/A _83333_/Q _56659_/Y _56836_/Y sky130_fd_sc_hd__nand4_4
X_75670_ _75670_/A _75669_/Y _75674_/A sky130_fd_sc_hd__xor2_4
X_87656_ _86932_/CLK _42911_/X _87656_/Q sky130_fd_sc_hd__dfxtp_4
X_72882_ _56181_/X _83077_/Q _72880_/X _72881_/X _72883_/B sky130_fd_sc_hd__a211o_4
X_84868_ _84823_/CLK _58365_/X _84868_/Q sky130_fd_sc_hd__dfxtp_4
X_43801_ _43752_/A _43801_/X sky130_fd_sc_hd__buf_2
X_74621_ _58253_/A _74613_/X _56164_/A _74614_/X _74621_/X sky130_fd_sc_hd__a211o_4
X_86607_ _86610_/CLK _86607_/D _72336_/A sky130_fd_sc_hd__dfxtp_4
X_71833_ _71829_/X _71839_/B _70771_/A _71826_/X _71833_/X sky130_fd_sc_hd__and4_4
X_59555_ _59602_/A _61276_/B sky130_fd_sc_hd__buf_2
X_83819_ _83819_/CLK _70261_/X _74751_/A sky130_fd_sc_hd__dfxtp_4
X_44781_ _44780_/Y _86958_/D sky130_fd_sc_hd__inv_2
X_56767_ _83324_/Q _56767_/X sky130_fd_sc_hd__buf_2
X_87587_ _87588_/CLK _87587_/D _43070_/A sky130_fd_sc_hd__dfxtp_4
X_41993_ _41993_/A _41993_/X sky130_fd_sc_hd__buf_2
X_53979_ _53977_/Y _53948_/X _53978_/Y _85530_/D sky130_fd_sc_hd__a21boi_4
X_84799_ _84797_/CLK _58803_/Y _84799_/Q sky130_fd_sc_hd__dfxtp_4
X_46520_ _54058_/B _51358_/B sky130_fd_sc_hd__buf_2
X_58506_ _58506_/A _58502_/B _58506_/Y sky130_fd_sc_hd__nor2_4
X_77340_ _77339_/B _77339_/A _77340_/Y sky130_fd_sc_hd__nand2_4
X_43732_ _43732_/A _69885_/B sky130_fd_sc_hd__inv_2
X_55718_ _55710_/Y _55712_/Y _55717_/Y _56167_/B sky130_fd_sc_hd__a21oi_4
X_86538_ _86218_/CLK _86538_/D _66242_/B sky130_fd_sc_hd__dfxtp_4
X_74552_ _45932_/Y _74552_/X sky130_fd_sc_hd__buf_2
X_40944_ _40835_/A _40944_/X sky130_fd_sc_hd__buf_2
X_71764_ _71763_/X _71422_/C _70794_/X _71764_/X sky130_fd_sc_hd__and3_4
X_59486_ _63384_/B _58532_/X _59486_/Y sky130_fd_sc_hd__nor2_4
X_56698_ _83337_/Q _56698_/Y sky130_fd_sc_hd__inv_2
X_73503_ _48683_/A _73502_/Y _73503_/X sky130_fd_sc_hd__xor2_4
X_46451_ _50460_/A _53874_/A sky130_fd_sc_hd__buf_2
X_70715_ _52760_/B _70699_/X _70714_/Y _83719_/D sky130_fd_sc_hd__o21ai_4
X_58437_ _63209_/A _58438_/A sky130_fd_sc_hd__buf_2
X_77271_ _77269_/Y _77266_/X _77267_/Y _77274_/B sky130_fd_sc_hd__nand3_4
X_43663_ _43663_/A _43663_/Y sky130_fd_sc_hd__inv_2
X_55649_ _56564_/A _55624_/X _56564_/C _56564_/D _55648_/X _55649_/Y
+ sky130_fd_sc_hd__a41oi_4
X_74483_ _48634_/A _74501_/B _74478_/C _74483_/X sky130_fd_sc_hd__and3_4
X_86469_ _86499_/CLK _48860_/Y _86469_/Q sky130_fd_sc_hd__dfxtp_4
X_40875_ _40870_/X _40871_/X _40874_/X _69842_/B _40867_/X _40875_/Y
+ sky130_fd_sc_hd__o32ai_4
X_71695_ _71690_/Y _71695_/X sky130_fd_sc_hd__buf_2
X_79010_ _79010_/A _79010_/B _79011_/B sky130_fd_sc_hd__xor2_4
X_45402_ _55640_/A _44935_/X _45757_/A _45402_/X sky130_fd_sc_hd__o21a_4
X_76222_ _76221_/Y _76222_/Y sky130_fd_sc_hd__inv_2
X_88208_ _88208_/CLK _88208_/D _66656_/B sky130_fd_sc_hd__dfxtp_4
X_42614_ _42590_/A _42614_/X sky130_fd_sc_hd__buf_2
X_49170_ _81189_/Q _49161_/B _49170_/Y sky130_fd_sc_hd__nor2_4
X_73434_ _73432_/X _73434_/B _73434_/C _73434_/Y sky130_fd_sc_hd__nand3_4
X_46382_ _51294_/B _52478_/B sky130_fd_sc_hd__buf_2
X_70646_ _53021_/B _70632_/X _70645_/Y _83735_/D sky130_fd_sc_hd__o21ai_4
X_58368_ _63344_/A _58370_/A sky130_fd_sc_hd__buf_2
X_43594_ _40559_/X _43586_/X _43587_/Y _43593_/X _43595_/A sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_41_0_CLK clkbuf_7_41_0_CLK/A clkbuf_8_83_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_48121_ _48117_/Y _48109_/X _48120_/X _48121_/Y sky130_fd_sc_hd__a21oi_4
X_45333_ _45330_/X _45332_/Y _45275_/X _45333_/Y sky130_fd_sc_hd__a21oi_4
X_57319_ _56782_/X _57023_/X _56768_/Y _57319_/D _57319_/X sky130_fd_sc_hd__and4_4
X_76153_ _76152_/Y _76153_/Y sky130_fd_sc_hd__inv_2
X_88139_ _86824_/CLK _88139_/D _88139_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_181_0_CLK clkbuf_7_90_0_CLK/X clkbuf_9_363_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_42545_ _72769_/A _69583_/B sky130_fd_sc_hd__inv_2
X_73365_ _73363_/X _73365_/B _73365_/C _73365_/Y sky130_fd_sc_hd__nand3_4
X_70577_ MACRO_WR_SELECT _70578_/A sky130_fd_sc_hd__buf_2
X_58299_ _64536_/C _63694_/B sky130_fd_sc_hd__buf_2
X_75104_ _75104_/A _75104_/B _75104_/C _75105_/A sky130_fd_sc_hd__nand3_4
X_48052_ _48051_/Y _50341_/B sky130_fd_sc_hd__buf_2
X_60330_ _60263_/A _60331_/B _60324_/C _60344_/C _65296_/A _60330_/Y
+ sky130_fd_sc_hd__a41oi_4
X_72316_ _72240_/X _85681_/Q _72241_/X _72316_/X sky130_fd_sc_hd__o21a_4
X_45264_ _85257_/Q _45222_/X _45263_/X _45264_/Y sky130_fd_sc_hd__o21ai_4
X_76084_ _81721_/D _76085_/B _76096_/A sky130_fd_sc_hd__or2_4
X_42476_ _42460_/X _42472_/X _40626_/X _42475_/Y _42463_/X _42476_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73296_ _42600_/A _73053_/B _73296_/Y sky130_fd_sc_hd__nor2_4
X_47003_ _47003_/A _47004_/A sky130_fd_sc_hd__buf_2
X_44215_ _44208_/X _44211_/Y _44214_/X _44215_/X sky130_fd_sc_hd__o21a_4
X_75035_ _75031_/Y _75023_/B _75049_/A _75035_/Y sky130_fd_sc_hd__o21ai_4
X_79912_ _79912_/A _79911_/Y _79912_/Y sky130_fd_sc_hd__nor2_4
X_41427_ _41427_/A _41435_/B _41427_/X sky130_fd_sc_hd__or2_4
X_72247_ _72247_/A _72332_/B _72247_/Y sky130_fd_sc_hd__nor2_4
X_60261_ _60249_/X _60252_/X _60256_/X _60259_/Y _60260_/Y _60261_/Y
+ sky130_fd_sc_hd__a41oi_4
X_45195_ _55817_/B _45194_/X _45153_/X _45195_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_7_56_0_CLK clkbuf_7_57_0_CLK/A clkbuf_7_56_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_62000_ _61957_/A _62000_/B _62000_/C _62000_/D _62000_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_8_196_0_CLK clkbuf_7_98_0_CLK/X clkbuf_9_393_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_44146_ _44146_/A _44147_/A sky130_fd_sc_hd__buf_2
X_79843_ _79836_/X _79838_/B _79843_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_191_0_CLK clkbuf_9_95_0_CLK/X _81070_/CLK sky130_fd_sc_hd__clkbuf_1
X_41358_ _40878_/A _41358_/X sky130_fd_sc_hd__buf_2
X_60192_ _60263_/A _60344_/A _60324_/A _60268_/A _59980_/X _60192_/Y
+ sky130_fd_sc_hd__a41oi_4
X_72178_ _72165_/Y _72152_/X _72171_/X _72177_/X _83277_/D sky130_fd_sc_hd__a22oi_4
X_71129_ _71129_/A _71230_/B _70914_/D _71129_/Y sky130_fd_sc_hd__nand3_4
X_48954_ _83618_/Q _53819_/B sky130_fd_sc_hd__inv_2
X_44077_ _55761_/A _44077_/X sky130_fd_sc_hd__buf_2
X_79774_ _84223_/Q _72236_/A _79774_/X sky130_fd_sc_hd__xor2_4
X_41289_ _41288_/X _41283_/X _67338_/B _41284_/X _88243_/D sky130_fd_sc_hd__a2bb2o_4
X_76986_ _76986_/A _62442_/C _76986_/X sky130_fd_sc_hd__xor2_4
X_47905_ _47972_/A _47963_/B sky130_fd_sc_hd__buf_2
X_43028_ _42439_/X _43017_/X _40581_/X _73599_/A _43025_/X _43029_/A
+ sky130_fd_sc_hd__o32ai_4
X_78725_ _78725_/A _78725_/B _78725_/X sky130_fd_sc_hd__and2_4
X_63951_ _64364_/B _64029_/B _63951_/C _64015_/D _63951_/Y sky130_fd_sc_hd__nand4_4
X_75937_ _75933_/Y _75936_/Y _75939_/B sky130_fd_sc_hd__xnor2_4
X_48885_ _48885_/A _48894_/B _48894_/C _48885_/X sky130_fd_sc_hd__and3_4
X_62902_ _63306_/A _62930_/B sky130_fd_sc_hd__buf_2
X_47836_ _65908_/B _43756_/X _47835_/X _47836_/Y sky130_fd_sc_hd__o21ai_4
X_66670_ _87131_/Q _66593_/X _66594_/X _66669_/X _66670_/X sky130_fd_sc_hd__a211o_4
X_78656_ _78639_/Y _78642_/Y _78638_/B _78657_/B sky130_fd_sc_hd__o21ai_4
X_63882_ _60920_/A _63947_/C sky130_fd_sc_hd__buf_2
X_75868_ _75867_/Y _75852_/A _75868_/X sky130_fd_sc_hd__and2_4
X_65621_ _65621_/A _65559_/B _84189_/Q _65621_/X sky130_fd_sc_hd__and3_4
X_77607_ _77596_/B _77590_/A _77590_/B _77607_/Y sky130_fd_sc_hd__a21boi_4
X_62833_ _62869_/A _62812_/B _61969_/X _62833_/Y sky130_fd_sc_hd__nand3_4
X_74819_ _74818_/Y _80664_/D sky130_fd_sc_hd__inv_2
X_47767_ _81224_/Q _47768_/A sky130_fd_sc_hd__inv_2
X_78587_ _78586_/Y _78587_/Y sky130_fd_sc_hd__inv_2
X_44979_ _45197_/A _44979_/X sky130_fd_sc_hd__buf_2
X_75799_ _75787_/A _75786_/X _75798_/X _75800_/B sky130_fd_sc_hd__a21oi_4
X_49506_ _49500_/A _49516_/B _49493_/X _52720_/D _49506_/X sky130_fd_sc_hd__and4_4
X_68340_ _68319_/X _68077_/Y _68326_/X _68339_/Y _68340_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_8_134_0_CLK clkbuf_7_67_0_CLK/X clkbuf_9_269_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_46718_ _46713_/Y _46704_/X _46717_/X _46718_/Y sky130_fd_sc_hd__a21oi_4
X_65552_ _65503_/X _85593_/Q _65504_/X _65551_/X _65552_/X sky130_fd_sc_hd__a211o_4
X_77538_ _77537_/Y _77538_/B _77539_/A sky130_fd_sc_hd__nand2_4
X_62764_ _62731_/A _59390_/Y _62744_/X _62717_/X _62764_/X sky130_fd_sc_hd__and4_4
X_47698_ _47745_/A _47698_/X sky130_fd_sc_hd__buf_2
X_64503_ _61232_/X _61636_/B _61207_/X _64503_/Y sky130_fd_sc_hd__nand3_4
X_49437_ _49432_/Y _49434_/X _49436_/X _49437_/Y sky130_fd_sc_hd__a21oi_4
X_61715_ _61715_/A _61715_/B _61710_/Y _61714_/Y _61715_/Y sky130_fd_sc_hd__nand4_4
X_68271_ _82644_/D _68259_/X _68270_/X _83996_/D sky130_fd_sc_hd__a21bo_4
X_46649_ _83685_/Q _46650_/A sky130_fd_sc_hd__inv_2
X_65483_ _64665_/A _65484_/A sky130_fd_sc_hd__buf_2
X_77469_ _77455_/Y _77467_/Y _77468_/Y _77478_/A sky130_fd_sc_hd__o21a_4
X_62695_ _62669_/A _63044_/A _62704_/C _62669_/D _62695_/X sky130_fd_sc_hd__and4_4
X_67222_ _67222_/A _67248_/A sky130_fd_sc_hd__buf_2
X_79208_ _79205_/Y _79208_/B _79208_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_250_0_CLK clkbuf_9_251_0_CLK/A clkbuf_9_250_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_64434_ _64494_/A _64434_/B _64391_/X _64434_/X sky130_fd_sc_hd__and3_4
X_49368_ _49504_/A _49451_/A sky130_fd_sc_hd__buf_2
X_61646_ _61634_/A _61634_/B _79131_/B _61646_/Y sky130_fd_sc_hd__nor3_4
X_80480_ _80480_/A _80480_/B _82259_/D sky130_fd_sc_hd__xnor2_4
Xclkbuf_8_149_0_CLK clkbuf_7_74_0_CLK/X clkbuf_9_299_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_48319_ _48319_/A _50365_/B _48319_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_144_0_CLK clkbuf_9_72_0_CLK/X _83188_/CLK sky130_fd_sc_hd__clkbuf_1
X_67153_ _66794_/A _67153_/X sky130_fd_sc_hd__buf_2
X_79139_ _79139_/A _84471_/Q _79139_/X sky130_fd_sc_hd__xor2_4
X_64365_ _64306_/A _64379_/B sky130_fd_sc_hd__buf_2
X_49299_ _49002_/A _49415_/A sky130_fd_sc_hd__buf_2
X_61577_ _61546_/A _61546_/B _61577_/C _61577_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_10_774_0_CLK clkbuf_9_387_0_CLK/X _82518_/CLK sky130_fd_sc_hd__clkbuf_1
X_66104_ _66104_/A _66135_/B sky130_fd_sc_hd__buf_2
X_51330_ _51330_/A _51266_/B _51330_/C _51330_/X sky130_fd_sc_hd__and3_4
X_63316_ _63316_/A _63316_/B _60588_/X _63344_/D _63316_/X sky130_fd_sc_hd__or4_4
X_82150_ _84231_/CLK _84142_/Q _82150_/Q sky130_fd_sc_hd__dfxtp_4
X_60528_ _60528_/A _60529_/A sky130_fd_sc_hd__buf_2
X_67084_ _87422_/Q _67035_/X _66984_/X _67083_/X _67084_/X sky130_fd_sc_hd__a211o_4
X_64296_ _64287_/A _84850_/Q _64287_/C _64296_/Y sky130_fd_sc_hd__nand3_4
X_81101_ _80817_/CLK _79676_/X _75817_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_265_0_CLK clkbuf_8_132_0_CLK/X clkbuf_9_265_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_66035_ _65992_/A _73780_/B _66035_/X sky130_fd_sc_hd__and2_4
X_51261_ _51280_/A _51261_/B _51261_/Y sky130_fd_sc_hd__nand2_4
X_63247_ _63247_/A _63281_/D sky130_fd_sc_hd__buf_2
X_82081_ _81160_/CLK _82081_/D _82081_/Q sky130_fd_sc_hd__dfxtp_4
X_60459_ _60421_/B _60459_/B _60606_/A _60458_/X _60460_/A sky130_fd_sc_hd__nand4_4
X_53000_ _85715_/Q _52984_/X _52999_/Y _53000_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_159_0_CLK clkbuf_9_79_0_CLK/X _81269_/CLK sky130_fd_sc_hd__clkbuf_1
X_50212_ _50212_/A _50595_/A sky130_fd_sc_hd__buf_2
X_81032_ _81928_/CLK _81032_/D _81032_/Q sky130_fd_sc_hd__dfxtp_4
X_51192_ _51191_/X _51192_/B _51192_/C _51192_/D _51192_/X sky130_fd_sc_hd__and4_4
X_63178_ _60607_/A _63192_/D sky130_fd_sc_hd__buf_2
Xclkbuf_10_789_0_CLK clkbuf_9_394_0_CLK/X _82152_/CLK sky130_fd_sc_hd__clkbuf_1
X_50143_ _50140_/Y _50141_/X _50142_/X _86256_/D sky130_fd_sc_hd__a21oi_4
X_62129_ _58287_/A _62129_/X sky130_fd_sc_hd__buf_2
X_85840_ _85558_/CLK _85840_/D _85840_/Q sky130_fd_sc_hd__dfxtp_4
X_67986_ _87896_/Q _67888_/X _67984_/X _67985_/X _67986_/X sky130_fd_sc_hd__a211o_4
X_69725_ _69092_/A _69725_/B _69725_/X sky130_fd_sc_hd__and2_4
X_50074_ _50072_/Y _50068_/X _50073_/X _86270_/D sky130_fd_sc_hd__a21oi_4
X_54951_ _54955_/A _54955_/B _46617_/A _53257_/D _54951_/X sky130_fd_sc_hd__and4_4
X_66937_ _87876_/Q _66935_/X _66911_/X _66936_/X _66937_/X sky130_fd_sc_hd__a211o_4
X_85771_ _85773_/CLK _52699_/Y _85771_/Q sky130_fd_sc_hd__dfxtp_4
X_82983_ _85128_/CLK _74693_/Y _82983_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_712_0_CLK clkbuf_9_356_0_CLK/X _88245_/CLK sky130_fd_sc_hd__clkbuf_1
X_87510_ _87790_/CLK _87510_/D _87510_/Q sky130_fd_sc_hd__dfxtp_4
X_53902_ _53902_/A _53902_/B _53902_/Y sky130_fd_sc_hd__nand2_4
X_84722_ _83464_/CLK _84722_/D _84722_/Q sky130_fd_sc_hd__dfxtp_4
X_57670_ _57670_/A _57666_/B _57670_/Y sky130_fd_sc_hd__nor2_4
X_81934_ _81933_/CLK _81934_/D _77404_/A sky130_fd_sc_hd__dfxtp_4
X_69656_ _69650_/X _69653_/X _69655_/X _69656_/Y sky130_fd_sc_hd__a21oi_4
X_54882_ _54882_/A _54882_/X sky130_fd_sc_hd__buf_2
X_66868_ _66868_/A _66868_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_203_0_CLK clkbuf_9_203_0_CLK/A clkbuf_9_203_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_56621_ _55536_/A _55536_/C _56621_/X sky130_fd_sc_hd__and2_4
X_68607_ _68560_/A _68607_/B _68607_/X sky130_fd_sc_hd__and2_4
X_87441_ _87484_/CLK _87441_/D _87441_/Q sky130_fd_sc_hd__dfxtp_4
X_53833_ _85559_/Q _53816_/X _53832_/Y _53833_/Y sky130_fd_sc_hd__o21ai_4
X_65819_ _65702_/A _85863_/Q _65819_/X sky130_fd_sc_hd__and2_4
X_84653_ _84652_/CLK _60144_/Y _79936_/B sky130_fd_sc_hd__dfxtp_4
X_81865_ _84441_/CLK _78056_/X _81865_/Q sky130_fd_sc_hd__dfxtp_4
X_69587_ _44518_/A _69457_/X _69458_/X _69586_/X _69587_/X sky130_fd_sc_hd__a211o_4
X_66799_ _87370_/Q _66797_/X _66747_/X _66798_/X _66799_/X sky130_fd_sc_hd__a211o_4
X_59340_ _59326_/X _86341_/Q _59340_/Y sky130_fd_sc_hd__nor2_4
X_83604_ _86155_/CLK _83604_/D _49093_/A sky130_fd_sc_hd__dfxtp_4
X_56552_ _56549_/X _45882_/A _45898_/X _56550_/X _56551_/X _56552_/Y
+ sky130_fd_sc_hd__a41oi_4
X_80816_ _80821_/CLK _80816_/D _75851_/B sky130_fd_sc_hd__dfxtp_4
X_68538_ _68516_/X _68525_/Y _68447_/X _68537_/Y _68538_/X sky130_fd_sc_hd__a211o_4
X_87372_ _86834_/CLK _43535_/X _87372_/Q sky130_fd_sc_hd__dfxtp_4
X_53764_ _48680_/A _53774_/B _53774_/C _53764_/X sky130_fd_sc_hd__and3_4
X_84584_ _84564_/CLK _60685_/Y _84584_/Q sky130_fd_sc_hd__dfxtp_4
X_50976_ _50971_/A _50976_/B _50976_/Y sky130_fd_sc_hd__nand2_4
X_81796_ _81668_/CLK _81796_/D _47501_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_727_0_CLK clkbuf_9_363_0_CLK/X _86989_/CLK sky130_fd_sc_hd__clkbuf_1
X_55503_ _55467_/X _55646_/A _55491_/X _55503_/D _55503_/Y sky130_fd_sc_hd__nand4_4
X_86323_ _86322_/CLK _86323_/D _86323_/Q sky130_fd_sc_hd__dfxtp_4
X_52715_ _52770_/A _52724_/B sky130_fd_sc_hd__buf_2
X_59271_ _59133_/A _59271_/X sky130_fd_sc_hd__buf_2
X_83535_ _86535_/CLK _83535_/D _48105_/A sky130_fd_sc_hd__dfxtp_4
X_56483_ _56538_/A _56483_/X sky130_fd_sc_hd__buf_2
X_80747_ _80835_/CLK _80747_/D _81123_/D sky130_fd_sc_hd__dfxtp_4
X_68469_ _73653_/A _68467_/X _68385_/X _68468_/Y _68469_/X sky130_fd_sc_hd__a211o_4
X_53695_ _85586_/Q _53610_/X _53694_/Y _53695_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_218_0_CLK clkbuf_9_219_0_CLK/A clkbuf_9_218_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_70500_ _71136_/A _70500_/B _70758_/B _70500_/D _70500_/Y sky130_fd_sc_hd__nor4_4
X_58222_ _58221_/X _58238_/B _58222_/Y sky130_fd_sc_hd__nor2_4
X_55434_ _55415_/A _55434_/B _55415_/B _55415_/C _55434_/Y sky130_fd_sc_hd__nand4_4
X_86254_ _85554_/CLK _50152_/Y _65096_/B sky130_fd_sc_hd__dfxtp_4
X_40660_ _40577_/X _82868_/Q _40659_/X _40660_/X sky130_fd_sc_hd__o21a_4
X_52646_ _85780_/Q _52629_/X _52645_/Y _52646_/Y sky130_fd_sc_hd__o21ai_4
X_71480_ _71463_/Y _83484_/Q _71479_/X _83484_/D sky130_fd_sc_hd__a21o_4
X_83466_ _85955_/CLK _83466_/D _47817_/A sky130_fd_sc_hd__dfxtp_4
XPHY_502 sky130_fd_sc_hd__decap_3
X_80678_ _80679_/CLK _80710_/Q _80678_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_513 sky130_fd_sc_hd__decap_3
XPHY_524 sky130_fd_sc_hd__decap_3
X_85205_ _86900_/CLK _85205_/D _56407_/C sky130_fd_sc_hd__dfxtp_4
X_70431_ _70442_/A _70940_/B _70431_/C _70431_/Y sky130_fd_sc_hd__nand3_4
X_58153_ _72484_/A _58153_/X sky130_fd_sc_hd__buf_2
XPHY_535 sky130_fd_sc_hd__decap_3
X_82417_ _82820_/CLK _82449_/Q _78524_/A sky130_fd_sc_hd__dfxtp_4
X_55365_ _55336_/X _55365_/B _55366_/A sky130_fd_sc_hd__and2_4
X_86185_ _86500_/CLK _50520_/Y _86185_/Q sky130_fd_sc_hd__dfxtp_4
X_52577_ _52590_/A _52577_/B _52577_/Y sky130_fd_sc_hd__nand2_4
X_40591_ _40344_/A _40591_/B _40591_/C _40591_/X sky130_fd_sc_hd__and3_4
XPHY_546 sky130_fd_sc_hd__decap_3
X_83397_ _83431_/CLK _71728_/Y _83397_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_557 sky130_fd_sc_hd__decap_3
Xclkbuf_4_3_0_CLK clkbuf_4_3_0_CLK/A clkbuf_4_3_0_CLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_568 sky130_fd_sc_hd__decap_3
X_57104_ _57097_/X _56589_/X _45470_/A _57099_/X _57104_/X sky130_fd_sc_hd__a2bb2o_4
X_54316_ _54316_/A _54325_/A sky130_fd_sc_hd__buf_2
X_42330_ _42417_/A _42330_/X sky130_fd_sc_hd__buf_2
X_73150_ _43152_/Y _72895_/X _72858_/X _73149_/Y _73150_/X sky130_fd_sc_hd__a211o_4
XPHY_579 sky130_fd_sc_hd__decap_3
X_85136_ _85103_/CLK _85136_/D _56705_/B sky130_fd_sc_hd__dfxtp_4
X_51528_ _51525_/Y _51503_/X _51527_/X _51528_/Y sky130_fd_sc_hd__a21oi_4
X_58084_ _58079_/X _58081_/Y _58082_/Y _58028_/X _58083_/X _58084_/X
+ sky130_fd_sc_hd__o32a_4
X_70362_ _71003_/A _70361_/Y _70362_/X sky130_fd_sc_hd__and2_4
X_82348_ _82925_/CLK _77123_/X _48056_/A sky130_fd_sc_hd__dfxtp_4
X_55296_ _55296_/A _55296_/B _55297_/A sky130_fd_sc_hd__and2_4
X_72101_ _72091_/X _49176_/A _72101_/Y sky130_fd_sc_hd__nand2_4
X_57035_ _57032_/Y _57034_/Y _57084_/A _57035_/X sky130_fd_sc_hd__a21o_4
X_42261_ _41469_/X _42258_/X _87953_/Q _42259_/X _42261_/X sky130_fd_sc_hd__a2bb2o_4
X_54247_ _54255_/A _54246_/X _54237_/C _53078_/D _54247_/X sky130_fd_sc_hd__and4_4
X_73081_ _73081_/A _73124_/B _73081_/Y sky130_fd_sc_hd__nor2_4
X_85067_ _85067_/CLK _85067_/D _57179_/B sky130_fd_sc_hd__dfxtp_4
X_51459_ _51211_/A _51481_/A sky130_fd_sc_hd__buf_2
X_70293_ _70289_/X _74796_/A _70292_/X _83808_/D sky130_fd_sc_hd__a21o_4
X_82279_ _82284_/CLK _77036_/B _40901_/B sky130_fd_sc_hd__dfxtp_4
X_44000_ _59571_/C _59544_/B sky130_fd_sc_hd__buf_2
X_41212_ _41007_/A _40694_/A _41212_/X sky130_fd_sc_hd__or2_4
X_72032_ _83298_/Q _72016_/X _72031_/Y _72032_/Y sky130_fd_sc_hd__o21ai_4
X_84018_ _84020_/CLK _68183_/X _84018_/Q sky130_fd_sc_hd__dfxtp_4
X_42192_ _42137_/A _42192_/X sky130_fd_sc_hd__buf_2
X_54178_ _54176_/Y _54171_/X _54177_/X _54178_/Y sky130_fd_sc_hd__a21oi_4
X_41143_ _41143_/A _41143_/X sky130_fd_sc_hd__buf_2
X_53129_ _53133_/A _53133_/B _53133_/C _53129_/D _53129_/X sky130_fd_sc_hd__and4_4
X_76840_ _81671_/Q _76840_/B _76840_/Y sky130_fd_sc_hd__xnor2_4
X_58986_ _58982_/X _83437_/Q _58985_/Y _84781_/D sky130_fd_sc_hd__o21a_4
X_45951_ _45935_/X _45951_/Y sky130_fd_sc_hd__inv_2
X_41074_ _82280_/Q _41019_/B _41074_/X sky130_fd_sc_hd__or2_4
X_57937_ _57903_/X _85490_/Q _57849_/X _57937_/X sky130_fd_sc_hd__o21a_4
X_76771_ _76771_/A _76771_/B _76771_/X sky130_fd_sc_hd__xor2_4
X_73983_ _73980_/X _73981_/Y _73982_/X _73983_/X sky130_fd_sc_hd__a21o_4
X_85969_ _85969_/CLK _85969_/D _85969_/Q sky130_fd_sc_hd__dfxtp_4
X_78510_ _78505_/X _78508_/Y _78510_/C _78510_/Y sky130_fd_sc_hd__nand3_4
X_44902_ _44894_/Y _44899_/Y _44901_/X _44902_/X sky130_fd_sc_hd__o21a_4
X_75722_ _75722_/A _75722_/B _75723_/B sky130_fd_sc_hd__nand2_4
X_87708_ _87708_/CLK _87708_/D _67889_/B sky130_fd_sc_hd__dfxtp_4
X_48670_ _48613_/A _48695_/A sky130_fd_sc_hd__buf_2
X_72934_ _72930_/X _72933_/X _72812_/X _72934_/X sky130_fd_sc_hd__a21o_4
X_79490_ _84814_/Q _84134_/Q _79490_/Y sky130_fd_sc_hd__nand2_4
X_45882_ _45882_/A _45883_/B sky130_fd_sc_hd__buf_2
X_57868_ _58696_/A _57868_/X sky130_fd_sc_hd__buf_2
X_47621_ _47620_/X _47649_/A sky130_fd_sc_hd__buf_2
X_59607_ _59637_/A _59608_/A sky130_fd_sc_hd__buf_2
X_78441_ _78450_/A _78450_/B _78441_/X sky130_fd_sc_hd__or2_4
X_44833_ _43896_/X _44833_/X sky130_fd_sc_hd__buf_2
X_56819_ _56649_/X _57186_/B _56818_/X _56820_/A sky130_fd_sc_hd__o21ai_4
X_87639_ _87189_/CLK _87639_/D _87639_/Q sky130_fd_sc_hd__dfxtp_4
X_75653_ _75660_/A _75659_/A _75652_/Y _75653_/Y sky130_fd_sc_hd__a21oi_4
X_72865_ _72896_/B _72865_/X sky130_fd_sc_hd__buf_2
X_57799_ _57866_/A _57800_/A sky130_fd_sc_hd__buf_2
X_74604_ _45244_/Y _74598_/X _74603_/X _74604_/Y sky130_fd_sc_hd__o21ai_4
X_47552_ _47552_/A _53115_/B sky130_fd_sc_hd__buf_2
X_71816_ _71805_/X _83365_/Q _71815_/X _71816_/X sky130_fd_sc_hd__a21o_4
X_59538_ _43995_/A _59876_/B _59538_/C _59538_/D _61078_/B sky130_fd_sc_hd__nand4_4
X_78372_ _78371_/Y _78375_/A sky130_fd_sc_hd__inv_2
X_44764_ _44740_/X _44741_/X _41331_/X _86966_/Q _44742_/X _44765_/A
+ sky130_fd_sc_hd__o32ai_4
X_75584_ _75888_/A _75580_/Y _75584_/C _75584_/Y sky130_fd_sc_hd__nand3_4
X_41976_ _88085_/Q _41976_/Y sky130_fd_sc_hd__inv_2
X_72796_ _42548_/A _73000_/B _72796_/Y sky130_fd_sc_hd__nor2_4
X_46503_ _86731_/Q _46474_/X _46502_/Y _46503_/Y sky130_fd_sc_hd__o21ai_4
X_77323_ _77324_/A _82089_/D _77323_/Y sky130_fd_sc_hd__nor2_4
X_43715_ _43715_/A _43715_/Y sky130_fd_sc_hd__inv_2
X_74535_ _56460_/B _56460_/D _74614_/A sky130_fd_sc_hd__nand2_4
X_40927_ _40927_/A _40842_/X _40927_/X sky130_fd_sc_hd__or2_4
X_47483_ _86630_/Q _47478_/X _47482_/Y _47483_/Y sky130_fd_sc_hd__o21ai_4
X_71747_ _71173_/A _71753_/B _71744_/C _71744_/D _71747_/Y sky130_fd_sc_hd__nand4_4
X_59469_ _59462_/X _83460_/Q _59468_/Y _84724_/D sky130_fd_sc_hd__o21a_4
X_44695_ _86997_/Q _44695_/Y sky130_fd_sc_hd__inv_2
X_49222_ _48548_/A _49222_/X sky130_fd_sc_hd__buf_2
X_61500_ _84819_/Q _61500_/X sky130_fd_sc_hd__buf_2
X_46434_ _46434_/A _51316_/B _46434_/Y sky130_fd_sc_hd__nand2_4
X_77254_ _77254_/A _77254_/Y sky130_fd_sc_hd__inv_2
X_43646_ _43645_/X _87329_/D sky130_fd_sc_hd__inv_2
X_62480_ _61548_/B _62462_/X _62436_/X _62478_/X _62479_/X _62480_/X
+ sky130_fd_sc_hd__a41o_4
X_74466_ _74466_/A _48593_/A _74466_/Y sky130_fd_sc_hd__nand2_4
X_40858_ _40784_/A _40883_/B sky130_fd_sc_hd__buf_2
X_71678_ _71680_/A _71671_/X _71302_/X _71678_/Y sky130_fd_sc_hd__nand3_4
X_76205_ _76205_/A _76205_/Y sky130_fd_sc_hd__inv_2
X_49153_ _49052_/A _49153_/X sky130_fd_sc_hd__buf_2
X_61431_ _59388_/A _61452_/B _61452_/C _61391_/D _61431_/Y sky130_fd_sc_hd__nand4_4
X_73417_ _87289_/Q _73530_/B _73417_/Y sky130_fd_sc_hd__nor2_4
X_46365_ _46290_/A _46366_/A sky130_fd_sc_hd__buf_2
X_70629_ _70668_/D _71735_/C sky130_fd_sc_hd__buf_2
X_77185_ _77184_/X _77185_/Y sky130_fd_sc_hd__inv_2
X_43577_ _43577_/A _87351_/D sky130_fd_sc_hd__inv_2
X_74397_ _74394_/Y _74370_/X _74396_/X _83075_/D sky130_fd_sc_hd__a21oi_4
X_40789_ _40788_/Y _88335_/D sky130_fd_sc_hd__inv_2
X_48104_ _48731_/A _48142_/A sky130_fd_sc_hd__buf_2
X_45316_ _45313_/Y _45315_/Y _45287_/X _45316_/X sky130_fd_sc_hd__a21o_4
X_76136_ _76136_/A _76136_/B _76136_/X sky130_fd_sc_hd__xor2_4
X_64150_ _61652_/B _64161_/B _64150_/C _64161_/D _64150_/Y sky130_fd_sc_hd__nand4_4
X_42528_ _74164_/A _42528_/Y sky130_fd_sc_hd__inv_2
X_49084_ _49056_/A _50153_/B _49084_/Y sky130_fd_sc_hd__nand2_4
X_61362_ _61384_/A _61384_/B _84487_/Q _61362_/Y sky130_fd_sc_hd__nor3_4
X_73348_ _73342_/X _73346_/X _73347_/X _73365_/B sky130_fd_sc_hd__a21o_4
X_46296_ _46421_/A _46295_/X _46296_/Y sky130_fd_sc_hd__nand2_4
X_63101_ _63095_/Y _63097_/X _63098_/X _63100_/X _63067_/X _63101_/Y
+ sky130_fd_sc_hd__o41ai_4
X_48035_ _46493_/X _82350_/Q _48034_/Y _48036_/A sky130_fd_sc_hd__o21ai_4
X_60313_ _60312_/Y _60313_/Y sky130_fd_sc_hd__inv_2
X_45247_ _64466_/B _61590_/B sky130_fd_sc_hd__buf_2
X_64081_ _64458_/B _64179_/B _64081_/C _64179_/D _64081_/Y sky130_fd_sc_hd__nand4_4
X_76067_ _76064_/Y _76066_/X _76067_/Y sky130_fd_sc_hd__nand2_4
X_42459_ _42458_/Y _87857_/D sky130_fd_sc_hd__inv_2
X_61293_ _61293_/A _61293_/B _61278_/B _61295_/A sky130_fd_sc_hd__nand3_4
X_73279_ _74246_/B _73279_/X sky130_fd_sc_hd__buf_2
X_63032_ _60508_/A _63033_/D sky130_fd_sc_hd__buf_2
X_75018_ _75018_/A _75017_/Y _75023_/A sky130_fd_sc_hd__nor2_4
X_60244_ _60244_/A _60244_/B _79863_/A _60244_/Y sky130_fd_sc_hd__nor3_4
X_45178_ _56424_/C _45176_/X _45177_/X _45178_/Y sky130_fd_sc_hd__o21ai_4
X_44129_ _72838_/A _73284_/A sky130_fd_sc_hd__buf_2
X_67840_ _67909_/A _67840_/B _67840_/X sky130_fd_sc_hd__and2_4
X_79826_ _79826_/A _84260_/Q _79834_/B sky130_fd_sc_hd__xor2_4
X_60175_ _60175_/A _60312_/C _60312_/D _61286_/B sky130_fd_sc_hd__nand3_4
X_49986_ _49906_/A _49986_/X sky130_fd_sc_hd__buf_2
X_48937_ _48881_/X _81788_/Q _48936_/Y _48938_/A sky130_fd_sc_hd__o21ai_4
X_67771_ _67793_/A _87649_/Q _67771_/X sky130_fd_sc_hd__and2_4
X_79757_ _79757_/A _79756_/Y _79767_/B sky130_fd_sc_hd__xor2_4
X_64983_ _64978_/X _65056_/B _64982_/X _64995_/A sky130_fd_sc_hd__nand3_4
X_76969_ _76969_/A _81349_/D sky130_fd_sc_hd__inv_2
X_69510_ _87512_/Q _69442_/X _69396_/X _69509_/X _69510_/X sky130_fd_sc_hd__a211o_4
X_66722_ _87885_/Q _66697_/X _66675_/X _66721_/X _66722_/X sky130_fd_sc_hd__a211o_4
X_78708_ _78700_/Y _78706_/B _78722_/A _78721_/A sky130_fd_sc_hd__o21a_4
X_63934_ _64026_/A _63934_/X sky130_fd_sc_hd__buf_2
X_48868_ _50056_/A _48695_/B _48868_/Y sky130_fd_sc_hd__nand2_4
X_79688_ _84214_/Q _83262_/Q _79688_/Y sky130_fd_sc_hd__nand2_4
X_69441_ _88029_/Q _69315_/X _69393_/X _69440_/X _69441_/X sky130_fd_sc_hd__a211o_4
X_47819_ _47819_/A _53259_/B _47819_/Y sky130_fd_sc_hd__nand2_4
X_66653_ _66602_/A _86803_/Q _66653_/X sky130_fd_sc_hd__and2_4
X_78639_ _78639_/A _78639_/Y sky130_fd_sc_hd__inv_2
X_63865_ _63863_/X _63833_/X _63864_/Y _84290_/D sky130_fd_sc_hd__a21oi_4
X_48799_ _48793_/A _48551_/X _48799_/Y sky130_fd_sc_hd__nand2_4
X_65604_ _84190_/Q _65605_/C sky130_fd_sc_hd__inv_2
X_50830_ _52524_/A _50825_/B _50830_/C _50830_/X sky130_fd_sc_hd__and3_4
X_62816_ _62792_/X _62839_/B _62816_/C _62816_/Y sky130_fd_sc_hd__nor3_4
X_81650_ _81362_/CLK _81682_/Q _81650_/Q sky130_fd_sc_hd__dfxtp_4
X_69372_ _69383_/A _69372_/B _69372_/X sky130_fd_sc_hd__and2_4
X_66584_ _44225_/B _88403_/Q _46212_/A _66583_/X _66584_/X sky130_fd_sc_hd__a211o_4
X_63796_ _61780_/X _63860_/B _63738_/C _63738_/D _63796_/Y sky130_fd_sc_hd__nand4_4
X_80601_ _80601_/A _80600_/Y _82270_/D sky130_fd_sc_hd__xor2_4
X_68323_ _67990_/X _67993_/X _68295_/X _68323_/Y sky130_fd_sc_hd__a21oi_4
X_65535_ _65667_/A _72957_/B _65535_/X sky130_fd_sc_hd__and2_4
X_50761_ _50771_/A _49241_/B _50761_/Y sky130_fd_sc_hd__nand2_4
X_62747_ _62766_/A _62766_/B _84386_/Q _62747_/Y sky130_fd_sc_hd__nor3_4
X_81581_ _81587_/CLK _84181_/Q _76753_/A sky130_fd_sc_hd__dfxtp_4
X_52500_ _52438_/A _52500_/X sky130_fd_sc_hd__buf_2
X_83320_ _83325_/CLK _71944_/X _83320_/Q sky130_fd_sc_hd__dfxtp_4
X_80532_ _80531_/B _80531_/A _80532_/X sky130_fd_sc_hd__and2_4
X_68254_ _68097_/A _68254_/X sky130_fd_sc_hd__buf_2
X_53480_ _47886_/X _50475_/B _53697_/C _53480_/Y sky130_fd_sc_hd__nand3_4
X_65466_ _65449_/A _65546_/B _65466_/C _65466_/X sky130_fd_sc_hd__and3_4
X_50692_ _50718_/A _50695_/A sky130_fd_sc_hd__buf_2
X_62678_ _62678_/A _60273_/X _61762_/X _62678_/Y sky130_fd_sc_hd__nand3_4
X_67205_ _67199_/X _67202_/X _67204_/X _67205_/X sky130_fd_sc_hd__a21o_4
X_52431_ _52431_/A _52436_/A sky130_fd_sc_hd__buf_2
X_64417_ _79700_/B _64373_/X _64416_/X _64417_/X sky130_fd_sc_hd__a21o_4
X_83251_ _84192_/CLK _72474_/Y _72465_/A sky130_fd_sc_hd__dfxtp_4
X_61629_ _61608_/X _61629_/B _61619_/C _61629_/Y sky130_fd_sc_hd__nand3_4
X_80463_ _84762_/Q _66138_/A _80472_/A sky130_fd_sc_hd__xor2_4
X_68185_ _68155_/X _67151_/Y _68168_/X _68184_/Y _68185_/X sky130_fd_sc_hd__a211o_4
X_65397_ _65397_/A _65397_/B _65397_/C _65397_/Y sky130_fd_sc_hd__nor3_4
X_82202_ _82961_/CLK _82202_/D _82202_/Q sky130_fd_sc_hd__dfxtp_4
X_55150_ _55224_/A _85066_/Q _55150_/X sky130_fd_sc_hd__and2_4
X_67136_ _67087_/A _67136_/B _67136_/X sky130_fd_sc_hd__and2_4
X_52362_ _52349_/A _50153_/B _52362_/Y sky130_fd_sc_hd__nand2_4
X_64348_ _64342_/X _64343_/X _64345_/X _64347_/Y _64326_/X _64348_/X
+ sky130_fd_sc_hd__o41a_4
X_83182_ _81696_/CLK _83182_/D _83182_/Q sky130_fd_sc_hd__dfxtp_4
X_80394_ _80394_/A _80394_/B _80394_/X sky130_fd_sc_hd__or2_4
X_54101_ _54098_/Y _53437_/X _54100_/X _85504_/D sky130_fd_sc_hd__a21oi_4
X_51313_ _51263_/A _51313_/X sky130_fd_sc_hd__buf_2
X_82133_ _82133_/CLK _82133_/D _82089_/D sky130_fd_sc_hd__dfxtp_4
X_55081_ _85322_/Q _55072_/X _55080_/Y _55081_/Y sky130_fd_sc_hd__o21ai_4
X_67067_ _66899_/X _67054_/Y _67031_/X _67066_/Y _67067_/X sky130_fd_sc_hd__a211o_4
X_52293_ _52293_/A _48944_/B _52293_/Y sky130_fd_sc_hd__nand2_4
X_64279_ _64273_/X _64275_/X _64276_/X _64278_/Y _64267_/X _64279_/X
+ sky130_fd_sc_hd__o41a_4
X_87990_ _87990_/CLK _42187_/X _87990_/Q sky130_fd_sc_hd__dfxtp_4
X_54032_ _54029_/Y _54006_/X _54031_/Y _54032_/Y sky130_fd_sc_hd__a21boi_4
X_66018_ _66015_/Y _65987_/X _66017_/Y _84162_/D sky130_fd_sc_hd__a21o_4
X_51244_ _51240_/A _50738_/B _51244_/Y sky130_fd_sc_hd__nand2_4
X_86941_ _86941_/CLK _86941_/D _67381_/B sky130_fd_sc_hd__dfxtp_4
X_82064_ _80928_/CLK _84024_/Q _77851_/A sky130_fd_sc_hd__dfxtp_4
X_81015_ _84150_/CLK _84223_/Q _81015_/Q sky130_fd_sc_hd__dfxtp_4
X_58840_ _58787_/X _86092_/Q _58839_/X _58840_/Y sky130_fd_sc_hd__o21ai_4
X_51175_ _51147_/A _51175_/X sky130_fd_sc_hd__buf_2
X_86872_ _84418_/CLK _45514_/Y _63089_/B sky130_fd_sc_hd__dfxtp_4
X_50126_ _50106_/A _53854_/B _50126_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_651_0_CLK clkbuf_9_325_0_CLK/X _88224_/CLK sky130_fd_sc_hd__clkbuf_1
X_85823_ _85535_/CLK _85823_/D _85823_/Q sky130_fd_sc_hd__dfxtp_4
X_58771_ _58740_/X _85457_/Q _58770_/X _58771_/Y sky130_fd_sc_hd__o21ai_4
X_67969_ _67966_/X _67968_/X _67875_/X _67969_/Y sky130_fd_sc_hd__a21oi_4
X_55983_ _55983_/A _55983_/B _55984_/A sky130_fd_sc_hd__and2_4
X_57722_ _57722_/A _57697_/X _57722_/Y sky130_fd_sc_hd__nor2_4
X_69708_ _69685_/A _73056_/A _69708_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_142_0_CLK clkbuf_8_71_0_CLK/X clkbuf_9_142_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_50057_ _64627_/B _48861_/X _50056_/Y _50057_/Y sky130_fd_sc_hd__o21ai_4
X_54934_ _54919_/X _47780_/A _54934_/Y sky130_fd_sc_hd__nand2_4
X_85754_ _85754_/CLK _52791_/Y _85754_/Q sky130_fd_sc_hd__dfxtp_4
X_70980_ _50799_/B _70961_/A _70979_/Y _83642_/D sky130_fd_sc_hd__o21ai_4
X_82966_ _82965_/CLK _82966_/D _46727_/A sky130_fd_sc_hd__dfxtp_4
X_84705_ _84329_/CLK _59748_/Y _80539_/A sky130_fd_sc_hd__dfxtp_4
X_57653_ _57652_/X _57657_/B _57653_/Y sky130_fd_sc_hd__nor2_4
X_81917_ _82008_/CLK _77650_/Y _82293_/D sky130_fd_sc_hd__dfxtp_4
X_69639_ _87066_/Q _66550_/X _66552_/X _69638_/X _69639_/X sky130_fd_sc_hd__a211o_4
X_54865_ _54892_/A _54865_/X sky130_fd_sc_hd__buf_2
X_85685_ _84787_/CLK _53166_/Y _85685_/Q sky130_fd_sc_hd__dfxtp_4
X_82897_ _82896_/CLK _78189_/B _82897_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_666_0_CLK clkbuf_9_333_0_CLK/X _88208_/CLK sky130_fd_sc_hd__clkbuf_1
X_56604_ _56602_/X _56604_/B _56696_/B _56604_/Y sky130_fd_sc_hd__nor3_4
X_87424_ _86814_/CLK _87424_/D _87424_/Q sky130_fd_sc_hd__dfxtp_4
X_53816_ _53846_/A _53816_/X sky130_fd_sc_hd__buf_2
X_41830_ _41824_/X _41825_/X _40459_/X _88132_/Q _41821_/X _41830_/Y
+ sky130_fd_sc_hd__o32ai_4
X_72650_ _72656_/A _72656_/B _56597_/X _72650_/Y sky130_fd_sc_hd__nand3_4
X_84636_ _83216_/CLK _60316_/Y _79742_/A sky130_fd_sc_hd__dfxtp_4
X_57584_ _57564_/X _53552_/B _57584_/Y sky130_fd_sc_hd__nand2_4
X_81848_ _81928_/CLK _81880_/Q _77551_/A sky130_fd_sc_hd__dfxtp_4
X_54796_ _54790_/A _47536_/A _54796_/Y sky130_fd_sc_hd__nand2_4
X_71601_ _71581_/A _83442_/Q _71600_/Y _71601_/X sky130_fd_sc_hd__a21o_4
X_59323_ _59320_/Y _59322_/Y _59278_/X _59323_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_9_157_0_CLK clkbuf_8_78_0_CLK/X clkbuf_9_157_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_56535_ _46187_/A _56535_/X sky130_fd_sc_hd__buf_2
X_41761_ _41603_/X _82888_/Q _41760_/X _41761_/X sky130_fd_sc_hd__o21a_4
X_87355_ _81182_/CLK _87355_/D _87355_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_2_0_2_CLK clkbuf_2_0_2_CLK/A clkbuf_2_0_2_CLK/X sky130_fd_sc_hd__clkbuf_1
X_53747_ _53747_/A _53747_/X sky130_fd_sc_hd__buf_2
X_72581_ _72581_/A _72573_/B _79372_/B _72581_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_9_84_0_CLK clkbuf_8_42_0_CLK/X clkbuf_9_84_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_84567_ _84562_/CLK _84567_/D _60789_/C sky130_fd_sc_hd__dfxtp_4
X_50959_ _50963_/A _50963_/B _50963_/C _46744_/X _50959_/X sky130_fd_sc_hd__and4_4
X_81779_ _88121_/CLK _76100_/X _81779_/Q sky130_fd_sc_hd__dfxtp_4
X_43500_ _41741_/X _43498_/X _87390_/Q _43499_/X _87390_/D sky130_fd_sc_hd__a2bb2o_4
X_74320_ _70304_/C _74314_/X _74319_/Y _83100_/D sky130_fd_sc_hd__a21bo_4
X_86306_ _86303_/CLK _49885_/Y _58135_/B sky130_fd_sc_hd__dfxtp_4
X_40712_ _40712_/A _40712_/X sky130_fd_sc_hd__buf_2
X_59254_ _58697_/A _59255_/A sky130_fd_sc_hd__buf_2
X_71532_ _71527_/Y _71602_/C sky130_fd_sc_hd__buf_2
X_83518_ _83521_/CLK _71384_/X _83518_/Q sky130_fd_sc_hd__dfxtp_4
X_56466_ _56462_/X _55987_/X _56465_/Y _85185_/D sky130_fd_sc_hd__o21ai_4
X_44480_ _41203_/A _44474_/X _87086_/Q _44475_/X _44480_/X sky130_fd_sc_hd__a2bb2o_4
X_87286_ _87542_/CLK _43747_/X _73487_/A sky130_fd_sc_hd__dfxtp_4
X_53678_ _53662_/X _53678_/B _53678_/Y sky130_fd_sc_hd__nand2_4
X_41692_ _41659_/X _81750_/Q _41691_/X _41692_/Y sky130_fd_sc_hd__o21ai_4
X_84498_ _84498_/CLK _84498_/D _61250_/C sky130_fd_sc_hd__dfxtp_4
X_58205_ _64534_/C _58207_/A sky130_fd_sc_hd__buf_2
XPHY_310 sky130_fd_sc_hd__decap_3
X_55417_ _55417_/A _55417_/Y sky130_fd_sc_hd__inv_2
X_43431_ _43396_/A _43431_/X sky130_fd_sc_hd__buf_2
X_74251_ _74038_/A _66334_/B _74251_/X sky130_fd_sc_hd__and2_4
X_86237_ _86237_/CLK _50259_/Y _86237_/Q sky130_fd_sc_hd__dfxtp_4
X_40643_ _40643_/A _40643_/Y sky130_fd_sc_hd__inv_2
XPHY_321 sky130_fd_sc_hd__decap_3
X_52629_ _52515_/X _52629_/X sky130_fd_sc_hd__buf_2
X_59185_ _59105_/X _85746_/Q _59106_/X _59185_/X sky130_fd_sc_hd__o21a_4
X_71463_ _71463_/A _71463_/Y sky130_fd_sc_hd__inv_2
X_83449_ _83480_/CLK _83449_/D _83449_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_332 sky130_fd_sc_hd__decap_3
X_56397_ _56435_/A _56397_/X sky130_fd_sc_hd__buf_2
XPHY_343 sky130_fd_sc_hd__decap_3
XPHY_354 sky130_fd_sc_hd__decap_3
X_73202_ _73704_/A _73202_/X sky130_fd_sc_hd__buf_2
X_46150_ _46144_/X _46150_/B _46149_/Y _86771_/D sky130_fd_sc_hd__and3_4
X_58136_ _58136_/A _58136_/B _58136_/Y sky130_fd_sc_hd__nor2_4
X_70414_ HASH_ADDR[4] _70700_/B sky130_fd_sc_hd__buf_2
XPHY_365 sky130_fd_sc_hd__decap_3
X_43362_ _41371_/X _43356_/X _87459_/Q _43357_/X _43362_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_9_99_0_CLK clkbuf_9_99_0_CLK/A clkbuf_9_99_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_55348_ _55344_/X _55347_/X _55309_/X _55352_/A sky130_fd_sc_hd__a21o_4
X_74182_ _74202_/A _74181_/Y _74182_/Y sky130_fd_sc_hd__nor2_4
X_86168_ _85562_/CLK _50611_/Y _86168_/Q sky130_fd_sc_hd__dfxtp_4
X_40574_ _40550_/X _40556_/X _40573_/X _88370_/Q _40568_/X _40574_/Y
+ sky130_fd_sc_hd__o32ai_4
XPHY_376 sky130_fd_sc_hd__decap_3
X_71394_ _71372_/Y _83514_/Q _71393_/Y _71394_/X sky130_fd_sc_hd__a21o_4
XPHY_387 sky130_fd_sc_hd__decap_3
X_45101_ _85268_/Q _45073_/X _45100_/X _45101_/Y sky130_fd_sc_hd__o21ai_4
XPHY_398 sky130_fd_sc_hd__decap_3
Xclkbuf_10_604_0_CLK clkbuf_9_302_0_CLK/X _81975_/CLK sky130_fd_sc_hd__clkbuf_1
X_42313_ _42307_/X _42297_/X _41616_/X _87926_/Q _42298_/X _42314_/A
+ sky130_fd_sc_hd__o32ai_4
X_73133_ _73062_/X _86195_/Q _72955_/X _73132_/X _73133_/X sky130_fd_sc_hd__a211o_4
X_85119_ _85152_/CLK _85119_/D _85119_/Q sky130_fd_sc_hd__dfxtp_4
X_58067_ _58043_/X _85992_/Q _58066_/X _58067_/Y sky130_fd_sc_hd__o21ai_4
X_70345_ _70337_/X _74769_/A _70344_/X _70345_/X sky130_fd_sc_hd__a21o_4
X_46081_ _46067_/X _43046_/A _41620_/X _67296_/B _46068_/X _46082_/A
+ sky130_fd_sc_hd__o32ai_4
X_43293_ _41179_/X _43287_/X _87494_/Q _43288_/X _87494_/D sky130_fd_sc_hd__a2bb2o_4
X_55279_ _57058_/B _55126_/X _55134_/X _55278_/Y _55279_/X sky130_fd_sc_hd__a211o_4
X_78990_ _78976_/Y _78978_/B _78966_/A _82516_/D _78990_/X sky130_fd_sc_hd__a2bb2o_4
X_86099_ _86100_/CLK _50964_/Y _86099_/Q sky130_fd_sc_hd__dfxtp_4
X_45032_ _83033_/Q _74564_/C sky130_fd_sc_hd__inv_2
X_57018_ _56782_/X _56785_/B _56785_/D _57024_/D _56767_/X _57019_/C
+ sky130_fd_sc_hd__a41o_4
X_42244_ _42276_/A _42244_/X sky130_fd_sc_hd__buf_2
X_73064_ _73062_/X _86198_/Q _72955_/X _73063_/X _73064_/X sky130_fd_sc_hd__a211o_4
X_77941_ _77941_/A _77940_/Y _77942_/B sky130_fd_sc_hd__xnor2_4
X_70276_ _70269_/X _74781_/A _70275_/X _70276_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_9_22_0_CLK clkbuf_9_23_0_CLK/A clkbuf_9_22_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_72015_ _72013_/Y _72009_/X _72014_/Y _72015_/Y sky130_fd_sc_hd__a21boi_4
X_49840_ _49838_/Y _49815_/X _49839_/X _86314_/D sky130_fd_sc_hd__a21oi_4
X_42175_ _42175_/A _42175_/Y sky130_fd_sc_hd__inv_2
X_77872_ _82242_/Q _77872_/B _77872_/Y sky130_fd_sc_hd__xnor2_4
Xclkbuf_10_619_0_CLK clkbuf_9_309_0_CLK/X _82317_/CLK sky130_fd_sc_hd__clkbuf_1
X_79611_ _79611_/A _79611_/B _79611_/Y sky130_fd_sc_hd__nand2_4
X_41126_ _41112_/X _41113_/X _41125_/X _88273_/Q _41088_/X _41127_/A
+ sky130_fd_sc_hd__o32ai_4
X_76823_ _76818_/A _76818_/B _76823_/X sky130_fd_sc_hd__or2_4
X_49771_ _57891_/B _49768_/X _49770_/Y _49771_/Y sky130_fd_sc_hd__o21ai_4
X_46983_ _46983_/A _54478_/B sky130_fd_sc_hd__inv_2
X_58969_ _84785_/Q _58970_/A sky130_fd_sc_hd__inv_2
X_48722_ _65455_/B _48150_/X _48721_/Y _48722_/Y sky130_fd_sc_hd__o21ai_4
X_79542_ _79542_/A _79542_/Y sky130_fd_sc_hd__inv_2
X_45934_ _45890_/X _44228_/X _45933_/Y _45935_/A sky130_fd_sc_hd__and3_4
X_41057_ _41057_/A _41091_/B _41057_/X sky130_fd_sc_hd__or2_4
Xclkbuf_9_37_0_CLK clkbuf_9_37_0_CLK/A clkbuf_9_37_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_76754_ _81486_/Q _76768_/A sky130_fd_sc_hd__inv_2
X_61980_ _61980_/A _63562_/A sky130_fd_sc_hd__inv_2
X_73966_ _43641_/Y _73872_/X _73894_/X _73965_/Y _73966_/X sky130_fd_sc_hd__a211o_4
X_75705_ _81008_/Q _75705_/B _80976_/D sky130_fd_sc_hd__xor2_4
X_48653_ _48653_/A _48654_/A sky130_fd_sc_hd__inv_2
X_60931_ _60826_/A _60838_/X _60931_/C _60931_/Y sky130_fd_sc_hd__nor3_4
X_72917_ _74389_/B _72917_/B _72917_/X sky130_fd_sc_hd__xor2_4
X_79473_ _84813_/Q _84133_/Q _79473_/Y sky130_fd_sc_hd__nand2_4
X_45865_ _45819_/X _61685_/A _45836_/X _45865_/Y sky130_fd_sc_hd__o21ai_4
X_76685_ _76969_/A _76686_/A _76685_/Y sky130_fd_sc_hd__nand2_4
X_73897_ _73893_/X _73896_/X _73799_/X _73913_/B sky130_fd_sc_hd__a21o_4
X_47604_ _47792_/A _47645_/B sky130_fd_sc_hd__buf_2
X_78424_ _78422_/X _78423_/Y _78450_/C sky130_fd_sc_hd__nand2_4
X_44816_ _44816_/A _44816_/Y sky130_fd_sc_hd__inv_2
X_75636_ _80906_/Q _75638_/A sky130_fd_sc_hd__inv_2
X_63650_ _58970_/A _60667_/A _60724_/A _62557_/Y _60671_/B _63650_/Y
+ sky130_fd_sc_hd__o32ai_4
X_48584_ _86509_/Q _48536_/X _48583_/Y _48584_/Y sky130_fd_sc_hd__o21ai_4
X_60862_ _61293_/A _60861_/X _60863_/A sky130_fd_sc_hd__and2_4
X_72848_ _72846_/X _72848_/B _72835_/X _72848_/Y sky130_fd_sc_hd__nand3_4
X_45796_ _57349_/B _44933_/X _45795_/X _45796_/Y sky130_fd_sc_hd__o21ai_4
X_62601_ _62623_/A _62151_/X _62601_/C _62623_/D _62601_/X sky130_fd_sc_hd__and4_4
X_47535_ _47535_/A _47536_/A sky130_fd_sc_hd__inv_2
X_78355_ _78356_/B _78355_/Y sky130_fd_sc_hd__inv_2
X_44747_ _44747_/A _44747_/Y sky130_fd_sc_hd__inv_2
X_63581_ _63413_/A _63581_/X sky130_fd_sc_hd__buf_2
X_75567_ _75567_/A _75567_/B _80769_/D sky130_fd_sc_hd__nand2_4
X_41959_ _40716_/X _41907_/X _74095_/A _41912_/X _88092_/D sky130_fd_sc_hd__a2bb2o_4
X_60793_ _60772_/Y _60791_/X _60749_/Y _60781_/Y _60792_/Y _84566_/D
+ sky130_fd_sc_hd__a41oi_4
X_72779_ _72929_/A _65439_/B _72779_/X sky130_fd_sc_hd__and2_4
X_65320_ _64704_/X _83286_/Q _64980_/X _65319_/X _65320_/X sky130_fd_sc_hd__a211o_4
X_77306_ _77305_/A _82132_/Q _77307_/A sky130_fd_sc_hd__nand2_4
X_62532_ _62532_/A _62532_/X sky130_fd_sc_hd__buf_2
X_74518_ _70368_/X _74518_/B _70880_/C _74518_/D _74518_/Y sky130_fd_sc_hd__nand4_4
X_47466_ _47437_/X _47463_/X _47466_/C _53063_/D _47466_/X sky130_fd_sc_hd__and4_4
X_78286_ _78279_/X _78286_/B _78287_/B sky130_fd_sc_hd__xor2_4
X_44678_ _44677_/Y _44678_/Y sky130_fd_sc_hd__inv_2
X_75498_ _75498_/A _75495_/Y _75497_/Y _75503_/A sky130_fd_sc_hd__or3_4
X_49205_ _49205_/A _49232_/A sky130_fd_sc_hd__buf_2
X_46417_ _46408_/A _46417_/B _46417_/Y sky130_fd_sc_hd__nand2_4
X_65251_ _65248_/X _65250_/X _65122_/X _65255_/A sky130_fd_sc_hd__a21o_4
X_77237_ _77236_/A _82083_/D _77239_/C sky130_fd_sc_hd__nand2_4
X_43629_ _43628_/X _87335_/D sky130_fd_sc_hd__inv_2
X_62463_ _62463_/A _62463_/X sky130_fd_sc_hd__buf_2
X_74449_ _46347_/A _52188_/B _74449_/Y sky130_fd_sc_hd__nand2_4
X_47397_ _86639_/Q _47382_/X _47396_/Y _47397_/Y sky130_fd_sc_hd__o21ai_4
X_64202_ _59450_/Y _61086_/X _64202_/Y sky130_fd_sc_hd__nor2_4
X_49136_ _49117_/A _49135_/X _49136_/Y sky130_fd_sc_hd__nand2_4
X_61414_ _61414_/A _61434_/B sky130_fd_sc_hd__buf_2
X_46348_ _46348_/A _46348_/X sky130_fd_sc_hd__buf_2
X_65182_ _64902_/A _65182_/X sky130_fd_sc_hd__buf_2
X_77168_ _82105_/Q _77168_/B _77168_/X sky130_fd_sc_hd__xor2_4
X_62394_ _62385_/X _62389_/Y _62393_/X _84741_/Q _62367_/X _62394_/Y
+ sky130_fd_sc_hd__o32ai_4
X_64133_ _59430_/Y _61003_/Y _62129_/X _60962_/Y _64133_/X sky130_fd_sc_hd__a2bb2o_4
X_76119_ _76112_/B _76112_/A _76118_/Y _76119_/Y sky130_fd_sc_hd__a21boi_4
X_61345_ _61344_/Y _61345_/Y sky130_fd_sc_hd__inv_2
X_49067_ _48976_/A _49067_/B _49067_/Y sky130_fd_sc_hd__nand2_4
X_46279_ _46279_/A _46279_/X sky130_fd_sc_hd__buf_2
X_69990_ _69943_/X _68446_/Y _69984_/X _69989_/Y _69990_/X sky130_fd_sc_hd__a211o_4
X_77099_ _77098_/A _82287_/D _77099_/Y sky130_fd_sc_hd__nand2_4
X_48018_ _48018_/A _47973_/B _48018_/X sky130_fd_sc_hd__or2_4
X_68941_ _68987_/A _68941_/B _68941_/X sky130_fd_sc_hd__and2_4
X_64064_ _64058_/Y _64059_/Y _64064_/C _64064_/D _64064_/X sky130_fd_sc_hd__and4_4
X_61276_ _72625_/B _61276_/B _60402_/A _61287_/A _61278_/A sky130_fd_sc_hd__and4_4
X_63015_ _60410_/B _63342_/C sky130_fd_sc_hd__buf_2
X_60227_ _60227_/A _60228_/A sky130_fd_sc_hd__buf_2
X_68872_ _68759_/A _87231_/Q _68872_/X sky130_fd_sc_hd__and2_4
X_67823_ _87391_/Q _67751_/X _67821_/X _67822_/X _67823_/X sky130_fd_sc_hd__a211o_4
X_79809_ _79786_/X _79799_/X _79809_/Y sky130_fd_sc_hd__nand2_4
X_60158_ _60251_/A _60159_/A sky130_fd_sc_hd__buf_2
X_49969_ _49973_/A _49973_/B _49973_/C _53181_/D _49969_/X sky130_fd_sc_hd__and4_4
X_82820_ _82820_/CLK _82820_/D _82820_/Q sky130_fd_sc_hd__dfxtp_4
X_67754_ _67750_/X _67753_/X _67681_/X _67754_/X sky130_fd_sc_hd__a21o_4
X_52980_ _85719_/Q _52957_/X _52979_/Y _52980_/Y sky130_fd_sc_hd__o21ai_4
X_64966_ _60151_/X _64953_/Y _64965_/Y _64966_/Y sky130_fd_sc_hd__o21ai_4
X_60089_ _60081_/A _60103_/B _60089_/C _60089_/Y sky130_fd_sc_hd__nor3_4
X_66705_ _88398_/Q _66633_/X _66682_/X _66704_/X _66705_/X sky130_fd_sc_hd__a211o_4
X_51931_ _53199_/A _53259_/A sky130_fd_sc_hd__buf_2
X_63917_ _60996_/B _63949_/C sky130_fd_sc_hd__buf_2
X_82751_ _84115_/CLK _84135_/Q _82751_/Q sky130_fd_sc_hd__dfxtp_4
X_67685_ _67682_/X _67684_/X _67637_/X _67685_/Y sky130_fd_sc_hd__a21oi_4
X_64897_ _64894_/X _64896_/X _64701_/X _64897_/X sky130_fd_sc_hd__a21o_4
X_81702_ _82053_/CLK _81702_/D _81702_/Q sky130_fd_sc_hd__dfxtp_4
X_69424_ _69162_/A _69424_/X sky130_fd_sc_hd__buf_2
X_54650_ _54649_/X _54125_/B _54650_/Y sky130_fd_sc_hd__nand2_4
X_66636_ _66632_/X _66635_/X _66366_/A _66636_/Y sky130_fd_sc_hd__a21oi_4
X_85470_ _82206_/CLK _54287_/Y _85470_/Q sky130_fd_sc_hd__dfxtp_4
X_51862_ _51853_/A _50998_/B _51862_/Y sky130_fd_sc_hd__nand2_4
X_63848_ _63644_/A _63848_/X sky130_fd_sc_hd__buf_2
X_82682_ _81190_/CLK _82694_/Q _82682_/Q sky130_fd_sc_hd__dfxtp_4
X_53601_ _53601_/A _57637_/B _53601_/Y sky130_fd_sc_hd__nand2_4
X_84421_ _84421_/CLK _62284_/Y _84421_/Q sky130_fd_sc_hd__dfxtp_4
X_50813_ _50811_/Y _50801_/X _50812_/X _50813_/Y sky130_fd_sc_hd__a21oi_4
X_81633_ _81695_/CLK _76643_/A _81825_/D sky130_fd_sc_hd__dfxtp_4
X_69355_ _88035_/Q _69121_/X _69232_/X _69354_/X _69355_/X sky130_fd_sc_hd__a211o_4
X_54581_ _54579_/Y _54558_/X _54580_/X _54581_/Y sky130_fd_sc_hd__a21oi_4
X_66567_ _69454_/A _66567_/B _66567_/X sky130_fd_sc_hd__and2_4
X_51793_ _51793_/A _51793_/X sky130_fd_sc_hd__buf_2
X_63779_ _63772_/Y _63775_/Y _63777_/Y _63779_/D _63779_/X sky130_fd_sc_hd__and4_4
X_56320_ _56070_/X _56305_/X _56319_/Y _85237_/D sky130_fd_sc_hd__o21ai_4
X_68306_ _68272_/X _67862_/Y _68287_/X _68305_/Y _68306_/X sky130_fd_sc_hd__a211o_4
X_87140_ _88220_/CLK _87140_/D _87140_/Q sky130_fd_sc_hd__dfxtp_4
X_53532_ _85618_/Q _53466_/X _53531_/Y _53532_/Y sky130_fd_sc_hd__o21ai_4
X_65518_ _65791_/A _65777_/A sky130_fd_sc_hd__buf_2
X_84352_ _83227_/CLK _84352_/D _79414_/A sky130_fd_sc_hd__dfxtp_4
X_50744_ _50771_/A _50744_/B _50744_/Y sky130_fd_sc_hd__nand2_4
X_81564_ _84064_/CLK _76891_/X _81564_/Q sky130_fd_sc_hd__dfxtp_4
X_69286_ _69286_/A _87784_/Q _69286_/X sky130_fd_sc_hd__and2_4
X_66498_ _68823_/A _66499_/B sky130_fd_sc_hd__buf_2
X_83303_ _83303_/CLK _72011_/Y _83303_/Q sky130_fd_sc_hd__dfxtp_4
X_80515_ _80505_/X _80506_/X _80514_/Y _80531_/A sky130_fd_sc_hd__a21boi_4
X_56251_ _56130_/X _56242_/X _56250_/Y _85259_/D sky130_fd_sc_hd__o21ai_4
X_68237_ _82652_/D _68220_/X _68236_/X _68237_/X sky130_fd_sc_hd__a21bo_4
X_87071_ _83115_/CLK _87071_/D _44514_/A sky130_fd_sc_hd__dfxtp_4
X_53463_ _53461_/Y _53455_/X _53462_/Y _53463_/Y sky130_fd_sc_hd__a21boi_4
X_65449_ _65449_/A _65294_/B _65449_/C _65449_/X sky130_fd_sc_hd__and3_4
X_84283_ _84668_/CLK _63977_/Y _80102_/B sky130_fd_sc_hd__dfxtp_4
X_50675_ _86155_/Q _50654_/X _50674_/Y _50675_/Y sky130_fd_sc_hd__o21ai_4
X_81495_ _81431_/CLK _84063_/Q _76839_/A sky130_fd_sc_hd__dfxtp_4
X_55202_ _55710_/B _45823_/Y _55202_/Y sky130_fd_sc_hd__nor2_4
X_86022_ _86118_/CLK _86022_/D _86022_/Q sky130_fd_sc_hd__dfxtp_4
X_52414_ _65384_/B _52397_/X _52413_/Y _52414_/Y sky130_fd_sc_hd__o21ai_4
X_83234_ _84350_/CLK _72560_/Y _79436_/B sky130_fd_sc_hd__dfxtp_4
X_56182_ _56181_/X _56182_/X sky130_fd_sc_hd__buf_2
X_80446_ _80435_/X _80446_/B _80446_/X sky130_fd_sc_hd__and2_4
X_68168_ _68168_/A _68168_/X sky130_fd_sc_hd__buf_2
X_53394_ _53391_/Y _53382_/X _53393_/X _53394_/Y sky130_fd_sc_hd__a21oi_4
X_67119_ _87932_/Q _67117_/X _67046_/X _67118_/X _67119_/X sky130_fd_sc_hd__a211o_4
X_55133_ _55133_/A _55133_/X sky130_fd_sc_hd__buf_2
X_52345_ _50645_/A _50645_/B _52280_/X _52345_/X sky130_fd_sc_hd__o21a_4
X_83165_ _86570_/CLK _73103_/X _83165_/Q sky130_fd_sc_hd__dfxtp_4
X_80377_ _59291_/Y _66264_/C _80376_/Y _80394_/A sky130_fd_sc_hd__o21a_4
X_68099_ _68097_/X _66623_/Y _68089_/X _68098_/Y _68099_/X sky130_fd_sc_hd__a211o_4
X_70130_ _70130_/A _70130_/B _70131_/C sky130_fd_sc_hd__nor2_4
X_82116_ _82116_/CLK _82116_/D _82116_/Q sky130_fd_sc_hd__dfxtp_4
X_55064_ _85325_/Q _55046_/X _55063_/Y _55064_/Y sky130_fd_sc_hd__o21ai_4
X_59941_ _62288_/A _62504_/A sky130_fd_sc_hd__buf_2
X_52276_ _52273_/Y _52262_/X _52275_/X _85855_/D sky130_fd_sc_hd__a21oi_4
X_87973_ _87149_/CLK _87973_/D _87973_/Q sky130_fd_sc_hd__dfxtp_4
X_83096_ _83846_/CLK _83096_/D _70315_/C sky130_fd_sc_hd__dfxtp_4
X_54015_ _53773_/A _54015_/X sky130_fd_sc_hd__buf_2
X_51227_ _51212_/A _52918_/B _51227_/Y sky130_fd_sc_hd__nand2_4
X_70061_ _69855_/Y _59834_/A _70056_/X _70060_/Y _70061_/X sky130_fd_sc_hd__a211o_4
X_86924_ _87652_/CLK _86924_/D _86924_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_590_0_CLK clkbuf_9_295_0_CLK/X _83957_/CLK sky130_fd_sc_hd__clkbuf_1
X_82047_ _82047_/CLK _78003_/Y _82015_/D sky130_fd_sc_hd__dfxtp_4
X_59872_ _59852_/A _59873_/B sky130_fd_sc_hd__buf_2
X_58823_ _58813_/X _85773_/Q _58706_/X _58823_/X sky130_fd_sc_hd__o21a_4
X_51158_ _51167_/A _52850_/B _51158_/Y sky130_fd_sc_hd__nand2_4
X_86855_ _86855_/CLK _86855_/D _62094_/D sky130_fd_sc_hd__dfxtp_4
X_50109_ _86262_/Q _50088_/X _50108_/Y _50109_/Y sky130_fd_sc_hd__o21ai_4
X_73820_ _73820_/A _73624_/X _73820_/Y sky130_fd_sc_hd__nor2_4
X_85806_ _86040_/CLK _52521_/Y _65103_/B sky130_fd_sc_hd__dfxtp_4
X_58754_ _58738_/Y _58739_/X _58745_/X _58753_/X _84803_/D sky130_fd_sc_hd__a22oi_4
X_51089_ _51084_/A _51071_/B _51110_/C _52779_/D _51089_/X sky130_fd_sc_hd__and4_4
X_55966_ _55966_/A _55966_/X sky130_fd_sc_hd__buf_2
X_43980_ _86840_/Q _43987_/B _43955_/Y _43979_/Y _59899_/D sky130_fd_sc_hd__a211o_4
X_86786_ _86784_/CLK _86786_/D _67049_/B sky130_fd_sc_hd__dfxtp_4
X_83998_ _82642_/CLK _68263_/X _83998_/Q sky130_fd_sc_hd__dfxtp_4
X_57705_ _44181_/X _57705_/X sky130_fd_sc_hd__buf_2
X_54917_ _54913_/Y _54909_/X _54916_/X _85354_/D sky130_fd_sc_hd__a21oi_4
X_42931_ _42951_/A _42931_/X sky130_fd_sc_hd__buf_2
X_73751_ _41914_/Y _73529_/X _73698_/X _73750_/Y _73751_/X sky130_fd_sc_hd__a211o_4
X_85737_ _85738_/CLK _52884_/Y _85737_/Q sky130_fd_sc_hd__dfxtp_4
X_70963_ _49245_/B _70961_/X _70962_/Y _70963_/Y sky130_fd_sc_hd__o21ai_4
X_58685_ _58681_/Y _58684_/Y _58610_/X _58685_/X sky130_fd_sc_hd__a21o_4
X_82949_ _86697_/CLK _82757_/Q _82949_/Q sky130_fd_sc_hd__dfxtp_4
X_55897_ _85207_/Q _44070_/B _55627_/X _55896_/X _55897_/X sky130_fd_sc_hd__a211o_4
X_72702_ _72686_/A _72702_/X sky130_fd_sc_hd__buf_2
X_45650_ _45646_/X _45649_/X _45602_/X _45650_/X sky130_fd_sc_hd__a21o_4
X_57636_ _72017_/A _71972_/A sky130_fd_sc_hd__buf_2
X_76470_ _76470_/A _76474_/A sky130_fd_sc_hd__inv_2
X_42862_ _41556_/X _42852_/X _87681_/Q _42853_/X _42862_/X sky130_fd_sc_hd__a2bb2o_4
X_54848_ _54857_/A _54857_/B _54857_/C _53155_/D _54848_/X sky130_fd_sc_hd__and4_4
X_73682_ _87002_/Q _56550_/X _73681_/X _73694_/C sky130_fd_sc_hd__o21ai_4
X_85668_ _85471_/CLK _85668_/D _85668_/Q sky130_fd_sc_hd__dfxtp_4
X_70894_ _50981_/B _70885_/X _70893_/Y _70894_/Y sky130_fd_sc_hd__o21ai_4
X_44601_ _44593_/X _44594_/X _40929_/A _44600_/Y _44596_/X _44601_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75421_ _75419_/X _75420_/Y _75421_/X sky130_fd_sc_hd__xor2_4
X_87407_ _87472_/CLK _87407_/D _87407_/Q sky130_fd_sc_hd__dfxtp_4
X_41813_ _48164_/A _41813_/X sky130_fd_sc_hd__buf_2
X_72633_ _72687_/A _72633_/X sky130_fd_sc_hd__buf_2
X_84619_ _84590_/CLK _60373_/X _79538_/A sky130_fd_sc_hd__dfxtp_4
X_57567_ _57567_/A _49317_/X _46603_/X _57567_/X sky130_fd_sc_hd__and3_4
X_45581_ _85077_/Q _45581_/Y sky130_fd_sc_hd__inv_2
X_88387_ _88387_/CLK _40470_/X _88387_/Q sky130_fd_sc_hd__dfxtp_4
X_42793_ _42774_/X _42775_/X _41376_/X _87714_/Q _42781_/X _42794_/A
+ sky130_fd_sc_hd__o32ai_4
X_54779_ _54807_/A _54798_/A sky130_fd_sc_hd__buf_2
X_85599_ _85599_/CLK _53632_/Y _85599_/Q sky130_fd_sc_hd__dfxtp_4
X_59306_ _86664_/Q _59306_/B _59306_/Y sky130_fd_sc_hd__nor2_4
X_47320_ _47320_/A _52982_/D sky130_fd_sc_hd__buf_2
X_78140_ _82571_/Q _82483_/Q _78143_/A sky130_fd_sc_hd__xor2_4
X_44532_ _44532_/A _44533_/A sky130_fd_sc_hd__buf_2
X_56518_ _56523_/A _56520_/B _56518_/C _56518_/Y sky130_fd_sc_hd__nand3_4
X_75352_ _75348_/Y _75349_/Y _75351_/Y _75354_/A sky130_fd_sc_hd__or3_4
X_87338_ _86988_/CLK _43622_/Y _87338_/Q sky130_fd_sc_hd__dfxtp_4
X_41744_ _41577_/X _82891_/Q _41743_/X _41744_/Y sky130_fd_sc_hd__o21ai_4
X_72564_ _72564_/A _72573_/B sky130_fd_sc_hd__buf_2
X_57498_ _57496_/Y _46576_/X _57497_/Y _84992_/D sky130_fd_sc_hd__a21boi_4
X_74303_ _74342_/A _74310_/B sky130_fd_sc_hd__buf_2
X_47251_ _83390_/Q _54106_/B sky130_fd_sc_hd__inv_2
X_59237_ _58864_/A _59237_/X sky130_fd_sc_hd__buf_2
X_71515_ _71521_/A _70714_/A _71515_/Y sky130_fd_sc_hd__nand2_4
X_78071_ _60746_/C _78071_/B _78071_/X sky130_fd_sc_hd__xor2_4
X_44463_ _41151_/A _44453_/X _87096_/Q _44454_/X _87096_/D sky130_fd_sc_hd__a2bb2o_4
X_56449_ _56448_/X _56454_/B sky130_fd_sc_hd__buf_2
X_75283_ _75248_/Y _75279_/Y _75282_/Y _75283_/Y sky130_fd_sc_hd__a21oi_4
X_41675_ _41628_/X _41326_/A _41674_/X _41675_/X sky130_fd_sc_hd__o21a_4
X_87269_ _87525_/CLK _87269_/D _69332_/B sky130_fd_sc_hd__dfxtp_4
X_72495_ _72484_/X _83381_/Q _72494_/Y _72495_/X sky130_fd_sc_hd__o21a_4
X_46202_ _58425_/A _58273_/A sky130_fd_sc_hd__buf_2
XPHY_140 sky130_fd_sc_hd__decap_3
X_77022_ _82085_/Q _77022_/B _82366_/D sky130_fd_sc_hd__xor2_4
X_43414_ _41511_/X _43412_/X _87433_/Q _43413_/X _87433_/D sky130_fd_sc_hd__a2bb2o_4
X_74234_ _73165_/A _74234_/B _74234_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_543_0_CLK clkbuf_9_271_0_CLK/X _80928_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_151 sky130_fd_sc_hd__decap_3
X_40626_ _40625_/Y _40626_/X sky130_fd_sc_hd__buf_2
X_59168_ _86676_/Q _59189_/B _59168_/Y sky130_fd_sc_hd__nor2_4
X_47182_ _47176_/Y _47177_/X _47181_/X _47182_/Y sky130_fd_sc_hd__a21oi_4
X_71446_ _71238_/B _71446_/X sky130_fd_sc_hd__buf_2
Xclkbuf_6_34_0_CLK clkbuf_6_35_0_CLK/A clkbuf_7_69_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_44394_ _44363_/X _44394_/X sky130_fd_sc_hd__buf_2
XPHY_162 sky130_fd_sc_hd__decap_3
XPHY_173 sky130_fd_sc_hd__decap_3
XPHY_184 sky130_fd_sc_hd__decap_3
X_46133_ _46133_/A _46133_/B _46133_/C _46207_/B _46134_/A sky130_fd_sc_hd__and4_4
X_58119_ _58108_/Y _57981_/X _58115_/X _58118_/X _84924_/D sky130_fd_sc_hd__a22oi_4
XPHY_195 sky130_fd_sc_hd__decap_3
X_43345_ _43344_/Y _87468_/D sky130_fd_sc_hd__inv_2
X_74165_ _41966_/Y _73930_/X _73551_/X _74164_/Y _74165_/X sky130_fd_sc_hd__a211o_4
X_40557_ _48135_/A _48606_/A sky130_fd_sc_hd__buf_2
X_59099_ _59061_/X _86073_/Q _59098_/X _59099_/Y sky130_fd_sc_hd__o21ai_4
X_71377_ _70670_/A _71377_/B _71377_/C _71377_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_opt_2_CLK _83246_/CLK _84894_/CLK sky130_fd_sc_hd__clkbuf_16
X_61130_ _64523_/B _61202_/B sky130_fd_sc_hd__buf_2
X_73116_ _73113_/X _73115_/X _72739_/X _73116_/X sky130_fd_sc_hd__a21o_4
X_46064_ _46046_/X _46054_/X _41564_/X _67049_/B _46047_/X _46065_/A
+ sky130_fd_sc_hd__o32ai_4
X_70328_ _70328_/A _70328_/B _70328_/C _70328_/D _70328_/X sky130_fd_sc_hd__and4_4
X_43276_ _41130_/X _43264_/X _87504_/Q _43265_/X _43276_/X sky130_fd_sc_hd__a2bb2o_4
X_74096_ _42518_/Y _73319_/X _73551_/X _74095_/Y _74096_/X sky130_fd_sc_hd__a211o_4
X_78973_ _78957_/B _78970_/X _78972_/Y _78979_/B sky130_fd_sc_hd__a21oi_4
X_40488_ _44382_/A _40488_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_558_0_CLK clkbuf_9_279_0_CLK/X _87408_/CLK sky130_fd_sc_hd__clkbuf_1
X_45015_ _85178_/Q _44982_/X _44959_/X _45015_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_6_49_0_CLK clkbuf_6_49_0_CLK/A clkbuf_7_98_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_42227_ _41881_/A _42276_/A sky130_fd_sc_hd__buf_2
X_73047_ _73044_/X _73046_/X _73048_/B sky130_fd_sc_hd__nand2_4
X_61061_ _60946_/X _61138_/B _76971_/A _61061_/Y sky130_fd_sc_hd__nor3_4
X_77924_ _82167_/Q _82039_/D _82135_/D sky130_fd_sc_hd__xor2_4
X_70259_ _70255_/X _74764_/B _70258_/X _83820_/D sky130_fd_sc_hd__a21o_4
X_60012_ _62515_/C _62548_/D sky130_fd_sc_hd__buf_2
X_49823_ _49830_/A _49830_/B _49830_/C _53036_/D _49823_/X sky130_fd_sc_hd__and4_4
X_42158_ _41189_/X _42148_/X _88005_/Q _42150_/X _88005_/D sky130_fd_sc_hd__a2bb2o_4
X_77855_ _77841_/Y _77854_/X _77855_/Y sky130_fd_sc_hd__nand2_4
X_41109_ _40941_/A _41109_/X sky130_fd_sc_hd__buf_2
X_64820_ _64804_/A _64820_/B _64820_/X sky130_fd_sc_hd__and2_4
X_76806_ _76806_/A _76792_/Y _76806_/Y sky130_fd_sc_hd__nor2_4
X_49754_ _86329_/Q _49742_/X _49753_/Y _49754_/Y sky130_fd_sc_hd__o21ai_4
X_46966_ _46960_/Y _46940_/X _46965_/X _86685_/D sky130_fd_sc_hd__a21oi_4
X_42089_ _42088_/Y _88040_/D sky130_fd_sc_hd__inv_2
X_77786_ _82265_/Q _81977_/Q _77786_/X sky130_fd_sc_hd__xor2_4
X_74998_ _80951_/Q _74998_/B _74998_/X sky130_fd_sc_hd__xor2_4
X_48705_ _48704_/Y _48872_/B sky130_fd_sc_hd__buf_2
X_79525_ _79161_/Y _79525_/B _82818_/D sky130_fd_sc_hd__xnor2_4
X_45917_ _69626_/A _65381_/A sky130_fd_sc_hd__buf_2
X_64751_ _64747_/X _64712_/B _64750_/X _64751_/Y sky130_fd_sc_hd__nand3_4
X_76737_ _76725_/A _76732_/A _76737_/X sky130_fd_sc_hd__and2_4
X_49685_ _49685_/A _49669_/B _49685_/C _52900_/D _49685_/X sky130_fd_sc_hd__and4_4
X_61963_ _61962_/X _61945_/X _58533_/A _61947_/D _61963_/X sky130_fd_sc_hd__and4_4
X_73949_ _73949_/A _66141_/B _73949_/X sky130_fd_sc_hd__and2_4
X_46897_ _46889_/Y _46891_/X _46896_/X _46897_/Y sky130_fd_sc_hd__a21oi_4
X_63702_ _63700_/Y _63679_/X _63701_/Y _63702_/Y sky130_fd_sc_hd__a21oi_4
X_48636_ _48841_/A _48657_/B _48657_/C _48636_/X sky130_fd_sc_hd__and3_4
X_60914_ _60909_/X _60865_/B _64081_/C _60910_/B _60988_/A sky130_fd_sc_hd__nand4_4
X_67470_ _67465_/X _67469_/X _67423_/X _67470_/Y sky130_fd_sc_hd__a21oi_4
X_79456_ _79456_/A _79456_/B _79457_/B sky130_fd_sc_hd__xor2_4
X_45848_ _74700_/B _45832_/B _45848_/Y sky130_fd_sc_hd__nand2_4
X_64682_ _64677_/X _64681_/X _64629_/X _64682_/X sky130_fd_sc_hd__a21o_4
X_76668_ _81684_/Q _76667_/Y _76668_/X sky130_fd_sc_hd__or2_4
X_61894_ _61879_/A _61889_/Y _61890_/Y _61893_/Y _61894_/Y sky130_fd_sc_hd__nand4_4
X_66421_ _66418_/Y _66414_/X _66420_/X _84127_/D sky130_fd_sc_hd__a21o_4
X_78407_ _78402_/Y _78407_/Y sky130_fd_sc_hd__inv_2
X_63633_ _58461_/A _63600_/X _63661_/C _63661_/D _63633_/Y sky130_fd_sc_hd__nand4_4
X_75619_ _75619_/A _80776_/D _75632_/A sky130_fd_sc_hd__xnor2_4
X_60845_ _61075_/B _60845_/Y sky130_fd_sc_hd__inv_2
X_48567_ _48567_/A _52194_/A sky130_fd_sc_hd__buf_2
X_79387_ _79387_/A _79386_/Y _79387_/X sky130_fd_sc_hd__xor2_4
X_45779_ _45773_/X _45776_/X _45778_/Y _86855_/D sky130_fd_sc_hd__a21oi_4
X_76599_ _76572_/Y _76576_/B _76574_/Y _76599_/X sky130_fd_sc_hd__o21a_4
X_69140_ _69128_/X _88307_/Q _69140_/X sky130_fd_sc_hd__and2_4
X_47518_ _58136_/A _47478_/X _47517_/Y _47518_/Y sky130_fd_sc_hd__o21ai_4
X_66352_ _66348_/X _66351_/X _58882_/A _66352_/X sky130_fd_sc_hd__a21o_4
X_78338_ _78338_/A _78339_/B sky130_fd_sc_hd__inv_2
X_63564_ _63443_/A _63575_/C sky130_fd_sc_hd__buf_2
X_48498_ _48498_/A _52161_/A sky130_fd_sc_hd__buf_2
X_60776_ _60804_/C _70021_/C _60736_/X _60776_/Y sky130_fd_sc_hd__nand3_4
X_65303_ _65300_/X _85510_/Q _65301_/X _65302_/X _65303_/X sky130_fd_sc_hd__a211o_4
X_62515_ _62515_/A _59995_/A _62515_/C _61580_/X _62515_/X sky130_fd_sc_hd__and4_4
X_69071_ _69068_/X _69070_/X _68748_/X _69071_/X sky130_fd_sc_hd__a21o_4
X_47449_ _47445_/Y _47414_/X _47448_/X _86634_/D sky130_fd_sc_hd__a21oi_4
X_66283_ _64826_/A _66283_/B _66283_/X sky130_fd_sc_hd__and2_4
X_78269_ _78262_/X _78268_/Y _78270_/B sky130_fd_sc_hd__xor2_4
X_63495_ _63368_/A _63495_/X sky130_fd_sc_hd__buf_2
X_80300_ _80302_/B _80299_/Y _80300_/Y sky130_fd_sc_hd__nor2_4
X_68022_ _68019_/X _68021_/X _67977_/X _68027_/A sky130_fd_sc_hd__a21o_4
X_65234_ _65155_/A _65234_/B _65234_/X sky130_fd_sc_hd__and2_4
X_50460_ _50460_/A _50496_/A sky130_fd_sc_hd__buf_2
X_62446_ _61528_/A _62472_/B _62490_/C _62431_/D _62446_/Y sky130_fd_sc_hd__nand4_4
X_81280_ _81682_/CLK _81280_/D _76620_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_2_0_CLK clkbuf_8_3_0_CLK/A clkbuf_9_5_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_49119_ _49119_/A _49029_/B _49119_/Y sky130_fd_sc_hd__nor2_4
X_80231_ _84951_/Q _65466_/C _80233_/A sky130_fd_sc_hd__xor2_4
X_65165_ _65065_/X _83292_/Q _65108_/X _65164_/X _65165_/X sky130_fd_sc_hd__a211o_4
X_50391_ _50391_/A _50475_/B _50257_/X _50391_/Y sky130_fd_sc_hd__nand3_4
X_62377_ _61461_/X _62420_/B _62420_/C _62334_/D _62378_/D sky130_fd_sc_hd__nand4_4
X_52130_ _48744_/A _52135_/B _52097_/X _52130_/X sky130_fd_sc_hd__and3_4
X_64116_ _64116_/A _64087_/X _79998_/B _64116_/Y sky130_fd_sc_hd__nor3_4
X_61328_ _72515_/D _61375_/C sky130_fd_sc_hd__buf_2
X_80162_ _80156_/Y _80162_/B _80162_/X sky130_fd_sc_hd__xor2_4
X_65096_ _64948_/A _65096_/B _65096_/X sky130_fd_sc_hd__and2_4
X_69973_ _87040_/Q _66550_/X _66552_/X _69972_/X _69973_/X sky130_fd_sc_hd__a211o_4
X_52061_ _85896_/Q _52013_/X _52060_/Y _52061_/Y sky130_fd_sc_hd__o21ai_4
X_68924_ _68994_/A _68924_/B _68924_/X sky130_fd_sc_hd__and2_4
X_64047_ _64040_/Y _64042_/Y _64044_/Y _64047_/D _64047_/X sky130_fd_sc_hd__and4_4
X_61259_ _61293_/A _61293_/B _72625_/A _61260_/A sky130_fd_sc_hd__and3_4
X_84970_ _84970_/CLK _57610_/Y _84970_/Q sky130_fd_sc_hd__dfxtp_4
X_80093_ _80089_/X _80105_/B _80098_/A sky130_fd_sc_hd__xor2_4
X_51012_ _51012_/A _51013_/A sky130_fd_sc_hd__buf_2
X_83921_ _81507_/CLK _83921_/D _81385_/D sky130_fd_sc_hd__dfxtp_4
X_68855_ _68852_/X _68854_/X _68661_/X _68855_/Y sky130_fd_sc_hd__a21oi_4
X_55820_ _55819_/X _56108_/A sky130_fd_sc_hd__buf_2
X_67806_ _67806_/A _67806_/X sky130_fd_sc_hd__buf_2
X_86640_ _86640_/CLK _86640_/D _86640_/Q sky130_fd_sc_hd__dfxtp_4
X_83852_ _82536_/CLK _70091_/X _83852_/Q sky130_fd_sc_hd__dfxtp_4
X_68786_ _44709_/A _68707_/X _68762_/X _68785_/X _68786_/X sky130_fd_sc_hd__a211o_4
X_65998_ _65824_/X _84987_/Q _65707_/X _65997_/X _65999_/B sky130_fd_sc_hd__a211o_4
X_82803_ _82803_/CLK _82835_/Q _78552_/A sky130_fd_sc_hd__dfxtp_4
X_55751_ _56442_/C _55272_/X _55168_/X _55750_/X _55752_/B sky130_fd_sc_hd__a211o_4
X_67737_ _67690_/X _87650_/Q _67737_/X sky130_fd_sc_hd__and2_4
X_86571_ _85601_/CLK _48070_/Y _74083_/B sky130_fd_sc_hd__dfxtp_4
X_52963_ _52947_/X _52982_/B _52977_/C _52963_/D _52963_/X sky130_fd_sc_hd__and4_4
X_64949_ _64846_/X _85556_/Q _64919_/X _64948_/X _64949_/X sky130_fd_sc_hd__a211o_4
X_83783_ _83783_/CLK _70380_/Y _46545_/A sky130_fd_sc_hd__dfxtp_4
X_80995_ _82610_/CLK _84203_/Q _80995_/Q sky130_fd_sc_hd__dfxtp_4
X_88310_ _87851_/CLK _88310_/D _88310_/Q sky130_fd_sc_hd__dfxtp_4
X_54702_ _54698_/Y _54694_/X _54701_/X _85394_/D sky130_fd_sc_hd__a21oi_4
X_85522_ _86139_/CLK _85522_/D _85522_/Q sky130_fd_sc_hd__dfxtp_4
X_51914_ _51914_/A _51898_/B _51893_/C _52742_/D _51914_/X sky130_fd_sc_hd__and4_4
X_58470_ _63557_/B _58474_/B _58470_/Y sky130_fd_sc_hd__nor2_4
X_82734_ _82147_/CLK _84118_/Q _82734_/Q sky130_fd_sc_hd__dfxtp_4
X_55682_ _55681_/X _55683_/D sky130_fd_sc_hd__inv_2
X_67668_ _87461_/Q _67594_/X _67595_/X _67667_/X _67668_/X sky130_fd_sc_hd__a211o_4
X_52894_ _52893_/X _52895_/A sky130_fd_sc_hd__buf_2
X_57421_ _57440_/A _57445_/B sky130_fd_sc_hd__buf_2
X_69407_ _69300_/X _69403_/Y _69405_/X _69406_/Y _69407_/X sky130_fd_sc_hd__a211o_4
X_88241_ _87408_/CLK _88241_/D _67399_/B sky130_fd_sc_hd__dfxtp_4
X_54633_ _85406_/Q _54621_/X _54632_/Y _54633_/Y sky130_fd_sc_hd__o21ai_4
X_66619_ _87377_/Q _66538_/X _66540_/X _66618_/X _66619_/X sky130_fd_sc_hd__a211o_4
X_85453_ _85773_/CLK _85453_/D _85453_/Q sky130_fd_sc_hd__dfxtp_4
X_51845_ _51841_/Y _51823_/X _51844_/X _51845_/Y sky130_fd_sc_hd__a21oi_4
X_82665_ _82665_/CLK _82709_/Q _78128_/A sky130_fd_sc_hd__dfxtp_4
X_67599_ _67126_/X _67696_/A sky130_fd_sc_hd__buf_2
X_84404_ _84418_/CLK _62528_/Y _62527_/C sky130_fd_sc_hd__dfxtp_4
X_57352_ _57289_/B _56862_/Y _57346_/C _57337_/Y _57352_/X sky130_fd_sc_hd__o22a_4
X_81616_ _81808_/CLK _76363_/B _81808_/D sky130_fd_sc_hd__dfxtp_4
X_69338_ _69329_/X _68725_/Y _69325_/X _69337_/Y _69338_/X sky130_fd_sc_hd__a211o_4
X_88172_ _83987_/CLK _41670_/Y _88172_/Q sky130_fd_sc_hd__dfxtp_4
X_54564_ _54537_/A _54565_/C sky130_fd_sc_hd__buf_2
X_85384_ _85379_/CLK _85384_/D _85384_/Q sky130_fd_sc_hd__dfxtp_4
X_51776_ _51747_/A _51794_/A sky130_fd_sc_hd__buf_2
X_82596_ _82596_/CLK _78831_/B _82564_/D sky130_fd_sc_hd__dfxtp_4
X_56303_ _56296_/A _56298_/X _56303_/C _56303_/Y sky130_fd_sc_hd__nand3_4
X_87123_ _87137_/CLK _87123_/D _87123_/Q sky130_fd_sc_hd__dfxtp_4
X_53515_ _85622_/Q _53506_/X _53514_/Y _53515_/Y sky130_fd_sc_hd__o21ai_4
X_84335_ _83227_/CLK _63308_/Y _79231_/A sky130_fd_sc_hd__dfxtp_4
X_50727_ _50506_/A _50727_/X sky130_fd_sc_hd__buf_2
X_57283_ _57049_/A _57283_/B _57326_/C _57283_/Y sky130_fd_sc_hd__nor3_4
X_81547_ _81412_/CLK _81547_/D _76595_/B sky130_fd_sc_hd__dfxtp_4
X_69269_ _69216_/X _69267_/Y _69231_/X _69268_/Y _69269_/X sky130_fd_sc_hd__a211o_4
X_54495_ _54492_/Y _54475_/X _54494_/X _85432_/D sky130_fd_sc_hd__a21oi_4
X_59022_ _58925_/X _85439_/Q _59021_/X _59022_/Y sky130_fd_sc_hd__o21ai_4
X_71300_ _71303_/A _71303_/B _70472_/X _71300_/Y sky130_fd_sc_hd__nand3_4
X_56234_ _56085_/X _56225_/X _56233_/Y _56234_/Y sky130_fd_sc_hd__o21ai_4
X_87054_ _88062_/CLK _44562_/Y _87054_/Q sky130_fd_sc_hd__dfxtp_4
X_41460_ _41449_/X _82337_/Q _41459_/X _41460_/Y sky130_fd_sc_hd__o21ai_4
X_53446_ _53445_/Y _85633_/D sky130_fd_sc_hd__inv_2
X_72280_ _72196_/X _85332_/Q _72255_/X _72280_/X sky130_fd_sc_hd__o21a_4
X_84266_ _84652_/CLK _64201_/Y _64200_/C sky130_fd_sc_hd__dfxtp_4
X_50658_ _86159_/Q _50654_/X _50657_/Y _50658_/Y sky130_fd_sc_hd__o21ai_4
X_81478_ _88116_/CLK _81478_/D _76692_/B sky130_fd_sc_hd__dfxtp_4
X_86005_ _86005_/CLK _86005_/D _86005_/Q sky130_fd_sc_hd__dfxtp_4
X_40411_ _40354_/X _40411_/X sky130_fd_sc_hd__buf_2
X_71231_ _48684_/B _71231_/A2 _71230_/Y _71231_/Y sky130_fd_sc_hd__o21ai_4
X_83217_ _83218_/CLK _72611_/X _83217_/Q sky130_fd_sc_hd__dfxtp_4
X_56165_ _56169_/A _56150_/B _56165_/C _56165_/Y sky130_fd_sc_hd__nand3_4
X_80429_ _80446_/B _80429_/B _80429_/X sky130_fd_sc_hd__xor2_4
X_41391_ _81741_/Q _41325_/X _41391_/X sky130_fd_sc_hd__or2_4
X_53377_ _53374_/Y _53355_/X _53376_/X _85645_/D sky130_fd_sc_hd__a21oi_4
X_84197_ _84197_/CLK _84197_/D _84197_/Q sky130_fd_sc_hd__dfxtp_4
X_50589_ _50587_/Y _50551_/X _50588_/X _86172_/D sky130_fd_sc_hd__a21oi_4
X_43130_ _43189_/A _43130_/X sky130_fd_sc_hd__buf_2
X_55116_ _55112_/A _47877_/A _55120_/C _47814_/A _55116_/X sky130_fd_sc_hd__and4_4
X_52328_ _52320_/A _52328_/B _52328_/X sky130_fd_sc_hd__and2_4
X_40342_ _74492_/A _40342_/X sky130_fd_sc_hd__buf_2
X_71162_ _70758_/A _71162_/B _70827_/C _70578_/A _71163_/A sky130_fd_sc_hd__nand4_4
X_83148_ _86218_/CLK _73506_/X _83148_/Q sky130_fd_sc_hd__dfxtp_4
X_56096_ _56100_/A _56115_/B _85297_/Q _56096_/Y sky130_fd_sc_hd__nand3_4
X_70113_ _70113_/A _70117_/A sky130_fd_sc_hd__inv_2
X_43061_ _43121_/A _43061_/X sky130_fd_sc_hd__buf_2
X_55047_ _47838_/X _55054_/A sky130_fd_sc_hd__buf_2
X_59924_ _59923_/Y _62237_/A sky130_fd_sc_hd__buf_2
X_52259_ _52250_/A _48878_/B _52259_/Y sky130_fd_sc_hd__nand2_4
X_71093_ _70905_/D _70959_/B _71093_/C _71115_/D _71093_/X sky130_fd_sc_hd__and4_4
X_75970_ _75970_/A _75969_/Y _81737_/D sky130_fd_sc_hd__xor2_4
X_83079_ _83589_/CLK _74376_/Y _83079_/Q sky130_fd_sc_hd__dfxtp_4
X_87956_ _87126_/CLK _87956_/D _87956_/Q sky130_fd_sc_hd__dfxtp_4
X_42012_ _41998_/X _42010_/X _40820_/X _42011_/Y _42000_/X _42012_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74921_ _80757_/Q _74921_/B _74923_/A sky130_fd_sc_hd__or2_4
X_70044_ _69655_/A _70044_/X sky130_fd_sc_hd__buf_2
X_86907_ _84420_/CLK _44978_/Y _63049_/B sky130_fd_sc_hd__dfxtp_4
X_59855_ _59855_/A _59855_/B _80347_/A _59855_/Y sky130_fd_sc_hd__nor3_4
X_87887_ _88144_/CLK _87887_/D _87887_/Q sky130_fd_sc_hd__dfxtp_4
X_46820_ _82956_/Q _46820_/Y sky130_fd_sc_hd__inv_2
X_58806_ _58897_/A _58873_/B sky130_fd_sc_hd__buf_2
X_77640_ _77638_/Y _77639_/Y _77645_/B sky130_fd_sc_hd__and2_4
X_74852_ _74850_/Y _74852_/B _74853_/B sky130_fd_sc_hd__xnor2_4
X_86838_ _87225_/CLK _45965_/X _66577_/B sky130_fd_sc_hd__dfxtp_4
X_59786_ _59743_/B _59688_/X _59783_/Y _59763_/X _59785_/Y _59786_/Y
+ sky130_fd_sc_hd__a41oi_4
X_56998_ _45673_/A _56997_/X _56998_/Y sky130_fd_sc_hd__nor2_4
X_73803_ _44695_/Y _73728_/X _73802_/Y _73815_/C sky130_fd_sc_hd__a21o_4
X_46751_ _46751_/A _46751_/X sky130_fd_sc_hd__buf_2
X_58737_ _84804_/Q _58725_/X _58729_/X _58736_/X _84804_/D sky130_fd_sc_hd__a2bb2oi_4
X_77571_ _77567_/Y _77570_/C _77570_/A _77571_/Y sky130_fd_sc_hd__o21ai_4
X_43963_ _44053_/A _43944_/A _43945_/Y _43962_/X _43963_/X sky130_fd_sc_hd__a211o_4
X_55949_ _55949_/A _55949_/B _55949_/X sky130_fd_sc_hd__and2_4
X_74783_ _74783_/A _74796_/B _74796_/C _71016_/A _74783_/Y sky130_fd_sc_hd__nand4_4
X_86769_ _84970_/CLK _86769_/D _44131_/A sky130_fd_sc_hd__dfxtp_4
X_71995_ _71992_/Y _71969_/X _71994_/Y _71995_/Y sky130_fd_sc_hd__a21boi_4
X_79310_ _79310_/A _79310_/B _79311_/B sky130_fd_sc_hd__xor2_4
X_45702_ _85069_/Q _55186_/B sky130_fd_sc_hd__inv_2
X_76522_ _76522_/A _76522_/B _76522_/Y sky130_fd_sc_hd__nand2_4
X_42914_ _42895_/X _42896_/X _41705_/X _67675_/B _42905_/X _42914_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49470_ _49496_/A _49470_/X sky130_fd_sc_hd__buf_2
X_73734_ _73731_/X _86234_/Q _73683_/X _73733_/X _73734_/X sky130_fd_sc_hd__a211o_4
X_58668_ _58125_/X _85785_/Q _58126_/X _58668_/X sky130_fd_sc_hd__o21a_4
X_70946_ _50738_/B _70937_/X _70945_/Y _70946_/Y sky130_fd_sc_hd__o21ai_4
X_46682_ _46717_/A _46682_/B _46682_/C _50919_/D _46682_/X sky130_fd_sc_hd__and4_4
X_43894_ _41328_/X _43886_/X _67527_/B _43887_/X _43894_/X sky130_fd_sc_hd__a2bb2o_4
X_48421_ _48613_/A _48469_/A sky130_fd_sc_hd__buf_2
X_79241_ _79238_/Y _79240_/Y _79251_/B sky130_fd_sc_hd__nand2_4
X_45633_ _55483_/A _45354_/X _45633_/Y sky130_fd_sc_hd__nor2_4
X_57619_ _57619_/A _57619_/B _71960_/C _57619_/X sky130_fd_sc_hd__and3_4
X_76453_ _76453_/A _76453_/Y sky130_fd_sc_hd__inv_2
X_42845_ _42845_/A _87688_/D sky130_fd_sc_hd__inv_2
X_73665_ _72829_/A _73665_/X sky130_fd_sc_hd__buf_2
X_70877_ _50961_/B _70855_/A _70876_/Y _70877_/Y sky130_fd_sc_hd__o21ai_4
X_58599_ _58599_/A _58599_/X sky130_fd_sc_hd__buf_2
X_75404_ _75404_/A _75404_/B _75383_/X _75386_/B _75404_/X sky130_fd_sc_hd__and4_4
X_48352_ _48392_/A _50389_/B _48352_/Y sky130_fd_sc_hd__nand2_4
X_60630_ _60630_/A _60620_/C _60630_/C _60620_/B _60631_/D sky130_fd_sc_hd__and4_4
X_72616_ _60053_/X _72614_/X _72625_/B _72607_/Y _72615_/Y _72616_/Y
+ sky130_fd_sc_hd__a41oi_4
X_79172_ _84787_/Q _82723_/D _79174_/A sky130_fd_sc_hd__nor2_4
X_45564_ _45511_/X _61451_/A _45530_/X _45564_/Y sky130_fd_sc_hd__o21ai_4
X_76384_ _76369_/X _76370_/Y _76364_/X _76384_/Y sky130_fd_sc_hd__a21boi_4
X_42776_ _42774_/X _42775_/X _41321_/X _87724_/Q _42750_/X _42776_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73596_ _68415_/Y _73250_/X _73344_/X _73595_/Y _73596_/X sky130_fd_sc_hd__a211o_4
X_47303_ _47330_/A _47311_/B _47321_/C _52971_/D _47303_/X sky130_fd_sc_hd__and4_4
X_78123_ _82664_/Q _78123_/B _78123_/X sky130_fd_sc_hd__xor2_4
X_44515_ _44532_/A _44516_/A sky130_fd_sc_hd__buf_2
X_75335_ _75331_/Y _75333_/Y _75330_/Y _75339_/C sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_482_0_CLK clkbuf_9_241_0_CLK/X _86282_/CLK sky130_fd_sc_hd__clkbuf_1
X_41727_ _41727_/A _41727_/X sky130_fd_sc_hd__buf_2
X_48283_ _48280_/Y _48273_/X _48282_/Y _86543_/D sky130_fd_sc_hd__a21boi_4
X_60561_ _60465_/Y _60481_/A _60471_/X _60557_/Y _60560_/Y _60561_/Y
+ sky130_fd_sc_hd__a41oi_4
X_72547_ _72573_/A _72544_/B _79456_/B _72547_/Y sky130_fd_sc_hd__nor3_4
X_45495_ _45495_/A _45381_/B _45495_/Y sky130_fd_sc_hd__nand2_4
X_62300_ _62214_/A _62300_/X sky130_fd_sc_hd__buf_2
X_47234_ _47140_/A _47234_/X sky130_fd_sc_hd__buf_2
X_78054_ _60817_/C _78054_/B _78054_/X sky130_fd_sc_hd__xor2_4
X_44446_ _44587_/A _44547_/A sky130_fd_sc_hd__buf_2
X_63280_ _63272_/A _63280_/B _63280_/C _63280_/Y sky130_fd_sc_hd__nand3_4
X_75266_ _80783_/Q _81039_/D _80751_/D sky130_fd_sc_hd__xor2_4
X_41658_ _41658_/A _88174_/D sky130_fd_sc_hd__inv_2
X_60492_ _79151_/A _60246_/X _60488_/Y _60491_/X _60492_/Y sky130_fd_sc_hd__a2bb2oi_4
X_72478_ _64758_/X _85314_/Q _57763_/X _72478_/X sky130_fd_sc_hd__o21a_4
X_77005_ _77013_/A _77013_/B _77006_/B sky130_fd_sc_hd__xor2_4
X_62231_ _59918_/Y _62471_/A sky130_fd_sc_hd__buf_2
X_74217_ _74237_/A _86533_/Q _74217_/X sky130_fd_sc_hd__and2_4
X_40609_ _40601_/X _81148_/Q _40608_/X _40610_/A sky130_fd_sc_hd__o21a_4
X_47165_ _83695_/Q _47165_/Y sky130_fd_sc_hd__inv_2
X_71429_ _71429_/A _71432_/D sky130_fd_sc_hd__buf_2
X_44377_ _44363_/X _44377_/X sky130_fd_sc_hd__buf_2
X_75197_ _75217_/A _75196_/Y _81034_/D sky130_fd_sc_hd__xnor2_4
X_41589_ _41482_/A _41624_/B sky130_fd_sc_hd__buf_2
X_46116_ _46141_/A _80653_/Q _46204_/D sky130_fd_sc_hd__nor2_4
Xclkbuf_10_497_0_CLK clkbuf_9_248_0_CLK/X _83673_/CLK sky130_fd_sc_hd__clkbuf_1
X_43328_ _41272_/X _43325_/X _87478_/Q _43326_/X _43328_/X sky130_fd_sc_hd__a2bb2o_4
X_62162_ _58987_/A _62162_/X sky130_fd_sc_hd__buf_2
X_74148_ _74141_/Y _74142_/Y _74147_/X _74148_/Y sky130_fd_sc_hd__o21ai_4
X_47096_ _47004_/A _47096_/X sky130_fd_sc_hd__buf_2
X_61113_ _61066_/Y _61205_/A sky130_fd_sc_hd__buf_2
X_46047_ _45981_/X _46047_/X sky130_fd_sc_hd__buf_2
X_43259_ _43259_/A _87513_/D sky130_fd_sc_hd__inv_2
X_66970_ _80913_/D _66850_/X _66969_/X _84089_/D sky130_fd_sc_hd__a21bo_4
X_62093_ _59858_/A _61618_/X _62092_/X _62093_/X sky130_fd_sc_hd__a21o_4
X_78956_ _78956_/A _78956_/B _78957_/B sky130_fd_sc_hd__nand2_4
X_74079_ _74079_/A _74078_/X _74079_/Y sky130_fd_sc_hd__nand2_4
X_65921_ _44263_/X _65921_/B _65921_/X sky130_fd_sc_hd__and2_4
X_61044_ _60993_/B _60954_/X _60908_/A _61044_/X sky130_fd_sc_hd__o21a_4
X_77907_ _82246_/Q _81958_/Q _77907_/Y sky130_fd_sc_hd__xnor2_4
Xclkbuf_10_420_0_CLK clkbuf_9_210_0_CLK/X _83508_/CLK sky130_fd_sc_hd__clkbuf_1
X_78887_ _78880_/Y _78881_/A _78886_/Y _78888_/B sky130_fd_sc_hd__a21oi_4
X_49806_ _49861_/A _49830_/B sky130_fd_sc_hd__buf_2
X_68640_ _68640_/A _68640_/X sky130_fd_sc_hd__buf_2
X_65852_ _65811_/X _83053_/Q _65768_/X _65851_/X _65852_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_4_12_1_CLK clkbuf_4_12_1_CLK/A clkbuf_4_12_1_CLK/X sky130_fd_sc_hd__clkbuf_1
X_77838_ _77814_/Y _77838_/Y sky130_fd_sc_hd__inv_2
X_47998_ _47840_/A _47998_/X sky130_fd_sc_hd__buf_2
X_64803_ _64803_/A _64804_/A sky130_fd_sc_hd__buf_2
X_49737_ _86332_/Q _49715_/X _49736_/Y _49737_/Y sky130_fd_sc_hd__o21ai_4
X_68571_ _69797_/A _68571_/X sky130_fd_sc_hd__buf_2
X_46949_ _59030_/A _46908_/X _46948_/Y _46949_/Y sky130_fd_sc_hd__o21ai_4
X_65783_ _65812_/A _86506_/Q _65783_/X sky130_fd_sc_hd__and2_4
X_77769_ _82263_/Q _81975_/Q _81927_/D sky130_fd_sc_hd__xor2_4
X_62995_ _63285_/A _63285_/B _62995_/C _62995_/Y sky130_fd_sc_hd__nor3_4
X_67522_ _66898_/X _67522_/X sky130_fd_sc_hd__buf_2
X_79508_ _79505_/Y _79488_/Y _79507_/X _79510_/A sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_435_0_CLK clkbuf_9_217_0_CLK/X _84223_/CLK sky130_fd_sc_hd__clkbuf_1
X_64734_ _64684_/A _86461_/Q _64734_/X sky130_fd_sc_hd__and2_4
X_61946_ _61787_/X _61947_/D sky130_fd_sc_hd__buf_2
X_49668_ _49641_/A _49669_/B sky130_fd_sc_hd__buf_2
X_80780_ _80849_/CLK _80780_/D _80780_/Q sky130_fd_sc_hd__dfxtp_4
X_48619_ _48618_/Y _48565_/B _48619_/Y sky130_fd_sc_hd__nand2_4
X_67453_ _67381_/A _67453_/B _67453_/X sky130_fd_sc_hd__and2_4
X_79439_ _79439_/A _79429_/X _79439_/Y sky130_fd_sc_hd__nand2_4
X_64665_ _64665_/A _64666_/A sky130_fd_sc_hd__buf_2
X_49599_ _49595_/Y _49596_/X _49598_/X _86358_/D sky130_fd_sc_hd__a21oi_4
X_61877_ _61777_/A _61878_/C sky130_fd_sc_hd__buf_2
X_66404_ _64822_/X _66417_/B _64824_/X _66404_/Y sky130_fd_sc_hd__nand3_4
X_51630_ _51629_/X _51619_/B _51608_/X _53155_/D _51630_/X sky130_fd_sc_hd__and4_4
X_63616_ _63614_/Y _63578_/X _63615_/Y _63616_/Y sky130_fd_sc_hd__a21oi_4
X_82450_ _82822_/CLK _79142_/X _82450_/Q sky130_fd_sc_hd__dfxtp_4
X_60828_ _64738_/A _72592_/A sky130_fd_sc_hd__buf_2
X_67384_ _67379_/X _67382_/X _67383_/X _67387_/A sky130_fd_sc_hd__a21o_4
X_64596_ _64731_/A _64683_/A sky130_fd_sc_hd__buf_2
X_81401_ _81351_/CLK _83937_/Q _76707_/B sky130_fd_sc_hd__dfxtp_4
X_69123_ _87988_/Q _69121_/X _69051_/X _69122_/X _69123_/X sky130_fd_sc_hd__a211o_4
X_66335_ _65300_/X _86211_/Q _64692_/X _66334_/X _66335_/X sky130_fd_sc_hd__a211o_4
X_51561_ _51545_/A _53086_/B _51561_/Y sky130_fd_sc_hd__nand2_4
X_82381_ _82381_/CLK _82189_/Q _47111_/A sky130_fd_sc_hd__dfxtp_4
X_63547_ _58562_/A _63497_/X _61513_/A _63498_/X _63547_/X sky130_fd_sc_hd__a2bb2o_4
X_60759_ _63389_/D _60804_/B _59512_/X _60758_/X _60690_/X _60759_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_53300_ _51822_/A _53355_/A sky130_fd_sc_hd__buf_2
X_84120_ _81019_/CLK _84120_/D _84120_/Q sky130_fd_sc_hd__dfxtp_4
X_50512_ _50509_/Y _50491_/X _50511_/X _86187_/D sky130_fd_sc_hd__a21oi_4
X_81332_ _81755_/CLK _76424_/X _81708_/D sky130_fd_sc_hd__dfxtp_4
X_69054_ _74204_/A _69007_/X _69051_/X _69053_/Y _69054_/X sky130_fd_sc_hd__a211o_4
X_54280_ _54278_/Y _54051_/X _54279_/X _54280_/Y sky130_fd_sc_hd__a21oi_4
X_66266_ _65484_/A _66266_/X sky130_fd_sc_hd__buf_2
X_51492_ _86000_/Q _51485_/X _51491_/Y _51492_/Y sky130_fd_sc_hd__o21ai_4
X_63478_ _63478_/A _63491_/B sky130_fd_sc_hd__buf_2
X_68005_ _68002_/X _68004_/X _68005_/Y sky130_fd_sc_hd__nand2_4
X_53231_ _53228_/Y _53215_/X _53230_/X _53231_/Y sky130_fd_sc_hd__a21oi_4
X_65217_ _65178_/X _86730_/Q _65108_/X _65216_/X _65217_/X sky130_fd_sc_hd__a211o_4
X_84051_ _84049_/CLK _84051_/D _81483_/D sky130_fd_sc_hd__dfxtp_4
X_50443_ _50443_/A _50456_/B _50462_/C _50443_/X sky130_fd_sc_hd__and3_4
X_62429_ _62415_/X _57683_/X _62565_/C _62608_/D _62429_/X sky130_fd_sc_hd__and4_4
X_81263_ _81296_/CLK _81295_/Q _76332_/A sky130_fd_sc_hd__dfxtp_4
X_66197_ _64598_/X _86221_/Q _65761_/X _66196_/X _66197_/X sky130_fd_sc_hd__a211o_4
X_83002_ _82998_/CLK _83002_/D _83002_/Q sky130_fd_sc_hd__dfxtp_4
X_80214_ _84950_/Q _65481_/C _80216_/A sky130_fd_sc_hd__xor2_4
X_53162_ _85685_/Q _53146_/X _53161_/Y _53162_/Y sky130_fd_sc_hd__o21ai_4
X_65148_ _65118_/X _85516_/Q _65146_/X _65147_/X _65148_/X sky130_fd_sc_hd__a211o_4
X_50374_ _50383_/A _48335_/B _50374_/Y sky130_fd_sc_hd__nand2_4
X_81194_ _84115_/CLK _81194_/D _49119_/A sky130_fd_sc_hd__dfxtp_4
X_52113_ _53636_/A _52135_/B _52097_/X _52113_/X sky130_fd_sc_hd__and3_4
X_87810_ _87553_/CLK _42588_/Y _69790_/A sky130_fd_sc_hd__dfxtp_4
X_80145_ _80143_/X _80144_/X _80145_/Y sky130_fd_sc_hd__xnor2_4
X_53093_ _53172_/A _53093_/X sky130_fd_sc_hd__buf_2
X_57970_ _84936_/Q _57896_/X _57961_/X _57969_/X _57970_/Y sky130_fd_sc_hd__a2bb2oi_4
X_65079_ _65381_/A _86415_/Q _65079_/X sky130_fd_sc_hd__and2_4
X_69956_ _69956_/A _73509_/A _69956_/X sky130_fd_sc_hd__and2_4
X_52044_ _66209_/B _52041_/X _52043_/Y _52044_/Y sky130_fd_sc_hd__o21ai_4
X_56921_ _56917_/Y _56921_/B _56921_/C _85123_/D sky130_fd_sc_hd__nand3_4
X_68907_ _69146_/A _68907_/X sky130_fd_sc_hd__buf_2
X_87741_ _88001_/CLK _42747_/X _68918_/B sky130_fd_sc_hd__dfxtp_4
X_84953_ _85404_/CLK _84953_/D _84953_/Q sky130_fd_sc_hd__dfxtp_4
X_80076_ _80063_/X _80074_/X _80075_/X _80076_/Y sky130_fd_sc_hd__a21oi_4
X_69887_ _69884_/X _69886_/X _69624_/X _69887_/X sky130_fd_sc_hd__a21o_4
X_83904_ _81928_/CLK _83904_/D _81976_/D sky130_fd_sc_hd__dfxtp_4
X_59640_ _59640_/A _60402_/A sky130_fd_sc_hd__buf_2
X_56852_ _56852_/A _56730_/X _56851_/X _56852_/X sky130_fd_sc_hd__or3_4
X_68838_ _68586_/A _68838_/X sky130_fd_sc_hd__buf_2
X_87672_ _87675_/CLK _87672_/D _67223_/B sky130_fd_sc_hd__dfxtp_4
X_84884_ _84884_/CLK _84884_/D _64536_/C sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_509_0_CLK clkbuf_9_509_0_CLK/A clkbuf_9_509_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_55803_ _44077_/X _56341_/C _55803_/X sky130_fd_sc_hd__and2_4
X_86623_ _84922_/CLK _47550_/Y _86623_/Q sky130_fd_sc_hd__dfxtp_4
X_59571_ _59562_/B _59571_/B _59571_/C _59741_/C _60160_/B sky130_fd_sc_hd__nand4_4
X_83835_ _83835_/CLK _83835_/D _83835_/Q sky130_fd_sc_hd__dfxtp_4
X_56783_ _83324_/Q _56783_/X sky130_fd_sc_hd__buf_2
X_68769_ _88003_/Q _68715_/X _68540_/X _68768_/X _68769_/X sky130_fd_sc_hd__a211o_4
X_53995_ _53991_/A _46376_/Y _53995_/Y sky130_fd_sc_hd__nand2_4
X_70800_ _71221_/A _70712_/A _70800_/X sky130_fd_sc_hd__and2_4
X_58522_ _58522_/A _58522_/Y sky130_fd_sc_hd__inv_2
X_55734_ _55731_/X _55733_/X _44108_/X _55734_/Y sky130_fd_sc_hd__a21oi_4
X_86554_ _86554_/CLK _48218_/Y _86554_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_62_0_CLK clkbuf_8_63_0_CLK/A clkbuf_8_62_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_40960_ _40944_/X _40946_/X _40959_/X _88303_/Q _40916_/X _40960_/Y
+ sky130_fd_sc_hd__o32ai_4
X_52946_ _52892_/A _52946_/X sky130_fd_sc_hd__buf_2
X_71780_ _71761_/Y _83378_/Q _71779_/X _83378_/D sky130_fd_sc_hd__a21o_4
X_83766_ _83766_/CLK _83766_/D _58356_/B sky130_fd_sc_hd__dfxtp_4
X_80978_ _81059_/CLK _75724_/X _75124_/B sky130_fd_sc_hd__dfxtp_4
X_85505_ _85505_/CLK _85505_/D _85505_/Q sky130_fd_sc_hd__dfxtp_4
X_70731_ _70358_/X _70827_/B _71735_/D sky130_fd_sc_hd__nor2_4
X_58453_ _58448_/X _83477_/Q _58452_/Y _84845_/D sky130_fd_sc_hd__o21a_4
X_82717_ _82503_/CLK _82717_/D _82673_/D sky130_fd_sc_hd__dfxtp_4
X_55665_ _55243_/A _83317_/Q _55243_/B _55665_/Y sky130_fd_sc_hd__nand3_4
X_86485_ _86196_/CLK _86485_/D _65612_/B sky130_fd_sc_hd__dfxtp_4
X_40891_ _40890_/X _40821_/X _88316_/Q _40822_/X _40891_/X sky130_fd_sc_hd__a2bb2o_4
X_52877_ _85738_/Q _52874_/X _52876_/Y _52877_/Y sky130_fd_sc_hd__o21ai_4
X_83697_ _83699_/CLK _70808_/Y _83697_/Q sky130_fd_sc_hd__dfxtp_4
X_57404_ _57394_/X _56634_/X _45584_/A _57395_/X _85013_/D sky130_fd_sc_hd__a2bb2o_4
X_88224_ _88224_/CLK _88224_/D _67801_/B sky130_fd_sc_hd__dfxtp_4
X_42630_ _52754_/A _53189_/A sky130_fd_sc_hd__buf_2
X_54616_ _54344_/A _54616_/X sky130_fd_sc_hd__buf_2
X_73450_ _72909_/A _73450_/X sky130_fd_sc_hd__buf_2
X_85436_ _85436_/CLK _85436_/D _85436_/Q sky130_fd_sc_hd__dfxtp_4
X_51828_ _51805_/A _51815_/B _51810_/C _52654_/D _51828_/X sky130_fd_sc_hd__and4_4
X_70662_ _70500_/B _70662_/X sky130_fd_sc_hd__buf_2
X_82648_ _82648_/CLK _82648_/D _82648_/Q sky130_fd_sc_hd__dfxtp_4
X_58384_ _58366_/X _83351_/Q _58383_/Y _84863_/D sky130_fd_sc_hd__o21a_4
X_55596_ _44064_/X _55596_/B _55596_/Y sky130_fd_sc_hd__nor2_4
X_72401_ _86602_/Q _72401_/B _72401_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_8_77_0_CLK clkbuf_8_77_0_CLK/A clkbuf_8_77_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_57335_ _57331_/Y _57335_/B _57335_/Y sky130_fd_sc_hd__nand2_4
X_88155_ _88220_/CLK _41759_/Y _88155_/Q sky130_fd_sc_hd__dfxtp_4
X_42561_ _42554_/X _40802_/A _42477_/X _69661_/B _42556_/X _87820_/D
+ sky130_fd_sc_hd__o32ai_4
X_54547_ _85422_/Q _54540_/X _54546_/Y _54547_/Y sky130_fd_sc_hd__o21ai_4
X_73381_ _73381_/A _86473_/Q _73381_/X sky130_fd_sc_hd__and2_4
X_85367_ _83275_/CLK _54849_/Y _85367_/Q sky130_fd_sc_hd__dfxtp_4
X_51759_ _85951_/Q _51387_/X _51758_/Y _51759_/Y sky130_fd_sc_hd__o21ai_4
X_70593_ _74716_/A _70620_/D sky130_fd_sc_hd__buf_2
Xclkbuf_7_9_0_CLK clkbuf_6_4_0_CLK/X clkbuf_7_9_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_82579_ _82711_/CLK _82611_/Q _78198_/A sky130_fd_sc_hd__dfxtp_4
X_44300_ _64619_/A _58020_/A _59238_/A _44265_/D _44300_/Y sky130_fd_sc_hd__nor4_4
X_75120_ _75120_/A _75120_/B _75116_/X _75121_/B sky130_fd_sc_hd__nand3_4
X_87106_ _87926_/CLK _87106_/D _87106_/Q sky130_fd_sc_hd__dfxtp_4
X_41512_ _41511_/X _41486_/X _88201_/Q _41487_/X _41512_/X sky130_fd_sc_hd__a2bb2o_4
X_72332_ _72332_/A _72332_/B _72332_/Y sky130_fd_sc_hd__nor2_4
X_84318_ _84321_/CLK _84318_/D _80506_/B sky130_fd_sc_hd__dfxtp_4
X_45280_ _45268_/X _45276_/Y _45279_/Y _45280_/Y sky130_fd_sc_hd__a21oi_4
X_57266_ _45631_/Y _57247_/Y _57265_/X _85042_/D sky130_fd_sc_hd__o21ai_4
X_88086_ _88086_/CLK _41974_/Y _41973_/A sky130_fd_sc_hd__dfxtp_4
X_54478_ _54478_/A _54478_/B _54478_/Y sky130_fd_sc_hd__nand2_4
X_42492_ _42492_/A _87847_/D sky130_fd_sc_hd__inv_2
X_85298_ _85279_/CLK _56087_/Y _55851_/B sky130_fd_sc_hd__dfxtp_4
X_59005_ _84777_/Q _58956_/X _58998_/X _59004_/X _84777_/D sky130_fd_sc_hd__a2bb2oi_4
X_56217_ _56055_/X _56210_/X _56216_/Y _85272_/D sky130_fd_sc_hd__o21ai_4
X_44231_ _44231_/A _44242_/C sky130_fd_sc_hd__buf_2
X_75051_ _75051_/A _75051_/B _75050_/Y _75051_/X sky130_fd_sc_hd__and3_4
X_87037_ _87032_/CLK _87037_/D _87037_/Q sky130_fd_sc_hd__dfxtp_4
X_53429_ _53420_/A _53428_/X _53410_/C _51225_/D _53429_/X sky130_fd_sc_hd__and4_4
X_41443_ _41399_/X _41400_/X _41442_/X _88214_/Q _41388_/X _41444_/A
+ sky130_fd_sc_hd__o32ai_4
X_72263_ _83269_/Q _72263_/Y sky130_fd_sc_hd__inv_2
X_84249_ _84849_/CLK _64408_/X _79713_/B sky130_fd_sc_hd__dfxtp_4
X_57197_ _56848_/X _57196_/Y _57198_/B sky130_fd_sc_hd__nor2_4
X_74002_ _73992_/Y _74002_/B _74002_/X sky130_fd_sc_hd__xor2_4
X_71214_ _52216_/B _71190_/A _71213_/Y _71214_/Y sky130_fd_sc_hd__o21ai_4
X_44162_ _43957_/B _44160_/A _59901_/C _44025_/X _44162_/Y sky130_fd_sc_hd__a22oi_4
X_56148_ _56148_/A _56148_/X sky130_fd_sc_hd__buf_2
X_41374_ _41374_/A _41275_/B _41374_/X sky130_fd_sc_hd__or2_4
X_72194_ _59133_/A _72194_/X sky130_fd_sc_hd__buf_2
X_43113_ _87571_/Q _43113_/Y sky130_fd_sc_hd__inv_2
X_78810_ _78807_/Y _78809_/Y _78802_/Y _78810_/Y sky130_fd_sc_hd__a21oi_4
X_40325_ _40324_/X _40325_/X sky130_fd_sc_hd__buf_2
X_71145_ _71145_/A _71225_/A sky130_fd_sc_hd__buf_2
X_48970_ _48908_/A _71998_/B _48970_/X sky130_fd_sc_hd__and2_4
X_56079_ _56079_/A _56079_/X sky130_fd_sc_hd__buf_2
X_44093_ _55158_/A _55140_/A sky130_fd_sc_hd__buf_2
X_79790_ _79776_/Y _79790_/B _79790_/X sky130_fd_sc_hd__and2_4
X_47921_ _47913_/Y _47903_/X _47920_/X _47921_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_8_15_0_CLK clkbuf_7_7_0_CLK/X clkbuf_9_31_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_59907_ _59906_/X _63632_/A sky130_fd_sc_hd__buf_2
X_43044_ _42060_/X _43031_/X _40626_/X _43043_/Y _43034_/X _87596_/D
+ sky130_fd_sc_hd__o32ai_4
X_78741_ _78722_/A _78697_/X _78717_/X _78718_/Y _78742_/A sky130_fd_sc_hd__nand4_4
X_71076_ _71078_/A _71076_/B _71078_/C _71076_/Y sky130_fd_sc_hd__nand3_4
X_87939_ _88386_/CLK _87939_/D _87939_/Q sky130_fd_sc_hd__dfxtp_4
X_75953_ _75948_/Y _75949_/A _75952_/Y _75953_/Y sky130_fd_sc_hd__a21boi_4
X_74904_ _74904_/A _74904_/B _74904_/Y sky130_fd_sc_hd__nand2_4
X_70027_ _69520_/X _69727_/Y _70012_/X _70026_/Y _70027_/X sky130_fd_sc_hd__a211o_4
X_47852_ _47845_/Y _47846_/X _47851_/X _86592_/D sky130_fd_sc_hd__a21oi_4
X_59838_ _59758_/X _59654_/X _59724_/Y _59836_/Y _59837_/Y _59839_/A
+ sky130_fd_sc_hd__a41o_4
X_78672_ _78671_/X _78672_/Y sky130_fd_sc_hd__inv_2
X_75884_ _75762_/Y _80791_/D sky130_fd_sc_hd__inv_2
X_46803_ _46797_/Y _46798_/X _46802_/X _86702_/D sky130_fd_sc_hd__a21oi_4
X_77623_ _77605_/X _77623_/Y sky130_fd_sc_hd__inv_2
X_74835_ _74835_/A _74835_/Y sky130_fd_sc_hd__inv_2
X_47783_ _81222_/Q _47784_/A sky130_fd_sc_hd__inv_2
X_59769_ _44173_/X _59772_/A sky130_fd_sc_hd__buf_2
X_44995_ _45219_/A _44995_/X sky130_fd_sc_hd__buf_2
X_61800_ _61789_/X _61792_/X _61799_/Y _58162_/A _61719_/X _61800_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49522_ _49537_/A _49516_/B _49522_/C _52735_/D _49522_/X sky130_fd_sc_hd__and4_4
X_46734_ _58722_/A _46719_/X _46733_/Y _46734_/Y sky130_fd_sc_hd__o21ai_4
X_77554_ _77553_/B _77552_/Y _77553_/A _77558_/C sky130_fd_sc_hd__o21ai_4
X_43946_ _80667_/Q _43979_/A sky130_fd_sc_hd__buf_2
X_62780_ _62766_/A _62766_/B _84383_/Q _62780_/Y sky130_fd_sc_hd__nor3_4
X_74766_ _74735_/X _83844_/Q _74763_/X _74764_/X _74765_/X _74766_/X
+ sky130_fd_sc_hd__a2111o_4
X_71978_ _71978_/A _71978_/X sky130_fd_sc_hd__buf_2
Xclkbuf_3_1_1_CLK clkbuf_3_1_0_CLK/X clkbuf_4_3_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_76505_ _76501_/Y _76502_/Y _76504_/Y _76510_/A sky130_fd_sc_hd__or3_4
X_49453_ _49450_/Y _49434_/X _49452_/X _86385_/D sky130_fd_sc_hd__a21oi_4
X_61731_ _59684_/X _61791_/B sky130_fd_sc_hd__buf_2
X_73717_ _73717_/A _73717_/B _73717_/X sky130_fd_sc_hd__xor2_4
X_46665_ _46616_/A _46902_/A sky130_fd_sc_hd__buf_2
X_70929_ _46899_/X _70909_/A _70928_/Y _70929_/Y sky130_fd_sc_hd__o21ai_4
X_77485_ _77485_/A _82195_/D _81907_/D sky130_fd_sc_hd__xor2_4
X_43877_ _43862_/X _43876_/X _41277_/X _69100_/B _43863_/X _43877_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74697_ _74691_/A _45832_/A _74697_/Y sky130_fd_sc_hd__nand2_4
X_48404_ _49215_/A _48557_/A sky130_fd_sc_hd__buf_2
X_79224_ _79224_/A _79224_/B _79251_/A sky130_fd_sc_hd__nand2_4
X_45616_ _45395_/X _45616_/X sky130_fd_sc_hd__buf_2
X_64450_ _58264_/Y _64423_/X _64449_/Y _64450_/Y sky130_fd_sc_hd__o21ai_4
X_76436_ _81365_/Q _76435_/Y _81333_/D sky130_fd_sc_hd__xor2_4
X_42828_ _42816_/X _42817_/X _41473_/X _66651_/B _42805_/X _42828_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49384_ _49520_/A _49493_/A sky130_fd_sc_hd__buf_2
X_61662_ _61658_/X _61645_/X _61661_/Y _84462_/D sky130_fd_sc_hd__a21oi_4
X_73648_ _70122_/Y _86754_/D _73647_/X _73648_/Y sky130_fd_sc_hd__o21ai_4
X_46596_ _46491_/A _51394_/B _46596_/Y sky130_fd_sc_hd__nand2_4
X_63401_ _61364_/B _60834_/X _63399_/X _63400_/X _63401_/X sky130_fd_sc_hd__a211o_4
X_48335_ _48401_/A _48335_/B _48335_/Y sky130_fd_sc_hd__nand2_4
X_60613_ _60359_/X _60524_/Y _60392_/B _60598_/Y _60612_/Y _60613_/Y
+ sky130_fd_sc_hd__a41oi_4
X_79155_ _79155_/A _84487_/Q _79155_/X sky130_fd_sc_hd__xor2_4
X_45547_ _85079_/Q _55520_/B sky130_fd_sc_hd__inv_2
X_64381_ _64323_/A _64381_/X sky130_fd_sc_hd__buf_2
X_76367_ _76366_/A _76366_/B _76368_/A sky130_fd_sc_hd__nand2_4
X_42759_ _42822_/A _42759_/X sky130_fd_sc_hd__buf_2
X_61593_ _61541_/A _61593_/B _61619_/C _61593_/Y sky130_fd_sc_hd__nand3_4
X_73579_ _73576_/X _73578_/X _73489_/X _73582_/A sky130_fd_sc_hd__a21o_4
X_66120_ _66117_/X _84979_/Q _66118_/X _66119_/X _66120_/X sky130_fd_sc_hd__a211o_4
X_78106_ _78130_/A _78105_/Y _78107_/B sky130_fd_sc_hd__xor2_4
X_63332_ _63289_/X _64536_/C _63341_/C _63332_/D _63332_/X sky130_fd_sc_hd__and4_4
X_75318_ _75314_/Y _75319_/B _75317_/Y _75318_/X sky130_fd_sc_hd__o21a_4
X_48266_ _86545_/Q _48263_/X _48265_/Y _48266_/Y sky130_fd_sc_hd__o21ai_4
X_60544_ _60541_/Y _60475_/A _60543_/Y _79143_/A _60341_/X _60544_/X
+ sky130_fd_sc_hd__o32a_4
X_79086_ _79086_/A _79086_/B _79095_/A sky130_fd_sc_hd__xnor2_4
X_45478_ _45473_/X _45477_/X _45446_/X _45478_/X sky130_fd_sc_hd__a21o_4
X_76298_ _76289_/A _81560_/Q _76298_/Y sky130_fd_sc_hd__nand2_4
X_47217_ _54612_/D _47218_/D sky130_fd_sc_hd__buf_2
X_66051_ _65990_/X _86231_/Q _66021_/X _66050_/X _66051_/X sky130_fd_sc_hd__a211o_4
X_78037_ _78037_/A _78037_/B _82145_/D sky130_fd_sc_hd__nand2_4
X_44429_ _44425_/X _44427_/X _41574_/X _87113_/Q _44428_/X _44430_/A
+ sky130_fd_sc_hd__o32ai_4
X_75249_ _75241_/Y _75248_/Y _75249_/Y sky130_fd_sc_hd__xnor2_4
X_63263_ _63203_/X _64467_/C _63204_/X _63332_/D _63263_/X sky130_fd_sc_hd__and4_4
X_48197_ _48191_/Y _48194_/X _48196_/X _48197_/Y sky130_fd_sc_hd__a21oi_4
X_60475_ _60475_/A _60586_/A sky130_fd_sc_hd__inv_2
X_65002_ _65002_/A _65002_/B _65002_/X sky130_fd_sc_hd__and2_4
X_62214_ _62214_/A _62214_/X sky130_fd_sc_hd__buf_2
X_47148_ _83697_/Q _53395_/B sky130_fd_sc_hd__inv_2
X_63194_ _63144_/X _84841_/Q _63146_/C _63239_/D _63194_/X sky130_fd_sc_hd__and4_4
X_69810_ _69806_/X _69809_/X _69768_/X _69810_/X sky130_fd_sc_hd__a21o_4
X_62145_ _62143_/Y _62101_/X _62144_/Y _62145_/Y sky130_fd_sc_hd__a21oi_4
X_47079_ _47063_/A _52843_/B _47079_/Y sky130_fd_sc_hd__nand2_4
X_79988_ _79988_/A _79988_/B _79989_/A sky130_fd_sc_hd__and2_4
X_69741_ _73104_/A _69690_/X _68473_/X _69740_/X _69741_/X sky130_fd_sc_hd__a211o_4
X_50090_ _50103_/A _48955_/X _50090_/Y sky130_fd_sc_hd__nand2_4
X_66953_ _68342_/A _66953_/X sky130_fd_sc_hd__buf_2
X_62076_ _63629_/B _61999_/B _62046_/C _62046_/D _62077_/D sky130_fd_sc_hd__nand4_4
X_78939_ _78939_/A _78939_/B _82704_/D sky130_fd_sc_hd__xor2_4
X_65904_ _65790_/A _65904_/X sky130_fd_sc_hd__buf_2
X_61027_ _60915_/A _60892_/Y _60853_/X _61027_/X sky130_fd_sc_hd__and3_4
X_69672_ _69733_/A _69672_/X sky130_fd_sc_hd__buf_2
X_81950_ _82047_/CLK _78013_/Y _77671_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_480_0_CLK clkbuf_8_240_0_CLK/X clkbuf_9_480_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_66884_ _66956_/A _88198_/Q _66884_/X sky130_fd_sc_hd__and2_4
X_80901_ _82067_/CLK _80901_/D _75598_/A sky130_fd_sc_hd__dfxtp_4
X_68623_ _68620_/X _68622_/X _68477_/X _68623_/Y sky130_fd_sc_hd__a21oi_4
X_65835_ _64691_/X _86182_/Q _64972_/X _65834_/X _65835_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_374_0_CLK clkbuf_9_187_0_CLK/X _85433_/CLK sky130_fd_sc_hd__clkbuf_1
X_81881_ _82531_/CLK _78072_/X _81881_/Q sky130_fd_sc_hd__dfxtp_4
X_52800_ _85752_/Q _52792_/X _52799_/Y _52800_/Y sky130_fd_sc_hd__o21ai_4
X_83620_ _85561_/CLK _83620_/D _48930_/A sky130_fd_sc_hd__dfxtp_4
X_80832_ _81065_/CLK _83976_/Q _75695_/B sky130_fd_sc_hd__dfxtp_4
X_68554_ _43043_/A _68527_/X _68552_/X _68553_/X _68554_/X sky130_fd_sc_hd__a211o_4
X_53780_ _53766_/A _48876_/Y _53780_/Y sky130_fd_sc_hd__nand2_4
X_65766_ _65733_/X _85579_/Q _65734_/X _65765_/X _65766_/X sky130_fd_sc_hd__a211o_4
X_50992_ _51101_/A _50992_/X sky130_fd_sc_hd__buf_2
X_62978_ _62976_/X _62942_/X _62977_/Y _62978_/Y sky130_fd_sc_hd__a21oi_4
X_67505_ _87160_/Q _67432_/X _67433_/X _67504_/X _67506_/B sky130_fd_sc_hd__a211o_4
X_52731_ _52727_/Y _52728_/X _52730_/X _52731_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_495_0_CLK clkbuf_9_495_0_CLK/A clkbuf_9_495_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_64717_ _64717_/A _64903_/A sky130_fd_sc_hd__buf_2
X_83551_ _83550_/CLK _83551_/D _47694_/A sky130_fd_sc_hd__dfxtp_4
X_61929_ _61915_/A _61915_/B _63520_/B _61915_/D _61929_/X sky130_fd_sc_hd__and4_4
X_80763_ _80854_/CLK _80763_/D _80763_/Q sky130_fd_sc_hd__dfxtp_4
X_68485_ _68409_/A _68485_/B _68485_/X sky130_fd_sc_hd__and2_4
X_65697_ _65929_/A _65775_/B sky130_fd_sc_hd__buf_2
X_82502_ _82675_/CLK _78839_/X _78370_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_389_0_CLK clkbuf_9_194_0_CLK/X _83227_/CLK sky130_fd_sc_hd__clkbuf_1
X_55450_ _55330_/X _55448_/Y _55449_/Y _55451_/B sky130_fd_sc_hd__o21a_4
X_67436_ _67436_/A _67435_/X _67436_/Y sky130_fd_sc_hd__nand2_4
X_86270_ _85561_/CLK _86270_/D _86270_/Q sky130_fd_sc_hd__dfxtp_4
X_52662_ _52659_/Y _52647_/X _52661_/X _52662_/Y sky130_fd_sc_hd__a21oi_4
X_64648_ _64577_/X _86751_/Q _64579_/X _64647_/X _64648_/X sky130_fd_sc_hd__a211o_4
X_83482_ _83482_/CLK _83482_/D _83482_/Q sky130_fd_sc_hd__dfxtp_4
X_80694_ _81104_/CLK _80694_/D _80694_/Q sky130_fd_sc_hd__dfxtp_4
X_54401_ _54401_/A _54402_/C sky130_fd_sc_hd__buf_2
X_85221_ _85221_/CLK _85221_/D _55730_/B sky130_fd_sc_hd__dfxtp_4
X_51613_ _51639_/A _51613_/X sky130_fd_sc_hd__buf_2
X_82433_ _82248_/CLK _82465_/Q _82433_/Q sky130_fd_sc_hd__dfxtp_4
X_55381_ _55316_/X _55328_/C _55382_/A sky130_fd_sc_hd__and2_4
X_67367_ _67367_/A _67366_/X _67367_/Y sky130_fd_sc_hd__nand2_4
XPHY_706 sky130_fd_sc_hd__decap_3
X_52593_ _52593_/A _52614_/A sky130_fd_sc_hd__buf_2
X_64579_ _64772_/A _64579_/X sky130_fd_sc_hd__buf_2
XPHY_717 sky130_fd_sc_hd__decap_3
X_57120_ _57109_/X _56639_/X _45595_/A _57110_/X _85076_/D sky130_fd_sc_hd__a2bb2o_4
X_69106_ _69102_/X _69105_/X _69017_/X _69106_/Y sky130_fd_sc_hd__a21oi_4
X_54332_ _54332_/A _54332_/B _54332_/Y sky130_fd_sc_hd__nand2_4
X_66318_ _65307_/A _66318_/X sky130_fd_sc_hd__buf_2
X_85152_ _85152_/CLK _56573_/X _85152_/Q sky130_fd_sc_hd__dfxtp_4
X_51544_ _51542_/Y _51531_/X _51543_/X _85991_/D sky130_fd_sc_hd__a21oi_4
X_82364_ _82925_/CLK _77007_/X _47893_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_312_0_CLK clkbuf_9_156_0_CLK/X _83380_/CLK sky130_fd_sc_hd__clkbuf_1
X_67298_ _67295_/X _67297_/X _67204_/X _67298_/X sky130_fd_sc_hd__a21o_4
X_84103_ _81169_/CLK _84103_/D _80927_/D sky130_fd_sc_hd__dfxtp_4
X_81315_ _84079_/CLK _76170_/X _81723_/D sky130_fd_sc_hd__dfxtp_4
X_57051_ _57051_/A _57051_/Y sky130_fd_sc_hd__inv_2
X_69037_ _69059_/A _88248_/Q _69037_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_942_0_CLK clkbuf_9_471_0_CLK/X _88060_/CLK sky130_fd_sc_hd__clkbuf_1
X_54263_ _54316_/A _54286_/A sky130_fd_sc_hd__buf_2
X_66249_ _66181_/A _74127_/B _66249_/X sky130_fd_sc_hd__and2_4
X_85083_ _85083_/CLK _85083_/D _85083_/Q sky130_fd_sc_hd__dfxtp_4
X_51475_ _51481_/A _52999_/B _51475_/Y sky130_fd_sc_hd__nand2_4
X_82295_ _82103_/CLK _77157_/B _82295_/Q sky130_fd_sc_hd__dfxtp_4
X_56002_ _56002_/A _56002_/Y sky130_fd_sc_hd__inv_2
X_53214_ _85675_/Q _53198_/X _53213_/Y _53214_/Y sky130_fd_sc_hd__o21ai_4
X_84034_ _81160_/CLK _68119_/X _82074_/D sky130_fd_sc_hd__dfxtp_4
X_50426_ _50424_/Y _50395_/X _50425_/X _86203_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_433_0_CLK clkbuf_8_216_0_CLK/X clkbuf_9_433_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_81246_ _85378_/CLK _81054_/Q _81246_/Q sky130_fd_sc_hd__dfxtp_4
X_54194_ _54194_/A _54215_/A sky130_fd_sc_hd__buf_2
Xclkbuf_opt_25_CLK _86505_/CLK _86473_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_10_327_0_CLK clkbuf_9_163_0_CLK/X _86342_/CLK sky130_fd_sc_hd__clkbuf_1
X_53145_ _53142_/Y _53137_/X _53144_/X _53145_/Y sky130_fd_sc_hd__a21oi_4
X_50357_ _50355_/Y _50351_/X _50356_/Y _50357_/Y sky130_fd_sc_hd__a21boi_4
X_81177_ _86758_/CLK _75014_/B _81177_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_957_0_CLK clkbuf_9_478_0_CLK/X _85895_/CLK sky130_fd_sc_hd__clkbuf_1
X_80128_ _80114_/Y _80119_/Y _80127_/X _80129_/B sky130_fd_sc_hd__o21ai_4
X_41090_ _41090_/A _41090_/Y sky130_fd_sc_hd__inv_2
X_57953_ _64621_/A _58721_/A sky130_fd_sc_hd__buf_2
X_53076_ _53080_/A _53076_/B _53076_/Y sky130_fd_sc_hd__nand2_4
X_69939_ _70001_/A _69939_/X sky130_fd_sc_hd__buf_2
X_50288_ _50286_/Y _50274_/X _50287_/Y _86231_/D sky130_fd_sc_hd__a21boi_4
X_85985_ _85697_/CLK _51576_/Y _85985_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_448_0_CLK clkbuf_8_224_0_CLK/X clkbuf_9_448_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_52027_ _52027_/A _48024_/B _52027_/Y sky130_fd_sc_hd__nand2_4
X_56904_ _56647_/X _56898_/Y _56725_/B _56903_/X _85124_/D sky130_fd_sc_hd__a2bb2o_4
X_87724_ _87708_/CLK _87724_/D _87724_/Q sky130_fd_sc_hd__dfxtp_4
X_72950_ _72949_/X _72951_/A sky130_fd_sc_hd__buf_2
X_84936_ _86317_/CLK _57970_/Y _84936_/Q sky130_fd_sc_hd__dfxtp_4
X_80059_ _84935_/Q _65713_/C _80059_/X sky130_fd_sc_hd__xor2_4
X_57884_ _45926_/X _57884_/X sky130_fd_sc_hd__buf_2
X_71901_ _56857_/X _71892_/X _71900_/Y _71901_/Y sky130_fd_sc_hd__o21ai_4
X_59623_ _60615_/A _59753_/B sky130_fd_sc_hd__buf_2
X_56835_ _56660_/A _56866_/A sky130_fd_sc_hd__buf_2
X_87655_ _86932_/CLK _42912_/X _87655_/Q sky130_fd_sc_hd__dfxtp_4
X_72881_ _72881_/A _86525_/Q _72881_/X sky130_fd_sc_hd__and2_4
X_84867_ _84250_/CLK _84867_/D _84867_/Q sky130_fd_sc_hd__dfxtp_4
X_43800_ _41059_/X _43770_/X _69443_/B _43772_/X _43800_/X sky130_fd_sc_hd__a2bb2o_4
X_74620_ _45331_/Y _74612_/X _74619_/X _83013_/D sky130_fd_sc_hd__o21ai_4
X_86606_ _86610_/CLK _86606_/D _86606_/Q sky130_fd_sc_hd__dfxtp_4
X_71832_ _71825_/X _83360_/Q _71831_/X _83360_/D sky130_fd_sc_hd__a21o_4
X_59554_ _59520_/A _59535_/A _59602_/A sky130_fd_sc_hd__and2_4
X_83818_ _83842_/CLK _70266_/X _74720_/B sky130_fd_sc_hd__dfxtp_4
X_44780_ _44766_/X _44767_/X _41376_/A _86958_/Q _44768_/X _44780_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56766_ _57023_/A _56766_/X sky130_fd_sc_hd__buf_2
X_87586_ _88111_/CLK _87586_/D _87586_/Q sky130_fd_sc_hd__dfxtp_4
X_41992_ _41992_/A _41993_/A sky130_fd_sc_hd__buf_2
X_53978_ _53978_/A _53978_/B _53978_/Y sky130_fd_sc_hd__nand2_4
X_84798_ _84797_/CLK _84798_/D _84798_/Q sky130_fd_sc_hd__dfxtp_4
X_58505_ _84832_/Q _58506_/A sky130_fd_sc_hd__buf_2
X_43731_ _40890_/X _43695_/X _87292_/Q _43696_/X _43731_/X sky130_fd_sc_hd__a2bb2o_4
X_55717_ _55714_/X _55716_/X _44108_/X _55717_/Y sky130_fd_sc_hd__a21oi_4
X_74551_ _74625_/A _74551_/X sky130_fd_sc_hd__buf_2
X_86537_ _86218_/CLK _48314_/Y _66256_/B sky130_fd_sc_hd__dfxtp_4
X_52929_ _52821_/A _52929_/X sky130_fd_sc_hd__buf_2
X_40943_ _40939_/X _40941_/X _88306_/Q _40942_/X _88306_/D sky130_fd_sc_hd__a2bb2o_4
X_71763_ _70504_/A _71763_/X sky130_fd_sc_hd__buf_2
X_83749_ _83749_/CLK _83749_/D _83749_/Q sky130_fd_sc_hd__dfxtp_4
X_59485_ _64236_/C _63384_/B sky130_fd_sc_hd__buf_2
X_56697_ _56725_/B _56687_/X _56696_/Y _56697_/X sky130_fd_sc_hd__o21a_4
X_73502_ _73502_/A _73501_/X _73502_/Y sky130_fd_sc_hd__nand2_4
X_70714_ _70714_/A _70713_/X _70710_/C _70710_/D _70714_/Y sky130_fd_sc_hd__nand4_4
X_46450_ _46450_/A _50460_/A sky130_fd_sc_hd__buf_2
X_58436_ _84848_/Q _63209_/A sky130_fd_sc_hd__inv_2
X_77270_ _77266_/X _77267_/Y _77269_/Y _77270_/X sky130_fd_sc_hd__a21o_4
X_43662_ _40723_/X _43659_/X _68959_/B _43661_/X _43663_/A sky130_fd_sc_hd__a2bb2o_4
X_55648_ _55647_/X _55676_/B _55648_/X sky130_fd_sc_hd__and2_4
X_74482_ _46725_/A _74501_/B sky130_fd_sc_hd__buf_2
X_86468_ _83311_/CLK _86468_/D _86468_/Q sky130_fd_sc_hd__dfxtp_4
X_40874_ _40873_/X _40874_/X sky130_fd_sc_hd__buf_2
X_71694_ _71691_/Y _83409_/Q _71693_/Y _83409_/D sky130_fd_sc_hd__a21o_4
X_45401_ _45596_/A _45401_/X sky130_fd_sc_hd__buf_2
X_76221_ _76219_/Y _76217_/X _76221_/C _76221_/Y sky130_fd_sc_hd__nand3_4
X_88207_ _87950_/CLK _41480_/X _88207_/Q sky130_fd_sc_hd__dfxtp_4
X_42613_ _49210_/B _40903_/A _41888_/X _42611_/Y _42612_/X _42613_/Y
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_5_12_0_CLK clkbuf_4_6_1_CLK/X clkbuf_6_25_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_73433_ _73434_/B _73434_/C _73432_/X _73433_/X sky130_fd_sc_hd__a21o_4
X_85419_ _85643_/CLK _54566_/Y _85419_/Q sky130_fd_sc_hd__dfxtp_4
X_46381_ _46348_/X _48996_/A _46380_/X _51294_/B sky130_fd_sc_hd__o21ai_4
X_70645_ _70714_/A _70639_/B _70642_/X _70638_/X _70645_/Y sky130_fd_sc_hd__nand4_4
X_58367_ _84867_/Q _63344_/A sky130_fd_sc_hd__inv_2
X_55579_ _45479_/A _44086_/A _55533_/X _55578_/X _55580_/B sky130_fd_sc_hd__a211o_4
X_43593_ _43611_/A _43593_/X sky130_fd_sc_hd__buf_2
X_86399_ _86398_/CLK _49375_/Y _58587_/B sky130_fd_sc_hd__dfxtp_4
X_48120_ _48138_/A _48329_/A _48120_/X sky130_fd_sc_hd__and2_4
X_57318_ _56766_/X _56782_/X _56810_/X _57318_/D _57318_/Y sky130_fd_sc_hd__nand4_4
X_45332_ _45331_/Y _45272_/X _45332_/Y sky130_fd_sc_hd__nand2_4
X_76152_ _76150_/A _81537_/Q _76150_/B _76152_/Y sky130_fd_sc_hd__nand3_4
X_88138_ _88394_/CLK _88138_/D _66802_/B sky130_fd_sc_hd__dfxtp_4
X_42544_ _42536_/X _42527_/X _40767_/X _42543_/Y _42538_/X _87827_/D
+ sky130_fd_sc_hd__o32ai_4
X_73364_ _73365_/B _73365_/C _73363_/X _73364_/X sky130_fd_sc_hd__a21o_4
X_70576_ _71162_/B _70412_/X _70933_/B _70423_/X _70576_/X sky130_fd_sc_hd__and4_4
X_58298_ _58298_/A _58298_/Y sky130_fd_sc_hd__inv_2
X_75103_ _75104_/C _75104_/B _75104_/A _75106_/A sky130_fd_sc_hd__a21oi_4
X_48051_ _83540_/Q _48051_/Y sky130_fd_sc_hd__inv_2
X_72315_ _72264_/X _85361_/Q _72314_/X _72315_/Y sky130_fd_sc_hd__o21ai_4
X_45263_ _55764_/B _45206_/X _45237_/X _45263_/X sky130_fd_sc_hd__o21a_4
X_57249_ _57340_/C _57249_/X sky130_fd_sc_hd__buf_2
X_76083_ _81528_/Q _76083_/B _81777_/D sky130_fd_sc_hd__xor2_4
X_88069_ _87813_/CLK _88069_/D _73124_/A sky130_fd_sc_hd__dfxtp_4
X_42475_ _42475_/A _42475_/Y sky130_fd_sc_hd__inv_2
X_73295_ _83157_/Q _73193_/X _73294_/Y _73295_/X sky130_fd_sc_hd__a21o_4
X_47002_ _47002_/A _47003_/A sky130_fd_sc_hd__buf_2
Xclkbuf_5_27_0_CLK clkbuf_5_27_0_CLK/A clkbuf_6_55_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_44214_ _44213_/X _44214_/X sky130_fd_sc_hd__buf_2
X_75034_ _75016_/Y _75032_/Y _75033_/Y _75049_/A sky130_fd_sc_hd__a21o_4
X_79911_ _79911_/A _79911_/Y sky130_fd_sc_hd__inv_2
X_41426_ _41425_/Y _88218_/D sky130_fd_sc_hd__inv_2
X_60260_ _60244_/A _60244_/B _79837_/A _60260_/Y sky130_fd_sc_hd__nor3_4
X_72246_ _57790_/X _72332_/B sky130_fd_sc_hd__buf_2
X_45194_ _45709_/A _45194_/X sky130_fd_sc_hd__buf_2
Xclkbuf_opt_16_CLK _84518_/CLK _84634_/CLK sky130_fd_sc_hd__clkbuf_16
X_44145_ _44143_/Y _44144_/Y _44163_/B _87186_/D sky130_fd_sc_hd__a21oi_4
X_79842_ _79839_/X _79842_/B _79842_/X sky130_fd_sc_hd__xor2_4
X_41357_ _41356_/X _41307_/X _67647_/B _41308_/X _88230_/D sky130_fd_sc_hd__a2bb2o_4
X_60191_ _60324_/B _60268_/A sky130_fd_sc_hd__buf_2
X_72177_ _72172_/X _72174_/Y _72175_/Y _59301_/X _72176_/X _72177_/X
+ sky130_fd_sc_hd__o32a_4
X_71128_ _50708_/B _71117_/X _71127_/Y _83597_/D sky130_fd_sc_hd__o21ai_4
X_48953_ _48898_/A _48964_/A sky130_fd_sc_hd__buf_2
X_44076_ _55159_/A _55761_/A sky130_fd_sc_hd__buf_2
X_79773_ _79763_/X _79765_/B _79772_/Y _79790_/B sky130_fd_sc_hd__a21boi_4
X_41288_ _41287_/Y _41288_/X sky130_fd_sc_hd__buf_2
X_76985_ _76985_/A _76985_/B _76985_/X sky130_fd_sc_hd__xor2_4
X_47904_ _47904_/A _47904_/X sky130_fd_sc_hd__buf_2
X_43027_ _43027_/A _43027_/Y sky130_fd_sc_hd__inv_2
X_78724_ _78722_/Y _78723_/Y _78720_/A _78725_/B sky130_fd_sc_hd__o21ai_4
X_63950_ _60871_/Y _64029_/B sky130_fd_sc_hd__buf_2
X_71059_ _48912_/B _71047_/X _71058_/Y _71059_/Y sky130_fd_sc_hd__o21ai_4
X_75936_ _75928_/A _75934_/Y _75935_/Y _75936_/Y sky130_fd_sc_hd__o21ai_4
X_48884_ _48884_/A _48885_/A sky130_fd_sc_hd__buf_2
X_62901_ _62791_/X _62930_/A sky130_fd_sc_hd__buf_2
X_47835_ _43585_/X _57491_/C _47834_/Y _47835_/X sky130_fd_sc_hd__o21a_4
X_78655_ _78653_/X _78655_/B _78655_/X sky130_fd_sc_hd__and2_4
X_63881_ _63879_/X _63833_/X _63880_/Y _84289_/D sky130_fd_sc_hd__a21oi_4
X_75867_ _75867_/A _75867_/Y sky130_fd_sc_hd__inv_2
X_65620_ _64967_/X _65621_/A sky130_fd_sc_hd__buf_2
X_77606_ _77606_/A _77605_/X _77622_/A sky130_fd_sc_hd__xnor2_4
X_62832_ _60362_/A _62869_/A sky130_fd_sc_hd__buf_2
X_74818_ _59426_/X _46111_/A _74818_/Y sky130_fd_sc_hd__nand2_4
X_47766_ _49379_/A _47804_/A sky130_fd_sc_hd__buf_2
X_78586_ _78586_/A _82677_/D _78586_/Y sky130_fd_sc_hd__nand2_4
X_44978_ _44962_/X _44974_/Y _44977_/Y _44978_/Y sky130_fd_sc_hd__a21oi_4
X_75798_ _75793_/B _75793_/A _75798_/X sky130_fd_sc_hd__and2_4
X_49505_ _49614_/A _49516_/B sky130_fd_sc_hd__buf_2
X_46717_ _46717_/A _46717_/B _46717_/C _46716_/X _46717_/X sky130_fd_sc_hd__and4_4
X_65551_ _65387_/A _65551_/B _65551_/X sky130_fd_sc_hd__and2_4
X_77537_ _77537_/A _77537_/B _77537_/Y sky130_fd_sc_hd__nor2_4
X_43929_ _43869_/X _43929_/X sky130_fd_sc_hd__buf_2
X_74749_ _74731_/A _74764_/A sky130_fd_sc_hd__buf_2
X_62763_ _61438_/X _62743_/B _62742_/X _62729_/D _62763_/Y sky130_fd_sc_hd__nand4_4
X_47697_ _72336_/A _47666_/X _47696_/Y _47697_/Y sky130_fd_sc_hd__o21ai_4
X_64502_ _64474_/X _64525_/B _62129_/X _64504_/C sky130_fd_sc_hd__nand3_4
X_49436_ _49447_/A _49447_/B _49420_/C _46744_/X _49436_/X sky130_fd_sc_hd__and4_4
X_61714_ _61714_/A _62128_/B _59608_/A _59761_/B _61714_/Y sky130_fd_sc_hd__nand4_4
X_68270_ _68246_/X _67649_/Y _68268_/X _68269_/Y _68270_/X sky130_fd_sc_hd__a211o_4
X_46648_ _46644_/Y _46598_/X _46647_/X _46648_/Y sky130_fd_sc_hd__a21oi_4
X_65482_ _65480_/Y _65448_/X _65481_/X _84198_/D sky130_fd_sc_hd__a21o_4
X_77468_ _77468_/A _77468_/B _77468_/Y sky130_fd_sc_hd__nand2_4
X_62694_ _61365_/X _62694_/B _62694_/C _62664_/D _62694_/Y sky130_fd_sc_hd__nand4_4
X_67221_ _67816_/A _67222_/A sky130_fd_sc_hd__buf_2
X_79207_ _79206_/Y _79207_/B _79208_/B sky130_fd_sc_hd__nand2_4
X_64433_ _64377_/A _64494_/A sky130_fd_sc_hd__buf_2
X_76419_ _76418_/X _76419_/Y sky130_fd_sc_hd__inv_2
X_49367_ _58576_/B _49360_/X _49366_/Y _49367_/Y sky130_fd_sc_hd__o21ai_4
X_61645_ _61645_/A _61645_/X sky130_fd_sc_hd__buf_2
X_46579_ _47972_/A _46579_/X sky130_fd_sc_hd__buf_2
X_77399_ _77386_/B _77398_/Y _77399_/Y sky130_fd_sc_hd__nand2_4
X_48318_ _48316_/Y _48302_/X _48317_/X _48318_/Y sky130_fd_sc_hd__a21oi_4
X_67152_ _66910_/A _67152_/X sky130_fd_sc_hd__buf_2
X_79138_ _79138_/A _79138_/B _79138_/X sky130_fd_sc_hd__xor2_4
X_64364_ _64319_/X _64364_/B _64333_/X _64364_/X sky130_fd_sc_hd__and3_4
X_49298_ _49296_/Y _49271_/X _49297_/Y _86415_/D sky130_fd_sc_hd__a21boi_4
X_61576_ _61394_/A _61576_/X sky130_fd_sc_hd__buf_2
X_66103_ _66099_/X _66102_/X _66103_/Y sky130_fd_sc_hd__nand2_4
X_63315_ _63311_/Y _63312_/X _63313_/X _63314_/X _63242_/X _63315_/Y
+ sky130_fd_sc_hd__o41ai_4
X_48249_ _48244_/A _47969_/B _48249_/Y sky130_fd_sc_hd__nand2_4
X_60527_ _60523_/X _60481_/X _60524_/Y _60491_/X _60526_/Y _60527_/Y
+ sky130_fd_sc_hd__a41oi_4
X_67083_ _67133_/A _86785_/Q _67083_/X sky130_fd_sc_hd__and2_4
X_79069_ _79027_/B _79066_/X _79068_/X _79070_/B sky130_fd_sc_hd__a21boi_4
X_64295_ _64295_/A _64248_/B _64295_/C _64295_/X sky130_fd_sc_hd__and3_4
X_81100_ _82220_/CLK _79667_/X _81100_/Q sky130_fd_sc_hd__dfxtp_4
X_66034_ _66032_/Y _65987_/X _66033_/X _84161_/D sky130_fd_sc_hd__a21o_4
X_51260_ _51286_/A _51280_/A sky130_fd_sc_hd__buf_2
X_63246_ _79301_/A _63189_/X _63245_/Y _63246_/X sky130_fd_sc_hd__a21o_4
X_82080_ _81169_/CLK _84040_/Q _78009_/A sky130_fd_sc_hd__dfxtp_4
X_60458_ _60447_/A _60458_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_110_0_CLK clkbuf_6_55_0_CLK/X clkbuf_8_221_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_50211_ _50523_/A _50473_/A sky130_fd_sc_hd__buf_2
X_81031_ _81061_/CLK _81031_/D _81031_/Q sky130_fd_sc_hd__dfxtp_4
X_51191_ _51191_/A _51191_/X sky130_fd_sc_hd__buf_2
X_63177_ _58562_/A _63131_/X _63175_/X _58338_/Y _63176_/X _63177_/Y
+ sky130_fd_sc_hd__o32ai_4
X_60389_ _60606_/A _60473_/C sky130_fd_sc_hd__buf_2
Xclkbuf_10_80_0_CLK clkbuf_9_40_0_CLK/X _86772_/CLK sky130_fd_sc_hd__clkbuf_1
X_50142_ _50142_/A _50082_/B _50059_/C _50142_/X sky130_fd_sc_hd__and3_4
X_62128_ _62948_/C _62128_/B _62128_/C _59761_/B _62131_/C sky130_fd_sc_hd__nand4_4
X_67985_ _68028_/A _67985_/B _67985_/X sky130_fd_sc_hd__and2_4
X_69724_ _69720_/X _69723_/X _68697_/X _69727_/A sky130_fd_sc_hd__a21o_4
X_50073_ _50578_/A _50578_/B _47848_/X _50073_/X sky130_fd_sc_hd__o21a_4
X_54950_ _54927_/A _54955_/B sky130_fd_sc_hd__buf_2
X_66936_ _66912_/A _87620_/Q _66936_/X sky130_fd_sc_hd__and2_4
X_85770_ _85770_/CLK _52705_/Y _85770_/Q sky130_fd_sc_hd__dfxtp_4
X_62059_ _61704_/Y _62088_/B sky130_fd_sc_hd__buf_2
Xclkbuf_7_125_0_CLK clkbuf_6_62_0_CLK/X clkbuf_8_251_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_82982_ _83012_/CLK _82982_/D _82982_/Q sky130_fd_sc_hd__dfxtp_4
X_53901_ _53929_/A _53902_/A sky130_fd_sc_hd__buf_2
X_84721_ _83464_/CLK _84721_/D _84721_/Q sky130_fd_sc_hd__dfxtp_4
X_81933_ _81933_/CLK _81933_/D _77390_/A sky130_fd_sc_hd__dfxtp_4
X_69655_ _69655_/A _69655_/X sky130_fd_sc_hd__buf_2
X_54881_ _85360_/Q _54865_/X _54880_/Y _54881_/Y sky130_fd_sc_hd__o21ai_4
X_66867_ _69751_/A _66868_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_95_0_CLK clkbuf_9_47_0_CLK/X _84914_/CLK sky130_fd_sc_hd__clkbuf_1
X_56620_ _56587_/X _56619_/X _85144_/Q _56590_/X _56620_/X sky130_fd_sc_hd__a2bb2o_4
X_68606_ _68600_/X _68605_/X _68558_/X _68606_/X sky130_fd_sc_hd__a21o_4
X_87440_ _87952_/CLK _87440_/D _87440_/Q sky130_fd_sc_hd__dfxtp_4
X_53832_ _53819_/A _72007_/B _53832_/Y sky130_fd_sc_hd__nand2_4
X_65818_ _65815_/Y _65757_/X _65817_/X _84176_/D sky130_fd_sc_hd__a21o_4
X_84652_ _84652_/CLK _60146_/Y _60145_/A sky130_fd_sc_hd__dfxtp_4
X_81864_ _84375_/CLK _78055_/X _81864_/Q sky130_fd_sc_hd__dfxtp_4
X_69586_ _69586_/A _88338_/Q _69586_/X sky130_fd_sc_hd__and2_4
Xclkbuf_8_241_0_CLK clkbuf_8_241_0_CLK/A clkbuf_9_483_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_66798_ _66819_/A _86829_/Q _66798_/X sky130_fd_sc_hd__and2_4
X_83603_ _86155_/CLK _71111_/Y _49106_/A sky130_fd_sc_hd__dfxtp_4
X_56551_ _44037_/X _56551_/X sky130_fd_sc_hd__buf_2
X_80815_ _80991_/CLK _83959_/Q _75839_/B sky130_fd_sc_hd__dfxtp_4
X_87371_ _87373_/CLK _87371_/D _87371_/Q sky130_fd_sc_hd__dfxtp_4
X_68537_ _68532_/X _68536_/X _68512_/X _68537_/Y sky130_fd_sc_hd__a21oi_4
X_53763_ _53763_/A _53774_/C sky130_fd_sc_hd__buf_2
X_65749_ _65654_/X _86188_/Q _65576_/X _65748_/X _65749_/X sky130_fd_sc_hd__a211o_4
X_84583_ _84583_/CLK _60701_/Y _60700_/C sky130_fd_sc_hd__dfxtp_4
X_50975_ _50972_/Y _50957_/X _50974_/X _86097_/D sky130_fd_sc_hd__a21oi_4
X_81795_ _81284_/CLK _81795_/D _81795_/Q sky130_fd_sc_hd__dfxtp_4
X_55502_ _55501_/X _55503_/D sky130_fd_sc_hd__buf_2
X_86322_ _86322_/CLK _86322_/D _57934_/B sky130_fd_sc_hd__dfxtp_4
X_52714_ _85768_/Q _52711_/X _52713_/Y _52714_/Y sky130_fd_sc_hd__o21ai_4
X_59270_ _59270_/A _59282_/B _59270_/Y sky130_fd_sc_hd__nor2_4
X_83534_ _86534_/CLK _83534_/D _83534_/Q sky130_fd_sc_hd__dfxtp_4
X_56482_ _56035_/X _56468_/X _56481_/Y _85179_/D sky130_fd_sc_hd__o21ai_4
X_80746_ _80746_/CLK _75198_/X _81122_/D sky130_fd_sc_hd__dfxtp_4
X_68468_ _57804_/A _68468_/B _68468_/Y sky130_fd_sc_hd__nor2_4
X_53694_ _53611_/X _74437_/B _53694_/Y sky130_fd_sc_hd__nand2_4
X_58221_ _63376_/B _58221_/X sky130_fd_sc_hd__buf_2
X_55433_ _55423_/Y _55427_/Y _55421_/Y _55434_/B sky130_fd_sc_hd__a21boi_4
X_67419_ _67416_/X _67418_/X _67322_/X _67419_/X sky130_fd_sc_hd__a21o_4
X_86253_ _83303_/CLK _50157_/Y _86253_/Q sky130_fd_sc_hd__dfxtp_4
X_52645_ _52637_/A _52645_/B _52645_/Y sky130_fd_sc_hd__nand2_4
X_83465_ _83464_/CLK _83465_/D _83465_/Q sky130_fd_sc_hd__dfxtp_4
X_80677_ _82211_/CLK _80709_/Q _75109_/A sky130_fd_sc_hd__dfxtp_4
X_68399_ _67013_/X _70001_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_251_0_CLK clkbuf_9_125_0_CLK/X _81839_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_503 sky130_fd_sc_hd__decap_3
XPHY_514 sky130_fd_sc_hd__decap_3
X_85204_ _85168_/CLK _85204_/D _85204_/Q sky130_fd_sc_hd__dfxtp_4
X_70430_ _71196_/A _70431_/C sky130_fd_sc_hd__buf_2
X_58152_ _46158_/B _63380_/A _58151_/Y _84920_/D sky130_fd_sc_hd__a21oi_4
X_82416_ _82462_/CLK _82448_/Q _78503_/A sky130_fd_sc_hd__dfxtp_4
XPHY_525 sky130_fd_sc_hd__decap_3
Xclkbuf_10_881_0_CLK clkbuf_9_440_0_CLK/X _86029_/CLK sky130_fd_sc_hd__clkbuf_1
X_55364_ _56708_/A _56708_/C _55392_/B sky130_fd_sc_hd__nand2_4
X_86184_ _86500_/CLK _50527_/Y _86184_/Q sky130_fd_sc_hd__dfxtp_4
X_40590_ _40590_/A _40590_/X sky130_fd_sc_hd__buf_2
X_52576_ _52602_/A _52590_/A sky130_fd_sc_hd__buf_2
XPHY_536 sky130_fd_sc_hd__decap_3
X_83396_ _83431_/CLK _83396_/D _83396_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_547 sky130_fd_sc_hd__decap_3
XPHY_558 sky130_fd_sc_hd__decap_3
Xclkbuf_10_33_0_CLK clkbuf_9_16_0_CLK/X _85114_/CLK sky130_fd_sc_hd__clkbuf_1
X_57103_ _57097_/X _56584_/X _45455_/A _57099_/X _85085_/D sky130_fd_sc_hd__a2bb2o_4
X_54315_ _85464_/Q _54294_/X _54314_/Y _54315_/Y sky130_fd_sc_hd__o21ai_4
XPHY_569 sky130_fd_sc_hd__decap_3
X_85135_ _85067_/CLK _85135_/D _85135_/Q sky130_fd_sc_hd__dfxtp_4
X_51527_ _51521_/X _51527_/B _51533_/C _53052_/D _51527_/X sky130_fd_sc_hd__and4_4
X_58083_ _58701_/A _58083_/X sky130_fd_sc_hd__buf_2
X_70361_ _70361_/A _70361_/Y sky130_fd_sc_hd__inv_2
X_82347_ _82859_/CLK _77118_/X _48064_/A sky130_fd_sc_hd__dfxtp_4
X_55295_ _55156_/X _55160_/X _83746_/Q _55296_/A sky130_fd_sc_hd__a21o_4
Xclkbuf_9_372_0_CLK clkbuf_9_373_0_CLK/A clkbuf_9_372_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_72100_ _72097_/Y _72083_/X _72099_/Y _83285_/D sky130_fd_sc_hd__a21boi_4
X_57034_ _57019_/A _57024_/Y _57034_/C _57034_/Y sky130_fd_sc_hd__nand3_4
X_42260_ _41465_/X _42258_/X _87954_/Q _42259_/X _87954_/D sky130_fd_sc_hd__a2bb2o_4
X_54246_ _54329_/A _54246_/X sky130_fd_sc_hd__buf_2
X_85066_ _83335_/CLK _57190_/Y _85066_/Q sky130_fd_sc_hd__dfxtp_4
X_73080_ _57376_/X _73104_/B sky130_fd_sc_hd__buf_2
X_51458_ _51539_/A _51458_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_266_0_CLK clkbuf_9_133_0_CLK/X _84714_/CLK sky130_fd_sc_hd__clkbuf_1
X_70292_ _70292_/A _70292_/B _70292_/C _70292_/D _70292_/X sky130_fd_sc_hd__and4_4
X_82278_ _82284_/CLK _77023_/B _41085_/A sky130_fd_sc_hd__dfxtp_4
X_41211_ _41210_/Y _88257_/D sky130_fd_sc_hd__inv_2
X_72031_ _72017_/X _53856_/B _72031_/Y sky130_fd_sc_hd__nand2_4
X_84017_ _84014_/CLK _84017_/D _82057_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_896_0_CLK clkbuf_9_448_0_CLK/X _87345_/CLK sky130_fd_sc_hd__clkbuf_1
X_50409_ _50406_/Y _50395_/X _50408_/X _86207_/D sky130_fd_sc_hd__a21oi_4
X_81229_ _81227_/CLK _81229_/D _81229_/Q sky130_fd_sc_hd__dfxtp_4
X_42191_ _41288_/X _42183_/X _87987_/Q _42184_/X _87987_/D sky130_fd_sc_hd__a2bb2o_4
X_54177_ _54160_/A _54186_/B _54191_/C _53008_/D _54177_/X sky130_fd_sc_hd__and4_4
X_51389_ _51758_/A _51389_/B _51389_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_48_0_CLK clkbuf_9_24_0_CLK/X _85074_/CLK sky130_fd_sc_hd__clkbuf_1
X_41142_ _40380_/A _41143_/A sky130_fd_sc_hd__buf_2
X_53128_ _85692_/Q _53120_/X _53127_/Y _53128_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_387_0_CLK clkbuf_9_387_0_CLK/A clkbuf_9_387_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_58985_ _58985_/A _58988_/B _58985_/Y sky130_fd_sc_hd__nand2_4
X_45950_ _45950_/A _45950_/B _44210_/X _45950_/Y sky130_fd_sc_hd__nor3_4
X_41073_ _41072_/X _41073_/X sky130_fd_sc_hd__buf_2
X_53059_ _53055_/Y _53056_/X _53058_/X _53059_/Y sky130_fd_sc_hd__a21oi_4
X_57936_ _57868_/X _57934_/Y _57935_/Y _57899_/X _57872_/X _57936_/X
+ sky130_fd_sc_hd__o32a_4
X_76770_ _76770_/A _76769_/Y _76771_/B sky130_fd_sc_hd__xnor2_4
X_73982_ _73367_/A _73982_/X sky130_fd_sc_hd__buf_2
X_85968_ _85679_/CLK _51670_/Y _85968_/Q sky130_fd_sc_hd__dfxtp_4
X_44901_ _45819_/A _44901_/X sky130_fd_sc_hd__buf_2
X_75721_ _80913_/Q _80785_/D _75720_/X _75722_/B sky130_fd_sc_hd__o21ai_4
X_87707_ _87195_/CLK _42810_/X _67901_/B sky130_fd_sc_hd__dfxtp_4
X_72933_ _72750_/X _85595_/Q _72839_/X _72932_/X _72933_/X sky130_fd_sc_hd__a211o_4
X_84919_ _84905_/CLK _84919_/D _58154_/A sky130_fd_sc_hd__dfxtp_4
X_45881_ _44196_/A _45882_/A sky130_fd_sc_hd__buf_2
X_57867_ _58827_/A _58696_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_310_0_CLK clkbuf_9_311_0_CLK/A clkbuf_9_310_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_85899_ _86210_/CLK _52051_/Y _85899_/Q sky130_fd_sc_hd__dfxtp_4
X_47620_ _57563_/A _47620_/X sky130_fd_sc_hd__buf_2
X_59606_ _59605_/Y _59637_/A sky130_fd_sc_hd__buf_2
X_78440_ _78439_/Y _78450_/B sky130_fd_sc_hd__inv_2
Xclkbuf_8_209_0_CLK clkbuf_8_209_0_CLK/A clkbuf_9_419_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_44832_ _45980_/A _44832_/X sky130_fd_sc_hd__buf_2
X_56818_ _45882_/A _56670_/A _56817_/X _56818_/X sky130_fd_sc_hd__a21o_4
X_75652_ _75638_/A _75637_/Y _75652_/Y sky130_fd_sc_hd__nor2_4
X_87638_ _87189_/CLK _87638_/D _68018_/B sky130_fd_sc_hd__dfxtp_4
X_72864_ _73124_/B _73370_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_204_0_CLK clkbuf_9_102_0_CLK/X _84269_/CLK sky130_fd_sc_hd__clkbuf_1
X_57798_ _46210_/A _57866_/A sky130_fd_sc_hd__buf_2
X_74603_ _74591_/X _74599_/X _56130_/A _74600_/X _74603_/X sky130_fd_sc_hd__a211o_4
X_47551_ _83710_/Q _47552_/A sky130_fd_sc_hd__inv_2
Xclkbuf_10_834_0_CLK clkbuf_9_417_0_CLK/X _84231_/CLK sky130_fd_sc_hd__clkbuf_1
X_71815_ _71813_/A _71815_/B _71049_/A _71815_/X sky130_fd_sc_hd__and3_4
X_59537_ _59537_/A _59662_/B sky130_fd_sc_hd__inv_2
X_78371_ _78373_/A _82663_/D _78371_/Y sky130_fd_sc_hd__nor2_4
X_44763_ _41327_/Y _44754_/X _86967_/Q _44755_/X _86967_/D sky130_fd_sc_hd__a2bb2o_4
X_56749_ _56713_/A _57149_/D _56739_/A _56749_/X sky130_fd_sc_hd__a21o_4
X_75583_ _75583_/A _75583_/Y sky130_fd_sc_hd__inv_2
X_87569_ _85895_/CLK _43118_/Y _87569_/Q sky130_fd_sc_hd__dfxtp_4
X_41975_ _42477_/A _41975_/X sky130_fd_sc_hd__buf_2
X_72795_ _72795_/A _73000_/B sky130_fd_sc_hd__buf_2
X_46502_ _46491_/A _51350_/B _46502_/Y sky130_fd_sc_hd__nand2_4
X_77322_ _81928_/Q _82184_/D _77322_/X sky130_fd_sc_hd__xor2_4
X_43714_ _40853_/X _43698_/X _69793_/B _43700_/X _43715_/A sky130_fd_sc_hd__a2bb2o_4
X_74534_ _52833_/B _74516_/X _74533_/Y _74534_/Y sky130_fd_sc_hd__o21ai_4
X_40926_ _40925_/X _40904_/X _69961_/B _40905_/X _40926_/X sky130_fd_sc_hd__a2bb2o_4
X_47482_ _47517_/A _53072_/B _47482_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_325_0_CLK clkbuf_9_325_0_CLK/A clkbuf_9_325_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_71746_ _70635_/A _71753_/B sky130_fd_sc_hd__buf_2
X_59468_ _59467_/Y _59478_/B _59468_/Y sky130_fd_sc_hd__nand2_4
X_44694_ _44694_/A _44694_/Y sky130_fd_sc_hd__inv_2
X_49221_ _49219_/Y _49214_/X _49220_/Y _86431_/D sky130_fd_sc_hd__a21boi_4
X_46433_ _46433_/A _51316_/B sky130_fd_sc_hd__buf_2
X_58419_ _58406_/X _83365_/Q _58418_/Y _58419_/X sky130_fd_sc_hd__o21a_4
X_77253_ _77253_/A _77253_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_219_0_CLK clkbuf_9_109_0_CLK/X _84507_/CLK sky130_fd_sc_hd__clkbuf_1
X_43645_ _40691_/A _43634_/X _43644_/Y _43636_/X _43645_/X sky130_fd_sc_hd__a2bb2o_4
X_74465_ _74462_/Y _74463_/X _74464_/X _83061_/D sky130_fd_sc_hd__a21oi_4
X_40857_ _40783_/A _40857_/X sky130_fd_sc_hd__buf_2
X_71677_ _58476_/Y _71669_/X _71676_/Y _83415_/D sky130_fd_sc_hd__o21ai_4
X_59399_ _59399_/A _59399_/B _59399_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_849_0_CLK clkbuf_9_424_0_CLK/X _82206_/CLK sky130_fd_sc_hd__clkbuf_1
X_76204_ _76189_/A _76189_/B _76187_/Y _76205_/A sky130_fd_sc_hd__a21boi_4
X_49152_ _49146_/Y _49138_/X _49151_/X _86439_/D sky130_fd_sc_hd__a21oi_4
X_61430_ _61430_/A _61404_/X _61406_/C _61390_/D _61430_/Y sky130_fd_sc_hd__nand4_4
X_73416_ _42050_/Y _72974_/X _73393_/X _73415_/Y _73416_/X sky130_fd_sc_hd__a211o_4
X_46364_ _46279_/A _46364_/X sky130_fd_sc_hd__buf_2
X_70628_ HASH_ADDR[5] HASH_ADDR[4] _70668_/D sky130_fd_sc_hd__nor2_4
X_77184_ _77184_/A _77177_/A _77184_/X sky130_fd_sc_hd__and2_4
X_43576_ _43557_/X _43563_/X _40532_/X _87351_/Q _43058_/A _43577_/A
+ sky130_fd_sc_hd__o32ai_4
X_74396_ _74396_/A _74395_/X _74366_/C _74396_/X sky130_fd_sc_hd__and3_4
X_40788_ _40758_/X _40759_/X _40787_/X _69627_/B _40744_/X _40788_/Y
+ sky130_fd_sc_hd__o32ai_4
X_48103_ _48781_/A _48103_/X sky130_fd_sc_hd__buf_2
X_45315_ _85190_/Q _45252_/X _45314_/X _45315_/Y sky130_fd_sc_hd__o21ai_4
X_76135_ _76135_/A _76134_/Y _76136_/B sky130_fd_sc_hd__xor2_4
X_42527_ _42547_/A _42527_/X sky130_fd_sc_hd__buf_2
X_61361_ _61354_/Y _61357_/Y _61334_/X _61358_/Y _61360_/Y _61361_/X
+ sky130_fd_sc_hd__a41o_4
X_49083_ _49083_/A _50153_/B sky130_fd_sc_hd__buf_2
X_73347_ _72951_/A _73347_/X sky130_fd_sc_hd__buf_2
X_46295_ _46295_/A _46295_/X sky130_fd_sc_hd__buf_2
X_70559_ _70558_/X _70549_/X _70568_/C _70550_/D _70559_/Y sky130_fd_sc_hd__nor4_4
X_63100_ _63100_/A _63100_/B _63079_/C _63066_/D _63100_/X sky130_fd_sc_hd__and4_4
X_60312_ _59755_/A _59716_/A _60312_/C _60312_/D _60312_/Y sky130_fd_sc_hd__nand4_4
X_48034_ _48044_/A _48034_/B _48034_/Y sky130_fd_sc_hd__nand2_4
X_45246_ _45243_/X _45245_/Y _45200_/X _45246_/Y sky130_fd_sc_hd__a21oi_4
X_64080_ _60926_/X _64179_/D sky130_fd_sc_hd__buf_2
X_76066_ _76065_/Y _76063_/C _76066_/X sky130_fd_sc_hd__and2_4
X_42458_ _51238_/B _42430_/X _40581_/X _87857_/Q _42453_/X _42458_/Y
+ sky130_fd_sc_hd__o32ai_4
X_61292_ _61292_/A _61329_/A sky130_fd_sc_hd__buf_2
X_73278_ _44189_/X _74246_/B sky130_fd_sc_hd__buf_2
X_63031_ _63025_/Y _63026_/X _63029_/X _63030_/X _63020_/X _63031_/Y
+ sky130_fd_sc_hd__o41ai_4
X_75017_ _75016_/Y _75017_/Y sky130_fd_sc_hd__inv_2
X_41409_ _41399_/X _41400_/X _41408_/X _88220_/Q _41388_/X _41410_/A
+ sky130_fd_sc_hd__o32ai_4
X_60243_ _60525_/A _60244_/B sky130_fd_sc_hd__buf_2
X_72229_ _72155_/X _85688_/Q _72156_/X _72229_/X sky130_fd_sc_hd__o21a_4
X_45177_ _55823_/B _45134_/X _45116_/X _45177_/X sky130_fd_sc_hd__o21a_4
X_42389_ _41911_/A _42389_/X sky130_fd_sc_hd__buf_2
X_44128_ _44127_/X _44128_/X sky130_fd_sc_hd__buf_2
X_79825_ _84228_/Q _83276_/Q _79825_/X sky130_fd_sc_hd__xor2_4
X_60174_ _72625_/B _72625_/A _60174_/C _60174_/D _60174_/X sky130_fd_sc_hd__and4_4
X_49985_ _49982_/Y _49977_/X _49984_/X _49985_/Y sky130_fd_sc_hd__a21oi_4
X_48936_ _48936_/A _48699_/B _48936_/Y sky130_fd_sc_hd__nand2_4
X_44059_ _44059_/A _44059_/X sky130_fd_sc_hd__buf_2
X_67770_ _68402_/A _67770_/X sky130_fd_sc_hd__buf_2
X_79756_ _79761_/A _79761_/B _79756_/Y sky130_fd_sc_hd__xnor2_4
X_64982_ _44150_/X _86739_/Q _64980_/X _64981_/X _64982_/X sky130_fd_sc_hd__a211o_4
X_76968_ _76967_/Y _76968_/Y sky130_fd_sc_hd__inv_2
X_66721_ _66651_/A _87629_/Q _66721_/X sky130_fd_sc_hd__and2_4
X_78707_ _78707_/A _82780_/D _82492_/D sky130_fd_sc_hd__xor2_4
X_63933_ _61483_/A _63947_/B _63947_/C _63866_/X _63933_/Y sky130_fd_sc_hd__nand4_4
X_75919_ _84517_/Q _84389_/Q _80733_/D sky130_fd_sc_hd__xor2_4
X_48867_ _48864_/Y _48865_/X _48866_/X _86468_/D sky130_fd_sc_hd__a21oi_4
X_79687_ _79704_/B _79686_/Y _79687_/X sky130_fd_sc_hd__xor2_4
X_76899_ _76899_/A _76899_/B _76899_/Y sky130_fd_sc_hd__nor2_4
X_69440_ _69286_/A _87773_/Q _69440_/X sky130_fd_sc_hd__and2_4
X_47818_ _47818_/A _53259_/B sky130_fd_sc_hd__buf_2
X_78638_ _78638_/A _78638_/B _78639_/A sky130_fd_sc_hd__and2_4
X_66652_ _87952_/Q _66562_/X _66564_/X _66651_/X _66652_/X sky130_fd_sc_hd__a211o_4
X_63864_ _63848_/X _63849_/X _63864_/C _63864_/Y sky130_fd_sc_hd__nor3_4
X_48798_ _48794_/Y _48785_/X _48797_/X _86481_/D sky130_fd_sc_hd__a21oi_4
X_65603_ _64739_/A _65634_/A sky130_fd_sc_hd__buf_2
X_62815_ _62810_/Y _62772_/X _62812_/Y _62813_/Y _62814_/X _62815_/X
+ sky130_fd_sc_hd__a41o_4
X_69371_ _69371_/A _69371_/X sky130_fd_sc_hd__buf_2
X_47749_ _47758_/A _47777_/B _47749_/C _53223_/D _47749_/X sky130_fd_sc_hd__and4_4
X_66583_ _66683_/A _66583_/B _66583_/X sky130_fd_sc_hd__and2_4
X_78569_ _78569_/A _78569_/B _78569_/C _78569_/X sky130_fd_sc_hd__or3_4
X_63795_ _64032_/A _63860_/B sky130_fd_sc_hd__buf_2
X_80600_ _80554_/Y _80594_/X _80599_/Y _80600_/Y sky130_fd_sc_hd__a21oi_4
X_68322_ _83983_/Q _68318_/X _68321_/X _83983_/D sky130_fd_sc_hd__a21bo_4
X_65534_ _65400_/A _65534_/X sky130_fd_sc_hd__buf_2
X_50760_ _50758_/Y _50735_/X _50759_/Y _86139_/D sky130_fd_sc_hd__a21boi_4
X_62746_ _62739_/Y _62713_/X _62740_/Y _62743_/Y _62745_/X _62746_/X
+ sky130_fd_sc_hd__a41o_4
X_81580_ _81352_/CLK _84180_/Q _76745_/A sky130_fd_sc_hd__dfxtp_4
X_49419_ _58687_/B _49415_/X _49418_/Y _49419_/Y sky130_fd_sc_hd__o21ai_4
X_80531_ _80531_/A _80531_/B _80531_/X sky130_fd_sc_hd__or2_4
X_68253_ _82648_/D _68238_/X _68252_/X _68253_/X sky130_fd_sc_hd__a21bo_4
X_65465_ _65929_/A _65546_/B sky130_fd_sc_hd__buf_2
X_50691_ _86152_/Q _50680_/X _50690_/Y _50691_/Y sky130_fd_sc_hd__o21ai_4
X_62677_ _58225_/X _60221_/A _60205_/X _60263_/C _62676_/X _62677_/Y
+ sky130_fd_sc_hd__a41oi_4
X_67204_ _67203_/X _67204_/X sky130_fd_sc_hd__buf_2
X_52430_ _52462_/A _52430_/X sky130_fd_sc_hd__buf_2
X_64416_ _64409_/Y _64415_/X _64386_/X _64416_/X sky130_fd_sc_hd__o21a_4
X_83250_ _85317_/CLK _83250_/D _83250_/Q sky130_fd_sc_hd__dfxtp_4
X_61628_ _59427_/A _61629_/B sky130_fd_sc_hd__buf_2
X_80462_ _80456_/A _80456_/B _80461_/Y _80478_/A sky130_fd_sc_hd__a21boi_4
X_68184_ _67159_/X _67162_/X _68173_/X _68184_/Y sky130_fd_sc_hd__a21oi_4
X_65396_ _84203_/Q _65397_/C sky130_fd_sc_hd__inv_2
X_82201_ _86104_/CLK _82201_/D _82393_/D sky130_fd_sc_hd__dfxtp_4
X_67135_ _67132_/X _67134_/X _67085_/X _67135_/X sky130_fd_sc_hd__a21o_4
X_52361_ _52358_/Y _52340_/X _52360_/X _85838_/D sky130_fd_sc_hd__a21oi_4
X_64347_ _58322_/Y _64308_/X _64346_/Y _64347_/Y sky130_fd_sc_hd__o21ai_4
X_83181_ _81696_/CLK _72713_/X _83181_/Q sky130_fd_sc_hd__dfxtp_4
X_80393_ _80406_/B _80406_/A _80393_/X sky130_fd_sc_hd__xor2_4
X_61559_ _84862_/Q _61560_/B sky130_fd_sc_hd__buf_2
X_54100_ _54123_/A _53428_/X _54111_/C _52934_/D _54100_/X sky130_fd_sc_hd__and4_4
X_51312_ _65002_/B _51309_/X _51311_/Y _51312_/Y sky130_fd_sc_hd__o21ai_4
X_82132_ _81970_/CLK _82132_/D _82132_/Q sky130_fd_sc_hd__dfxtp_4
X_55080_ _55093_/A _47741_/Y _55080_/Y sky130_fd_sc_hd__nand2_4
X_67066_ _67061_/X _67065_/X _66871_/X _67066_/Y sky130_fd_sc_hd__a21oi_4
X_52292_ _52288_/Y _52289_/X _52291_/X _52292_/Y sky130_fd_sc_hd__a21oi_4
X_64278_ _59467_/Y _64249_/X _64277_/Y _64278_/Y sky130_fd_sc_hd__o21ai_4
X_54031_ _54031_/A _50816_/B _54031_/Y sky130_fd_sc_hd__nand2_4
X_66017_ _65888_/A _65888_/B _66016_/Y _66017_/Y sky130_fd_sc_hd__nor3_4
X_51243_ _51241_/Y _51237_/X _51242_/X _51243_/Y sky130_fd_sc_hd__a21oi_4
X_63229_ _63053_/A _63316_/B sky130_fd_sc_hd__buf_2
X_86940_ _87922_/CLK _44813_/X _67417_/B sky130_fd_sc_hd__dfxtp_4
X_82063_ _83933_/CLK _84023_/Q _82063_/Q sky130_fd_sc_hd__dfxtp_4
X_81014_ _84197_/CLK _84222_/Q _81014_/Q sky130_fd_sc_hd__dfxtp_4
X_51174_ _86060_/Q _51156_/X _51173_/Y _51174_/Y sky130_fd_sc_hd__o21ai_4
X_86871_ _86882_/CLK _45532_/Y _63100_/B sky130_fd_sc_hd__dfxtp_4
X_50125_ _86259_/Q _50113_/X _50124_/Y _50125_/Y sky130_fd_sc_hd__o21ai_4
X_85822_ _85822_/CLK _52443_/Y _85822_/Q sky130_fd_sc_hd__dfxtp_4
X_58770_ _58756_/X _85937_/Q _58664_/X _58770_/X sky130_fd_sc_hd__o21a_4
X_55982_ _44917_/A _55690_/X _44102_/X _55981_/X _55983_/B sky130_fd_sc_hd__a211o_4
X_67968_ _87141_/Q _67942_/X _67872_/X _67967_/X _67968_/X sky130_fd_sc_hd__a211o_4
X_57721_ _44151_/X _57721_/B _57721_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_7_40_0_CLK clkbuf_7_41_0_CLK/A clkbuf_8_81_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_69707_ _81975_/D _69696_/X _69706_/X _83903_/D sky130_fd_sc_hd__a21bo_4
X_50056_ _50056_/A _48889_/B _50056_/Y sky130_fd_sc_hd__nand2_4
X_54933_ _54931_/Y _54909_/X _54932_/X _85351_/D sky130_fd_sc_hd__a21oi_4
X_66919_ _57866_/A _66919_/X sky130_fd_sc_hd__buf_2
X_85753_ _85754_/CLK _52798_/Y _85753_/Q sky130_fd_sc_hd__dfxtp_4
X_82965_ _82965_/CLK _82773_/Q _46735_/A sky130_fd_sc_hd__dfxtp_4
X_67899_ _67782_/X _67887_/Y _67863_/X _67898_/Y _67899_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_8_180_0_CLK clkbuf_7_90_0_CLK/X clkbuf_8_180_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_84704_ _84713_/CLK _84704_/D _80526_/A sky130_fd_sc_hd__dfxtp_4
X_57652_ _84961_/Q _57652_/X sky130_fd_sc_hd__buf_2
X_81916_ _82008_/CLK _81916_/D _81916_/Q sky130_fd_sc_hd__dfxtp_4
X_69638_ _69586_/A _88334_/Q _69638_/X sky130_fd_sc_hd__and2_4
X_54864_ _54860_/Y _54856_/X _54863_/X _85364_/D sky130_fd_sc_hd__a21oi_4
X_85684_ _84787_/CLK _85684_/D _85684_/Q sky130_fd_sc_hd__dfxtp_4
X_82896_ _82896_/CLK _78182_/B _41719_/A sky130_fd_sc_hd__dfxtp_4
X_56603_ _44135_/X _56696_/B sky130_fd_sc_hd__buf_2
X_87423_ _87421_/CLK _87423_/D _87423_/Q sky130_fd_sc_hd__dfxtp_4
X_53815_ _53813_/Y _53799_/X _53814_/Y _53815_/Y sky130_fd_sc_hd__a21boi_4
X_84635_ _84645_/CLK _60318_/Y _79733_/A sky130_fd_sc_hd__dfxtp_4
X_57583_ _57579_/Y _57581_/X _57582_/Y _57583_/Y sky130_fd_sc_hd__a21boi_4
X_81847_ _82221_/CLK _81879_/Q _77532_/A sky130_fd_sc_hd__dfxtp_4
X_69569_ _41980_/A _69442_/X _69567_/X _69568_/Y _69569_/X sky130_fd_sc_hd__a211o_4
X_54795_ _54791_/Y _54774_/X _54794_/X _85377_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_7_55_0_CLK clkbuf_7_55_0_CLK/A clkbuf_7_55_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_59322_ _59286_/X _86055_/Q _59321_/X _59322_/Y sky130_fd_sc_hd__o21ai_4
X_71600_ _71576_/X _71626_/B _71598_/C _71600_/Y sky130_fd_sc_hd__nor3_4
X_56534_ _56148_/X _56528_/X _56533_/Y _56534_/Y sky130_fd_sc_hd__o21ai_4
X_87354_ _81182_/CLK _87354_/D _87354_/Q sky130_fd_sc_hd__dfxtp_4
X_41760_ _40414_/X _41422_/A _41760_/X sky130_fd_sc_hd__or2_4
X_53746_ _85576_/Q _53729_/X _53745_/Y _53746_/Y sky130_fd_sc_hd__o21ai_4
X_72580_ _64561_/A _72581_/A sky130_fd_sc_hd__buf_2
X_84566_ _84583_/CLK _84566_/D _84566_/Q sky130_fd_sc_hd__dfxtp_4
X_50958_ _50929_/A _50963_/B sky130_fd_sc_hd__buf_2
Xclkbuf_8_195_0_CLK clkbuf_7_97_0_CLK/X clkbuf_9_391_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_81778_ _82053_/CLK _76090_/X _81778_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_190_0_CLK clkbuf_9_95_0_CLK/X _81038_/CLK sky130_fd_sc_hd__clkbuf_1
X_86305_ _86303_/CLK _49890_/Y _72116_/B sky130_fd_sc_hd__dfxtp_4
X_40711_ _40670_/X _40883_/A _40710_/X _40712_/A sky130_fd_sc_hd__o21ai_4
X_59253_ _58918_/A _59253_/X sky130_fd_sc_hd__buf_2
X_71531_ _71530_/Y _71531_/X sky130_fd_sc_hd__buf_2
X_83517_ _83520_/CLK _83517_/D _83517_/Q sky130_fd_sc_hd__dfxtp_4
X_56465_ _56545_/A _56454_/B _85185_/Q _56465_/Y sky130_fd_sc_hd__nand3_4
X_80729_ _80728_/CLK _75915_/X _80729_/Q sky130_fd_sc_hd__dfxtp_4
X_41691_ _82902_/Q _41660_/X _41691_/X sky130_fd_sc_hd__or2_4
X_87285_ _87285_/CLK _43748_/X _73509_/A sky130_fd_sc_hd__dfxtp_4
X_53677_ _53675_/Y _53653_/X _53676_/X _53677_/Y sky130_fd_sc_hd__a21oi_4
X_84497_ _84559_/CLK _61255_/X _75899_/A sky130_fd_sc_hd__dfxtp_4
X_50889_ _86112_/Q _50882_/X _50888_/Y _50889_/Y sky130_fd_sc_hd__o21ai_4
X_58204_ _83372_/Q _58204_/Y sky130_fd_sc_hd__inv_2
XPHY_300 sky130_fd_sc_hd__decap_3
X_43430_ _41556_/X _43412_/X _87425_/Q _43413_/X _87425_/D sky130_fd_sc_hd__a2bb2o_4
X_55416_ _55373_/Y _55297_/X _55416_/Y sky130_fd_sc_hd__nand2_4
X_74250_ _44747_/Y _56183_/X _74249_/Y _74250_/X sky130_fd_sc_hd__a21o_4
X_86236_ _84991_/CLK _50263_/Y _86236_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_311 sky130_fd_sc_hd__decap_3
X_40642_ _40635_/X _40638_/X _40641_/X _68595_/B _40612_/X _40643_/A
+ sky130_fd_sc_hd__o32ai_4
X_52628_ _52625_/Y _52619_/X _52627_/X _85784_/D sky130_fd_sc_hd__a21oi_4
X_59184_ _59146_/X _85426_/Q _59183_/X _59184_/Y sky130_fd_sc_hd__o21ai_4
X_71462_ _70426_/A _71462_/B _71463_/A sky130_fd_sc_hd__and2_4
X_83448_ _83480_/CLK _83448_/D _83448_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_322 sky130_fd_sc_hd__decap_3
X_56396_ _56040_/X _56394_/X _56395_/Y _85210_/D sky130_fd_sc_hd__o21ai_4
XPHY_333 sky130_fd_sc_hd__decap_3
XPHY_344 sky130_fd_sc_hd__decap_3
X_73201_ _73197_/X _73199_/X _73200_/X _73220_/B sky130_fd_sc_hd__a21o_4
X_58135_ _58576_/A _58135_/B _58135_/Y sky130_fd_sc_hd__nor2_4
X_70413_ HASH_ADDR[3] _70694_/A sky130_fd_sc_hd__buf_2
XPHY_355 sky130_fd_sc_hd__decap_3
X_43361_ _41367_/X _43356_/X _87460_/Q _43357_/X _87460_/D sky130_fd_sc_hd__a2bb2o_4
X_55347_ _45647_/A _44060_/X _55301_/X _55346_/Y _55347_/X sky130_fd_sc_hd__a211o_4
X_86167_ _85561_/CLK _50616_/Y _86167_/Q sky130_fd_sc_hd__dfxtp_4
X_74181_ _74181_/A _74181_/B _74181_/Y sky130_fd_sc_hd__xnor2_4
X_40573_ _40573_/A _40573_/X sky130_fd_sc_hd__buf_2
XPHY_366 sky130_fd_sc_hd__decap_3
X_52559_ _52567_/A _54077_/B _52559_/Y sky130_fd_sc_hd__nand2_4
X_83379_ _83414_/CLK _83379_/D _83379_/Q sky130_fd_sc_hd__dfxtp_4
X_71393_ _70692_/A _71386_/B _71399_/C _71393_/Y sky130_fd_sc_hd__nor3_4
XPHY_377 sky130_fd_sc_hd__decap_3
X_45100_ _55865_/B _45056_/X _45087_/X _45100_/X sky130_fd_sc_hd__o21a_4
XPHY_388 sky130_fd_sc_hd__decap_3
X_42312_ _42312_/A _87927_/D sky130_fd_sc_hd__inv_2
X_73132_ _73132_/A _85875_/Q _73132_/X sky130_fd_sc_hd__and2_4
X_85118_ _85152_/CLK _85118_/D _45440_/A sky130_fd_sc_hd__dfxtp_4
XPHY_399 sky130_fd_sc_hd__decap_3
X_46080_ _46080_/A _46080_/Y sky130_fd_sc_hd__inv_2
X_58066_ _58065_/X _85704_/Q _58020_/X _58066_/X sky130_fd_sc_hd__o21a_4
X_70344_ _70348_/A _70348_/B _83085_/Q _70348_/D _70344_/X sky130_fd_sc_hd__and4_4
X_43292_ _43292_/A _87495_/D sky130_fd_sc_hd__inv_2
X_55278_ _55278_/A _45792_/Y _55278_/Y sky130_fd_sc_hd__nor2_4
X_86098_ _85459_/CLK _50970_/Y _86098_/Q sky130_fd_sc_hd__dfxtp_4
X_45031_ _55913_/B _44963_/X _45004_/X _45031_/X sky130_fd_sc_hd__o21a_4
X_57017_ _57017_/A _85101_/D sky130_fd_sc_hd__inv_2
X_42243_ _42199_/X _42243_/X sky130_fd_sc_hd__buf_2
X_54229_ _54224_/Y _54226_/X _54228_/X _85481_/D sky130_fd_sc_hd__a21oi_4
X_73063_ _73132_/A _85878_/Q _73063_/X sky130_fd_sc_hd__and2_4
X_77940_ _82072_/Q _81944_/D _77939_/Y _77940_/Y sky130_fd_sc_hd__a21oi_4
X_85049_ _85049_/CLK _57255_/Y _57254_/B sky130_fd_sc_hd__dfxtp_4
X_70275_ _70267_/A _70267_/B _70275_/C _70264_/X _70275_/X sky130_fd_sc_hd__and4_4
Xclkbuf_8_133_0_CLK clkbuf_7_66_0_CLK/X clkbuf_9_267_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_72014_ _71993_/X _72014_/B _72014_/Y sky130_fd_sc_hd__nand2_4
X_42174_ _42173_/X _42169_/X _41225_/X _87998_/Q _42170_/X _42175_/A
+ sky130_fd_sc_hd__o32ai_4
X_77871_ _82066_/Q _77885_/A sky130_fd_sc_hd__inv_2
X_79610_ _79610_/A _79599_/Y _79611_/B sky130_fd_sc_hd__nand2_4
X_41125_ _41124_/X _41125_/X sky130_fd_sc_hd__buf_2
X_76822_ _76822_/A _76821_/Y _76825_/A sky130_fd_sc_hd__xor2_4
X_49770_ _49769_/X _52986_/B _49770_/Y sky130_fd_sc_hd__nand2_4
X_46982_ _46978_/Y _46940_/X _46981_/X _46982_/Y sky130_fd_sc_hd__a21oi_4
X_58968_ _84786_/Q _58956_/X _58960_/X _58967_/X _84786_/D sky130_fd_sc_hd__a2bb2oi_4
X_48721_ _48725_/A _48380_/X _48721_/Y sky130_fd_sc_hd__nand2_4
X_79541_ _84203_/Q _72465_/A _79543_/A sky130_fd_sc_hd__nor2_4
X_57919_ _57919_/A _57791_/X _57919_/Y sky130_fd_sc_hd__nor2_4
X_45933_ _45932_/Y _45933_/Y sky130_fd_sc_hd__inv_2
X_41056_ _41056_/A _41056_/Y sky130_fd_sc_hd__inv_2
X_76753_ _76753_/A _76753_/B _76753_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_8_148_0_CLK clkbuf_7_74_0_CLK/X clkbuf_9_296_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_73965_ _87586_/Q _73873_/B _73965_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_143_0_CLK clkbuf_9_71_0_CLK/X _81362_/CLK sky130_fd_sc_hd__clkbuf_1
X_58899_ _58828_/X _58896_/Y _58898_/Y _58874_/X _58832_/X _58899_/X
+ sky130_fd_sc_hd__o32a_4
X_75704_ _75696_/X _75704_/B _75705_/B sky130_fd_sc_hd__xor2_4
X_48652_ _48471_/A _48652_/X sky130_fd_sc_hd__buf_2
X_60930_ _60930_/A _60926_/X _60930_/C _60962_/A sky130_fd_sc_hd__nand3_4
X_72916_ _72916_/A _72916_/B _72917_/B sky130_fd_sc_hd__nand2_4
X_79472_ _79480_/A _79471_/Y _82845_/D sky130_fd_sc_hd__xor2_4
Xclkbuf_10_773_0_CLK clkbuf_9_386_0_CLK/X _82665_/CLK sky130_fd_sc_hd__clkbuf_1
X_45864_ _63342_/B _61685_/A sky130_fd_sc_hd__buf_2
X_76684_ _76692_/B _81350_/D _76688_/A sky130_fd_sc_hd__xnor2_4
X_73896_ _68732_/B _73872_/X _73894_/X _73895_/Y _73896_/X sky130_fd_sc_hd__a211o_4
X_47603_ _49504_/A _47792_/A sky130_fd_sc_hd__buf_2
X_78423_ _78423_/A _78421_/Y _78423_/C _78423_/Y sky130_fd_sc_hd__nand3_4
X_44815_ _44807_/X _43924_/X _41655_/X _86938_/Q _44808_/X _44816_/A
+ sky130_fd_sc_hd__o32ai_4
X_75635_ _75635_/A _75635_/B _75635_/X sky130_fd_sc_hd__xor2_4
X_60861_ _59540_/Y _61278_/B _60615_/A _61075_/C _60861_/X sky130_fd_sc_hd__and4_4
X_48583_ _48604_/A _48816_/B _48583_/Y sky130_fd_sc_hd__nand2_4
X_72847_ _72848_/B _72835_/X _72846_/X _72847_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_9_264_0_CLK clkbuf_8_132_0_CLK/X clkbuf_9_264_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_45795_ _84999_/Q _44935_/X _45389_/X _45795_/X sky130_fd_sc_hd__o21a_4
X_62600_ _62622_/A _62600_/B _62600_/C _62600_/D _62600_/Y sky130_fd_sc_hd__nand4_4
X_47534_ _47529_/Y _47509_/X _47533_/X _47534_/Y sky130_fd_sc_hd__a21oi_4
X_78354_ _78352_/X _78354_/B _78356_/B sky130_fd_sc_hd__nand2_4
X_44746_ _49210_/A _50731_/B _40749_/X _44745_/Y _44736_/X _86978_/D
+ sky130_fd_sc_hd__o32ai_4
X_63580_ _63576_/Y _63578_/X _63579_/Y _63580_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_158_0_CLK clkbuf_9_79_0_CLK/X _81680_/CLK sky130_fd_sc_hd__clkbuf_1
X_75566_ _75561_/Y _80801_/Q _75563_/B _75567_/B sky130_fd_sc_hd__nand3_4
X_41958_ _41937_/X _41956_/X _40712_/X _41957_/Y _41939_/X _88093_/D
+ sky130_fd_sc_hd__o32ai_4
X_60792_ _60792_/A _60761_/B _84566_/Q _60792_/Y sky130_fd_sc_hd__nor3_4
X_72778_ _44518_/Y _72775_/X _72777_/Y _72791_/C sky130_fd_sc_hd__a21o_4
X_77305_ _77305_/A _82132_/Q _77310_/A sky130_fd_sc_hd__nor2_4
Xclkbuf_10_788_0_CLK clkbuf_9_394_0_CLK/X _82740_/CLK sky130_fd_sc_hd__clkbuf_1
X_62531_ _61597_/A _62566_/B _62501_/X _62566_/D _62536_/B sky130_fd_sc_hd__nand4_4
X_74517_ _74516_/X _74517_/X sky130_fd_sc_hd__buf_2
X_40909_ _40908_/X _40909_/X sky130_fd_sc_hd__buf_2
X_47465_ _47465_/A _53063_/D sky130_fd_sc_hd__buf_2
X_71729_ _71729_/A _71256_/B _71724_/X _71729_/Y sky130_fd_sc_hd__nand3_4
X_78285_ _78280_/Y _78256_/B _78284_/X _78286_/B sky130_fd_sc_hd__o21ai_4
X_44677_ _44658_/X _44659_/X _40605_/X _87003_/Q _44660_/X _44677_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75497_ _75497_/A _75497_/Y sky130_fd_sc_hd__inv_2
X_41889_ _88112_/Q _41889_/Y sky130_fd_sc_hd__inv_2
X_49204_ _49052_/A _49204_/X sky130_fd_sc_hd__buf_2
X_46416_ _46416_/A _46417_/B sky130_fd_sc_hd__buf_2
X_65250_ _65118_/X _85544_/Q _65146_/X _65249_/X _65250_/X sky130_fd_sc_hd__a211o_4
X_77236_ _77236_/A _82083_/D _77239_/A sky130_fd_sc_hd__or2_4
X_43628_ _40656_/A _43609_/X _68672_/B _43611_/X _43628_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_9_279_0_CLK clkbuf_9_278_0_CLK/A clkbuf_9_279_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_62462_ _62623_/C _62462_/X sky130_fd_sc_hd__buf_2
X_74448_ _83064_/Q _74387_/X _74447_/Y _74448_/Y sky130_fd_sc_hd__o21ai_4
X_47396_ _47404_/A _53021_/B _47396_/Y sky130_fd_sc_hd__nand2_4
X_64201_ _64197_/X _64186_/X _64200_/Y _64201_/Y sky130_fd_sc_hd__a21oi_4
X_49135_ _49135_/A _49135_/X sky130_fd_sc_hd__buf_2
X_61413_ _61413_/A _61434_/A sky130_fd_sc_hd__buf_2
X_46347_ _46347_/A _46362_/A sky130_fd_sc_hd__buf_2
X_65181_ _65177_/X _65056_/B _65180_/X _65181_/Y sky130_fd_sc_hd__nand3_4
X_77167_ _77167_/A _77167_/B _77168_/B sky130_fd_sc_hd__xor2_4
X_43559_ _43558_/Y _87361_/D sky130_fd_sc_hd__inv_2
Xclkbuf_10_711_0_CLK clkbuf_9_355_0_CLK/X _88268_/CLK sky130_fd_sc_hd__clkbuf_1
X_62393_ _61479_/B _62390_/X _62363_/X _62323_/X _62392_/X _62393_/X
+ sky130_fd_sc_hd__a41o_4
X_74379_ _74408_/A _48391_/A _74379_/Y sky130_fd_sc_hd__nand2_4
X_64132_ _58976_/A _64102_/B _64132_/Y sky130_fd_sc_hd__nor2_4
X_76118_ _81724_/D _76126_/C _76118_/Y sky130_fd_sc_hd__nand2_4
X_49066_ _65087_/B _49052_/X _49065_/Y _49066_/Y sky130_fd_sc_hd__o21ai_4
X_61344_ _63380_/A _61368_/B _61368_/C _61368_/D _61344_/Y sky130_fd_sc_hd__nand4_4
X_46278_ _46273_/Y _46258_/X _46277_/Y _46278_/Y sky130_fd_sc_hd__a21boi_4
X_77098_ _77098_/A _82287_/D _77098_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_9_202_0_CLK clkbuf_9_203_0_CLK/A clkbuf_9_202_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_48017_ _66155_/B _47998_/X _48016_/Y _48017_/Y sky130_fd_sc_hd__o21ai_4
X_45229_ _45651_/A _45229_/X sky130_fd_sc_hd__buf_2
X_64063_ _83245_/Q _64158_/B _64158_/C _64045_/X _64064_/D sky130_fd_sc_hd__nand4_4
X_68940_ _68937_/X _68940_/B _68940_/Y sky130_fd_sc_hd__nand2_4
X_76049_ _81339_/Q _76041_/B _76049_/Y sky130_fd_sc_hd__nor2_4
X_61275_ _60440_/X _61272_/B _61264_/B _61202_/Y _61274_/Y _61275_/Y
+ sky130_fd_sc_hd__a41oi_4
X_63014_ _60595_/C _64225_/C _60399_/B _63014_/D _63014_/X sky130_fd_sc_hd__and4_4
X_60226_ _60255_/B _60331_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_726_0_CLK clkbuf_9_363_0_CLK/X _88301_/CLK sky130_fd_sc_hd__clkbuf_1
X_68871_ _69371_/A _68871_/X sky130_fd_sc_hd__buf_2
X_67822_ _67891_/A _86923_/Q _67822_/X sky130_fd_sc_hd__and2_4
X_79808_ _79804_/X _79820_/B _79829_/A sky130_fd_sc_hd__xor2_4
X_60157_ _60156_/Y _60251_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_217_0_CLK clkbuf_9_217_0_CLK/A clkbuf_9_217_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_49968_ _49915_/A _49973_/B sky130_fd_sc_hd__buf_2
X_48919_ _48913_/Y _48880_/X _48918_/X _48919_/Y sky130_fd_sc_hd__a21oi_4
X_79739_ _79732_/X _79739_/B _79739_/Y sky130_fd_sc_hd__nand2_4
X_67753_ _87458_/Q _67751_/X _67702_/X _67752_/X _67753_/X sky130_fd_sc_hd__a211o_4
X_64965_ _64960_/X _65111_/B _64964_/X _64965_/Y sky130_fd_sc_hd__nand3_4
X_60088_ _59852_/A _60103_/B sky130_fd_sc_hd__buf_2
X_49899_ _49904_/A _49893_/B _49893_/C _53113_/D _49899_/X sky130_fd_sc_hd__and4_4
X_66704_ _66728_/A _66704_/B _66704_/X sky130_fd_sc_hd__and2_4
Xclkbuf_4_2_0_CLK clkbuf_4_3_0_CLK/A clkbuf_4_2_1_CLK/A sky130_fd_sc_hd__clkbuf_1
X_51930_ _52322_/A _53199_/A sky130_fd_sc_hd__buf_2
X_63916_ _61468_/A _63853_/B _63947_/C _63866_/X _63916_/Y sky130_fd_sc_hd__nand4_4
X_82750_ _84161_/CLK _84134_/Q _79071_/A sky130_fd_sc_hd__dfxtp_4
X_67684_ _87153_/Q _67585_/X _67633_/X _67683_/X _67684_/X sky130_fd_sc_hd__a211o_4
X_64896_ _64696_/X _85526_/Q _64697_/X _64895_/X _64896_/X sky130_fd_sc_hd__a211o_4
X_81701_ _82053_/CLK _81701_/D _41266_/A sky130_fd_sc_hd__dfxtp_4
X_69423_ _69746_/A _69423_/X sky130_fd_sc_hd__buf_2
X_66635_ _87133_/Q _66633_/X _46212_/A _66634_/X _66635_/X sky130_fd_sc_hd__a211o_4
X_51861_ _51858_/Y _51850_/X _51860_/X _51861_/Y sky130_fd_sc_hd__a21oi_4
X_63847_ _63842_/X _63810_/X _63843_/Y _63844_/Y _63846_/X _63847_/X
+ sky130_fd_sc_hd__a41o_4
X_82681_ _81198_/CLK _82681_/D _78247_/A sky130_fd_sc_hd__dfxtp_4
X_53600_ _53598_/Y _53574_/X _53599_/Y _85605_/D sky130_fd_sc_hd__a21boi_4
X_84420_ _84420_/CLK _62303_/Y _62302_/C sky130_fd_sc_hd__dfxtp_4
X_50812_ _50812_/A _50751_/B _50751_/C _50812_/X sky130_fd_sc_hd__and3_4
X_81632_ _81632_/CLK _76628_/Y _81632_/Q sky130_fd_sc_hd__dfxtp_4
X_69354_ _69234_/A _69354_/B _69354_/X sky130_fd_sc_hd__and2_4
X_54580_ _54565_/A _54585_/B _54565_/C _54580_/D _54580_/X sky130_fd_sc_hd__and4_4
X_66566_ _69178_/A _69454_/A sky130_fd_sc_hd__buf_2
X_51792_ _85945_/Q _51789_/X _51791_/Y _51792_/Y sky130_fd_sc_hd__o21ai_4
X_63778_ _58225_/X _64189_/C _60908_/A _63731_/D _63779_/D sky130_fd_sc_hd__nand4_4
X_68305_ _67871_/X _67874_/X _68295_/X _68305_/Y sky130_fd_sc_hd__a21oi_4
X_53531_ _53468_/A _53531_/B _53531_/Y sky130_fd_sc_hd__nand2_4
X_65517_ _65790_/A _65517_/X sky130_fd_sc_hd__buf_2
X_84351_ _84350_/CLK _84351_/D _84351_/Q sky130_fd_sc_hd__dfxtp_4
X_50743_ _50596_/A _50771_/A sky130_fd_sc_hd__buf_2
X_62729_ _61399_/X _62694_/B _62694_/C _62729_/D _62729_/Y sky130_fd_sc_hd__nand4_4
X_81563_ _84064_/CLK _76879_/X _81563_/Q sky130_fd_sc_hd__dfxtp_4
X_69285_ _69190_/A _69286_/A sky130_fd_sc_hd__buf_2
X_66497_ _64636_/A _68823_/A sky130_fd_sc_hd__buf_2
X_83302_ _83303_/CLK _72015_/Y _83302_/Q sky130_fd_sc_hd__dfxtp_4
X_80514_ _84766_/Q _84158_/Q _80514_/Y sky130_fd_sc_hd__nand2_4
X_68236_ _68188_/X _67458_/Y _68228_/X _68235_/Y _68236_/X sky130_fd_sc_hd__a211o_4
X_56250_ _56250_/A _56253_/B _56250_/C _56250_/Y sky130_fd_sc_hd__nand3_4
X_87070_ _87070_/CLK _87070_/D _44518_/A sky130_fd_sc_hd__dfxtp_4
X_53462_ _53458_/A _50234_/B _53462_/Y sky130_fd_sc_hd__nand2_4
X_65448_ _65529_/A _65448_/X sky130_fd_sc_hd__buf_2
X_84282_ _84280_/CLK _84282_/D _63995_/C sky130_fd_sc_hd__dfxtp_4
X_50674_ _50657_/A _50674_/B _50674_/Y sky130_fd_sc_hd__nand2_4
X_81494_ _81333_/CLK _81494_/D _81494_/Q sky130_fd_sc_hd__dfxtp_4
X_55201_ _55201_/A _55196_/B _55201_/C _55201_/Y sky130_fd_sc_hd__nand3_4
X_86021_ _86121_/CLK _51381_/Y _65337_/B sky130_fd_sc_hd__dfxtp_4
X_52413_ _52400_/X _50716_/B _52413_/Y sky130_fd_sc_hd__nand2_4
X_83233_ _83227_/CLK _72566_/Y _79427_/B sky130_fd_sc_hd__dfxtp_4
X_56181_ _73163_/A _56181_/X sky130_fd_sc_hd__buf_2
X_80445_ _80467_/A _80445_/Y sky130_fd_sc_hd__inv_2
X_68167_ _67388_/X _68168_/A sky130_fd_sc_hd__buf_2
X_53393_ _53397_/A _53388_/B _53388_/C _52879_/D _53393_/X sky130_fd_sc_hd__and4_4
X_65379_ _65376_/X _65378_/X _64574_/X _65379_/X sky130_fd_sc_hd__a21o_4
X_55132_ _85035_/Q _55126_/X _55128_/X _55131_/X _55132_/X sky130_fd_sc_hd__a211o_4
X_67118_ _67095_/A _67118_/B _67118_/X sky130_fd_sc_hd__and2_4
X_52344_ _65032_/B _52324_/X _52343_/Y _52344_/Y sky130_fd_sc_hd__o21ai_4
X_83164_ _86570_/CLK _73123_/X _83164_/Q sky130_fd_sc_hd__dfxtp_4
X_80376_ _80370_/X _80372_/B _80376_/Y sky130_fd_sc_hd__nand2_4
X_68098_ _66632_/X _66635_/X _68062_/X _68098_/Y sky130_fd_sc_hd__a21oi_4
X_82115_ _82104_/CLK _82115_/D _82103_/D sky130_fd_sc_hd__dfxtp_4
X_55063_ _55054_/A _54898_/B _55063_/Y sky130_fd_sc_hd__nand2_4
X_59940_ _59938_/Y _59910_/X _62463_/A _59951_/B sky130_fd_sc_hd__nand3_4
X_67049_ _67023_/A _67049_/B _67049_/X sky130_fd_sc_hd__and2_4
X_52275_ _52295_/A _52275_/B _52275_/X sky130_fd_sc_hd__and2_4
X_87972_ _87150_/CLK _42221_/X _87972_/Q sky130_fd_sc_hd__dfxtp_4
X_83095_ _83095_/CLK _74333_/X _70318_/A sky130_fd_sc_hd__dfxtp_4
X_54014_ _85522_/Q _53940_/X _54013_/Y _54014_/Y sky130_fd_sc_hd__o21ai_4
X_51226_ _51223_/Y _51201_/X _51225_/X _86051_/D sky130_fd_sc_hd__a21oi_4
X_70060_ _68890_/X _68893_/X _70044_/X _70060_/Y sky130_fd_sc_hd__a21oi_4
X_86923_ _87144_/CLK _86923_/D _86923_/Q sky130_fd_sc_hd__dfxtp_4
X_82046_ _82047_/CLK _77994_/B _82046_/Q sky130_fd_sc_hd__dfxtp_4
X_59871_ _59651_/A _59797_/Y _59825_/X _59847_/Y _59870_/Y _59871_/Y
+ sky130_fd_sc_hd__a41oi_4
X_58822_ _58703_/X _85453_/Q _58821_/X _58822_/Y sky130_fd_sc_hd__o21ai_4
X_51157_ _51129_/A _51167_/A sky130_fd_sc_hd__buf_2
X_86854_ _84408_/CLK _86854_/D _63292_/B sky130_fd_sc_hd__dfxtp_4
X_50108_ _50103_/A _48992_/X _50108_/Y sky130_fd_sc_hd__nand2_4
X_85805_ _86040_/CLK _52525_/Y _65115_/B sky130_fd_sc_hd__dfxtp_4
X_58753_ _58748_/X _58750_/Y _58751_/Y _58650_/X _58752_/X _58753_/X
+ sky130_fd_sc_hd__o32a_4
X_51088_ _51141_/A _51110_/C sky130_fd_sc_hd__buf_2
X_55965_ _55965_/A _55965_/B _55966_/A sky130_fd_sc_hd__and2_4
X_86785_ _82317_/CLK _86785_/D _86785_/Q sky130_fd_sc_hd__dfxtp_4
X_83997_ _82642_/CLK _68266_/X _83997_/Q sky130_fd_sc_hd__dfxtp_4
X_57704_ _46213_/X _57692_/Y _57698_/Y _57700_/X _57703_/X _57704_/X
+ sky130_fd_sc_hd__o32a_4
X_42930_ _42962_/A _42930_/X sky130_fd_sc_hd__buf_2
X_50039_ _72461_/B _48170_/X _50038_/Y _50039_/Y sky130_fd_sc_hd__o21ai_4
X_54916_ _54932_/A _54910_/B _54932_/C _53223_/D _54916_/X sky130_fd_sc_hd__and4_4
X_73750_ _73750_/A _73624_/X _73750_/Y sky130_fd_sc_hd__nor2_4
X_85736_ _85738_/CLK _52888_/Y _85736_/Q sky130_fd_sc_hd__dfxtp_4
X_58684_ _58618_/X _86104_/Q _58683_/X _58684_/Y sky130_fd_sc_hd__o21ai_4
X_70962_ _70969_/A _70940_/B _70962_/C _70962_/Y sky130_fd_sc_hd__nand3_4
X_82948_ _82768_/CLK _82948_/D _82948_/Q sky130_fd_sc_hd__dfxtp_4
X_55896_ _55903_/A _55896_/B _55896_/X sky130_fd_sc_hd__and2_4
X_72701_ _83184_/Q _72699_/X _72700_/X _72701_/X sky130_fd_sc_hd__a21o_4
X_57635_ _71985_/A _57635_/X sky130_fd_sc_hd__buf_2
X_42861_ _41552_/X _42852_/X _66982_/B _42853_/X _42861_/X sky130_fd_sc_hd__a2bb2o_4
X_54847_ _54900_/A _54857_/B sky130_fd_sc_hd__buf_2
X_85667_ _85471_/CLK _85667_/D _85667_/Q sky130_fd_sc_hd__dfxtp_4
X_73681_ _68498_/B _73279_/X _73656_/X _73681_/X sky130_fd_sc_hd__o21a_4
X_70893_ _70867_/A _70890_/B _70890_/C _70899_/D _70893_/Y sky130_fd_sc_hd__nand4_4
X_82879_ _82879_/CLK _78296_/B _82879_/Q sky130_fd_sc_hd__dfxtp_4
X_44600_ _87040_/Q _44600_/Y sky130_fd_sc_hd__inv_2
X_87406_ _88171_/CLK _43470_/Y _87406_/Q sky130_fd_sc_hd__dfxtp_4
X_75420_ _75403_/Y _75406_/Y _75401_/Y _75420_/Y sky130_fd_sc_hd__o21ai_4
X_41812_ _48192_/A _48164_/A sky130_fd_sc_hd__buf_2
X_72632_ _45891_/X _72687_/A sky130_fd_sc_hd__buf_2
X_84618_ _84620_/CLK _84618_/D _60374_/C sky130_fd_sc_hd__dfxtp_4
X_45580_ _45574_/X _45577_/X _45579_/Y _86868_/D sky130_fd_sc_hd__a21oi_4
X_57566_ _84978_/Q _57562_/X _57565_/Y _57566_/Y sky130_fd_sc_hd__o21ai_4
X_42792_ _41371_/X _42787_/X _67727_/B _42788_/X _87715_/D sky130_fd_sc_hd__a2bb2o_4
X_88386_ _88386_/CLK _88386_/D _88386_/Q sky130_fd_sc_hd__dfxtp_4
X_54778_ _85379_/Q _54757_/X _54777_/Y _54778_/Y sky130_fd_sc_hd__o21ai_4
X_85598_ _85590_/CLK _53637_/Y _85598_/Q sky130_fd_sc_hd__dfxtp_4
X_59305_ _57696_/X _59306_/B sky130_fd_sc_hd__buf_2
X_44531_ _44531_/A _44531_/Y sky130_fd_sc_hd__inv_2
X_56517_ _56109_/X _56515_/X _56516_/Y _85166_/D sky130_fd_sc_hd__o21ai_4
X_75351_ _75351_/A _75351_/Y sky130_fd_sc_hd__inv_2
X_41743_ _40620_/X _41743_/B _41743_/X sky130_fd_sc_hd__or2_4
X_87337_ _87595_/CLK _87337_/D _73797_/A sky130_fd_sc_hd__dfxtp_4
X_53729_ _53729_/A _53729_/X sky130_fd_sc_hd__buf_2
X_72563_ _72525_/A _72563_/B _72563_/C _72570_/C sky130_fd_sc_hd__nand3_4
X_84549_ _84549_/CLK _84549_/D _60947_/C sky130_fd_sc_hd__dfxtp_4
X_57497_ _57497_/A _48178_/X _57497_/Y sky130_fd_sc_hd__nand2_4
X_74302_ _72704_/A _74302_/X sky130_fd_sc_hd__buf_2
X_47250_ _47245_/Y _47224_/X _47249_/X _86655_/D sky130_fd_sc_hd__a21oi_4
X_71514_ _71525_/A _71521_/A sky130_fd_sc_hd__buf_2
X_59236_ _59233_/Y _59235_/Y _59165_/X _59236_/X sky130_fd_sc_hd__a21o_4
X_78070_ _84575_/Q _78070_/B _78070_/X sky130_fd_sc_hd__xor2_4
X_44462_ _41147_/A _44453_/X _87097_/Q _44454_/X _44462_/X sky130_fd_sc_hd__a2bb2o_4
X_56448_ _44207_/A _56448_/X sky130_fd_sc_hd__buf_2
X_75282_ _75280_/X _75263_/X _75281_/Y _75282_/Y sky130_fd_sc_hd__a21oi_4
X_87268_ _87525_/CLK _87268_/D _87268_/Q sky130_fd_sc_hd__dfxtp_4
X_41674_ _41674_/A _41653_/X _41674_/X sky130_fd_sc_hd__or2_4
X_72494_ _63611_/A _72488_/B _72494_/Y sky130_fd_sc_hd__nand2_4
X_46201_ _44228_/X _58425_/A sky130_fd_sc_hd__buf_2
XPHY_130 sky130_fd_sc_hd__decap_3
X_77021_ _77021_/A _77020_/Y _77022_/B sky130_fd_sc_hd__xor2_4
X_43413_ _43397_/A _43413_/X sky130_fd_sc_hd__buf_2
X_74233_ _45931_/X _86212_/Q _72985_/X _74232_/X _74233_/X sky130_fd_sc_hd__a211o_4
X_86219_ _85599_/CLK _86219_/D _86219_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_141 sky130_fd_sc_hd__decap_3
X_40625_ _40621_/X _82874_/Q _40624_/X _40625_/Y sky130_fd_sc_hd__o21ai_4
X_47181_ _47152_/X _47181_/B _47143_/C _52900_/D _47181_/X sky130_fd_sc_hd__and4_4
X_59167_ _59154_/A _59167_/B _59167_/Y sky130_fd_sc_hd__nor2_4
X_71445_ _71444_/Y _71445_/X sky130_fd_sc_hd__buf_2
X_44393_ _41479_/X _44377_/X _87131_/Q _44379_/X _44393_/X sky130_fd_sc_hd__a2bb2o_4
X_56379_ _56458_/A _56363_/B _56379_/C _56379_/Y sky130_fd_sc_hd__nand3_4
XPHY_152 sky130_fd_sc_hd__decap_3
X_87199_ _87720_/CLK _43920_/X _67810_/B sky130_fd_sc_hd__dfxtp_4
XPHY_163 sky130_fd_sc_hd__decap_3
XPHY_174 sky130_fd_sc_hd__decap_3
X_46132_ _46111_/B _74846_/B _46207_/B sky130_fd_sc_hd__nor2_4
X_58118_ _57989_/X _58116_/Y _58117_/Y _58007_/X _57993_/X _58118_/X
+ sky130_fd_sc_hd__o32a_4
XPHY_185 sky130_fd_sc_hd__decap_3
X_43344_ _43316_/X _43319_/X _41321_/X _87468_/Q _43330_/X _43344_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74164_ _74164_/A _73152_/X _74164_/Y sky130_fd_sc_hd__nor2_4
XPHY_196 sky130_fd_sc_hd__decap_3
X_40556_ _40556_/A _40556_/X sky130_fd_sc_hd__buf_2
X_71376_ _71458_/C _71377_/C sky130_fd_sc_hd__buf_2
X_59098_ _59073_/X _85753_/Q _59037_/X _59098_/X sky130_fd_sc_hd__o21a_4
X_73115_ _72988_/X _85588_/Q _73092_/A _73114_/X _73115_/X sky130_fd_sc_hd__a211o_4
X_46063_ _41559_/Y _46061_/X _86787_/Q _46062_/X _46063_/X sky130_fd_sc_hd__a2bb2o_4
X_58049_ _57997_/X _85481_/Q _57923_/X _58049_/X sky130_fd_sc_hd__o21a_4
X_70327_ _70325_/Y _70157_/A _70326_/Y _83796_/D sky130_fd_sc_hd__o21ai_4
X_43275_ _43274_/Y _43275_/Y sky130_fd_sc_hd__inv_2
X_74095_ _74095_/A _74095_/B _74095_/Y sky130_fd_sc_hd__nor2_4
X_78972_ _78959_/Y _78960_/Y _78971_/X _78972_/Y sky130_fd_sc_hd__a21oi_4
X_40487_ _40362_/X _44382_/A sky130_fd_sc_hd__buf_2
X_45014_ _56211_/C _44998_/X _45013_/X _45014_/Y sky130_fd_sc_hd__o21ai_4
X_42226_ _42199_/X _42226_/X sky130_fd_sc_hd__buf_2
X_61060_ _84524_/Q _60349_/X _61059_/X _84524_/D sky130_fd_sc_hd__o21a_4
X_73046_ _56181_/X _83071_/Q _72880_/X _73045_/X _73046_/X sky130_fd_sc_hd__a211o_4
X_77923_ _77923_/A _77922_/Y _82039_/D sky130_fd_sc_hd__xnor2_4
X_70258_ _70260_/A _70260_/B _83180_/Q _70260_/D _70258_/X sky130_fd_sc_hd__and4_4
X_60011_ _62478_/A _60011_/X sky130_fd_sc_hd__buf_2
X_49822_ _49794_/X _49830_/C sky130_fd_sc_hd__buf_2
X_42157_ _41179_/X _42148_/X _88006_/Q _42150_/X _88006_/D sky130_fd_sc_hd__a2bb2o_4
X_77854_ _77842_/A _77849_/A _77854_/X sky130_fd_sc_hd__and2_4
X_70189_ _70169_/X _83844_/Q _70188_/X _83844_/D sky130_fd_sc_hd__a21o_4
X_41108_ _41107_/Y _41108_/X sky130_fd_sc_hd__buf_2
X_76805_ _76805_/A _76804_/Y _76808_/A sky130_fd_sc_hd__xor2_4
X_49753_ _49757_/A _52969_/B _49753_/Y sky130_fd_sc_hd__nand2_4
X_46965_ _46981_/A _46944_/B _46981_/C _52775_/D _46965_/X sky130_fd_sc_hd__and4_4
X_42088_ _42083_/X _42077_/X _40994_/X _88040_/Q _42078_/X _42088_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77785_ _82152_/Q _77785_/B _82120_/D sky130_fd_sc_hd__xor2_4
X_74997_ _74994_/X _74996_/Y _74998_/B sky130_fd_sc_hd__xnor2_4
X_48704_ _48704_/A _48704_/Y sky130_fd_sc_hd__inv_2
X_79524_ _79524_/A _79163_/Y _79525_/B sky130_fd_sc_hd__nand2_4
X_41039_ _41039_/A _41039_/Y sky130_fd_sc_hd__inv_2
X_45916_ _45915_/X _69626_/A sky130_fd_sc_hd__buf_2
X_64750_ _64657_/X _86748_/Q _64733_/X _64749_/X _64750_/X sky130_fd_sc_hd__a211o_4
X_76736_ _76736_/A _76735_/Y _76744_/A sky130_fd_sc_hd__xor2_4
X_61962_ _59721_/X _61962_/X sky130_fd_sc_hd__buf_2
X_49684_ _49657_/A _49685_/C sky130_fd_sc_hd__buf_2
X_73948_ _73948_/A _73948_/X sky130_fd_sc_hd__buf_2
X_46896_ _46868_/A _46896_/B _46868_/C _52735_/D _46896_/X sky130_fd_sc_hd__and4_4
X_63701_ _63701_/A _63701_/B _80293_/A _63701_/Y sky130_fd_sc_hd__nor3_4
X_60913_ _60908_/X _60911_/X _60994_/A _60913_/Y sky130_fd_sc_hd__o21ai_4
X_48635_ _48635_/A _48657_/B sky130_fd_sc_hd__buf_2
X_79455_ _58623_/A _79455_/B _79455_/X sky130_fd_sc_hd__xor2_4
X_45847_ _45847_/A _74700_/B sky130_fd_sc_hd__inv_2
X_64681_ _64678_/X _85566_/Q _64679_/X _64680_/X _64681_/X sky130_fd_sc_hd__a211o_4
X_76667_ _76967_/B _76667_/Y sky130_fd_sc_hd__inv_2
X_61893_ _61891_/X _61846_/B _61878_/C _61910_/D _61893_/Y sky130_fd_sc_hd__nand4_4
X_73879_ _73850_/X _86228_/Q _73804_/X _73878_/X _73879_/X sky130_fd_sc_hd__a211o_4
X_66420_ _66433_/A _66419_/X _66420_/C _66420_/X sky130_fd_sc_hd__and3_4
X_78406_ _78402_/Y _78404_/Y _78405_/Y _78411_/A sky130_fd_sc_hd__o21ai_4
X_63632_ _63632_/A _63661_/C sky130_fd_sc_hd__buf_2
X_75618_ _81112_/Q _80824_/Q _80776_/D sky130_fd_sc_hd__xor2_4
X_48566_ _48563_/X _82351_/Q _48565_/Y _48567_/A sky130_fd_sc_hd__o21ai_4
X_60844_ _60843_/X _60844_/X sky130_fd_sc_hd__buf_2
X_79386_ _79384_/X _79391_/B _79386_/Y sky130_fd_sc_hd__xnor2_4
X_45778_ _45748_/X _63280_/B _45765_/X _45778_/Y sky130_fd_sc_hd__o21ai_4
X_76598_ _76597_/B _76596_/Y _76593_/Y _76598_/Y sky130_fd_sc_hd__o21ai_4
X_47517_ _47517_/A _53095_/B _47517_/Y sky130_fd_sc_hd__nand2_4
X_66351_ _58697_/A _85602_/Q _66349_/X _66350_/X _66351_/X sky130_fd_sc_hd__a211o_4
X_78337_ _78335_/Y _78334_/Y _78337_/C _78338_/A sky130_fd_sc_hd__nand3_4
X_44729_ _44712_/X _44713_/X _40724_/X _74119_/A _44714_/X _44730_/A
+ sky130_fd_sc_hd__o32ai_4
X_63563_ _61521_/B _63548_/X _63561_/X _63562_/Y _63563_/X sky130_fd_sc_hd__a211o_4
X_75549_ _75546_/Y _75562_/A _75551_/B sky130_fd_sc_hd__nand2_4
X_48497_ _48471_/X _47963_/A _48496_/Y _48498_/A sky130_fd_sc_hd__o21ai_4
X_60775_ _60267_/A _70021_/C sky130_fd_sc_hd__buf_2
X_65302_ _57694_/X _86022_/Q _65302_/X sky130_fd_sc_hd__and2_4
X_62514_ _62512_/Y _62467_/X _62513_/Y _84405_/D sky130_fd_sc_hd__a21oi_4
X_69070_ _41973_/A _68958_/X _68745_/X _69069_/Y _69070_/X sky130_fd_sc_hd__a211o_4
X_47448_ _47437_/X _47415_/X _47466_/C _53052_/D _47448_/X sky130_fd_sc_hd__and4_4
X_66282_ _65516_/A _66282_/X sky130_fd_sc_hd__buf_2
X_78268_ _78264_/Y _78256_/B _78282_/A _78268_/Y sky130_fd_sc_hd__o21ai_4
X_63494_ _63492_/Y _63455_/X _63493_/Y _84319_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_650_0_CLK clkbuf_9_325_0_CLK/X _88232_/CLK sky130_fd_sc_hd__clkbuf_1
X_68021_ _87382_/Q _67953_/X _67954_/X _68020_/X _68021_/X sky130_fd_sc_hd__a211o_4
X_65233_ _65233_/A _65233_/B _65233_/Y sky130_fd_sc_hd__nand2_4
X_77219_ _77219_/A _77219_/B _77220_/B sky130_fd_sc_hd__xor2_4
X_62445_ _62198_/Y _62493_/A sky130_fd_sc_hd__buf_2
X_47379_ _47379_/A _53015_/D sky130_fd_sc_hd__buf_2
X_78199_ _78199_/A _78199_/B _78199_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_141_0_CLK clkbuf_8_70_0_CLK/X clkbuf_9_141_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_49118_ _86442_/Q _49104_/X _49117_/Y _49118_/Y sky130_fd_sc_hd__o21ai_4
X_80230_ _80216_/A _80215_/X _80229_/Y _80230_/Y sky130_fd_sc_hd__a21boi_4
X_65164_ _65164_/A _65164_/B _65164_/X sky130_fd_sc_hd__and2_4
X_50390_ _86210_/Q _50387_/X _50389_/Y _50390_/Y sky130_fd_sc_hd__o21ai_4
X_62376_ _62522_/B _62420_/C sky130_fd_sc_hd__buf_2
X_64115_ _64077_/Y _64110_/Y _64111_/X _64113_/X _64114_/X _64115_/Y
+ sky130_fd_sc_hd__o41ai_4
X_49049_ _49049_/A _48959_/B _50645_/B sky130_fd_sc_hd__nor2_4
X_61327_ _59829_/X _61325_/Y _61326_/X _84489_/D sky130_fd_sc_hd__o21a_4
X_80161_ _80139_/Y _80157_/X _80160_/Y _80162_/B sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_665_0_CLK clkbuf_9_332_0_CLK/X _87684_/CLK sky130_fd_sc_hd__clkbuf_1
X_65095_ _64944_/X _86158_/Q _65022_/X _65094_/X _65095_/X sky130_fd_sc_hd__a211o_4
X_69972_ _69853_/A _69972_/B _69972_/X sky130_fd_sc_hd__and2_4
X_52060_ _52014_/X _50358_/B _52060_/Y sky130_fd_sc_hd__nand2_4
X_68923_ _68919_/X _68921_/X _68922_/X _68923_/X sky130_fd_sc_hd__a21o_4
X_64046_ _62022_/A _64046_/B _64046_/C _64045_/X _64047_/D sky130_fd_sc_hd__nand4_4
X_61258_ _61258_/A _61258_/Y sky130_fd_sc_hd__inv_2
X_80092_ _80092_/A _80091_/X _80105_/B sky130_fd_sc_hd__xnor2_4
Xclkbuf_9_156_0_CLK clkbuf_8_78_0_CLK/X clkbuf_9_156_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_51011_ _51039_/A _51011_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_83_0_CLK clkbuf_9_83_0_CLK/A clkbuf_9_83_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_60209_ _62644_/A _60211_/A sky130_fd_sc_hd__buf_2
X_83920_ _81507_/CLK _83920_/D _81384_/D sky130_fd_sc_hd__dfxtp_4
X_68854_ _87084_/Q _68832_/X _68762_/X _68853_/X _68854_/X sky130_fd_sc_hd__a211o_4
X_61189_ _84511_/Q _60719_/X _59753_/Y _61188_/Y _61189_/X sky130_fd_sc_hd__o22a_4
X_67805_ _81486_/D _67688_/X _67804_/X _84054_/D sky130_fd_sc_hd__a21bo_4
X_83851_ _86988_/CLK _70094_/X _82531_/D sky130_fd_sc_hd__dfxtp_4
X_68785_ _68785_/A _88355_/Q _68785_/X sky130_fd_sc_hd__and2_4
X_65997_ _65980_/X _65997_/B _65997_/X sky130_fd_sc_hd__and2_4
X_82802_ _84177_/CLK _82834_/Q _82802_/Q sky130_fd_sc_hd__dfxtp_4
X_55750_ _55252_/A _85160_/Q _55750_/X sky130_fd_sc_hd__and2_4
X_67736_ _84057_/Q _67688_/X _67735_/X _67736_/X sky130_fd_sc_hd__a21bo_4
X_86570_ _86570_/CLK _86570_/D _66238_/B sky130_fd_sc_hd__dfxtp_4
X_64948_ _64948_/A _64948_/B _64948_/X sky130_fd_sc_hd__and2_4
X_52962_ _53069_/A _52982_/B sky130_fd_sc_hd__buf_2
X_83782_ _83783_/CLK _70385_/Y _83782_/Q sky130_fd_sc_hd__dfxtp_4
X_80994_ _81985_/CLK _65421_/C _75571_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_98_0_CLK clkbuf_9_99_0_CLK/A clkbuf_9_98_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_54701_ _54699_/X _54707_/B _54721_/C _47369_/A _54701_/X sky130_fd_sc_hd__and4_4
X_85521_ _85815_/CLK _85521_/D _85521_/Q sky130_fd_sc_hd__dfxtp_4
X_51913_ _51804_/A _51914_/A sky130_fd_sc_hd__buf_2
X_82733_ _82692_/CLK _66469_/C _82733_/Q sky130_fd_sc_hd__dfxtp_4
X_55681_ _55681_/A _55680_/Y _55681_/X sky130_fd_sc_hd__xor2_4
X_67667_ _67615_/X _67667_/B _67667_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_603_0_CLK clkbuf_9_301_0_CLK/X _81989_/CLK sky130_fd_sc_hd__clkbuf_1
X_52893_ _52620_/A _52893_/X sky130_fd_sc_hd__buf_2
X_64879_ _64809_/X _86743_/Q _64864_/X _64878_/X _64879_/X sky130_fd_sc_hd__a211o_4
X_57420_ _57275_/X _56727_/X _57419_/X _57420_/X sky130_fd_sc_hd__o21a_4
X_69406_ _68852_/X _68854_/X _69295_/X _69406_/Y sky130_fd_sc_hd__a21oi_4
X_88240_ _87408_/CLK _88240_/D _67411_/B sky130_fd_sc_hd__dfxtp_4
X_54632_ _54636_/A _54106_/B _54632_/Y sky130_fd_sc_hd__nand2_4
X_66618_ _68999_/A _66618_/B _66618_/X sky130_fd_sc_hd__and2_4
X_85452_ _85773_/CLK _85452_/D _85452_/Q sky130_fd_sc_hd__dfxtp_4
X_51844_ _51851_/A _51851_/B _51851_/C _46783_/X _51844_/X sky130_fd_sc_hd__and4_4
X_82664_ _82879_/CLK _82664_/D _82664_/Q sky130_fd_sc_hd__dfxtp_4
X_67598_ _67593_/X _67597_/X _67502_/X _67602_/A sky130_fd_sc_hd__a21o_4
Xclkbuf_9_21_0_CLK clkbuf_8_10_0_CLK/X clkbuf_9_21_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_84403_ _84403_/CLK _84403_/D _62541_/C sky130_fd_sc_hd__dfxtp_4
X_81615_ _81615_/CLK _81615_/D _81807_/D sky130_fd_sc_hd__dfxtp_4
X_57351_ _57351_/A _57351_/B _57351_/Y sky130_fd_sc_hd__nand2_4
X_69337_ _69334_/X _69336_/X _69142_/X _69337_/Y sky130_fd_sc_hd__a21oi_4
X_88171_ _88171_/CLK _41678_/Y _88171_/Q sky130_fd_sc_hd__dfxtp_4
X_54563_ _54481_/A _54565_/A sky130_fd_sc_hd__buf_2
X_66549_ _68342_/A _69457_/A sky130_fd_sc_hd__buf_2
X_85383_ _85379_/CLK _85383_/D _85383_/Q sky130_fd_sc_hd__dfxtp_4
X_51775_ _85948_/Q _51763_/X _51774_/Y _51775_/Y sky130_fd_sc_hd__o21ai_4
X_82595_ _82595_/CLK _78821_/B _82595_/Q sky130_fd_sc_hd__dfxtp_4
X_56302_ _56031_/X _56290_/X _56301_/Y _56302_/Y sky130_fd_sc_hd__o21ai_4
X_87122_ _88201_/CLK _87122_/D _87122_/Q sky130_fd_sc_hd__dfxtp_4
X_53514_ _53509_/A _53514_/B _53514_/Y sky130_fd_sc_hd__nand2_4
X_84334_ _82272_/CLK _63319_/Y _79211_/B sky130_fd_sc_hd__dfxtp_4
X_50726_ _50722_/Y _50676_/X _50725_/X _50726_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_618_0_CLK clkbuf_9_309_0_CLK/X _81182_/CLK sky130_fd_sc_hd__clkbuf_1
X_57282_ _57281_/X _57273_/Y _56704_/X _57282_/Y sky130_fd_sc_hd__a21oi_4
X_81546_ _81344_/CLK _76726_/X _81546_/Q sky130_fd_sc_hd__dfxtp_4
X_69268_ _68606_/X _68608_/X _69212_/X _69268_/Y sky130_fd_sc_hd__a21oi_4
X_54494_ _54483_/A _54503_/B _54483_/C _54494_/D _54494_/X sky130_fd_sc_hd__and4_4
X_59021_ _58961_/X _85663_/Q _59010_/X _59021_/X sky130_fd_sc_hd__o21a_4
X_56233_ _56233_/A _56243_/B _56233_/C _56233_/Y sky130_fd_sc_hd__nand3_4
X_68219_ _82657_/D _68200_/X _68218_/X _68219_/X sky130_fd_sc_hd__a21bo_4
X_87053_ _88062_/CLK _44564_/Y _87053_/Q sky130_fd_sc_hd__dfxtp_4
X_53445_ _85633_/Q _43021_/X _53444_/X _53445_/Y sky130_fd_sc_hd__o21ai_4
X_84265_ _84623_/CLK _64216_/Y _79883_/B sky130_fd_sc_hd__dfxtp_4
X_50657_ _50657_/A _50144_/B _50657_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_109_0_CLK clkbuf_8_54_0_CLK/X clkbuf_9_109_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_81477_ _88121_/CLK _81477_/D _81477_/Q sky130_fd_sc_hd__dfxtp_4
X_69199_ _68484_/X _68486_/X _69061_/X _69199_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_36_0_CLK clkbuf_9_37_0_CLK/A clkbuf_9_36_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_86004_ _85718_/CLK _51474_/Y _86004_/Q sky130_fd_sc_hd__dfxtp_4
X_40410_ _40409_/X _40410_/X sky130_fd_sc_hd__buf_2
X_71230_ _71232_/A _71230_/B _71232_/C _71230_/Y sky130_fd_sc_hd__nand3_4
X_83216_ _83216_/CLK _72613_/X _79245_/B sky130_fd_sc_hd__dfxtp_4
X_80428_ _80425_/Y _80408_/Y _80427_/X _80429_/B sky130_fd_sc_hd__o21ai_4
X_56164_ _56164_/A _56164_/X sky130_fd_sc_hd__buf_2
X_41390_ _41389_/Y _88224_/D sky130_fd_sc_hd__inv_2
X_53376_ _53371_/A _53388_/B _53371_/C _52861_/D _53376_/X sky130_fd_sc_hd__and4_4
X_84196_ _85315_/CLK _84196_/D _84196_/Q sky130_fd_sc_hd__dfxtp_4
X_50588_ _52291_/A _50560_/X _50568_/C _50588_/X sky130_fd_sc_hd__and3_4
X_55115_ _85315_/Q _55098_/X _55114_/Y _55115_/Y sky130_fd_sc_hd__o21ai_4
X_40341_ _47363_/A _74492_/A sky130_fd_sc_hd__buf_2
X_52327_ _85845_/Q _52324_/X _52326_/Y _52327_/Y sky130_fd_sc_hd__o21ai_4
X_71161_ _48435_/B _71138_/A _71160_/Y _83586_/D sky130_fd_sc_hd__o21ai_4
X_83147_ _86218_/CLK _83147_/D _83147_/Q sky130_fd_sc_hd__dfxtp_4
X_56095_ _45765_/A _56115_/B sky130_fd_sc_hd__buf_2
X_80359_ _80360_/B _80350_/B _80358_/Y _80361_/A sky130_fd_sc_hd__a21o_4
X_70112_ _70108_/Y _70109_/Y _70112_/C _70111_/Y _70118_/C sky130_fd_sc_hd__nand4_4
X_55046_ _55072_/A _55046_/X sky130_fd_sc_hd__buf_2
X_59923_ _59909_/Y _59923_/Y sky130_fd_sc_hd__inv_2
X_43060_ _43024_/A _43121_/A sky130_fd_sc_hd__buf_2
X_71092_ _52338_/B _71070_/A _71091_/Y _71092_/Y sky130_fd_sc_hd__o21ai_4
X_52258_ _52256_/Y _52117_/X _52257_/Y _52258_/Y sky130_fd_sc_hd__a21boi_4
X_83078_ _86523_/CLK _74382_/Y _83078_/Q sky130_fd_sc_hd__dfxtp_4
X_87955_ _87126_/CLK _87955_/D _87955_/Q sky130_fd_sc_hd__dfxtp_4
X_42011_ _88072_/Q _42011_/Y sky130_fd_sc_hd__inv_2
X_51209_ _51128_/A _51209_/X sky130_fd_sc_hd__buf_2
X_86906_ _84420_/CLK _44997_/Y _64275_/B sky130_fd_sc_hd__dfxtp_4
X_74920_ _74920_/A _74920_/B _81189_/D sky130_fd_sc_hd__xor2_4
X_82029_ _82131_/CLK _77831_/B _82029_/Q sky130_fd_sc_hd__dfxtp_4
X_70043_ _82545_/D _70029_/X _70042_/X _70043_/X sky130_fd_sc_hd__a21bo_4
X_59854_ _59727_/X _59850_/Y _59762_/Y _59733_/Y _59853_/Y _59854_/Y
+ sky130_fd_sc_hd__a41oi_4
X_52189_ _52187_/Y _52117_/X _52188_/Y _85872_/D sky130_fd_sc_hd__a21boi_4
X_87886_ _87625_/CLK _87886_/D _87886_/Q sky130_fd_sc_hd__dfxtp_4
X_58805_ _58805_/A _58897_/A sky130_fd_sc_hd__buf_2
X_74851_ _81123_/D _80835_/Q _74852_/B sky130_fd_sc_hd__xor2_4
X_86837_ _87995_/CLK _45966_/X _66602_/B sky130_fd_sc_hd__dfxtp_4
X_59785_ _59737_/A _59848_/B _80497_/A _59785_/Y sky130_fd_sc_hd__nor3_4
X_56997_ _44184_/X _56997_/X sky130_fd_sc_hd__buf_2
X_73802_ _88361_/Q _73801_/X _73704_/X _73802_/Y sky130_fd_sc_hd__o21ai_4
X_46750_ _58751_/A _46719_/X _46749_/Y _46750_/Y sky130_fd_sc_hd__o21ai_4
X_58736_ _58732_/Y _58734_/Y _58735_/X _58736_/X sky130_fd_sc_hd__a21o_4
X_77570_ _77570_/A _77567_/Y _77570_/C _77575_/A sky130_fd_sc_hd__or3_4
X_43962_ _43957_/A _87178_/Q _43962_/X sky130_fd_sc_hd__and2_4
X_55948_ _56203_/C _55605_/X _44090_/B _55947_/X _55948_/X sky130_fd_sc_hd__a211o_4
X_86768_ _86218_/CLK _46172_/Y _72838_/A sky130_fd_sc_hd__dfxtp_4
X_74782_ _74723_/X _74782_/B _74745_/D _74782_/Y sky130_fd_sc_hd__nand3_4
X_71994_ _71993_/X _71994_/B _71994_/Y sky130_fd_sc_hd__nand2_4
X_45701_ _45694_/X _45698_/Y _45700_/Y _45701_/Y sky130_fd_sc_hd__a21oi_4
X_76521_ _76522_/A _76522_/B _76521_/Y sky130_fd_sc_hd__nor2_4
X_42913_ _41701_/X _42900_/X _67652_/B _42901_/X _42913_/X sky130_fd_sc_hd__a2bb2o_4
X_73733_ _73733_/A _66006_/B _73733_/X sky130_fd_sc_hd__and2_4
X_85719_ _85718_/CLK _52983_/Y _85719_/Q sky130_fd_sc_hd__dfxtp_4
X_46681_ _46680_/Y _50919_/D sky130_fd_sc_hd__buf_2
X_58667_ _58796_/A _58667_/X sky130_fd_sc_hd__buf_2
X_70945_ _70947_/A _70945_/B _70947_/C _70945_/Y sky130_fd_sc_hd__nand3_4
X_43893_ _43892_/Y _87212_/D sky130_fd_sc_hd__inv_2
X_55879_ _44081_/X _55879_/B _55879_/X sky130_fd_sc_hd__and2_4
X_86699_ _86701_/CLK _86699_/D _58853_/A sky130_fd_sc_hd__dfxtp_4
X_48420_ _48897_/A _48613_/A sky130_fd_sc_hd__buf_2
X_79240_ _79248_/C _79240_/B _79235_/B _79240_/Y sky130_fd_sc_hd__nand3_4
X_45632_ _45734_/A _45632_/X sky130_fd_sc_hd__buf_2
X_57618_ _84968_/Q _57615_/X _57617_/Y _57618_/Y sky130_fd_sc_hd__o21ai_4
X_76452_ _76451_/Y _76455_/B sky130_fd_sc_hd__inv_2
X_42844_ _42816_/X _42817_/X _41515_/X _66828_/B _42836_/X _42845_/A
+ sky130_fd_sc_hd__o32ai_4
X_73664_ _73660_/X _73663_/X _73612_/X _73668_/A sky130_fd_sc_hd__a21o_4
X_70876_ _70903_/A _70869_/B _70869_/C _70875_/X _70876_/Y sky130_fd_sc_hd__nand4_4
X_58598_ _84815_/Q _58095_/X _58590_/X _58597_/X _84815_/D sky130_fd_sc_hd__a2bb2oi_4
X_75403_ _75403_/A _75403_/Y sky130_fd_sc_hd__inv_2
X_48351_ _48163_/X _48392_/A sky130_fd_sc_hd__buf_2
X_72615_ _72581_/A _72604_/B _79231_/B _72615_/Y sky130_fd_sc_hd__nor3_4
X_79171_ _79171_/A _79171_/B _79171_/C _79171_/Y sky130_fd_sc_hd__nand3_4
X_45563_ _63124_/B _61451_/A sky130_fd_sc_hd__buf_2
X_57549_ _57547_/Y _57543_/X _57548_/Y _84981_/D sky130_fd_sc_hd__a21boi_4
X_76383_ _76347_/A _76348_/X _76371_/X _76383_/X sky130_fd_sc_hd__a21bo_4
X_88369_ _86982_/CLK _40583_/Y _88369_/Q sky130_fd_sc_hd__dfxtp_4
X_42775_ _42723_/A _42775_/X sky130_fd_sc_hd__buf_2
X_73595_ _73595_/A _73228_/B _73595_/Y sky130_fd_sc_hd__nor2_4
X_47302_ _47302_/A _52971_/D sky130_fd_sc_hd__buf_2
X_78122_ _78121_/X _78123_/B sky130_fd_sc_hd__buf_2
X_44514_ _44514_/A _44514_/Y sky130_fd_sc_hd__inv_2
X_75334_ _75330_/Y _75331_/Y _75333_/Y _75334_/X sky130_fd_sc_hd__or3_4
X_41726_ _41717_/X _81743_/Q _41725_/X _41727_/A sky130_fd_sc_hd__o21ai_4
X_48282_ _48275_/X _50326_/B _48282_/Y sky130_fd_sc_hd__nand2_4
X_60560_ _60612_/A _60526_/B _79140_/A _60560_/Y sky130_fd_sc_hd__nor3_4
X_72546_ _72528_/Y _72575_/A _72555_/B _65307_/A _64789_/A _72546_/Y
+ sky130_fd_sc_hd__a32oi_4
X_45494_ _45494_/A _45495_/A sky130_fd_sc_hd__inv_2
X_47233_ _57722_/A _47192_/X _47232_/Y _47233_/Y sky130_fd_sc_hd__o21ai_4
X_59219_ _58846_/A _59219_/X sky130_fd_sc_hd__buf_2
X_78053_ _60822_/C _78053_/B _78053_/X sky130_fd_sc_hd__xor2_4
X_44445_ _41626_/X _44431_/X _87104_/Q _44432_/X _87104_/D sky130_fd_sc_hd__a2bb2o_4
X_75265_ _75279_/B _75265_/B _81039_/D sky130_fd_sc_hd__xor2_4
X_41657_ _41611_/X _41613_/X _41656_/X _67468_/B _41608_/X _41658_/A
+ sky130_fd_sc_hd__o32ai_4
X_72477_ _72413_/X _72475_/Y _72476_/Y _57793_/X _72417_/X _72477_/X
+ sky130_fd_sc_hd__o32a_4
X_60491_ _60476_/D _63004_/C _60341_/A _60491_/X sky130_fd_sc_hd__o21a_4
X_77004_ _81986_/Q _82274_/D _77004_/Y sky130_fd_sc_hd__nand2_4
X_74216_ _74213_/X _74215_/X _56547_/X _74216_/X sky130_fd_sc_hd__a21o_4
X_62230_ _62522_/B _62233_/C sky130_fd_sc_hd__buf_2
X_40608_ _47943_/A _82876_/Q _40608_/X sky130_fd_sc_hd__or2_4
X_47164_ _47160_/Y _47128_/X _47163_/X _47164_/Y sky130_fd_sc_hd__a21oi_4
X_71428_ _71420_/X _83503_/Q _71427_/X _83503_/D sky130_fd_sc_hd__a21o_4
X_44376_ _41778_/X _44364_/X _87139_/Q _44365_/X _87139_/D sky130_fd_sc_hd__a2bb2o_4
X_75196_ _75192_/Y _75135_/Y _75195_/X _75196_/Y sky130_fd_sc_hd__o21ai_4
X_41588_ _41411_/X _41588_/X sky130_fd_sc_hd__buf_2
X_46115_ _46115_/A _46094_/A _46204_/C sky130_fd_sc_hd__nor2_4
X_43327_ _41268_/X _43325_/X _87479_/Q _43326_/X _87479_/D sky130_fd_sc_hd__a2bb2o_4
X_62161_ _61673_/B _62161_/B _62187_/C _61706_/X _62161_/Y sky130_fd_sc_hd__nand4_4
X_74147_ _74144_/X _74146_/X _72737_/A _74147_/X sky130_fd_sc_hd__a21o_4
X_40539_ _40538_/X _40508_/X _88374_/Q _40510_/X _88374_/D sky130_fd_sc_hd__a2bb2o_4
X_47095_ _47090_/Y _47081_/X _47094_/X _86671_/D sky130_fd_sc_hd__a21oi_4
X_71359_ _71504_/C _71351_/X _70778_/A _71363_/D _71359_/X sky130_fd_sc_hd__and4_4
X_61112_ _61112_/A _61112_/X sky130_fd_sc_hd__buf_2
X_46046_ _40556_/A _46046_/X sky130_fd_sc_hd__buf_2
X_43258_ _43241_/X _43244_/X _41082_/X _87513_/Q _43250_/X _43259_/A
+ sky130_fd_sc_hd__o32ai_4
X_62092_ _62055_/A _84913_/Q _61755_/X _61728_/A _62092_/X sky130_fd_sc_hd__and4_4
X_78955_ _78940_/A _82513_/D _78954_/X _78956_/B sky130_fd_sc_hd__o21ai_4
X_74078_ _44725_/Y _73491_/X _74077_/Y _74078_/X sky130_fd_sc_hd__a21o_4
X_42209_ _42258_/A _42209_/X sky130_fd_sc_hd__buf_2
X_65920_ _65654_/X _86240_/Q _65761_/X _65919_/X _65920_/X sky130_fd_sc_hd__a211o_4
X_61043_ _61004_/Y _61030_/Y _61042_/Y _84530_/Q _59509_/X _61043_/X
+ sky130_fd_sc_hd__o32a_4
X_77906_ _77906_/A _77908_/A sky130_fd_sc_hd__inv_2
X_73029_ _88329_/Q _73026_/X _73028_/X _73029_/Y sky130_fd_sc_hd__o21ai_4
X_43189_ _43189_/A _53944_/A sky130_fd_sc_hd__buf_2
X_78886_ _78886_/A _78896_/A _78886_/Y sky130_fd_sc_hd__nor2_4
X_49805_ _57958_/B _49798_/X _49804_/Y _49805_/Y sky130_fd_sc_hd__o21ai_4
X_65851_ _65812_/A _86501_/Q _65851_/X sky130_fd_sc_hd__and2_4
X_77837_ _77826_/Y _81933_/D sky130_fd_sc_hd__inv_2
X_47997_ _47989_/Y _47954_/X _47996_/X _47997_/Y sky130_fd_sc_hd__a21oi_4
X_64802_ _64650_/X _86170_/Q _64776_/X _64801_/X _64802_/X sky130_fd_sc_hd__a211o_4
X_49736_ _49716_/X _52950_/B _49736_/Y sky130_fd_sc_hd__nand2_4
X_68570_ _69796_/A _68570_/X sky130_fd_sc_hd__buf_2
X_46948_ _46948_/A _52768_/B _46948_/Y sky130_fd_sc_hd__nand2_4
X_65782_ _65782_/A _65812_/A sky130_fd_sc_hd__buf_2
X_77768_ _82150_/Q _77768_/B _77768_/X sky130_fd_sc_hd__xor2_4
X_62994_ _63306_/A _63285_/B sky130_fd_sc_hd__buf_2
X_67521_ _81498_/D _67449_/X _67520_/X _84066_/D sky130_fd_sc_hd__a21bo_4
X_79507_ _79491_/Y _79494_/Y _79506_/X _79507_/X sky130_fd_sc_hd__a21o_4
X_64733_ _64600_/A _64733_/X sky130_fd_sc_hd__buf_2
X_76719_ _76719_/A _76718_/Y _76719_/Y sky130_fd_sc_hd__nand2_4
X_49667_ _86345_/Q _49660_/X _49666_/Y _49667_/Y sky130_fd_sc_hd__o21ai_4
X_61945_ _59765_/A _61945_/X sky130_fd_sc_hd__buf_2
X_46879_ _52726_/B _51037_/B sky130_fd_sc_hd__buf_2
X_77699_ _77712_/A _82124_/Q _77699_/X sky130_fd_sc_hd__xor2_4
X_48618_ _81770_/Q _48618_/Y sky130_fd_sc_hd__inv_2
X_67452_ _87982_/Q _67355_/X _67405_/X _67451_/X _67452_/X sky130_fd_sc_hd__a211o_4
X_79438_ _79438_/A _79438_/B _79459_/A sky130_fd_sc_hd__xor2_4
X_64664_ _64661_/Y _64662_/X _64663_/X _84231_/D sky130_fd_sc_hd__a21o_4
X_49598_ _49610_/A _49592_/B _49577_/C _52811_/D _49598_/X sky130_fd_sc_hd__and4_4
X_61876_ _84880_/Q _61876_/X sky130_fd_sc_hd__buf_2
X_66403_ _66399_/Y _66377_/X _66402_/Y _84130_/D sky130_fd_sc_hd__a21o_4
X_63615_ _63615_/A _63615_/B _80413_/B _63615_/Y sky130_fd_sc_hd__nor3_4
X_48549_ _49223_/A _49212_/A sky130_fd_sc_hd__buf_2
X_60827_ _60692_/X _60825_/Y _60708_/Y _60795_/X _60826_/Y _84557_/D
+ sky130_fd_sc_hd__a41oi_4
X_67383_ _67025_/X _67383_/X sky130_fd_sc_hd__buf_2
X_79369_ _79362_/X _79369_/B _79369_/Y sky130_fd_sc_hd__nand2_4
X_64595_ _64588_/X _64594_/X _59297_/A _64595_/X sky130_fd_sc_hd__a21o_4
X_81400_ _81351_/CLK _81400_/D _76696_/B sky130_fd_sc_hd__dfxtp_4
X_69122_ _69134_/A _69122_/B _69122_/X sky130_fd_sc_hd__and2_4
X_66334_ _57694_/X _66334_/B _66334_/X sky130_fd_sc_hd__and2_4
X_51560_ _51556_/Y _51557_/X _51559_/X _85988_/D sky130_fd_sc_hd__a21oi_4
X_63546_ _63546_/A _58533_/A _63520_/C _63546_/D _63546_/X sky130_fd_sc_hd__and4_4
X_82380_ _82381_/CLK _82188_/Q _82380_/Q sky130_fd_sc_hd__dfxtp_4
X_60758_ _60703_/Y _60758_/X sky130_fd_sc_hd__buf_2
X_50511_ _50511_/A _50526_/B _50526_/C _50511_/X sky130_fd_sc_hd__and3_4
X_81331_ _83926_/CLK _76407_/X _81707_/D sky130_fd_sc_hd__dfxtp_4
X_69053_ _69735_/A _69053_/B _69053_/Y sky130_fd_sc_hd__nor2_4
X_66265_ _66261_/Y _66205_/X _66264_/Y _84145_/D sky130_fd_sc_hd__a21o_4
X_51491_ _51491_/A _53017_/B _51491_/Y sky130_fd_sc_hd__nand2_4
X_63477_ _61437_/B _63426_/X _63474_/X _63476_/X _63477_/X sky130_fd_sc_hd__a211o_4
X_60689_ _60632_/X _60714_/A _60713_/A _60689_/Y sky130_fd_sc_hd__o21ai_4
X_68004_ _86947_/Q _67906_/X _67908_/X _68003_/X _68004_/X sky130_fd_sc_hd__a211o_4
X_53230_ _53217_/A _53244_/B _53222_/X _53230_/D _53230_/X sky130_fd_sc_hd__and4_4
X_65216_ _65164_/A _86410_/Q _65216_/X sky130_fd_sc_hd__and2_4
X_84050_ _84049_/CLK _84050_/D _81482_/D sky130_fd_sc_hd__dfxtp_4
X_50442_ _50510_/A _50462_/C sky130_fd_sc_hd__buf_2
X_62428_ _62193_/A _62608_/D sky130_fd_sc_hd__buf_2
X_81262_ _81296_/CLK _81262_/D _76328_/A sky130_fd_sc_hd__dfxtp_4
X_66196_ _65763_/A _85901_/Q _66196_/X sky130_fd_sc_hd__and2_4
X_83001_ _83001_/CLK _83001_/D _45526_/A sky130_fd_sc_hd__dfxtp_4
X_80213_ _57753_/Y _65498_/C _80212_/Y _80213_/X sky130_fd_sc_hd__o21a_4
X_53161_ _53147_/X _53161_/B _53161_/Y sky130_fd_sc_hd__nand2_4
X_65147_ _65227_/A _65147_/B _65147_/X sky130_fd_sc_hd__and2_4
X_50373_ _50371_/Y _50351_/X _50372_/Y _50373_/Y sky130_fd_sc_hd__a21boi_4
X_62359_ _62319_/A _58511_/A _62319_/C _62359_/Y sky130_fd_sc_hd__nand3_4
X_81193_ _81190_/CLK _74949_/X _49129_/A sky130_fd_sc_hd__dfxtp_4
X_52112_ _72836_/B _52089_/X _52111_/Y _52112_/Y sky130_fd_sc_hd__o21ai_4
X_80144_ _60047_/C _63914_/C _80144_/X sky130_fd_sc_hd__xor2_4
X_53092_ _52126_/A _53172_/A sky130_fd_sc_hd__buf_2
X_65078_ _65075_/X _65077_/X _64574_/X _65078_/X sky130_fd_sc_hd__a21o_4
X_69955_ _69988_/A _69955_/X sky130_fd_sc_hd__buf_2
X_52043_ _52070_/A _50341_/B _52043_/Y sky130_fd_sc_hd__nand2_4
X_56920_ _56552_/Y _56920_/B _56921_/C sky130_fd_sc_hd__nand2_4
X_68906_ _83956_/Q _68838_/X _68905_/X _83956_/D sky130_fd_sc_hd__a21bo_4
X_64029_ _64420_/B _64029_/B _64029_/C _64029_/D _64029_/Y sky130_fd_sc_hd__nand4_4
X_87740_ _87487_/CLK _42749_/Y _68941_/B sky130_fd_sc_hd__dfxtp_4
X_84952_ _85404_/CLK _84952_/D _84952_/Q sky130_fd_sc_hd__dfxtp_4
X_80075_ _80074_/B _80058_/X _80075_/X sky130_fd_sc_hd__and2_4
X_69886_ _73374_/A _69837_/X _69779_/X _69885_/Y _69886_/X sky130_fd_sc_hd__a211o_4
X_83903_ _81975_/CLK _83903_/D _81975_/D sky130_fd_sc_hd__dfxtp_4
X_56851_ _56848_/X _56850_/X _56842_/X _56851_/X sky130_fd_sc_hd__o21a_4
X_68837_ _83959_/Q _68713_/X _68836_/X _68837_/X sky130_fd_sc_hd__a21bo_4
X_87671_ _87671_/CLK _87671_/D _67248_/B sky130_fd_sc_hd__dfxtp_4
X_84883_ _84883_/CLK _58306_/Y _64546_/C sky130_fd_sc_hd__dfxtp_4
X_55802_ _55802_/A _55802_/X sky130_fd_sc_hd__buf_2
X_86622_ _85981_/CLK _47560_/Y _72162_/A sky130_fd_sc_hd__dfxtp_4
X_59570_ _59570_/A _60639_/A sky130_fd_sc_hd__inv_2
X_83834_ _83191_/CLK _83834_/D _83834_/Q sky130_fd_sc_hd__dfxtp_4
X_56782_ _56729_/X _56782_/X sky130_fd_sc_hd__buf_2
X_68768_ _68542_/X _68768_/B _68768_/X sky130_fd_sc_hd__and2_4
X_53994_ _53992_/Y _53982_/X _53993_/Y _53994_/Y sky130_fd_sc_hd__a21boi_4
Xclkbuf_10_542_0_CLK clkbuf_9_271_0_CLK/X _84020_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_33_0_CLK clkbuf_6_33_0_CLK/A clkbuf_7_67_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_58521_ _58517_/X _58518_/Y _58520_/Y _58521_/Y sky130_fd_sc_hd__a21oi_4
X_55733_ _56450_/C _55126_/A _55128_/A _55732_/X _55733_/X sky130_fd_sc_hd__a211o_4
X_67719_ _67615_/X _67719_/B _67719_/X sky130_fd_sc_hd__and2_4
X_86553_ _86553_/CLK _86553_/D _66028_/B sky130_fd_sc_hd__dfxtp_4
X_52945_ _85725_/Q _52929_/X _52944_/Y _52945_/Y sky130_fd_sc_hd__o21ai_4
X_83765_ _83763_/CLK _70481_/X _83765_/Q sky130_fd_sc_hd__dfxtp_4
X_80977_ _81061_/CLK _75712_/X _75109_/B sky130_fd_sc_hd__dfxtp_4
X_68699_ _69092_/A _68699_/B _68699_/X sky130_fd_sc_hd__and2_4
X_85504_ _85505_/CLK _85504_/D _85504_/Q sky130_fd_sc_hd__dfxtp_4
X_70730_ _71266_/A _70730_/X sky130_fd_sc_hd__buf_2
X_58452_ _58452_/A _58498_/B _58452_/Y sky130_fd_sc_hd__nand2_4
X_82716_ _82715_/CLK _82716_/D _82672_/D sky130_fd_sc_hd__dfxtp_4
X_55664_ _55662_/Y _55663_/Y _55664_/Y sky130_fd_sc_hd__nand2_4
X_86484_ _86196_/CLK _48780_/Y _86484_/Q sky130_fd_sc_hd__dfxtp_4
X_40890_ _40889_/Y _40890_/X sky130_fd_sc_hd__buf_2
X_52876_ _52885_/A _52876_/B _52876_/Y sky130_fd_sc_hd__nand2_4
X_83696_ _85645_/CLK _70811_/Y _47157_/A sky130_fd_sc_hd__dfxtp_4
X_57403_ _57394_/X _56630_/X _85014_/Q _57395_/X _57403_/X sky130_fd_sc_hd__a2bb2o_4
X_88223_ _88232_/CLK _88223_/D _67813_/B sky130_fd_sc_hd__dfxtp_4
X_54615_ _85409_/Q _54593_/X _54614_/Y _54615_/Y sky130_fd_sc_hd__o21ai_4
X_85435_ _85754_/CLK _85435_/D _85435_/Q sky130_fd_sc_hd__dfxtp_4
X_51827_ _85939_/Q _51817_/X _51826_/Y _51827_/Y sky130_fd_sc_hd__o21ai_4
X_70661_ _70886_/A _70884_/A sky130_fd_sc_hd__buf_2
X_58383_ _58383_/A _58369_/X _58383_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_557_0_CLK clkbuf_9_278_0_CLK/X _87922_/CLK sky130_fd_sc_hd__clkbuf_1
X_82647_ _84003_/CLK _83999_/Q _82647_/Q sky130_fd_sc_hd__dfxtp_4
X_55595_ _45440_/A _55571_/X _44049_/X _55594_/Y _55595_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_6_48_0_CLK clkbuf_6_49_0_CLK/A clkbuf_7_96_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_72400_ _72461_/A _72400_/B _72400_/Y sky130_fd_sc_hd__nor2_4
X_57334_ _45947_/B _85033_/Q _57333_/X _57331_/B _57335_/B sky130_fd_sc_hd__a211o_4
X_88154_ _88220_/CLK _41764_/Y _67932_/B sky130_fd_sc_hd__dfxtp_4
X_54546_ _54546_/A _53369_/B _54546_/Y sky130_fd_sc_hd__nand2_4
X_42560_ _72945_/A _69661_/B sky130_fd_sc_hd__inv_2
X_73380_ _73378_/X _86185_/Q _72905_/X _73379_/X _73380_/X sky130_fd_sc_hd__a211o_4
X_85366_ _83630_/CLK _54853_/Y _85366_/Q sky130_fd_sc_hd__dfxtp_4
X_51758_ _51758_/A _50893_/B _51758_/Y sky130_fd_sc_hd__nand2_4
X_70592_ _74731_/A _74716_/A sky130_fd_sc_hd__buf_2
X_82578_ _82610_/CLK _82578_/D _78199_/A sky130_fd_sc_hd__dfxtp_4
X_87105_ _87926_/CLK _87105_/D _87105_/Q sky130_fd_sc_hd__dfxtp_4
X_41511_ _41510_/Y _41511_/X sky130_fd_sc_hd__buf_2
X_72331_ _72366_/A _86288_/Q _72331_/Y sky130_fd_sc_hd__nor2_4
X_84317_ _84321_/CLK _63518_/Y _63517_/C sky130_fd_sc_hd__dfxtp_4
X_50709_ _86149_/Q _50706_/X _50708_/Y _50709_/Y sky130_fd_sc_hd__o21ai_4
X_81529_ _82053_/CLK _81541_/Q _81529_/Q sky130_fd_sc_hd__dfxtp_4
X_57265_ _57331_/B _57264_/Y _56664_/Y _56972_/Y _57265_/X sky130_fd_sc_hd__a2bb2o_4
X_42491_ _42466_/X _42467_/X _40656_/X _68668_/A _42480_/X _42492_/A
+ sky130_fd_sc_hd__o32ai_4
X_88085_ _88085_/CLK _88085_/D _88085_/Q sky130_fd_sc_hd__dfxtp_4
X_54477_ _54474_/Y _54475_/X _54476_/X _85435_/D sky130_fd_sc_hd__a21oi_4
X_85297_ _85297_/CLK _56097_/Y _85297_/Q sky130_fd_sc_hd__dfxtp_4
X_51689_ _51695_/A _51684_/B _51695_/C _53211_/D _51689_/X sky130_fd_sc_hd__and4_4
X_59004_ _59000_/Y _59003_/Y _58966_/X _59004_/X sky130_fd_sc_hd__a21o_4
X_44230_ _56995_/A _44231_/A sky130_fd_sc_hd__buf_2
X_56216_ _56214_/A _56205_/X _56216_/C _56216_/Y sky130_fd_sc_hd__nand3_4
X_75050_ _75039_/X _75042_/A _75042_/B _75050_/Y sky130_fd_sc_hd__nand3_4
X_41442_ _41441_/X _41442_/X sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_0 _46167_/Y _86769_/D sky130_fd_sc_hd__buf_8
X_87036_ _86989_/CLK _44608_/X _87036_/Q sky130_fd_sc_hd__dfxtp_4
X_53428_ _53347_/A _53428_/X sky130_fd_sc_hd__buf_2
X_72262_ _83270_/Q _72250_/X _72254_/X _72261_/X _83270_/D sky130_fd_sc_hd__a2bb2oi_4
X_84248_ _84849_/CLK _64417_/X _79700_/B sky130_fd_sc_hd__dfxtp_4
X_57196_ _56859_/X _56675_/X _56876_/X _57196_/Y sky130_fd_sc_hd__nand3_4
X_74001_ _48022_/Y _74001_/B _74002_/B sky130_fd_sc_hd__xor2_4
X_71213_ _71211_/A _71091_/B _71219_/C _71213_/Y sky130_fd_sc_hd__nand3_4
X_56147_ _56147_/A _56117_/A _56148_/A sky130_fd_sc_hd__xor2_4
X_44161_ _44159_/X _44160_/Y _44163_/B _87185_/D sky130_fd_sc_hd__a21oi_4
X_41373_ _41072_/X _41373_/X sky130_fd_sc_hd__buf_2
X_53359_ _53354_/Y _53355_/X _53358_/X _85649_/D sky130_fd_sc_hd__a21oi_4
X_72193_ _72193_/A _72193_/B _72193_/Y sky130_fd_sc_hd__nor2_4
X_84179_ _84175_/CLK _84179_/D _84179_/Q sky130_fd_sc_hd__dfxtp_4
X_43112_ _43112_/A _87572_/D sky130_fd_sc_hd__inv_2
X_40324_ _49140_/B _40324_/X sky130_fd_sc_hd__buf_2
X_71144_ _48368_/X _71138_/X _71143_/Y _83592_/D sky130_fd_sc_hd__o21ai_4
X_44092_ _80666_/Q _55158_/A sky130_fd_sc_hd__inv_2
X_56078_ _55863_/X _55995_/X _56079_/A sky130_fd_sc_hd__xnor2_4
X_47920_ _50270_/A _49312_/C _47919_/X _47920_/X sky130_fd_sc_hd__and3_4
X_43043_ _43043_/A _43043_/Y sky130_fd_sc_hd__inv_2
X_55029_ _85332_/Q _55020_/X _55028_/Y _55029_/Y sky130_fd_sc_hd__o21ai_4
X_59906_ _60418_/D _61070_/B _59906_/X sky130_fd_sc_hd__and2_4
X_78740_ _78701_/A _78701_/B _78700_/A _78720_/A _78740_/X sky130_fd_sc_hd__and4_4
X_71075_ _70809_/A _71076_/B sky130_fd_sc_hd__buf_2
X_75952_ _81702_/D _75952_/B _75952_/Y sky130_fd_sc_hd__nand2_4
X_87938_ _88128_/CLK _87938_/D _87938_/Q sky130_fd_sc_hd__dfxtp_4
X_74903_ _74887_/C _74899_/Y _74902_/Y _74904_/B sky130_fd_sc_hd__o21a_4
X_70026_ _68674_/X _68677_/X _70005_/X _70026_/Y sky130_fd_sc_hd__a21oi_4
X_47851_ _47848_/X _47851_/B _47851_/X sky130_fd_sc_hd__and2_4
X_59837_ _59772_/A _59837_/B _80391_/A _59837_/Y sky130_fd_sc_hd__nor3_4
X_78671_ _78638_/A _78653_/X _78638_/B _78655_/B _78671_/X sky130_fd_sc_hd__and4_4
X_87869_ _82888_/CLK _42427_/Y _87869_/Q sky130_fd_sc_hd__dfxtp_4
X_75883_ _75750_/Y _75883_/Y sky130_fd_sc_hd__inv_2
X_46802_ _46784_/A _46830_/B _46784_/C _52681_/D _46802_/X sky130_fd_sc_hd__and4_4
X_77622_ _77622_/A _77596_/A _77622_/X sky130_fd_sc_hd__and2_4
X_74834_ _74844_/A _46114_/A _74835_/A sky130_fd_sc_hd__nand2_4
X_47782_ _86598_/Q _47760_/X _47781_/Y _47782_/Y sky130_fd_sc_hd__o21ai_4
X_59768_ _61770_/B _59731_/Y _61770_/D _59836_/D _59816_/A _59768_/Y
+ sky130_fd_sc_hd__a41oi_4
X_44994_ _45835_/A _45219_/A sky130_fd_sc_hd__buf_2
X_49521_ _49548_/A _49522_/C sky130_fd_sc_hd__buf_2
X_46733_ _46733_/A _51812_/B _46733_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_1_0_CLK clkbuf_8_1_0_CLK/A clkbuf_9_3_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_58719_ _58713_/Y _58718_/Y _58646_/X _58719_/X sky130_fd_sc_hd__a21o_4
X_77553_ _77553_/A _77553_/B _77552_/Y _77553_/X sky130_fd_sc_hd__or3_4
X_43945_ _43945_/A _43945_/Y sky130_fd_sc_hd__inv_2
X_74765_ _70576_/X _83828_/Q _74764_/A _74765_/X sky130_fd_sc_hd__and3_4
X_71977_ _83309_/Q _57615_/X _71976_/Y _71977_/Y sky130_fd_sc_hd__o21ai_4
X_59699_ _59699_/A _59722_/A _61755_/A _59797_/A sky130_fd_sc_hd__and3_4
X_76504_ _76503_/Y _76504_/Y sky130_fd_sc_hd__inv_2
X_49452_ _49447_/A _49456_/B _49447_/C _46775_/X _49452_/X sky130_fd_sc_hd__and4_4
X_73716_ _73716_/A _73715_/X _73717_/B sky130_fd_sc_hd__nand2_4
X_61730_ _59806_/A _61730_/X sky130_fd_sc_hd__buf_2
X_46664_ _58634_/A _46622_/X _46663_/Y _46664_/Y sky130_fd_sc_hd__o21ai_4
X_70928_ _70903_/A _70863_/C _70925_/X _70919_/D _70928_/Y sky130_fd_sc_hd__nand4_4
X_77484_ _77481_/Y _77484_/B _82195_/D sky130_fd_sc_hd__xor2_4
X_43876_ _43854_/A _43876_/X sky130_fd_sc_hd__buf_2
X_74696_ _74695_/X _82982_/D sky130_fd_sc_hd__inv_2
X_48403_ _49247_/A _48403_/X sky130_fd_sc_hd__buf_2
X_79223_ _79221_/Y _79217_/Y _79218_/X _79224_/B sky130_fd_sc_hd__nand3_4
X_45615_ _85011_/Q _45615_/Y sky130_fd_sc_hd__inv_2
X_76435_ _76433_/X _76435_/B _76435_/Y sky130_fd_sc_hd__xnor2_4
X_42827_ _41469_/X _42821_/X _66626_/B _42822_/X _87697_/D sky130_fd_sc_hd__a2bb2o_4
X_49383_ _58613_/B _49360_/X _49382_/Y _49383_/Y sky130_fd_sc_hd__o21ai_4
X_61661_ _61690_/A _61690_/B _79130_/B _61661_/Y sky130_fd_sc_hd__nor3_4
X_73647_ _73645_/X _73646_/Y _73546_/X _73647_/X sky130_fd_sc_hd__a21o_4
X_70859_ _70866_/A _70863_/C sky130_fd_sc_hd__buf_2
X_46595_ _52571_/B _51394_/B sky130_fd_sc_hd__buf_2
X_63400_ _63400_/A _63400_/B _63400_/C _63400_/X sky130_fd_sc_hd__and3_4
X_48334_ _49223_/A _48401_/A sky130_fd_sc_hd__buf_2
X_60612_ _60612_/A _60612_/B _60612_/C _60612_/Y sky130_fd_sc_hd__nor3_4
X_79154_ _79154_/A _79154_/B _82462_/D sky130_fd_sc_hd__xor2_4
X_45546_ _45540_/X _45543_/X _45545_/Y _45546_/Y sky130_fd_sc_hd__a21oi_4
X_76366_ _76366_/A _76366_/B _76369_/B sky130_fd_sc_hd__nor2_4
X_64380_ _64263_/A _64380_/X sky130_fd_sc_hd__buf_2
X_42758_ _42680_/A _42822_/A sky130_fd_sc_hd__buf_2
X_73578_ _68387_/B _73030_/X _73486_/X _73577_/Y _73578_/X sky130_fd_sc_hd__a211o_4
X_61592_ _61400_/X _61619_/C sky130_fd_sc_hd__buf_2
X_78105_ _78103_/Y _78099_/Y _78104_/Y _78105_/Y sky130_fd_sc_hd__o21ai_4
X_75317_ _81075_/Q _75317_/Y sky130_fd_sc_hd__inv_2
X_63331_ _60454_/A _64535_/B _60441_/B _60473_/B _63331_/X sky130_fd_sc_hd__and4_4
X_41709_ _41628_/X _81746_/Q _41708_/X _41709_/X sky130_fd_sc_hd__o21a_4
X_48265_ _48264_/X _50310_/B _48265_/Y sky130_fd_sc_hd__nand2_4
X_60543_ _60481_/A _60543_/B _60542_/Y _60543_/Y sky130_fd_sc_hd__nand3_4
X_72529_ _72528_/Y _72550_/C _72529_/C _72530_/A sky130_fd_sc_hd__nand3_4
X_79085_ _82800_/D _82544_/Q _79086_/B sky130_fd_sc_hd__xnor2_4
X_45477_ _45474_/Y _45412_/X _45443_/X _45476_/Y _45477_/X sky130_fd_sc_hd__a211o_4
X_76297_ _81356_/Q _76297_/B _76297_/X sky130_fd_sc_hd__xor2_4
X_42689_ _42687_/X _42688_/X _41082_/X _87769_/Q _42673_/X _42689_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47216_ _82370_/Q _54612_/D sky130_fd_sc_hd__inv_2
X_66050_ _65992_/A _85911_/Q _66050_/X sky130_fd_sc_hd__and2_4
X_78036_ _78033_/A _82177_/Q _78033_/B _78037_/B sky130_fd_sc_hd__nand3_4
X_44428_ _44352_/X _44428_/X sky130_fd_sc_hd__buf_2
X_63262_ _60458_/X _63332_/D sky130_fd_sc_hd__buf_2
X_75248_ _75243_/Y _75219_/Y _75247_/X _75248_/Y sky130_fd_sc_hd__o21ai_4
X_60474_ _60493_/A _60556_/B _60475_/A sky130_fd_sc_hd__nand2_4
X_48196_ _48196_/A _46487_/B _48195_/X _48196_/X sky130_fd_sc_hd__and3_4
X_65001_ _64999_/X _86130_/Q _64927_/X _65000_/X _65001_/X sky130_fd_sc_hd__a211o_4
X_62213_ _62572_/A _62214_/A sky130_fd_sc_hd__buf_2
X_47147_ _47147_/A _47150_/A sky130_fd_sc_hd__buf_2
X_44359_ _41731_/X _44345_/X _87148_/Q _44346_/X _87148_/D sky130_fd_sc_hd__a2bb2o_4
X_63193_ _60458_/X _63239_/D sky130_fd_sc_hd__buf_2
X_75179_ _75179_/A _75179_/Y sky130_fd_sc_hd__inv_2
X_62144_ _62144_/A _62121_/X _78053_/B _62144_/Y sky130_fd_sc_hd__nor3_4
X_47078_ _53360_/B _52843_/B sky130_fd_sc_hd__buf_2
X_79987_ _79985_/Y _79972_/Y _79973_/Y _79988_/B sky130_fd_sc_hd__nand3_4
X_46029_ _45962_/X _46029_/X sky130_fd_sc_hd__buf_2
X_69740_ _69680_/A _69740_/B _69740_/X sky130_fd_sc_hd__and2_4
X_66952_ _66949_/X _66951_/X _66905_/X _66952_/X sky130_fd_sc_hd__a21o_4
X_62075_ _84891_/Q _63629_/B sky130_fd_sc_hd__buf_2
X_78938_ _78938_/A _78952_/A _78939_/B sky130_fd_sc_hd__xor2_4
X_65903_ _65516_/A _65903_/X sky130_fd_sc_hd__buf_2
X_61026_ _60968_/X _61024_/Y _61025_/X _84536_/Q _61020_/X _84536_/D
+ sky130_fd_sc_hd__o32a_4
X_69671_ _81978_/D _69632_/X _69670_/X _83906_/D sky130_fd_sc_hd__a21bo_4
X_66883_ _66647_/A _66956_/A sky130_fd_sc_hd__buf_2
X_78869_ _78869_/A _78869_/B _78869_/X sky130_fd_sc_hd__xor2_4
X_80900_ _84074_/CLK _80900_/D _80900_/Q sky130_fd_sc_hd__dfxtp_4
X_68622_ _86997_/Q _68472_/X _68473_/X _68621_/X _68622_/X sky130_fd_sc_hd__a211o_4
X_65834_ _57788_/X _85862_/Q _65834_/X sky130_fd_sc_hd__and2_4
X_81880_ _81928_/CLK _78071_/X _81880_/Q sky130_fd_sc_hd__dfxtp_4
X_49719_ _49708_/A _49697_/B _49724_/C _52934_/D _49719_/X sky130_fd_sc_hd__and4_4
X_80831_ _81065_/CLK _83975_/Q _80831_/Q sky130_fd_sc_hd__dfxtp_4
X_68553_ _68553_/A _87340_/Q _68553_/X sky130_fd_sc_hd__and2_4
X_65765_ _65735_/A _86475_/Q _65765_/X sky130_fd_sc_hd__and2_4
X_50991_ _50991_/A _51101_/A sky130_fd_sc_hd__buf_2
X_62977_ _62988_/A _62988_/B _84364_/Q _62977_/Y sky130_fd_sc_hd__nor3_4
X_67504_ _67575_/A _88172_/Q _67504_/X sky130_fd_sc_hd__and2_4
X_52730_ _52729_/X _52724_/B _52708_/X _52730_/D _52730_/X sky130_fd_sc_hd__and4_4
X_64716_ _65790_/A _64716_/X sky130_fd_sc_hd__buf_2
X_83550_ _83550_/CLK _83550_/D _47704_/A sky130_fd_sc_hd__dfxtp_4
X_61928_ _61926_/Y _61881_/X _61927_/Y _84445_/D sky130_fd_sc_hd__a21oi_4
X_68484_ _68481_/X _68483_/X _68429_/X _68484_/X sky130_fd_sc_hd__a21o_4
X_80762_ _81994_/CLK _75440_/X _80762_/Q sky130_fd_sc_hd__dfxtp_4
X_65696_ _65533_/X _65694_/Y _65695_/Y _65696_/Y sky130_fd_sc_hd__o21ai_4
X_82501_ _82942_/CLK _82501_/D _78356_/A sky130_fd_sc_hd__dfxtp_4
X_67435_ _87163_/Q _67432_/X _67433_/X _67434_/X _67435_/X sky130_fd_sc_hd__a211o_4
X_52661_ _52648_/X _52661_/B _52654_/C _52661_/D _52661_/X sky130_fd_sc_hd__and4_4
X_64647_ _64773_/A _64647_/B _64647_/X sky130_fd_sc_hd__and2_4
X_83481_ _83415_/CLK _71490_/X _83481_/Q sky130_fd_sc_hd__dfxtp_4
X_61859_ _59823_/X _61860_/D sky130_fd_sc_hd__buf_2
X_80693_ _80697_/CLK _80725_/Q _80693_/Q sky130_fd_sc_hd__dfxtp_4
X_54400_ _54400_/A _54401_/A sky130_fd_sc_hd__buf_2
X_85220_ _85186_/CLK _85220_/D _55722_/B sky130_fd_sc_hd__dfxtp_4
X_51612_ _85978_/Q _51594_/X _51611_/Y _51612_/Y sky130_fd_sc_hd__o21ai_4
X_82432_ _82462_/CLK _82464_/Q _78788_/A sky130_fd_sc_hd__dfxtp_4
X_55380_ _55383_/A _55377_/Y _55379_/Y _55380_/Y sky130_fd_sc_hd__a21oi_4
X_67366_ _87166_/Q _67311_/X _67313_/X _67365_/X _67366_/X sky130_fd_sc_hd__a211o_4
X_52592_ _52496_/A _52592_/X sky130_fd_sc_hd__buf_2
X_64578_ _44170_/A _64772_/A sky130_fd_sc_hd__buf_2
XPHY_707 sky130_fd_sc_hd__decap_3
X_69105_ _87073_/Q _69058_/X _69103_/X _69104_/X _69105_/X sky130_fd_sc_hd__a211o_4
X_54331_ _54328_/Y _54311_/X _54330_/X _85462_/D sky130_fd_sc_hd__a21oi_4
X_66317_ _66294_/X _66315_/Y _66316_/Y _66317_/Y sky130_fd_sc_hd__o21ai_4
X_85151_ _85213_/CLK _85151_/D _55622_/B sky130_fd_sc_hd__dfxtp_4
X_51543_ _51521_/X _51553_/B _51533_/C _53070_/D _51543_/X sky130_fd_sc_hd__and4_4
X_63529_ _63468_/A _63554_/B sky130_fd_sc_hd__buf_2
X_82363_ _84981_/CLK _82363_/D _82363_/Q sky130_fd_sc_hd__dfxtp_4
X_67297_ _87413_/Q _67274_/X _67226_/X _67296_/X _67297_/X sky130_fd_sc_hd__a211o_4
X_84102_ _81169_/CLK _84102_/D _84102_/Q sky130_fd_sc_hd__dfxtp_4
X_57050_ _57050_/A _56953_/A _57051_/A sky130_fd_sc_hd__nand2_4
X_81314_ _84020_/CLK _76157_/X _81722_/D sky130_fd_sc_hd__dfxtp_4
X_69036_ _69032_/X _69034_/X _69035_/X _69036_/X sky130_fd_sc_hd__a21o_4
X_54262_ _85474_/Q _54249_/X _54261_/Y _54262_/Y sky130_fd_sc_hd__o21ai_4
X_66248_ _66246_/Y _66205_/X _66247_/X _84146_/D sky130_fd_sc_hd__a21o_4
X_85082_ _85083_/CLK _85082_/D _45500_/A sky130_fd_sc_hd__dfxtp_4
X_51474_ _51470_/Y _51448_/X _51473_/X _51474_/Y sky130_fd_sc_hd__a21oi_4
X_82294_ _82103_/CLK _81918_/Q _82294_/Q sky130_fd_sc_hd__dfxtp_4
X_56001_ _56001_/A _55927_/X _55956_/B _74297_/C _56002_/A sky130_fd_sc_hd__nand4_4
X_53213_ _53219_/A _53213_/B _53213_/Y sky130_fd_sc_hd__nand2_4
X_84033_ _81154_/CLK _84033_/D _82073_/D sky130_fd_sc_hd__dfxtp_4
X_50425_ _48744_/A _50430_/B _50435_/C _50425_/X sky130_fd_sc_hd__and3_4
X_81245_ _85342_/CLK _81053_/Q _81245_/Q sky130_fd_sc_hd__dfxtp_4
X_54193_ _54249_/A _54193_/X sky130_fd_sc_hd__buf_2
X_66179_ _66366_/A _66179_/X sky130_fd_sc_hd__buf_2
X_53144_ _53139_/A _53133_/B _53143_/X _53144_/D _53144_/X sky130_fd_sc_hd__and4_4
X_50356_ _50356_/A _50356_/B _50356_/Y sky130_fd_sc_hd__nand2_4
X_81176_ _82335_/CLK _75007_/B _81176_/Q sky130_fd_sc_hd__dfxtp_4
X_80127_ _80109_/X _80112_/Y _80127_/X sky130_fd_sc_hd__or2_4
X_53075_ _53073_/Y _53056_/X _53074_/X _85702_/D sky130_fd_sc_hd__a21oi_4
X_57952_ _57952_/A _57952_/B _57952_/Y sky130_fd_sc_hd__nor2_4
X_69938_ _70012_/A _69938_/X sky130_fd_sc_hd__buf_2
X_50287_ _48234_/A _50475_/B _50257_/X _50287_/Y sky130_fd_sc_hd__nand3_4
X_85984_ _85697_/CLK _51581_/Y _85984_/Q sky130_fd_sc_hd__dfxtp_4
X_52026_ _52020_/Y _52022_/X _52025_/Y _85904_/D sky130_fd_sc_hd__a21boi_4
X_56903_ _46237_/A _56901_/Y _56902_/Y _56903_/X sky130_fd_sc_hd__o21a_4
X_87723_ _86930_/CLK _42778_/X _87723_/Q sky130_fd_sc_hd__dfxtp_4
X_84935_ _86317_/CLK _84935_/D _84935_/Q sky130_fd_sc_hd__dfxtp_4
X_80058_ _57980_/Y _65728_/C _80057_/Y _80058_/X sky130_fd_sc_hd__o21a_4
X_57883_ _84942_/Q _57883_/Y sky130_fd_sc_hd__inv_2
X_69869_ _81963_/D _69831_/X _69868_/X _69869_/X sky130_fd_sc_hd__a21bo_4
Xclkbuf_10_481_0_CLK clkbuf_9_240_0_CLK/X _86610_/CLK sky130_fd_sc_hd__clkbuf_1
X_71900_ _74523_/A _71893_/X _71755_/X _71898_/D _71900_/Y sky130_fd_sc_hd__nand4_4
X_59622_ _59622_/A _60615_/A sky130_fd_sc_hd__inv_2
X_56834_ _56832_/X _55681_/X _56833_/Y _56838_/A sky130_fd_sc_hd__a21o_4
X_87654_ _86930_/CLK _42913_/X _67652_/B sky130_fd_sc_hd__dfxtp_4
X_72880_ _72880_/A _72880_/X sky130_fd_sc_hd__buf_2
X_84866_ _84299_/CLK _84866_/D _84866_/Q sky130_fd_sc_hd__dfxtp_4
X_86605_ _86610_/CLK _86605_/D _72368_/A sky130_fd_sc_hd__dfxtp_4
X_71831_ _71829_/X _71839_/B _70768_/A _71826_/X _71831_/X sky130_fd_sc_hd__and4_4
X_83817_ _83842_/CLK _83817_/D _74807_/A sky130_fd_sc_hd__dfxtp_4
X_59553_ _59552_/Y _59661_/D sky130_fd_sc_hd__inv_2
X_56765_ _56765_/A _56753_/Y _56764_/Y _56765_/Y sky130_fd_sc_hd__nand3_4
X_41991_ _41990_/Y _41991_/Y sky130_fd_sc_hd__inv_2
X_87585_ _88108_/CLK _87585_/D _73989_/A sky130_fd_sc_hd__dfxtp_4
X_53977_ _85530_/Q _53955_/X _53976_/Y _53977_/Y sky130_fd_sc_hd__o21ai_4
X_84797_ _84797_/CLK _84797_/D _84797_/Q sky130_fd_sc_hd__dfxtp_4
X_58504_ _83424_/Q _58504_/Y sky130_fd_sc_hd__inv_2
X_43730_ _43729_/X _43730_/Y sky130_fd_sc_hd__inv_2
X_55716_ _56454_/C _55126_/A _55128_/A _55715_/X _55716_/X sky130_fd_sc_hd__a211o_4
X_74550_ _74549_/Y _74625_/A sky130_fd_sc_hd__buf_2
X_86536_ _86210_/CLK _48318_/Y _86536_/Q sky130_fd_sc_hd__dfxtp_4
X_40942_ _40756_/A _40942_/X sky130_fd_sc_hd__buf_2
X_52928_ _52925_/Y _52920_/X _52927_/X _85729_/D sky130_fd_sc_hd__a21oi_4
X_59484_ _59484_/A _59484_/Y sky130_fd_sc_hd__inv_2
X_71762_ _71761_/Y _71762_/X sky130_fd_sc_hd__buf_2
X_83748_ _83749_/CLK _83748_/D _83748_/Q sky130_fd_sc_hd__dfxtp_4
X_56696_ _56696_/A _56696_/B _56696_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_496_0_CLK clkbuf_9_248_0_CLK/X _86384_/CLK sky130_fd_sc_hd__clkbuf_1
X_73501_ _73163_/X _83052_/Q _73385_/X _73500_/X _73501_/X sky130_fd_sc_hd__a211o_4
X_70713_ _70848_/A _70713_/X sky130_fd_sc_hd__buf_2
X_58435_ _58423_/X _83481_/Q _58434_/Y _84849_/D sky130_fd_sc_hd__o21a_4
X_55647_ _56650_/B _55467_/X _55646_/X _55503_/D _55647_/X sky130_fd_sc_hd__and4_4
X_43661_ _43611_/A _43661_/X sky130_fd_sc_hd__buf_2
X_74481_ _83057_/Q _74474_/X _74480_/Y _74481_/Y sky130_fd_sc_hd__o21ai_4
X_86467_ _83311_/CLK _86467_/D _86467_/Q sky130_fd_sc_hd__dfxtp_4
X_40873_ _40857_/X _41048_/A _40872_/X _40873_/X sky130_fd_sc_hd__o21a_4
X_52859_ _52850_/A _52859_/B _52859_/Y sky130_fd_sc_hd__nand2_4
X_83679_ _86104_/CLK _70868_/Y _83679_/Q sky130_fd_sc_hd__dfxtp_4
X_71693_ _71626_/A _71690_/A _71874_/D _71693_/Y sky130_fd_sc_hd__nor3_4
X_45400_ _45392_/X _45399_/X _45361_/X _45400_/X sky130_fd_sc_hd__a21o_4
X_76220_ _76217_/X _76221_/C _76219_/Y _76220_/Y sky130_fd_sc_hd__a21oi_4
X_88206_ _87950_/CLK _88206_/D _66694_/B sky130_fd_sc_hd__dfxtp_4
X_42612_ _42612_/A _42612_/X sky130_fd_sc_hd__buf_2
X_73432_ _48647_/Y _73432_/B _73432_/X sky130_fd_sc_hd__xor2_4
X_85418_ _85643_/CLK _54572_/Y _85418_/Q sky130_fd_sc_hd__dfxtp_4
X_46380_ _46380_/A _46380_/B _46380_/X sky130_fd_sc_hd__or2_4
X_70644_ _53017_/B _70632_/X _70643_/Y _83736_/D sky130_fd_sc_hd__o21ai_4
X_58366_ _58328_/A _58366_/X sky130_fd_sc_hd__buf_2
X_43592_ _43605_/A _43611_/A sky130_fd_sc_hd__buf_2
X_55578_ _44081_/X _85148_/Q _55578_/X sky130_fd_sc_hd__and2_4
X_86398_ _86398_/CLK _86398_/D _86398_/Q sky130_fd_sc_hd__dfxtp_4
X_45331_ _45331_/A _45331_/Y sky130_fd_sc_hd__inv_2
X_57317_ _57317_/A _57317_/Y sky130_fd_sc_hd__inv_2
X_76151_ _76150_/A _76150_/B _81537_/Q _76151_/Y sky130_fd_sc_hd__a21oi_4
X_88137_ _88398_/CLK _41818_/Y _88137_/Q sky130_fd_sc_hd__dfxtp_4
X_42543_ _72728_/A _42543_/Y sky130_fd_sc_hd__inv_2
X_54529_ _85425_/Q _54512_/X _54528_/Y _54529_/Y sky130_fd_sc_hd__o21ai_4
X_73363_ _48615_/A _73363_/B _73363_/X sky130_fd_sc_hd__xor2_4
X_85349_ _85957_/CLK _54943_/Y _85349_/Q sky130_fd_sc_hd__dfxtp_4
X_70575_ HASH_ADDR[4] _70933_/B sky130_fd_sc_hd__inv_2
X_58297_ _58282_/X _58294_/Y _58296_/Y _84885_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_4_11_1_CLK clkbuf_4_11_0_CLK/X clkbuf_5_23_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_75102_ _75102_/A _75102_/B _75104_/A sky130_fd_sc_hd__nand2_4
X_72314_ _72287_/X _85329_/Q _72225_/X _72314_/X sky130_fd_sc_hd__o21a_4
X_48050_ _48731_/A _48092_/A sky130_fd_sc_hd__buf_2
X_45262_ _45255_/X _45259_/Y _45261_/Y _45262_/Y sky130_fd_sc_hd__a21oi_4
X_76082_ _76082_/A _76081_/Y _76083_/B sky130_fd_sc_hd__xor2_4
X_57248_ _57327_/B _57340_/C sky130_fd_sc_hd__buf_2
X_88068_ _87820_/CLK _42021_/Y _88068_/Q sky130_fd_sc_hd__dfxtp_4
X_42474_ _42460_/X _42472_/X _40617_/X _68520_/B _42463_/X _42474_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73294_ _73292_/X _73293_/Y _73221_/X _73294_/Y sky130_fd_sc_hd__a21oi_4
X_47001_ _46996_/Y _46987_/X _47000_/X _86681_/D sky130_fd_sc_hd__a21oi_4
X_44213_ _57019_/A _44213_/X sky130_fd_sc_hd__buf_2
X_79910_ _84923_/Q _84171_/Q _79912_/A sky130_fd_sc_hd__nor2_4
X_75033_ _81147_/D _75032_/B _75033_/Y sky130_fd_sc_hd__nor2_4
X_87019_ _88301_/CLK _44645_/X _87019_/Q sky130_fd_sc_hd__dfxtp_4
X_41425_ _41399_/X _41400_/X _41424_/X _88218_/Q _41388_/X _41425_/Y
+ sky130_fd_sc_hd__o32ai_4
X_72245_ _72220_/A _86295_/Q _72245_/Y sky130_fd_sc_hd__nor2_4
X_45193_ _45193_/A _45709_/A sky130_fd_sc_hd__buf_2
X_57179_ _57179_/A _57179_/B _57179_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_434_0_CLK clkbuf_9_217_0_CLK/X _84228_/CLK sky130_fd_sc_hd__clkbuf_1
X_44144_ _44160_/A _87186_/Q _44144_/Y sky130_fd_sc_hd__nand2_4
X_79841_ _79828_/Y _79832_/Y _79840_/X _79842_/B sky130_fd_sc_hd__o21ai_4
X_41356_ _41355_/Y _41356_/X sky130_fd_sc_hd__buf_2
X_60190_ _60189_/Y _60324_/B sky130_fd_sc_hd__buf_2
X_72176_ _72176_/A _72176_/X sky130_fd_sc_hd__buf_2
X_71127_ _71129_/A _71082_/B _71119_/C _71127_/Y sky130_fd_sc_hd__nand3_4
X_48952_ _48612_/A _48952_/X sky130_fd_sc_hd__buf_2
X_44075_ _55741_/A _55159_/A sky130_fd_sc_hd__buf_2
X_79772_ _84222_/Q _83270_/Q _79772_/Y sky130_fd_sc_hd__nand2_4
X_41287_ _41255_/X _82913_/Q _41286_/X _41287_/Y sky130_fd_sc_hd__o21ai_4
X_76984_ _84536_/Q _76984_/B _76984_/X sky130_fd_sc_hd__xor2_4
X_47903_ _47846_/A _47903_/X sky130_fd_sc_hd__buf_2
X_43026_ _42439_/X _43017_/X _40573_/X _73577_/A _43025_/X _43027_/A
+ sky130_fd_sc_hd__o32ai_4
X_78723_ _78700_/Y _78706_/B _78723_/Y sky130_fd_sc_hd__nor2_4
X_71058_ _71058_/A _71080_/B _71055_/C _71058_/Y sky130_fd_sc_hd__nand3_4
X_75935_ _81699_/D _75927_/B _75935_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_449_0_CLK clkbuf_9_224_0_CLK/X _86303_/CLK sky130_fd_sc_hd__clkbuf_1
X_48883_ _48881_/X _81793_/Q _48882_/Y _48884_/A sky130_fd_sc_hd__o21ai_4
X_62900_ _62897_/Y _60337_/A _62650_/X _62898_/X _62899_/Y _62900_/X
+ sky130_fd_sc_hd__a41o_4
X_70009_ _70009_/A _70048_/A sky130_fd_sc_hd__buf_2
X_47834_ _47834_/A _57489_/B _47841_/A _47834_/Y sky130_fd_sc_hd__nand3_4
X_78654_ _78654_/A _78652_/Y _78654_/C _78655_/B sky130_fd_sc_hd__nand3_4
X_63880_ _63848_/X _63849_/X _84289_/Q _63880_/Y sky130_fd_sc_hd__nor3_4
X_75866_ _75863_/Y _75865_/Y _80992_/D sky130_fd_sc_hd__nor2_4
X_77605_ _77603_/X _77604_/Y _77605_/X sky130_fd_sc_hd__and2_4
X_74817_ _74817_/A _74817_/Y sky130_fd_sc_hd__inv_2
X_62831_ _62886_/A _62831_/X sky130_fd_sc_hd__buf_2
X_47765_ _86600_/Q _47760_/X _47764_/Y _47765_/Y sky130_fd_sc_hd__o21ai_4
X_78585_ _78586_/A _82677_/D _78585_/Y sky130_fd_sc_hd__nor2_4
X_44977_ _44975_/X _61375_/B _44907_/X _44977_/Y sky130_fd_sc_hd__o21ai_4
X_75797_ _75802_/B _75796_/Y _75800_/A sky130_fd_sc_hd__xor2_4
X_49504_ _49504_/A _49614_/A sky130_fd_sc_hd__buf_2
X_46716_ _54325_/D _46716_/X sky130_fd_sc_hd__buf_2
X_65550_ _65438_/X _86201_/Q _65182_/X _65549_/X _65550_/X sky130_fd_sc_hd__a211o_4
X_77536_ _77537_/A _77537_/B _77535_/Y _77540_/B sky130_fd_sc_hd__o21a_4
X_43928_ _43927_/X _43928_/X sky130_fd_sc_hd__buf_2
X_62762_ _62727_/A _62762_/B _61876_/X _62762_/Y sky130_fd_sc_hd__nand3_4
X_74748_ _74748_/A _70638_/A _74797_/C _74769_/D _74748_/Y sky130_fd_sc_hd__nand4_4
X_47696_ _47696_/A _53193_/B _47696_/Y sky130_fd_sc_hd__nand2_4
X_64501_ _61140_/X _64523_/B _58194_/A _64523_/D _64501_/X sky130_fd_sc_hd__and4_4
X_61713_ _61712_/X _62128_/B sky130_fd_sc_hd__buf_2
X_49435_ _49407_/A _49447_/A sky130_fd_sc_hd__buf_2
X_46647_ _46670_/A _46647_/B _46659_/C _51768_/D _46647_/X sky130_fd_sc_hd__and4_4
X_65481_ _65449_/A _65546_/B _65481_/C _65481_/X sky130_fd_sc_hd__and3_4
X_77467_ _77468_/A _77468_/B _77467_/Y sky130_fd_sc_hd__nor2_4
X_43859_ _43846_/X _43854_/X _41225_/X _68898_/B _43847_/X _43859_/Y
+ sky130_fd_sc_hd__o32ai_4
X_62693_ _62678_/A _62727_/B _61780_/X _62693_/Y sky130_fd_sc_hd__nand3_4
X_74679_ _74679_/A _74679_/B _74679_/Y sky130_fd_sc_hd__nand2_4
X_67220_ _67220_/A _67219_/X _67220_/Y sky130_fd_sc_hd__nand2_4
X_79206_ _79205_/C _79205_/B _79206_/Y sky130_fd_sc_hd__nand2_4
X_64432_ _63598_/A _64419_/B _64432_/Y sky130_fd_sc_hd__nor2_4
X_76418_ _76418_/A _76417_/Y _76418_/X sky130_fd_sc_hd__and2_4
X_49366_ _49382_/A _46625_/X _49366_/Y sky130_fd_sc_hd__nand2_4
X_61644_ _61348_/A _61645_/A sky130_fd_sc_hd__buf_2
X_46578_ _47904_/A _46578_/X sky130_fd_sc_hd__buf_2
X_77398_ _77386_/A _77398_/Y sky130_fd_sc_hd__inv_2
X_48317_ _50360_/A _48286_/X _48287_/C _48317_/X sky130_fd_sc_hd__and3_4
X_67151_ _67148_/X _67150_/X _67151_/Y sky130_fd_sc_hd__nand2_4
X_79137_ _79137_/A _61577_/C _79137_/X sky130_fd_sc_hd__xor2_4
X_45529_ _63100_/B _61430_/A sky130_fd_sc_hd__buf_2
X_64363_ _64363_/A _64363_/B _63524_/B _64318_/D _64363_/X sky130_fd_sc_hd__and4_4
X_76349_ _76348_/B _76348_/C _76344_/Y _76349_/Y sky130_fd_sc_hd__o21ai_4
X_61575_ _61568_/Y _61570_/Y _61525_/X _61572_/Y _61574_/Y _61575_/X
+ sky130_fd_sc_hd__a41o_4
X_49297_ _49273_/A _50816_/B _49297_/Y sky130_fd_sc_hd__nand2_4
X_66102_ _66040_/X _84980_/Q _66027_/X _66101_/X _66102_/X sky130_fd_sc_hd__a211o_4
X_63314_ _60433_/A _63314_/B _63333_/C _63240_/X _63314_/X sky130_fd_sc_hd__and4_4
X_48248_ _48245_/Y _48226_/X _48247_/Y _86549_/D sky130_fd_sc_hd__a21boi_4
X_60526_ _60526_/A _60526_/B _79146_/A _60526_/Y sky130_fd_sc_hd__nor3_4
X_67082_ _67082_/A _67133_/A sky130_fd_sc_hd__buf_2
X_79068_ _79055_/B _79055_/A _79044_/C _79044_/B _79067_/Y _79068_/X
+ sky130_fd_sc_hd__o41a_4
Xclkbuf_9_508_0_CLK clkbuf_9_509_0_CLK/A clkbuf_9_508_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_64294_ _64275_/A _64294_/B _64274_/X _64294_/X sky130_fd_sc_hd__and3_4
X_66033_ _65970_/A _66004_/B _84161_/Q _66033_/X sky130_fd_sc_hd__and3_4
X_78019_ _78018_/B _78018_/A _78021_/C sky130_fd_sc_hd__nand2_4
X_63245_ _63243_/Y _63244_/X _63231_/X _63245_/Y sky130_fd_sc_hd__a21oi_4
X_48179_ _48184_/A _48178_/X _48179_/Y sky130_fd_sc_hd__nand2_4
X_60457_ _60456_/X _60457_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_61_0_CLK clkbuf_8_61_0_CLK/A clkbuf_8_61_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_50210_ _50208_/Y _50191_/X _50209_/X _50210_/Y sky130_fd_sc_hd__a21oi_4
X_81030_ _81061_/CLK _81030_/D _81222_/D sky130_fd_sc_hd__dfxtp_4
X_51190_ _86057_/Q _51183_/X _51189_/Y _51190_/Y sky130_fd_sc_hd__o21ai_4
X_63176_ _63118_/A _63176_/X sky130_fd_sc_hd__buf_2
X_60388_ _60387_/X _60606_/A sky130_fd_sc_hd__buf_2
X_50141_ _50092_/A _50141_/X sky130_fd_sc_hd__buf_2
X_62127_ _61716_/X _61636_/B _62126_/X _62127_/X sky130_fd_sc_hd__a21o_4
X_67984_ _68651_/A _67984_/X sky130_fd_sc_hd__buf_2
X_69723_ _73083_/A _68640_/X _68070_/X _69722_/Y _69723_/X sky130_fd_sc_hd__a211o_4
X_50072_ _86270_/Q _50061_/X _50071_/Y _50072_/Y sky130_fd_sc_hd__o21ai_4
X_66935_ _69582_/A _66935_/X sky130_fd_sc_hd__buf_2
X_62058_ _61716_/X _61579_/B _62057_/X _62058_/X sky130_fd_sc_hd__a21o_4
X_82981_ _82987_/CLK _82981_/D _82981_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_76_0_CLK clkbuf_8_77_0_CLK/A clkbuf_8_76_0_CLK/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_7_8_0_CLK clkbuf_6_4_0_CLK/X clkbuf_7_8_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_53900_ _53900_/A _53929_/A sky130_fd_sc_hd__buf_2
X_61009_ _61004_/Y _61008_/Y _60938_/A _76990_/A _60898_/X _84542_/D
+ sky130_fd_sc_hd__o32a_4
X_84720_ _84727_/CLK _84720_/D _64225_/C sky130_fd_sc_hd__dfxtp_4
X_81932_ _83906_/CLK _77838_/Y _81932_/Q sky130_fd_sc_hd__dfxtp_4
X_69654_ _69654_/A _69655_/A sky130_fd_sc_hd__buf_2
X_54880_ _54885_/A _54880_/B _54880_/Y sky130_fd_sc_hd__nand2_4
X_66866_ _66862_/X _66865_/X _66843_/X _66866_/X sky130_fd_sc_hd__a21o_4
X_68605_ _87498_/Q _68504_/X _68601_/X _68604_/X _68605_/X sky130_fd_sc_hd__a211o_4
X_53831_ _53828_/Y _53829_/X _53830_/X _53831_/Y sky130_fd_sc_hd__a21oi_4
X_65817_ _65855_/A _65916_/B _65817_/C _65817_/X sky130_fd_sc_hd__and3_4
X_84651_ _84652_/CLK _60149_/X _79907_/B sky130_fd_sc_hd__dfxtp_4
X_81863_ _84375_/CLK _78054_/X _81863_/Q sky130_fd_sc_hd__dfxtp_4
X_69585_ _69581_/X _69584_/X _69570_/X _69585_/X sky130_fd_sc_hd__a21o_4
X_66797_ _69162_/A _66797_/X sky130_fd_sc_hd__buf_2
X_83602_ _85557_/CLK _71114_/Y _49115_/A sky130_fd_sc_hd__dfxtp_4
X_56550_ _72973_/B _56550_/X sky130_fd_sc_hd__buf_2
X_80814_ _80821_/CLK _83958_/Q _75829_/B sky130_fd_sc_hd__dfxtp_4
X_68536_ _87097_/Q _68455_/X _68509_/X _68535_/X _68536_/X sky130_fd_sc_hd__a211o_4
X_87370_ _87373_/CLK _87370_/D _87370_/Q sky130_fd_sc_hd__dfxtp_4
X_53762_ _85573_/Q _53754_/X _53761_/Y _53762_/Y sky130_fd_sc_hd__o21ai_4
X_65748_ _65731_/A _85868_/Q _65748_/X sky130_fd_sc_hd__and2_4
X_84582_ _84590_/CLK _60706_/Y _84582_/Q sky130_fd_sc_hd__dfxtp_4
X_50974_ _50973_/X _50963_/B _50963_/C _46775_/X _50974_/X sky130_fd_sc_hd__and4_4
X_81794_ _81794_/CLK _81602_/Q _81794_/Q sky130_fd_sc_hd__dfxtp_4
X_55501_ _55501_/A _55500_/X _55501_/X sky130_fd_sc_hd__and2_4
X_86321_ _86640_/CLK _86321_/D _57952_/B sky130_fd_sc_hd__dfxtp_4
X_52713_ _52718_/A _52713_/B _52713_/Y sky130_fd_sc_hd__nand2_4
X_83533_ _86213_/CLK _83533_/D _83533_/Q sky130_fd_sc_hd__dfxtp_4
X_56481_ _56474_/X _56472_/B _55931_/B _56481_/Y sky130_fd_sc_hd__nand3_4
X_80745_ _80962_/CLK _75183_/X _81153_/D sky130_fd_sc_hd__dfxtp_4
X_68467_ _68384_/A _68467_/X sky130_fd_sc_hd__buf_2
X_53693_ _53690_/Y _53680_/X _53692_/X _85587_/D sky130_fd_sc_hd__a21oi_4
X_65679_ _65533_/X _65676_/Y _65678_/Y _65679_/Y sky130_fd_sc_hd__o21ai_4
X_58220_ _83400_/Q _58220_/Y sky130_fd_sc_hd__inv_2
X_55432_ _56777_/A _55405_/X _55411_/Y _55432_/Y sky130_fd_sc_hd__a21boi_4
X_67418_ _87408_/Q _67394_/X _67344_/X _67417_/X _67418_/X sky130_fd_sc_hd__a211o_4
X_86252_ _85554_/CLK _86252_/D _86252_/Q sky130_fd_sc_hd__dfxtp_4
X_52644_ _52642_/Y _52619_/X _52643_/X _85781_/D sky130_fd_sc_hd__a21oi_4
X_83464_ _83464_/CLK _83464_/D _83464_/Q sky130_fd_sc_hd__dfxtp_4
X_80676_ _80676_/CLK _80676_/D _80676_/Q sky130_fd_sc_hd__dfxtp_4
X_68398_ _87006_/Q _68394_/X _44246_/A _68397_/X _68398_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_8_14_0_CLK clkbuf_7_7_0_CLK/X clkbuf_9_29_0_CLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_504 sky130_fd_sc_hd__decap_3
X_85203_ _85168_/CLK _85203_/D _56414_/C sky130_fd_sc_hd__dfxtp_4
X_58151_ _58151_/A _58151_/B _58151_/Y sky130_fd_sc_hd__nor2_4
XPHY_515 sky130_fd_sc_hd__decap_3
X_82415_ _82828_/CLK _82447_/Q _78489_/A sky130_fd_sc_hd__dfxtp_4
X_55363_ _55329_/Y _55363_/B _55330_/X _56708_/C sky130_fd_sc_hd__nand3_4
X_67349_ _67324_/A _67349_/B _67349_/X sky130_fd_sc_hd__and2_4
X_86183_ _86505_/CLK _86183_/D _86183_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_526 sky130_fd_sc_hd__decap_3
X_52575_ _52515_/X _52575_/X sky130_fd_sc_hd__buf_2
X_83395_ _83756_/CLK _71732_/Y _58240_/A sky130_fd_sc_hd__dfxtp_4
XPHY_537 sky130_fd_sc_hd__decap_3
XPHY_548 sky130_fd_sc_hd__decap_3
X_57102_ _57097_/X _56578_/X _85086_/Q _57099_/X _85086_/D sky130_fd_sc_hd__a2bb2o_4
X_54314_ _54314_/A _54314_/B _54314_/Y sky130_fd_sc_hd__nand2_4
XPHY_559 sky130_fd_sc_hd__decap_3
X_85134_ _85134_/CLK _56765_/Y _85134_/Q sky130_fd_sc_hd__dfxtp_4
X_51526_ _51552_/A _51533_/C sky130_fd_sc_hd__buf_2
X_58082_ _86630_/Q _58136_/B _58082_/Y sky130_fd_sc_hd__nor2_4
X_70360_ _70827_/C _70358_/X _70907_/B _70361_/A sky130_fd_sc_hd__nand3_4
X_82346_ _86753_/CLK _82346_/D _48077_/A sky130_fd_sc_hd__dfxtp_4
X_55294_ _55293_/X _55162_/Y _55417_/A sky130_fd_sc_hd__and2_4
X_57033_ _56787_/X _56994_/D _56732_/X _56788_/X _56821_/X _57034_/C
+ sky130_fd_sc_hd__a41o_4
X_69019_ _68907_/X _68882_/X _69006_/Y _69018_/Y _69019_/X sky130_fd_sc_hd__a211o_4
X_54245_ _54245_/A _54329_/A sky130_fd_sc_hd__buf_2
X_85065_ _84998_/CLK _57195_/Y _85065_/Q sky130_fd_sc_hd__dfxtp_4
X_51457_ _51455_/Y _51448_/X _51456_/X _51457_/Y sky130_fd_sc_hd__a21oi_4
X_70291_ _70289_/X _74809_/A _70290_/X _83809_/D sky130_fd_sc_hd__a21o_4
Xclkbuf_8_29_0_CLK clkbuf_8_29_0_CLK/A clkbuf_9_59_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_82277_ _82339_/CLK _82277_/D _40912_/B sky130_fd_sc_hd__dfxtp_4
X_41210_ _41205_/X _41206_/X _41209_/X _68820_/B _41194_/X _41210_/Y
+ sky130_fd_sc_hd__o32ai_4
X_72030_ _72028_/Y _72009_/X _72029_/Y _83299_/D sky130_fd_sc_hd__a21boi_4
X_84016_ _84014_/CLK _84016_/D _84016_/Q sky130_fd_sc_hd__dfxtp_4
X_50408_ _48388_/A _50430_/B _50435_/C _50408_/X sky130_fd_sc_hd__and3_4
X_81228_ _81227_/CLK _81036_/Q _81228_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_3_0_1_CLK clkbuf_3_0_1_CLK/A clkbuf_3_0_1_CLK/X sky130_fd_sc_hd__clkbuf_1
X_42190_ _41282_/X _42183_/X _87988_/Q _42184_/X _87988_/D sky130_fd_sc_hd__a2bb2o_4
X_54176_ _85490_/Q _54167_/X _54175_/Y _54176_/Y sky130_fd_sc_hd__o21ai_4
X_51388_ _51790_/A _51758_/A sky130_fd_sc_hd__buf_2
X_41141_ _41141_/A _41141_/Y sky130_fd_sc_hd__inv_2
X_53127_ _53121_/X _53127_/B _53127_/Y sky130_fd_sc_hd__nand2_4
X_50339_ _52039_/A _50331_/B _50338_/X _50339_/X sky130_fd_sc_hd__and3_4
X_81159_ _81160_/CLK _74879_/B _81159_/Q sky130_fd_sc_hd__dfxtp_4
X_58984_ _58984_/A _58988_/B sky130_fd_sc_hd__buf_2
X_53058_ _53074_/A _53063_/B _53058_/C _53058_/D _53058_/X sky130_fd_sc_hd__and4_4
X_57935_ _86642_/Q _57845_/X _57935_/Y sky130_fd_sc_hd__nor2_4
X_41072_ _47825_/A _41072_/X sky130_fd_sc_hd__buf_2
X_73981_ _73979_/X _73967_/X _73981_/C _73981_/Y sky130_fd_sc_hd__nand3_4
X_85967_ _85679_/CLK _85967_/D _85967_/Q sky130_fd_sc_hd__dfxtp_4
X_52009_ _51947_/A _50306_/B _52009_/Y sky130_fd_sc_hd__nand2_4
X_44900_ _44904_/A _45819_/A sky130_fd_sc_hd__buf_2
X_75720_ _75708_/A _75707_/Y _75694_/A _75719_/Y _75720_/X sky130_fd_sc_hd__a2bb2o_4
X_87706_ _87446_/CLK _87706_/D _87706_/Q sky130_fd_sc_hd__dfxtp_4
X_72932_ _73093_/A _65521_/B _72932_/X sky130_fd_sc_hd__and2_4
X_84918_ _84905_/CLK _58161_/X _84918_/Q sky130_fd_sc_hd__dfxtp_4
X_45880_ _45873_/X _45877_/Y _45879_/Y _45880_/Y sky130_fd_sc_hd__a21oi_4
X_57866_ _57866_/A _58827_/A sky130_fd_sc_hd__buf_2
X_85898_ _84970_/CLK _85898_/D _74104_/B sky130_fd_sc_hd__dfxtp_4
X_59605_ _59604_/X _59605_/Y sky130_fd_sc_hd__inv_2
X_44831_ _41700_/Y _44817_/X _67654_/B _44818_/X _44831_/X sky130_fd_sc_hd__a2bb2o_4
X_56817_ _56816_/Y _56713_/A _56817_/X sky130_fd_sc_hd__xor2_4
X_75651_ _75649_/Y _75650_/Y _75659_/B sky130_fd_sc_hd__xor2_4
X_87637_ _87636_/CLK _87637_/D _68051_/B sky130_fd_sc_hd__dfxtp_4
X_72863_ _72856_/X _72860_/X _72862_/X _72869_/A sky130_fd_sc_hd__a21o_4
X_84849_ _84849_/CLK _84849_/D _84849_/Q sky130_fd_sc_hd__dfxtp_4
X_57797_ _57753_/Y _57758_/X _57780_/X _57796_/X _84949_/D sky130_fd_sc_hd__a22oi_4
X_74602_ _45232_/A _74598_/X _74601_/X _74602_/Y sky130_fd_sc_hd__o21ai_4
X_47550_ _47546_/Y _47509_/X _47549_/X _47550_/Y sky130_fd_sc_hd__a21oi_4
X_71814_ _71805_/X _83366_/Q _71813_/X _83366_/D sky130_fd_sc_hd__a21o_4
X_59536_ _59536_/A _60175_/A _59716_/B _61285_/C _59537_/A sky130_fd_sc_hd__nand4_4
X_78370_ _78370_/A _82758_/D _82470_/D sky130_fd_sc_hd__xor2_4
X_44762_ _44762_/A _44762_/Y sky130_fd_sc_hd__inv_2
X_56748_ _56721_/Y _56750_/B sky130_fd_sc_hd__inv_2
X_75582_ _75888_/A _75580_/Y _75584_/C _75583_/A sky130_fd_sc_hd__a21oi_4
X_87568_ _86534_/CLK _43120_/Y _87568_/Q sky130_fd_sc_hd__dfxtp_4
X_41974_ _41965_/X _41956_/X _40749_/X _41973_/Y _41967_/X _41974_/Y
+ sky130_fd_sc_hd__o32ai_4
X_72794_ _72943_/A _72794_/X sky130_fd_sc_hd__buf_2
X_46501_ _46500_/Y _51350_/B sky130_fd_sc_hd__buf_2
X_77321_ _77317_/X _77320_/Y _82184_/D sky130_fd_sc_hd__xor2_4
X_43713_ _43713_/A _69793_/B sky130_fd_sc_hd__inv_2
X_74533_ _74533_/A _74531_/B _74531_/C _74533_/D _74533_/Y sky130_fd_sc_hd__nand4_4
X_86519_ _86516_/CLK _48477_/Y _65584_/B sky130_fd_sc_hd__dfxtp_4
X_40925_ _40924_/Y _40925_/X sky130_fd_sc_hd__buf_2
X_47481_ _47481_/A _53072_/B sky130_fd_sc_hd__buf_2
X_71745_ _52931_/B _71737_/X _71744_/Y _83392_/D sky130_fd_sc_hd__o21ai_4
X_59467_ _84724_/Q _59467_/Y sky130_fd_sc_hd__inv_2
X_44693_ _44679_/X _44680_/X _40641_/X _86998_/Q _44681_/X _44694_/A
+ sky130_fd_sc_hd__o32ai_4
X_56679_ _56674_/X _56679_/B _57140_/B _83336_/Q _56680_/A sky130_fd_sc_hd__and4_4
X_87499_ _87757_/CLK _87499_/D _87499_/Q sky130_fd_sc_hd__dfxtp_4
X_49220_ _49220_/A _53953_/B _49220_/Y sky130_fd_sc_hd__nand2_4
X_46432_ _83641_/Q _46433_/A sky130_fd_sc_hd__inv_2
X_58418_ _58418_/A _58415_/B _58418_/Y sky130_fd_sc_hd__nand2_4
X_77252_ _77252_/A _77254_/A _77253_/A _77252_/Y sky130_fd_sc_hd__nand3_4
X_43644_ _87329_/Q _43644_/Y sky130_fd_sc_hd__inv_2
X_74464_ _48589_/A _74478_/B _74478_/C _74464_/X sky130_fd_sc_hd__and3_4
X_40856_ _40855_/Y _88322_/D sky130_fd_sc_hd__inv_2
X_71676_ _71680_/A _71671_/X _70472_/X _71676_/Y sky130_fd_sc_hd__nand3_4
X_59398_ _59398_/A _59399_/B sky130_fd_sc_hd__buf_2
X_76203_ _76200_/X _81638_/Q _76201_/Y _76219_/A sky130_fd_sc_hd__nand3_4
X_49151_ _49080_/A _50183_/B _49151_/X sky130_fd_sc_hd__and2_4
X_73415_ _73415_/A _73053_/B _73415_/Y sky130_fd_sc_hd__nor2_4
X_46363_ _46358_/Y _46346_/X _46362_/Y _86744_/D sky130_fd_sc_hd__a21boi_4
X_70627_ _70627_/A _71115_/D sky130_fd_sc_hd__buf_2
X_58349_ _58328_/X _83768_/Q _58348_/Y _58349_/X sky130_fd_sc_hd__o21a_4
X_77183_ _82012_/Q _82300_/D _77202_/A sky130_fd_sc_hd__xor2_4
X_43575_ _40528_/X _53455_/A _87352_/Q _43185_/A _87352_/D sky130_fd_sc_hd__a2bb2o_4
X_74395_ _74453_/A _74395_/X sky130_fd_sc_hd__buf_2
X_40787_ _40787_/A _40787_/X sky130_fd_sc_hd__buf_2
X_48102_ _47838_/X _48781_/A sky130_fd_sc_hd__buf_2
X_45314_ _56536_/C _45284_/X _45265_/X _45314_/X sky130_fd_sc_hd__o21a_4
X_76134_ _76129_/B _76132_/X _76133_/Y _76134_/Y sky130_fd_sc_hd__a21boi_4
X_42526_ _42517_/X _42501_/X _40729_/X _42525_/Y _42519_/X _87834_/D
+ sky130_fd_sc_hd__o32ai_4
X_49082_ _49082_/A _49083_/A sky130_fd_sc_hd__inv_2
X_61360_ _61359_/Y _61360_/Y sky130_fd_sc_hd__inv_2
X_73346_ _42041_/Y _73298_/X _73344_/X _73345_/Y _73346_/X sky130_fd_sc_hd__a211o_4
X_46294_ _46294_/A _46295_/A sky130_fd_sc_hd__inv_2
X_70558_ _71883_/A _70558_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_373_0_CLK clkbuf_9_186_0_CLK/X _85751_/CLK sky130_fd_sc_hd__clkbuf_1
X_48033_ _66183_/B _47998_/X _48032_/Y _48033_/Y sky130_fd_sc_hd__o21ai_4
X_60311_ _79755_/A _59822_/X _60300_/Y _60310_/X _84637_/D sky130_fd_sc_hd__o22a_4
X_45245_ _45244_/Y _45199_/B _45245_/Y sky130_fd_sc_hd__nand2_4
X_76065_ _76063_/B _81716_/D _76058_/B _76065_/Y sky130_fd_sc_hd__nand3_4
X_42457_ _42456_/Y _87858_/D sky130_fd_sc_hd__inv_2
X_61291_ _61290_/X _61292_/A sky130_fd_sc_hd__buf_2
X_73277_ _73274_/X _73276_/X _73200_/X _73277_/X sky130_fd_sc_hd__a21o_4
X_70489_ _71323_/A _71500_/C _71779_/B _70489_/Y sky130_fd_sc_hd__nand3_4
X_63030_ _60476_/A _63030_/B _63030_/C _60541_/C _63030_/X sky130_fd_sc_hd__and4_4
X_75016_ _81146_/D _75016_/B _75016_/Y sky130_fd_sc_hd__nand2_4
X_41408_ _41407_/X _41408_/X sky130_fd_sc_hd__buf_2
X_72228_ _59085_/A _72228_/X sky130_fd_sc_hd__buf_2
X_60242_ _60036_/A _60525_/A sky130_fd_sc_hd__buf_2
X_45176_ _45252_/A _45176_/X sky130_fd_sc_hd__buf_2
X_42388_ _42373_/X _42388_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_494_0_CLK clkbuf_9_495_0_CLK/A clkbuf_9_494_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_44127_ _44126_/X _44127_/X sky130_fd_sc_hd__buf_2
X_79824_ _79816_/X _79817_/X _79823_/Y _79840_/A sky130_fd_sc_hd__a21boi_4
X_41339_ _41686_/B _41275_/B _41339_/X sky130_fd_sc_hd__or2_4
X_60173_ _60406_/B _72625_/A sky130_fd_sc_hd__buf_2
X_72159_ _72154_/Y _72158_/Y _59297_/X _72159_/X sky130_fd_sc_hd__a21o_4
X_49984_ _49995_/A _49973_/B _50005_/C _53196_/D _49984_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_388_0_CLK clkbuf_9_194_0_CLK/X _84350_/CLK sky130_fd_sc_hd__clkbuf_1
X_48935_ _48985_/A _48935_/X sky130_fd_sc_hd__buf_2
X_44058_ _44058_/A _44059_/A sky130_fd_sc_hd__buf_2
X_79755_ _79755_/A _79755_/B _79761_/B sky130_fd_sc_hd__xor2_4
X_64981_ _65319_/A _86419_/Q _64981_/X sky130_fd_sc_hd__and2_4
X_76967_ _81684_/Q _76967_/B _76967_/Y sky130_fd_sc_hd__xnor2_4
X_43009_ _40538_/X _51934_/A _67259_/B _42634_/A _87606_/D sky130_fd_sc_hd__a2bb2o_4
X_78706_ _78700_/Y _78706_/B _82780_/D sky130_fd_sc_hd__xor2_4
X_66720_ _66720_/A _66719_/X _66720_/Y sky130_fd_sc_hd__nand2_4
X_63932_ _63749_/A _63947_/B sky130_fd_sc_hd__buf_2
X_75918_ _61165_/C _75918_/B _75918_/X sky130_fd_sc_hd__xor2_4
X_48866_ _48691_/A _48859_/B _48854_/C _48866_/X sky130_fd_sc_hd__and3_4
X_79686_ _79683_/Y _79666_/Y _79685_/X _79686_/Y sky130_fd_sc_hd__o21ai_4
X_76898_ _76897_/Y _76899_/B sky130_fd_sc_hd__inv_2
Xclkbuf_10_311_0_CLK clkbuf_9_155_0_CLK/X _85489_/CLK sky130_fd_sc_hd__clkbuf_1
X_47817_ _47817_/A _47818_/A sky130_fd_sc_hd__inv_2
X_66651_ _66651_/A _66651_/B _66651_/X sky130_fd_sc_hd__and2_4
X_78637_ _78632_/X _78637_/B _78637_/C _78638_/B sky130_fd_sc_hd__nand3_4
X_63863_ _63859_/X _63810_/X _63860_/Y _63861_/Y _63862_/X _63863_/X
+ sky130_fd_sc_hd__a41o_4
X_75849_ _75846_/A _81023_/Q _75849_/Y sky130_fd_sc_hd__nand2_4
X_48797_ _52182_/A _48829_/B _48814_/C _48797_/X sky130_fd_sc_hd__and3_4
Xclkbuf_10_941_0_CLK clkbuf_9_470_0_CLK/X _87542_/CLK sky130_fd_sc_hd__clkbuf_1
X_65602_ _65529_/A _65602_/X sky130_fd_sc_hd__buf_2
X_62814_ _62789_/A _63161_/A _62848_/C _62789_/D _62814_/X sky130_fd_sc_hd__and4_4
X_69370_ _88034_/Q _69368_/X _69232_/X _69369_/X _69370_/X sky130_fd_sc_hd__a211o_4
X_47748_ _55083_/D _53223_/D sky130_fd_sc_hd__buf_2
X_66582_ _68474_/A _66683_/A sky130_fd_sc_hd__buf_2
X_78568_ _78568_/A _78569_/C sky130_fd_sc_hd__inv_2
X_63794_ _63787_/Y _63789_/Y _63791_/Y _63794_/D _63794_/X sky130_fd_sc_hd__and4_4
Xclkbuf_9_432_0_CLK clkbuf_8_216_0_CLK/X clkbuf_9_432_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_68321_ _68319_/X _67961_/Y _68308_/X _68320_/Y _68321_/X sky130_fd_sc_hd__a211o_4
X_65533_ _65198_/A _65533_/X sky130_fd_sc_hd__buf_2
X_77519_ _77519_/A _77518_/X _77520_/B sky130_fd_sc_hd__xor2_4
X_62745_ _62731_/A _58177_/Y _62744_/X _62717_/X _62745_/X sky130_fd_sc_hd__and4_4
X_47679_ _47679_/A _53183_/B sky130_fd_sc_hd__buf_2
X_78499_ _78499_/A _78498_/Y _82767_/D sky130_fd_sc_hd__xor2_4
Xclkbuf_10_326_0_CLK clkbuf_9_163_0_CLK/X _86340_/CLK sky130_fd_sc_hd__clkbuf_1
X_49418_ _49418_/A _51800_/B _49418_/Y sky130_fd_sc_hd__nand2_4
X_80530_ _80530_/A _80513_/A _80530_/X sky130_fd_sc_hd__and2_4
X_68252_ _68246_/X _67555_/Y _68247_/X _68251_/Y _68252_/X sky130_fd_sc_hd__a211o_4
X_65464_ _65464_/A _65929_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_956_0_CLK clkbuf_9_478_0_CLK/X _86534_/CLK sky130_fd_sc_hd__clkbuf_1
X_50690_ _50682_/A _49135_/X _50690_/Y sky130_fd_sc_hd__nand2_4
X_62676_ _62658_/A _64236_/C _62676_/C _62657_/X _62676_/X sky130_fd_sc_hd__and4_4
X_67203_ _68389_/A _67203_/X sky130_fd_sc_hd__buf_2
X_64415_ _64410_/Y _64411_/X _64412_/X _64414_/Y _64384_/X _64415_/X
+ sky130_fd_sc_hd__o41a_4
X_49349_ _65367_/B _49334_/X _49348_/Y _49349_/Y sky130_fd_sc_hd__o21ai_4
X_61627_ _61636_/A _61627_/B _61590_/C _61627_/Y sky130_fd_sc_hd__nand3_4
X_80461_ _84761_/Q _84153_/Q _80461_/Y sky130_fd_sc_hd__nand2_4
X_68183_ _84018_/Q _68180_/X _68182_/X _68183_/X sky130_fd_sc_hd__a21bo_4
X_65395_ _65395_/A _65394_/Y _65395_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_447_0_CLK clkbuf_9_446_0_CLK/A clkbuf_9_447_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_82200_ _83681_/CLK _82200_/D _82392_/D sky130_fd_sc_hd__dfxtp_4
X_67134_ _87356_/Q _67035_/X _67106_/X _67133_/X _67134_/X sky130_fd_sc_hd__a211o_4
X_52360_ _52385_/A _49079_/A _52360_/X sky130_fd_sc_hd__and2_4
X_64346_ _64336_/A _58546_/A _64323_/X _64346_/Y sky130_fd_sc_hd__nand3_4
X_83180_ _83820_/CLK _83180_/D _83180_/Q sky130_fd_sc_hd__dfxtp_4
X_61558_ _61558_/A _61558_/B _61538_/C _61558_/Y sky130_fd_sc_hd__nand3_4
X_80392_ _80390_/X _80391_/X _80406_/A sky130_fd_sc_hd__xnor2_4
X_51311_ _51310_/X _50799_/B _51311_/Y sky130_fd_sc_hd__nand2_4
X_82131_ _82131_/CLK _82131_/D _77294_/B sky130_fd_sc_hd__dfxtp_4
X_60509_ _61287_/A _60509_/Y sky130_fd_sc_hd__inv_2
X_67065_ _88383_/Q _66988_/X _67040_/X _67064_/X _67065_/X sky130_fd_sc_hd__a211o_4
X_52291_ _52291_/A _52267_/B _52291_/C _52291_/X sky130_fd_sc_hd__and3_4
X_64277_ _64287_/A _84852_/Q _64287_/C _64277_/Y sky130_fd_sc_hd__nand3_4
X_61489_ _61437_/A _61489_/B _61459_/X _61489_/Y sky130_fd_sc_hd__nand3_4
X_54030_ _53929_/A _54031_/A sky130_fd_sc_hd__buf_2
X_66016_ _84162_/Q _66016_/Y sky130_fd_sc_hd__inv_2
X_51242_ _51242_/A _46267_/A _51242_/X sky130_fd_sc_hd__and2_4
X_63228_ _63223_/Y _63225_/X _63226_/X _63227_/X _63183_/X _63228_/Y
+ sky130_fd_sc_hd__o41ai_4
X_82062_ _84105_/CLK _82062_/D _77832_/A sky130_fd_sc_hd__dfxtp_4
X_81013_ _84150_/CLK _84221_/Q _81013_/Q sky130_fd_sc_hd__dfxtp_4
X_51173_ _51167_/A _52863_/B _51173_/Y sky130_fd_sc_hd__nand2_4
X_63159_ _63153_/Y _63155_/X _63156_/X _63158_/X _63125_/X _63159_/Y
+ sky130_fd_sc_hd__o41ai_4
X_86870_ _86873_/CLK _45546_/Y _63110_/B sky130_fd_sc_hd__dfxtp_4
X_50124_ _50120_/A _49025_/X _50124_/Y sky130_fd_sc_hd__nand2_4
X_85821_ _86045_/CLK _85821_/D _64694_/B sky130_fd_sc_hd__dfxtp_4
X_55981_ _55698_/A _85312_/Q _55981_/X sky130_fd_sc_hd__and2_4
X_67967_ _67992_/A _88153_/Q _67967_/X sky130_fd_sc_hd__and2_4
Xclkbuf_5_11_0_CLK clkbuf_4_5_1_CLK/X clkbuf_6_23_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_57720_ _84953_/Q _57691_/X _57704_/X _57719_/X _84953_/D sky130_fd_sc_hd__a2bb2oi_4
X_69706_ _69281_/Y _69644_/X _69672_/X _69705_/Y _69706_/X sky130_fd_sc_hd__a211o_4
X_50055_ _50053_/Y _48865_/X _50054_/X _86273_/D sky130_fd_sc_hd__a21oi_4
X_54932_ _54932_/A _54942_/B _54932_/C _53238_/D _54932_/X sky130_fd_sc_hd__and4_4
X_66918_ _66913_/X _66917_/X _66843_/X _66918_/X sky130_fd_sc_hd__a21o_4
X_85752_ _85751_/CLK _85752_/D _85752_/Q sky130_fd_sc_hd__dfxtp_4
X_82964_ _82774_/CLK _82964_/D _82964_/Q sky130_fd_sc_hd__dfxtp_4
X_67898_ _67893_/X _67896_/X _67897_/X _67898_/Y sky130_fd_sc_hd__a21oi_4
X_84703_ _84713_/CLK _59774_/Y _80517_/A sky130_fd_sc_hd__dfxtp_4
X_57651_ _83761_/Q _57651_/Y sky130_fd_sc_hd__inv_2
X_81915_ _82008_/CLK _81915_/D _77127_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_909_0_CLK clkbuf_9_454_0_CLK/X _87851_/CLK sky130_fd_sc_hd__clkbuf_1
X_69637_ _69634_/X _69636_/X _69570_/X _69637_/X sky130_fd_sc_hd__a21o_4
X_54863_ _54883_/A _54857_/B _54883_/C _53170_/D _54863_/X sky130_fd_sc_hd__and4_4
X_66849_ _80918_/D _66734_/X _66848_/X _66849_/X sky130_fd_sc_hd__a21bo_4
X_85683_ _84787_/CLK _85683_/D _85683_/Q sky130_fd_sc_hd__dfxtp_4
X_82895_ _86941_/CLK _78173_/B _41725_/A sky130_fd_sc_hd__dfxtp_4
X_56602_ _56774_/A _56602_/X sky130_fd_sc_hd__buf_2
X_87422_ _82317_/CLK _43437_/X _87422_/Q sky130_fd_sc_hd__dfxtp_4
X_53814_ _53825_/A _71989_/B _53814_/Y sky130_fd_sc_hd__nand2_4
X_84634_ _84634_/CLK _84634_/D _79722_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_5_26_0_CLK clkbuf_5_27_0_CLK/A clkbuf_6_53_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_57582_ _57597_/A _50326_/B _57582_/Y sky130_fd_sc_hd__nand2_4
X_81846_ _82221_/CLK _81846_/D _77518_/A sky130_fd_sc_hd__dfxtp_4
X_69568_ _68934_/X _42543_/Y _69568_/Y sky130_fd_sc_hd__nor2_4
X_54794_ _54798_/A _54816_/B _54798_/C _53103_/D _54794_/X sky130_fd_sc_hd__and4_4
X_59321_ _59311_/X _85735_/Q _59263_/X _59321_/X sky130_fd_sc_hd__o21a_4
X_56533_ _56533_/A _56533_/B _85159_/Q _56533_/Y sky130_fd_sc_hd__nand3_4
X_68519_ _87597_/Q _68066_/X _68517_/X _68518_/X _68519_/X sky130_fd_sc_hd__a211o_4
X_87353_ _81182_/CLK _87353_/D _87353_/Q sky130_fd_sc_hd__dfxtp_4
X_53745_ _53750_/A _48639_/A _53745_/Y sky130_fd_sc_hd__nand2_4
X_84565_ _84603_/CLK _84565_/D _84565_/Q sky130_fd_sc_hd__dfxtp_4
X_50957_ _50957_/A _50957_/X sky130_fd_sc_hd__buf_2
X_69499_ _69496_/X _69498_/X _69499_/Y sky130_fd_sc_hd__nand2_4
X_81777_ _83133_/CLK _81777_/D _49048_/B sky130_fd_sc_hd__dfxtp_4
X_86304_ _86303_/CLK _49894_/Y _72128_/B sky130_fd_sc_hd__dfxtp_4
X_40710_ _40710_/A _40710_/B _40710_/X sky130_fd_sc_hd__or2_4
X_59252_ _84757_/Q _59129_/X _59246_/X _59251_/X _59252_/Y sky130_fd_sc_hd__a2bb2oi_4
X_71530_ _71530_/A _71530_/Y sky130_fd_sc_hd__inv_2
X_83516_ _83520_/CLK _83516_/D _83516_/Q sky130_fd_sc_hd__dfxtp_4
X_56464_ _56525_/A _56545_/A sky130_fd_sc_hd__buf_2
X_80728_ _80728_/CLK _75914_/X _80696_/D sky130_fd_sc_hd__dfxtp_4
X_87284_ _87824_/CLK _87284_/D _69967_/B sky130_fd_sc_hd__dfxtp_4
X_41690_ _41690_/A _41690_/Y sky130_fd_sc_hd__inv_2
X_53676_ _52156_/A _53666_/X _53692_/C _53676_/X sky130_fd_sc_hd__and3_4
X_84496_ _84501_/CLK _61258_/Y _75898_/A sky130_fd_sc_hd__dfxtp_4
X_50888_ _50906_/A _46625_/X _50888_/Y sky130_fd_sc_hd__nand2_4
X_58203_ _58191_/X _58200_/Y _58202_/Y _84909_/D sky130_fd_sc_hd__a21oi_4
X_55415_ _55415_/A _55415_/B _55415_/C _55683_/A sky130_fd_sc_hd__and3_4
X_86235_ _86235_/CLK _86235_/D _86235_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_301 sky130_fd_sc_hd__decap_3
X_40641_ _40640_/X _40641_/X sky130_fd_sc_hd__buf_2
X_52627_ _52643_/A _52605_/X _52643_/C _46707_/X _52627_/X sky130_fd_sc_hd__and4_4
X_59183_ _59160_/X _85650_/Q _59081_/X _59183_/X sky130_fd_sc_hd__o21a_4
X_71461_ _71444_/Y _83490_/Q _71460_/Y _71461_/X sky130_fd_sc_hd__a21o_4
X_83447_ _83480_/CLK _83447_/D _83447_/Q sky130_fd_sc_hd__dfxtp_4
X_56395_ _56383_/X _56386_/B _56395_/C _56395_/Y sky130_fd_sc_hd__nand3_4
XPHY_312 sky130_fd_sc_hd__decap_3
X_80659_ _80657_/CLK _74822_/Y _46141_/A sky130_fd_sc_hd__dfxtp_4
XPHY_323 sky130_fd_sc_hd__decap_3
XPHY_334 sky130_fd_sc_hd__decap_3
X_73200_ _72951_/A _73200_/X sky130_fd_sc_hd__buf_2
X_58134_ _79903_/A _57981_/X _58129_/X _58133_/X _84923_/D sky130_fd_sc_hd__a22oi_4
X_70412_ _70412_/A _70412_/X sky130_fd_sc_hd__buf_2
XPHY_345 sky130_fd_sc_hd__decap_3
X_43360_ _41361_/X _43356_/X _87461_/Q _43357_/X _87461_/D sky130_fd_sc_hd__a2bb2o_4
X_55346_ _55305_/X _55346_/B _55346_/Y sky130_fd_sc_hd__nor2_4
X_74180_ _53588_/B _74180_/B _74181_/B sky130_fd_sc_hd__xor2_4
X_86166_ _83303_/CLK _50621_/Y _86166_/Q sky130_fd_sc_hd__dfxtp_4
X_52558_ _52556_/Y _52541_/X _52557_/Y _85798_/D sky130_fd_sc_hd__a21boi_4
X_40572_ _40380_/X _82880_/Q _40571_/X _40573_/A sky130_fd_sc_hd__o21a_4
XPHY_356 sky130_fd_sc_hd__decap_3
X_71392_ _71372_/Y _83515_/Q _71391_/Y _71392_/X sky130_fd_sc_hd__a21o_4
X_83378_ _83380_/CLK _83378_/D _83378_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_367 sky130_fd_sc_hd__decap_3
XPHY_378 sky130_fd_sc_hd__decap_3
X_42311_ _42307_/X _42297_/X _41606_/X _87927_/Q _42298_/X _42312_/A
+ sky130_fd_sc_hd__o32ai_4
X_73131_ _87057_/Q _73129_/X _73130_/X _73131_/Y sky130_fd_sc_hd__o21ai_4
X_85117_ _85114_/CLK _85117_/D _85117_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_389 sky130_fd_sc_hd__decap_3
X_51509_ _51509_/A _51527_/B _51522_/C _53036_/D _51509_/X sky130_fd_sc_hd__and4_4
X_70343_ _70337_/X _74780_/A _70342_/X _83790_/D sky130_fd_sc_hd__a21o_4
X_58065_ _58813_/A _58065_/X sky130_fd_sc_hd__buf_2
X_82329_ _82327_/CLK _77168_/B _82329_/Q sky130_fd_sc_hd__dfxtp_4
X_43291_ _43260_/X _43269_/X _41174_/X _87495_/Q _43273_/X _43292_/A
+ sky130_fd_sc_hd__o32ai_4
X_55277_ _57349_/B _55272_/A _55128_/X _55276_/X _55277_/X sky130_fd_sc_hd__a211o_4
X_86097_ _86096_/CLK _86097_/D _86097_/Q sky130_fd_sc_hd__dfxtp_4
X_52489_ _52485_/Y _52486_/X _52488_/Y _52489_/Y sky130_fd_sc_hd__a21boi_4
X_45030_ _45026_/Y _45029_/Y _44986_/X _45030_/X sky130_fd_sc_hd__a21o_4
X_57016_ _56966_/X _57007_/X _57015_/Y _57017_/A sky130_fd_sc_hd__o21ai_4
X_42242_ _41416_/X _42222_/X _87963_/Q _42224_/X _87963_/D sky130_fd_sc_hd__a2bb2o_4
X_54228_ _54208_/X _54237_/B _54237_/C _53058_/D _54228_/X sky130_fd_sc_hd__and4_4
X_73062_ _72806_/A _73062_/X sky130_fd_sc_hd__buf_2
X_85048_ _85083_/CLK _85048_/D _85048_/Q sky130_fd_sc_hd__dfxtp_4
X_70274_ _74788_/A _70157_/X _70273_/Y _83815_/D sky130_fd_sc_hd__o21ai_4
X_72013_ _83302_/Q _71985_/X _72012_/Y _72013_/Y sky130_fd_sc_hd__o21ai_4
X_54159_ _85493_/Q _54140_/X _54158_/Y _54159_/Y sky130_fd_sc_hd__o21ai_4
X_42173_ _42083_/A _42173_/X sky130_fd_sc_hd__buf_2
X_77870_ _82161_/Q _82033_/D _82129_/D sky130_fd_sc_hd__xor2_4
X_41124_ _41073_/X _40579_/A _41123_/X _41124_/X sky130_fd_sc_hd__o21a_4
X_76821_ _81637_/D _76821_/B _76821_/Y sky130_fd_sc_hd__xnor2_4
X_46981_ _46981_/A _46944_/B _46981_/C _52785_/D _46981_/X sky130_fd_sc_hd__and4_4
X_58967_ _58963_/Y _58965_/Y _58966_/X _58967_/X sky130_fd_sc_hd__a21o_4
X_86999_ _88363_/CLK _44692_/Y _44691_/A sky130_fd_sc_hd__dfxtp_4
X_48720_ _48718_/Y _48156_/X _48719_/X _86496_/D sky130_fd_sc_hd__a21oi_4
X_79540_ _79536_/Y _79544_/A _79540_/C _79546_/A sky130_fd_sc_hd__nand3_4
X_45932_ _45930_/X _72739_/A _45931_/X _45932_/Y sky130_fd_sc_hd__nand3_4
X_41055_ _41040_/X _41041_/X _41054_/X _69431_/B _41037_/X _41056_/A
+ sky130_fd_sc_hd__o32ai_4
X_57918_ _57952_/A _57918_/B _57918_/Y sky130_fd_sc_hd__nor2_4
X_76752_ _76757_/B _76751_/Y _76753_/B sky130_fd_sc_hd__xnor2_4
X_73964_ _68802_/B _73891_/X _73962_/X _73963_/Y _73964_/X sky130_fd_sc_hd__a211o_4
X_58898_ _86695_/Q _58898_/B _58898_/Y sky130_fd_sc_hd__nor2_4
X_75703_ _75703_/A _75702_/Y _75704_/B sky130_fd_sc_hd__nand2_4
X_48651_ _48651_/A _48651_/X sky130_fd_sc_hd__buf_2
X_72915_ _56181_/X _83076_/Q _72880_/X _72914_/X _72916_/B sky130_fd_sc_hd__a211o_4
X_79471_ _79481_/A _79462_/Y _79470_/X _79471_/Y sky130_fd_sc_hd__o21ai_4
X_45863_ _45860_/X _45862_/Y _45803_/X _45863_/Y sky130_fd_sc_hd__a21oi_4
X_57849_ _58679_/A _57849_/X sky130_fd_sc_hd__buf_2
X_76683_ _81686_/Q _76683_/B _81350_/D sky130_fd_sc_hd__xor2_4
X_73895_ _73895_/A _73873_/B _73895_/Y sky130_fd_sc_hd__nor2_4
X_47602_ _47745_/A _47602_/X sky130_fd_sc_hd__buf_2
X_78422_ _78423_/A _78423_/C _78421_/Y _78422_/X sky130_fd_sc_hd__a21o_4
X_44814_ _41651_/A _43939_/X _67429_/B _43941_/X _86939_/D sky130_fd_sc_hd__a2bb2o_4
X_75634_ _75639_/B _75633_/Y _75635_/B sky130_fd_sc_hd__xor2_4
X_48582_ _48582_/A _48816_/B sky130_fd_sc_hd__buf_2
X_60860_ _61277_/B _61277_/C _61293_/A sky130_fd_sc_hd__nor2_4
X_72846_ _48391_/A _72846_/B _72846_/X sky130_fd_sc_hd__xor2_4
X_45794_ _45792_/Y _45394_/X _45720_/X _45793_/Y _45794_/X sky130_fd_sc_hd__a211o_4
X_47533_ _47530_/X _47549_/B _47519_/X _53103_/D _47533_/X sky130_fd_sc_hd__and4_4
X_59519_ _59557_/A _59562_/B _59519_/C _59520_/A sky130_fd_sc_hd__nand3_4
X_78353_ _78353_/A _78353_/B _78353_/C _78354_/B sky130_fd_sc_hd__nand3_4
X_44745_ _44745_/A _44745_/Y sky130_fd_sc_hd__inv_2
X_75565_ _81057_/D _75564_/Y _75567_/A sky130_fd_sc_hd__nand2_4
X_60791_ _60785_/Y _60820_/A _60708_/Y _60791_/X sky130_fd_sc_hd__and3_4
X_41957_ _41957_/A _41957_/Y sky130_fd_sc_hd__inv_2
X_72777_ _88338_/Q _56939_/X _72776_/X _72777_/Y sky130_fd_sc_hd__o21ai_4
X_77304_ _81927_/Q _82183_/D _81895_/D sky130_fd_sc_hd__xor2_4
X_62530_ _62198_/Y _62622_/A sky130_fd_sc_hd__buf_2
X_74516_ _74515_/X _74516_/X sky130_fd_sc_hd__buf_2
X_40908_ _40931_/A _41085_/A _40907_/X _40908_/X sky130_fd_sc_hd__o21a_4
X_47464_ _47464_/A _47465_/A sky130_fd_sc_hd__inv_2
X_71728_ _58233_/Y _71718_/X _71727_/Y _71728_/Y sky130_fd_sc_hd__o21ai_4
X_78284_ _78282_/X _78284_/B _78283_/Y _78284_/X sky130_fd_sc_hd__and3_4
X_44676_ _44593_/X _44594_/X _40590_/A _44675_/Y _44596_/X _87004_/D
+ sky130_fd_sc_hd__o32ai_4
X_75496_ _80702_/Q _80958_/D _75497_/A sky130_fd_sc_hd__nand2_4
X_41888_ _42547_/A _41888_/X sky130_fd_sc_hd__buf_2
X_49203_ _49198_/Y _49189_/X _49202_/X _86434_/D sky130_fd_sc_hd__a21oi_4
X_46415_ _46403_/X _49029_/A _46414_/X _46416_/A sky130_fd_sc_hd__o21ai_4
X_77235_ _81922_/Q _82178_/D _77235_/X sky130_fd_sc_hd__xor2_4
X_43627_ _87335_/Q _68672_/B sky130_fd_sc_hd__inv_2
X_62461_ _62493_/A _62458_/Y _62461_/C _62461_/D _62461_/Y sky130_fd_sc_hd__nand4_4
X_74447_ _74466_/A _48550_/Y _74447_/Y sky130_fd_sc_hd__nand2_4
X_40839_ _40839_/A _40839_/X sky130_fd_sc_hd__buf_2
X_47395_ _47394_/Y _53021_/B sky130_fd_sc_hd__buf_2
X_71659_ _58513_/Y _71649_/X _71658_/Y _71659_/Y sky130_fd_sc_hd__o21ai_4
X_64200_ _64490_/A _64490_/B _64200_/C _64200_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_7_124_0_CLK clkbuf_6_62_0_CLK/X clkbuf_8_249_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_49134_ _83600_/Q _49135_/A sky130_fd_sc_hd__inv_2
X_61412_ _61412_/A _61413_/A sky130_fd_sc_hd__buf_2
X_46346_ _46258_/A _46346_/X sky130_fd_sc_hd__buf_2
X_65180_ _65178_/X _86731_/Q _65108_/X _65179_/X _65180_/X sky130_fd_sc_hd__a211o_4
X_77166_ _77174_/B _81920_/Q _77165_/Y _77167_/B sky130_fd_sc_hd__a21oi_4
X_43558_ _43557_/X _43546_/X _40480_/X _87361_/Q _43549_/X _43558_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74378_ _57563_/X _74408_/A sky130_fd_sc_hd__buf_2
X_62392_ _62337_/A _61922_/X _62364_/X _62392_/D _62392_/X sky130_fd_sc_hd__and4_4
X_76117_ _76126_/A _76127_/B _76117_/Y sky130_fd_sc_hd__nand2_4
X_64131_ _64128_/X _64129_/X _64130_/Y _84272_/D sky130_fd_sc_hd__a21oi_4
X_42509_ _74005_/A _42509_/Y sky130_fd_sc_hd__inv_2
X_49065_ _49056_/A _50144_/B _49065_/Y sky130_fd_sc_hd__nand2_4
X_73329_ _73495_/A _85867_/Q _73329_/X sky130_fd_sc_hd__and2_4
X_61343_ _61342_/X _61368_/D sky130_fd_sc_hd__buf_2
Xclkbuf_10_94_0_CLK clkbuf_9_47_0_CLK/X _84915_/CLK sky130_fd_sc_hd__clkbuf_1
X_46277_ _46288_/A _53953_/B _46277_/Y sky130_fd_sc_hd__nand2_4
X_77097_ _77097_/A _77097_/B _77097_/Y sky130_fd_sc_hd__nand2_4
X_43489_ _43472_/X _43475_/X _41710_/X _87396_/Q _43479_/X _43490_/A
+ sky130_fd_sc_hd__o32ai_4
X_48016_ _48004_/A _48016_/B _48016_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_240_0_CLK clkbuf_8_241_0_CLK/A clkbuf_8_240_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_45228_ _80672_/Q _45651_/A sky130_fd_sc_hd__buf_2
X_64062_ _60906_/X _64158_/C sky130_fd_sc_hd__buf_2
X_76048_ _76039_/B _76048_/B _76048_/Y sky130_fd_sc_hd__nand2_4
X_61274_ _61262_/A _72544_/B _84490_/Q _61274_/Y sky130_fd_sc_hd__nor3_4
X_63013_ _60383_/A _63014_/D sky130_fd_sc_hd__buf_2
X_60225_ _60291_/C _60255_/B sky130_fd_sc_hd__buf_2
X_45159_ _45127_/X _61521_/B _45144_/X _45159_/Y sky130_fd_sc_hd__o21ai_4
X_68870_ _68757_/A _68870_/X sky130_fd_sc_hd__buf_2
X_79807_ _79807_/A _79807_/B _79820_/B sky130_fd_sc_hd__xnor2_4
X_67821_ _68450_/A _67821_/X sky130_fd_sc_hd__buf_2
X_60156_ _60193_/A _60156_/Y sky130_fd_sc_hd__inv_2
X_49967_ _72301_/B _49960_/X _49966_/Y _49967_/Y sky130_fd_sc_hd__o21ai_4
X_77999_ _77999_/A _77999_/B _78000_/A sky130_fd_sc_hd__nor2_4
Xclkbuf_8_255_0_CLK clkbuf_8_255_0_CLK/A clkbuf_9_510_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_250_0_CLK clkbuf_9_125_0_CLK/X _81872_/CLK sky130_fd_sc_hd__clkbuf_1
X_48918_ _50578_/A _50578_/B _48917_/X _48918_/X sky130_fd_sc_hd__o21a_4
X_67752_ _67678_/X _67752_/B _67752_/X sky130_fd_sc_hd__and2_4
X_79738_ _79735_/X _79737_/Y _79738_/Y sky130_fd_sc_hd__xnor2_4
X_64964_ _64934_/X _86740_/Q _64864_/X _64963_/X _64964_/X sky130_fd_sc_hd__a211o_4
X_60087_ _62548_/B _62576_/C _70056_/A _60087_/Y sky130_fd_sc_hd__a21oi_4
X_49898_ _49925_/A _49904_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_880_0_CLK clkbuf_9_440_0_CLK/X _86733_/CLK sky130_fd_sc_hd__clkbuf_1
X_66703_ _68474_/A _66728_/A sky130_fd_sc_hd__buf_2
X_63915_ _63911_/X _63913_/X _63914_/Y _84287_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_32_0_CLK clkbuf_9_16_0_CLK/X _85152_/CLK sky130_fd_sc_hd__clkbuf_1
X_48849_ _48849_/A _48849_/B _48849_/C _48849_/X sky130_fd_sc_hd__and3_4
X_67683_ _67658_/X _67683_/B _67683_/X sky130_fd_sc_hd__and2_4
X_79669_ _65170_/C _72371_/Y _79668_/Y _79669_/X sky130_fd_sc_hd__o21a_4
X_64895_ _65836_/A _86038_/Q _64895_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_371_0_CLK clkbuf_9_370_0_CLK/A clkbuf_9_371_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_81700_ _84014_/CLK _81700_/D _41096_/B sky130_fd_sc_hd__dfxtp_4
X_69422_ _64636_/A _69746_/A sky130_fd_sc_hd__buf_2
X_66634_ _66683_/A _66634_/B _66634_/X sky130_fd_sc_hd__and2_4
X_51860_ _51870_/A _51851_/B _51851_/C _46810_/X _51860_/X sky130_fd_sc_hd__and4_4
X_63846_ _63831_/A _64282_/A _63862_/C _63846_/X sky130_fd_sc_hd__and3_4
X_82680_ _81216_/CLK _82692_/Q _78240_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_265_0_CLK clkbuf_9_132_0_CLK/X _84869_/CLK sky130_fd_sc_hd__clkbuf_1
X_50811_ _86128_/Q _50727_/X _50810_/Y _50811_/Y sky130_fd_sc_hd__o21ai_4
X_81631_ _81631_/CLK _81631_/D _81631_/Q sky130_fd_sc_hd__dfxtp_4
X_69353_ _83930_/Q _69299_/X _69352_/X _69353_/X sky130_fd_sc_hd__a21bo_4
X_66565_ _66565_/A _69178_/A sky130_fd_sc_hd__buf_2
X_51791_ _51796_/A _51791_/B _51791_/Y sky130_fd_sc_hd__nand2_4
X_63777_ _61354_/B _64192_/B _63757_/C _63776_/X _63777_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_10_895_0_CLK clkbuf_9_447_0_CLK/X _85535_/CLK sky130_fd_sc_hd__clkbuf_1
X_60989_ _60950_/Y _60993_/B _60988_/Y _60989_/X sky130_fd_sc_hd__a21o_4
X_68304_ _83988_/Q _68299_/X _68303_/X _83988_/D sky130_fd_sc_hd__a21bo_4
X_65516_ _65516_/A _65516_/X sky130_fd_sc_hd__buf_2
X_53530_ _53528_/Y _53524_/X _53529_/Y _53530_/Y sky130_fd_sc_hd__a21boi_4
Xclkbuf_10_47_0_CLK clkbuf_9_23_0_CLK/X _83191_/CLK sky130_fd_sc_hd__clkbuf_1
X_84350_ _84350_/CLK _63141_/X _79394_/A sky130_fd_sc_hd__dfxtp_4
X_50742_ _50742_/A _50742_/X sky130_fd_sc_hd__buf_2
X_62728_ _60274_/X _62729_/D sky130_fd_sc_hd__buf_2
X_81562_ _84064_/CLK _81562_/D _81518_/D sky130_fd_sc_hd__dfxtp_4
X_69284_ _83935_/Q _69230_/X _69283_/X _69284_/X sky130_fd_sc_hd__a21bo_4
X_66496_ _66494_/Y _66483_/X _66495_/X _84112_/D sky130_fd_sc_hd__a21o_4
Xclkbuf_9_386_0_CLK clkbuf_9_387_0_CLK/A clkbuf_9_386_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_83301_ _85555_/CLK _72021_/Y _83301_/Q sky130_fd_sc_hd__dfxtp_4
X_80513_ _80513_/A _80512_/Y _82262_/D sky130_fd_sc_hd__xor2_4
X_68235_ _67465_/X _67469_/X _68216_/X _68235_/Y sky130_fd_sc_hd__a21oi_4
X_53461_ _85631_/Q _53449_/X _53460_/Y _53461_/Y sky130_fd_sc_hd__o21ai_4
X_65447_ _65447_/A _65446_/Y _65447_/Y sky130_fd_sc_hd__nand2_4
X_84281_ _84668_/CLK _64010_/Y _80082_/B sky130_fd_sc_hd__dfxtp_4
X_50673_ _50671_/Y _50609_/X _50672_/X _50673_/Y sky130_fd_sc_hd__a21oi_4
X_62659_ _58221_/X _60221_/A _60205_/X _60263_/C _62658_/X _62659_/Y
+ sky130_fd_sc_hd__a41oi_4
X_81493_ _81492_/CLK _84061_/Q _81493_/Q sky130_fd_sc_hd__dfxtp_4
X_55200_ _55196_/A _83748_/Q _55200_/C _55201_/C sky130_fd_sc_hd__nand3_4
X_86020_ _86118_/CLK _86020_/D _86020_/Q sky130_fd_sc_hd__dfxtp_4
X_52412_ _52410_/Y _52390_/X _52411_/X _52412_/Y sky130_fd_sc_hd__a21oi_4
X_83232_ _83229_/CLK _72568_/Y _79414_/B sky130_fd_sc_hd__dfxtp_4
X_80444_ _80458_/A _80458_/B _80467_/A sky130_fd_sc_hd__xor2_4
X_56180_ _73378_/A _73163_/A sky130_fd_sc_hd__buf_2
X_68166_ _82062_/D _68160_/X _68165_/X _68166_/X sky130_fd_sc_hd__a21bo_4
X_53392_ _53311_/A _53397_/A sky130_fd_sc_hd__buf_2
X_65378_ _44149_/X _85507_/Q _64571_/X _65377_/X _65378_/X sky130_fd_sc_hd__a211o_4
X_55131_ _55135_/A _85003_/Q _55131_/X sky130_fd_sc_hd__and2_4
X_67117_ _66758_/X _67117_/X sky130_fd_sc_hd__buf_2
X_52343_ _52334_/A _50133_/B _52343_/Y sky130_fd_sc_hd__nand2_4
X_64329_ _64316_/Y _64327_/X _64328_/X _64329_/X sky130_fd_sc_hd__o21a_4
X_83163_ _86570_/CLK _73145_/X _83163_/Q sky130_fd_sc_hd__dfxtp_4
X_80375_ _80375_/A _80375_/B _80375_/X sky130_fd_sc_hd__xor2_4
X_68097_ _68097_/A _68097_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_208_0_CLK clkbuf_8_209_0_CLK/A clkbuf_8_208_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_203_0_CLK clkbuf_9_101_0_CLK/X _81117_/CLK sky130_fd_sc_hd__clkbuf_1
X_82114_ _82145_/CLK _77728_/X _82114_/Q sky130_fd_sc_hd__dfxtp_4
X_55062_ _55060_/Y _55050_/X _55061_/X _85326_/D sky130_fd_sc_hd__a21oi_4
X_67048_ _87935_/Q _66994_/X _67046_/X _67047_/X _67048_/X sky130_fd_sc_hd__a211o_4
X_52274_ _52274_/A _52295_/A sky130_fd_sc_hd__buf_2
X_87971_ _87720_/CLK _87971_/D _87971_/Q sky130_fd_sc_hd__dfxtp_4
X_83094_ _83846_/CLK _74335_/X _70321_/C sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_833_0_CLK clkbuf_9_416_0_CLK/X _85315_/CLK sky130_fd_sc_hd__clkbuf_1
X_54013_ _53942_/A _52494_/B _54013_/Y sky130_fd_sc_hd__nand2_4
X_51225_ _51220_/A _51203_/B _51225_/C _51225_/D _51225_/X sky130_fd_sc_hd__and4_4
X_86922_ _87652_/CLK _86922_/D _67836_/B sky130_fd_sc_hd__dfxtp_4
X_82045_ _82047_/CLK _77981_/Y _82013_/D sky130_fd_sc_hd__dfxtp_4
X_59870_ _59873_/A _59855_/B _80277_/B _59870_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_9_324_0_CLK clkbuf_9_325_0_CLK/A clkbuf_9_324_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_58821_ _58730_/X _85933_/Q _58810_/X _58821_/X sky130_fd_sc_hd__o21a_4
X_51156_ _51128_/A _51156_/X sky130_fd_sc_hd__buf_2
X_86853_ _86855_/CLK _45807_/Y _62126_/D sky130_fd_sc_hd__dfxtp_4
X_68999_ _68999_/A _74166_/A _68999_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_218_0_CLK clkbuf_9_109_0_CLK/X _84375_/CLK sky130_fd_sc_hd__clkbuf_1
X_50107_ _50104_/Y _50092_/X _50106_/X _86263_/D sky130_fd_sc_hd__a21oi_4
X_85804_ _86040_/CLK _52529_/Y _65144_/B sky130_fd_sc_hd__dfxtp_4
X_58752_ _58868_/A _58752_/X sky130_fd_sc_hd__buf_2
X_51087_ _86076_/Q _51073_/X _51086_/Y _51087_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_848_0_CLK clkbuf_9_424_0_CLK/X _82394_/CLK sky130_fd_sc_hd__clkbuf_1
X_55964_ _74547_/C _55690_/X _44102_/X _55963_/X _55965_/B sky130_fd_sc_hd__a211o_4
X_86784_ _86784_/CLK _46070_/Y _86784_/Q sky130_fd_sc_hd__dfxtp_4
X_83996_ _82642_/CLK _83996_/D _82644_/D sky130_fd_sc_hd__dfxtp_4
X_57703_ _57872_/A _57703_/X sky130_fd_sc_hd__buf_2
X_50038_ _50048_/A _51728_/B _50038_/Y sky130_fd_sc_hd__nand2_4
X_54915_ _54889_/A _54932_/C sky130_fd_sc_hd__buf_2
X_85735_ _85735_/CLK _52896_/Y _85735_/Q sky130_fd_sc_hd__dfxtp_4
X_58683_ _58682_/X _85784_/Q _58594_/X _58683_/X sky130_fd_sc_hd__o21a_4
X_70961_ _70961_/A _70961_/X sky130_fd_sc_hd__buf_2
X_82947_ _82961_/CLK _82755_/Q _82947_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_339_0_CLK clkbuf_9_339_0_CLK/A clkbuf_9_339_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_55895_ _56219_/C _44070_/B _44051_/A _55894_/X _55895_/X sky130_fd_sc_hd__a211o_4
X_72700_ _72710_/A _56824_/X _55254_/A _55253_/X _72700_/X sky130_fd_sc_hd__and4_4
X_57634_ _46249_/A _71985_/A sky130_fd_sc_hd__buf_2
X_42860_ _42860_/A _42860_/Y sky130_fd_sc_hd__inv_2
X_54846_ _85367_/Q _54839_/X _54845_/Y _54846_/Y sky130_fd_sc_hd__o21ai_4
X_73680_ _73676_/X _73678_/X _73679_/X _73694_/B sky130_fd_sc_hd__a21o_4
X_85666_ _85471_/CLK _53262_/Y _85666_/Q sky130_fd_sc_hd__dfxtp_4
X_70892_ _70905_/D _70899_/D sky130_fd_sc_hd__buf_2
X_82878_ _82942_/CLK _78290_/B _82878_/Q sky130_fd_sc_hd__dfxtp_4
X_87405_ _87471_/CLK _87405_/D _87405_/Q sky130_fd_sc_hd__dfxtp_4
X_41811_ _40404_/X _41799_/X _88140_/Q _41800_/X _88140_/D sky130_fd_sc_hd__a2bb2o_4
X_72631_ _72630_/X _72631_/X sky130_fd_sc_hd__buf_2
X_84617_ _83218_/CLK _60424_/X _79157_/A sky130_fd_sc_hd__dfxtp_4
X_57565_ _57564_/X _53531_/B _57565_/Y sky130_fd_sc_hd__nand2_4
X_81829_ _80708_/CLK _81861_/Q _77265_/A sky130_fd_sc_hd__dfxtp_4
X_88385_ _88386_/CLK _88385_/D _88385_/Q sky130_fd_sc_hd__dfxtp_4
X_42791_ _41367_/X _42787_/X _67700_/B _42788_/X _87716_/D sky130_fd_sc_hd__a2bb2o_4
X_54777_ _54758_/X _47506_/A _54777_/Y sky130_fd_sc_hd__nand2_4
X_85597_ _85596_/CLK _53642_/Y _85597_/Q sky130_fd_sc_hd__dfxtp_4
X_51989_ _51986_/Y _51987_/X _51988_/X _85911_/D sky130_fd_sc_hd__a21oi_4
X_59304_ _59256_/A _86344_/Q _59304_/Y sky130_fd_sc_hd__nor2_4
X_44530_ _44530_/A _44530_/X sky130_fd_sc_hd__buf_2
X_56516_ _56523_/A _56520_/B _55814_/B _56516_/Y sky130_fd_sc_hd__nand3_4
X_75350_ _80693_/Q _80949_/D _75351_/A sky130_fd_sc_hd__nand2_4
X_87336_ _87045_/CLK _43626_/X _73822_/A sky130_fd_sc_hd__dfxtp_4
X_41742_ _41741_/X _41722_/X _67840_/B _41723_/X _88158_/D sky130_fd_sc_hd__a2bb2o_4
X_53728_ _53990_/A _53729_/A sky130_fd_sc_hd__buf_2
X_72562_ _72562_/A _72562_/Y sky130_fd_sc_hd__inv_2
X_84548_ _84529_/CLK _84548_/D _60959_/C sky130_fd_sc_hd__dfxtp_4
X_57496_ _84992_/Q _57493_/X _57495_/Y _57496_/Y sky130_fd_sc_hd__o21ai_4
X_74301_ _72686_/A _74301_/X sky130_fd_sc_hd__buf_2
X_59235_ _59208_/X _86062_/Q _59234_/X _59235_/Y sky130_fd_sc_hd__o21ai_4
X_71513_ _53232_/B _71508_/X _71512_/Y _83472_/D sky130_fd_sc_hd__o21ai_4
X_44461_ _44461_/A _44461_/Y sky130_fd_sc_hd__inv_2
X_56447_ _56153_/X _56439_/X _56446_/Y _56447_/Y sky130_fd_sc_hd__o21ai_4
X_75281_ _75258_/X _75259_/Y _75261_/A _75281_/Y sky130_fd_sc_hd__a21boi_4
X_87267_ _88034_/CLK _43788_/X _69358_/B sky130_fd_sc_hd__dfxtp_4
X_53659_ _53657_/Y _53653_/X _53658_/X _85593_/D sky130_fd_sc_hd__a21oi_4
X_41673_ _41825_/A _41673_/X sky130_fd_sc_hd__buf_2
X_72493_ _72484_/X _83382_/Q _72492_/Y _83246_/D sky130_fd_sc_hd__o21a_4
X_84479_ _84481_/CLK _61457_/Y _84479_/Q sky130_fd_sc_hd__dfxtp_4
X_46200_ _46199_/X _72527_/B sky130_fd_sc_hd__buf_2
XPHY_120 sky130_fd_sc_hd__decap_3
X_77020_ _77014_/Y _77019_/Y _77011_/B _77020_/Y sky130_fd_sc_hd__a21oi_4
X_43412_ _43396_/A _43412_/X sky130_fd_sc_hd__buf_2
X_74232_ _74232_/A _74232_/B _74232_/X sky130_fd_sc_hd__and2_4
X_86218_ _86218_/CLK _50353_/Y _86218_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_131 sky130_fd_sc_hd__decap_3
X_40624_ _40624_/A _40623_/X _40624_/X sky130_fd_sc_hd__or2_4
X_47180_ _47180_/A _52900_/D sky130_fd_sc_hd__buf_2
X_71444_ _71444_/A _71444_/Y sky130_fd_sc_hd__inv_2
X_59166_ _59162_/Y _59164_/Y _59165_/X _59166_/X sky130_fd_sc_hd__a21o_4
X_44392_ _44392_/A _87132_/D sky130_fd_sc_hd__inv_2
XPHY_142 sky130_fd_sc_hd__decap_3
X_56378_ _56377_/X _56378_/X sky130_fd_sc_hd__buf_2
X_87198_ _87720_/CLK _87198_/D _67845_/B sky130_fd_sc_hd__dfxtp_4
XPHY_153 sky130_fd_sc_hd__decap_3
XPHY_164 sky130_fd_sc_hd__decap_3
X_46131_ _46107_/A _46115_/A _46133_/C sky130_fd_sc_hd__nor2_4
X_58117_ _86628_/Q _57954_/X _58117_/Y sky130_fd_sc_hd__nor2_4
XPHY_175 sky130_fd_sc_hd__decap_3
X_43343_ _43342_/Y _87469_/D sky130_fd_sc_hd__inv_2
X_55329_ _55201_/Y _55299_/Y _55328_/X _55329_/Y sky130_fd_sc_hd__o21ai_4
X_74163_ _83120_/Q _74139_/X _74162_/Y _83120_/D sky130_fd_sc_hd__a21o_4
X_86149_ _86149_/CLK _86149_/D _86149_/Q sky130_fd_sc_hd__dfxtp_4
X_40555_ _40554_/X _40556_/A sky130_fd_sc_hd__buf_2
XPHY_186 sky130_fd_sc_hd__decap_3
X_59097_ _59033_/X _85433_/Q _59096_/X _59097_/Y sky130_fd_sc_hd__o21ai_4
X_71375_ _71485_/B _71458_/C sky130_fd_sc_hd__buf_2
XPHY_197 sky130_fd_sc_hd__decap_3
X_73114_ _73183_/A _86484_/Q _73114_/X sky130_fd_sc_hd__and2_4
X_58048_ _84929_/Q _58048_/Y sky130_fd_sc_hd__inv_2
X_70326_ _70326_/A _70183_/A _70183_/B _70183_/D _70326_/Y sky130_fd_sc_hd__nand4_4
X_46062_ _43611_/A _46062_/X sky130_fd_sc_hd__buf_2
X_43274_ _43260_/X _43269_/X _41125_/X _87505_/Q _43273_/X _43274_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74094_ _70128_/A _73549_/X _74093_/Y _83123_/D sky130_fd_sc_hd__a21o_4
X_78971_ _78948_/Y _79115_/A _78959_/Y _78960_/Y _78971_/X sky130_fd_sc_hd__o22a_4
X_40486_ _40485_/X _40410_/X _88384_/Q _40411_/X _40486_/X sky130_fd_sc_hd__a2bb2o_4
X_45013_ _56306_/C _44979_/X _45012_/X _45013_/X sky130_fd_sc_hd__o21a_4
X_42225_ _41371_/X _42222_/X _87971_/Q _42224_/X _87971_/D sky130_fd_sc_hd__a2bb2o_4
X_77922_ _77916_/B _77916_/A _77921_/Y _77922_/Y sky130_fd_sc_hd__a21oi_4
X_73045_ _72881_/A _65584_/B _73045_/X sky130_fd_sc_hd__and2_4
X_70257_ _70255_/X _74771_/A _70256_/X _70257_/X sky130_fd_sc_hd__a21o_4
X_60010_ _62504_/A _62478_/A sky130_fd_sc_hd__buf_2
X_49821_ _86317_/Q _49798_/X _49820_/Y _49821_/Y sky130_fd_sc_hd__o21ai_4
X_42156_ _42155_/Y _88007_/D sky130_fd_sc_hd__inv_2
X_77853_ _77851_/Y _77852_/Y _77861_/A sky130_fd_sc_hd__xor2_4
X_70188_ _70200_/A _70200_/B _70188_/C _70200_/D _70188_/X sky130_fd_sc_hd__and4_4
X_59999_ _59931_/X _60000_/A sky130_fd_sc_hd__inv_2
X_41107_ _41100_/X _81698_/Q _41106_/X _41107_/Y sky130_fd_sc_hd__o21ai_4
X_76804_ _81667_/Q _76804_/B _76804_/Y sky130_fd_sc_hd__xnor2_4
X_49752_ _49749_/Y _49732_/X _49751_/X _49752_/Y sky130_fd_sc_hd__a21oi_4
X_46964_ _46964_/A _52775_/D sky130_fd_sc_hd__buf_2
X_42087_ _40986_/X _42072_/X _88041_/Q _42073_/X _42087_/X sky130_fd_sc_hd__a2bb2o_4
X_77784_ _77796_/A _77783_/Y _77785_/B sky130_fd_sc_hd__xor2_4
X_74996_ _75001_/A _74986_/X _74995_/Y _74996_/Y sky130_fd_sc_hd__a21boi_4
X_48703_ _48696_/Y _48651_/X _48702_/X _48703_/Y sky130_fd_sc_hd__a21oi_4
X_79523_ _79164_/Y _79523_/B _79523_/X sky130_fd_sc_hd__xor2_4
X_41038_ _40999_/X _41000_/X _41036_/X _88289_/Q _41037_/X _41039_/A
+ sky130_fd_sc_hd__o32ai_4
X_45915_ _44020_/A _45915_/X sky130_fd_sc_hd__buf_2
X_76735_ _81692_/Q _76735_/B _76735_/Y sky130_fd_sc_hd__xnor2_4
X_49683_ _59327_/B _49660_/X _49682_/Y _49683_/Y sky130_fd_sc_hd__o21ai_4
X_61961_ _61958_/Y _61959_/X _61960_/Y _84443_/D sky130_fd_sc_hd__a21oi_4
X_73947_ _44709_/Y _73728_/X _73946_/Y _73947_/X sky130_fd_sc_hd__a21o_4
X_46895_ _46894_/Y _52735_/D sky130_fd_sc_hd__buf_2
X_63700_ _63624_/X _63694_/X _63695_/X _63698_/X _63699_/Y _63700_/Y
+ sky130_fd_sc_hd__o41ai_4
X_48634_ _48634_/A _48841_/A sky130_fd_sc_hd__buf_2
X_60912_ _60870_/X _60994_/A sky130_fd_sc_hd__buf_2
X_79454_ _58639_/Y _66395_/C _79453_/Y _79470_/A sky130_fd_sc_hd__o21a_4
X_45846_ _56898_/A _45798_/X _44889_/A _45846_/X sky130_fd_sc_hd__o21a_4
X_64680_ _64680_/A _86270_/Q _64680_/X sky130_fd_sc_hd__and2_4
X_76666_ _76664_/A _76662_/Y _76661_/A _76666_/Y sky130_fd_sc_hd__a21oi_4
X_73878_ _73949_/A _66094_/B _73878_/X sky130_fd_sc_hd__and2_4
X_61892_ _61747_/X _61910_/D sky130_fd_sc_hd__buf_2
X_78405_ _78405_/A _78405_/Y sky130_fd_sc_hd__inv_2
X_63631_ _61590_/B _63609_/X _63629_/X _63630_/Y _63631_/X sky130_fd_sc_hd__a211o_4
X_75617_ _75617_/A _75617_/B _80967_/D sky130_fd_sc_hd__xor2_4
X_72829_ _72829_/A _72829_/X sky130_fd_sc_hd__buf_2
X_48565_ _49067_/B _48565_/B _48565_/Y sky130_fd_sc_hd__nand2_4
X_60843_ _60843_/A _61071_/A _59602_/A _60406_/B _60843_/X sky130_fd_sc_hd__and4_4
X_79385_ _79385_/A _79385_/B _79391_/B sky130_fd_sc_hd__xor2_4
X_45777_ _62094_/D _63280_/B sky130_fd_sc_hd__buf_2
X_76597_ _76593_/Y _76597_/B _76596_/Y _76597_/X sky130_fd_sc_hd__or3_4
X_42989_ _42988_/Y _87617_/D sky130_fd_sc_hd__inv_2
X_47516_ _47516_/A _53095_/B sky130_fd_sc_hd__buf_2
X_66350_ _64923_/A _86562_/Q _66350_/X sky130_fd_sc_hd__and2_4
X_78336_ _78337_/C _78334_/Y _78335_/Y _78339_/A sky130_fd_sc_hd__a21oi_4
X_44728_ _44707_/X _44708_/X _40716_/A _44727_/Y _44710_/X _86984_/D
+ sky130_fd_sc_hd__o32ai_4
X_63562_ _63562_/A _60712_/B _60739_/X _63562_/Y sky130_fd_sc_hd__nor3_4
X_75548_ _75547_/Y _75544_/X _75562_/A sky130_fd_sc_hd__nand2_4
X_48496_ _48495_/Y _48485_/B _48496_/Y sky130_fd_sc_hd__nand2_4
X_60774_ _63374_/A _60758_/X _60773_/Y _84570_/Q _60341_/X _60774_/X
+ sky130_fd_sc_hd__o32a_4
X_65301_ _64642_/A _65301_/X sky130_fd_sc_hd__buf_2
X_62513_ _62483_/X _62541_/B _76981_/B _62513_/Y sky130_fd_sc_hd__nor3_4
X_47447_ _54743_/D _53052_/D sky130_fd_sc_hd__buf_2
X_66281_ _66277_/Y _66278_/X _66280_/X _84144_/D sky130_fd_sc_hd__a21o_4
XPHY_0 sky130_fd_sc_hd__decap_3
X_78267_ _78250_/A _78265_/Y _78266_/Y _78282_/A sky130_fd_sc_hd__a21o_4
X_44659_ _44567_/A _44659_/X sky130_fd_sc_hd__buf_2
X_63493_ _63517_/A _63517_/B _63493_/C _63493_/Y sky130_fd_sc_hd__nor3_4
X_75479_ _75457_/A _75457_/B _75456_/A _75479_/X sky130_fd_sc_hd__o21a_4
X_68020_ _68044_/A _68020_/B _68020_/X sky130_fd_sc_hd__and2_4
X_65232_ _65099_/X _83289_/Q _65230_/X _65231_/X _65233_/B sky130_fd_sc_hd__a211o_4
X_77218_ _77216_/Y _77212_/Y _77217_/Y _77219_/B sky130_fd_sc_hd__o21ai_4
X_62444_ _62415_/X _61980_/A _62618_/D _62194_/D _62444_/X sky130_fd_sc_hd__and4_4
X_47378_ _47378_/A _47379_/A sky130_fd_sc_hd__inv_2
X_78198_ _78198_/A _82491_/Q _78204_/B sky130_fd_sc_hd__xor2_4
X_49117_ _49117_/A _50169_/B _49117_/Y sky130_fd_sc_hd__nand2_4
X_46329_ _46262_/X _48947_/A _46328_/X _46330_/A sky130_fd_sc_hd__o21ai_4
X_65163_ _64683_/A _65631_/B sky130_fd_sc_hd__buf_2
X_77149_ _77149_/A _81918_/Q _77149_/Y sky130_fd_sc_hd__nand2_4
X_62375_ _62319_/A _63496_/B _62375_/C _62378_/C sky130_fd_sc_hd__nand3_4
X_64114_ _84873_/Q _64136_/B _64114_/X sky130_fd_sc_hd__or2_4
X_61326_ _59834_/A _61587_/B _84489_/Q _61326_/X sky130_fd_sc_hd__or3_4
X_49048_ _49048_/A _49048_/B _50645_/A sky130_fd_sc_hd__nor2_4
X_80160_ _80147_/X _80158_/X _80159_/X _80160_/Y sky130_fd_sc_hd__a21oi_4
X_65094_ _64946_/A _65094_/B _65094_/X sky130_fd_sc_hd__and2_4
X_69971_ _69968_/X _69970_/X _66547_/X _69971_/X sky130_fd_sc_hd__a21o_4
X_64045_ _64045_/A _64045_/X sky130_fd_sc_hd__buf_2
X_68922_ _69035_/A _68922_/X sky130_fd_sc_hd__buf_2
X_61257_ _64689_/A _72604_/B _75898_/A _61218_/Y _61256_/Y _61258_/A
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_7_54_0_CLK clkbuf_7_55_0_CLK/A clkbuf_7_54_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_80091_ _80091_/A _63995_/C _80091_/X sky130_fd_sc_hd__xor2_4
X_51010_ _51010_/A _51039_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_194_0_CLK clkbuf_7_97_0_CLK/X clkbuf_9_389_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_60208_ _60387_/A _60164_/Y _60166_/X _61316_/A _60174_/X _62644_/A
+ sky130_fd_sc_hd__a32oi_4
X_68853_ _68785_/A _88256_/Q _68853_/X sky130_fd_sc_hd__and2_4
X_61188_ _61105_/X _61188_/B _61188_/C _61188_/Y sky130_fd_sc_hd__nand3_4
X_67804_ _67782_/X _67792_/Y _67747_/X _67803_/Y _67804_/X sky130_fd_sc_hd__a211o_4
X_60139_ _60125_/A _60214_/B _60139_/C _60139_/Y sky130_fd_sc_hd__nor3_4
X_83850_ _82536_/CLK _70097_/X _82530_/D sky130_fd_sc_hd__dfxtp_4
X_68784_ _69014_/A _68785_/A sky130_fd_sc_hd__buf_2
X_65996_ _65993_/X _65995_/X _65880_/X _65999_/A sky130_fd_sc_hd__a21o_4
X_82801_ _82833_/CLK _82833_/Q _82801_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_69_0_CLK clkbuf_7_69_0_CLK/A clkbuf_7_69_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_67735_ _67496_/X _67726_/Y _67624_/X _67734_/Y _67735_/X sky130_fd_sc_hd__a211o_4
X_52961_ _53097_/A _53069_/A sky130_fd_sc_hd__buf_2
X_64947_ _64944_/X _86164_/Q _64766_/X _64946_/X _64947_/X sky130_fd_sc_hd__a211o_4
X_83781_ _85953_/CLK _70390_/Y _83781_/Q sky130_fd_sc_hd__dfxtp_4
X_80993_ _81990_/CLK _75880_/Y _80949_/D sky130_fd_sc_hd__dfxtp_4
X_54700_ _54672_/X _54721_/C sky130_fd_sc_hd__buf_2
X_85520_ _86246_/CLK _54027_/Y _85520_/Q sky130_fd_sc_hd__dfxtp_4
X_51912_ _85923_/Q _51900_/X _51911_/Y _51912_/Y sky130_fd_sc_hd__o21ai_4
X_82732_ _82692_/CLK _84116_/Q _82732_/Q sky130_fd_sc_hd__dfxtp_4
X_67666_ _87973_/Q _67591_/X _67641_/X _67665_/X _67666_/X sky130_fd_sc_hd__a211o_4
X_55680_ _55290_/Y _55680_/B _55680_/Y sky130_fd_sc_hd__nor2_4
X_52892_ _52892_/A _52892_/X sky130_fd_sc_hd__buf_2
X_64878_ _64877_/X _86423_/Q _64878_/X sky130_fd_sc_hd__and2_4
X_69405_ _69733_/A _69405_/X sky130_fd_sc_hd__buf_2
X_54631_ _54628_/Y _54611_/X _54630_/X _54631_/Y sky130_fd_sc_hd__a21oi_4
X_85451_ _85773_/CLK _85451_/D _85451_/Q sky130_fd_sc_hd__dfxtp_4
X_66617_ _87889_/Q _66529_/X _66531_/X _66616_/X _66617_/X sky130_fd_sc_hd__a211o_4
X_51843_ _51843_/A _51851_/B sky130_fd_sc_hd__buf_2
X_63829_ _63734_/A _64184_/A sky130_fd_sc_hd__buf_2
X_82663_ _82665_/CLK _82663_/D _78112_/A sky130_fd_sc_hd__dfxtp_4
X_67597_ _87464_/Q _67594_/X _67595_/X _67596_/X _67597_/X sky130_fd_sc_hd__a211o_4
X_84402_ _84293_/CLK _62555_/Y _84402_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_132_0_CLK clkbuf_7_66_0_CLK/X clkbuf_8_132_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_57350_ _57348_/X _57349_/Y _57331_/B _57351_/B sky130_fd_sc_hd__a21o_4
X_81614_ _81296_/CLK _76326_/B _81614_/Q sky130_fd_sc_hd__dfxtp_4
X_69336_ _87025_/Q _69239_/X _69103_/X _69335_/X _69336_/X sky130_fd_sc_hd__a211o_4
X_88170_ _87471_/CLK _88170_/D _67563_/B sky130_fd_sc_hd__dfxtp_4
X_54562_ _85419_/Q _54540_/X _54561_/Y _54562_/Y sky130_fd_sc_hd__o21ai_4
X_66548_ _66536_/X _66545_/X _66547_/X _66548_/X sky130_fd_sc_hd__a21o_4
X_85382_ _85379_/CLK _85382_/D _85382_/Q sky130_fd_sc_hd__dfxtp_4
X_51774_ _51779_/A _46662_/X _51774_/Y sky130_fd_sc_hd__nand2_4
X_82594_ _82595_/CLK _78805_/B _82562_/D sky130_fd_sc_hd__dfxtp_4
X_56301_ _56296_/A _56298_/X _85244_/Q _56301_/Y sky130_fd_sc_hd__nand3_4
X_87121_ _87686_/CLK _44414_/X _87121_/Q sky130_fd_sc_hd__dfxtp_4
X_53513_ _53510_/Y _53498_/X _53512_/Y _53513_/Y sky130_fd_sc_hd__a21boi_4
X_84333_ _84333_/CLK _63328_/Y _79197_/B sky130_fd_sc_hd__dfxtp_4
X_50725_ _50209_/A _50751_/B _50668_/C _50725_/X sky130_fd_sc_hd__and3_4
X_81545_ _81344_/CLK _81545_/D _81545_/Q sky130_fd_sc_hd__dfxtp_4
X_57281_ _57268_/X _57149_/B _56733_/X _56735_/X _57270_/X _57281_/X
+ sky130_fd_sc_hd__a41o_4
X_69267_ _69264_/X _69266_/X _69267_/Y sky130_fd_sc_hd__nand2_4
X_54493_ _54385_/A _54503_/B sky130_fd_sc_hd__buf_2
X_66479_ _66445_/A _66514_/B _66478_/Y _66479_/Y sky130_fd_sc_hd__nor3_4
X_59020_ _58918_/X _59018_/Y _59019_/Y _58959_/X _58923_/X _59020_/X
+ sky130_fd_sc_hd__o32a_4
X_56232_ _56245_/A _56243_/B sky130_fd_sc_hd__buf_2
X_68218_ _68188_/X _67340_/Y _68207_/X _68217_/Y _68218_/X sky130_fd_sc_hd__a211o_4
X_87052_ _87813_/CLK _44570_/Y _87052_/Q sky130_fd_sc_hd__dfxtp_4
X_53444_ _53443_/A _47829_/A _53443_/Y _53444_/X sky130_fd_sc_hd__o21a_4
X_84264_ _84263_/CLK _64232_/X _79872_/B sky130_fd_sc_hd__dfxtp_4
X_50656_ _50728_/A _50657_/A sky130_fd_sc_hd__buf_2
X_81476_ _88121_/CLK _84044_/Q _81476_/Q sky130_fd_sc_hd__dfxtp_4
X_69198_ _69195_/X _69197_/X _69198_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_147_0_CLK clkbuf_7_73_0_CLK/X clkbuf_9_295_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_86003_ _85712_/CLK _86003_/D _86003_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_142_0_CLK clkbuf_9_71_0_CLK/X _81811_/CLK sky130_fd_sc_hd__clkbuf_1
X_83215_ _84350_/CLK _72616_/Y _79231_/B sky130_fd_sc_hd__dfxtp_4
X_56163_ _56163_/A _56162_/X _56164_/A sky130_fd_sc_hd__xnor2_4
X_80427_ _80411_/Y _80414_/Y _80426_/X _80427_/X sky130_fd_sc_hd__a21o_4
X_68149_ _66940_/X _66943_/X _68133_/X _68149_/Y sky130_fd_sc_hd__a21oi_4
X_53375_ _53347_/A _53388_/B sky130_fd_sc_hd__buf_2
X_84195_ _84192_/CLK _84195_/D _65531_/C sky130_fd_sc_hd__dfxtp_4
X_50587_ _86172_/Q _50563_/X _50586_/Y _50587_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_772_0_CLK clkbuf_9_386_0_CLK/X _82610_/CLK sky130_fd_sc_hd__clkbuf_1
X_55114_ _55118_/A _47809_/A _55114_/Y sky130_fd_sc_hd__nand2_4
X_40340_ _44362_/A _47363_/A sky130_fd_sc_hd__buf_2
X_52326_ _52334_/A _49006_/X _52326_/Y sky130_fd_sc_hd__nand2_4
X_71160_ _71041_/X _71173_/B _71160_/C _71160_/D _71160_/Y sky130_fd_sc_hd__nand4_4
X_83146_ _86218_/CLK _73548_/X _83146_/Q sky130_fd_sc_hd__dfxtp_4
X_80358_ _80358_/A _80357_/X _80358_/Y sky130_fd_sc_hd__xnor2_4
X_56094_ _56094_/A _56094_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_263_0_CLK clkbuf_9_262_0_CLK/A clkbuf_9_263_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_70111_ _83124_/Q _70111_/Y sky130_fd_sc_hd__inv_2
X_55045_ _55042_/Y _55024_/X _55044_/X _55045_/Y sky130_fd_sc_hd__a21oi_4
X_59922_ _60058_/B _59913_/X _59922_/C _59922_/X sky130_fd_sc_hd__and3_4
X_52257_ _52188_/A _50556_/B _52257_/Y sky130_fd_sc_hd__nand2_4
X_71091_ _71088_/A _71091_/B _71088_/C _71091_/Y sky130_fd_sc_hd__nand3_4
X_83077_ _83282_/CLK _83077_/D _83077_/Q sky130_fd_sc_hd__dfxtp_4
X_87954_ _87950_/CLK _87954_/D _87954_/Q sky130_fd_sc_hd__dfxtp_4
X_80289_ _80284_/Y _80273_/Y _80282_/Y _80302_/B sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_157_0_CLK clkbuf_9_78_0_CLK/X _81304_/CLK sky130_fd_sc_hd__clkbuf_1
X_42010_ _41993_/A _42010_/X sky130_fd_sc_hd__buf_2
X_51208_ _51206_/Y _51201_/X _51207_/X _51208_/Y sky130_fd_sc_hd__a21oi_4
X_70042_ _70040_/X _69785_/Y _70033_/X _70041_/Y _70042_/X sky130_fd_sc_hd__a211o_4
X_86905_ _86882_/CLK _45011_/Y _64284_/B sky130_fd_sc_hd__dfxtp_4
X_82028_ _81989_/CLK _77824_/B _81996_/D sky130_fd_sc_hd__dfxtp_4
X_59853_ _59855_/A _59855_/B _84688_/Q _59853_/Y sky130_fd_sc_hd__nor3_4
X_52188_ _52188_/A _52188_/B _52188_/Y sky130_fd_sc_hd__nand2_4
X_87885_ _88144_/CLK _42393_/X _87885_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_787_0_CLK clkbuf_9_393_0_CLK/X _82743_/CLK sky130_fd_sc_hd__clkbuf_1
X_58804_ _58699_/A _58804_/B _58804_/Y sky130_fd_sc_hd__nor2_4
X_51139_ _51130_/A _52833_/B _51139_/Y sky130_fd_sc_hd__nand2_4
X_86836_ _87625_/CLK _86836_/D _66618_/B sky130_fd_sc_hd__dfxtp_4
X_74850_ _81122_/D _74848_/B _74850_/Y sky130_fd_sc_hd__nand2_4
X_59784_ _66262_/A _59848_/B sky130_fd_sc_hd__buf_2
X_56996_ _56993_/X _56994_/Y _56995_/X _56996_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_278_0_CLK clkbuf_9_278_0_CLK/A clkbuf_9_278_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_73801_ _74244_/B _73801_/X sky130_fd_sc_hd__buf_2
X_58735_ _58610_/A _58735_/X sky130_fd_sc_hd__buf_2
X_43961_ _44003_/A _59901_/C sky130_fd_sc_hd__inv_2
X_55947_ _55947_/A _85245_/Q _55947_/X sky130_fd_sc_hd__and2_4
X_74781_ _74781_/A _74775_/A _70884_/A _70662_/X _74781_/Y sky130_fd_sc_hd__nand4_4
X_86767_ _84980_/CLK _86767_/D _44187_/A sky130_fd_sc_hd__dfxtp_4
X_71993_ _71993_/A _71993_/X sky130_fd_sc_hd__buf_2
X_83979_ _87671_/CLK _83979_/D _83979_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_710_0_CLK clkbuf_9_355_0_CLK/X _87103_/CLK sky130_fd_sc_hd__clkbuf_1
X_45700_ _45668_/X _61561_/A _45685_/X _45700_/Y sky130_fd_sc_hd__o21ai_4
X_76520_ _81659_/Q _76520_/Y sky130_fd_sc_hd__inv_2
X_42912_ _41697_/X _42900_/X _87655_/Q _42901_/X _42912_/X sky130_fd_sc_hd__a2bb2o_4
X_73732_ _73709_/X _73733_/A sky130_fd_sc_hd__buf_2
X_85718_ _85718_/CLK _52990_/Y _85718_/Q sky130_fd_sc_hd__dfxtp_4
X_70944_ _70944_/A _70947_/A sky130_fd_sc_hd__buf_2
X_46680_ _46680_/A _46680_/Y sky130_fd_sc_hd__inv_2
X_58666_ _58625_/X _85465_/Q _58665_/X _58666_/Y sky130_fd_sc_hd__o21ai_4
X_43892_ _43862_/X _43876_/X _41321_/X _87212_/Q _43863_/X _43892_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55878_ _55875_/X _55877_/X _55517_/X _55881_/A sky130_fd_sc_hd__a21o_4
X_86698_ _86701_/CLK _86698_/D _58867_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_201_0_CLK clkbuf_9_201_0_CLK/A clkbuf_9_201_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_45631_ _85042_/Q _45631_/Y sky130_fd_sc_hd__inv_2
X_57617_ _71957_/A _57617_/B _57617_/Y sky130_fd_sc_hd__nand2_4
X_76451_ _81271_/Q _81539_/Q _76451_/Y sky130_fd_sc_hd__nand2_4
X_42843_ _41511_/X _42830_/X _66817_/B _42832_/X _87689_/D sky130_fd_sc_hd__a2bb2o_4
X_54829_ _54284_/A _54882_/A sky130_fd_sc_hd__buf_2
X_73663_ _73609_/X _85629_/Q _73661_/X _73662_/X _73663_/X sky130_fd_sc_hd__a211o_4
X_85649_ _85651_/CLK _85649_/D _85649_/Q sky130_fd_sc_hd__dfxtp_4
X_70875_ _70862_/A _70875_/X sky130_fd_sc_hd__buf_2
X_58597_ _58593_/Y _58596_/Y _58105_/X _58597_/X sky130_fd_sc_hd__a21o_4
X_75402_ _75400_/X _75401_/Y _75403_/A sky130_fd_sc_hd__and2_4
X_48350_ _48478_/A _48350_/X sky130_fd_sc_hd__buf_2
X_72614_ _72562_/Y _72570_/C _72614_/X sky130_fd_sc_hd__and2_4
X_79170_ _63338_/Y _79168_/A _79171_/C sky130_fd_sc_hd__nand2_4
X_57548_ _57531_/A _53520_/B _57548_/Y sky130_fd_sc_hd__nand2_4
X_45562_ _45557_/X _45560_/Y _45561_/X _45562_/Y sky130_fd_sc_hd__a21oi_4
X_76382_ _76382_/A _76382_/Y sky130_fd_sc_hd__inv_2
X_88368_ _83139_/CLK _40600_/X _88368_/Q sky130_fd_sc_hd__dfxtp_4
X_42774_ _42720_/X _42774_/X sky130_fd_sc_hd__buf_2
X_73594_ _83144_/Q _73549_/X _73593_/Y _73594_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_10_725_0_CLK clkbuf_9_362_0_CLK/X _82339_/CLK sky130_fd_sc_hd__clkbuf_1
X_47301_ _81817_/Q _47302_/A sky130_fd_sc_hd__inv_2
X_78121_ _78119_/X _78120_/Y _78121_/X sky130_fd_sc_hd__and2_4
X_44513_ _44530_/A _44513_/X sky130_fd_sc_hd__buf_2
X_75333_ _75333_/A _75333_/Y sky130_fd_sc_hd__inv_2
X_87319_ _88084_/CLK _87319_/D _43667_/A sky130_fd_sc_hd__dfxtp_4
X_41725_ _41725_/A _41718_/X _41725_/X sky130_fd_sc_hd__or2_4
X_48281_ _48028_/B _50326_/B sky130_fd_sc_hd__buf_2
X_72545_ _60053_/X _72537_/Y _72539_/Y _72584_/A _72544_/Y _83237_/D
+ sky130_fd_sc_hd__a41oi_4
X_45493_ _56604_/B _45343_/X _45378_/X _45493_/X sky130_fd_sc_hd__o21a_4
X_57479_ _45947_/B _84996_/Q _56646_/Y _57470_/B _57479_/X sky130_fd_sc_hd__a211o_4
X_88299_ _87790_/CLK _40979_/Y _88299_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_216_0_CLK clkbuf_9_217_0_CLK/A clkbuf_9_216_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_47232_ _47196_/A _52931_/B _47232_/Y sky130_fd_sc_hd__nand2_4
X_59218_ _59146_/X _85423_/Q _59217_/X _59218_/Y sky130_fd_sc_hd__o21ai_4
X_78052_ _60826_/C _78052_/B _81861_/D sky130_fd_sc_hd__xor2_4
X_44444_ _44444_/A _87105_/D sky130_fd_sc_hd__inv_2
X_75264_ _75248_/Y _75262_/X _75263_/X _75265_/B sky130_fd_sc_hd__a21boi_4
X_41656_ _41655_/X _41656_/X sky130_fd_sc_hd__buf_2
X_60490_ _60489_/X _63004_/C sky130_fd_sc_hd__buf_2
X_72476_ _72476_/A _72476_/B _72476_/Y sky130_fd_sc_hd__nor2_4
X_77003_ _82082_/Q _77002_/X _82363_/D sky130_fd_sc_hd__xor2_4
X_74215_ _44270_/X _85605_/Q _44272_/X _74214_/X _74215_/X sky130_fd_sc_hd__a211o_4
X_40607_ _40607_/A _40607_/Y sky130_fd_sc_hd__inv_2
X_59149_ _59105_/X _85749_/Q _59106_/X _59149_/X sky130_fd_sc_hd__o21a_4
X_47163_ _47152_/X _47133_/B _47143_/C _52887_/D _47163_/X sky130_fd_sc_hd__and4_4
X_71427_ _71432_/A _71432_/B _71427_/C _71365_/X _71427_/X sky130_fd_sc_hd__and4_4
X_44375_ _44374_/Y _87140_/D sky130_fd_sc_hd__inv_2
X_75195_ _75165_/X _75193_/Y _75194_/X _75195_/X sky130_fd_sc_hd__o21a_4
X_41587_ _41586_/X _41581_/X _67161_/B _41582_/X _88187_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_4_1_0_CLK clkbuf_3_0_1_CLK/X clkbuf_4_1_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_46114_ _46114_/A _80656_/Q _80655_/Q _74846_/B _46204_/B sky130_fd_sc_hd__nor4_4
X_43326_ _43302_/A _43326_/X sky130_fd_sc_hd__buf_2
X_62160_ _61675_/B _62149_/B _61765_/C _61749_/B _62160_/Y sky130_fd_sc_hd__nand4_4
X_74146_ _43094_/Y _72722_/X _72798_/X _74145_/Y _74146_/X sky130_fd_sc_hd__a211o_4
X_40538_ _40537_/Y _40538_/X sky130_fd_sc_hd__buf_2
X_47094_ _47067_/A _47082_/X _47091_/X _52853_/D _47094_/X sky130_fd_sc_hd__and4_4
X_71358_ _71344_/X _83527_/Q _71357_/X _71358_/X sky130_fd_sc_hd__a21o_4
X_61111_ _61101_/A _61122_/C _61122_/B _61195_/A sky130_fd_sc_hd__nand3_4
X_46045_ _41510_/Y _46043_/X _66819_/B _46044_/X _86796_/D sky130_fd_sc_hd__a2bb2o_4
X_70309_ _70303_/X _74729_/A _70308_/X _70309_/X sky130_fd_sc_hd__a21o_4
X_43257_ _43256_/Y _87514_/D sky130_fd_sc_hd__inv_2
X_62091_ _62089_/Y _62033_/X _62090_/Y _62091_/Y sky130_fd_sc_hd__a21oi_4
X_78954_ _78942_/A _78953_/A _78928_/A _82512_/D _78954_/X sky130_fd_sc_hd__a2bb2o_4
X_74077_ _88349_/Q _73153_/X _72901_/X _74077_/Y sky130_fd_sc_hd__o21ai_4
X_40469_ _40468_/Y _40469_/X sky130_fd_sc_hd__buf_2
X_71289_ _71137_/A _71289_/B _71289_/Y sky130_fd_sc_hd__nor2_4
X_42208_ _51584_/A _42258_/A sky130_fd_sc_hd__buf_2
X_61042_ _60918_/X _60957_/B _61041_/Y _61042_/Y sky130_fd_sc_hd__o21ai_4
X_77905_ _82165_/Q _82037_/D _82133_/D sky130_fd_sc_hd__xor2_4
X_73028_ _73704_/A _73028_/X sky130_fd_sc_hd__buf_2
X_43188_ _43188_/A _87547_/D sky130_fd_sc_hd__inv_2
X_78885_ _78885_/A _78885_/B _78888_/A sky130_fd_sc_hd__xor2_4
X_49804_ _49809_/A _53017_/B _49804_/Y sky130_fd_sc_hd__nand2_4
X_42139_ _41130_/X _42137_/X _88016_/Q _42138_/X _88016_/D sky130_fd_sc_hd__a2bb2o_4
X_65850_ _65847_/X _65849_/X _65809_/X _65850_/X sky130_fd_sc_hd__a21o_4
X_77836_ _77822_/Y _77836_/B _77841_/A sky130_fd_sc_hd__nand2_4
X_47996_ _50308_/A _48069_/B _47919_/X _47996_/X sky130_fd_sc_hd__and3_4
X_64801_ _64778_/A _85850_/Q _64801_/X sky130_fd_sc_hd__and2_4
X_49735_ _49731_/Y _49732_/X _49734_/X _49735_/Y sky130_fd_sc_hd__a21oi_4
X_46947_ _54460_/B _52768_/B sky130_fd_sc_hd__buf_2
X_65781_ _65778_/X _65780_/X _65566_/X _65781_/X sky130_fd_sc_hd__a21o_4
X_77767_ _77763_/Y _77766_/Y _77768_/B sky130_fd_sc_hd__xor2_4
X_74979_ _81141_/D _74980_/B _74987_/B sky130_fd_sc_hd__or2_4
X_62993_ _62791_/X _63285_/A sky130_fd_sc_hd__buf_2
X_67520_ _67496_/X _67506_/Y _67507_/X _67519_/Y _67520_/X sky130_fd_sc_hd__a211o_4
X_79506_ _79474_/Y _79496_/B _79491_/Y _79494_/Y _79506_/X sky130_fd_sc_hd__o22a_4
X_64732_ _64732_/A _64761_/B sky130_fd_sc_hd__buf_2
X_76718_ _76688_/A _76694_/A _76718_/Y sky130_fd_sc_hd__nor2_4
X_49666_ _49661_/X _52881_/B _49666_/Y sky130_fd_sc_hd__nand2_4
X_61944_ _61942_/Y _61881_/X _61943_/Y _84444_/D sky130_fd_sc_hd__a21oi_4
X_46878_ _83661_/Q _52726_/B sky130_fd_sc_hd__inv_2
X_77698_ _82240_/Q _77698_/Y sky130_fd_sc_hd__inv_2
X_48617_ _86506_/Q _48612_/X _48616_/Y _48617_/Y sky130_fd_sc_hd__o21ai_4
X_67451_ _67497_/A _67451_/B _67451_/X sky130_fd_sc_hd__and2_4
X_79437_ _79444_/A _79444_/B _79438_/B sky130_fd_sc_hd__xnor2_4
X_45829_ _45825_/X _45828_/X _44898_/X _45829_/X sky130_fd_sc_hd__a21o_4
X_64663_ _64637_/X _64638_/B _64663_/C _64663_/X sky130_fd_sc_hd__and3_4
X_76649_ _81570_/Q _76649_/B _81538_/D sky130_fd_sc_hd__xor2_4
X_49597_ _49571_/A _49610_/A sky130_fd_sc_hd__buf_2
X_61875_ _61437_/B _61843_/B _61860_/C _61860_/D _61875_/Y sky130_fd_sc_hd__nand4_4
X_66402_ _66389_/A _66402_/B _66402_/C _66402_/Y sky130_fd_sc_hd__nor3_4
X_63614_ _63556_/X _63607_/X _63608_/X _63612_/X _63613_/Y _63614_/Y
+ sky130_fd_sc_hd__o41ai_4
X_60826_ _60826_/A _60810_/B _60826_/C _60826_/Y sky130_fd_sc_hd__nor3_4
X_48548_ _48548_/A _48548_/X sky130_fd_sc_hd__buf_2
X_79368_ _79365_/X _79368_/B _82835_/D sky130_fd_sc_hd__xnor2_4
X_67382_ _87409_/Q _67358_/X _67360_/X _67381_/X _67382_/X sky130_fd_sc_hd__a211o_4
X_64594_ _64589_/X _85569_/Q _64591_/X _64593_/X _64594_/X sky130_fd_sc_hd__a211o_4
X_69121_ _69645_/A _69121_/X sky130_fd_sc_hd__buf_2
X_66333_ _66330_/Y _66278_/X _66332_/Y _84140_/D sky130_fd_sc_hd__a21o_4
X_78319_ _78312_/A _82658_/D _78320_/A sky130_fd_sc_hd__nor2_4
X_63545_ _63484_/A _63546_/A sky130_fd_sc_hd__buf_2
X_48479_ _48613_/A _48515_/A sky130_fd_sc_hd__buf_2
X_60757_ _63417_/A _63389_/D sky130_fd_sc_hd__buf_2
X_79299_ _79287_/X _79288_/X _79298_/Y _79303_/A sky130_fd_sc_hd__a21boi_4
X_50510_ _50510_/A _50526_/C sky130_fd_sc_hd__buf_2
X_81330_ _81330_/CLK _76388_/X _81706_/D sky130_fd_sc_hd__dfxtp_4
X_69052_ _69052_/A _69053_/B sky130_fd_sc_hd__inv_2
X_66264_ _66177_/A _66389_/B _66264_/C _66264_/Y sky130_fd_sc_hd__nor3_4
X_51490_ _51488_/Y _51477_/X _51489_/X _86001_/D sky130_fd_sc_hd__a21oi_4
X_63476_ _63463_/A _84960_/Q _63476_/C _63476_/X sky130_fd_sc_hd__and3_4
X_60688_ _60720_/A _60711_/A _60714_/A sky130_fd_sc_hd__nand2_4
X_68003_ _68025_/A _88215_/Q _68003_/X sky130_fd_sc_hd__and2_4
X_65215_ _65210_/X _65214_/X _65161_/X _65215_/X sky130_fd_sc_hd__a21o_4
X_50441_ _86200_/Q _50437_/X _50440_/Y _50441_/Y sky130_fd_sc_hd__o21ai_4
X_62427_ _62425_/Y _62396_/X _62426_/Y _84411_/D sky130_fd_sc_hd__a21oi_4
X_81261_ _81260_/CLK _81261_/D _76301_/A sky130_fd_sc_hd__dfxtp_4
X_66195_ _65737_/X _66195_/B _65740_/X _66204_/A sky130_fd_sc_hd__nand3_4
X_83000_ _83843_/CLK _74649_/X _83000_/Q sky130_fd_sc_hd__dfxtp_4
X_80212_ _80205_/X _80207_/B _80212_/Y sky130_fd_sc_hd__nand2_4
X_53160_ _53158_/Y _53137_/X _53159_/X _85686_/D sky130_fd_sc_hd__a21oi_4
X_65146_ _65669_/A _65146_/X sky130_fd_sc_hd__buf_2
X_50372_ _50381_/A _50372_/B _50372_/Y sky130_fd_sc_hd__nand2_4
X_62358_ _61451_/A _62332_/B _62386_/C _62332_/D _62358_/Y sky130_fd_sc_hd__nand4_4
X_81192_ _81195_/CLK _74940_/X _49140_/A sky130_fd_sc_hd__dfxtp_4
X_52111_ _52100_/A _48391_/X _52111_/Y sky130_fd_sc_hd__nand2_4
X_61309_ _72507_/A _61686_/A sky130_fd_sc_hd__buf_2
X_80143_ _84943_/Q _84191_/Q _80143_/X sky130_fd_sc_hd__xor2_4
X_65077_ _44149_/X _85519_/Q _64571_/X _65076_/X _65077_/X sky130_fd_sc_hd__a211o_4
X_53091_ _53087_/Y _53082_/X _53090_/X _53091_/Y sky130_fd_sc_hd__a21oi_4
X_69954_ _81956_/D _69894_/X _69953_/X _83884_/D sky130_fd_sc_hd__a21bo_4
X_62289_ _62288_/X _62285_/X _64275_/B _60025_/X _62289_/X sky130_fd_sc_hd__and4_4
X_52042_ _52185_/A _52070_/A sky130_fd_sc_hd__buf_2
X_68905_ _68666_/X _68882_/X _68894_/Y _68904_/Y _68905_/X sky130_fd_sc_hd__a211o_4
X_64028_ _60926_/X _64029_/D sky130_fd_sc_hd__buf_2
X_84951_ _84951_/CLK _84951_/D _84951_/Q sky130_fd_sc_hd__dfxtp_4
X_80074_ _80058_/X _80074_/B _80074_/X sky130_fd_sc_hd__or2_4
X_69885_ _69897_/A _69885_/B _69885_/Y sky130_fd_sc_hd__nor2_4
X_83902_ _82234_/CLK _83902_/D _83902_/Q sky130_fd_sc_hd__dfxtp_4
X_56850_ _56849_/X _56850_/X sky130_fd_sc_hd__buf_2
X_68836_ _68822_/Y _68823_/X _68824_/X _68835_/Y _68836_/X sky130_fd_sc_hd__a211o_4
X_87670_ _87671_/CLK _42883_/Y _87670_/Q sky130_fd_sc_hd__dfxtp_4
X_84882_ _84921_/CLK _84882_/D _84882_/Q sky130_fd_sc_hd__dfxtp_4
X_55801_ _55801_/A _55801_/B _55801_/C _55801_/D _55802_/A sky130_fd_sc_hd__and4_4
X_86621_ _85981_/CLK _47569_/Y _86621_/Q sky130_fd_sc_hd__dfxtp_4
X_83833_ _83191_/CLK _83833_/D _83833_/Q sky130_fd_sc_hd__dfxtp_4
X_56781_ _56780_/X _85133_/D sky130_fd_sc_hd__inv_2
X_68767_ _80818_/D _68713_/X _68766_/X _83962_/D sky130_fd_sc_hd__a21bo_4
X_53993_ _53978_/A _53993_/B _53993_/Y sky130_fd_sc_hd__nand2_4
X_65979_ _65973_/X _65978_/X _65880_/X _65983_/A sky130_fd_sc_hd__a21o_4
X_58520_ _58520_/A _58510_/X _58520_/Y sky130_fd_sc_hd__nor2_4
X_55732_ _55235_/A _55732_/B _55732_/X sky130_fd_sc_hd__and2_4
X_67718_ _67359_/X _67718_/X sky130_fd_sc_hd__buf_2
X_86552_ _85915_/CLK _86552_/D _66041_/B sky130_fd_sc_hd__dfxtp_4
X_52944_ _52944_/A _52944_/B _52944_/Y sky130_fd_sc_hd__nand2_4
X_83764_ _83482_/CLK _83764_/D _83764_/Q sky130_fd_sc_hd__dfxtp_4
X_80976_ _82084_/CLK _80976_/D _80932_/D sky130_fd_sc_hd__dfxtp_4
X_68698_ _68694_/X _68696_/X _68697_/X _68698_/X sky130_fd_sc_hd__a21o_4
X_85503_ _85505_/CLK _85503_/D _85503_/Q sky130_fd_sc_hd__dfxtp_4
X_58451_ _58984_/A _58498_/B sky130_fd_sc_hd__buf_2
X_82715_ _82715_/CLK _79035_/X _82671_/D sky130_fd_sc_hd__dfxtp_4
X_55663_ _83317_/Q _55663_/Y sky130_fd_sc_hd__inv_2
X_67649_ _67649_/A _67649_/B _67649_/Y sky130_fd_sc_hd__nand2_4
X_86483_ _86193_/CLK _48787_/Y _86483_/Q sky130_fd_sc_hd__dfxtp_4
X_52875_ _52767_/A _52885_/A sky130_fd_sc_hd__buf_2
X_83695_ _83699_/CLK _83695_/D _83695_/Q sky130_fd_sc_hd__dfxtp_4
X_57402_ _56626_/X _57391_/Y _57401_/Y _85015_/D sky130_fd_sc_hd__a21oi_4
X_88222_ _88232_/CLK _88222_/D _67848_/B sky130_fd_sc_hd__dfxtp_4
X_54614_ _54600_/A _47221_/A _54614_/Y sky130_fd_sc_hd__nand2_4
X_85434_ _85433_/CLK _54484_/Y _85434_/Q sky130_fd_sc_hd__dfxtp_4
X_51826_ _51820_/A _50961_/B _51826_/Y sky130_fd_sc_hd__nand2_4
X_70660_ _70423_/X _70886_/A sky130_fd_sc_hd__buf_2
X_82646_ _82648_/CLK _83998_/Q _82646_/Q sky130_fd_sc_hd__dfxtp_4
X_58382_ _58382_/A _58383_/A sky130_fd_sc_hd__inv_2
X_55594_ _55572_/X _45438_/Y _55594_/Y sky130_fd_sc_hd__nor2_4
X_57333_ _56732_/X _57290_/A _57332_/Y _57333_/X sky130_fd_sc_hd__o21a_4
X_69319_ _87526_/Q _69261_/X _69248_/X _69318_/X _69319_/X sky130_fd_sc_hd__a211o_4
X_88153_ _87141_/CLK _88153_/D _88153_/Q sky130_fd_sc_hd__dfxtp_4
X_54545_ _54543_/Y _54530_/X _54544_/X _54545_/Y sky130_fd_sc_hd__a21oi_4
X_85365_ _83630_/CLK _54858_/Y _85365_/Q sky130_fd_sc_hd__dfxtp_4
X_51757_ _51753_/Y _51391_/X _51756_/X _85952_/D sky130_fd_sc_hd__a21oi_4
X_70591_ _70591_/A _74533_/D sky130_fd_sc_hd__buf_2
X_82577_ _82702_/CLK _82609_/Q _78183_/A sky130_fd_sc_hd__dfxtp_4
X_87104_ _87110_/CLK _87104_/D _87104_/Q sky130_fd_sc_hd__dfxtp_4
X_41510_ _41481_/X _82327_/Q _41509_/X _41510_/Y sky130_fd_sc_hd__o21ai_4
X_72330_ _72326_/Y _72329_/Y _72292_/X _72330_/X sky130_fd_sc_hd__a21o_4
X_84316_ _84314_/CLK _63531_/Y _84316_/Q sky130_fd_sc_hd__dfxtp_4
X_50708_ _50738_/A _50708_/B _50708_/Y sky130_fd_sc_hd__nand2_4
X_57264_ _45947_/B _56971_/B _56899_/Y _57264_/Y sky130_fd_sc_hd__nor3_4
X_81528_ _84014_/CLK _81528_/D _81528_/Q sky130_fd_sc_hd__dfxtp_4
X_88084_ _88084_/CLK _88084_/D _88084_/Q sky130_fd_sc_hd__dfxtp_4
X_42490_ _42486_/X _42472_/X _40650_/X _68641_/B _42489_/X _42490_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54476_ _54453_/X _54471_/B _54471_/C _46979_/Y _54476_/X sky130_fd_sc_hd__and4_4
X_85296_ _85279_/CLK _85296_/D _85296_/Q sky130_fd_sc_hd__dfxtp_4
X_51688_ _51608_/A _51695_/C sky130_fd_sc_hd__buf_2
X_59003_ _59001_/X _86081_/Q _59002_/X _59003_/Y sky130_fd_sc_hd__o21ai_4
X_56215_ _56188_/X _56050_/X _56214_/Y _56215_/Y sky130_fd_sc_hd__o21ai_4
X_87035_ _87333_/CLK _87035_/D _87035_/Q sky130_fd_sc_hd__dfxtp_4
X_41441_ _41421_/X _82884_/Q _41440_/X _41441_/X sky130_fd_sc_hd__o21a_4
X_53427_ _85635_/Q _53404_/X _53426_/Y _53427_/Y sky130_fd_sc_hd__o21ai_4
X_72261_ _72257_/Y _72260_/Y _72201_/X _72261_/X sky130_fd_sc_hd__a21o_4
X_84247_ _84849_/CLK _84247_/D _79691_/B sky130_fd_sc_hd__dfxtp_4
X_50639_ _50718_/A _50640_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_1 _44265_/Y _44267_/A sky130_fd_sc_hd__buf_8
X_57195_ _57195_/A _57195_/B _57195_/C _57195_/Y sky130_fd_sc_hd__nand3_4
X_81459_ _81461_/CLK _76809_/B _81459_/Q sky130_fd_sc_hd__dfxtp_4
X_74000_ _74000_/A _73999_/X _74001_/B sky130_fd_sc_hd__nand2_4
X_71212_ _50508_/B _71190_/A _71211_/Y _71212_/Y sky130_fd_sc_hd__o21ai_4
X_44160_ _44160_/A _44160_/B _44160_/Y sky130_fd_sc_hd__nand2_4
X_56146_ _56142_/X _56144_/X _56145_/Y _85288_/D sky130_fd_sc_hd__o21ai_4
X_41372_ _41371_/X _41362_/X _67732_/B _41363_/X _88227_/D sky130_fd_sc_hd__a2bb2o_4
X_53358_ _53339_/A _53371_/B _53371_/C _52841_/D _53358_/X sky130_fd_sc_hd__and4_4
X_72192_ _72277_/A _72192_/B _72192_/Y sky130_fd_sc_hd__nor2_4
X_84178_ _84175_/CLK _84178_/D _84178_/Q sky130_fd_sc_hd__dfxtp_4
X_43111_ _43100_/X _43110_/X _40762_/X _74266_/A _43080_/X _43112_/A
+ sky130_fd_sc_hd__o32ai_4
X_40323_ _48135_/A _49140_/B sky130_fd_sc_hd__buf_2
X_52309_ _52309_/A _52310_/B sky130_fd_sc_hd__buf_2
X_71143_ _71171_/A _71141_/B _71152_/C _70875_/X _71143_/Y sky130_fd_sc_hd__nand4_4
X_83129_ _83561_/CLK _83129_/D _70115_/A sky130_fd_sc_hd__dfxtp_4
X_44091_ _44052_/X _44068_/Y _44071_/X _44085_/Y _44090_/Y _44091_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56077_ _56058_/X _56074_/X _56076_/Y _85300_/D sky130_fd_sc_hd__o21ai_4
X_53289_ _53287_/Y _53272_/X _53288_/X _53289_/Y sky130_fd_sc_hd__a21oi_4
X_43042_ _42060_/X _43031_/X _40617_/X _43041_/Y _43034_/X _87597_/D
+ sky130_fd_sc_hd__o32ai_4
X_55028_ _55037_/A _54859_/B _55028_/Y sky130_fd_sc_hd__nand2_4
X_59905_ _59570_/A _59905_/B _61070_/B sky130_fd_sc_hd__nor2_4
X_71074_ _48963_/X _71070_/X _71073_/Y _71074_/Y sky130_fd_sc_hd__o21ai_4
X_75951_ _75957_/A _75957_/B _75954_/A sky130_fd_sc_hd__xor2_4
X_87937_ _82888_/CLK _42292_/X _87937_/Q sky130_fd_sc_hd__dfxtp_4
X_74902_ _81129_/D _74891_/B _74901_/X _74902_/Y sky130_fd_sc_hd__a21oi_4
X_70025_ _82550_/D _70010_/X _70024_/X _83870_/D sky130_fd_sc_hd__a21bo_4
X_47850_ _46578_/X _46265_/A _47849_/X _47851_/B sky130_fd_sc_hd__o21ai_4
X_59836_ _59689_/B _59731_/Y _59631_/B _59836_/D _59836_/Y sky130_fd_sc_hd__nand4_4
X_78670_ _78669_/X _78701_/B sky130_fd_sc_hd__buf_2
X_75882_ _75726_/Y _80787_/D sky130_fd_sc_hd__inv_2
X_87868_ _82899_/CLK _42428_/X _87868_/Q sky130_fd_sc_hd__dfxtp_4
X_46801_ _46800_/Y _52681_/D sky130_fd_sc_hd__buf_2
X_77621_ _77621_/A _77627_/A sky130_fd_sc_hd__inv_2
X_74833_ _74832_/Y _74833_/Y sky130_fd_sc_hd__inv_2
X_86819_ _87077_/CLK _86819_/D _67023_/B sky130_fd_sc_hd__dfxtp_4
X_47781_ _47799_/A _53240_/B _47781_/Y sky130_fd_sc_hd__nand2_4
X_59767_ _59766_/X _61770_/D sky130_fd_sc_hd__buf_2
X_44993_ _56670_/A _45835_/A sky130_fd_sc_hd__buf_2
X_56979_ _45643_/Y _56671_/X _56979_/Y sky130_fd_sc_hd__nand2_4
X_87799_ _87544_/CLK _42619_/Y _69929_/A sky130_fd_sc_hd__dfxtp_4
X_49520_ _49520_/A _49548_/A sky130_fd_sc_hd__buf_2
X_46732_ _54332_/B _51812_/B sky130_fd_sc_hd__buf_2
X_58718_ _58667_/X _86101_/Q _58717_/X _58718_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_140_0_CLK clkbuf_8_70_0_CLK/X clkbuf_9_140_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_77552_ _77552_/A _77552_/Y sky130_fd_sc_hd__inv_2
X_43944_ _43944_/A _43987_/B sky130_fd_sc_hd__buf_2
X_74764_ _74764_/A _74764_/B _71010_/X _70732_/X _74764_/X sky130_fd_sc_hd__and4_4
X_71976_ _71957_/A _48920_/Y _71976_/Y sky130_fd_sc_hd__nand2_4
X_59698_ _59605_/Y _59722_/A sky130_fd_sc_hd__buf_2
X_76503_ _76503_/A _81542_/Q _76503_/Y sky130_fd_sc_hd__nand2_4
X_49451_ _49451_/A _49456_/B sky130_fd_sc_hd__buf_2
X_73715_ _73665_/X _84987_/Q _73614_/X _73714_/X _73715_/X sky130_fd_sc_hd__a211o_4
X_70927_ _51043_/B _70909_/A _70926_/Y _70927_/Y sky130_fd_sc_hd__o21ai_4
X_46663_ _46651_/A _46662_/X _46663_/Y sky130_fd_sc_hd__nand2_4
X_58649_ _58649_/A _58649_/B _58649_/Y sky130_fd_sc_hd__nor2_4
X_77483_ _77454_/X _77458_/B _77482_/Y _77484_/B sky130_fd_sc_hd__o21a_4
X_43875_ _41272_/X _43868_/X _87222_/Q _43870_/X _87222_/D sky130_fd_sc_hd__a2bb2o_4
X_74695_ _56886_/B _74656_/X _74694_/Y _74695_/X sky130_fd_sc_hd__a21bo_4
Xclkbuf_10_664_0_CLK clkbuf_9_332_0_CLK/X _82629_/CLK sky130_fd_sc_hd__clkbuf_1
X_48402_ _86525_/Q _48333_/X _48401_/Y _48402_/Y sky130_fd_sc_hd__o21ai_4
X_79222_ _79217_/Y _79218_/X _79221_/Y _79224_/A sky130_fd_sc_hd__a21o_4
X_45614_ _55470_/B _45596_/X _45548_/X _45613_/Y _45614_/X sky130_fd_sc_hd__a211o_4
X_76434_ _76419_/Y _76422_/Y _76417_/Y _76435_/B sky130_fd_sc_hd__o21ai_4
X_42826_ _41465_/X _42821_/X _87698_/Q _42822_/X _42826_/X sky130_fd_sc_hd__a2bb2o_4
X_49382_ _49382_/A _51770_/B _49382_/Y sky130_fd_sc_hd__nand2_4
X_61660_ _61476_/A _61690_/B sky130_fd_sc_hd__buf_2
X_73646_ _73644_/X _73646_/B _73635_/X _73646_/Y sky130_fd_sc_hd__nand3_4
X_46594_ _83778_/Q _52571_/B sky130_fd_sc_hd__inv_2
X_70858_ _71072_/A _71088_/C sky130_fd_sc_hd__buf_2
Xclkbuf_9_155_0_CLK clkbuf_8_77_0_CLK/X clkbuf_9_155_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_48333_ _48548_/A _48333_/X sky130_fd_sc_hd__buf_2
X_60611_ _60376_/X _60532_/A _60571_/Y _60609_/X _60610_/X _60611_/X
+ sky130_fd_sc_hd__o41a_4
X_79153_ _79153_/A _79153_/B _79153_/X sky130_fd_sc_hd__xor2_4
X_45545_ _45511_/X _61440_/A _45530_/X _45545_/Y sky130_fd_sc_hd__o21ai_4
X_76365_ _76365_/A _76369_/A sky130_fd_sc_hd__inv_2
Xclkbuf_9_82_0_CLK clkbuf_9_83_0_CLK/A clkbuf_9_82_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_42757_ _42745_/A _42757_/X sky130_fd_sc_hd__buf_2
X_61591_ _84859_/Q _61593_/B sky130_fd_sc_hd__buf_2
X_73577_ _73577_/A _73577_/B _73577_/Y sky130_fd_sc_hd__nor2_4
X_70789_ _70400_/A _70790_/A sky130_fd_sc_hd__buf_2
X_78104_ _82565_/Q _78103_/B _78104_/Y sky130_fd_sc_hd__nand2_4
X_63330_ _59439_/Y _63259_/X _60523_/A _58987_/Y _63060_/A _63330_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75316_ _75315_/Y _75319_/B sky130_fd_sc_hd__inv_2
X_41708_ _82898_/Q _41653_/X _41708_/X sky130_fd_sc_hd__or2_4
X_60542_ _60566_/A _60476_/A _60488_/C _60542_/Y sky130_fd_sc_hd__nand3_4
X_48264_ _48163_/X _48264_/X sky130_fd_sc_hd__buf_2
X_72528_ _72528_/A _72528_/Y sky130_fd_sc_hd__inv_2
X_79084_ _79084_/A _79083_/Y _82719_/D sky130_fd_sc_hd__nand2_4
X_45476_ _85052_/Q _45490_/B _45476_/Y sky130_fd_sc_hd__nor2_4
X_76296_ _76296_/A _76295_/Y _76297_/B sky130_fd_sc_hd__xor2_4
X_42688_ _42592_/A _42688_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_679_0_CLK clkbuf_9_339_0_CLK/X _86920_/CLK sky130_fd_sc_hd__clkbuf_1
X_47215_ _59377_/A _47192_/X _47214_/Y _47215_/Y sky130_fd_sc_hd__o21ai_4
X_78035_ _78033_/Y _78034_/Y _78037_/A sky130_fd_sc_hd__nand2_4
X_44427_ _44548_/A _44427_/X sky130_fd_sc_hd__buf_2
X_63261_ _63288_/A _64466_/B _63312_/C _63237_/X _63261_/X sky130_fd_sc_hd__and4_4
X_75247_ _75233_/X _75245_/Y _75246_/Y _75247_/X sky130_fd_sc_hd__a21o_4
X_41639_ _41457_/A _41639_/X sky130_fd_sc_hd__buf_2
X_48195_ _52309_/A _48195_/X sky130_fd_sc_hd__buf_2
X_60473_ _60421_/B _60473_/B _60473_/C _60438_/A _60556_/B sky130_fd_sc_hd__nand4_4
X_72459_ _72327_/X _85956_/Q _72458_/X _72459_/Y sky130_fd_sc_hd__o21ai_4
X_65000_ _64929_/A _65000_/B _65000_/X sky130_fd_sc_hd__and2_4
X_62212_ _62212_/A _62202_/Y _62206_/Y _62211_/Y _62212_/Y sky130_fd_sc_hd__nand4_4
X_47146_ _57563_/A _47147_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_97_0_CLK clkbuf_9_97_0_CLK/A clkbuf_9_97_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_44358_ _41727_/X _44345_/X _87149_/Q _44346_/X _44358_/X sky130_fd_sc_hd__a2bb2o_4
X_63192_ _63154_/X _64401_/B _63165_/X _63192_/D _63192_/X sky130_fd_sc_hd__and4_4
X_75178_ _75178_/A _75178_/B _75178_/C _75179_/A sky130_fd_sc_hd__nand3_4
Xclkbuf_10_602_0_CLK clkbuf_9_301_0_CLK/X _81990_/CLK sky130_fd_sc_hd__clkbuf_1
X_43309_ _43296_/X _43305_/X _41214_/X _87488_/Q _43308_/X _43309_/Y
+ sky130_fd_sc_hd__o32ai_4
X_62143_ _62135_/X _62137_/X _62142_/Y _84870_/Q _62117_/X _62143_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74129_ _74152_/A _74129_/B _74129_/X sky130_fd_sc_hd__and2_4
X_47077_ _47077_/A _53360_/B sky130_fd_sc_hd__inv_2
X_44289_ _44284_/Y _44285_/Y _44288_/X _44289_/X sky130_fd_sc_hd__o21a_4
X_79986_ _79972_/Y _79973_/Y _79985_/Y _79988_/A sky130_fd_sc_hd__a21o_4
X_46028_ _41464_/Y _46022_/X _86805_/Q _46023_/X _86805_/D sky130_fd_sc_hd__a2bb2o_4
X_66951_ _87363_/Q _66878_/X _66879_/X _66950_/X _66951_/X sky130_fd_sc_hd__a211o_4
X_62074_ _61590_/B _61995_/X _62010_/X _62011_/X _62077_/C sky130_fd_sc_hd__nand4_4
X_78937_ _78937_/A _78937_/B _78952_/A sky130_fd_sc_hd__nand2_4
Xclkbuf_9_20_0_CLK clkbuf_8_10_0_CLK/X clkbuf_9_20_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_65902_ _65899_/Y _65830_/X _65901_/X _84170_/D sky130_fd_sc_hd__a21o_4
X_61025_ _60994_/A _60994_/B _60951_/Y _61025_/X sky130_fd_sc_hd__a21o_4
X_69670_ _69579_/X _69668_/Y _69604_/X _69669_/Y _69670_/X sky130_fd_sc_hd__a211o_4
X_66882_ _66877_/X _66881_/X _66787_/X _66886_/A sky130_fd_sc_hd__a21o_4
X_78868_ _78868_/A _78867_/Y _78869_/B sky130_fd_sc_hd__xor2_4
Xclkbuf_10_617_0_CLK clkbuf_9_308_0_CLK/X _81179_/CLK sky130_fd_sc_hd__clkbuf_1
X_68621_ _69004_/A _88361_/Q _68621_/X sky130_fd_sc_hd__and2_4
X_65833_ _65317_/X _65833_/B _65320_/X _65833_/Y sky130_fd_sc_hd__nand3_4
X_77819_ _77819_/A _77819_/Y sky130_fd_sc_hd__inv_2
X_47979_ _47988_/A _50302_/B _47979_/Y sky130_fd_sc_hd__nand2_4
X_78799_ _82785_/D _78799_/B _78801_/A sky130_fd_sc_hd__nand2_4
Xclkbuf_9_108_0_CLK clkbuf_8_54_0_CLK/X clkbuf_9_108_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_49718_ _57721_/B _49715_/X _49717_/Y _49718_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_35_0_CLK clkbuf_9_35_0_CLK/A clkbuf_9_35_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_80830_ _83944_/CLK _83974_/Q _75677_/B sky130_fd_sc_hd__dfxtp_4
X_68552_ _66540_/A _68552_/X sky130_fd_sc_hd__buf_2
X_65764_ _65654_/X _86187_/Q _65761_/X _65763_/X _65764_/X sky130_fd_sc_hd__a211o_4
X_50990_ _50988_/Y _50983_/X _50989_/X _50990_/Y sky130_fd_sc_hd__a21oi_4
X_62976_ _62972_/Y _62642_/B _62973_/Y _62974_/Y _62975_/X _62976_/X
+ sky130_fd_sc_hd__a41o_4
X_67503_ _67498_/X _67501_/X _67502_/X _67506_/A sky130_fd_sc_hd__a21o_4
X_64715_ _64565_/A _65790_/A sky130_fd_sc_hd__buf_2
X_61927_ _61960_/A _61960_/B _78068_/B _61927_/Y sky130_fd_sc_hd__nor3_4
X_49649_ _59256_/B _49632_/X _49648_/Y _49649_/Y sky130_fd_sc_hd__o21ai_4
X_80761_ _80968_/CLK _80761_/D _81137_/D sky130_fd_sc_hd__dfxtp_4
X_68483_ _87503_/Q _68365_/X _68450_/X _68482_/X _68483_/X sky130_fd_sc_hd__a211o_4
X_65695_ _65063_/X _65828_/B _65067_/X _65695_/Y sky130_fd_sc_hd__nand3_4
X_82500_ _82942_/CLK _79124_/Y _78341_/A sky130_fd_sc_hd__dfxtp_4
X_67434_ _67364_/X _67434_/B _67434_/X sky130_fd_sc_hd__and2_4
X_52660_ _52605_/A _52661_/B sky130_fd_sc_hd__buf_2
X_64646_ _64923_/A _64773_/A sky130_fd_sc_hd__buf_2
X_83480_ _83480_/CLK _83480_/D _83480_/Q sky130_fd_sc_hd__dfxtp_4
X_61858_ _61708_/X _61860_/C sky130_fd_sc_hd__buf_2
X_80692_ _81104_/CLK _80692_/D _80692_/Q sky130_fd_sc_hd__dfxtp_4
X_51611_ _51617_/A _53135_/B _51611_/Y sky130_fd_sc_hd__nand2_4
X_82431_ _83167_/CLK _82463_/Q _78750_/A sky130_fd_sc_hd__dfxtp_4
X_60809_ _60765_/Y _60809_/Y sky130_fd_sc_hd__inv_2
X_67365_ _67364_/X _67365_/B _67365_/X sky130_fd_sc_hd__and2_4
X_64577_ _64797_/A _64577_/X sky130_fd_sc_hd__buf_2
X_52591_ _85790_/Q _52575_/X _52590_/Y _52591_/Y sky130_fd_sc_hd__o21ai_4
X_61789_ _61770_/A _61823_/B _63410_/B _61788_/X _61789_/X sky130_fd_sc_hd__and4_4
XPHY_708 sky130_fd_sc_hd__decap_3
X_69104_ _69059_/A _69104_/B _69104_/X sky130_fd_sc_hd__and2_4
X_54330_ _54325_/A _54353_/B _54317_/X _46727_/Y _54330_/X sky130_fd_sc_hd__and4_4
X_66316_ _65850_/X _66276_/B _65852_/X _66316_/Y sky130_fd_sc_hd__nand3_4
X_85150_ _85152_/CLK _85150_/D _55599_/B sky130_fd_sc_hd__dfxtp_4
X_51542_ _85991_/Q _51539_/X _51541_/Y _51542_/Y sky130_fd_sc_hd__o21ai_4
X_63528_ _63528_/A _63554_/A sky130_fd_sc_hd__buf_2
X_82362_ _84980_/CLK _77232_/Y _82362_/Q sky130_fd_sc_hd__dfxtp_4
X_67296_ _67250_/A _67296_/B _67296_/X sky130_fd_sc_hd__and2_4
X_84101_ _80928_/CLK _66687_/X _84101_/Q sky130_fd_sc_hd__dfxtp_4
X_81313_ _81801_/CLK _77001_/X _81313_/Q sky130_fd_sc_hd__dfxtp_4
X_69035_ _69035_/A _69035_/X sky130_fd_sc_hd__buf_2
X_54261_ _54961_/A _53095_/B _54261_/Y sky130_fd_sc_hd__nand2_4
X_66247_ _66231_/X _66151_/B _66247_/C _66247_/X sky130_fd_sc_hd__and3_4
X_85081_ _85089_/CLK _85081_/D _57113_/B sky130_fd_sc_hd__dfxtp_4
X_51473_ _51473_/A _51473_/B _51494_/C _52997_/D _51473_/X sky130_fd_sc_hd__and4_4
X_63459_ _63448_/A _63459_/B _63458_/X _63410_/D _63459_/X sky130_fd_sc_hd__and4_4
X_82293_ _82103_/CLK _82293_/D _82293_/Q sky130_fd_sc_hd__dfxtp_4
X_56000_ _55999_/X _56001_/A sky130_fd_sc_hd__buf_2
X_53212_ _53210_/Y _53189_/X _53211_/X _85676_/D sky130_fd_sc_hd__a21oi_4
X_84032_ _81160_/CLK _68127_/X _82072_/D sky130_fd_sc_hd__dfxtp_4
X_50424_ _86203_/Q _50403_/X _50423_/Y _50424_/Y sky130_fd_sc_hd__o21ai_4
X_81244_ _85372_/CLK _81052_/Q _81244_/Q sky130_fd_sc_hd__dfxtp_4
X_54192_ _54189_/Y _54171_/X _54191_/X _54192_/Y sky130_fd_sc_hd__a21oi_4
X_66178_ _66174_/Y _66137_/X _66177_/Y _84151_/D sky130_fd_sc_hd__a21o_4
X_53143_ _53195_/A _53143_/X sky130_fd_sc_hd__buf_2
X_65129_ _65791_/A _65155_/A sky130_fd_sc_hd__buf_2
X_50355_ _86217_/Q _50316_/X _50354_/Y _50355_/Y sky130_fd_sc_hd__o21ai_4
X_81175_ _82335_/CLK _74998_/B _81175_/Q sky130_fd_sc_hd__dfxtp_4
Xpsn_inst_psn_buff_30 _40351_/Y _47002_/A sky130_fd_sc_hd__buf_8
X_80126_ _80122_/X _80125_/Y _80126_/X sky130_fd_sc_hd__xor2_4
X_53074_ _53074_/A _53069_/X _53074_/C _53074_/D _53074_/X sky130_fd_sc_hd__and4_4
X_57951_ _57946_/Y _57950_/Y _57889_/X _57951_/X sky130_fd_sc_hd__a21o_4
X_69937_ _69937_/A _69937_/B _69937_/Y sky130_fd_sc_hd__nand2_4
X_50286_ _86231_/Q _50282_/X _50285_/Y _50286_/Y sky130_fd_sc_hd__o21ai_4
X_85983_ _85697_/CLK _85983_/D _85983_/Q sky130_fd_sc_hd__dfxtp_4
X_52025_ _52058_/A _50322_/B _52025_/Y sky130_fd_sc_hd__nand2_4
X_56902_ _55657_/Y _56688_/X _56902_/Y sky130_fd_sc_hd__nand2_4
X_87722_ _87708_/CLK _87722_/D _87722_/Q sky130_fd_sc_hd__dfxtp_4
X_84934_ _85381_/CLK _84934_/D _84934_/Q sky130_fd_sc_hd__dfxtp_4
X_80057_ _80048_/X _80057_/B _80057_/Y sky130_fd_sc_hd__nand2_4
X_57882_ _84943_/Q _57819_/X _57873_/X _57881_/X _84943_/D sky130_fd_sc_hd__a2bb2oi_4
X_69868_ _69448_/Y _69732_/X _69815_/X _69867_/Y _69868_/X sky130_fd_sc_hd__a211o_4
X_59621_ _61276_/B _59639_/A _59640_/A _60175_/A _59621_/X sky130_fd_sc_hd__and4_4
X_56833_ _56832_/X _55681_/X _56777_/B _56833_/Y sky130_fd_sc_hd__o21ai_4
X_68819_ _64980_/A _68819_/X sky130_fd_sc_hd__buf_2
X_87653_ _87653_/CLK _87653_/D _67675_/B sky130_fd_sc_hd__dfxtp_4
X_84865_ _84344_/CLK _84865_/D _84865_/Q sky130_fd_sc_hd__dfxtp_4
X_69799_ _87054_/Q _69796_/X _69797_/X _69798_/X _69800_/B sky130_fd_sc_hd__a211o_4
X_86604_ _85962_/CLK _86604_/D _72378_/A sky130_fd_sc_hd__dfxtp_4
X_71830_ _71714_/Y _71839_/B sky130_fd_sc_hd__buf_2
X_59552_ _60407_/A _59552_/B _59552_/C _60407_/C _59552_/Y sky130_fd_sc_hd__nand4_4
X_83816_ _83813_/CLK _83816_/D _74801_/B sky130_fd_sc_hd__dfxtp_4
X_56764_ _59498_/A _56764_/B _56764_/C _56764_/D _56764_/Y sky130_fd_sc_hd__nand4_4
X_87584_ _87595_/CLK _43079_/Y _87584_/Q sky130_fd_sc_hd__dfxtp_4
X_53976_ _53956_/X _53976_/B _53976_/Y sky130_fd_sc_hd__nand2_4
X_41990_ _41960_/X _41951_/X _40787_/X _72855_/A _41953_/X _41990_/Y
+ sky130_fd_sc_hd__o32ai_4
X_84796_ _86701_/CLK _84796_/D _84796_/Q sky130_fd_sc_hd__dfxtp_4
X_58503_ _58492_/X _58500_/Y _58502_/Y _58503_/Y sky130_fd_sc_hd__a21oi_4
X_55715_ _55245_/A _55715_/B _55715_/X sky130_fd_sc_hd__and2_4
X_86535_ _86535_/CLK _48326_/Y _74177_/B sky130_fd_sc_hd__dfxtp_4
X_40941_ _40941_/A _40941_/X sky130_fd_sc_hd__buf_2
X_52927_ _52922_/A _52916_/B _52926_/X _52927_/D _52927_/X sky130_fd_sc_hd__and4_4
X_71761_ _71761_/A _71761_/Y sky130_fd_sc_hd__inv_2
X_83747_ _83753_/CLK _83747_/D _83747_/Q sky130_fd_sc_hd__dfxtp_4
X_59483_ _58517_/X _59480_/Y _59482_/Y _84720_/D sky130_fd_sc_hd__a21oi_4
X_56695_ _56694_/Y _56696_/A sky130_fd_sc_hd__buf_2
X_80959_ _81994_/CLK _80959_/D _80959_/Q sky130_fd_sc_hd__dfxtp_4
X_73500_ _73386_/A _86500_/Q _73500_/X sky130_fd_sc_hd__and2_4
X_70712_ _70712_/A _70848_/A sky130_fd_sc_hd__buf_2
X_58434_ _58434_/A _58426_/X _58434_/Y sky130_fd_sc_hd__nand2_4
X_43660_ _43660_/A _68959_/B sky130_fd_sc_hd__inv_2
X_55646_ _55646_/A _55646_/X sky130_fd_sc_hd__buf_2
X_74480_ _74490_/A _48627_/A _74480_/Y sky130_fd_sc_hd__nand2_4
X_86466_ _83310_/CLK _86466_/D _86466_/Q sky130_fd_sc_hd__dfxtp_4
X_40872_ _82861_/Q _40883_/B _40872_/X sky130_fd_sc_hd__or2_4
X_52858_ _52856_/Y _52839_/X _52857_/X _52858_/Y sky130_fd_sc_hd__a21oi_4
X_71692_ _71319_/B _71874_/D sky130_fd_sc_hd__buf_2
X_83678_ _86104_/CLK _70870_/Y _46721_/A sky130_fd_sc_hd__dfxtp_4
X_88205_ _87436_/CLK _88205_/D _66718_/B sky130_fd_sc_hd__dfxtp_4
X_42611_ _73415_/A _42611_/Y sky130_fd_sc_hd__inv_2
X_73431_ _73428_/X _73430_/X _73432_/B sky130_fd_sc_hd__nand2_4
X_85417_ _85735_/CLK _54577_/Y _85417_/Q sky130_fd_sc_hd__dfxtp_4
X_51809_ _51781_/A _51810_/C sky130_fd_sc_hd__buf_2
X_70643_ _70710_/A _70639_/B _70642_/X _70638_/X _70643_/Y sky130_fd_sc_hd__nand4_4
X_58365_ _58328_/X _83764_/Q _58364_/Y _58365_/X sky130_fd_sc_hd__o21a_4
X_82629_ _82629_/CLK _82629_/D _82629_/Q sky130_fd_sc_hd__dfxtp_4
X_43591_ _43591_/A _43605_/A sky130_fd_sc_hd__buf_2
X_55577_ _55574_/X _55576_/X _55517_/X _55580_/A sky130_fd_sc_hd__a21o_4
X_86397_ _84807_/CLK _86397_/D _58613_/B sky130_fd_sc_hd__dfxtp_4
X_52789_ _52708_/A _52789_/X sky130_fd_sc_hd__buf_2
X_45330_ _85285_/Q _45269_/X _45303_/X _45330_/X sky130_fd_sc_hd__o21a_4
X_57316_ _57280_/X _57312_/Y _57313_/Y _57315_/Y _57317_/A sky130_fd_sc_hd__a211o_4
X_88136_ _88133_/CLK _88136_/D _66845_/B sky130_fd_sc_hd__dfxtp_4
X_76150_ _76150_/A _76150_/B _76150_/X sky130_fd_sc_hd__and2_4
X_42542_ _42542_/A _87828_/D sky130_fd_sc_hd__inv_2
X_54528_ _54518_/A _53353_/B _54528_/Y sky130_fd_sc_hd__nand2_4
X_73362_ _73362_/A _73361_/X _73363_/B sky130_fd_sc_hd__nand2_4
X_85348_ _85346_/CLK _85348_/D _85348_/Q sky130_fd_sc_hd__dfxtp_4
X_70574_ _70532_/Y _83746_/Q _70573_/Y _83746_/D sky130_fd_sc_hd__a21o_4
X_58296_ _58296_/A _58248_/B _58296_/Y sky130_fd_sc_hd__nor2_4
X_75101_ _75096_/A _75099_/Y _75100_/Y _75104_/B sky130_fd_sc_hd__o21ai_4
X_72313_ _72313_/A _72313_/Y sky130_fd_sc_hd__inv_2
X_45261_ _45202_/X _61607_/B _45219_/X _45261_/Y sky130_fd_sc_hd__o21ai_4
X_57247_ _57244_/X _57247_/Y sky130_fd_sc_hd__inv_2
X_76081_ _76077_/Y _76080_/X _76081_/Y sky130_fd_sc_hd__nand2_4
X_88067_ _87553_/CLK _42023_/Y _73175_/A sky130_fd_sc_hd__dfxtp_4
X_42473_ _73699_/A _68520_/B sky130_fd_sc_hd__inv_2
X_54459_ _54486_/A _54478_/A sky130_fd_sc_hd__buf_2
X_73293_ _73291_/X _73277_/X _73281_/Y _73293_/Y sky130_fd_sc_hd__nand3_4
X_85279_ _85279_/CLK _85279_/D _56198_/C sky130_fd_sc_hd__dfxtp_4
X_47000_ _46981_/A _47029_/B _47029_/C _52797_/D _47000_/X sky130_fd_sc_hd__and4_4
X_44212_ _44196_/X _57019_/A sky130_fd_sc_hd__inv_2
X_75032_ _81147_/D _75032_/B _75032_/Y sky130_fd_sc_hd__nand2_4
X_87018_ _87026_/CLK _44647_/Y _87018_/Q sky130_fd_sc_hd__dfxtp_4
X_41424_ _41423_/X _41424_/X sky130_fd_sc_hd__buf_2
X_72244_ _72239_/Y _72243_/Y _72185_/X _72244_/X sky130_fd_sc_hd__a21o_4
X_45192_ _45188_/Y _45191_/Y _45137_/X _45192_/X sky130_fd_sc_hd__a21o_4
X_57178_ _56801_/X _57141_/X _57177_/Y _57178_/Y sky130_fd_sc_hd__o21ai_4
X_44143_ _44139_/X _44141_/X _44025_/X _44142_/X _44143_/Y sky130_fd_sc_hd__nand4_4
X_56129_ _55801_/C _56128_/Y _56130_/A sky130_fd_sc_hd__xor2_4
X_79840_ _79840_/A _79827_/Y _79840_/X sky130_fd_sc_hd__or2_4
X_41355_ _41261_/X _41699_/B _41354_/X _41355_/Y sky130_fd_sc_hd__o21ai_4
X_72175_ _86621_/Q _72162_/B _72175_/Y sky130_fd_sc_hd__nor2_4
X_71126_ _50188_/B _71117_/X _71125_/Y _71126_/Y sky130_fd_sc_hd__o21ai_4
X_48951_ _48945_/Y _48935_/X _48950_/X _86459_/D sky130_fd_sc_hd__a21oi_4
X_44074_ _55129_/A _55741_/A sky130_fd_sc_hd__buf_2
X_79771_ _79766_/X _79770_/Y _79771_/X sky130_fd_sc_hd__xor2_4
X_41286_ _41286_/A _41280_/B _41286_/X sky130_fd_sc_hd__or2_4
X_76983_ _76983_/A _62485_/C _76983_/X sky130_fd_sc_hd__xor2_4
X_47902_ _73711_/B _47897_/X _47901_/Y _47902_/Y sky130_fd_sc_hd__o21ai_4
X_43025_ _43127_/A _43025_/X sky130_fd_sc_hd__buf_2
X_78722_ _78722_/A _78722_/Y sky130_fd_sc_hd__inv_2
X_71057_ _71071_/A _71058_/A sky130_fd_sc_hd__buf_2
X_75934_ _81699_/D _75927_/B _75934_/Y sky130_fd_sc_hd__nor2_4
X_48882_ _48882_/A _48699_/B _48882_/Y sky130_fd_sc_hd__nand2_4
X_70008_ _83874_/Q _69988_/X _70007_/X _70008_/X sky130_fd_sc_hd__a21bo_4
X_47833_ _47832_/X _47841_/A sky130_fd_sc_hd__buf_2
X_59819_ _58094_/A _72381_/A sky130_fd_sc_hd__buf_2
X_78653_ _78654_/A _78654_/C _78652_/Y _78653_/X sky130_fd_sc_hd__a21o_4
X_75865_ _75865_/A _75865_/Y sky130_fd_sc_hd__inv_2
X_77604_ _77600_/Y _77603_/C _77603_/A _77604_/Y sky130_fd_sc_hd__o21ai_4
X_62830_ _57683_/X _62808_/X _62827_/X _62818_/X _62829_/X _62830_/Y
+ sky130_fd_sc_hd__a41oi_4
X_74816_ _59426_/X _46107_/A _74817_/A sky130_fd_sc_hd__nand2_4
X_47764_ _47799_/A _53232_/B _47764_/Y sky130_fd_sc_hd__nand2_4
X_78584_ _82805_/Q _78584_/Y sky130_fd_sc_hd__inv_2
X_44976_ _63049_/B _61375_/B sky130_fd_sc_hd__buf_2
X_75796_ _81099_/Q _75796_/B _75796_/Y sky130_fd_sc_hd__xnor2_4
X_49503_ _58896_/B _49496_/X _49502_/Y _49503_/Y sky130_fd_sc_hd__o21ai_4
X_46715_ _46715_/A _54325_/D sky130_fd_sc_hd__inv_2
X_77535_ _77538_/B _77535_/Y sky130_fd_sc_hd__inv_2
X_43927_ _43602_/X _43927_/X sky130_fd_sc_hd__buf_2
X_62761_ _57656_/X _62749_/X _62708_/X _62759_/X _62760_/X _62761_/Y
+ sky130_fd_sc_hd__a41oi_4
X_74747_ _70735_/X _74769_/D sky130_fd_sc_hd__buf_2
X_47695_ _54885_/B _53193_/B sky130_fd_sc_hd__buf_2
X_71959_ _71959_/A _71959_/X sky130_fd_sc_hd__buf_2
X_64500_ _84240_/Q _64429_/X _64499_/X _84240_/D sky130_fd_sc_hd__a21o_4
X_49434_ _49434_/A _49434_/X sky130_fd_sc_hd__buf_2
X_61712_ _61711_/X _61712_/X sky130_fd_sc_hd__buf_2
X_46646_ _54286_/D _51768_/D sky130_fd_sc_hd__buf_2
X_65480_ _65399_/X _65477_/Y _65479_/Y _65480_/Y sky130_fd_sc_hd__o21ai_4
X_77466_ _81938_/Q _82194_/D _81906_/D sky130_fd_sc_hd__xor2_4
X_43858_ _43858_/A _43858_/Y sky130_fd_sc_hd__inv_2
X_62692_ _60273_/A _62727_/B sky130_fd_sc_hd__buf_2
X_74678_ _74678_/A _74678_/Y sky130_fd_sc_hd__inv_2
X_79205_ _79195_/Y _79205_/B _79205_/C _79205_/Y sky130_fd_sc_hd__nand3_4
X_64431_ _58446_/A _64511_/B _64431_/Y sky130_fd_sc_hd__nor2_4
X_76417_ _76412_/X _76415_/Y _76417_/C _76417_/Y sky130_fd_sc_hd__nand3_4
X_42809_ _42808_/Y _87708_/D sky130_fd_sc_hd__inv_2
X_61643_ _61636_/Y _61638_/Y _61583_/Y _61640_/Y _61642_/Y _61643_/X
+ sky130_fd_sc_hd__a41o_4
X_49365_ _49363_/Y _49316_/X _49364_/X _49365_/Y sky130_fd_sc_hd__a21oi_4
X_73629_ _87344_/Q _73701_/B _73629_/Y sky130_fd_sc_hd__nor2_4
X_46577_ _46401_/A _57497_/A sky130_fd_sc_hd__buf_2
X_77397_ _77396_/Y _77397_/Y sky130_fd_sc_hd__inv_2
X_43789_ _41032_/X _43770_/X _69372_/B _43772_/X _43789_/X sky130_fd_sc_hd__a2bb2o_4
X_48316_ _86536_/Q _48263_/X _48315_/Y _48316_/Y sky130_fd_sc_hd__o21ai_4
X_67150_ _88379_/Q _67074_/X _67075_/X _67149_/X _67150_/X sky130_fd_sc_hd__a211o_4
X_79136_ _79136_/A _79136_/B _79136_/X sky130_fd_sc_hd__xor2_4
X_45528_ _45525_/X _45527_/Y _45348_/X _45528_/Y sky130_fd_sc_hd__a21oi_4
X_64362_ _64303_/A _64363_/B sky130_fd_sc_hd__buf_2
X_76348_ _76344_/Y _76348_/B _76348_/C _76348_/X sky130_fd_sc_hd__or3_4
X_49296_ _86415_/Q _49285_/X _49295_/Y _49296_/Y sky130_fd_sc_hd__o21ai_4
X_61574_ _61574_/A _61574_/Y sky130_fd_sc_hd__inv_2
X_66101_ _66226_/A _66101_/B _66101_/X sky130_fd_sc_hd__and2_4
X_63313_ _63289_/X _84886_/Q _63341_/C _63332_/D _63313_/X sky130_fd_sc_hd__and4_4
X_48247_ _48229_/A _53520_/B _48247_/Y sky130_fd_sc_hd__nand2_4
X_60525_ _60525_/A _60526_/B sky130_fd_sc_hd__buf_2
X_67081_ _66553_/X _67082_/A sky130_fd_sc_hd__buf_2
X_79067_ _79049_/A _79054_/A _79055_/A _79067_/Y sky130_fd_sc_hd__a21oi_4
X_45459_ _85021_/Q _55585_/B sky130_fd_sc_hd__inv_2
X_64293_ _64273_/A _64273_/B _84898_/Q _64304_/D _64293_/X sky130_fd_sc_hd__and4_4
X_76279_ _76260_/X _81642_/Q _76278_/Y _76281_/A sky130_fd_sc_hd__a21boi_4
X_66032_ _66020_/X _66030_/Y _66031_/Y _66032_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_541_0_CLK clkbuf_9_270_0_CLK/X _84105_/CLK sky130_fd_sc_hd__clkbuf_1
X_78018_ _78018_/A _78018_/B _78021_/A sky130_fd_sc_hd__or2_4
Xclkbuf_6_32_0_CLK clkbuf_6_33_0_CLK/A clkbuf_6_32_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_63244_ _63244_/A _63316_/B _63295_/C _63267_/D _63244_/X sky130_fd_sc_hd__or4_4
X_48178_ _47851_/B _48178_/X sky130_fd_sc_hd__buf_2
X_60456_ _79155_/A _60132_/X _60445_/Y _60455_/Y _60456_/X sky130_fd_sc_hd__a2bb2o_4
X_47129_ _46892_/A _47130_/A sky130_fd_sc_hd__buf_2
X_63175_ _60522_/A _63175_/X sky130_fd_sc_hd__buf_2
X_60387_ _60387_/A _60404_/C _60387_/C _60387_/X sky130_fd_sc_hd__and3_4
X_50140_ _65061_/B _50137_/X _50139_/Y _50140_/Y sky130_fd_sc_hd__o21ai_4
X_62126_ _61730_/X _62094_/B _59722_/X _62126_/D _62126_/X sky130_fd_sc_hd__and4_4
X_67983_ _68089_/A _67983_/X sky130_fd_sc_hd__buf_2
X_79969_ _79968_/Y _79977_/A sky130_fd_sc_hd__inv_2
Xclkbuf_10_556_0_CLK clkbuf_9_278_0_CLK/X _86941_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_47_0_CLK clkbuf_6_47_0_CLK/A clkbuf_7_95_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_69722_ _69766_/A _69722_/B _69722_/Y sky130_fd_sc_hd__nor2_4
X_50071_ _50084_/A _48912_/B _50071_/Y sky130_fd_sc_hd__nand2_4
X_66934_ _66931_/X _66933_/X _66934_/Y sky130_fd_sc_hd__nand2_4
X_62057_ _59761_/A _62094_/B _59722_/X _62057_/D _62057_/X sky130_fd_sc_hd__and4_4
X_82980_ _82980_/CLK _82980_/D _45847_/A sky130_fd_sc_hd__dfxtp_4
X_61008_ _61008_/A _61008_/Y sky130_fd_sc_hd__inv_2
X_81931_ _82234_/CLK _77818_/Y _81931_/Q sky130_fd_sc_hd__dfxtp_4
X_69653_ _44531_/A _69485_/X _69611_/X _69652_/X _69653_/X sky130_fd_sc_hd__a211o_4
X_66865_ _87367_/Q _66797_/X _66863_/X _66864_/X _66865_/X sky130_fd_sc_hd__a211o_4
X_68604_ _68604_/A _68604_/B _68604_/X sky130_fd_sc_hd__and2_4
X_53830_ _48979_/A _53806_/B _53806_/C _53830_/X sky130_fd_sc_hd__and3_4
X_65816_ _65929_/A _65916_/B sky130_fd_sc_hd__buf_2
X_84650_ _84652_/CLK _84650_/D _60152_/A sky130_fd_sc_hd__dfxtp_4
X_81862_ _81859_/CLK _78053_/X _81862_/Q sky130_fd_sc_hd__dfxtp_4
X_69584_ _88082_/Q _69582_/X _69567_/X _69583_/Y _69584_/X sky130_fd_sc_hd__a211o_4
X_66796_ _87882_/Q _66697_/X _66794_/X _66795_/X _66796_/X sky130_fd_sc_hd__a211o_4
X_83601_ _86145_/CLK _71120_/Y _83601_/Q sky130_fd_sc_hd__dfxtp_4
X_80813_ _80813_/CLK _83957_/Q _75817_/B sky130_fd_sc_hd__dfxtp_4
X_68535_ _68560_/A _88269_/Q _68535_/X sky130_fd_sc_hd__and2_4
X_53761_ _53766_/A _48672_/A _53761_/Y sky130_fd_sc_hd__nand2_4
X_65747_ _65162_/X _65653_/B _65165_/X _65747_/Y sky130_fd_sc_hd__nand3_4
X_84581_ _84562_/CLK _84581_/D _60717_/C sky130_fd_sc_hd__dfxtp_4
X_50973_ _50973_/A _50973_/X sky130_fd_sc_hd__buf_2
X_62959_ _62967_/A _63316_/A _62939_/X _62967_/D _62959_/X sky130_fd_sc_hd__and4_4
X_81793_ _82369_/CLK _75966_/X _81793_/Q sky130_fd_sc_hd__dfxtp_4
X_55500_ _82997_/Q _55498_/X _44096_/X _55499_/X _55500_/X sky130_fd_sc_hd__a211o_4
X_86320_ _86640_/CLK _49808_/Y _57958_/B sky130_fd_sc_hd__dfxtp_4
X_52712_ _52657_/A _52718_/A sky130_fd_sc_hd__buf_2
X_83532_ _86490_/CLK _71334_/Y _48130_/A sky130_fd_sc_hd__dfxtp_4
X_56480_ _56031_/X _56468_/X _56479_/Y _85180_/D sky130_fd_sc_hd__o21ai_4
X_80744_ _81994_/CLK _75168_/X _80744_/Q sky130_fd_sc_hd__dfxtp_4
X_68466_ _73650_/A _68463_/X _68439_/X _68465_/Y _68466_/X sky130_fd_sc_hd__a211o_4
X_53692_ _50469_/A _53720_/B _53692_/C _53692_/X sky130_fd_sc_hd__and3_4
X_65678_ _65039_/X _65828_/B _65041_/X _65678_/Y sky130_fd_sc_hd__nand3_4
X_55431_ _55415_/B _55431_/Y sky130_fd_sc_hd__inv_2
X_67417_ _67320_/A _67417_/B _67417_/X sky130_fd_sc_hd__and2_4
X_86251_ _86154_/CLK _86251_/D _86251_/Q sky130_fd_sc_hd__dfxtp_4
X_52643_ _52643_/A _52654_/B _52643_/C _46736_/X _52643_/X sky130_fd_sc_hd__and4_4
X_64629_ _64629_/A _64629_/X sky130_fd_sc_hd__buf_2
X_83463_ _83495_/CLK _83463_/D _59457_/B sky130_fd_sc_hd__dfxtp_4
X_80675_ _80679_/CLK _80675_/D _80675_/Q sky130_fd_sc_hd__dfxtp_4
X_68397_ _69877_/A _88370_/Q _68397_/X sky130_fd_sc_hd__and2_4
X_85202_ _85297_/CLK _56417_/Y _85202_/Q sky130_fd_sc_hd__dfxtp_4
X_58150_ _63022_/A _63380_/A sky130_fd_sc_hd__buf_2
XPHY_505 sky130_fd_sc_hd__decap_3
X_82414_ _82248_/CLK _82446_/Q _78472_/A sky130_fd_sc_hd__dfxtp_4
X_55362_ _55362_/A _55363_/B sky130_fd_sc_hd__inv_2
X_67348_ _66868_/A _67348_/X sky130_fd_sc_hd__buf_2
X_86182_ _85859_/CLK _86182_/D _86182_/Q sky130_fd_sc_hd__dfxtp_4
X_52574_ _52572_/Y _52532_/X _52573_/X _85794_/D sky130_fd_sc_hd__a21oi_4
XPHY_516 sky130_fd_sc_hd__decap_3
X_83394_ _83756_/CLK _71734_/Y _58246_/A sky130_fd_sc_hd__dfxtp_4
XPHY_527 sky130_fd_sc_hd__decap_3
XPHY_538 sky130_fd_sc_hd__decap_3
X_57101_ _57097_/X _56575_/X _45422_/A _57099_/X _57101_/X sky130_fd_sc_hd__a2bb2o_4
X_54313_ _54310_/Y _54311_/X _54312_/X _85465_/D sky130_fd_sc_hd__a21oi_4
XPHY_549 sky130_fd_sc_hd__decap_3
X_85133_ _85071_/CLK _85133_/D _85133_/Q sky130_fd_sc_hd__dfxtp_4
X_51525_ _85994_/Q _51511_/X _51524_/Y _51525_/Y sky130_fd_sc_hd__o21ai_4
X_58081_ _58576_/A _58081_/B _58081_/Y sky130_fd_sc_hd__nor2_4
X_82345_ _82369_/CLK _77103_/X _48086_/A sky130_fd_sc_hd__dfxtp_4
X_67279_ _67183_/A _67279_/B _67279_/X sky130_fd_sc_hd__and2_4
X_55293_ _55139_/X _55146_/X _83747_/Q _55293_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_10_509_0_CLK clkbuf_9_254_0_CLK/X _82956_/CLK sky130_fd_sc_hd__clkbuf_1
X_57032_ _56820_/A _57043_/B _57032_/Y sky130_fd_sc_hd__nand2_4
X_69018_ _69013_/X _69016_/X _69017_/X _69018_/Y sky130_fd_sc_hd__a21oi_4
X_54244_ _85477_/Q _54220_/X _54243_/Y _54244_/Y sky130_fd_sc_hd__o21ai_4
X_85064_ _84998_/CLK _85064_/D _57199_/A sky130_fd_sc_hd__dfxtp_4
X_51456_ _51456_/A _51473_/B _51467_/C _52982_/D _51456_/X sky130_fd_sc_hd__and4_4
X_70290_ _70292_/A _70292_/B _83105_/Q _70292_/D _70290_/X sky130_fd_sc_hd__and4_4
X_82276_ _82103_/CLK _82276_/D _40919_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_0_0_CLK clkbuf_8_1_0_CLK/A clkbuf_8_0_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_84015_ _84074_/CLK _68195_/X _82055_/D sky130_fd_sc_hd__dfxtp_4
X_50407_ _50510_/A _50435_/C sky130_fd_sc_hd__buf_2
X_81227_ _81227_/CLK _81035_/Q _81227_/Q sky130_fd_sc_hd__dfxtp_4
X_54175_ _54184_/A _47360_/A _54175_/Y sky130_fd_sc_hd__nand2_4
X_51387_ _51789_/A _51387_/X sky130_fd_sc_hd__buf_2
X_53126_ _53123_/Y _53111_/X _53125_/X _53126_/Y sky130_fd_sc_hd__a21oi_4
X_41140_ _41112_/X _41113_/X _41139_/X _88270_/Q _41088_/X _41141_/A
+ sky130_fd_sc_hd__o32ai_4
X_50338_ _50510_/A _50338_/X sky130_fd_sc_hd__buf_2
X_81158_ _81160_/CLK _74874_/B _81158_/Q sky130_fd_sc_hd__dfxtp_4
X_58983_ _58983_/A _58985_/A sky130_fd_sc_hd__inv_2
X_80109_ _57922_/Y _65651_/C _80108_/Y _80109_/X sky130_fd_sc_hd__o21a_4
X_41071_ _41070_/X _41065_/X _69472_/B _41066_/X _41071_/X sky130_fd_sc_hd__a2bb2o_4
X_53057_ _53112_/A _53074_/A sky130_fd_sc_hd__buf_2
X_57934_ _57971_/A _57934_/B _57934_/Y sky130_fd_sc_hd__nor2_4
X_50269_ _86234_/Q _50238_/X _50268_/Y _50269_/Y sky130_fd_sc_hd__o21ai_4
X_73980_ _73967_/X _73981_/C _73979_/X _73980_/X sky130_fd_sc_hd__a21o_4
X_85966_ _85679_/CLK _85966_/D _85966_/Q sky130_fd_sc_hd__dfxtp_4
X_81089_ _81121_/CLK _81121_/Q _81089_/Q sky130_fd_sc_hd__dfxtp_4
X_52008_ _52006_/Y _51981_/X _52007_/Y _85907_/D sky130_fd_sc_hd__a21boi_4
X_87705_ _87446_/CLK _87705_/D _87705_/Q sky130_fd_sc_hd__dfxtp_4
X_72931_ _73306_/A _73093_/A sky130_fd_sc_hd__buf_2
X_84917_ _84906_/CLK _58165_/X _58162_/A sky130_fd_sc_hd__dfxtp_4
X_57865_ _84944_/Q _57819_/X _57859_/X _57864_/X _57865_/Y sky130_fd_sc_hd__a2bb2oi_4
X_85897_ _86218_/CLK _52059_/Y _74127_/B sky130_fd_sc_hd__dfxtp_4
X_59604_ _59600_/X _72569_/C _59604_/X sky130_fd_sc_hd__and2_4
X_44830_ _41697_/A _44817_/X _67629_/B _44818_/X _86931_/D sky130_fd_sc_hd__a2bb2o_4
X_56816_ _56816_/A _56816_/Y sky130_fd_sc_hd__inv_2
X_75650_ _75650_/A _75650_/B _75650_/Y sky130_fd_sc_hd__xnor2_4
X_87636_ _87636_/CLK _42949_/Y _68078_/B sky130_fd_sc_hd__dfxtp_4
X_84848_ _83457_/CLK _58439_/X _84848_/Q sky130_fd_sc_hd__dfxtp_4
X_72862_ _72861_/X _72862_/X sky130_fd_sc_hd__buf_2
X_57796_ _57781_/X _57786_/Y _57792_/Y _57793_/X _57795_/X _57796_/X
+ sky130_fd_sc_hd__o32a_4
X_74601_ _74591_/X _74599_/X _56121_/A _74600_/X _74601_/X sky130_fd_sc_hd__a211o_4
X_71813_ _71813_/A _70476_/X _70852_/C _71813_/X sky130_fd_sc_hd__and3_4
X_59535_ _59535_/A _61285_/C sky130_fd_sc_hd__buf_2
X_44761_ _44740_/X _44741_/X _41320_/X _86968_/Q _44742_/X _44762_/A
+ sky130_fd_sc_hd__o32ai_4
X_56747_ _55383_/A _56707_/X _55377_/Y _57427_/A sky130_fd_sc_hd__nand3_4
X_75581_ _80899_/Q _75584_/C sky130_fd_sc_hd__inv_2
X_87567_ _87288_/CLK _43123_/Y _72859_/A sky130_fd_sc_hd__dfxtp_4
X_41973_ _41973_/A _41973_/Y sky130_fd_sc_hd__inv_2
X_53959_ _53949_/A _53959_/B _53959_/Y sky130_fd_sc_hd__nand2_4
X_72793_ _83176_/Q _72709_/X _72792_/Y _72793_/X sky130_fd_sc_hd__a21o_4
X_84779_ _83464_/CLK _58992_/X _58990_/A sky130_fd_sc_hd__dfxtp_4
X_46500_ _83635_/Q _46500_/Y sky130_fd_sc_hd__inv_2
X_77320_ _77318_/Y _77290_/B _77319_/X _77320_/Y sky130_fd_sc_hd__o21ai_4
X_43712_ _43712_/A _43712_/Y sky130_fd_sc_hd__inv_2
X_74532_ _52829_/B _74516_/X _74531_/Y _74532_/Y sky130_fd_sc_hd__o21ai_4
X_86518_ _86516_/CLK _86518_/D _73070_/B sky130_fd_sc_hd__dfxtp_4
X_40924_ _40817_/X _82275_/Q _40923_/X _40924_/Y sky130_fd_sc_hd__o21ai_4
X_71744_ _71171_/A _70656_/B _71744_/C _71744_/D _71744_/Y sky130_fd_sc_hd__nand4_4
X_47480_ _47480_/A _47481_/A sky130_fd_sc_hd__inv_2
X_59466_ _59462_/X _83461_/Q _59465_/Y _84725_/D sky130_fd_sc_hd__o21a_4
X_44692_ _44686_/X _44687_/X _40633_/X _44691_/Y _44689_/X _44692_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56678_ _83337_/Q _57140_/B sky130_fd_sc_hd__buf_2
X_87498_ _88012_/CLK _43285_/X _87498_/Q sky130_fd_sc_hd__dfxtp_4
X_46431_ _46366_/A _46434_/A sky130_fd_sc_hd__buf_2
X_58417_ _84853_/Q _58418_/A sky130_fd_sc_hd__inv_2
X_77251_ _77249_/A _82084_/D _77253_/A sky130_fd_sc_hd__nand2_4
X_43643_ _43642_/X _87330_/D sky130_fd_sc_hd__inv_2
X_55629_ _45413_/A _44116_/B _55627_/X _55628_/Y _55629_/X sky130_fd_sc_hd__a211o_4
X_86449_ _85557_/CLK _49051_/Y _86449_/Q sky130_fd_sc_hd__dfxtp_4
X_74463_ _74492_/A _74463_/X sky130_fd_sc_hd__buf_2
X_40855_ _40835_/X _40836_/X _40854_/X _88322_/Q _40832_/X _40855_/Y
+ sky130_fd_sc_hd__o32ai_4
X_71675_ _58472_/Y _71669_/X _71674_/Y _83416_/D sky130_fd_sc_hd__o21ai_4
X_59397_ _58425_/A _59398_/A sky130_fd_sc_hd__buf_2
X_76202_ _76200_/X _76201_/Y _81638_/Q _76202_/X sky130_fd_sc_hd__a21o_4
X_49150_ _52395_/B _50183_/B sky130_fd_sc_hd__buf_2
X_73414_ _83152_/Q _73318_/X _73413_/Y _73414_/X sky130_fd_sc_hd__a21o_4
X_46362_ _46362_/A _52468_/B _46362_/Y sky130_fd_sc_hd__nand2_4
X_70626_ _70625_/Y _70630_/B sky130_fd_sc_hd__buf_2
X_58348_ _58348_/A _58364_/B _58348_/Y sky130_fd_sc_hd__nand2_4
X_77182_ _82107_/Q _77182_/B _77182_/X sky130_fd_sc_hd__xor2_4
X_43574_ _53443_/A _53455_/A sky130_fd_sc_hd__buf_2
X_74394_ _83075_/Q _74377_/X _74393_/Y _74394_/Y sky130_fd_sc_hd__o21ai_4
X_40786_ _40783_/X _82301_/Q _40785_/X _40787_/A sky130_fd_sc_hd__o21a_4
X_48101_ _48093_/Y _48055_/X _48100_/X _48101_/Y sky130_fd_sc_hd__a21oi_4
X_45313_ _85254_/Q _45297_/X _45312_/X _45313_/Y sky130_fd_sc_hd__o21ai_4
X_76133_ _81726_/D _76133_/B _76133_/Y sky130_fd_sc_hd__nand2_4
X_88119_ _87417_/CLK _88119_/D _67245_/B sky130_fd_sc_hd__dfxtp_4
X_42525_ _74143_/A _42525_/Y sky130_fd_sc_hd__inv_2
X_49081_ _49075_/Y _49038_/X _49080_/X _86446_/D sky130_fd_sc_hd__a21oi_4
X_73345_ _73345_/A _73003_/B _73345_/Y sky130_fd_sc_hd__nor2_4
X_46293_ _46623_/A _46421_/A sky130_fd_sc_hd__buf_2
X_70557_ DATA_TO_HASH[3] _71883_/A sky130_fd_sc_hd__inv_2
X_58279_ _58279_/A _58279_/Y sky130_fd_sc_hd__inv_2
X_48032_ _48004_/A _50328_/B _48032_/Y sky130_fd_sc_hd__nand2_4
X_60310_ _60275_/X _60344_/B _59789_/A _60259_/A _60309_/X _60310_/X
+ sky130_fd_sc_hd__a2111o_4
X_45244_ _45244_/A _45244_/Y sky130_fd_sc_hd__inv_2
X_76064_ _76052_/Y _76064_/B _76064_/Y sky130_fd_sc_hd__nand2_4
X_42456_ _51238_/B _42430_/X _40573_/X _68380_/A _42453_/X _42456_/Y
+ sky130_fd_sc_hd__o32ai_4
X_61290_ _61290_/A _61290_/X sky130_fd_sc_hd__buf_2
X_73276_ _69838_/B _73250_/X _73251_/X _73275_/Y _73276_/X sky130_fd_sc_hd__a211o_4
X_70488_ _71090_/A _71779_/B sky130_fd_sc_hd__buf_2
X_75015_ _81146_/D _75016_/B _75018_/A sky130_fd_sc_hd__nor2_4
X_41407_ _41373_/X _41747_/A _41406_/X _41407_/X sky130_fd_sc_hd__o21a_4
X_60241_ _60241_/A _60367_/B sky130_fd_sc_hd__buf_2
X_72227_ _72166_/X _85368_/Q _72226_/X _72227_/Y sky130_fd_sc_hd__o21ai_4
X_45175_ _85263_/Q _45147_/X _45174_/X _45175_/Y sky130_fd_sc_hd__o21ai_4
X_42387_ _40387_/X _42374_/X _87888_/Q _42375_/X _42387_/X sky130_fd_sc_hd__a2bb2o_4
X_44126_ _73352_/A _44126_/X sky130_fd_sc_hd__buf_2
X_79823_ _84227_/Q _83275_/Q _79823_/Y sky130_fd_sc_hd__nand2_4
X_41338_ _41490_/A _41338_/X sky130_fd_sc_hd__buf_2
X_60172_ _60172_/A _60406_/B sky130_fd_sc_hd__buf_2
X_72158_ _59368_/X _85982_/Q _72157_/X _72158_/Y sky130_fd_sc_hd__o21ai_4
X_49983_ _49930_/X _50005_/C sky130_fd_sc_hd__buf_2
X_71109_ _52367_/B _71095_/A _71108_/Y _83604_/D sky130_fd_sc_hd__o21ai_4
X_48934_ _48934_/A _48985_/A sky130_fd_sc_hd__buf_2
X_44057_ _55152_/A _44058_/A sky130_fd_sc_hd__buf_2
X_79754_ _84221_/Q _83269_/Q _79761_/A sky130_fd_sc_hd__xor2_4
X_41269_ _41268_/X _41251_/X _69048_/B _41253_/X _41269_/X sky130_fd_sc_hd__a2bb2o_4
X_64980_ _64980_/A _64980_/X sky130_fd_sc_hd__buf_2
X_72089_ _72087_/Y _72083_/X _72088_/Y _83287_/D sky130_fd_sc_hd__a21boi_4
X_76966_ _76662_/A _76658_/Y _76966_/Y sky130_fd_sc_hd__nand2_4
X_43008_ _52021_/A _51934_/A sky130_fd_sc_hd__buf_2
X_78705_ _78675_/B _78701_/X _78742_/B _78706_/B sky130_fd_sc_hd__a21boi_4
X_63931_ _63927_/X _63913_/X _63930_/Y _84286_/D sky130_fd_sc_hd__a21oi_4
X_75917_ _84515_/Q _84387_/Q _75917_/X sky130_fd_sc_hd__xor2_4
X_48865_ _48840_/A _48865_/X sky130_fd_sc_hd__buf_2
X_79685_ _79669_/X _79672_/Y _79684_/X _79685_/X sky130_fd_sc_hd__a21o_4
X_76897_ _76895_/Y _76894_/Y _76897_/Y sky130_fd_sc_hd__nand2_4
X_47816_ _47811_/Y _47791_/X _47815_/X _86595_/D sky130_fd_sc_hd__a21oi_4
X_66650_ _66646_/X _66649_/X _66650_/Y sky130_fd_sc_hd__nand2_4
X_78636_ _78632_/X _78637_/C _78637_/B _78638_/A sky130_fd_sc_hd__a21o_4
X_63862_ _63831_/A _64292_/A _63862_/C _63862_/X sky130_fd_sc_hd__and3_4
X_75848_ _80895_/D _75848_/B _75850_/A sky130_fd_sc_hd__nand2_4
X_48796_ _48833_/A _48829_/B sky130_fd_sc_hd__buf_2
X_65601_ _65533_/X _65599_/Y _65600_/Y _65601_/Y sky130_fd_sc_hd__o21ai_4
X_62813_ _61490_/X _62834_/B _62801_/X _62834_/D _62813_/Y sky130_fd_sc_hd__nand4_4
X_47747_ _47747_/A _55083_/D sky130_fd_sc_hd__inv_2
X_66581_ _45915_/X _68474_/A sky130_fd_sc_hd__buf_2
X_78567_ _78566_/A _82720_/Q _78568_/A sky130_fd_sc_hd__nand2_4
X_44959_ _45720_/A _44959_/X sky130_fd_sc_hd__buf_2
X_63793_ _58228_/X _64189_/C _60908_/A _63793_/D _63794_/D sky130_fd_sc_hd__nand4_4
X_75779_ _81097_/Q _80809_/Q _75779_/Y sky130_fd_sc_hd__xnor2_4
X_68320_ _67966_/X _67968_/X _68295_/X _68320_/Y sky130_fd_sc_hd__a21oi_4
X_65532_ _65528_/Y _65529_/X _65531_/X _84195_/D sky130_fd_sc_hd__a21o_4
X_77518_ _77518_/A _82114_/Q _77518_/X sky130_fd_sc_hd__xor2_4
X_62744_ _62667_/X _62744_/X sky130_fd_sc_hd__buf_2
X_47678_ _83553_/Q _47679_/A sky130_fd_sc_hd__inv_2
X_78498_ _78482_/B _78496_/X _78497_/X _78498_/Y sky130_fd_sc_hd__a21boi_4
X_49417_ _49444_/A _49418_/A sky130_fd_sc_hd__buf_2
X_68251_ _67562_/X _67564_/X _68216_/X _68251_/Y sky130_fd_sc_hd__a21oi_4
X_46629_ _46629_/A _54275_/D sky130_fd_sc_hd__inv_2
X_65463_ _65399_/X _65461_/Y _65462_/Y _65463_/Y sky130_fd_sc_hd__o21ai_4
X_77449_ _77447_/X _77448_/Y _77449_/X sky130_fd_sc_hd__and2_4
X_62675_ _62737_/A _62676_/C sky130_fd_sc_hd__buf_2
X_67202_ _87353_/Q _67156_/X _67106_/X _67201_/X _67202_/X sky130_fd_sc_hd__a211o_4
X_64414_ _58254_/Y _64367_/X _64413_/Y _64414_/Y sky130_fd_sc_hd__o21ai_4
X_49348_ _49352_/A _50870_/B _49348_/Y sky130_fd_sc_hd__nand2_4
X_61626_ _61374_/A _61636_/A sky130_fd_sc_hd__buf_2
X_80460_ _80457_/X _80460_/B _82257_/D sky130_fd_sc_hd__xor2_4
X_68182_ _68144_/X _67130_/Y _68168_/X _68181_/Y _68182_/X sky130_fd_sc_hd__a211o_4
X_65394_ _65390_/X _65192_/B _65393_/X _65394_/Y sky130_fd_sc_hd__nand3_4
X_67133_ _67133_/A _67133_/B _67133_/X sky130_fd_sc_hd__and2_4
X_79119_ _79031_/B _79119_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_480_0_CLK clkbuf_9_240_0_CLK/X _86289_/CLK sky130_fd_sc_hd__clkbuf_1
X_64345_ _64344_/X _64307_/B _84830_/Q _64345_/X sky130_fd_sc_hd__and3_4
X_49279_ _49232_/A _50799_/B _49279_/Y sky130_fd_sc_hd__nand2_4
X_61557_ _61374_/A _61558_/A sky130_fd_sc_hd__buf_2
X_80391_ _80391_/A _63636_/C _80391_/X sky130_fd_sc_hd__xor2_4
X_51310_ _51286_/A _51310_/X sky130_fd_sc_hd__buf_2
X_82130_ _81970_/CLK _82130_/D _82086_/D sky130_fd_sc_hd__dfxtp_4
X_60508_ _60508_/A _63252_/B sky130_fd_sc_hd__buf_2
X_67064_ _67087_/A _88127_/Q _67064_/X sky130_fd_sc_hd__and2_4
X_52290_ _52247_/A _52291_/C sky130_fd_sc_hd__buf_2
X_64276_ _64248_/A _64248_/B _64276_/C _64276_/X sky130_fd_sc_hd__and3_4
X_61488_ _61486_/X _61455_/X _61487_/Y _84477_/D sky130_fd_sc_hd__a21oi_4
X_66015_ _65903_/X _65543_/Y _66014_/Y _66015_/Y sky130_fd_sc_hd__o21ai_4
X_51241_ _64617_/B _51233_/X _51240_/Y _51241_/Y sky130_fd_sc_hd__o21ai_4
X_63227_ _63216_/X _63227_/B _63241_/C _63181_/X _63227_/X sky130_fd_sc_hd__and4_4
X_82061_ _84105_/CLK _82061_/D _77825_/A sky130_fd_sc_hd__dfxtp_4
X_60439_ _60501_/A _60439_/X sky130_fd_sc_hd__buf_2
X_81012_ _85315_/CLK _84220_/Q _81012_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_495_0_CLK clkbuf_9_247_0_CLK/X _83685_/CLK sky130_fd_sc_hd__clkbuf_1
X_51172_ _51168_/Y _51147_/X _51171_/X _51172_/Y sky130_fd_sc_hd__a21oi_4
X_63158_ _63157_/X _63158_/B _63147_/C _63124_/D _63158_/X sky130_fd_sc_hd__and4_4
X_50123_ _50121_/Y _50117_/X _50122_/X _86260_/D sky130_fd_sc_hd__a21oi_4
X_62109_ _58187_/X _62105_/X _61916_/X _61948_/X _62108_/X _62109_/X
+ sky130_fd_sc_hd__a41o_4
X_85820_ _86045_/CLK _52451_/Y _64743_/B sky130_fd_sc_hd__dfxtp_4
X_55980_ _55977_/X _55979_/X _55615_/X _55983_/A sky130_fd_sc_hd__a21o_4
X_67966_ _67963_/X _67965_/X _67917_/X _67966_/X sky130_fd_sc_hd__a21o_4
X_63089_ _63041_/A _63089_/B _63079_/C _63066_/D _63089_/X sky130_fd_sc_hd__and4_4
X_69705_ _69702_/X _69704_/X _69655_/X _69705_/Y sky130_fd_sc_hd__a21oi_4
X_50054_ _48885_/A _48859_/B _48854_/C _50054_/X sky130_fd_sc_hd__and3_4
X_54931_ _85351_/Q _54918_/X _54930_/Y _54931_/Y sky130_fd_sc_hd__o21ai_4
X_66917_ _87365_/Q _66915_/X _66863_/X _66916_/X _66917_/X sky130_fd_sc_hd__a211o_4
X_85751_ _85751_/CLK _52806_/Y _85751_/Q sky130_fd_sc_hd__dfxtp_4
X_82963_ _82965_/CLK _82771_/Q _82963_/Q sky130_fd_sc_hd__dfxtp_4
X_67897_ _67014_/X _67897_/X sky130_fd_sc_hd__buf_2
X_84702_ _84713_/CLK _59780_/Y _80506_/A sky130_fd_sc_hd__dfxtp_4
X_57650_ _57650_/A _57650_/X sky130_fd_sc_hd__buf_2
Xclkbuf_4_10_1_CLK clkbuf_4_10_1_CLK/A clkbuf_4_10_1_CLK/X sky130_fd_sc_hd__clkbuf_1
X_81914_ _82008_/CLK _81914_/D _82290_/D sky130_fd_sc_hd__dfxtp_4
X_69636_ _88078_/Q _69582_/X _69567_/X _69635_/Y _69636_/X sky130_fd_sc_hd__a211o_4
X_54862_ _54889_/A _54883_/C sky130_fd_sc_hd__buf_2
X_66848_ _66757_/X _66837_/Y _66793_/X _66847_/Y _66848_/X sky130_fd_sc_hd__a211o_4
X_85682_ _84797_/CLK _85682_/D _85682_/Q sky130_fd_sc_hd__dfxtp_4
X_82894_ _87473_/CLK _78168_/B _41729_/A sky130_fd_sc_hd__dfxtp_4
X_56601_ _56551_/X _56774_/A sky130_fd_sc_hd__buf_2
X_87421_ _87421_/CLK _43439_/Y _87421_/Q sky130_fd_sc_hd__dfxtp_4
X_53813_ _85563_/Q _53722_/X _53812_/Y _53813_/Y sky130_fd_sc_hd__o21ai_4
X_84633_ _84487_/CLK _60322_/X _79713_/A sky130_fd_sc_hd__dfxtp_4
X_57581_ _72009_/A _57581_/X sky130_fd_sc_hd__buf_2
X_81845_ _81839_/CLK _81877_/Q _77507_/A sky130_fd_sc_hd__dfxtp_4
X_69567_ _69567_/A _69567_/X sky130_fd_sc_hd__buf_2
X_54793_ _54900_/A _54816_/B sky130_fd_sc_hd__buf_2
X_66779_ _66776_/X _66778_/X _66706_/X _66779_/Y sky130_fd_sc_hd__a21oi_4
X_59320_ _59260_/X _85415_/Q _59319_/X _59320_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_433_0_CLK clkbuf_9_216_0_CLK/X _83498_/CLK sky130_fd_sc_hd__clkbuf_1
X_56532_ _56144_/X _56528_/X _56531_/Y _56532_/Y sky130_fd_sc_hd__o21ai_4
X_68518_ _68437_/A _87341_/Q _68518_/X sky130_fd_sc_hd__and2_4
X_87352_ _81154_/CLK _87352_/D _87352_/Q sky130_fd_sc_hd__dfxtp_4
X_53744_ _53742_/Y _53715_/X _53743_/X _53744_/Y sky130_fd_sc_hd__a21oi_4
X_84564_ _84564_/CLK _84564_/D _78059_/A sky130_fd_sc_hd__dfxtp_4
X_50956_ _86100_/Q _50936_/X _50955_/Y _50956_/Y sky130_fd_sc_hd__o21ai_4
X_69498_ _87013_/Q _69457_/X _69458_/X _69497_/X _69498_/X sky130_fd_sc_hd__a211o_4
X_81776_ _86753_/CLK _76074_/X _81776_/Q sky130_fd_sc_hd__dfxtp_4
X_86303_ _86303_/CLK _49900_/Y _72139_/B sky130_fd_sc_hd__dfxtp_4
X_59251_ _59248_/Y _59250_/Y _59140_/X _59251_/X sky130_fd_sc_hd__a21o_4
X_83515_ _83515_/CLK _71392_/X _83515_/Q sky130_fd_sc_hd__dfxtp_4
X_56463_ _56463_/A _56525_/A sky130_fd_sc_hd__buf_2
X_68449_ _88016_/Q _68402_/X _68359_/X _68448_/X _68449_/X sky130_fd_sc_hd__a211o_4
X_80727_ _80708_/CLK _75913_/X _80695_/D sky130_fd_sc_hd__dfxtp_4
X_87283_ _87285_/CLK _87283_/D _87283_/Q sky130_fd_sc_hd__dfxtp_4
X_53675_ _85590_/Q _53660_/X _53674_/Y _53675_/Y sky130_fd_sc_hd__o21ai_4
X_84495_ _84649_/CLK _84495_/D _61262_/C sky130_fd_sc_hd__dfxtp_4
X_50887_ _50885_/Y _50839_/X _50886_/X _86113_/D sky130_fd_sc_hd__a21oi_4
X_58202_ _58201_/X _58184_/B _58202_/Y sky130_fd_sc_hd__nor2_4
X_55414_ _55411_/Y _55414_/B _55415_/C sky130_fd_sc_hd__and2_4
X_86234_ _86238_/CLK _50271_/Y _86234_/Q sky130_fd_sc_hd__dfxtp_4
X_52626_ _52626_/A _52643_/C sky130_fd_sc_hd__buf_2
X_40640_ _40577_/X _82872_/Q _40639_/X _40640_/X sky130_fd_sc_hd__o21a_4
X_71460_ _70692_/A _71446_/X _71458_/C _71460_/Y sky130_fd_sc_hd__nor3_4
X_59182_ _84762_/Q _59182_/Y sky130_fd_sc_hd__inv_2
X_83446_ _83480_/CLK _83446_/D _83446_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_302 sky130_fd_sc_hd__decap_3
X_56394_ _56377_/X _56394_/X sky130_fd_sc_hd__buf_2
X_80658_ _80657_/CLK _80658_/D _46115_/A sky130_fd_sc_hd__dfxtp_4
XPHY_313 sky130_fd_sc_hd__decap_3
Xclkbuf_10_448_0_CLK clkbuf_9_224_0_CLK/X _83711_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_324 sky130_fd_sc_hd__decap_3
X_70411_ _70410_/Y _71012_/A sky130_fd_sc_hd__buf_2
X_58133_ _57989_/X _58130_/Y _58132_/Y _58007_/X _57993_/X _58133_/X
+ sky130_fd_sc_hd__o32a_4
XPHY_335 sky130_fd_sc_hd__decap_3
X_55345_ _57409_/A _55346_/B sky130_fd_sc_hd__inv_2
X_86165_ _85557_/CLK _86165_/D _86165_/Q sky130_fd_sc_hd__dfxtp_4
X_40571_ _40571_/A _48606_/A _40571_/X sky130_fd_sc_hd__or2_4
X_52557_ _52542_/X _54075_/B _52557_/Y sky130_fd_sc_hd__nand2_4
XPHY_346 sky130_fd_sc_hd__decap_3
X_71391_ _70689_/A _71386_/B _71399_/C _71391_/Y sky130_fd_sc_hd__nor3_4
X_83377_ _83372_/CLK _83377_/D _83377_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_357 sky130_fd_sc_hd__decap_3
X_80589_ _80587_/X _80589_/B _80608_/B sky130_fd_sc_hd__xnor2_4
XPHY_368 sky130_fd_sc_hd__decap_3
X_42310_ _41601_/X _42303_/X _87928_/Q _42305_/X _87928_/D sky130_fd_sc_hd__a2bb2o_4
X_73130_ _69756_/B _73086_/X _73087_/X _73130_/X sky130_fd_sc_hd__o21a_4
XPHY_379 sky130_fd_sc_hd__decap_3
X_85116_ _85114_/CLK _85116_/D _85116_/Q sky130_fd_sc_hd__dfxtp_4
X_51508_ _85997_/Q _51485_/X _51507_/Y _51508_/Y sky130_fd_sc_hd__o21ai_4
X_58064_ _58017_/X _85384_/Q _58063_/X _58064_/Y sky130_fd_sc_hd__o21ai_4
X_70342_ _70338_/A _70333_/B _83086_/Q _70332_/X _70342_/X sky130_fd_sc_hd__and4_4
X_82328_ _82327_/CLK _77161_/B _82328_/Q sky130_fd_sc_hd__dfxtp_4
X_55276_ _55276_/A _84999_/Q _55276_/X sky130_fd_sc_hd__and2_4
X_43290_ _41169_/X _43287_/X _87496_/Q _43288_/X _87496_/D sky130_fd_sc_hd__a2bb2o_4
X_86096_ _86096_/CLK _86096_/D _86096_/Q sky130_fd_sc_hd__dfxtp_4
X_52488_ _52487_/X _46407_/X _52488_/Y sky130_fd_sc_hd__nand2_4
X_57015_ _57013_/X _57014_/Y _44213_/X _57015_/Y sky130_fd_sc_hd__o21ai_4
X_54227_ _54254_/A _54237_/C sky130_fd_sc_hd__buf_2
X_42241_ _42241_/A _42241_/Y sky130_fd_sc_hd__inv_2
X_73061_ _44543_/Y _73006_/X _73060_/Y _73075_/C sky130_fd_sc_hd__a21o_4
X_85047_ _85013_/CLK _57258_/Y _45553_/A sky130_fd_sc_hd__dfxtp_4
X_51439_ _51436_/Y _51420_/X _51438_/X _86010_/D sky130_fd_sc_hd__a21oi_4
X_82259_ _84223_/CLK _82259_/D _82259_/Q sky130_fd_sc_hd__dfxtp_4
X_70273_ _70273_/A _70160_/X _70162_/X _70164_/X _70273_/Y sky130_fd_sc_hd__nand4_4
X_72012_ _72007_/A _72012_/B _72012_/Y sky130_fd_sc_hd__nand2_4
X_42172_ _42172_/A _42172_/Y sky130_fd_sc_hd__inv_2
X_54158_ _54149_/A _47334_/Y _54158_/Y sky130_fd_sc_hd__nand2_4
X_41123_ _81727_/Q _41079_/X _41123_/X sky130_fd_sc_hd__or2_4
X_53109_ _53115_/A _53109_/B _53109_/Y sky130_fd_sc_hd__nand2_4
X_76820_ _81493_/Q _76822_/A sky130_fd_sc_hd__inv_2
X_46980_ _46979_/Y _52785_/D sky130_fd_sc_hd__buf_2
X_58966_ _59053_/A _58966_/X sky130_fd_sc_hd__buf_2
X_54089_ _54037_/A _52571_/B _54089_/Y sky130_fd_sc_hd__nand2_4
X_86998_ _86998_/CLK _44694_/Y _86998_/Q sky130_fd_sc_hd__dfxtp_4
X_45931_ _72908_/A _45931_/X sky130_fd_sc_hd__buf_2
X_41054_ _41053_/X _41054_/X sky130_fd_sc_hd__buf_2
X_57917_ _57914_/Y _57916_/Y _57889_/X _57917_/X sky130_fd_sc_hd__a21o_4
X_76751_ _76734_/A _76749_/Y _76750_/Y _76751_/Y sky130_fd_sc_hd__a21oi_4
X_85949_ _82394_/CLK _51773_/Y _85949_/Q sky130_fd_sc_hd__dfxtp_4
X_73963_ _73963_/A _73869_/X _73963_/Y sky130_fd_sc_hd__nor2_4
X_58897_ _58897_/A _58898_/B sky130_fd_sc_hd__buf_2
X_75702_ _75687_/A _80783_/D _75701_/X _75702_/Y sky130_fd_sc_hd__o21ai_4
X_48650_ _86503_/Q _48612_/X _48649_/Y _48650_/Y sky130_fd_sc_hd__o21ai_4
X_72914_ _72881_/A _86524_/Q _72914_/X sky130_fd_sc_hd__and2_4
X_79470_ _79470_/A _79470_/B _79470_/X sky130_fd_sc_hd__or2_4
X_45862_ _74702_/B _45832_/B _45862_/Y sky130_fd_sc_hd__nand2_4
X_57848_ _57848_/A _58679_/A sky130_fd_sc_hd__buf_2
X_76682_ _76682_/A _81445_/D _76682_/X sky130_fd_sc_hd__xor2_4
X_73894_ _72979_/X _73894_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_507_0_CLK clkbuf_9_506_0_CLK/A clkbuf_9_507_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_47601_ _47363_/A _47745_/A sky130_fd_sc_hd__buf_2
X_78421_ _78420_/X _78421_/Y sky130_fd_sc_hd__inv_2
X_44813_ _41646_/Y _43939_/X _67417_/B _43941_/X _44813_/X sky130_fd_sc_hd__a2bb2o_4
X_75633_ _75631_/X _75633_/B _75633_/Y sky130_fd_sc_hd__nor2_4
X_87619_ _88387_/CLK _87619_/D _66948_/B sky130_fd_sc_hd__dfxtp_4
X_48581_ _48581_/A _48582_/A sky130_fd_sc_hd__inv_2
X_72845_ _72845_/A _72844_/X _72846_/B sky130_fd_sc_hd__nand2_4
X_45793_ _57058_/B _45793_/B _45793_/Y sky130_fd_sc_hd__nor2_4
X_57779_ _72201_/A _57779_/X sky130_fd_sc_hd__buf_2
X_47532_ _47532_/A _53103_/D sky130_fd_sc_hd__buf_2
X_59518_ _59517_/Y _59519_/C sky130_fd_sc_hd__inv_2
Xclkbuf_8_60_0_CLK clkbuf_8_61_0_CLK/A clkbuf_8_60_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_78352_ _78353_/C _78353_/B _78353_/A _78352_/X sky130_fd_sc_hd__a21o_4
X_44744_ _44744_/A _44744_/Y sky130_fd_sc_hd__inv_2
X_75564_ _80801_/Q _75564_/Y sky130_fd_sc_hd__inv_2
X_41956_ _42477_/A _41956_/X sky130_fd_sc_hd__buf_2
X_60790_ _61075_/B _60782_/Y _60403_/C _60697_/Y _60789_/Y _84567_/D
+ sky130_fd_sc_hd__a41oi_4
X_72776_ _73007_/A _72776_/X sky130_fd_sc_hd__buf_2
X_77303_ _77318_/B _77302_/Y _82183_/D sky130_fd_sc_hd__xor2_4
X_74515_ _70506_/A _70701_/A _74515_/C _74515_/X sky130_fd_sc_hd__and3_4
X_40907_ _82854_/Q _40907_/B _40907_/X sky130_fd_sc_hd__or2_4
X_47463_ _47556_/A _47463_/X sky130_fd_sc_hd__buf_2
X_71727_ _71729_/A _71680_/C _71724_/X _71727_/Y sky130_fd_sc_hd__nand3_4
X_59449_ _59442_/X _83338_/Q _59448_/Y _59449_/X sky130_fd_sc_hd__o21a_4
X_78283_ _78274_/A _78262_/A _78262_/B _78283_/Y sky130_fd_sc_hd__nand3_4
X_44675_ _44675_/A _44675_/Y sky130_fd_sc_hd__inv_2
X_75495_ _80702_/Q _80958_/D _75495_/Y sky130_fd_sc_hd__nor2_4
X_41887_ _41887_/A _41887_/X sky130_fd_sc_hd__buf_2
X_49202_ _50209_/A _49113_/B _49091_/C _49202_/X sky130_fd_sc_hd__and3_4
X_46414_ _82931_/Q _46459_/B _46414_/X sky130_fd_sc_hd__or2_4
X_77234_ _77234_/A _77233_/X _82178_/D sky130_fd_sc_hd__xor2_4
X_43626_ _40650_/X _43624_/X _73822_/A _43625_/X _43626_/X sky130_fd_sc_hd__a2bb2o_4
X_74446_ _74444_/Y _74430_/X _74445_/X _74446_/Y sky130_fd_sc_hd__a21oi_4
X_62460_ _61541_/B _62492_/B _62449_/X _62404_/X _62461_/D sky130_fd_sc_hd__nand4_4
X_40838_ _40783_/X _41014_/A _40837_/X _40839_/A sky130_fd_sc_hd__o21a_4
X_47394_ _83735_/Q _47394_/Y sky130_fd_sc_hd__inv_2
X_71658_ _71660_/A _71226_/B _71660_/C _71658_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_8_75_0_CLK clkbuf_8_75_0_CLK/A clkbuf_8_75_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_49133_ _49127_/Y _49086_/X _49132_/X _49133_/Y sky130_fd_sc_hd__a21oi_4
X_61411_ _61398_/Y _61402_/Y _61403_/X _61406_/Y _61410_/Y _61411_/X
+ sky130_fd_sc_hd__a41o_4
X_46345_ _86745_/Q _46279_/X _46344_/Y _46345_/Y sky130_fd_sc_hd__o21ai_4
X_70609_ _70609_/A _70627_/A sky130_fd_sc_hd__buf_2
X_77165_ _77159_/A _77159_/B _77173_/A _77165_/Y sky130_fd_sc_hd__a21boi_4
X_43557_ _40363_/X _43557_/X sky130_fd_sc_hd__buf_2
X_62391_ _62463_/A _62392_/D sky130_fd_sc_hd__buf_2
X_74377_ _72001_/A _74377_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_7_0_CLK clkbuf_7_6_0_CLK/A clkbuf_7_7_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_40769_ _82880_/Q _40765_/B _40769_/X sky130_fd_sc_hd__or2_4
X_71589_ _71581_/X _83447_/Q _71588_/Y _83447_/D sky130_fd_sc_hd__a21o_4
Xclkbuf_opt_5_CLK _83248_/CLK _84841_/CLK sky130_fd_sc_hd__clkbuf_16
X_64130_ _64116_/A _64087_/X _64130_/C _64130_/Y sky130_fd_sc_hd__nor3_4
X_76116_ _81725_/D _76116_/B _76127_/B sky130_fd_sc_hd__nand2_4
X_42508_ _42508_/A _42508_/Y sky130_fd_sc_hd__inv_2
X_49064_ _49064_/A _50144_/B sky130_fd_sc_hd__buf_2
X_61342_ _61313_/A _61342_/X sky130_fd_sc_hd__buf_2
X_73328_ _73325_/X _73327_/Y _73328_/Y sky130_fd_sc_hd__nand2_4
X_46276_ _46276_/A _53953_/B sky130_fd_sc_hd__buf_2
X_77096_ _77096_/A _77096_/B _77097_/B sky130_fd_sc_hd__and2_4
X_43488_ _43488_/A _43488_/Y sky130_fd_sc_hd__inv_2
X_48015_ _48014_/Y _48016_/B sky130_fd_sc_hd__buf_2
X_45227_ _45224_/Y _45226_/Y _45212_/X _45227_/X sky130_fd_sc_hd__a21o_4
X_76047_ _76047_/A _76047_/B _76048_/B sky130_fd_sc_hd__and2_4
X_64061_ _63724_/A _64158_/B sky130_fd_sc_hd__buf_2
X_42439_ _43146_/A _42439_/X sky130_fd_sc_hd__buf_2
X_61273_ _84491_/Q _61252_/X _61272_/Y _61238_/Y _61273_/X sky130_fd_sc_hd__o22a_4
X_73259_ _73257_/X _86190_/Q _73205_/X _73258_/X _73259_/X sky130_fd_sc_hd__a211o_4
X_63012_ _60562_/B _64223_/B _63347_/C _60541_/B _63012_/X sky130_fd_sc_hd__and4_4
X_60224_ _60408_/A _60095_/X _60155_/D _60185_/X _60166_/X _60224_/Y
+ sky130_fd_sc_hd__a32oi_4
X_45158_ _64401_/B _61521_/B sky130_fd_sc_hd__buf_2
X_44109_ _44108_/X _44109_/X sky130_fd_sc_hd__buf_2
X_67820_ _66572_/X _68450_/A sky130_fd_sc_hd__buf_2
X_79806_ _79806_/A _79806_/B _79807_/B sky130_fd_sc_hd__xor2_4
X_60155_ _60095_/X _60402_/A _60155_/C _60155_/D _60193_/A sky130_fd_sc_hd__and4_4
X_49966_ _49981_/A _53179_/B _49966_/Y sky130_fd_sc_hd__nand2_4
X_45089_ _56223_/C _45073_/X _45088_/X _45089_/Y sky130_fd_sc_hd__o21ai_4
X_77998_ _77998_/A _78002_/A sky130_fd_sc_hd__inv_2
Xclkbuf_8_13_0_CLK clkbuf_7_6_0_CLK/X clkbuf_9_27_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_48917_ _48995_/A _48917_/X sky130_fd_sc_hd__buf_2
X_67751_ _67987_/A _67751_/X sky130_fd_sc_hd__buf_2
X_79737_ _79728_/Y _79724_/X _79736_/X _79737_/Y sky130_fd_sc_hd__a21boi_4
X_64963_ _64877_/X _86420_/Q _64963_/X sky130_fd_sc_hd__and2_4
X_60086_ _59896_/X _62548_/B sky130_fd_sc_hd__buf_2
X_76949_ _81681_/Q _76949_/B _76949_/X sky130_fd_sc_hd__xor2_4
X_49897_ _49924_/A _49897_/X sky130_fd_sc_hd__buf_2
X_66702_ _66699_/X _66701_/X _66606_/X _66702_/X sky130_fd_sc_hd__a21o_4
X_63914_ _63848_/X _63849_/X _63914_/C _63914_/Y sky130_fd_sc_hd__nor3_4
X_48848_ _86471_/Q _48836_/X _48847_/Y _48848_/Y sky130_fd_sc_hd__o21ai_4
X_67682_ _67676_/X _67680_/X _67681_/X _67682_/X sky130_fd_sc_hd__a21o_4
X_79668_ _79657_/X _79668_/B _79668_/Y sky130_fd_sc_hd__nand2_4
X_64894_ _64691_/X _86134_/Q _64692_/X _64893_/X _64894_/X sky130_fd_sc_hd__a211o_4
X_69421_ _83925_/Q _69367_/X _69420_/X _83925_/D sky130_fd_sc_hd__a21bo_4
X_66633_ _66608_/A _66633_/X sky130_fd_sc_hd__buf_2
X_78619_ _78610_/X _78615_/X _78618_/Y _78640_/C sky130_fd_sc_hd__or3_4
X_63845_ _64184_/C _63862_/C sky130_fd_sc_hd__buf_2
X_48779_ _52166_/A _48770_/X _48786_/C _48779_/X sky130_fd_sc_hd__and3_4
X_79599_ _79588_/A _79586_/A _79585_/Y _79599_/Y sky130_fd_sc_hd__a21boi_4
Xclkbuf_8_28_0_CLK clkbuf_8_29_0_CLK/A clkbuf_9_57_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_50810_ _50799_/A _51320_/B _50810_/Y sky130_fd_sc_hd__nand2_4
X_81630_ _81275_/CLK _76591_/X _81630_/Q sky130_fd_sc_hd__dfxtp_4
X_69352_ _69300_/X _69340_/X _69350_/Y _69351_/Y _69352_/X sky130_fd_sc_hd__a211o_4
X_66564_ _69567_/A _66564_/X sky130_fd_sc_hd__buf_2
X_51790_ _51790_/A _51796_/A sky130_fd_sc_hd__buf_2
X_63776_ _64045_/A _63776_/X sky130_fd_sc_hd__buf_2
X_60988_ _60988_/A _60988_/Y sky130_fd_sc_hd__inv_2
X_68303_ _68301_/X _67842_/Y _68287_/X _68302_/Y _68303_/X sky130_fd_sc_hd__a211o_4
X_65515_ _65515_/A _65516_/A sky130_fd_sc_hd__buf_2
X_50741_ _50739_/Y _50735_/X _50740_/Y _86143_/D sky130_fd_sc_hd__a21boi_4
X_62727_ _62727_/A _62727_/B _61831_/X _62727_/Y sky130_fd_sc_hd__nand3_4
X_81561_ _81433_/CLK _81561_/D _81561_/Q sky130_fd_sc_hd__dfxtp_4
X_69283_ _69216_/X _69281_/Y _69231_/X _69282_/Y _69283_/X sky130_fd_sc_hd__a211o_4
X_66495_ _66501_/A _66501_/B _66495_/C _66495_/X sky130_fd_sc_hd__and3_4
X_83300_ _83300_/CLK _72026_/Y _83300_/Q sky130_fd_sc_hd__dfxtp_4
X_80512_ _80509_/Y _80492_/Y _80511_/X _80512_/Y sky130_fd_sc_hd__o21ai_4
X_68234_ _82653_/D _68220_/X _68233_/X _84005_/D sky130_fd_sc_hd__a21bo_4
X_53460_ _53460_/A _47853_/Y _53460_/Y sky130_fd_sc_hd__nand2_4
X_65446_ _65446_/A _65192_/B _65445_/X _65446_/Y sky130_fd_sc_hd__nand3_4
X_84280_ _84280_/CLK _64023_/Y _64022_/C sky130_fd_sc_hd__dfxtp_4
X_50672_ _52370_/A _50651_/X _50668_/C _50672_/X sky130_fd_sc_hd__and3_4
X_62658_ _62658_/A _64225_/C _60197_/C _62657_/X _62658_/X sky130_fd_sc_hd__and4_4
X_81492_ _81492_/CLK _81492_/D _76810_/A sky130_fd_sc_hd__dfxtp_4
X_52411_ _52407_/A _49181_/A _52411_/X sky130_fd_sc_hd__and2_4
X_83231_ _83231_/CLK _83231_/D _79405_/B sky130_fd_sc_hd__dfxtp_4
X_61609_ _58399_/A _61609_/X sky130_fd_sc_hd__buf_2
X_80443_ _80452_/A _80452_/B _80458_/B sky130_fd_sc_hd__xnor2_4
X_68165_ _68155_/X _67030_/Y _68148_/X _68164_/Y _68165_/X sky130_fd_sc_hd__a211o_4
X_53391_ _85642_/Q _53378_/X _53390_/Y _53391_/Y sky130_fd_sc_hd__o21ai_4
X_65377_ _58785_/A _86019_/Q _65377_/X sky130_fd_sc_hd__and2_4
X_62589_ _62622_/A _62586_/Y _62587_/Y _62589_/D _62589_/Y sky130_fd_sc_hd__nand4_4
X_55130_ _55149_/A _55135_/A sky130_fd_sc_hd__buf_2
X_67116_ _80907_/D _67092_/X _67115_/X _67116_/X sky130_fd_sc_hd__a21bo_4
X_52342_ _52339_/Y _52340_/X _52341_/X _52342_/Y sky130_fd_sc_hd__a21oi_4
X_64328_ _64328_/A _64328_/X sky130_fd_sc_hd__buf_2
X_83162_ _86570_/CLK _83162_/D _83162_/Q sky130_fd_sc_hd__dfxtp_4
X_80374_ _80366_/A _80366_/B _80361_/A _80375_/B sky130_fd_sc_hd__o21ai_4
X_68096_ _69156_/A _68097_/A sky130_fd_sc_hd__buf_2
X_82113_ _82485_/CLK _82125_/Q _77230_/B sky130_fd_sc_hd__dfxtp_4
X_55061_ _55043_/X _55056_/X _55070_/C _47710_/A _55061_/X sky130_fd_sc_hd__and4_4
X_67047_ _66972_/X _67047_/B _67047_/X sky130_fd_sc_hd__and2_4
X_52273_ _85855_/Q _52269_/X _52272_/Y _52273_/Y sky130_fd_sc_hd__o21ai_4
X_64259_ _64273_/A _64273_/B _58232_/A _64304_/D _64259_/X sky130_fd_sc_hd__and4_4
X_83093_ _83846_/CLK _74337_/X _70323_/C sky130_fd_sc_hd__dfxtp_4
X_87970_ _87720_/CLK _87970_/D _87970_/Q sky130_fd_sc_hd__dfxtp_4
X_54012_ _54010_/Y _54006_/X _54011_/Y _54012_/Y sky130_fd_sc_hd__a21boi_4
X_51224_ _51170_/A _51225_/C sky130_fd_sc_hd__buf_2
X_86921_ _86920_/CLK _86921_/D _86921_/Q sky130_fd_sc_hd__dfxtp_4
X_82044_ _82047_/CLK _77970_/B _82044_/Q sky130_fd_sc_hd__dfxtp_4
X_58820_ _58696_/X _58818_/Y _58819_/Y _58728_/X _58701_/X _58820_/X
+ sky130_fd_sc_hd__o32a_4
X_51155_ _51153_/Y _51147_/X _51154_/X _51155_/Y sky130_fd_sc_hd__a21oi_4
X_86852_ _86869_/CLK _86852_/D _63314_/B sky130_fd_sc_hd__dfxtp_4
X_68998_ _80808_/D _68954_/X _68997_/X _83952_/D sky130_fd_sc_hd__a21bo_4
X_50106_ _50106_/A _53834_/B _50106_/X sky130_fd_sc_hd__and2_4
X_85803_ _86122_/CLK _85803_/D _85803_/Q sky130_fd_sc_hd__dfxtp_4
X_58751_ _58751_/A _58764_/B _58751_/Y sky130_fd_sc_hd__nor2_4
X_51086_ _51097_/A _52777_/B _51086_/Y sky130_fd_sc_hd__nand2_4
X_55963_ _55698_/A _55963_/B _55963_/X sky130_fd_sc_hd__and2_4
X_67949_ _68714_/A _69747_/A sky130_fd_sc_hd__buf_2
X_86783_ _82317_/CLK _86783_/D _67123_/B sky130_fd_sc_hd__dfxtp_4
X_83995_ _84003_/CLK _83995_/D _82643_/D sky130_fd_sc_hd__dfxtp_4
X_57702_ _58635_/A _57872_/A sky130_fd_sc_hd__buf_2
X_50037_ _50034_/Y _50029_/X _50036_/X _86277_/D sky130_fd_sc_hd__a21oi_4
X_54914_ _54888_/A _54932_/A sky130_fd_sc_hd__buf_2
X_85734_ _85735_/CLK _52901_/Y _85734_/Q sky130_fd_sc_hd__dfxtp_4
X_70960_ _70959_/X _70961_/A sky130_fd_sc_hd__buf_2
X_82946_ _82961_/CLK _82946_/D _82946_/Q sky130_fd_sc_hd__dfxtp_4
X_58682_ _58813_/A _58682_/X sky130_fd_sc_hd__buf_2
X_55894_ _55620_/A _85239_/Q _55894_/X sky130_fd_sc_hd__and2_4
X_57633_ _57631_/Y _57627_/X _57632_/Y _84965_/D sky130_fd_sc_hd__a21boi_4
X_69619_ _64696_/A _69619_/B _69619_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_372_0_CLK clkbuf_9_186_0_CLK/X _85431_/CLK sky130_fd_sc_hd__clkbuf_1
X_54845_ _54850_/A _47623_/A _54845_/Y sky130_fd_sc_hd__nand2_4
X_85665_ _85444_/CLK _53267_/Y _85665_/Q sky130_fd_sc_hd__dfxtp_4
X_70891_ _50976_/B _70885_/X _70890_/Y _70891_/Y sky130_fd_sc_hd__o21ai_4
X_82877_ _82859_/CLK _78273_/B _82877_/Q sky130_fd_sc_hd__dfxtp_4
X_87404_ _83987_/CLK _87404_/D _87404_/Q sky130_fd_sc_hd__dfxtp_4
X_41810_ _40400_/X _41799_/X _88141_/Q _41800_/X _41810_/X sky130_fd_sc_hd__a2bb2o_4
X_72630_ _73078_/A _72630_/X sky130_fd_sc_hd__buf_2
X_84616_ _83216_/CLK _84616_/D _79156_/A sky130_fd_sc_hd__dfxtp_4
X_57564_ _57563_/X _57564_/X sky130_fd_sc_hd__buf_2
X_81828_ _82211_/CLK _81828_/D _77249_/A sky130_fd_sc_hd__dfxtp_4
X_88384_ _86796_/CLK _40486_/X _88384_/Q sky130_fd_sc_hd__dfxtp_4
X_54776_ _54773_/Y _54774_/X _54775_/X _85380_/D sky130_fd_sc_hd__a21oi_4
X_42790_ _41361_/X _42787_/X _87717_/Q _42788_/X _42790_/X sky130_fd_sc_hd__a2bb2o_4
X_85596_ _85596_/CLK _85596_/D _85596_/Q sky130_fd_sc_hd__dfxtp_4
X_51988_ _51988_/A _51972_/X _51958_/C _51988_/X sky130_fd_sc_hd__and3_4
X_59303_ _59291_/Y _59230_/X _59298_/X _59302_/X _59303_/Y sky130_fd_sc_hd__a22oi_4
X_56515_ _56528_/A _56515_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_493_0_CLK clkbuf_9_493_0_CLK/A clkbuf_9_493_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_87335_ _87345_/CLK _87335_/D _87335_/Q sky130_fd_sc_hd__dfxtp_4
X_53727_ _53725_/Y _53696_/X _53726_/Y _53727_/Y sky130_fd_sc_hd__a21boi_4
X_41741_ _41741_/A _41741_/X sky130_fd_sc_hd__buf_2
X_72561_ _72539_/B _72510_/C _72561_/C _72562_/A sky130_fd_sc_hd__and3_4
X_84547_ _84529_/CLK _84547_/D _60970_/C sky130_fd_sc_hd__dfxtp_4
X_50939_ _50938_/X _51800_/B _50939_/Y sky130_fd_sc_hd__nand2_4
X_57495_ _57499_/A _73591_/A _57495_/Y sky130_fd_sc_hd__nand2_4
X_81759_ _81783_/CLK _76136_/B _81759_/Q sky130_fd_sc_hd__dfxtp_4
X_74300_ _70285_/C _74288_/X _74299_/Y _83107_/D sky130_fd_sc_hd__a21bo_4
Xclkbuf_10_387_0_CLK clkbuf_9_193_0_CLK/X _84487_/CLK sky130_fd_sc_hd__clkbuf_1
X_59234_ _59219_/X _85742_/Q _59220_/X _59234_/X sky130_fd_sc_hd__o21a_4
X_71512_ _71512_/A _70710_/A _71512_/Y sky130_fd_sc_hd__nand2_4
X_44460_ _44447_/X _44448_/X _41138_/X _87098_/Q _44449_/X _44461_/A
+ sky130_fd_sc_hd__o32ai_4
X_56446_ _56446_/A _56446_/B _85190_/Q _56446_/Y sky130_fd_sc_hd__nand3_4
X_75280_ _75252_/Y _75251_/Y _75261_/B _75280_/X sky130_fd_sc_hd__a21bo_4
X_41672_ _41802_/A _41672_/X sky130_fd_sc_hd__buf_2
X_87266_ _88034_/CLK _43789_/X _69372_/B sky130_fd_sc_hd__dfxtp_4
X_53658_ _48752_/A _53658_/B _53667_/C _53658_/X sky130_fd_sc_hd__and3_4
X_72492_ _63598_/A _72488_/B _72492_/Y sky130_fd_sc_hd__nand2_4
X_84478_ _84481_/CLK _84478_/D _84478_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_110 sky130_fd_sc_hd__decap_3
X_43411_ _41507_/X _43396_/X _87434_/Q _43397_/X _43411_/X sky130_fd_sc_hd__a2bb2o_4
X_74231_ _74228_/X _74230_/X _74241_/A sky130_fd_sc_hd__nand2_4
X_86217_ _86218_/CLK _50357_/Y _86217_/Q sky130_fd_sc_hd__dfxtp_4
X_40623_ _48904_/A _40623_/X sky130_fd_sc_hd__buf_2
XPHY_121 sky130_fd_sc_hd__decap_3
X_52609_ _85787_/Q _52601_/X _52608_/Y _52609_/Y sky130_fd_sc_hd__o21ai_4
X_59165_ _58939_/A _59165_/X sky130_fd_sc_hd__buf_2
X_71443_ _58145_/Y _71444_/A _71442_/Y _71443_/Y sky130_fd_sc_hd__o21ai_4
X_83429_ _82386_/CLK _71640_/Y _59493_/A sky130_fd_sc_hd__dfxtp_4
X_56377_ _56370_/Y _56377_/X sky130_fd_sc_hd__buf_2
X_44391_ _44381_/X _44382_/X _41473_/X _87132_/Q _44383_/X _44392_/A
+ sky130_fd_sc_hd__o32ai_4
XPHY_132 sky130_fd_sc_hd__decap_3
X_87197_ _87446_/CLK _87197_/D _67856_/B sky130_fd_sc_hd__dfxtp_4
X_53589_ _85607_/Q _53586_/X _53588_/Y _53589_/Y sky130_fd_sc_hd__o21ai_4
XPHY_143 sky130_fd_sc_hd__decap_3
XPHY_154 sky130_fd_sc_hd__decap_3
X_58116_ _57991_/A _58116_/B _58116_/Y sky130_fd_sc_hd__nor2_4
X_46130_ _46164_/A _46087_/A _46133_/B sky130_fd_sc_hd__nor2_4
XPHY_165 sky130_fd_sc_hd__decap_3
X_43342_ _43316_/X _43319_/X _41316_/X _87469_/Q _43330_/X _43342_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74162_ _74202_/A _74161_/Y _74162_/Y sky130_fd_sc_hd__nor2_4
X_55328_ _55316_/X _55325_/X _55328_/C _55384_/A _55328_/X sky130_fd_sc_hd__and4_4
X_86148_ _83594_/CLK _86148_/D _86148_/Q sky130_fd_sc_hd__dfxtp_4
X_40554_ _40636_/A _40554_/X sky130_fd_sc_hd__buf_2
XPHY_176 sky130_fd_sc_hd__decap_3
Xclkbuf_10_310_0_CLK clkbuf_9_155_0_CLK/X _84939_/CLK sky130_fd_sc_hd__clkbuf_1
X_59096_ _59048_/X _85657_/Q _59070_/X _59096_/X sky130_fd_sc_hd__o21a_4
X_71374_ _71164_/B _71377_/B sky130_fd_sc_hd__buf_2
XPHY_187 sky130_fd_sc_hd__decap_3
XPHY_198 sky130_fd_sc_hd__decap_3
X_73113_ _72988_/X _86196_/Q _72985_/X _73112_/X _73113_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_940_0_CLK clkbuf_9_470_0_CLK/X _87577_/CLK sky130_fd_sc_hd__clkbuf_1
X_46061_ _43585_/X _46061_/X sky130_fd_sc_hd__buf_2
X_58047_ _84930_/Q _58025_/X _58040_/X _58046_/X _84930_/D sky130_fd_sc_hd__a2bb2oi_4
X_70325_ _83796_/Q _70325_/Y sky130_fd_sc_hd__inv_2
X_43273_ _43212_/A _43273_/X sky130_fd_sc_hd__buf_2
X_55259_ _57039_/A _44058_/A _55134_/X _55258_/X _55259_/X sky130_fd_sc_hd__a211o_4
X_74093_ _74117_/A _74093_/B _74093_/Y sky130_fd_sc_hd__nor2_4
X_78970_ _78957_/A _78970_/B _78970_/X sky130_fd_sc_hd__and2_4
X_86079_ _85761_/CLK _51072_/Y _86079_/Q sky130_fd_sc_hd__dfxtp_4
X_40485_ _40484_/Y _40485_/X sky130_fd_sc_hd__buf_2
X_45012_ _45237_/A _45012_/X sky130_fd_sc_hd__buf_2
X_42224_ _42259_/A _42224_/X sky130_fd_sc_hd__buf_2
X_73044_ _73041_/X _73043_/X _72877_/X _73044_/X sky130_fd_sc_hd__a21o_4
X_77921_ _77908_/A _77907_/Y _77921_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_9_431_0_CLK clkbuf_9_430_0_CLK/A clkbuf_9_431_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_70256_ _70260_/A _70260_/B _83181_/Q _70260_/D _70256_/X sky130_fd_sc_hd__and4_4
X_49820_ _49809_/A _53033_/B _49820_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_325_0_CLK clkbuf_9_162_0_CLK/X _85635_/CLK sky130_fd_sc_hd__clkbuf_1
X_42155_ _42154_/X _42141_/X _41174_/X _88007_/Q _42142_/X _42155_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77852_ _82272_/Q _81984_/Q _77852_/Y sky130_fd_sc_hd__xnor2_4
X_70187_ _70233_/A _70200_/D sky130_fd_sc_hd__buf_2
X_59998_ _60543_/B _59998_/B _59951_/C _59977_/Y _59998_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_10_955_0_CLK clkbuf_9_477_0_CLK/X _87821_/CLK sky130_fd_sc_hd__clkbuf_1
X_41106_ _82274_/Q _41102_/B _41106_/X sky130_fd_sc_hd__or2_4
X_76803_ _81491_/Q _76805_/A sky130_fd_sc_hd__inv_2
X_49751_ _49751_/A _49750_/X _49761_/C _52967_/D _49751_/X sky130_fd_sc_hd__and4_4
X_46963_ _82397_/Q _46964_/A sky130_fd_sc_hd__inv_2
X_42086_ _40982_/X _42072_/X _88042_/Q _42073_/X _42086_/X sky130_fd_sc_hd__a2bb2o_4
X_58949_ _58846_/X _85763_/Q _58847_/X _58949_/X sky130_fd_sc_hd__o21a_4
X_77783_ _77777_/Y _77778_/X _77782_/Y _77783_/Y sky130_fd_sc_hd__a21oi_4
X_74995_ _80766_/Q _74995_/B _74995_/Y sky130_fd_sc_hd__nand2_4
X_48702_ _48702_/A _48894_/B _48894_/C _48702_/X sky130_fd_sc_hd__and3_4
Xclkbuf_9_446_0_CLK clkbuf_9_446_0_CLK/A clkbuf_9_446_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_79522_ _79522_/A _79522_/B _82849_/D sky130_fd_sc_hd__nand2_4
X_45914_ DATA_AVAILABLE _80673_/Q _45913_/Y _86843_/D sky130_fd_sc_hd__o21a_4
X_41037_ _40995_/A _41037_/X sky130_fd_sc_hd__buf_2
X_76734_ _76734_/A _76736_/A sky130_fd_sc_hd__inv_2
X_49682_ _49661_/X _47174_/X _49682_/Y sky130_fd_sc_hd__nand2_4
X_61960_ _61960_/A _61960_/B _78066_/B _61960_/Y sky130_fd_sc_hd__nor3_4
X_73946_ _88355_/Q _73801_/X _73087_/X _73946_/Y sky130_fd_sc_hd__o21ai_4
X_46894_ _82948_/Q _46894_/Y sky130_fd_sc_hd__inv_2
X_48633_ _48563_/X _48086_/A _48632_/Y _48634_/A sky130_fd_sc_hd__o21ai_4
X_60911_ _60910_/X _60911_/X sky130_fd_sc_hd__buf_2
X_79453_ _79446_/X _79453_/B _79453_/Y sky130_fd_sc_hd__nand2_4
X_45845_ _45841_/X _45844_/X _44898_/X _45845_/X sky130_fd_sc_hd__a21o_4
X_76665_ _76665_/A _81443_/D _81539_/D sky130_fd_sc_hd__xor2_4
X_61891_ _58319_/A _61891_/X sky130_fd_sc_hd__buf_2
X_73877_ _86994_/Q _73776_/X _73876_/X _73888_/C sky130_fd_sc_hd__o21ai_4
X_78404_ _78408_/C _78404_/Y sky130_fd_sc_hd__inv_2
X_63630_ _63630_/A _63630_/B _63630_/C _63630_/Y sky130_fd_sc_hd__nor3_4
X_75616_ _75616_/A _75615_/Y _75617_/B sky130_fd_sc_hd__xnor2_4
X_48564_ _81775_/Q _49067_/B sky130_fd_sc_hd__inv_2
X_60842_ _59539_/A _59557_/X _59564_/B _59901_/C _59877_/X _61071_/A
+ sky130_fd_sc_hd__a41oi_4
X_72828_ _74012_/A _72829_/A sky130_fd_sc_hd__buf_2
X_79384_ _84805_/Q _84125_/Q _79384_/X sky130_fd_sc_hd__xor2_4
X_45776_ _45775_/Y _44975_/A _45776_/X sky130_fd_sc_hd__and2_4
X_76596_ _76595_/Y _76596_/Y sky130_fd_sc_hd__inv_2
X_42988_ _42984_/X _42985_/X _40480_/X _66995_/B _42976_/X _42988_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47515_ _47515_/A _47516_/A sky130_fd_sc_hd__inv_2
X_78335_ _78335_/A _78335_/B _78335_/Y sky130_fd_sc_hd__nand2_4
X_44727_ _44727_/A _44727_/Y sky130_fd_sc_hd__inv_2
X_75547_ _75537_/Y _75538_/B _75539_/X _75547_/Y sky130_fd_sc_hd__o21ai_4
X_63561_ _63523_/A _63561_/B _63561_/X sky130_fd_sc_hd__and2_4
X_41939_ _41967_/A _41939_/X sky130_fd_sc_hd__buf_2
X_48495_ _81781_/Q _48495_/Y sky130_fd_sc_hd__inv_2
X_60773_ _60543_/B _60727_/A _60772_/Y _60725_/B _60773_/Y sky130_fd_sc_hd__nand4_4
X_72759_ _72758_/X _86529_/Q _72759_/X sky130_fd_sc_hd__and2_4
X_65300_ _57965_/A _65300_/X sky130_fd_sc_hd__buf_2
X_62512_ _62500_/X _62506_/Y _62510_/X _84845_/Q _62511_/X _62512_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47446_ _81802_/Q _54743_/D sky130_fd_sc_hd__inv_2
X_66280_ _66231_/X _66319_/B _84144_/Q _66280_/X sky130_fd_sc_hd__and3_4
X_78266_ _78265_/A _82467_/Q _78266_/Y sky130_fd_sc_hd__nor2_4
X_44658_ _44679_/A _44658_/X sky130_fd_sc_hd__buf_2
X_63492_ _63434_/X _63485_/X _63486_/X _63490_/X _63491_/Y _63492_/Y
+ sky130_fd_sc_hd__o41ai_4
XPHY_1 sky130_fd_sc_hd__decap_3
X_75478_ _75477_/B _75477_/C _75477_/A _75478_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_5_10_0_CLK clkbuf_4_5_1_CLK/X clkbuf_6_21_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_65231_ _65206_/A _86441_/Q _65231_/X sky130_fd_sc_hd__and2_4
X_77217_ _77217_/A _77217_/B _77217_/Y sky130_fd_sc_hd__nand2_4
X_43609_ _43585_/X _43609_/X sky130_fd_sc_hd__buf_2
X_62443_ _62441_/Y _62396_/X _62442_/Y _84410_/D sky130_fd_sc_hd__a21oi_4
X_74429_ _83068_/Q _74412_/X _74428_/Y _74429_/Y sky130_fd_sc_hd__o21ai_4
X_47377_ _47565_/A _47377_/X sky130_fd_sc_hd__buf_2
X_78197_ _78197_/A _78197_/B _78197_/X sky130_fd_sc_hd__xor2_4
X_44589_ _44567_/A _44589_/X sky130_fd_sc_hd__buf_2
X_49116_ _72072_/B _50169_/B sky130_fd_sc_hd__buf_2
X_46328_ _82939_/Q _46328_/B _46328_/X sky130_fd_sc_hd__or2_4
X_65162_ _65156_/X _65160_/X _65161_/X _65162_/X sky130_fd_sc_hd__a21o_4
X_77148_ _77157_/A _77157_/B _77151_/A sky130_fd_sc_hd__xor2_4
X_62374_ _62532_/A _62375_/C sky130_fd_sc_hd__buf_2
Xclkbuf_10_908_0_CLK clkbuf_9_454_0_CLK/X _88345_/CLK sky130_fd_sc_hd__clkbuf_1
X_64113_ _63280_/B _60967_/X _64112_/Y _64113_/X sky130_fd_sc_hd__a21bo_4
X_49047_ _86449_/Q _49003_/X _49046_/Y _49047_/Y sky130_fd_sc_hd__o21ai_4
X_61325_ _61298_/Y _61305_/Y _61315_/Y _61320_/Y _61324_/Y _61325_/Y
+ sky130_fd_sc_hd__a41oi_4
X_46259_ _46259_/A _46347_/A sky130_fd_sc_hd__buf_2
X_65093_ _65090_/Y _65070_/X _65092_/X _84215_/D sky130_fd_sc_hd__a21o_4
X_69970_ _42063_/A _69582_/X _66564_/X _69969_/Y _69970_/X sky130_fd_sc_hd__a211o_4
X_77079_ _77084_/A _77073_/A _77078_/Y _77079_/Y sky130_fd_sc_hd__a21boi_4
Xclkbuf_5_25_0_CLK clkbuf_4_12_1_CLK/X clkbuf_6_51_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_68921_ _87485_/Q _68870_/X _68871_/X _68920_/X _68921_/X sky130_fd_sc_hd__a211o_4
X_64044_ _64434_/B _64145_/B _64029_/C _64029_/D _64044_/Y sky130_fd_sc_hd__nand4_4
X_61256_ _64203_/B _61256_/Y sky130_fd_sc_hd__inv_2
X_80090_ _84938_/Q _84186_/Q _80092_/A sky130_fd_sc_hd__xor2_4
X_60207_ _60159_/A _60324_/C _60218_/A _60205_/X _61286_/A _60207_/Y
+ sky130_fd_sc_hd__a41oi_4
X_68852_ _68849_/X _68851_/X _68806_/X _68852_/X sky130_fd_sc_hd__a21o_4
X_61187_ _61107_/X _61109_/X _61172_/A _61188_/C sky130_fd_sc_hd__nand3_4
X_67803_ _67800_/X _67802_/X _67709_/X _67803_/Y sky130_fd_sc_hd__a21oi_4
X_60138_ _59985_/X _60091_/A _59966_/Y _60138_/Y sky130_fd_sc_hd__o21ai_4
X_49949_ _49955_/A _53161_/B _49949_/Y sky130_fd_sc_hd__nand2_4
X_68783_ _68780_/X _68782_/X _68684_/X _68783_/X sky130_fd_sc_hd__a21o_4
X_65995_ _65876_/X _85627_/Q _65976_/X _65994_/X _65995_/X sky130_fd_sc_hd__a211o_4
X_82800_ _82833_/CLK _82800_/D _82800_/Q sky130_fd_sc_hd__dfxtp_4
X_67734_ _67731_/X _67733_/X _67709_/X _67734_/Y sky130_fd_sc_hd__a21oi_4
X_52960_ _85723_/Q _52957_/X _52959_/Y _52960_/Y sky130_fd_sc_hd__o21ai_4
X_64946_ _64946_/A _85844_/Q _64946_/X sky130_fd_sc_hd__and2_4
X_60069_ _45943_/A _59901_/A _59901_/C _63001_/A _57754_/X _60069_/Y
+ sky130_fd_sc_hd__a41oi_4
X_83780_ _83783_/CLK _83780_/D _83780_/Q sky130_fd_sc_hd__dfxtp_4
X_80992_ _80821_/CLK _80992_/D _80948_/D sky130_fd_sc_hd__dfxtp_4
X_51911_ _51902_/A _46899_/X _51911_/Y sky130_fd_sc_hd__nand2_4
X_82731_ _84115_/CLK _84115_/Q _78889_/A sky130_fd_sc_hd__dfxtp_4
X_67665_ _67569_/X _87717_/Q _67665_/X sky130_fd_sc_hd__and2_4
X_52891_ _52754_/A _52892_/A sky130_fd_sc_hd__buf_2
X_64877_ _64602_/A _64877_/X sky130_fd_sc_hd__buf_2
X_69404_ _69814_/A _69733_/A sky130_fd_sc_hd__buf_2
X_54630_ _54625_/A _54645_/B _54618_/X _54630_/D _54630_/X sky130_fd_sc_hd__and4_4
X_66616_ _66689_/A _66616_/B _66616_/X sky130_fd_sc_hd__and2_4
X_85450_ _85773_/CLK _85450_/D _85450_/Q sky130_fd_sc_hd__dfxtp_4
X_51842_ _51842_/A _51843_/A sky130_fd_sc_hd__buf_2
X_63828_ _61387_/X _63877_/B _63814_/C _63877_/D _63828_/Y sky130_fd_sc_hd__nand4_4
X_82662_ _82665_/CLK _78358_/B _78107_/A sky130_fd_sc_hd__dfxtp_4
X_67596_ _67572_/A _67596_/B _67596_/X sky130_fd_sc_hd__and2_4
X_84401_ _83242_/CLK _84401_/D _84401_/Q sky130_fd_sc_hd__dfxtp_4
X_81613_ _81620_/CLK _76312_/B _81613_/Q sky130_fd_sc_hd__dfxtp_4
X_69335_ _69128_/X _88293_/Q _69335_/X sky130_fd_sc_hd__and2_4
X_54561_ _54546_/A _53386_/B _54561_/Y sky130_fd_sc_hd__nand2_4
X_66547_ _66547_/A _66547_/X sky130_fd_sc_hd__buf_2
X_85381_ _85381_/CLK _54771_/Y _85381_/Q sky130_fd_sc_hd__dfxtp_4
X_51773_ _51771_/Y _51767_/X _51772_/X _51773_/Y sky130_fd_sc_hd__a21oi_4
X_63759_ _63747_/Y _63759_/B _63757_/Y _63758_/Y _63759_/X sky130_fd_sc_hd__and4_4
X_82593_ _81216_/CLK _82625_/Q _82593_/Q sky130_fd_sc_hd__dfxtp_4
X_56300_ _56026_/X _56290_/X _56299_/Y _85245_/D sky130_fd_sc_hd__o21ai_4
X_87120_ _87137_/CLK _87120_/D _87120_/Q sky130_fd_sc_hd__dfxtp_4
X_53512_ _48234_/A _53697_/B _53697_/C _53512_/Y sky130_fd_sc_hd__nand3_4
X_84332_ _82272_/CLK _63337_/Y _79183_/B sky130_fd_sc_hd__dfxtp_4
X_50724_ _50724_/A _50751_/B sky130_fd_sc_hd__buf_2
X_57280_ _44286_/Y _57280_/X sky130_fd_sc_hd__buf_2
X_81544_ _81532_/CLK _81544_/D _76533_/B sky130_fd_sc_hd__dfxtp_4
X_69266_ _87030_/Q _69182_/X _69183_/X _69265_/X _69266_/X sky130_fd_sc_hd__a211o_4
X_54492_ _85432_/Q _54485_/X _54491_/Y _54492_/Y sky130_fd_sc_hd__o21ai_4
X_66478_ _84115_/Q _66478_/Y sky130_fd_sc_hd__inv_2
X_56231_ _45369_/A _56245_/A sky130_fd_sc_hd__buf_2
X_68217_ _67347_/X _67350_/X _68216_/X _68217_/Y sky130_fd_sc_hd__a21oi_4
X_87051_ _87553_/CLK _44572_/Y _87051_/Q sky130_fd_sc_hd__dfxtp_4
X_65429_ _65408_/A _86529_/Q _65429_/X sky130_fd_sc_hd__and2_4
X_53443_ _53443_/A _47830_/Y _54067_/A _53443_/Y sky130_fd_sc_hd__nand3_4
X_84263_ _84263_/CLK _84263_/D _79863_/B sky130_fd_sc_hd__dfxtp_4
X_50655_ _50655_/A _50728_/A sky130_fd_sc_hd__buf_2
X_81475_ _81475_/CLK _81475_/D _76659_/A sky130_fd_sc_hd__dfxtp_4
X_69197_ _87035_/Q _69182_/X _69183_/X _69196_/X _69197_/X sky130_fd_sc_hd__a211o_4
X_86002_ _85712_/CLK _86002_/D _86002_/Q sky130_fd_sc_hd__dfxtp_4
X_83214_ _83231_/CLK _72620_/Y _72617_/A sky130_fd_sc_hd__dfxtp_4
X_56162_ _56167_/B _56167_/A _56162_/X sky130_fd_sc_hd__and2_4
X_80426_ _80416_/A _80416_/B _80411_/Y _80414_/Y _80426_/X sky130_fd_sc_hd__o22a_4
X_68148_ _68089_/A _68148_/X sky130_fd_sc_hd__buf_2
X_53374_ _85645_/Q _53351_/X _53373_/Y _53374_/Y sky130_fd_sc_hd__o21ai_4
X_84194_ _84194_/CLK _65547_/X _65546_/C sky130_fd_sc_hd__dfxtp_4
X_50586_ _50607_/A _52287_/B _50586_/Y sky130_fd_sc_hd__nand2_4
X_55113_ _55111_/Y _55102_/X _55112_/X _55113_/Y sky130_fd_sc_hd__a21oi_4
X_52325_ _52271_/A _52334_/A sky130_fd_sc_hd__buf_2
X_83145_ _83145_/CLK _83145_/D _83145_/Q sky130_fd_sc_hd__dfxtp_4
X_56093_ _56171_/A _56171_/C _56093_/C _56094_/A sky130_fd_sc_hd__nand3_4
X_68079_ _87892_/Q _68006_/X _67984_/X _68078_/X _68079_/X sky130_fd_sc_hd__a211o_4
X_80357_ _84688_/Q _80357_/B _80357_/X sky130_fd_sc_hd__xor2_4
X_70110_ _70110_/A _70112_/C sky130_fd_sc_hd__inv_2
X_55044_ _55043_/X _55030_/X _55026_/C _47682_/Y _55044_/X sky130_fd_sc_hd__and4_4
X_59921_ _62515_/C _59922_/C sky130_fd_sc_hd__buf_2
X_52256_ _65890_/B _52184_/X _52255_/Y _52256_/Y sky130_fd_sc_hd__o21ai_4
X_71090_ _71090_/A _71091_/B sky130_fd_sc_hd__buf_2
X_83076_ _83313_/CLK _74392_/Y _83076_/Q sky130_fd_sc_hd__dfxtp_4
X_87953_ _87950_/CLK _42261_/X _87953_/Q sky130_fd_sc_hd__dfxtp_4
X_80288_ _80288_/A _80288_/B _80304_/A sky130_fd_sc_hd__nor2_4
X_51207_ _51191_/X _51203_/B _51197_/C _52900_/D _51207_/X sky130_fd_sc_hd__and4_4
X_70041_ _68783_/X _68786_/X _70005_/X _70041_/Y sky130_fd_sc_hd__a21oi_4
X_86904_ _84407_/CLK _45024_/Y _64294_/B sky130_fd_sc_hd__dfxtp_4
X_82027_ _81975_/CLK _77812_/B _82027_/Q sky130_fd_sc_hd__dfxtp_4
X_59852_ _59852_/A _59855_/B sky130_fd_sc_hd__buf_2
X_52187_ _85872_/Q _52184_/X _52186_/Y _52187_/Y sky130_fd_sc_hd__o21ai_4
X_87884_ _88144_/CLK _87884_/D _87884_/Q sky130_fd_sc_hd__dfxtp_4
X_58803_ _58792_/Y _58739_/X _58799_/X _58802_/X _58803_/Y sky130_fd_sc_hd__a22oi_4
X_51138_ _51135_/Y _51119_/X _51137_/X _51138_/Y sky130_fd_sc_hd__a21oi_4
X_86835_ _87995_/CLK _86835_/D _66644_/B sky130_fd_sc_hd__dfxtp_4
X_59783_ _59689_/B _59631_/B _59687_/A _59836_/D _59782_/X _59783_/Y
+ sky130_fd_sc_hd__a41oi_4
X_56995_ _56995_/A _56995_/X sky130_fd_sc_hd__buf_2
X_73800_ _73796_/X _73798_/X _73799_/X _73815_/B sky130_fd_sc_hd__a21o_4
X_58734_ _58618_/X _86100_/Q _58733_/X _58734_/Y sky130_fd_sc_hd__o21ai_4
X_43960_ _59538_/D _44003_/A sky130_fd_sc_hd__buf_2
X_51069_ _51058_/A _52760_/B _51069_/Y sky130_fd_sc_hd__nand2_4
X_55946_ _55946_/A _74297_/C sky130_fd_sc_hd__buf_2
Xclkbuf_7_123_0_CLK clkbuf_6_61_0_CLK/X clkbuf_8_247_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_74780_ _74780_/A _74720_/C _74744_/X _74780_/D _74784_/A sky130_fd_sc_hd__nand4_4
X_86766_ _84549_/CLK _46180_/Y _44008_/A sky130_fd_sc_hd__dfxtp_4
X_71992_ _83306_/Q _71985_/X _71991_/Y _71992_/Y sky130_fd_sc_hd__o21ai_4
X_83978_ _88376_/CLK _68341_/X _82626_/D sky130_fd_sc_hd__dfxtp_4
X_42911_ _41693_/X _42900_/X _87656_/Q _42901_/X _42911_/X sky130_fd_sc_hd__a2bb2o_4
X_73731_ _73355_/A _73731_/X sky130_fd_sc_hd__buf_2
X_85717_ _85718_/CLK _52994_/Y _85717_/Q sky130_fd_sc_hd__dfxtp_4
X_58665_ _58641_/X _85945_/Q _58664_/X _58665_/X sky130_fd_sc_hd__o21a_4
X_70943_ _49212_/B _70937_/X _70942_/Y _70943_/Y sky130_fd_sc_hd__o21ai_4
X_82929_ _81190_/CLK _78240_/X _46436_/A sky130_fd_sc_hd__dfxtp_4
X_43891_ _43890_/Y _43891_/Y sky130_fd_sc_hd__inv_2
X_55877_ _56407_/C _55505_/X _55513_/X _55876_/X _55877_/X sky130_fd_sc_hd__a211o_4
X_86697_ _86697_/CLK _86697_/D _86697_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_93_0_CLK clkbuf_9_46_0_CLK/X clkbuf_opt_9_CLK/A sky130_fd_sc_hd__clkbuf_1
X_57616_ _57563_/X _71957_/A sky130_fd_sc_hd__buf_2
X_45630_ _45626_/Y _45627_/X _45548_/X _45629_/Y _45630_/X sky130_fd_sc_hd__a211o_4
X_76450_ _81271_/Q _81539_/Q _76455_/A sky130_fd_sc_hd__nor2_4
X_42842_ _41507_/X _42830_/X _87690_/Q _42832_/X _42842_/X sky130_fd_sc_hd__a2bb2o_4
X_54828_ _85370_/Q _54812_/X _54827_/Y _54828_/Y sky130_fd_sc_hd__o21ai_4
X_73662_ _73638_/A _86589_/Q _73662_/X sky130_fd_sc_hd__and2_4
X_85648_ _85648_/CLK _85648_/D _85648_/Q sky130_fd_sc_hd__dfxtp_4
X_70874_ _46740_/X _70855_/A _70873_/Y _70874_/Y sky130_fd_sc_hd__o21ai_4
X_58596_ _58140_/X _86111_/Q _58595_/X _58596_/Y sky130_fd_sc_hd__o21ai_4
X_75401_ _75401_/A _75399_/Y _75397_/Y _75401_/Y sky130_fd_sc_hd__nand3_4
X_72613_ _79245_/B _72590_/X _72608_/Y _72612_/X _72613_/X sky130_fd_sc_hd__o22a_4
X_45561_ _45714_/A _45561_/X sky130_fd_sc_hd__buf_2
X_57547_ _84981_/Q _57527_/X _57546_/Y _57547_/Y sky130_fd_sc_hd__o21ai_4
X_76381_ _76381_/A _76381_/B _76382_/A sky130_fd_sc_hd__and2_4
X_42773_ _42773_/A _42773_/Y sky130_fd_sc_hd__inv_2
X_88367_ _86982_/CLK _40607_/Y _88367_/Q sky130_fd_sc_hd__dfxtp_4
X_54759_ _54758_/X _47469_/A _54759_/Y sky130_fd_sc_hd__nand2_4
X_73593_ _74117_/A _73592_/Y _73593_/Y sky130_fd_sc_hd__nor2_4
X_85579_ _86500_/CLK _53735_/Y _85579_/Q sky130_fd_sc_hd__dfxtp_4
X_47300_ _57846_/A _47286_/X _47299_/Y _47300_/Y sky130_fd_sc_hd__o21ai_4
X_78120_ _78120_/A _78120_/B _78120_/C _78120_/Y sky130_fd_sc_hd__nand3_4
X_44512_ _44512_/A _44512_/X sky130_fd_sc_hd__buf_2
X_75332_ _80692_/Q _80948_/D _75333_/A sky130_fd_sc_hd__nand2_4
X_41724_ _41721_/X _41722_/X _88162_/Q _41723_/X _88162_/D sky130_fd_sc_hd__a2bb2o_4
X_87318_ _87577_/CLK _87318_/D _74226_/A sky130_fd_sc_hd__dfxtp_4
X_48280_ _66171_/B _48241_/X _48279_/Y _48280_/Y sky130_fd_sc_hd__o21ai_4
X_72544_ _72573_/A _72544_/B _79467_/B _72544_/Y sky130_fd_sc_hd__nor3_4
X_45492_ _45487_/X _45491_/X _45446_/X _45492_/X sky130_fd_sc_hd__a21o_4
X_57478_ _57478_/A _57478_/Y sky130_fd_sc_hd__inv_2
X_88298_ _88301_/CLK _88298_/D _69265_/B sky130_fd_sc_hd__dfxtp_4
X_59217_ _59160_/X _85647_/Q _59205_/X _59217_/X sky130_fd_sc_hd__o21a_4
X_47231_ _54097_/B _52931_/B sky130_fd_sc_hd__buf_2
X_78051_ _84556_/Q _78051_/B _78051_/X sky130_fd_sc_hd__xor2_4
X_44443_ _44425_/X _44427_/X _41621_/X _87105_/Q _44428_/X _44444_/A
+ sky130_fd_sc_hd__o32ai_4
X_56429_ _56431_/A _56433_/B _85197_/Q _56429_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_8_254_0_CLK clkbuf_8_255_0_CLK/A clkbuf_9_509_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_75263_ _75226_/Y _75228_/X _75240_/X _75263_/X sky130_fd_sc_hd__a21o_4
X_87249_ _87249_/CLK _87249_/D _68427_/B sky130_fd_sc_hd__dfxtp_4
X_41655_ _41628_/X _41310_/A _41654_/X _41655_/X sky130_fd_sc_hd__o21a_4
X_72475_ _72414_/X _72475_/B _72475_/Y sky130_fd_sc_hd__nor2_4
X_77002_ _81986_/Q _82274_/D _77002_/X sky130_fd_sc_hd__xor2_4
X_74214_ _73165_/A _66310_/B _74214_/X sky130_fd_sc_hd__and2_4
X_40606_ _40550_/X _40556_/X _40605_/X _88367_/Q _40568_/X _40607_/A
+ sky130_fd_sc_hd__o32ai_4
X_47162_ _54580_/D _52887_/D sky130_fd_sc_hd__buf_2
X_59148_ _59146_/X _85429_/Q _59147_/X _59148_/Y sky130_fd_sc_hd__o21ai_4
X_71426_ _70370_/A _71432_/A sky130_fd_sc_hd__buf_2
X_44374_ _44350_/X _44351_/X _41773_/X _87140_/Q _44353_/X _44374_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75194_ _75162_/B _75180_/A _75179_/A _75194_/X sky130_fd_sc_hd__o21a_4
X_41586_ _41585_/Y _41586_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_31_0_CLK clkbuf_9_15_0_CLK/X _82980_/CLK sky130_fd_sc_hd__clkbuf_1
X_46113_ _46138_/A _46120_/A sky130_fd_sc_hd__buf_2
X_43325_ _43287_/A _43325_/X sky130_fd_sc_hd__buf_2
X_74145_ _74145_/A _72795_/A _74145_/Y sky130_fd_sc_hd__nor2_4
X_40537_ _40504_/X _82308_/Q _40536_/X _40537_/Y sky130_fd_sc_hd__o21ai_4
X_47093_ _47093_/A _52853_/D sky130_fd_sc_hd__buf_2
X_71357_ _71504_/C _71351_/X _71427_/C _71363_/D _71357_/X sky130_fd_sc_hd__and4_4
X_59079_ _64565_/A _64776_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_370_0_CLK clkbuf_9_370_0_CLK/A clkbuf_9_370_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_61110_ _61230_/C _61107_/X _61109_/X _61110_/Y sky130_fd_sc_hd__o21ai_4
X_70308_ _70296_/X _70297_/X _83098_/Q _70301_/D _70308_/X sky130_fd_sc_hd__and4_4
X_46044_ _45975_/X _46044_/X sky130_fd_sc_hd__buf_2
X_43256_ _43241_/X _43244_/X _41076_/X _87514_/Q _43250_/X _43256_/Y
+ sky130_fd_sc_hd__o32ai_4
X_62090_ _62050_/X _62090_/B _78057_/B _62090_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_10_264_0_CLK clkbuf_9_132_0_CLK/X _84829_/CLK sky130_fd_sc_hd__clkbuf_1
X_78953_ _78953_/A _82513_/D sky130_fd_sc_hd__inv_2
X_74076_ _74072_/X _74075_/X _73489_/X _74079_/A sky130_fd_sc_hd__a21o_4
X_40468_ _40463_/X _81169_/Q _40467_/X _40468_/Y sky130_fd_sc_hd__o21ai_4
X_71288_ _71287_/Y _71289_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_894_0_CLK clkbuf_9_447_0_CLK/X _85536_/CLK sky130_fd_sc_hd__clkbuf_1
X_42207_ _42206_/Y _87980_/D sky130_fd_sc_hd__inv_2
X_61041_ _64172_/C _64182_/C _60992_/X _60014_/X _60111_/X _61041_/Y
+ sky130_fd_sc_hd__a32oi_4
X_77904_ _77904_/A _77903_/Y _82037_/D sky130_fd_sc_hd__xor2_4
X_73027_ _73067_/A _73704_/A sky130_fd_sc_hd__buf_2
X_70239_ _70239_/A _70239_/B _70239_/C _70239_/D _70239_/X sky130_fd_sc_hd__and4_4
X_43187_ _43162_/X _43167_/X _40894_/X _73374_/A _43172_/X _43188_/A
+ sky130_fd_sc_hd__o32ai_4
X_78884_ _82843_/Q _82555_/Q _78885_/B sky130_fd_sc_hd__xnor2_4
X_40399_ _40381_/X _81179_/Q _40398_/X _40399_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_46_0_CLK clkbuf_9_23_0_CLK/X _83835_/CLK sky130_fd_sc_hd__clkbuf_1
X_49803_ _49801_/Y _49787_/X _49802_/X _86321_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_385_0_CLK clkbuf_8_192_0_CLK/X clkbuf_9_385_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_42138_ _41912_/A _42138_/X sky130_fd_sc_hd__buf_2
X_77835_ _77835_/A _77835_/B _77836_/B sky130_fd_sc_hd__and2_4
X_47995_ _52573_/B _48069_/B sky130_fd_sc_hd__buf_2
X_64800_ _64800_/A _64800_/B _64800_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_279_0_CLK clkbuf_9_139_0_CLK/X _85499_/CLK sky130_fd_sc_hd__clkbuf_1
X_49734_ _49751_/A _49724_/B _49724_/C _52948_/D _49734_/X sky130_fd_sc_hd__and4_4
X_46946_ _83718_/Q _54460_/B sky130_fd_sc_hd__inv_2
X_42069_ _40955_/X _41907_/X _88048_/Q _41912_/X _88048_/D sky130_fd_sc_hd__a2bb2o_4
X_65780_ _65717_/X _85578_/Q _65718_/X _65779_/X _65780_/X sky130_fd_sc_hd__a211o_4
X_77766_ _77759_/Y _77764_/Y _77765_/Y _77766_/Y sky130_fd_sc_hd__a21oi_4
X_62992_ _62642_/Y _62990_/Y _62991_/X _58374_/A _62650_/X _62992_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74978_ _80948_/Q _74978_/B _74978_/X sky130_fd_sc_hd__xor2_4
X_79505_ _79505_/A _79505_/B _79505_/Y sky130_fd_sc_hd__nand2_4
X_64731_ _64731_/A _64732_/A sky130_fd_sc_hd__buf_2
X_76717_ _76697_/Y _76712_/A _76719_/A sky130_fd_sc_hd__nor2_4
X_49665_ _49663_/Y _49650_/X _49664_/X _49665_/Y sky130_fd_sc_hd__a21oi_4
X_61943_ _61960_/A _61960_/B _78067_/B _61943_/Y sky130_fd_sc_hd__nor3_4
X_73929_ _73926_/X _73928_/X _72735_/X _73933_/A sky130_fd_sc_hd__a21o_4
X_46877_ _46873_/Y _46844_/X _46876_/X _86694_/D sky130_fd_sc_hd__a21oi_4
X_77697_ _77676_/A _77673_/Y _77675_/A _77701_/A sky130_fd_sc_hd__o21a_4
X_48616_ _48661_/A _52216_/B _48616_/Y sky130_fd_sc_hd__nand2_4
X_79436_ _79436_/A _79436_/B _79444_/B sky130_fd_sc_hd__xor2_4
Xclkbuf_8_207_0_CLK clkbuf_8_207_0_CLK/A clkbuf_9_415_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_67450_ _67093_/X _67497_/A sky130_fd_sc_hd__buf_2
X_45828_ _45826_/Y _45570_/X _44875_/X _45827_/Y _45828_/X sky130_fd_sc_hd__a211o_4
X_64662_ _64939_/A _64662_/X sky130_fd_sc_hd__buf_2
X_76648_ _76648_/A _76965_/A _76649_/B sky130_fd_sc_hd__xor2_4
Xclkbuf_10_202_0_CLK clkbuf_9_101_0_CLK/X _81084_/CLK sky130_fd_sc_hd__clkbuf_1
X_49596_ _49570_/A _49596_/X sky130_fd_sc_hd__buf_2
X_61874_ _61438_/X _61874_/B _61809_/C _61874_/D _61879_/B sky130_fd_sc_hd__nand4_4
X_66401_ _79435_/B _66402_/C sky130_fd_sc_hd__inv_2
Xclkbuf_10_832_0_CLK clkbuf_9_416_0_CLK/X _84220_/CLK sky130_fd_sc_hd__clkbuf_1
X_63613_ _58452_/A _63600_/X _63575_/C _63661_/D _63613_/Y sky130_fd_sc_hd__nand4_4
X_48547_ _48541_/Y _48517_/X _48546_/X _48547_/Y sky130_fd_sc_hd__a21oi_4
X_60825_ _60736_/X _60804_/C _63389_/B _63389_/D _63130_/A _60825_/Y
+ sky130_fd_sc_hd__a41oi_4
X_67381_ _67381_/A _67381_/B _67381_/X sky130_fd_sc_hd__and2_4
X_79367_ _79358_/Y _79354_/X _79366_/X _79368_/B sky130_fd_sc_hd__a21boi_4
X_45759_ _85130_/Q _45709_/X _45743_/X _45759_/X sky130_fd_sc_hd__o21a_4
X_64593_ _64593_/A _86273_/Q _64593_/X sky130_fd_sc_hd__and2_4
X_76579_ _76578_/X _76579_/Y sky130_fd_sc_hd__inv_2
X_69120_ _69117_/X _69119_/X _60014_/X _69120_/Y sky130_fd_sc_hd__a21oi_4
X_66332_ _66177_/A _66389_/B _66332_/C _66332_/Y sky130_fd_sc_hd__nor3_4
X_78318_ _78318_/A _78318_/B _78335_/B _78335_/A sky130_fd_sc_hd__nand3_4
X_63544_ _63542_/Y _63516_/X _63543_/Y _63544_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_323_0_CLK clkbuf_9_323_0_CLK/A clkbuf_9_323_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_60756_ _60707_/X _60692_/X _60732_/Y _60754_/X _60755_/Y _84574_/D
+ sky130_fd_sc_hd__a41oi_4
X_48478_ _48478_/A _48478_/X sky130_fd_sc_hd__buf_2
X_79298_ _84796_/Q _84116_/Q _79298_/Y sky130_fd_sc_hd__nand2_4
X_69051_ _69478_/A _69051_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_217_0_CLK clkbuf_9_108_0_CLK/X _84501_/CLK sky130_fd_sc_hd__clkbuf_1
X_47429_ _47382_/A _47429_/X sky130_fd_sc_hd__buf_2
X_66263_ _84145_/Q _66264_/C sky130_fd_sc_hd__inv_2
X_78249_ _78248_/A _78248_/B _78250_/A sky130_fd_sc_hd__nand2_4
X_63475_ _63413_/A _63476_/C sky130_fd_sc_hd__buf_2
X_60687_ _60687_/A _60711_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_847_0_CLK clkbuf_9_423_0_CLK/X _86119_/CLK sky130_fd_sc_hd__clkbuf_1
X_68002_ _67999_/X _68001_/X _67977_/X _68002_/X sky130_fd_sc_hd__a21o_4
X_65214_ _65211_/X _85514_/Q _65212_/X _65213_/X _65214_/X sky130_fd_sc_hd__a211o_4
X_50440_ _50439_/X _50440_/B _50440_/Y sky130_fd_sc_hd__nand2_4
X_62426_ _62411_/X _62412_/X _62426_/C _62426_/Y sky130_fd_sc_hd__nor3_4
X_81260_ _81260_/CLK _81260_/D _76289_/A sky130_fd_sc_hd__dfxtp_4
X_66194_ _66191_/Y _66137_/X _66193_/Y _84150_/D sky130_fd_sc_hd__a21o_4
X_80211_ _80208_/X _80210_/Y _80211_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_9_338_0_CLK clkbuf_9_339_0_CLK/A clkbuf_9_338_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_65145_ _64944_/X _86124_/Q _65022_/X _65144_/X _65145_/X sky130_fd_sc_hd__a211o_4
X_50371_ _86214_/Q _50363_/X _50370_/Y _50371_/Y sky130_fd_sc_hd__o21ai_4
X_81191_ _81216_/CLK _81191_/D _49148_/A sky130_fd_sc_hd__dfxtp_4
X_62357_ _62501_/A _62386_/C sky130_fd_sc_hd__buf_2
X_52110_ _52106_/Y _52108_/X _52109_/X _85887_/D sky130_fd_sc_hd__a21oi_4
X_61308_ _61308_/A _72550_/A sky130_fd_sc_hd__buf_2
X_80142_ _57883_/Y _65605_/C _80141_/Y _80142_/X sky130_fd_sc_hd__o21a_4
X_53090_ _53107_/A _53069_/X _53107_/C _53090_/D _53090_/X sky130_fd_sc_hd__and4_4
X_65076_ _58785_/A _86031_/Q _65076_/X sky130_fd_sc_hd__and2_4
X_69953_ _69943_/X _69951_/Y _69938_/X _69952_/Y _69953_/X sky130_fd_sc_hd__a211o_4
X_62288_ _62288_/A _62288_/X sky130_fd_sc_hd__buf_2
X_52041_ _51928_/X _52041_/X sky130_fd_sc_hd__buf_2
X_68904_ _68900_/X _68903_/X _68878_/X _68904_/Y sky130_fd_sc_hd__a21oi_4
X_64027_ _64422_/C _64091_/B _64091_/C _64027_/D _64027_/Y sky130_fd_sc_hd__nand4_4
X_61239_ _75903_/A _60719_/X _61237_/Y _61238_/Y _84501_/D sky130_fd_sc_hd__o22a_4
X_84950_ _85407_/CLK _84950_/D _84950_/Q sky130_fd_sc_hd__dfxtp_4
X_80073_ _80073_/A _80073_/B _80073_/X sky130_fd_sc_hd__and2_4
X_69884_ _73372_/A _69833_/X _69617_/X _69883_/Y _69884_/X sky130_fd_sc_hd__a211o_4
X_83901_ _81975_/CLK _83901_/D _83901_/Q sky130_fd_sc_hd__dfxtp_4
X_68835_ _68831_/X _68834_/X _68737_/X _68835_/Y sky130_fd_sc_hd__a21oi_4
X_84881_ _84877_/CLK _58315_/X _84881_/Q sky130_fd_sc_hd__dfxtp_4
X_55800_ _55800_/A _55801_/D sky130_fd_sc_hd__buf_2
X_86620_ _85981_/CLK _47580_/Y _72188_/A sky130_fd_sc_hd__dfxtp_4
X_83832_ _83191_/CLK _70222_/X _83832_/Q sky130_fd_sc_hd__dfxtp_4
X_56780_ _56764_/B _56773_/Y _56774_/Y _56779_/Y _56780_/X sky130_fd_sc_hd__a211o_4
X_68766_ _68666_/X _68612_/X _68752_/Y _68765_/Y _68766_/X sky130_fd_sc_hd__a211o_4
X_53992_ _85527_/Q _53989_/X _53991_/Y _53992_/Y sky130_fd_sc_hd__o21ai_4
X_65978_ _65876_/X _85628_/Q _65976_/X _65977_/X _65978_/X sky130_fd_sc_hd__a211o_4
X_55731_ _85253_/Q _55244_/A _44043_/X _55730_/X _55731_/X sky130_fd_sc_hd__a211o_4
X_67717_ _68640_/A _67717_/X sky130_fd_sc_hd__buf_2
X_86551_ _86554_/CLK _48235_/Y _86551_/Q sky130_fd_sc_hd__dfxtp_4
X_64929_ _64929_/A _85845_/Q _64929_/X sky130_fd_sc_hd__and2_4
X_52943_ _52941_/Y _52920_/X _52942_/X _85726_/D sky130_fd_sc_hd__a21oi_4
X_83763_ _83763_/CLK _83763_/D _83763_/Q sky130_fd_sc_hd__dfxtp_4
X_80975_ _81059_/CLK _75693_/X _75082_/B sky130_fd_sc_hd__dfxtp_4
X_68697_ _69768_/A _68697_/X sky130_fd_sc_hd__buf_2
X_85502_ _85505_/CLK _54112_/Y _85502_/Q sky130_fd_sc_hd__dfxtp_4
X_58450_ _63244_/A _58452_/A sky130_fd_sc_hd__buf_2
X_82714_ _82715_/CLK _79028_/X _82670_/D sky130_fd_sc_hd__dfxtp_4
X_55662_ _55243_/A _55243_/B _55662_/Y sky130_fd_sc_hd__nand2_4
X_67648_ _86962_/Q _67551_/X _67552_/X _67647_/X _67649_/B sky130_fd_sc_hd__a211o_4
X_86482_ _86193_/CLK _48792_/Y _86482_/Q sky130_fd_sc_hd__dfxtp_4
X_52874_ _52821_/A _52874_/X sky130_fd_sc_hd__buf_2
X_83694_ _82381_/CLK _70815_/Y _83694_/Q sky130_fd_sc_hd__dfxtp_4
X_57401_ _57650_/A _57401_/B _57400_/X _57401_/Y sky130_fd_sc_hd__nor3_4
X_88221_ _87141_/CLK _41405_/Y _67860_/B sky130_fd_sc_hd__dfxtp_4
X_54613_ _54610_/Y _54611_/X _54612_/X _54613_/Y sky130_fd_sc_hd__a21oi_4
X_85433_ _85433_/CLK _54490_/Y _85433_/Q sky130_fd_sc_hd__dfxtp_4
X_51825_ _51821_/Y _51823_/X _51824_/X _51825_/Y sky130_fd_sc_hd__a21oi_4
X_58381_ _58366_/X _83352_/Q _58380_/Y _58381_/X sky130_fd_sc_hd__o21a_4
X_82645_ _82642_/CLK _83997_/Q _82645_/Q sky130_fd_sc_hd__dfxtp_4
X_55593_ _55592_/X _72643_/C sky130_fd_sc_hd__buf_2
X_67579_ _67675_/A _87721_/Q _67579_/X sky130_fd_sc_hd__and2_4
X_57332_ _56785_/B _56787_/X _56788_/A _57319_/D _45955_/X _57332_/Y
+ sky130_fd_sc_hd__a41oi_4
X_69318_ _69288_/A _69318_/B _69318_/X sky130_fd_sc_hd__and2_4
X_88152_ _88208_/CLK _88152_/D _67992_/B sky130_fd_sc_hd__dfxtp_4
X_54544_ _54538_/A _54526_/B _54538_/C _47093_/A _54544_/X sky130_fd_sc_hd__and4_4
X_85364_ _83630_/CLK _85364_/D _85364_/Q sky130_fd_sc_hd__dfxtp_4
X_51756_ _51768_/A _51749_/X _51755_/X _51756_/D _51756_/X sky130_fd_sc_hd__and4_4
X_70590_ _70959_/C _70591_/A sky130_fd_sc_hd__buf_2
X_82576_ _82702_/CLK _82576_/D _78193_/B sky130_fd_sc_hd__dfxtp_4
X_87103_ _87103_/CLK _44451_/Y _87103_/Q sky130_fd_sc_hd__dfxtp_4
X_84315_ _84314_/CLK _63544_/Y _80475_/B sky130_fd_sc_hd__dfxtp_4
X_50707_ _50596_/A _50738_/A sky130_fd_sc_hd__buf_2
X_57263_ _57261_/X _56643_/X _45617_/A _57236_/X _85043_/D sky130_fd_sc_hd__a2bb2o_4
X_81527_ _84079_/CLK _81539_/Q _81527_/Q sky130_fd_sc_hd__dfxtp_4
X_69249_ _69179_/A _87275_/Q _69249_/X sky130_fd_sc_hd__and2_4
X_88083_ _87826_/CLK _88083_/D _41980_/A sky130_fd_sc_hd__dfxtp_4
X_54475_ _54475_/A _54475_/X sky130_fd_sc_hd__buf_2
X_85295_ _83022_/CLK _56106_/Y _55826_/B sky130_fd_sc_hd__dfxtp_4
X_51687_ _85964_/Q _51675_/X _51686_/Y _51687_/Y sky130_fd_sc_hd__o21ai_4
X_59002_ _58904_/X _85761_/Q _58928_/X _59002_/X sky130_fd_sc_hd__o21a_4
X_56214_ _56214_/A _56205_/X _85273_/Q _56214_/Y sky130_fd_sc_hd__nand3_4
X_41440_ _41440_/A _41471_/B _41440_/X sky130_fd_sc_hd__or2_4
X_87034_ _86989_/CLK _87034_/D _87034_/Q sky130_fd_sc_hd__dfxtp_4
X_53426_ _53405_/X _53426_/B _53426_/Y sky130_fd_sc_hd__nand2_4
X_72260_ _72209_/X _85974_/Q _72259_/X _72260_/Y sky130_fd_sc_hd__o21ai_4
X_84246_ _82436_/CLK _64444_/X _84246_/Q sky130_fd_sc_hd__dfxtp_4
X_50638_ _50638_/A _50718_/A sky130_fd_sc_hd__buf_2
X_81458_ _83926_/CLK _76802_/B _81426_/D sky130_fd_sc_hd__dfxtp_4
X_57194_ _56698_/Y _57193_/Y _56671_/X _57182_/X _44239_/A _57195_/C
+ sky130_fd_sc_hd__a2111o_4
Xpsn_inst_psn_buff_2 _44267_/A _44279_/D sky130_fd_sc_hd__buf_2
X_71211_ _71211_/A _71232_/B _71219_/C _71211_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_opt_28_CLK _86500_/CLK _85865_/CLK sky130_fd_sc_hd__clkbuf_16
X_80409_ _80409_/A _80408_/Y _80409_/X sky130_fd_sc_hd__xor2_4
X_56145_ _56140_/A _56140_/B _56145_/C _56145_/Y sky130_fd_sc_hd__nand3_4
X_41371_ _41370_/Y _41371_/X sky130_fd_sc_hd__buf_2
X_53357_ _53357_/A _53371_/C sky130_fd_sc_hd__buf_2
X_72191_ _72179_/Y _72152_/X _72186_/X _72190_/X _83276_/D sky130_fd_sc_hd__a22oi_4
X_84177_ _84177_/CLK _84177_/D _84177_/Q sky130_fd_sc_hd__dfxtp_4
X_50569_ _50566_/Y _50551_/X _50568_/X _50569_/Y sky130_fd_sc_hd__a21oi_4
X_81389_ _81265_/CLK _83925_/Q _76895_/B sky130_fd_sc_hd__dfxtp_4
X_43110_ _43017_/A _43110_/X sky130_fd_sc_hd__buf_2
X_40322_ _46526_/A _48135_/A sky130_fd_sc_hd__buf_2
X_52308_ _64844_/B _52297_/X _52307_/Y _52308_/Y sky130_fd_sc_hd__o21ai_4
X_71142_ _48358_/X _71138_/X _71141_/Y _71142_/Y sky130_fd_sc_hd__o21ai_4
X_83128_ _83561_/CLK _83128_/D _83128_/Q sky130_fd_sc_hd__dfxtp_4
X_44090_ _44090_/A _44090_/B _44090_/Y sky130_fd_sc_hd__nand2_4
X_56076_ _56100_/A _56086_/B _55870_/B _56076_/Y sky130_fd_sc_hd__nand3_4
X_53288_ _53293_/A _53274_/B _53293_/C _52775_/D _53288_/X sky130_fd_sc_hd__and4_4
X_55027_ _55023_/Y _55024_/X _55026_/X _55027_/Y sky130_fd_sc_hd__a21oi_4
X_59904_ _60162_/A _59904_/B _60403_/A _59909_/A sky130_fd_sc_hd__and3_4
X_43041_ _87597_/Q _43041_/Y sky130_fd_sc_hd__inv_2
X_52239_ _52214_/A _52239_/X sky130_fd_sc_hd__buf_2
X_71073_ _71078_/A _71073_/B _71078_/C _71073_/Y sky130_fd_sc_hd__nand3_4
X_75950_ _75950_/A _81734_/D _75950_/X sky130_fd_sc_hd__xor2_4
X_83059_ _83572_/CLK _83059_/D _83059_/Q sky130_fd_sc_hd__dfxtp_4
X_87936_ _82888_/CLK _87936_/D _87936_/Q sky130_fd_sc_hd__dfxtp_4
X_74901_ _81129_/D _74891_/B _74900_/Y _74901_/X sky130_fd_sc_hd__o21a_4
X_70024_ _70011_/X _68647_/Y _70012_/X _70023_/Y _70024_/X sky130_fd_sc_hd__a211o_4
X_59835_ _59829_/X _59830_/Y _59834_/X _59835_/X sky130_fd_sc_hd__o21a_4
X_75881_ _75714_/Y _80786_/D sky130_fd_sc_hd__inv_2
X_87867_ _87086_/CLK _42432_/Y _87867_/Q sky130_fd_sc_hd__dfxtp_4
X_46800_ _82958_/Q _46800_/Y sky130_fd_sc_hd__inv_2
X_77620_ _77664_/C _77666_/A _77621_/A sky130_fd_sc_hd__and2_4
X_74832_ _74844_/A _46115_/A _74832_/Y sky130_fd_sc_hd__nand2_4
X_86818_ _86814_/CLK _46006_/Y _86818_/Q sky130_fd_sc_hd__dfxtp_4
X_47780_ _47780_/A _53240_/B sky130_fd_sc_hd__buf_2
X_59766_ _59664_/A _59766_/X sky130_fd_sc_hd__buf_2
X_56978_ _56975_/Y _56977_/Y _45909_/A _56978_/Y sky130_fd_sc_hd__o21ai_4
X_44992_ _64275_/B _61386_/B sky130_fd_sc_hd__buf_2
X_87798_ _87285_/CLK _42621_/Y _73484_/A sky130_fd_sc_hd__dfxtp_4
X_58717_ _58714_/X _85781_/Q _58716_/X _58717_/X sky130_fd_sc_hd__o21a_4
X_46731_ _83677_/Q _54332_/B sky130_fd_sc_hd__inv_2
X_77551_ _77551_/A _82116_/Q _77552_/A sky130_fd_sc_hd__nand2_4
X_43943_ _80667_/Q _43944_/A sky130_fd_sc_hd__buf_2
X_74763_ _71735_/A _70630_/B _74763_/C _71010_/X _74763_/X sky130_fd_sc_hd__and4_4
X_55929_ _55947_/A _56303_/C _55929_/X sky130_fd_sc_hd__and2_4
X_86749_ _86749_/CLK _86749_/D _86749_/Q sky130_fd_sc_hd__dfxtp_4
X_71975_ _71973_/Y _71969_/X _71974_/Y _71975_/Y sky130_fd_sc_hd__a21boi_4
X_59697_ _59680_/Y _59688_/X _59689_/Y _59695_/Y _59696_/Y _59697_/Y
+ sky130_fd_sc_hd__a41oi_4
X_76502_ _76503_/A _81542_/Q _76502_/Y sky130_fd_sc_hd__nor2_4
X_49450_ _86385_/Q _49443_/X _49449_/Y _49450_/Y sky130_fd_sc_hd__o21ai_4
X_73714_ _73641_/A _65997_/B _73714_/X sky130_fd_sc_hd__and2_4
X_46662_ _46662_/A _46662_/X sky130_fd_sc_hd__buf_2
X_70926_ _70873_/A _70863_/C _70925_/X _70919_/D _70926_/Y sky130_fd_sc_hd__nand4_4
X_58648_ _58659_/A _86395_/Q _58648_/Y sky130_fd_sc_hd__nor2_4
X_77482_ _77465_/B _77458_/X _77482_/Y sky130_fd_sc_hd__nand2_4
X_43874_ _41268_/X _43868_/X _69045_/B _43870_/X _43874_/X sky130_fd_sc_hd__a2bb2o_4
X_74694_ _74694_/A _74694_/B _74694_/Y sky130_fd_sc_hd__nand2_4
X_48401_ _48401_/A _48401_/B _48401_/Y sky130_fd_sc_hd__nand2_4
X_79221_ _79220_/Y _79221_/Y sky130_fd_sc_hd__inv_2
X_45613_ _85107_/Q _45793_/B _45613_/Y sky130_fd_sc_hd__nor2_4
X_76433_ _76425_/X _76432_/X _76433_/X sky130_fd_sc_hd__xor2_4
X_42825_ _41461_/X _42821_/X _66535_/B _42822_/X _42825_/X sky130_fd_sc_hd__a2bb2o_4
X_49381_ _49377_/Y _49378_/X _49380_/X _86398_/D sky130_fd_sc_hd__a21oi_4
X_73645_ _73646_/B _73635_/X _73644_/X _73645_/X sky130_fd_sc_hd__a21o_4
X_46593_ _46588_/Y _46576_/X _46592_/Y _46593_/Y sky130_fd_sc_hd__a21boi_4
X_70857_ _71068_/B _71072_/A sky130_fd_sc_hd__buf_2
X_58579_ _58100_/X _85952_/Q _58568_/X _58579_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_7_53_0_CLK clkbuf_6_26_0_CLK/X clkbuf_7_53_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_60610_ _60610_/A _60513_/B _79127_/A _60610_/X sky130_fd_sc_hd__or3_4
X_48332_ _48897_/A _48548_/A sky130_fd_sc_hd__buf_2
X_79152_ _79152_/A _79152_/B _79152_/X sky130_fd_sc_hd__xor2_4
X_45544_ _63110_/B _61440_/A sky130_fd_sc_hd__buf_2
X_76364_ _76344_/Y _76348_/B _76347_/A _76364_/X sky130_fd_sc_hd__o21a_4
X_42756_ _41268_/X _42745_/X _69042_/B _42746_/X _42756_/X sky130_fd_sc_hd__a2bb2o_4
X_61590_ _61558_/A _61590_/B _61590_/C _61590_/Y sky130_fd_sc_hd__nand3_4
X_73576_ _68380_/Y _73319_/X _73551_/X _73575_/Y _73576_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_8_193_0_CLK clkbuf_7_96_0_CLK/X clkbuf_9_387_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_70788_ _52863_/B _70761_/A _70787_/Y _70788_/Y sky130_fd_sc_hd__o21ai_4
X_78103_ _82565_/Q _78103_/B _78103_/Y sky130_fd_sc_hd__nor2_4
X_75315_ _80691_/Q _80991_/Q _75315_/Y sky130_fd_sc_hd__nand2_4
X_41707_ _41707_/A _88165_/D sky130_fd_sc_hd__inv_2
X_48263_ _48478_/A _48263_/X sky130_fd_sc_hd__buf_2
X_60541_ _63301_/C _60541_/B _60541_/C _60541_/Y sky130_fd_sc_hd__nor3_4
X_72527_ _72527_/A _72527_/B _79493_/B _72527_/Y sky130_fd_sc_hd__nand3_4
X_79083_ _79080_/A _82751_/Q _79083_/Y sky130_fd_sc_hd__nand2_4
X_45475_ _44932_/A _45490_/B sky130_fd_sc_hd__buf_2
X_76295_ _76272_/Y _76293_/Y _76294_/Y _76295_/Y sky130_fd_sc_hd__a21oi_4
X_42687_ _42590_/A _42687_/X sky130_fd_sc_hd__buf_2
X_47214_ _47196_/A _52918_/B _47214_/Y sky130_fd_sc_hd__nand2_4
X_78034_ _82177_/Q _78034_/Y sky130_fd_sc_hd__inv_2
X_44426_ _40362_/X _44548_/A sky130_fd_sc_hd__buf_2
X_63260_ _58396_/Y _63259_/X _63234_/X _58274_/A _63235_/X _63260_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75246_ _75230_/B _75228_/X _75223_/Y _75246_/Y sky130_fd_sc_hd__a21boi_4
X_41638_ _41799_/A _41638_/X sky130_fd_sc_hd__buf_2
X_72458_ _72361_/X _85668_/Q _72362_/X _72458_/X sky130_fd_sc_hd__o21a_4
X_48194_ _48193_/X _48194_/X sky130_fd_sc_hd__buf_2
X_60472_ _60472_/A _60606_/A _60430_/Y _60443_/A _60493_/A sky130_fd_sc_hd__nand4_4
Xclkbuf_7_68_0_CLK clkbuf_7_69_0_CLK/A clkbuf_7_68_0_CLK/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_opt_19_CLK _85557_/CLK _83297_/CLK sky130_fd_sc_hd__clkbuf_16
X_62211_ _61301_/X _62560_/B _62560_/C _62211_/D _62211_/Y sky130_fd_sc_hd__nand4_4
X_47145_ _47004_/A _47145_/X sky130_fd_sc_hd__buf_2
X_71409_ _70682_/A _71411_/B _71411_/C _71409_/Y sky130_fd_sc_hd__nor3_4
X_44357_ _41721_/X _44345_/X _87150_/Q _44346_/X _44357_/X sky130_fd_sc_hd__a2bb2o_4
X_63191_ _58377_/A _63190_/X _63175_/X _58251_/A _63176_/X _63191_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75177_ _75178_/A _75178_/B _75178_/C _75180_/A sky130_fd_sc_hd__a21oi_4
X_41569_ _41548_/X _82316_/Q _41568_/X _41569_/Y sky130_fd_sc_hd__o21ai_4
X_72389_ _72123_/A _72389_/X sky130_fd_sc_hd__buf_2
X_43308_ _43212_/A _43308_/X sky130_fd_sc_hd__buf_2
X_62142_ _62142_/A _62138_/Y _62139_/Y _62141_/Y _62142_/Y sky130_fd_sc_hd__nand4_4
X_74128_ _74080_/X _86217_/Q _74103_/X _74127_/X _74128_/X sky130_fd_sc_hd__a211o_4
X_47076_ _47072_/Y _47035_/X _47075_/X _86673_/D sky130_fd_sc_hd__a21oi_4
X_44288_ _44287_/X _44288_/X sky130_fd_sc_hd__buf_2
X_79985_ _79985_/A _79985_/B _79985_/Y sky130_fd_sc_hd__xnor2_4
X_46027_ _41460_/Y _46022_/X _66544_/B _46023_/X _46027_/X sky130_fd_sc_hd__a2bb2o_4
X_43239_ _41028_/X _43216_/X _87523_/Q _43218_/X _87523_/D sky130_fd_sc_hd__a2bb2o_4
X_74059_ _74012_/X _86220_/Q _73948_/X _74058_/X _74059_/X sky130_fd_sc_hd__a211o_4
X_66950_ _66902_/X _86822_/Q _66950_/X sky130_fd_sc_hd__and2_4
X_62073_ _61593_/B _62007_/X _62149_/C _62008_/X _62077_/B sky130_fd_sc_hd__nand4_4
X_78936_ _78921_/A _82511_/D _78935_/X _78937_/B sky130_fd_sc_hd__o21ai_4
Xclkbuf_8_131_0_CLK clkbuf_7_65_0_CLK/X clkbuf_9_262_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_65901_ _65916_/A _65916_/B _65901_/C _65901_/X sky130_fd_sc_hd__and3_4
X_61024_ _60937_/B _61024_/B _61024_/Y sky130_fd_sc_hd__nand2_4
X_66881_ _87430_/Q _66878_/X _66879_/X _66880_/X _66881_/X sky130_fd_sc_hd__a211o_4
X_78867_ _78865_/X _78867_/B _78867_/Y sky130_fd_sc_hd__nor2_4
X_68620_ _68616_/X _68619_/X _68470_/X _68620_/X sky130_fd_sc_hd__a21o_4
X_65832_ _65829_/Y _65830_/X _65831_/X _65832_/X sky130_fd_sc_hd__a21o_4
X_77818_ _77807_/Y _77818_/Y sky130_fd_sc_hd__inv_2
X_47978_ _47978_/A _50302_/B sky130_fd_sc_hd__buf_2
X_78798_ _78798_/A _78799_/B sky130_fd_sc_hd__inv_2
X_49717_ _49716_/X _52931_/B _49717_/Y sky130_fd_sc_hd__nand2_4
X_68551_ _68548_/X _68551_/B _68551_/Y sky130_fd_sc_hd__nand2_4
X_46929_ _54446_/B _52752_/B sky130_fd_sc_hd__buf_2
Xclkbuf_8_146_0_CLK clkbuf_7_73_0_CLK/X clkbuf_8_146_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_65763_ _65763_/A _85867_/Q _65763_/X sky130_fd_sc_hd__and2_4
X_77749_ _82052_/Q _77751_/B sky130_fd_sc_hd__inv_2
X_62975_ _62967_/A _63335_/A _62939_/X _62975_/D _62975_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_141_0_CLK clkbuf_9_70_0_CLK/X _81259_/CLK sky130_fd_sc_hd__clkbuf_1
X_67502_ _67025_/X _67502_/X sky130_fd_sc_hd__buf_2
X_64714_ _64752_/A _64714_/X sky130_fd_sc_hd__buf_2
X_49648_ _49638_/A _52863_/B _49648_/Y sky130_fd_sc_hd__nand2_4
X_61926_ _61915_/X _61918_/X _61925_/Y _84741_/Q _61895_/X _61926_/Y
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_10_771_0_CLK clkbuf_9_385_0_CLK/X _82532_/CLK sky130_fd_sc_hd__clkbuf_1
X_80760_ _80792_/CLK _80760_/D _81136_/D sky130_fd_sc_hd__dfxtp_4
X_68482_ _68452_/A _87247_/Q _68482_/X sky130_fd_sc_hd__and2_4
X_65694_ _65694_/A _65694_/B _65694_/Y sky130_fd_sc_hd__nand2_4
X_67433_ _67312_/X _67433_/X sky130_fd_sc_hd__buf_2
X_79419_ _79419_/A _79419_/B _79419_/X sky130_fd_sc_hd__or2_4
X_64645_ _64641_/X _64644_/X _64619_/X _64649_/A sky130_fd_sc_hd__a21o_4
Xclkbuf_9_262_0_CLK clkbuf_9_262_0_CLK/A clkbuf_9_262_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_49579_ _49496_/A _49579_/X sky130_fd_sc_hd__buf_2
X_80691_ _80676_/CLK _80691_/D _80691_/Q sky130_fd_sc_hd__dfxtp_4
X_61857_ _61428_/X _61874_/B _61809_/C _61874_/D _61857_/Y sky130_fd_sc_hd__nand4_4
X_51610_ _51606_/Y _51585_/X _51609_/X _51610_/Y sky130_fd_sc_hd__a21oi_4
X_82430_ _84119_/CLK _82462_/Q _78729_/A sky130_fd_sc_hd__dfxtp_4
X_60808_ _60805_/Y _60743_/X _60696_/Y _60781_/Y _60807_/Y _84562_/D
+ sky130_fd_sc_hd__a41oi_4
X_67364_ _67126_/X _67364_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_156_0_CLK clkbuf_9_78_0_CLK/X _81279_/CLK sky130_fd_sc_hd__clkbuf_1
X_52590_ _52590_/A _52590_/B _52590_/Y sky130_fd_sc_hd__nand2_4
X_64576_ _58124_/A _64797_/A sky130_fd_sc_hd__buf_2
X_61788_ _61787_/X _61788_/X sky130_fd_sc_hd__buf_2
X_69103_ _69611_/A _69103_/X sky130_fd_sc_hd__buf_2
XPHY_709 sky130_fd_sc_hd__decap_3
X_66315_ _66312_/X _66314_/X _66315_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_786_0_CLK clkbuf_9_393_0_CLK/X _82624_/CLK sky130_fd_sc_hd__clkbuf_1
X_51541_ _51545_/A _53067_/B _51541_/Y sky130_fd_sc_hd__nand2_4
X_63527_ _63495_/X _63520_/X _63521_/X _63525_/X _63526_/Y _63527_/Y
+ sky130_fd_sc_hd__o41ai_4
X_82361_ _84981_/CLK _77220_/X _47926_/A sky130_fd_sc_hd__dfxtp_4
X_60739_ _60738_/Y _60739_/X sky130_fd_sc_hd__buf_2
X_67295_ _87925_/Q _67293_/X _67271_/X _67294_/X _67295_/X sky130_fd_sc_hd__a211o_4
X_84100_ _84105_/CLK _66709_/X _84100_/Q sky130_fd_sc_hd__dfxtp_4
X_81312_ _81801_/CLK _77000_/X _81280_/D sky130_fd_sc_hd__dfxtp_4
X_69034_ _87480_/Q _68989_/X _69010_/X _69033_/X _69034_/X sky130_fd_sc_hd__a211o_4
X_54260_ _54258_/Y _54253_/X _54259_/X _85475_/D sky130_fd_sc_hd__a21oi_4
X_66246_ _66179_/X _66244_/Y _66245_/Y _66246_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_277_0_CLK clkbuf_9_277_0_CLK/A clkbuf_9_277_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_85080_ _85083_/CLK _85080_/D _85080_/Q sky130_fd_sc_hd__dfxtp_4
X_51472_ _51552_/A _51494_/C sky130_fd_sc_hd__buf_2
X_63458_ _63458_/A _63458_/X sky130_fd_sc_hd__buf_2
X_82292_ _82103_/CLK _81916_/Q _40829_/B sky130_fd_sc_hd__dfxtp_4
X_53211_ _53211_/A _53211_/B _53195_/X _53211_/D _53211_/X sky130_fd_sc_hd__and4_4
X_84031_ _81154_/CLK _68132_/X _82071_/D sky130_fd_sc_hd__dfxtp_4
X_50423_ _50432_/A _52128_/B _50423_/Y sky130_fd_sc_hd__nand2_4
X_62409_ _61489_/B _62390_/X _62363_/X _62407_/X _62408_/X _62409_/X
+ sky130_fd_sc_hd__a41o_4
X_81243_ _85338_/CLK _81051_/Q _47585_/A sky130_fd_sc_hd__dfxtp_4
X_54191_ _54191_/A _54191_/B _54191_/C _53023_/D _54191_/X sky130_fd_sc_hd__and4_4
X_66177_ _66177_/A _66164_/B _66177_/C _66177_/Y sky130_fd_sc_hd__nor3_4
X_63389_ _63389_/A _63389_/B _63418_/C _63389_/D _63389_/Y sky130_fd_sc_hd__nand4_4
X_53142_ _85689_/Q _53120_/X _53141_/Y _53142_/Y sky130_fd_sc_hd__o21ai_4
X_65128_ _64584_/X _65791_/A sky130_fd_sc_hd__buf_2
X_50354_ _50317_/X _48310_/B _50354_/Y sky130_fd_sc_hd__nand2_4
X_81174_ _83974_/CLK _74993_/B _40430_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_200_0_CLK clkbuf_9_201_0_CLK/A clkbuf_9_200_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
Xpsn_inst_psn_buff_20 _43018_/Y _53441_/A sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_31 _47002_/A _40372_/B1 sky130_fd_sc_hd__buf_2
X_80125_ _80125_/A _80124_/X _80125_/Y sky130_fd_sc_hd__xnor2_4
X_53073_ _85702_/Q _53065_/X _53072_/Y _53073_/Y sky130_fd_sc_hd__o21ai_4
X_57950_ _57926_/X _86001_/Q _57949_/X _57950_/Y sky130_fd_sc_hd__o21ai_4
X_65059_ _64828_/A _65059_/X sky130_fd_sc_hd__buf_2
X_69936_ _87043_/Q _44225_/B _57800_/A _69935_/X _69937_/B sky130_fd_sc_hd__a211o_4
X_50285_ _50285_/A _48231_/B _50285_/Y sky130_fd_sc_hd__nand2_4
X_85982_ _85692_/CLK _51593_/Y _85982_/Q sky130_fd_sc_hd__dfxtp_4
X_52024_ _52431_/A _52058_/A sky130_fd_sc_hd__buf_2
X_56901_ _56900_/X _56901_/Y sky130_fd_sc_hd__inv_2
X_87721_ _87210_/CLK _87721_/D _87721_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_724_0_CLK clkbuf_9_362_0_CLK/X _82301_/CLK sky130_fd_sc_hd__clkbuf_1
X_84933_ _85379_/CLK _84933_/D _84933_/Q sky130_fd_sc_hd__dfxtp_4
X_80056_ _80073_/B _80056_/B _80056_/X sky130_fd_sc_hd__xor2_4
X_57881_ _57877_/Y _57880_/Y _57829_/X _57881_/X sky130_fd_sc_hd__a21o_4
X_69867_ _69864_/X _69866_/X _69742_/X _69867_/Y sky130_fd_sc_hd__a21oi_4
X_59620_ _60122_/A _60122_/C _59640_/A sky130_fd_sc_hd__and2_4
X_56832_ _56831_/X _56832_/X sky130_fd_sc_hd__buf_2
X_68818_ _69182_/A _68818_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_215_0_CLK clkbuf_9_214_0_CLK/A clkbuf_9_215_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_87652_ _87652_/CLK _87652_/D _67691_/B sky130_fd_sc_hd__dfxtp_4
X_84864_ _84344_/CLK _58381_/X _84864_/Q sky130_fd_sc_hd__dfxtp_4
X_69798_ _69770_/A _88322_/Q _69798_/X sky130_fd_sc_hd__and2_4
X_86603_ _85962_/CLK _47740_/Y _72384_/A sky130_fd_sc_hd__dfxtp_4
X_83815_ _83842_/CLK _83815_/D _83815_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_109_0_CLK clkbuf_9_54_0_CLK/X _84549_/CLK sky130_fd_sc_hd__clkbuf_1
X_59551_ _59551_/A _60407_/C sky130_fd_sc_hd__buf_2
X_56763_ _56740_/X _56756_/X _56758_/X _56761_/X _57003_/B _56764_/D
+ sky130_fd_sc_hd__a41o_4
X_68749_ _68744_/X _68747_/X _68748_/X _68749_/X sky130_fd_sc_hd__a21o_4
X_87583_ _88111_/CLK _43082_/Y _74033_/A sky130_fd_sc_hd__dfxtp_4
X_53975_ _53972_/Y _53948_/X _53974_/Y _85531_/D sky130_fd_sc_hd__a21boi_4
X_84795_ _86713_/CLK _84795_/D _84795_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_739_0_CLK clkbuf_9_369_0_CLK/X _87225_/CLK sky130_fd_sc_hd__clkbuf_1
X_58502_ _63459_/B _58502_/B _58502_/Y sky130_fd_sc_hd__nor2_4
X_55714_ _56270_/C _55244_/A _44043_/X _55713_/X _55714_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_4_0_0_CLK clkbuf_3_0_1_CLK/X clkbuf_4_0_1_CLK/A sky130_fd_sc_hd__clkbuf_1
X_86534_ _86534_/CLK _86534_/D _66301_/B sky130_fd_sc_hd__dfxtp_4
X_40940_ _40717_/X _40941_/A sky130_fd_sc_hd__buf_2
X_52926_ _52845_/A _52926_/X sky130_fd_sc_hd__buf_2
X_71760_ _70500_/D _70760_/B _71761_/A sky130_fd_sc_hd__nor2_4
X_59482_ _63369_/B _58532_/X _59482_/Y sky130_fd_sc_hd__nor2_4
X_83746_ _83749_/CLK _83746_/D _83746_/Q sky130_fd_sc_hd__dfxtp_4
X_56694_ _56694_/A _56664_/Y _56694_/C _56694_/Y sky130_fd_sc_hd__nand3_4
X_80958_ _83967_/CLK _80958_/D _80958_/Q sky130_fd_sc_hd__dfxtp_4
X_70711_ _52752_/B _70699_/X _70710_/Y _70711_/Y sky130_fd_sc_hd__o21ai_4
X_58433_ _63198_/A _58434_/A sky130_fd_sc_hd__buf_2
X_55645_ _55447_/Y _55451_/B _55491_/X _56650_/B sky130_fd_sc_hd__a21boi_4
X_86465_ _83311_/CLK _86465_/D _86465_/Q sky130_fd_sc_hd__dfxtp_4
X_40871_ _40836_/A _40871_/X sky130_fd_sc_hd__buf_2
X_52857_ _52853_/A _52853_/B _52853_/C _52857_/D _52857_/X sky130_fd_sc_hd__and4_4
X_71691_ _71690_/Y _71691_/Y sky130_fd_sc_hd__inv_2
X_83677_ _83681_/CLK _70872_/Y _83677_/Q sky130_fd_sc_hd__dfxtp_4
X_80889_ _80818_/CLK _80889_/D _80889_/Q sky130_fd_sc_hd__dfxtp_4
X_88204_ _87436_/CLK _41500_/Y _66752_/B sky130_fd_sc_hd__dfxtp_4
X_42610_ _42610_/A _49210_/B sky130_fd_sc_hd__buf_2
X_73430_ _73359_/X _83055_/Q _73406_/X _73429_/X _73430_/X sky130_fd_sc_hd__a211o_4
X_85416_ _85643_/CLK _54581_/Y _85416_/Q sky130_fd_sc_hd__dfxtp_4
X_51808_ _85942_/Q _51789_/X _51807_/Y _51808_/Y sky130_fd_sc_hd__o21ai_4
X_70642_ _70925_/A _70642_/X sky130_fd_sc_hd__buf_2
X_58364_ _58364_/A _58364_/B _58364_/Y sky130_fd_sc_hd__nand2_4
X_82628_ _87684_/CLK _82628_/D _82628_/Q sky130_fd_sc_hd__dfxtp_4
X_43590_ _47872_/A _43013_/X _47832_/A _43591_/A sky130_fd_sc_hd__a21oi_4
X_55576_ _85052_/Q _55571_/X _55513_/X _55575_/Y _55576_/X sky130_fd_sc_hd__a211o_4
X_86396_ _86398_/CLK _86396_/D _58633_/B sky130_fd_sc_hd__dfxtp_4
X_52788_ _85754_/Q _52765_/X _52787_/Y _52788_/Y sky130_fd_sc_hd__o21ai_4
X_57315_ _57315_/A _57315_/Y sky130_fd_sc_hd__inv_2
X_88135_ _88133_/CLK _88135_/D _88135_/Q sky130_fd_sc_hd__dfxtp_4
X_42541_ _42521_/X _42522_/X _40762_/X _69110_/A _42540_/X _42542_/A
+ sky130_fd_sc_hd__o32ai_4
X_54527_ _54525_/Y _54502_/X _54526_/X _54527_/Y sky130_fd_sc_hd__a21oi_4
X_73361_ _73359_/X _83058_/Q _73238_/X _73360_/X _73361_/X sky130_fd_sc_hd__a211o_4
X_85347_ _85346_/CLK _85347_/D _85347_/Q sky130_fd_sc_hd__dfxtp_4
X_51739_ _46616_/A _54400_/A sky130_fd_sc_hd__buf_2
X_70573_ _71867_/A _70573_/B _70568_/C _70568_/D _70573_/Y sky130_fd_sc_hd__nor4_4
X_82559_ _82557_/CLK _82559_/D _82559_/Q sky130_fd_sc_hd__dfxtp_4
X_58295_ _64525_/C _58296_/A sky130_fd_sc_hd__buf_2
X_75100_ _75100_/A _75100_/Y sky130_fd_sc_hd__inv_2
X_72312_ _83266_/Q _72250_/X _72304_/X _72311_/X _72312_/Y sky130_fd_sc_hd__a2bb2oi_4
X_45260_ _62544_/A _61607_/B sky130_fd_sc_hd__buf_2
X_57246_ _57243_/X _56589_/X _85052_/Q _57245_/X _85052_/D sky130_fd_sc_hd__a2bb2o_4
X_76080_ _76071_/Y _76078_/Y _76079_/Y _76080_/X sky130_fd_sc_hd__o21a_4
X_88066_ _87553_/CLK _42027_/Y _73196_/A sky130_fd_sc_hd__dfxtp_4
X_42472_ _41993_/A _42472_/X sky130_fd_sc_hd__buf_2
X_54458_ _54321_/A _54486_/A sky130_fd_sc_hd__buf_2
X_73292_ _73277_/X _73281_/Y _73291_/X _73292_/X sky130_fd_sc_hd__a21o_4
X_85278_ _85248_/CLK _85278_/D _85278_/Q sky130_fd_sc_hd__dfxtp_4
X_44211_ _45950_/A _44204_/Y _44210_/X _44211_/Y sky130_fd_sc_hd__nor3_4
X_75031_ _75047_/B _75031_/Y sky130_fd_sc_hd__inv_2
X_41423_ _41421_/X _82888_/Q _41422_/X _41423_/X sky130_fd_sc_hd__o21a_4
X_87017_ _87011_/CLK _87017_/D _87017_/Q sky130_fd_sc_hd__dfxtp_4
X_53409_ _53357_/A _53410_/C sky130_fd_sc_hd__buf_2
X_72243_ _72228_/X _85975_/Q _72242_/X _72243_/Y sky130_fd_sc_hd__o21ai_4
X_84229_ _85315_/CLK _84229_/D _79836_/A sky130_fd_sc_hd__dfxtp_4
X_45191_ _85198_/Q _45176_/X _45190_/X _45191_/Y sky130_fd_sc_hd__o21ai_4
X_57177_ _56801_/X _56738_/X _56821_/X _57156_/X _45957_/A _57177_/Y
+ sky130_fd_sc_hd__a41oi_4
X_54389_ _85451_/Q _54376_/X _54388_/Y _54389_/Y sky130_fd_sc_hd__o21ai_4
X_56128_ _56117_/B _56143_/B _55773_/D _55801_/B _56128_/Y sky130_fd_sc_hd__nand4_4
X_44142_ _44004_/Y _44142_/X sky130_fd_sc_hd__buf_2
X_41354_ _41159_/A _82900_/Q _41354_/X sky130_fd_sc_hd__or2_4
X_72174_ _72220_/A _72174_/B _72174_/Y sky130_fd_sc_hd__nor2_4
X_71125_ _71112_/X _71080_/B _71119_/C _71125_/Y sky130_fd_sc_hd__nand3_4
X_48950_ _48908_/A _71989_/B _48950_/X sky130_fd_sc_hd__and2_4
X_44073_ _86755_/Q _55129_/A sky130_fd_sc_hd__inv_2
X_56059_ _74310_/C _55928_/A _56059_/Y sky130_fd_sc_hd__xnor2_4
X_79770_ _79767_/Y _79750_/Y _79769_/X _79770_/Y sky130_fd_sc_hd__o21ai_4
X_41285_ _41282_/X _41283_/X _69129_/B _41284_/X _88244_/D sky130_fd_sc_hd__a2bb2o_4
X_76982_ _84534_/Q _62498_/C _76982_/X sky130_fd_sc_hd__xor2_4
X_47901_ _47912_/A _50264_/B _47901_/Y sky130_fd_sc_hd__nand2_4
X_43024_ _43024_/A _43127_/A sky130_fd_sc_hd__buf_2
X_78721_ _78721_/A _78721_/B _78725_/A sky130_fd_sc_hd__nand2_4
X_71056_ _48901_/B _71047_/X _71055_/Y _71056_/Y sky130_fd_sc_hd__o21ai_4
X_75933_ _75933_/A _75933_/B _75933_/Y sky130_fd_sc_hd__nor2_4
X_87919_ _87473_/CLK _87919_/D _87919_/Q sky130_fd_sc_hd__dfxtp_4
X_48881_ _48471_/A _48881_/X sky130_fd_sc_hd__buf_2
X_70007_ _69520_/X _69668_/Y _69984_/X _70006_/Y _70007_/X sky130_fd_sc_hd__a211o_4
X_47832_ _47832_/A _47832_/X sky130_fd_sc_hd__buf_2
X_59818_ _80433_/A _59339_/X _59688_/X _59817_/Y _84695_/D sky130_fd_sc_hd__a2bb2oi_4
X_78652_ _78651_/X _78652_/Y sky130_fd_sc_hd__inv_2
X_75864_ _75864_/A _81024_/Q _75862_/Y _75865_/A sky130_fd_sc_hd__nand3_4
X_77603_ _77603_/A _77600_/Y _77603_/C _77603_/X sky130_fd_sc_hd__or3_4
X_74815_ _46227_/A _80667_/D sky130_fd_sc_hd__inv_2
X_47763_ _47762_/Y _53232_/B sky130_fd_sc_hd__buf_2
X_59749_ _59629_/A _59755_/A sky130_fd_sc_hd__buf_2
X_78583_ _78569_/A _78569_/B _78568_/A _78591_/A sky130_fd_sc_hd__o21a_4
X_44975_ _44975_/A _44975_/X sky130_fd_sc_hd__buf_2
X_75795_ _80923_/Q _75802_/B sky130_fd_sc_hd__inv_2
X_49502_ _49502_/A _51026_/B _49502_/Y sky130_fd_sc_hd__nand2_4
X_46714_ _46667_/A _46717_/C sky130_fd_sc_hd__buf_2
X_77534_ _77533_/Y _77537_/B sky130_fd_sc_hd__inv_2
X_43926_ _43926_/A _87196_/D sky130_fd_sc_hd__inv_2
X_62760_ _62711_/A _84832_/Q _62737_/X _62738_/D _62760_/X sky130_fd_sc_hd__and4_4
X_74746_ _70730_/X _74797_/C sky130_fd_sc_hd__buf_2
X_71958_ _83313_/Q _57615_/X _71957_/Y _71958_/Y sky130_fd_sc_hd__o21ai_4
X_47694_ _47694_/A _54885_/B sky130_fd_sc_hd__inv_2
X_49433_ _49569_/A _49434_/A sky130_fd_sc_hd__buf_2
X_61711_ _59635_/Y _61711_/X sky130_fd_sc_hd__buf_2
X_70909_ _70909_/A _70909_/X sky130_fd_sc_hd__buf_2
X_46645_ _82974_/Q _54286_/D sky130_fd_sc_hd__inv_2
X_77465_ _77458_/X _77465_/B _82194_/D sky130_fd_sc_hd__xor2_4
X_43857_ _43846_/X _43854_/X _41220_/X _87231_/Q _43847_/X _43858_/A
+ sky130_fd_sc_hd__o32ai_4
X_62691_ _58228_/X _62689_/X _60205_/X _60263_/C _62690_/X _62691_/Y
+ sky130_fd_sc_hd__a41oi_4
X_74677_ _74675_/X _56798_/A _74676_/Y _74678_/A sky130_fd_sc_hd__o21ai_4
X_71889_ _71867_/A _71783_/A _71783_/C _71319_/B _71889_/Y sky130_fd_sc_hd__nor4_4
X_79204_ _79201_/Y _79202_/Y _79203_/A _79205_/C sky130_fd_sc_hd__a21o_4
X_64430_ _64267_/A _64511_/B sky130_fd_sc_hd__buf_2
X_76416_ _76412_/X _76417_/C _76415_/Y _76418_/A sky130_fd_sc_hd__a21o_4
X_42808_ _42795_/X _42796_/X _41408_/X _67889_/B _42805_/X _42808_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49364_ _49374_/A _49364_/B _49380_/C _52580_/D _49364_/X sky130_fd_sc_hd__and4_4
X_61642_ _61642_/A _61642_/Y sky130_fd_sc_hd__inv_2
X_73628_ _44189_/X _73701_/B sky130_fd_sc_hd__buf_2
X_46576_ _46399_/A _46576_/X sky130_fd_sc_hd__buf_2
X_77396_ _77396_/A _77396_/B _77396_/Y sky130_fd_sc_hd__nor2_4
X_43788_ _41028_/X _43770_/X _69358_/B _43772_/X _43788_/X sky130_fd_sc_hd__a2bb2o_4
X_48315_ _48264_/X _50358_/B _48315_/Y sky130_fd_sc_hd__nand2_4
X_79135_ _79135_/A _79135_/B _79135_/X sky130_fd_sc_hd__xor2_4
X_45527_ _45527_/A _45381_/B _45527_/Y sky130_fd_sc_hd__nand2_4
X_64361_ _64361_/A _64363_/A sky130_fd_sc_hd__buf_2
X_76347_ _76347_/A _76348_/C sky130_fd_sc_hd__inv_2
X_42739_ _42720_/X _42739_/X sky130_fd_sc_hd__buf_2
X_49295_ _49287_/A _51324_/B _49295_/Y sky130_fd_sc_hd__nand2_4
X_73559_ _73556_/X _73558_/Y _73559_/Y sky130_fd_sc_hd__nand2_4
X_61573_ _58452_/A _61563_/B _61563_/C _61563_/D _61574_/A sky130_fd_sc_hd__nand4_4
X_66100_ _64898_/A _66226_/A sky130_fd_sc_hd__buf_2
X_63312_ _60454_/A _63312_/B _63312_/C _63237_/X _63312_/X sky130_fd_sc_hd__and4_4
X_48246_ _47965_/B _53520_/B sky130_fd_sc_hd__buf_2
X_60524_ _60488_/B _60476_/D _60445_/A _60524_/Y sky130_fd_sc_hd__o21ai_4
X_67080_ _87934_/Q _67056_/X _67032_/X _67079_/X _67080_/X sky130_fd_sc_hd__a211o_4
X_79066_ _79027_/A _79042_/A _79034_/A _79057_/C _79066_/X sky130_fd_sc_hd__and4_4
X_45458_ _45455_/Y _45439_/X _45390_/X _45457_/Y _45458_/X sky130_fd_sc_hd__a211o_4
X_64292_ _64292_/A _64301_/B _64292_/Y sky130_fd_sc_hd__nor2_4
X_76278_ _81258_/Q _81514_/D _76278_/Y sky130_fd_sc_hd__nand2_4
X_66031_ _65553_/X _66062_/B _65556_/C _66031_/Y sky130_fd_sc_hd__nand3_4
X_78017_ _78018_/A _78018_/B _78017_/X sky130_fd_sc_hd__xor2_4
X_44409_ _44404_/X _44405_/X _41520_/X _87123_/Q _44406_/X _44410_/A
+ sky130_fd_sc_hd__o32ai_4
X_63243_ _63236_/Y _63238_/X _63239_/X _63241_/X _63242_/X _63243_/Y
+ sky130_fd_sc_hd__o41ai_4
X_75229_ _75225_/Y _75227_/Y _75224_/Y _75230_/B sky130_fd_sc_hd__o21ai_4
X_48177_ _49173_/A _48184_/A sky130_fd_sc_hd__buf_2
X_60455_ _60572_/A _60572_/B _60572_/C _60476_/D _60562_/B _60455_/Y
+ sky130_fd_sc_hd__a32oi_4
X_45389_ _45389_/A _45389_/X sky130_fd_sc_hd__buf_2
X_47128_ _47128_/A _47128_/X sky130_fd_sc_hd__buf_2
X_63174_ _79363_/A _63130_/X _63173_/Y _84347_/D sky130_fd_sc_hd__a21o_4
X_60386_ _60386_/A _60418_/D _60387_/C sky130_fd_sc_hd__and2_4
X_62125_ _59858_/A _61637_/X _62124_/X _62125_/X sky130_fd_sc_hd__a21o_4
X_47059_ _47067_/A _47039_/B _47048_/C _52831_/D _47059_/X sky130_fd_sc_hd__and4_4
X_67982_ _67388_/X _68089_/A sky130_fd_sc_hd__buf_2
X_79968_ _79957_/A _79957_/B _79957_/C _79968_/Y sky130_fd_sc_hd__a21boi_4
X_69721_ _44148_/A _69766_/A sky130_fd_sc_hd__buf_2
X_50070_ _50066_/Y _50068_/X _50069_/X _50070_/Y sky130_fd_sc_hd__a21oi_4
X_66933_ _87120_/Q _66833_/X _66834_/X _66932_/X _66933_/X sky130_fd_sc_hd__a211o_4
X_62056_ _59858_/A _61580_/X _62055_/X _62056_/X sky130_fd_sc_hd__a21o_4
X_78919_ _78919_/A _78918_/Y _78920_/B sky130_fd_sc_hd__xor2_4
X_79899_ _79899_/A _79898_/Y _80264_/A sky130_fd_sc_hd__nand2_4
X_61007_ _59875_/A _63765_/A _61008_/A sky130_fd_sc_hd__nor2_4
X_81930_ _82234_/CLK _77819_/Y _81930_/Q sky130_fd_sc_hd__dfxtp_4
X_69652_ _69680_/A _88333_/Q _69652_/X sky130_fd_sc_hd__and2_4
X_66864_ _66840_/X _86826_/Q _66864_/X sky130_fd_sc_hd__and2_4
X_68603_ _69357_/A _68604_/A sky130_fd_sc_hd__buf_2
X_65815_ _65789_/X _65255_/Y _65814_/Y _65815_/Y sky130_fd_sc_hd__o21ai_4
X_81861_ _80708_/CLK _81861_/D _81861_/Q sky130_fd_sc_hd__dfxtp_4
X_69583_ _68934_/X _69583_/B _69583_/Y sky130_fd_sc_hd__nor2_4
X_66795_ _66795_/A _66795_/B _66795_/X sky130_fd_sc_hd__and2_4
X_83600_ _86145_/CLK _83600_/D _83600_/Q sky130_fd_sc_hd__dfxtp_4
X_80812_ _81134_/CLK _83956_/Q _75806_/B sky130_fd_sc_hd__dfxtp_4
X_68534_ _69014_/A _68560_/A sky130_fd_sc_hd__buf_2
X_53760_ _53757_/Y _53747_/X _53759_/X _53760_/Y sky130_fd_sc_hd__a21oi_4
X_65746_ _65742_/Y _65681_/X _65745_/Y _65746_/X sky130_fd_sc_hd__a21o_4
X_84580_ _84583_/CLK _60728_/X _84580_/Q sky130_fd_sc_hd__dfxtp_4
X_50972_ _86097_/Q _50965_/X _50971_/Y _50972_/Y sky130_fd_sc_hd__o21ai_4
X_62958_ _61652_/B _62936_/X _62982_/C _62908_/X _62958_/Y sky130_fd_sc_hd__nand4_4
X_81792_ _86807_/CLK _75955_/X _48373_/A sky130_fd_sc_hd__dfxtp_4
X_52711_ _52684_/A _52711_/X sky130_fd_sc_hd__buf_2
X_83531_ _86203_/CLK _71336_/Y _83531_/Q sky130_fd_sc_hd__dfxtp_4
X_61909_ _58322_/A _61909_/X sky130_fd_sc_hd__buf_2
X_80743_ _80961_/CLK _80743_/D _75062_/A sky130_fd_sc_hd__dfxtp_4
X_68465_ _64615_/A _68465_/B _68465_/Y sky130_fd_sc_hd__nor2_4
X_53691_ _53733_/A _53720_/B sky130_fd_sc_hd__buf_2
X_65677_ _65984_/A _65828_/B sky130_fd_sc_hd__buf_2
X_62889_ _61570_/B _62858_/X _62859_/X _62889_/D _62889_/Y sky130_fd_sc_hd__nand4_4
X_55430_ _55683_/A _55429_/Y _55373_/Y _55430_/Y sky130_fd_sc_hd__nand3_4
X_67416_ _87920_/Q _67414_/X _67391_/X _67415_/X _67416_/X sky130_fd_sc_hd__a211o_4
X_86250_ _83613_/CLK _86250_/D _86250_/Q sky130_fd_sc_hd__dfxtp_4
X_52642_ _85781_/Q _52629_/X _52641_/Y _52642_/Y sky130_fd_sc_hd__o21ai_4
X_64628_ _64589_/X _85568_/Q _64591_/X _64627_/X _64628_/X sky130_fd_sc_hd__a211o_4
X_83462_ _83464_/CLK _83462_/D _83462_/Q sky130_fd_sc_hd__dfxtp_4
X_80674_ _81104_/CLK _80674_/D _75086_/A sky130_fd_sc_hd__dfxtp_4
X_68396_ _69651_/A _69877_/A sky130_fd_sc_hd__buf_2
X_85201_ _85297_/CLK _85201_/D _85201_/Q sky130_fd_sc_hd__dfxtp_4
X_82413_ _82248_/CLK _82445_/Q _78458_/A sky130_fd_sc_hd__dfxtp_4
X_55361_ _56689_/A _55360_/X _55443_/A sky130_fd_sc_hd__nand2_4
X_86181_ _86499_/CLK _86181_/D _86181_/Q sky130_fd_sc_hd__dfxtp_4
X_67347_ _67343_/X _67346_/X _67322_/X _67347_/X sky130_fd_sc_hd__a21o_4
XPHY_506 sky130_fd_sc_hd__decap_3
X_52573_ _51396_/A _52573_/B _50918_/A _52573_/X sky130_fd_sc_hd__and3_4
X_64559_ _64689_/A _64741_/B _79529_/B _64559_/Y sky130_fd_sc_hd__nor3_4
X_83393_ _85505_/CLK _71742_/Y _83393_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_517 sky130_fd_sc_hd__decap_3
XPHY_528 sky130_fd_sc_hd__decap_3
X_57100_ _57097_/X _56571_/X _45408_/A _57099_/X _57100_/X sky130_fd_sc_hd__a2bb2o_4
X_54312_ _54312_/A _54325_/B _54312_/C _54312_/D _54312_/X sky130_fd_sc_hd__and4_4
XPHY_539 sky130_fd_sc_hd__decap_3
X_85132_ _85067_/CLK _56799_/Y _85132_/Q sky130_fd_sc_hd__dfxtp_4
X_51524_ _51514_/A _53050_/B _51524_/Y sky130_fd_sc_hd__nand2_4
X_58080_ _58080_/A _58576_/A sky130_fd_sc_hd__buf_2
X_82344_ _82558_/CLK _77094_/X _48094_/A sky130_fd_sc_hd__dfxtp_4
X_55292_ _55265_/Y _55289_/X _55291_/Y _55292_/X sky130_fd_sc_hd__o21a_4
X_67278_ _67039_/X _67278_/X sky130_fd_sc_hd__buf_2
X_57031_ _57031_/A _57031_/Y sky130_fd_sc_hd__inv_2
X_69017_ _68660_/X _69017_/X sky130_fd_sc_hd__buf_2
X_54243_ _54230_/A _53076_/B _54243_/Y sky130_fd_sc_hd__nand2_4
X_66229_ _65767_/X _66135_/B _65770_/X _66229_/Y sky130_fd_sc_hd__nand3_4
X_85063_ _85128_/CLK _57207_/X _85063_/Q sky130_fd_sc_hd__dfxtp_4
X_51455_ _86007_/Q _51429_/X _51454_/Y _51455_/Y sky130_fd_sc_hd__o21ai_4
X_82275_ _82103_/CLK _77013_/B _82275_/Q sky130_fd_sc_hd__dfxtp_4
X_84014_ _84014_/CLK _68199_/X _84014_/Q sky130_fd_sc_hd__dfxtp_4
X_50406_ _86207_/Q _50403_/X _50405_/Y _50406_/Y sky130_fd_sc_hd__o21ai_4
X_81226_ _81224_/CLK _81034_/Q _47747_/A sky130_fd_sc_hd__dfxtp_4
X_54174_ _54170_/Y _54171_/X _54173_/X _85491_/D sky130_fd_sc_hd__a21oi_4
X_51386_ _48808_/A _51789_/A sky130_fd_sc_hd__buf_2
X_53125_ _53133_/A _53133_/B _53133_/C _53125_/D _53125_/X sky130_fd_sc_hd__and4_4
X_50337_ _50537_/A _50510_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_663_0_CLK clkbuf_9_331_0_CLK/X _88128_/CLK sky130_fd_sc_hd__clkbuf_1
X_81157_ _81179_/CLK _74868_/B _40530_/B sky130_fd_sc_hd__dfxtp_4
X_58982_ _58982_/A _58982_/X sky130_fd_sc_hd__buf_2
X_80108_ _80101_/X _80108_/B _80108_/Y sky130_fd_sc_hd__nand2_4
X_57933_ _57922_/Y _57758_/X _57929_/X _57932_/X _57933_/Y sky130_fd_sc_hd__a22oi_4
X_41070_ _41069_/Y _41070_/X sky130_fd_sc_hd__buf_2
X_53056_ _53111_/A _53056_/X sky130_fd_sc_hd__buf_2
X_69919_ _73438_/A _68463_/X _69478_/X _69918_/Y _69919_/X sky130_fd_sc_hd__a211o_4
X_50268_ _50240_/A _50268_/B _50268_/Y sky130_fd_sc_hd__nand2_4
X_85965_ _84802_/CLK _51685_/Y _85965_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_154_0_CLK clkbuf_8_77_0_CLK/X clkbuf_9_154_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_81088_ _80681_/CLK _81120_/Q _75541_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_81_0_CLK clkbuf_8_40_0_CLK/X clkbuf_9_81_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_52007_ _51982_/X _48257_/B _52007_/Y sky130_fd_sc_hd__nand2_4
X_87704_ _87221_/CLK _42814_/X _67972_/B sky130_fd_sc_hd__dfxtp_4
X_72930_ _72806_/X _86203_/Q _72746_/X _72929_/X _72930_/X sky130_fd_sc_hd__a211o_4
X_84916_ _84915_/CLK _58169_/X _58166_/A sky130_fd_sc_hd__dfxtp_4
X_80039_ _84933_/Q _84181_/Q _80039_/X sky130_fd_sc_hd__xor2_4
X_57864_ _57861_/Y _57863_/Y _57829_/X _57864_/X sky130_fd_sc_hd__a21o_4
X_50199_ _50187_/X _50712_/B _50199_/Y sky130_fd_sc_hd__nand2_4
X_85896_ _86210_/CLK _85896_/D _85896_/Q sky130_fd_sc_hd__dfxtp_4
X_59603_ _59603_/A _72569_/C sky130_fd_sc_hd__buf_2
Xclkbuf_10_678_0_CLK clkbuf_9_339_0_CLK/X _87898_/CLK sky130_fd_sc_hd__clkbuf_1
X_56815_ _56725_/B _56806_/Y _56814_/Y _85131_/D sky130_fd_sc_hd__o21ai_4
X_87635_ _87995_/CLK _87635_/D _66567_/B sky130_fd_sc_hd__dfxtp_4
X_72861_ _73067_/A _72861_/X sky130_fd_sc_hd__buf_2
X_84847_ _83457_/CLK _84847_/D _84847_/Q sky130_fd_sc_hd__dfxtp_4
X_57795_ _72417_/A _57795_/X sky130_fd_sc_hd__buf_2
X_74600_ _74600_/A _74600_/X sky130_fd_sc_hd__buf_2
X_71812_ _71805_/X _83367_/Q _71811_/X _83367_/D sky130_fd_sc_hd__a21o_4
X_59534_ _59546_/A _59563_/A _59519_/C _59535_/A sky130_fd_sc_hd__nand3_4
Xclkbuf_9_169_0_CLK clkbuf_8_84_0_CLK/X clkbuf_9_169_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_44760_ _44760_/A _86969_/D sky130_fd_sc_hd__inv_2
X_56746_ _56725_/Y _56745_/X _85135_/D sky130_fd_sc_hd__nand2_4
X_75580_ _75579_/Y _80819_/Q _75580_/Y sky130_fd_sc_hd__nand2_4
X_87566_ _87824_/CLK _87566_/D _43126_/A sky130_fd_sc_hd__dfxtp_4
X_41972_ _41972_/A _41972_/Y sky130_fd_sc_hd__inv_2
X_53958_ _85534_/Q _53955_/X _53957_/Y _53958_/Y sky130_fd_sc_hd__o21ai_4
X_72792_ _72790_/X _72791_/Y _72766_/X _72792_/Y sky130_fd_sc_hd__a21oi_4
X_84778_ _84778_/CLK _58995_/Y _62186_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_96_0_CLK clkbuf_9_97_0_CLK/A clkbuf_9_96_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_43711_ _40848_/X _43698_/X _69780_/B _43700_/X _43712_/A sky130_fd_sc_hd__a2bb2o_4
X_74531_ _74531_/A _74531_/B _74531_/C _74531_/D _74531_/Y sky130_fd_sc_hd__nand4_4
X_86517_ _85581_/CLK _86517_/D _73096_/B sky130_fd_sc_hd__dfxtp_4
X_40923_ _40923_/A _40842_/X _40923_/X sky130_fd_sc_hd__or2_4
X_52909_ _52906_/Y _52892_/X _52908_/X _85733_/D sky130_fd_sc_hd__a21oi_4
X_71743_ _71026_/A _71744_/C sky130_fd_sc_hd__buf_2
X_59465_ _59463_/Y _59478_/B _59465_/Y sky130_fd_sc_hd__nand2_4
X_83729_ _85379_/CLK _70671_/X _83729_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_601_0_CLK clkbuf_9_300_0_CLK/X _81985_/CLK sky130_fd_sc_hd__clkbuf_1
X_44691_ _44691_/A _44691_/Y sky130_fd_sc_hd__inv_2
X_56677_ _56700_/C _56676_/Y _56679_/B sky130_fd_sc_hd__nor2_4
X_87497_ _88012_/CLK _43289_/X _87497_/Q sky130_fd_sc_hd__dfxtp_4
X_53889_ _53887_/Y _53829_/X _53888_/X _85548_/D sky130_fd_sc_hd__a21oi_4
X_46430_ _46279_/A _46430_/X sky130_fd_sc_hd__buf_2
X_58416_ _58406_/X _83366_/Q _58415_/Y _84854_/D sky130_fd_sc_hd__o21a_4
X_77250_ _77250_/A _77252_/A sky130_fd_sc_hd__inv_2
X_55628_ _44070_/B _55628_/B _55628_/Y sky130_fd_sc_hd__nor2_4
X_43642_ _40682_/A _43634_/X _43641_/Y _43636_/X _43642_/X sky130_fd_sc_hd__a2bb2o_4
X_74462_ _83061_/Q _74441_/X _74461_/Y _74462_/Y sky130_fd_sc_hd__o21ai_4
X_86448_ _85554_/CLK _49062_/Y _65066_/B sky130_fd_sc_hd__dfxtp_4
X_40854_ _40853_/X _40854_/X sky130_fd_sc_hd__buf_2
X_71674_ _71680_/A _71671_/X _71297_/X _71674_/Y sky130_fd_sc_hd__nand3_4
X_59396_ _63127_/A _59399_/A sky130_fd_sc_hd__buf_2
X_76201_ _76200_/A _76200_/B _76201_/Y sky130_fd_sc_hd__nand2_4
X_73413_ _73411_/X _73412_/Y _73367_/X _73413_/Y sky130_fd_sc_hd__a21oi_4
X_46361_ _46361_/A _52468_/B sky130_fd_sc_hd__buf_2
X_70625_ _70423_/X _71162_/B _70625_/Y sky130_fd_sc_hd__nor2_4
X_58347_ _63295_/A _58348_/A sky130_fd_sc_hd__buf_2
X_77181_ _77184_/A _77181_/B _77182_/B sky130_fd_sc_hd__xor2_4
X_43573_ _40524_/X _43560_/X _87353_/Q _43561_/X _87353_/D sky130_fd_sc_hd__a2bb2o_4
X_55559_ _85115_/Q _55522_/X _55506_/X _55558_/Y _55559_/X sky130_fd_sc_hd__a211o_4
X_74393_ _74408_/A _53647_/B _74393_/Y sky130_fd_sc_hd__nand2_4
X_86379_ _86381_/CLK _86379_/D _86379_/Q sky130_fd_sc_hd__dfxtp_4
X_40785_ _82877_/Q _40847_/B _40785_/X sky130_fd_sc_hd__or2_4
X_48100_ _50360_/A _48099_/X _48723_/C _48100_/X sky130_fd_sc_hd__and3_4
X_45312_ _55702_/B _45281_/X _45311_/X _45312_/X sky130_fd_sc_hd__o21a_4
X_76132_ _81726_/D _76133_/B _76132_/X sky130_fd_sc_hd__or2_4
X_88118_ _88376_/CLK _88118_/D _88118_/Q sky130_fd_sc_hd__dfxtp_4
X_42524_ _42524_/A _87835_/D sky130_fd_sc_hd__inv_2
X_49080_ _49080_/A _53879_/B _49080_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_616_0_CLK clkbuf_9_308_0_CLK/X _81154_/CLK sky130_fd_sc_hd__clkbuf_1
X_73344_ _73343_/X _73344_/X sky130_fd_sc_hd__buf_2
X_46292_ _46719_/A _46292_/X sky130_fd_sc_hd__buf_2
X_70556_ _70533_/X _83750_/Q _70555_/Y _70556_/X sky130_fd_sc_hd__a21o_4
X_58278_ _58271_/X _83442_/Q _58277_/Y _84890_/D sky130_fd_sc_hd__o21a_4
X_48031_ _53552_/B _50328_/B sky130_fd_sc_hd__buf_2
X_57229_ _45883_/B _72710_/A sky130_fd_sc_hd__buf_2
X_45243_ _85291_/Q _45194_/X _45229_/X _45243_/X sky130_fd_sc_hd__o21a_4
X_76063_ _76063_/A _76063_/B _76063_/C _76064_/B sky130_fd_sc_hd__and3_4
X_88049_ _88056_/CLK _88049_/D _88049_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_107_0_CLK clkbuf_8_53_0_CLK/X clkbuf_9_107_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_42455_ _42454_/Y _87859_/D sky130_fd_sc_hd__inv_2
X_73275_ _73275_/A _73228_/B _73275_/Y sky130_fd_sc_hd__nor2_4
X_70487_ _70466_/Y _83763_/Q _70486_/X _83763_/D sky130_fd_sc_hd__a21o_4
Xclkbuf_9_34_0_CLK clkbuf_9_35_0_CLK/A clkbuf_9_34_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_75014_ _80953_/Q _75014_/B _75014_/X sky130_fd_sc_hd__xor2_4
X_41406_ _41406_/A _41379_/X _41406_/X sky130_fd_sc_hd__or2_4
X_60240_ _60239_/X _60241_/A sky130_fd_sc_hd__inv_2
X_72226_ _72180_/X _85336_/Q _72225_/X _72226_/X sky130_fd_sc_hd__o21a_4
X_45174_ _55821_/B _45131_/X _45161_/X _45174_/X sky130_fd_sc_hd__o21a_4
X_42386_ _42386_/A _87889_/D sky130_fd_sc_hd__inv_2
X_44125_ _72814_/A _73352_/A sky130_fd_sc_hd__buf_2
X_79822_ _79829_/B _79822_/B _79822_/Y sky130_fd_sc_hd__xnor2_4
X_41337_ _41336_/X _41337_/X sky130_fd_sc_hd__buf_2
X_60171_ _60171_/A _60171_/B _60172_/A sky130_fd_sc_hd__and2_4
X_72157_ _72155_/X _85694_/Q _72156_/X _72157_/X sky130_fd_sc_hd__o21a_4
X_49982_ _86287_/Q _49960_/X _49981_/Y _49982_/Y sky130_fd_sc_hd__o21ai_4
X_71108_ _71101_/X _71230_/B _70890_/D _71108_/Y sky130_fd_sc_hd__nand3_4
X_48933_ _64759_/B _48896_/X _48932_/Y _48933_/Y sky130_fd_sc_hd__o21ai_4
X_44056_ _55125_/A _55152_/A sky130_fd_sc_hd__buf_2
X_79753_ _79741_/X _79742_/X _79752_/Y _79757_/A sky130_fd_sc_hd__a21boi_4
X_41268_ _41267_/Y _41268_/X sky130_fd_sc_hd__buf_2
X_72088_ _72075_/A _50183_/B _72088_/Y sky130_fd_sc_hd__nand2_4
X_76965_ _76965_/A _76965_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_9_49_0_CLK clkbuf_9_49_0_CLK/A clkbuf_9_49_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_43007_ _43006_/Y _87607_/D sky130_fd_sc_hd__inv_2
X_78704_ _78685_/A _78702_/Y _78703_/Y _78742_/B sky130_fd_sc_hd__a21bo_4
X_63930_ _63960_/A _63960_/B _80133_/B _63930_/Y sky130_fd_sc_hd__nor3_4
X_71039_ _71183_/A _71030_/B _71030_/C _71039_/D _71039_/Y sky130_fd_sc_hd__nand4_4
X_75916_ _61174_/C _84386_/Q _75916_/X sky130_fd_sc_hd__xor2_4
X_48864_ _86468_/Q _48861_/X _48863_/Y _48864_/Y sky130_fd_sc_hd__o21ai_4
X_79684_ _79660_/A _79659_/Y _79669_/X _79672_/Y _79684_/X sky130_fd_sc_hd__o22a_4
X_41199_ _41198_/Y _41199_/X sky130_fd_sc_hd__buf_2
X_76896_ _76894_/Y _76895_/Y _76899_/A sky130_fd_sc_hd__nor2_4
Xclkbuf_3_7_0_CLK clkbuf_3_6_0_CLK/A clkbuf_3_7_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_47815_ _49374_/A _49364_/B _50886_/C _53257_/D _47815_/X sky130_fd_sc_hd__and4_4
X_78635_ _78634_/X _78637_/B sky130_fd_sc_hd__inv_2
X_63861_ _61419_/X _63877_/B _63814_/C _63877_/D _63861_/Y sky130_fd_sc_hd__nand4_4
X_75847_ _81023_/Q _75848_/B sky130_fd_sc_hd__inv_2
X_48795_ _52139_/A _48833_/A sky130_fd_sc_hd__buf_2
X_65600_ _64908_/X _65647_/B _64910_/X _65600_/Y sky130_fd_sc_hd__nand3_4
X_62812_ _62773_/X _62812_/B _61939_/X _62812_/Y sky130_fd_sc_hd__nand3_4
X_47746_ _47792_/A _47777_/B sky130_fd_sc_hd__buf_2
X_66580_ _66568_/X _66578_/X _66579_/X _66580_/X sky130_fd_sc_hd__a21o_4
X_78566_ _78566_/A _82720_/Q _78569_/B sky130_fd_sc_hd__nor2_4
X_44958_ _45389_/A _45720_/A sky130_fd_sc_hd__buf_2
X_63792_ _64012_/A _63793_/D sky130_fd_sc_hd__buf_2
X_75778_ _75778_/A _75778_/Y sky130_fd_sc_hd__inv_2
X_65531_ _65559_/A _65546_/B _65531_/C _65531_/X sky130_fd_sc_hd__and3_4
X_77517_ _77517_/A _77519_/A sky130_fd_sc_hd__inv_2
X_43909_ _41361_/X _43907_/X _67667_/B _43908_/X _43909_/X sky130_fd_sc_hd__a2bb2o_4
X_62743_ _61419_/X _62743_/B _62742_/X _62729_/D _62743_/Y sky130_fd_sc_hd__nand4_4
X_74729_ _74729_/A _74796_/B _74796_/C _71016_/A _74729_/Y sky130_fd_sc_hd__nand4_4
X_47677_ _47671_/Y _47651_/X _47676_/X _47677_/Y sky130_fd_sc_hd__a21oi_4
X_78497_ _78460_/A _78463_/A _78473_/X _78497_/X sky130_fd_sc_hd__a21o_4
X_44889_ _44889_/A _44889_/X sky130_fd_sc_hd__buf_2
X_49416_ _49416_/A _49444_/A sky130_fd_sc_hd__buf_2
X_68250_ _84001_/Q _68238_/X _68249_/X _68250_/X sky130_fd_sc_hd__a21bo_4
X_46628_ _74509_/B _46670_/A sky130_fd_sc_hd__buf_2
X_65462_ _64655_/X _65340_/X _64659_/X _65462_/Y sky130_fd_sc_hd__nand3_4
X_77448_ _77444_/Y _77446_/Y _77447_/A _77448_/Y sky130_fd_sc_hd__o21ai_4
X_62674_ _62670_/X _62652_/X _62673_/Y _62674_/Y sky130_fd_sc_hd__a21oi_4
X_67201_ _67250_/A _67201_/B _67201_/X sky130_fd_sc_hd__and2_4
X_64413_ _64380_/X _84864_/Q _64381_/X _64413_/Y sky130_fd_sc_hd__nand3_4
X_49347_ _49345_/Y _49326_/X _49346_/Y _86405_/D sky130_fd_sc_hd__a21boi_4
X_61625_ _61623_/X _61576_/X _61624_/Y _61625_/Y sky130_fd_sc_hd__a21oi_4
X_68181_ _67135_/X _67137_/X _68169_/X _68181_/Y sky130_fd_sc_hd__a21oi_4
X_46559_ _46525_/X _49161_/A _46558_/X _51376_/B sky130_fd_sc_hd__o21ai_4
X_65393_ _65342_/X _83283_/Q _65391_/X _65392_/X _65393_/X sky130_fd_sc_hd__a211o_4
X_77379_ _77380_/A _82093_/D _77382_/B sky130_fd_sc_hd__nor2_4
X_67132_ _87868_/Q _67056_/X _67032_/X _67131_/X _67132_/X sky130_fd_sc_hd__a211o_4
X_79118_ _78997_/B _82519_/D sky130_fd_sc_hd__inv_2
X_64344_ _64285_/A _64344_/X sky130_fd_sc_hd__buf_2
X_61556_ _61554_/X _61517_/X _61555_/Y _61556_/Y sky130_fd_sc_hd__a21oi_4
X_49278_ _49276_/Y _49271_/X _49277_/Y _86419_/D sky130_fd_sc_hd__a21boi_4
X_80390_ _84755_/Q _80397_/B _80390_/X sky130_fd_sc_hd__xor2_4
X_60507_ _63247_/A _60508_/A sky130_fd_sc_hd__buf_2
X_48229_ _48229_/A _53504_/B _48229_/Y sky130_fd_sc_hd__nand2_4
X_67063_ _67062_/X _67087_/A sky130_fd_sc_hd__buf_2
X_79049_ _79049_/A _79057_/B sky130_fd_sc_hd__inv_2
X_64275_ _64275_/A _64275_/B _64274_/X _64275_/X sky130_fd_sc_hd__and3_4
X_61487_ _61518_/A _61518_/B _84477_/Q _61487_/Y sky130_fd_sc_hd__nor3_4
X_66014_ _66010_/X _65967_/B _66013_/X _66014_/Y sky130_fd_sc_hd__nand3_4
X_51240_ _51240_/A _49212_/B _51240_/Y sky130_fd_sc_hd__nand2_4
X_63226_ _63203_/X _84838_/Q _63204_/X _63239_/D _63226_/X sky130_fd_sc_hd__and4_4
X_82060_ _81507_/CLK _82060_/D _77813_/A sky130_fd_sc_hd__dfxtp_4
X_60438_ _60438_/A _60583_/A sky130_fd_sc_hd__buf_2
X_81011_ _84223_/CLK _84219_/Q _81011_/Q sky130_fd_sc_hd__dfxtp_4
X_51171_ _51177_/A _51160_/B _51192_/C _52861_/D _51171_/X sky130_fd_sc_hd__and4_4
X_63157_ _60469_/X _63157_/X sky130_fd_sc_hd__buf_2
X_60369_ _79553_/A _60132_/X _60331_/D _60247_/Y _60369_/X sky130_fd_sc_hd__a2bb2o_4
X_50122_ _50106_/A _72025_/B _50122_/X sky130_fd_sc_hd__and2_4
X_62108_ _61949_/A _62170_/B _62158_/C _63292_/B _62108_/X sky130_fd_sc_hd__and4_4
X_67965_ _87385_/Q _67868_/X _67938_/X _67964_/X _67965_/X sky130_fd_sc_hd__a211o_4
X_63088_ _63088_/A _64295_/C _63087_/X _63077_/D _63088_/X sky130_fd_sc_hd__and4_4
X_69704_ _73024_/A _66608_/X _57800_/A _69703_/X _69704_/X sky130_fd_sc_hd__a211o_4
X_50053_ _86273_/Q _48861_/X _50052_/Y _50053_/Y sky130_fd_sc_hd__o21ai_4
X_54930_ _54919_/X _47771_/Y _54930_/Y sky130_fd_sc_hd__nand2_4
X_66916_ _66840_/X _86824_/Q _66916_/X sky130_fd_sc_hd__and2_4
X_62039_ _83245_/Q _63611_/A sky130_fd_sc_hd__inv_2
X_85750_ _85751_/CLK _52812_/Y _85750_/Q sky130_fd_sc_hd__dfxtp_4
X_82962_ _82774_/CLK _82770_/Q _46762_/A sky130_fd_sc_hd__dfxtp_4
X_67896_ _86952_/Q _67825_/X _67872_/X _67895_/X _67896_/X sky130_fd_sc_hd__a211o_4
X_84701_ _84713_/CLK _59786_/Y _80497_/A sky130_fd_sc_hd__dfxtp_4
X_81913_ _82005_/CLK _81913_/D _81913_/Q sky130_fd_sc_hd__dfxtp_4
X_69635_ _68360_/X _42555_/Y _69635_/Y sky130_fd_sc_hd__nor2_4
X_54861_ _54807_/A _54883_/A sky130_fd_sc_hd__buf_2
X_66847_ _66844_/X _66846_/X _66706_/X _66847_/Y sky130_fd_sc_hd__a21oi_4
X_85681_ _84797_/CLK _85681_/D _85681_/Q sky130_fd_sc_hd__dfxtp_4
X_82893_ _82906_/CLK _78160_/B _82893_/Q sky130_fd_sc_hd__dfxtp_4
X_56600_ _56600_/A _56600_/X sky130_fd_sc_hd__buf_2
X_87420_ _82317_/CLK _43440_/X _87420_/Q sky130_fd_sc_hd__dfxtp_4
X_53812_ _53791_/A _71987_/B _53812_/Y sky130_fd_sc_hd__nand2_4
X_84632_ _84620_/CLK _60326_/X _79700_/A sky130_fd_sc_hd__dfxtp_4
X_57580_ _46653_/A _72009_/A sky130_fd_sc_hd__buf_2
X_69566_ _87571_/Q _69506_/X _66349_/X _69565_/X _69566_/X sky130_fd_sc_hd__a211o_4
X_81844_ _81094_/CLK _81876_/Q _77488_/A sky130_fd_sc_hd__dfxtp_4
X_54792_ _51340_/A _54900_/A sky130_fd_sc_hd__buf_2
X_66778_ _88395_/Q _66751_/X _66682_/X _66777_/X _66778_/X sky130_fd_sc_hd__a211o_4
X_56531_ _56533_/A _56533_/B _85160_/Q _56531_/Y sky130_fd_sc_hd__nand3_4
X_68517_ _68517_/A _68517_/X sky130_fd_sc_hd__buf_2
X_87351_ _86814_/CLK _87351_/D _87351_/Q sky130_fd_sc_hd__dfxtp_4
X_53743_ _48841_/A _53748_/B _53748_/C _53743_/X sky130_fd_sc_hd__and3_4
X_65729_ _65726_/Y _65681_/X _65728_/Y _84182_/D sky130_fd_sc_hd__a21o_4
X_84563_ _84454_/CLK _60803_/Y _84563_/Q sky130_fd_sc_hd__dfxtp_4
X_50955_ _50938_/X _46740_/X _50955_/Y sky130_fd_sc_hd__nand2_4
X_81775_ _84014_/CLK _76069_/X _81775_/Q sky130_fd_sc_hd__dfxtp_4
X_69497_ _69322_/A _88281_/Q _69497_/X sky130_fd_sc_hd__and2_4
X_86302_ _86303_/CLK _49905_/Y _72160_/B sky130_fd_sc_hd__dfxtp_4
X_59250_ _59177_/X _86061_/Q _59249_/X _59250_/Y sky130_fd_sc_hd__o21ai_4
X_83514_ _83514_/CLK _71394_/X _83514_/Q sky130_fd_sc_hd__dfxtp_4
X_56462_ _56528_/A _56462_/X sky130_fd_sc_hd__buf_2
X_80726_ _80676_/CLK _75912_/X _80694_/D sky130_fd_sc_hd__dfxtp_4
X_68448_ _68403_/A _87760_/Q _68448_/X sky130_fd_sc_hd__and2_4
X_87282_ _88084_/CLK _87282_/D _87282_/Q sky130_fd_sc_hd__dfxtp_4
X_53674_ _53662_/X _73073_/A _53674_/Y sky130_fd_sc_hd__nand2_4
X_84494_ _84623_/CLK _61266_/X _61265_/C sky130_fd_sc_hd__dfxtp_4
X_50886_ _50257_/X _50045_/X _50886_/C _52580_/D _50886_/X sky130_fd_sc_hd__and4_4
X_58201_ _58201_/A _58201_/X sky130_fd_sc_hd__buf_2
X_55413_ _55399_/X _55412_/Y _55409_/Y _55414_/B sky130_fd_sc_hd__nand3_4
X_86233_ _86235_/CLK _50276_/Y _86233_/Q sky130_fd_sc_hd__dfxtp_4
X_52625_ _85784_/Q _52601_/X _52624_/Y _52625_/Y sky130_fd_sc_hd__o21ai_4
X_59181_ _84763_/Q _59129_/X _59174_/X _59180_/X _84763_/D sky130_fd_sc_hd__a2bb2oi_4
X_83445_ _83763_/CLK _83445_/D _83445_/Q sky130_fd_sc_hd__dfxtp_4
X_56393_ _56035_/X _56378_/X _56392_/Y _85211_/D sky130_fd_sc_hd__o21ai_4
X_80657_ _80657_/CLK _74833_/Y _46114_/A sky130_fd_sc_hd__dfxtp_4
X_68379_ _69088_/A _68379_/X sky130_fd_sc_hd__buf_2
XPHY_303 sky130_fd_sc_hd__decap_3
XPHY_314 sky130_fd_sc_hd__decap_3
X_58132_ _58132_/A _58649_/B _58132_/Y sky130_fd_sc_hd__nor2_4
X_70410_ _70609_/A _70410_/Y sky130_fd_sc_hd__inv_2
XPHY_325 sky130_fd_sc_hd__decap_3
X_55344_ _85105_/Q _55342_/X _44046_/X _55343_/X _55344_/X sky130_fd_sc_hd__a211o_4
X_86164_ _85557_/CLK _50631_/Y _86164_/Q sky130_fd_sc_hd__dfxtp_4
X_40570_ _40569_/Y _88371_/D sky130_fd_sc_hd__inv_2
XPHY_336 sky130_fd_sc_hd__decap_3
X_52556_ _65298_/B _52549_/X _52555_/Y _52556_/Y sky130_fd_sc_hd__o21ai_4
X_71390_ _71372_/Y _83516_/Q _71389_/Y _83516_/D sky130_fd_sc_hd__a21o_4
X_83376_ _83756_/CLK _83376_/D _83376_/Q sky130_fd_sc_hd__dfxtp_4
X_80588_ _80588_/A _80588_/B _80589_/B sky130_fd_sc_hd__xor2_4
XPHY_347 sky130_fd_sc_hd__decap_3
XPHY_358 sky130_fd_sc_hd__decap_3
X_85115_ _85089_/CLK _85115_/D _85115_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_369 sky130_fd_sc_hd__decap_3
X_51507_ _51491_/A _53033_/B _51507_/Y sky130_fd_sc_hd__nand2_4
X_58063_ _58030_/X _85480_/Q _58062_/X _58063_/X sky130_fd_sc_hd__o21a_4
X_70341_ _70337_/X _74786_/A _70340_/X _83791_/D sky130_fd_sc_hd__a21o_4
X_82327_ _82327_/CLK _77152_/B _82327_/Q sky130_fd_sc_hd__dfxtp_4
X_55275_ _55285_/A _55274_/X _83318_/Q _55287_/A sky130_fd_sc_hd__a21o_4
X_86095_ _85778_/CLK _86095_/D _86095_/Q sky130_fd_sc_hd__dfxtp_4
X_52487_ _52319_/A _52487_/X sky130_fd_sc_hd__buf_2
X_57014_ _85101_/Q _56997_/X _57014_/Y sky130_fd_sc_hd__nor2_4
X_42240_ _42231_/X _42226_/X _41408_/X _87964_/Q _42228_/X _42241_/A
+ sky130_fd_sc_hd__o32ai_4
X_54226_ _54253_/A _54226_/X sky130_fd_sc_hd__buf_2
X_73060_ _88328_/Q _73059_/X _73007_/X _73060_/Y sky130_fd_sc_hd__o21ai_4
X_85046_ _85050_/CLK _57259_/X _45567_/A sky130_fd_sc_hd__dfxtp_4
X_51438_ _51456_/A _51421_/X _51438_/C _52967_/D _51438_/X sky130_fd_sc_hd__and4_4
X_70272_ _83815_/Q _74788_/A sky130_fd_sc_hd__inv_2
X_82258_ _82436_/CLK _80471_/X _82258_/Q sky130_fd_sc_hd__dfxtp_4
X_72011_ _72008_/Y _72009_/X _72010_/Y _72011_/Y sky130_fd_sc_hd__a21boi_4
X_81209_ _81996_/CLK _75066_/X _48967_/A sky130_fd_sc_hd__dfxtp_4
X_42171_ _42154_/X _42169_/X _41220_/X _87999_/Q _42170_/X _42172_/A
+ sky130_fd_sc_hd__o32ai_4
X_54157_ _54154_/Y _54144_/X _54156_/X _85494_/D sky130_fd_sc_hd__a21oi_4
X_51369_ _51365_/Y _51366_/X _51368_/X _86024_/D sky130_fd_sc_hd__a21oi_4
X_82189_ _84945_/CLK _82189_/D _82189_/Q sky130_fd_sc_hd__dfxtp_4
X_41122_ _41121_/X _41109_/X _88274_/Q _41110_/X _41122_/X sky130_fd_sc_hd__a2bb2o_4
X_53108_ _53106_/Y _53082_/X _53107_/X _85696_/D sky130_fd_sc_hd__a21oi_4
X_58965_ _58891_/X _86082_/Q _58964_/X _58965_/Y sky130_fd_sc_hd__o21ai_4
X_54088_ _54086_/Y _53472_/X _54087_/Y _54088_/Y sky130_fd_sc_hd__a21boi_4
X_86997_ _88363_/CLK _44696_/Y _86997_/Q sky130_fd_sc_hd__dfxtp_4
X_45930_ _72905_/A _45930_/X sky130_fd_sc_hd__buf_2
X_41053_ _40991_/X _41223_/A _41052_/X _41053_/X sky130_fd_sc_hd__o21a_4
X_53039_ _52630_/A _53147_/A sky130_fd_sc_hd__buf_2
X_57916_ _72476_/B _86004_/Q _57915_/X _57916_/Y sky130_fd_sc_hd__o21ai_4
X_76750_ _76738_/Y _76742_/Y _76744_/A _76750_/Y sky130_fd_sc_hd__a21boi_4
X_73962_ _73343_/X _73962_/X sky130_fd_sc_hd__buf_2
X_85948_ _82394_/CLK _85948_/D _85948_/Q sky130_fd_sc_hd__dfxtp_4
X_58896_ _58872_/A _58896_/B _58896_/Y sky130_fd_sc_hd__nor2_4
X_75701_ _75689_/A _75688_/Y _80910_/Q _80782_/D _75701_/X sky130_fd_sc_hd__a2bb2o_4
X_72913_ _72907_/X _72912_/X _72877_/X _72916_/A sky130_fd_sc_hd__a21o_4
X_45861_ _45861_/A _74702_/B sky130_fd_sc_hd__inv_2
X_57847_ _57801_/X _57843_/Y _57846_/Y _57822_/X _57809_/X _57847_/X
+ sky130_fd_sc_hd__o32a_4
X_76681_ _76678_/X _76680_/Y _81445_/D sky130_fd_sc_hd__xor2_4
X_73893_ _68727_/Y _73891_/X _73819_/X _73892_/Y _73893_/X sky130_fd_sc_hd__a211o_4
X_85879_ _85879_/CLK _85879_/D _73040_/B sky130_fd_sc_hd__dfxtp_4
X_47600_ _86617_/Q _47570_/X _47599_/Y _47600_/Y sky130_fd_sc_hd__o21ai_4
X_78420_ _78405_/Y _78402_/Y _78408_/C _78420_/X sky130_fd_sc_hd__o21a_4
X_44812_ _41642_/Y _43939_/X _67381_/B _43941_/X _86941_/D sky130_fd_sc_hd__a2bb2o_4
X_75632_ _75632_/A _75632_/B _75633_/B sky130_fd_sc_hd__nor2_4
X_87618_ _88387_/CLK _42987_/Y _87618_/Q sky130_fd_sc_hd__dfxtp_4
X_48580_ _48574_/Y _48517_/X _48579_/X _48580_/Y sky130_fd_sc_hd__a21oi_4
X_72844_ _72755_/X _83078_/Q _72785_/X _72843_/X _72844_/X sky130_fd_sc_hd__a211o_4
X_45792_ _85063_/Q _45792_/Y sky130_fd_sc_hd__inv_2
X_57778_ _58002_/A _72201_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_540_0_CLK clkbuf_9_270_0_CLK/X _83933_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_31_0_CLK clkbuf_6_31_0_CLK/A clkbuf_7_63_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_47531_ _81249_/Q _47532_/A sky130_fd_sc_hd__inv_2
X_59517_ _43959_/A _45941_/A _43959_/B _59517_/Y sky130_fd_sc_hd__nand3_4
X_78351_ _78325_/B _78339_/A _78338_/A _78353_/A sky130_fd_sc_hd__o21ai_4
X_56729_ _57140_/A _56729_/X sky130_fd_sc_hd__buf_2
X_44743_ _44740_/X _44741_/X _40743_/X _86979_/Q _44742_/X _44744_/A
+ sky130_fd_sc_hd__o32ai_4
X_75563_ _75561_/Y _75563_/B _81057_/D sky130_fd_sc_hd__nand2_4
X_87549_ _87813_/CLK _43174_/Y _73323_/A sky130_fd_sc_hd__dfxtp_4
X_41955_ _41955_/A _41955_/Y sky130_fd_sc_hd__inv_2
X_72775_ _56274_/X _72775_/X sky130_fd_sc_hd__buf_2
X_77302_ _77287_/A _77290_/B _77286_/A _77302_/Y sky130_fd_sc_hd__o21ai_4
X_74514_ _74512_/Y _46300_/X _74513_/Y _83050_/D sky130_fd_sc_hd__a21boi_4
X_40906_ _40903_/X _40904_/X _88313_/Q _40905_/X _88313_/D sky130_fd_sc_hd__a2bb2o_4
X_47462_ _47414_/A _47462_/X sky130_fd_sc_hd__buf_2
X_71726_ _58229_/Y _71718_/X _71725_/Y _71726_/Y sky130_fd_sc_hd__o21ai_4
X_59448_ _59448_/A _59444_/X _59448_/Y sky130_fd_sc_hd__nand2_4
X_78282_ _78282_/A _78281_/Y _78282_/X sky130_fd_sc_hd__or2_4
X_44674_ _44674_/A _44674_/Y sky130_fd_sc_hd__inv_2
X_75494_ _81086_/Q _75498_/A sky130_fd_sc_hd__inv_2
X_41886_ _42059_/A _41887_/A sky130_fd_sc_hd__buf_2
X_49201_ _72113_/A _50209_/A sky130_fd_sc_hd__buf_2
X_46413_ _86739_/Q _46364_/X _46412_/Y _46413_/Y sky130_fd_sc_hd__o21ai_4
X_77233_ _77233_/A _82082_/D _77233_/X sky130_fd_sc_hd__xor2_4
X_43625_ _43607_/A _43625_/X sky130_fd_sc_hd__buf_2
X_74445_ _48544_/A _74420_/X _74425_/X _74445_/X sky130_fd_sc_hd__and3_4
X_40837_ _82867_/Q _40847_/B _40837_/X sky130_fd_sc_hd__or2_4
Xclkbuf_10_555_0_CLK clkbuf_9_277_0_CLK/X _87473_/CLK sky130_fd_sc_hd__clkbuf_1
X_47393_ _47388_/Y _47364_/X _47392_/X _86640_/D sky130_fd_sc_hd__a21oi_4
X_59379_ _59346_/X _85634_/Q _59308_/X _59379_/X sky130_fd_sc_hd__o21a_4
X_71657_ _58508_/Y _71649_/X _71656_/Y _71657_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_6_46_0_CLK clkbuf_6_47_0_CLK/A clkbuf_7_93_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_61410_ _61409_/Y _61410_/Y sky130_fd_sc_hd__inv_2
X_49132_ _49080_/A _72079_/B _49132_/X sky130_fd_sc_hd__and2_4
X_46344_ _46326_/A _49245_/B _46344_/Y sky130_fd_sc_hd__nand2_4
X_70608_ _70997_/A _70719_/A sky130_fd_sc_hd__buf_2
X_77164_ _77173_/B _77173_/C _77167_/A sky130_fd_sc_hd__nand2_4
X_43556_ _43555_/Y _87362_/D sky130_fd_sc_hd__inv_2
X_62390_ _62623_/C _62390_/X sky130_fd_sc_hd__buf_2
X_74376_ _74374_/Y _74370_/X _74375_/X _74376_/Y sky130_fd_sc_hd__a21oi_4
X_40768_ _40767_/X _40754_/X _88339_/Q _40756_/X _88339_/D sky130_fd_sc_hd__a2bb2o_4
X_71588_ _71698_/A _71590_/B _71582_/X _71588_/Y sky130_fd_sc_hd__nor3_4
X_76115_ _76114_/X _76126_/A sky130_fd_sc_hd__buf_2
X_42507_ _42495_/X _42496_/X _40691_/X _87841_/Q _42506_/X _42508_/A
+ sky130_fd_sc_hd__o32ai_4
X_49063_ _83607_/Q _49064_/A sky130_fd_sc_hd__inv_2
X_61341_ _61317_/X _61368_/C sky130_fd_sc_hd__buf_2
X_73327_ _87049_/Q _73370_/B _73326_/X _73327_/Y sky130_fd_sc_hd__o21ai_4
X_46275_ _46262_/X _81215_/Q _46274_/X _46276_/A sky130_fd_sc_hd__o21ai_4
X_70539_ _70361_/A _71215_/C sky130_fd_sc_hd__buf_2
X_77095_ _77114_/B _82288_/D _77112_/A sky130_fd_sc_hd__xor2_4
X_43487_ _43472_/X _43475_/X _41705_/X _87397_/Q _43479_/X _43488_/A
+ sky130_fd_sc_hd__o32ai_4
X_40699_ _40784_/A _40760_/B sky130_fd_sc_hd__buf_2
X_48014_ _83544_/Q _48014_/Y sky130_fd_sc_hd__inv_2
X_45226_ _85196_/Q _45176_/X _45225_/X _45226_/Y sky130_fd_sc_hd__o21ai_4
X_64060_ _63238_/B _64145_/B _64029_/C _64029_/D _64064_/C sky130_fd_sc_hd__nand4_4
X_76046_ _81716_/D _76058_/B _76063_/A sky130_fd_sc_hd__xor2_4
X_42438_ _43161_/A _43146_/A sky130_fd_sc_hd__buf_2
X_61272_ _60296_/X _61272_/B _61151_/Y _61271_/Y _61272_/Y sky130_fd_sc_hd__nand4_4
X_73258_ _73206_/X _85870_/Q _73258_/X sky130_fd_sc_hd__and2_4
X_63011_ _58409_/A _63010_/X _60523_/X _59454_/A _60412_/X _63011_/Y
+ sky130_fd_sc_hd__o32ai_4
X_72209_ _59286_/A _72209_/X sky130_fd_sc_hd__buf_2
X_60223_ _60222_/X _60408_/A sky130_fd_sc_hd__buf_2
X_45157_ _45154_/X _45156_/Y _45125_/X _45157_/Y sky130_fd_sc_hd__a21oi_4
X_42369_ _42397_/A _42369_/X sky130_fd_sc_hd__buf_2
X_73189_ _48538_/Y _73188_/Y _73189_/X sky130_fd_sc_hd__xor2_4
X_44108_ _80666_/Q _44108_/X sky130_fd_sc_hd__buf_2
X_79805_ _84226_/Q _83274_/Q _79807_/A sky130_fd_sc_hd__xor2_4
X_60154_ _59875_/X _60062_/X _60049_/A _60000_/Y _60153_/Y _84650_/D
+ sky130_fd_sc_hd__o41a_4
X_49965_ _49963_/Y _49951_/X _49964_/X _86291_/D sky130_fd_sc_hd__a21oi_4
X_45088_ _55874_/B _45056_/X _45087_/X _45088_/X sky130_fd_sc_hd__o21a_4
X_77997_ _77997_/A _78012_/A _77998_/A sky130_fd_sc_hd__xor2_4
X_48916_ _48903_/A _48995_/A sky130_fd_sc_hd__buf_2
X_67750_ _87970_/Q _67651_/X _67748_/X _67749_/X _67750_/X sky130_fd_sc_hd__a211o_4
X_44039_ _44038_/X _44039_/X sky130_fd_sc_hd__buf_2
X_79736_ _79720_/X _79724_/B _79736_/X sky130_fd_sc_hd__or2_4
X_64962_ _65984_/A _65111_/B sky130_fd_sc_hd__buf_2
X_76948_ _76953_/A _76953_/B _76948_/Y sky130_fd_sc_hd__nand2_4
X_60085_ _60085_/A _60092_/B sky130_fd_sc_hd__inv_2
X_49896_ _72139_/B _49880_/X _49895_/Y _49896_/Y sky130_fd_sc_hd__o21ai_4
X_66701_ _87374_/Q _66678_/X _66629_/X _66700_/X _66701_/X sky130_fd_sc_hd__a211o_4
X_63913_ _63912_/X _63913_/X sky130_fd_sc_hd__buf_2
X_48847_ _48851_/A _48847_/B _48847_/Y sky130_fd_sc_hd__nand2_4
X_67681_ _67203_/X _67681_/X sky130_fd_sc_hd__buf_2
X_79667_ _79667_/A _79666_/Y _79667_/X sky130_fd_sc_hd__xor2_4
X_64893_ _64694_/A _85814_/Q _64893_/X sky130_fd_sc_hd__and2_4
X_76879_ _81595_/Q _76879_/B _76879_/X sky130_fd_sc_hd__xor2_4
X_69420_ _69300_/X _69340_/X _69417_/Y _69419_/Y _69420_/X sky130_fd_sc_hd__a211o_4
X_66632_ _66627_/X _66631_/X _66606_/X _66632_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_10_508_0_CLK clkbuf_9_254_0_CLK/X _86104_/CLK sky130_fd_sc_hd__clkbuf_1
X_78618_ _78617_/Y _78618_/Y sky130_fd_sc_hd__inv_2
X_63844_ _61399_/X _63877_/B _63814_/C _63877_/D _63844_/Y sky130_fd_sc_hd__nand4_4
X_48778_ _86484_/Q _48754_/X _48777_/Y _48778_/Y sky130_fd_sc_hd__o21ai_4
X_79598_ _79598_/A _81094_/D sky130_fd_sc_hd__inv_2
X_69351_ _68761_/X _68764_/X _69295_/X _69351_/Y sky130_fd_sc_hd__a21oi_4
X_47729_ _81228_/Q _47729_/Y sky130_fd_sc_hd__inv_2
X_66563_ _66563_/A _69567_/A sky130_fd_sc_hd__buf_2
X_78549_ _78549_/A _82675_/D _78554_/A sky130_fd_sc_hd__nor2_4
X_63775_ _63384_/B _63820_/B _63753_/C _64177_/D _63775_/Y sky130_fd_sc_hd__nand4_4
X_60987_ _61012_/C _60918_/X _60987_/Y sky130_fd_sc_hd__nor2_4
X_68302_ _67847_/X _67849_/X _68283_/X _68302_/Y sky130_fd_sc_hd__a21oi_4
X_65514_ _65512_/Y _65448_/X _65513_/X _84196_/D sky130_fd_sc_hd__a21o_4
X_50740_ _50740_/A _53953_/B _50740_/Y sky130_fd_sc_hd__nand2_4
X_62726_ _58241_/X _62689_/X _62708_/X _62699_/X _62725_/X _62726_/Y
+ sky130_fd_sc_hd__a41oi_4
X_81560_ _81433_/CLK _81560_/D _81560_/Q sky130_fd_sc_hd__dfxtp_4
X_69282_ _68629_/X _68632_/X _69212_/X _69282_/Y sky130_fd_sc_hd__a21oi_4
X_66494_ _66475_/X _66275_/Y _66493_/Y _66494_/Y sky130_fd_sc_hd__o21ai_4
X_80511_ _80495_/X _80498_/Y _80510_/X _80511_/X sky130_fd_sc_hd__a21o_4
X_68233_ _68221_/X _67436_/Y _68228_/X _68232_/Y _68233_/X sky130_fd_sc_hd__a211o_4
X_65445_ _64835_/X _83080_/Q _65015_/X _65444_/X _65445_/X sky130_fd_sc_hd__a211o_4
X_50671_ _86156_/Q _50654_/X _50670_/Y _50671_/Y sky130_fd_sc_hd__o21ai_4
X_62657_ _60239_/A _62657_/X sky130_fd_sc_hd__buf_2
X_81491_ _81265_/CLK _84059_/Q _81491_/Q sky130_fd_sc_hd__dfxtp_4
X_52410_ _85828_/Q _52397_/X _52409_/Y _52410_/Y sky130_fd_sc_hd__o21ai_4
X_83230_ _83229_/CLK _72574_/Y _79394_/B sky130_fd_sc_hd__dfxtp_4
X_61608_ _61290_/X _61608_/X sky130_fd_sc_hd__buf_2
X_80442_ _80442_/A _80442_/B _80452_/B sky130_fd_sc_hd__xor2_4
X_68164_ _67038_/X _67042_/X _68129_/X _68164_/Y sky130_fd_sc_hd__a21oi_4
X_53390_ _53386_/A _53390_/B _53390_/Y sky130_fd_sc_hd__nand2_4
X_65376_ _64564_/X _86115_/Q _64566_/X _65375_/X _65376_/X sky130_fd_sc_hd__a211o_4
X_62588_ _61652_/B _62504_/X _62534_/X _62621_/D _62589_/D sky130_fd_sc_hd__nand4_4
X_67115_ _66899_/X _67102_/Y _67031_/X _67114_/Y _67115_/X sky130_fd_sc_hd__a211o_4
X_52341_ _52320_/A _49041_/A _52341_/X sky130_fd_sc_hd__and2_4
X_64327_ _64318_/X _64320_/X _64321_/X _64325_/Y _64326_/X _64327_/X
+ sky130_fd_sc_hd__o41a_4
X_83161_ _83161_/CLK _73192_/X _83161_/Q sky130_fd_sc_hd__dfxtp_4
X_61539_ _61355_/A _61541_/A sky130_fd_sc_hd__buf_2
X_80373_ _80383_/B _80372_/X _80375_/A sky130_fd_sc_hd__xor2_4
X_68095_ _84040_/Q _68040_/X _68094_/X _68095_/X sky130_fd_sc_hd__a21bo_4
X_82112_ _82580_/CLK _82124_/Q _82112_/Q sky130_fd_sc_hd__dfxtp_4
X_55060_ _85326_/Q _55046_/X _55059_/Y _55060_/Y sky130_fd_sc_hd__o21ai_4
X_67046_ _67046_/A _67046_/X sky130_fd_sc_hd__buf_2
X_52272_ _52293_/A _48901_/B _52272_/Y sky130_fd_sc_hd__nand2_4
X_64258_ _64221_/A _64304_/D sky130_fd_sc_hd__buf_2
X_83092_ _83095_/CLK _74339_/X _70326_/A sky130_fd_sc_hd__dfxtp_4
X_54011_ _53998_/A _46417_/B _54011_/Y sky130_fd_sc_hd__nand2_4
X_51223_ _86051_/Q _51209_/X _51222_/Y _51223_/Y sky130_fd_sc_hd__o21ai_4
X_86920_ _86920_/CLK _86920_/D _86920_/Q sky130_fd_sc_hd__dfxtp_4
X_82043_ _82139_/CLK _77958_/B _82043_/Q sky130_fd_sc_hd__dfxtp_4
X_63209_ _63209_/A _63170_/X _63161_/C _63267_/D _63209_/X sky130_fd_sc_hd__or4_4
X_64189_ _84730_/Q _64067_/A _64189_/C _64189_/D _64189_/Y sky130_fd_sc_hd__nand4_4
X_51154_ _51160_/A _51160_/B _51141_/X _52846_/D _51154_/X sky130_fd_sc_hd__and4_4
X_86851_ _86882_/CLK _45838_/Y _63324_/B sky130_fd_sc_hd__dfxtp_4
X_68997_ _68986_/Y _68823_/X _68824_/X _68996_/Y _68997_/X sky130_fd_sc_hd__a211o_4
X_50105_ _50105_/A _50106_/A sky130_fd_sc_hd__buf_2
X_85802_ _85514_/CLK _85802_/D _65209_/B sky130_fd_sc_hd__dfxtp_4
X_58750_ _58763_/A _58750_/B _58750_/Y sky130_fd_sc_hd__nor2_4
X_51085_ _51081_/Y _51065_/X _51084_/X _86077_/D sky130_fd_sc_hd__a21oi_4
X_55962_ _55959_/X _55961_/X _55615_/X _55965_/A sky130_fd_sc_hd__a21o_4
X_67948_ _66898_/X _67948_/X sky130_fd_sc_hd__buf_2
X_86782_ _82317_/CLK _86782_/D _86782_/Q sky130_fd_sc_hd__dfxtp_4
X_83994_ _82642_/CLK _68278_/X _83994_/Q sky130_fd_sc_hd__dfxtp_4
X_57701_ _57701_/A _58635_/A sky130_fd_sc_hd__buf_2
X_50036_ _50050_/A _50040_/B _51750_/C _53249_/D _50036_/X sky130_fd_sc_hd__and4_4
X_54913_ _85354_/Q _54892_/X _54912_/Y _54913_/Y sky130_fd_sc_hd__o21ai_4
X_85733_ _86342_/CLK _85733_/D _85733_/Q sky130_fd_sc_hd__dfxtp_4
X_58681_ _58591_/X _85464_/Q _58680_/X _58681_/Y sky130_fd_sc_hd__o21ai_4
X_82945_ _82369_/CLK _78123_/X _82945_/Q sky130_fd_sc_hd__dfxtp_4
X_55893_ _55892_/X _55928_/A sky130_fd_sc_hd__buf_2
X_67879_ _67997_/A _67879_/X sky130_fd_sc_hd__buf_2
X_57632_ _57608_/X _52079_/B _57632_/Y sky130_fd_sc_hd__nand2_4
X_69618_ _87823_/Q _69619_/B sky130_fd_sc_hd__inv_2
X_54844_ _54842_/Y _54830_/X _54843_/X _85368_/D sky130_fd_sc_hd__a21oi_4
X_85664_ _85439_/CLK _85664_/D _85664_/Q sky130_fd_sc_hd__dfxtp_4
X_70890_ _70863_/A _70890_/B _70890_/C _70890_/D _70890_/Y sky130_fd_sc_hd__nand4_4
X_82876_ _82942_/CLK _78262_/B _82876_/Q sky130_fd_sc_hd__dfxtp_4
X_87403_ _88171_/CLK _43477_/Y _87403_/Q sky130_fd_sc_hd__dfxtp_4
X_84615_ _84477_/CLK _60457_/Y _79155_/A sky130_fd_sc_hd__dfxtp_4
X_57563_ _57563_/A _57563_/X sky130_fd_sc_hd__buf_2
X_81827_ _82211_/CLK _81827_/D _77236_/A sky130_fd_sc_hd__dfxtp_4
X_69549_ _69546_/X _69548_/X _69433_/X _69549_/Y sky130_fd_sc_hd__a21oi_4
X_88383_ _87417_/CLK _40494_/Y _88383_/Q sky130_fd_sc_hd__dfxtp_4
X_54775_ _54775_/A _54788_/B _54775_/C _47502_/A _54775_/X sky130_fd_sc_hd__and4_4
X_85595_ _85590_/CLK _85595_/D _85595_/Q sky130_fd_sc_hd__dfxtp_4
X_51987_ _52486_/A _51987_/X sky130_fd_sc_hd__buf_2
X_59302_ _59237_/X _59299_/Y _59300_/Y _59301_/X _59241_/X _59302_/X
+ sky130_fd_sc_hd__o32a_4
X_56514_ _56103_/X _56499_/X _56513_/Y _56514_/Y sky130_fd_sc_hd__o21ai_4
X_41740_ _41717_/X _81740_/Q _41739_/X _41741_/A sky130_fd_sc_hd__o21ai_4
X_87334_ _87345_/CLK _43632_/Y _87334_/Q sky130_fd_sc_hd__dfxtp_4
X_53726_ _53778_/A _50503_/B _53726_/Y sky130_fd_sc_hd__nand2_4
X_72560_ _72559_/Y _72560_/Y sky130_fd_sc_hd__inv_2
X_84546_ _84529_/CLK _84546_/D _84546_/Q sky130_fd_sc_hd__dfxtp_4
X_50938_ _51021_/A _50938_/X sky130_fd_sc_hd__buf_2
X_57494_ _46366_/A _57499_/A sky130_fd_sc_hd__buf_2
X_81758_ _81783_/CLK _76130_/B _81758_/Q sky130_fd_sc_hd__dfxtp_4
X_59233_ _59231_/X _85422_/Q _59232_/X _59233_/Y sky130_fd_sc_hd__o21ai_4
X_71511_ _53227_/B _71508_/X _71510_/Y _83473_/D sky130_fd_sc_hd__o21ai_4
X_56445_ _56148_/X _56439_/X _56444_/Y _85191_/D sky130_fd_sc_hd__o21ai_4
X_80709_ _80676_/CLK _75895_/X _80709_/Q sky130_fd_sc_hd__dfxtp_4
X_87265_ _88036_/CLK _87265_/D _87265_/Q sky130_fd_sc_hd__dfxtp_4
X_41671_ _44587_/A _41802_/A sky130_fd_sc_hd__buf_2
X_53657_ _85593_/Q _53626_/X _53656_/Y _53657_/Y sky130_fd_sc_hd__o21ai_4
X_72491_ _72484_/X _83383_/Q _72490_/Y _83247_/D sky130_fd_sc_hd__o21a_4
X_84477_ _84477_/CLK _84477_/D _84477_/Q sky130_fd_sc_hd__dfxtp_4
X_50869_ _50867_/Y _50849_/X _50868_/Y _50869_/Y sky130_fd_sc_hd__a21boi_4
X_81689_ _81689_/CLK _80171_/X _76707_/A sky130_fd_sc_hd__dfxtp_4
XPHY_100 sky130_fd_sc_hd__decap_3
X_43410_ _41503_/X _43396_/X _87435_/Q _43397_/X _87435_/D sky130_fd_sc_hd__a2bb2o_4
X_86216_ _85599_/CLK _50361_/Y _86216_/Q sky130_fd_sc_hd__dfxtp_4
X_74230_ _44745_/Y _56274_/X _74229_/Y _74230_/X sky130_fd_sc_hd__a21o_4
X_40622_ _46526_/A _48904_/A sky130_fd_sc_hd__buf_2
XPHY_111 sky130_fd_sc_hd__decap_3
X_52608_ _52624_/A _46676_/A _52608_/Y sky130_fd_sc_hd__nand2_4
X_59164_ _59085_/X _86068_/Q _59163_/X _59164_/Y sky130_fd_sc_hd__o21ai_4
X_83428_ _82386_/CLK _71643_/Y _83428_/Q sky130_fd_sc_hd__dfxtp_4
X_71442_ _71258_/A _71217_/B _71500_/C _71442_/Y sky130_fd_sc_hd__nand3_4
XPHY_122 sky130_fd_sc_hd__decap_3
X_44390_ _41469_/X _44377_/X _87133_/Q _44379_/X _44390_/X sky130_fd_sc_hd__a2bb2o_4
X_56376_ _56372_/X _55987_/X _56375_/Y _85217_/D sky130_fd_sc_hd__o21ai_4
X_87196_ _87446_/CLK _87196_/D _67891_/B sky130_fd_sc_hd__dfxtp_4
X_53588_ _53601_/A _53588_/B _53588_/Y sky130_fd_sc_hd__nand2_4
XPHY_133 sky130_fd_sc_hd__decap_3
XPHY_144 sky130_fd_sc_hd__decap_3
X_58115_ _58111_/Y _58114_/Y _58003_/X _58115_/X sky130_fd_sc_hd__a21o_4
XPHY_155 sky130_fd_sc_hd__decap_3
X_43341_ _41312_/X _43336_/X _87470_/Q _43337_/X _87470_/D sky130_fd_sc_hd__a2bb2o_4
X_55327_ _55322_/X _83750_/Q _55324_/X _55384_/A sky130_fd_sc_hd__nand3_4
X_74161_ _74148_/Y _74161_/B _74161_/Y sky130_fd_sc_hd__xnor2_4
X_86147_ _83594_/CLK _86147_/D _86147_/Q sky130_fd_sc_hd__dfxtp_4
X_40553_ _42446_/A _40636_/A sky130_fd_sc_hd__inv_2
X_52539_ _52501_/X _54058_/B _52539_/Y sky130_fd_sc_hd__nand2_4
XPHY_166 sky130_fd_sc_hd__decap_3
X_59095_ _59027_/X _59093_/Y _59094_/Y _59046_/X _59031_/X _59095_/X
+ sky130_fd_sc_hd__o32a_4
X_71373_ _71372_/Y _71373_/X sky130_fd_sc_hd__buf_2
X_83359_ _83421_/CLK _83359_/D _83359_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_177 sky130_fd_sc_hd__decap_3
XPHY_188 sky130_fd_sc_hd__decap_3
X_73112_ _73181_/A _85876_/Q _73112_/X sky130_fd_sc_hd__and2_4
XPHY_199 sky130_fd_sc_hd__decap_3
X_70324_ _70320_/X _74768_/B _70323_/X _83797_/D sky130_fd_sc_hd__a21o_4
X_46060_ _41555_/Y _46043_/X _86788_/Q _46044_/X _46060_/X sky130_fd_sc_hd__a2bb2o_4
X_58046_ _58042_/Y _58045_/Y _58035_/X _58046_/X sky130_fd_sc_hd__a21o_4
X_43272_ _41121_/X _43264_/X _87506_/Q _43265_/X _87506_/D sky130_fd_sc_hd__a2bb2o_4
X_55258_ _55135_/A _85065_/Q _55258_/X sky130_fd_sc_hd__and2_4
X_86078_ _85757_/CLK _86078_/D _86078_/Q sky130_fd_sc_hd__dfxtp_4
X_74092_ _74079_/Y _74092_/B _74093_/B sky130_fd_sc_hd__xnor2_4
X_40484_ _40325_/X _82318_/Q _40483_/X _40484_/Y sky130_fd_sc_hd__o21ai_4
X_45011_ _45003_/X _45008_/Y _45010_/Y _45011_/Y sky130_fd_sc_hd__a21oi_4
X_42223_ _41909_/Y _42259_/A sky130_fd_sc_hd__buf_2
X_54209_ _54208_/X _54191_/B _54209_/C _53044_/D _54209_/X sky130_fd_sc_hd__and4_4
X_73043_ _72908_/X _85591_/Q _72909_/X _73042_/X _73043_/X sky130_fd_sc_hd__a211o_4
X_77920_ _77920_/A _77919_/Y _77923_/A sky130_fd_sc_hd__xor2_4
X_85029_ _85040_/CLK _85029_/D _85029_/Q sky130_fd_sc_hd__dfxtp_4
X_70255_ _70238_/A _70255_/X sky130_fd_sc_hd__buf_2
X_55189_ _55278_/A _55710_/B sky130_fd_sc_hd__buf_2
X_42154_ _42083_/A _42154_/X sky130_fd_sc_hd__buf_2
X_77851_ _77851_/A _77851_/Y sky130_fd_sc_hd__inv_2
X_70186_ _70232_/A _70200_/B sky130_fd_sc_hd__buf_2
X_59997_ _59995_/X _59950_/B _59977_/B _60091_/B _59998_/B sky130_fd_sc_hd__nand4_4
X_41105_ _41104_/X _41065_/X _69547_/B _41066_/X _88277_/D sky130_fd_sc_hd__a2bb2o_4
X_76802_ _76802_/A _76802_/B _76802_/X sky130_fd_sc_hd__xor2_4
X_49750_ _49641_/A _49750_/X sky130_fd_sc_hd__buf_2
X_46962_ _46961_/X _46981_/A sky130_fd_sc_hd__buf_2
X_42085_ _42084_/Y _42085_/Y sky130_fd_sc_hd__inv_2
X_58948_ _58858_/X _85443_/Q _58947_/X _58948_/Y sky130_fd_sc_hd__o21ai_4
X_77782_ _77782_/A _77782_/Y sky130_fd_sc_hd__inv_2
X_74994_ _81143_/D _75003_/B _74994_/X sky130_fd_sc_hd__xor2_4
X_48701_ _74509_/A _48702_/A sky130_fd_sc_hd__buf_2
X_79521_ _79510_/Y _79512_/B _79519_/A _79522_/B sky130_fd_sc_hd__nand3_4
X_45913_ MACRO_RD_SELECT _59498_/A _45913_/Y sky130_fd_sc_hd__nor2_4
X_41036_ _41035_/X _41036_/X sky130_fd_sc_hd__buf_2
X_76733_ _76733_/A _76733_/B _81547_/D sky130_fd_sc_hd__xor2_4
X_49681_ _49676_/Y _49677_/X _49680_/X _86343_/D sky130_fd_sc_hd__a21oi_4
X_73945_ _73941_/X _73943_/X _73944_/X _73945_/X sky130_fd_sc_hd__a21o_4
X_58879_ _58835_/X _85449_/Q _58878_/X _58879_/Y sky130_fd_sc_hd__o21ai_4
X_46893_ _46941_/A _46896_/B sky130_fd_sc_hd__buf_2
X_60910_ _60909_/X _60910_/B _60910_/X sky130_fd_sc_hd__and2_4
X_48632_ _48632_/A _48632_/B _48632_/Y sky130_fd_sc_hd__nand2_4
X_79452_ _79459_/B _79451_/Y _82843_/D sky130_fd_sc_hd__xnor2_4
X_45844_ _45842_/Y _45632_/X _44884_/X _45843_/Y _45844_/X sky130_fd_sc_hd__a211o_4
X_76664_ _76664_/A _76663_/Y _81443_/D sky130_fd_sc_hd__xnor2_4
X_61890_ _61447_/B _61843_/B _61860_/C _61860_/D _61890_/Y sky130_fd_sc_hd__nand4_4
X_73876_ _68699_/B _73777_/X _73656_/X _73876_/X sky130_fd_sc_hd__o21a_4
X_78403_ _78403_/A _82709_/Q _78408_/C sky130_fd_sc_hd__nand2_4
X_75615_ _75640_/A _75609_/Y _75622_/A _75615_/Y sky130_fd_sc_hd__o21ai_4
X_48563_ _48471_/A _48563_/X sky130_fd_sc_hd__buf_2
X_60841_ _60615_/A _59551_/A _60843_/A sky130_fd_sc_hd__and2_4
X_72827_ _44187_/A _74012_/A sky130_fd_sc_hd__buf_2
X_79383_ _79373_/A _79373_/B _79382_/Y _79387_/A sky130_fd_sc_hd__a21boi_4
X_45775_ _82985_/Q _45388_/X _45774_/X _45775_/Y sky130_fd_sc_hd__o21ai_4
X_76595_ _76595_/A _76595_/B _76595_/Y sky130_fd_sc_hd__nand2_4
X_42987_ _42986_/Y _42987_/Y sky130_fd_sc_hd__inv_2
X_47514_ _47508_/Y _47509_/X _47513_/X _86627_/D sky130_fd_sc_hd__a21oi_4
X_78334_ _78329_/A _78332_/Y _78333_/Y _78334_/Y sky130_fd_sc_hd__o21ai_4
X_44726_ _44707_/X _44708_/X _40712_/A _44725_/Y _44710_/X _44726_/Y
+ sky130_fd_sc_hd__o32ai_4
X_63560_ _58377_/A _63558_/X _61528_/A _63559_/X _63560_/X sky130_fd_sc_hd__a2bb2o_4
X_75546_ _75546_/A _75539_/X _75546_/C _75546_/Y sky130_fd_sc_hd__nand3_4
X_41938_ _41938_/A _41938_/Y sky130_fd_sc_hd__inv_2
X_60772_ _60711_/X _60660_/X _60697_/B _60772_/Y sky130_fd_sc_hd__nand3_4
X_48494_ _73096_/B _48478_/X _48493_/Y _48494_/Y sky130_fd_sc_hd__o21ai_4
X_72758_ _73638_/A _72758_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_494_0_CLK clkbuf_9_247_0_CLK/X _84815_/CLK sky130_fd_sc_hd__clkbuf_1
X_62511_ _62214_/A _62511_/X sky130_fd_sc_hd__buf_2
X_47445_ _86634_/Q _47429_/X _47444_/Y _47445_/Y sky130_fd_sc_hd__o21ai_4
X_71709_ _71691_/Y _83402_/Q _71708_/Y _83402_/D sky130_fd_sc_hd__a21o_4
X_78265_ _78265_/A _82467_/Q _78265_/Y sky130_fd_sc_hd__nand2_4
X_44657_ _44657_/A _44657_/Y sky130_fd_sc_hd__inv_2
X_63491_ _59399_/A _63491_/B _63465_/C _63491_/D _63491_/Y sky130_fd_sc_hd__nand4_4
X_75477_ _75477_/A _75477_/B _75477_/C _75477_/X sky130_fd_sc_hd__or3_4
X_41869_ _41869_/A _41869_/B _41869_/C _41869_/Y sky130_fd_sc_hd__nor3_4
X_72689_ _72697_/A _72697_/B _55405_/X _72689_/Y sky130_fd_sc_hd__nand3_4
XPHY_2 sky130_fd_sc_hd__decap_3
X_65230_ _64772_/A _65230_/X sky130_fd_sc_hd__buf_2
X_77216_ _77217_/A _77217_/B _77216_/Y sky130_fd_sc_hd__nor2_4
X_43608_ _40590_/X _43604_/X _87344_/Q _43607_/X _87344_/D sky130_fd_sc_hd__a2bb2o_4
X_62442_ _62411_/X _62412_/X _62442_/C _62442_/Y sky130_fd_sc_hd__nor3_4
X_74428_ _74413_/X _74428_/B _74428_/Y sky130_fd_sc_hd__nand2_4
X_47376_ _46902_/A _47565_/A sky130_fd_sc_hd__buf_2
X_78196_ _78204_/A _78205_/A _78197_/B sky130_fd_sc_hd__xor2_4
X_44588_ _44679_/A _44588_/X sky130_fd_sc_hd__buf_2
X_49115_ _49115_/A _72072_/B sky130_fd_sc_hd__inv_2
X_46327_ _86747_/Q _46279_/X _46326_/Y _46327_/Y sky130_fd_sc_hd__o21ai_4
X_65161_ _64807_/A _65161_/X sky130_fd_sc_hd__buf_2
X_77147_ _82102_/Q _77147_/B _77147_/X sky130_fd_sc_hd__xor2_4
X_43539_ _43538_/Y _87369_/D sky130_fd_sc_hd__inv_2
X_62373_ _61468_/A _62332_/B _62386_/C _62332_/D _62378_/B sky130_fd_sc_hd__nand4_4
X_74359_ _45954_/X _58334_/A _56167_/B _74359_/Y sky130_fd_sc_hd__nand3_4
X_64112_ _62557_/Y _60880_/X _84913_/Q _61028_/X _64112_/Y sky130_fd_sc_hd__a2bb2oi_4
X_49046_ _49007_/A _50133_/B _49046_/Y sky130_fd_sc_hd__nand2_4
X_61324_ _61323_/X _61324_/Y sky130_fd_sc_hd__inv_2
X_46258_ _46258_/A _46258_/X sky130_fd_sc_hd__buf_2
X_65092_ _65196_/A _65268_/B _84215_/Q _65092_/X sky130_fd_sc_hd__and3_4
X_77078_ _77066_/A _82284_/D _77078_/Y sky130_fd_sc_hd__nand2_4
X_45209_ _45284_/A _45209_/X sky130_fd_sc_hd__buf_2
X_68920_ _68759_/A _68920_/B _68920_/X sky130_fd_sc_hd__and2_4
X_64043_ _60871_/Y _64145_/B sky130_fd_sc_hd__buf_2
X_76029_ _76023_/A _76023_/B _76024_/A _76029_/Y sky130_fd_sc_hd__a21boi_4
X_61255_ _75899_/A _61252_/X _61208_/Y _61254_/Y _61255_/X sky130_fd_sc_hd__o22a_4
X_46189_ _46195_/A _46133_/C _46217_/B _46189_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_432_0_CLK clkbuf_9_216_0_CLK/X _83526_/CLK sky130_fd_sc_hd__clkbuf_1
X_60206_ _60182_/A _61286_/A sky130_fd_sc_hd__buf_2
X_68851_ _87488_/Q _68757_/X _68731_/X _68850_/X _68851_/X sky130_fd_sc_hd__a211o_4
X_61186_ _60933_/X _61110_/Y _61294_/D _59662_/C _61185_/Y _84512_/D
+ sky130_fd_sc_hd__a41oi_4
X_67802_ _86956_/Q _67706_/X _67755_/X _67801_/X _67802_/X sky130_fd_sc_hd__a211o_4
X_60137_ _60028_/Y _60102_/Y _60119_/Y _59988_/Y _60136_/Y _84655_/D
+ sky130_fd_sc_hd__a41oi_4
X_49948_ _49946_/Y _49924_/X _49947_/X _49948_/Y sky130_fd_sc_hd__a21oi_4
X_68782_ _41941_/A _68757_/X _68555_/X _68781_/Y _68782_/X sky130_fd_sc_hd__a211o_4
X_65994_ _65878_/A _73711_/B _65994_/X sky130_fd_sc_hd__and2_4
X_67733_ _86959_/Q _67706_/X _67633_/X _67732_/X _67733_/X sky130_fd_sc_hd__a211o_4
X_79719_ _79712_/X _79719_/B _79719_/Y sky130_fd_sc_hd__nand2_4
X_64945_ _64667_/A _64946_/A sky130_fd_sc_hd__buf_2
X_60068_ _59951_/B _60061_/Y _60000_/A _60129_/B _60067_/Y _84667_/D
+ sky130_fd_sc_hd__a41oi_4
Xclkbuf_10_447_0_CLK clkbuf_9_223_0_CLK/X _85317_/CLK sky130_fd_sc_hd__clkbuf_1
X_49879_ _48897_/A _49906_/A sky130_fd_sc_hd__buf_2
X_80991_ _80991_/CLK _75850_/Y _80991_/Q sky130_fd_sc_hd__dfxtp_4
X_51910_ _51908_/Y _51904_/X _51909_/X _51910_/Y sky130_fd_sc_hd__a21oi_4
X_82730_ _84111_/CLK _84114_/Q _82730_/Q sky130_fd_sc_hd__dfxtp_4
X_67664_ _66898_/X _67664_/X sky130_fd_sc_hd__buf_2
X_52890_ _85735_/Q _52874_/X _52889_/Y _52890_/Y sky130_fd_sc_hd__o21ai_4
X_64876_ _64873_/X _64875_/X _64807_/X _64876_/X sky130_fd_sc_hd__a21o_4
X_69403_ _69400_/X _69402_/X _69403_/Y sky130_fd_sc_hd__nand2_4
X_66615_ _66534_/A _66689_/A sky130_fd_sc_hd__buf_2
X_51841_ _85936_/Q _51817_/X _51840_/Y _51841_/Y sky130_fd_sc_hd__o21ai_4
X_63827_ _63761_/A _63877_/D sky130_fd_sc_hd__buf_2
X_82661_ _82879_/CLK _82661_/D _82661_/Q sky130_fd_sc_hd__dfxtp_4
X_67595_ _67359_/X _67595_/X sky130_fd_sc_hd__buf_2
X_84400_ _84400_/CLK _84400_/D _84400_/Q sky130_fd_sc_hd__dfxtp_4
X_81612_ _81259_/CLK _76297_/B _81612_/Q sky130_fd_sc_hd__dfxtp_4
X_69334_ _69331_/X _69333_/X _69138_/X _69334_/X sky130_fd_sc_hd__a21o_4
X_54560_ _54556_/Y _54558_/X _54559_/X _54560_/Y sky130_fd_sc_hd__a21oi_4
X_66546_ _57776_/A _66547_/A sky130_fd_sc_hd__buf_2
X_85380_ _85379_/CLK _85380_/D _85380_/Q sky130_fd_sc_hd__dfxtp_4
X_51772_ _51768_/A _51782_/B _51755_/X _51772_/D _51772_/X sky130_fd_sc_hd__and4_4
X_63758_ _58221_/X _64189_/C _60908_/A _63731_/D _63758_/Y sky130_fd_sc_hd__nand4_4
X_82592_ _82671_/CLK _82624_/Q _78301_/A sky130_fd_sc_hd__dfxtp_4
X_53511_ _53511_/A _53697_/B sky130_fd_sc_hd__buf_2
X_84331_ _84187_/CLK _63346_/Y _79169_/B sky130_fd_sc_hd__dfxtp_4
X_50723_ _50460_/A _50724_/A sky130_fd_sc_hd__buf_2
X_81543_ _81575_/CLK _81543_/D _76522_/B sky130_fd_sc_hd__dfxtp_4
X_62709_ _62655_/Y _62979_/A sky130_fd_sc_hd__buf_2
X_69265_ _69253_/A _69265_/B _69265_/X sky130_fd_sc_hd__and2_4
X_54491_ _54486_/X _47006_/Y _54491_/Y sky130_fd_sc_hd__nand2_4
X_66477_ _66475_/X _66228_/Y _66476_/Y _66477_/Y sky130_fd_sc_hd__o21ai_4
X_63689_ _63644_/A _63701_/A sky130_fd_sc_hd__buf_2
X_56230_ _56079_/X _56225_/X _56229_/Y _56230_/Y sky130_fd_sc_hd__o21ai_4
X_68216_ _68106_/A _68216_/X sky130_fd_sc_hd__buf_2
X_87050_ _88324_/CLK _44574_/Y _44573_/A sky130_fd_sc_hd__dfxtp_4
X_53442_ _53817_/A _54067_/A sky130_fd_sc_hd__buf_2
X_65428_ _64797_/A _65428_/X sky130_fd_sc_hd__buf_2
X_84262_ _83402_/CLK _64254_/X _79846_/B sky130_fd_sc_hd__dfxtp_4
X_50654_ _50506_/A _50654_/X sky130_fd_sc_hd__buf_2
X_81474_ _81352_/CLK _81474_/D _81474_/Q sky130_fd_sc_hd__dfxtp_4
X_69196_ _69027_/A _88303_/Q _69196_/X sky130_fd_sc_hd__and2_4
X_86001_ _85712_/CLK _86001_/D _86001_/Q sky130_fd_sc_hd__dfxtp_4
X_83213_ _83216_/CLK _72622_/X _79198_/B sky130_fd_sc_hd__dfxtp_4
X_80425_ _80425_/A _80425_/B _80425_/Y sky130_fd_sc_hd__nand2_4
X_68147_ _82067_/D _68140_/X _68146_/X _68147_/X sky130_fd_sc_hd__a21bo_4
X_56161_ _56142_/X _56159_/X _56160_/Y _56161_/Y sky130_fd_sc_hd__o21ai_4
X_53373_ _53353_/A _53373_/B _53373_/Y sky130_fd_sc_hd__nand2_4
X_65359_ _65359_/A _65358_/X _65359_/Y sky130_fd_sc_hd__nand2_4
X_84193_ _84192_/CLK _84193_/D _65559_/C sky130_fd_sc_hd__dfxtp_4
X_50585_ _50583_/Y _50551_/X _50584_/X _50585_/Y sky130_fd_sc_hd__a21oi_4
X_55112_ _55112_/A _47877_/A _55120_/C _47803_/A _55112_/X sky130_fd_sc_hd__and4_4
X_52324_ _52324_/A _52324_/X sky130_fd_sc_hd__buf_2
X_83144_ _83544_/CLK _73594_/X _83144_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_506_0_CLK clkbuf_9_506_0_CLK/A clkbuf_9_506_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_56092_ _56088_/X _56091_/X _55830_/X _56083_/C _56093_/C sky130_fd_sc_hd__a2bb2oi_4
X_80356_ _84752_/Q _84144_/Q _80358_/A sky130_fd_sc_hd__xor2_4
X_68078_ _68403_/A _68078_/B _68078_/X sky130_fd_sc_hd__and2_4
X_55043_ _46614_/X _55043_/X sky130_fd_sc_hd__buf_2
X_59920_ _62475_/A _62515_/C sky130_fd_sc_hd__buf_2
X_67029_ _88384_/Q _66954_/X _66955_/X _67028_/X _67030_/B sky130_fd_sc_hd__a211o_4
X_52255_ _52185_/X _48872_/B _52255_/Y sky130_fd_sc_hd__nand2_4
X_83075_ _86523_/CLK _83075_/D _83075_/Q sky130_fd_sc_hd__dfxtp_4
X_87952_ _87952_/CLK _42263_/Y _87952_/Q sky130_fd_sc_hd__dfxtp_4
X_80287_ _80288_/A _80288_/B _80287_/X sky130_fd_sc_hd__xor2_4
X_51206_ _86054_/Q _51183_/X _51205_/Y _51206_/Y sky130_fd_sc_hd__o21ai_4
X_70040_ _64732_/A _70040_/X sky130_fd_sc_hd__buf_2
X_86903_ _84421_/CLK _45037_/Y _64305_/B sky130_fd_sc_hd__dfxtp_4
X_82026_ _81954_/CLK _77805_/B _81994_/D sky130_fd_sc_hd__dfxtp_4
X_59851_ _60036_/A _59852_/A sky130_fd_sc_hd__buf_2
X_52186_ _52185_/X _48551_/X _52186_/Y sky130_fd_sc_hd__nand2_4
X_87883_ _87883_/CLK _87883_/D _87883_/Q sky130_fd_sc_hd__dfxtp_4
X_58802_ _58748_/X _58800_/Y _58801_/Y _58766_/X _58752_/X _58802_/X
+ sky130_fd_sc_hd__o32a_4
X_51137_ _51160_/A _51121_/B _51115_/C _52831_/D _51137_/X sky130_fd_sc_hd__and4_4
X_86834_ _86834_/CLK _86834_/D _86834_/Q sky130_fd_sc_hd__dfxtp_4
X_59782_ _70056_/A _59782_/X sky130_fd_sc_hd__buf_2
X_56994_ _56726_/X _56684_/B _56739_/X _56994_/D _56994_/Y sky130_fd_sc_hd__nand4_4
X_58733_ _58682_/X _85780_/Q _58706_/X _58733_/X sky130_fd_sc_hd__o21a_4
X_55945_ _55945_/A _55945_/B _55946_/A sky130_fd_sc_hd__and2_4
X_51068_ _51064_/Y _51065_/X _51067_/X _86080_/D sky130_fd_sc_hd__a21oi_4
X_86765_ _84409_/CLK _86765_/D _44904_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_74_0_CLK clkbuf_8_75_0_CLK/A clkbuf_8_74_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_71991_ _72007_/A _53819_/B _71991_/Y sky130_fd_sc_hd__nand2_4
X_83977_ _80740_/CLK _83977_/D _83977_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_6_0_CLK clkbuf_7_6_0_CLK/A clkbuf_7_6_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_42910_ _42909_/Y _42910_/Y sky130_fd_sc_hd__inv_2
X_50019_ _72415_/B _50012_/X _50018_/Y _50019_/Y sky130_fd_sc_hd__o21ai_4
X_85716_ _84757_/CLK _52998_/Y _85716_/Q sky130_fd_sc_hd__dfxtp_4
X_73730_ _44688_/Y _73728_/X _73729_/Y _73730_/X sky130_fd_sc_hd__a21o_4
X_58664_ _58793_/A _58664_/X sky130_fd_sc_hd__buf_2
X_70942_ _70942_/A _70942_/B _70947_/C _70942_/Y sky130_fd_sc_hd__nand3_4
X_82928_ _81190_/CLK _78231_/X _82928_/Q sky130_fd_sc_hd__dfxtp_4
X_43890_ _43862_/X _43876_/X _41316_/X _87213_/Q _43863_/X _43890_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55876_ _55549_/A _55876_/B _55876_/X sky130_fd_sc_hd__and2_4
X_86696_ _86697_/CLK _86696_/D _58887_/A sky130_fd_sc_hd__dfxtp_4
X_57615_ _47714_/A _57615_/X sky130_fd_sc_hd__buf_2
X_42841_ _41503_/X _42830_/X _87691_/Q _42832_/X _42841_/X sky130_fd_sc_hd__a2bb2o_4
X_54827_ _54823_/A _47589_/Y _54827_/Y sky130_fd_sc_hd__nand2_4
X_73661_ _73284_/A _73661_/X sky130_fd_sc_hd__buf_2
X_85647_ _85648_/CLK _53368_/Y _85647_/Q sky130_fd_sc_hd__dfxtp_4
X_70873_ _70873_/A _70869_/B _70869_/C _70869_/D _70873_/Y sky130_fd_sc_hd__nand4_4
X_58595_ _58571_/X _85791_/Q _58594_/X _58595_/X sky130_fd_sc_hd__o21a_4
X_82859_ _82859_/CLK _82483_/Q _40883_/A sky130_fd_sc_hd__dfxtp_4
X_75400_ _75401_/A _75397_/Y _75399_/Y _75400_/X sky130_fd_sc_hd__a21o_4
X_72612_ _72516_/B _72579_/A _59512_/X _72602_/X _72612_/X sky130_fd_sc_hd__a211o_4
X_45560_ _45560_/A _45654_/B _45560_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_89_0_CLK clkbuf_8_89_0_CLK/A clkbuf_8_89_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_57546_ _57528_/X _73864_/A _57546_/Y sky130_fd_sc_hd__nand2_4
X_76380_ _76376_/X _76379_/X _76387_/A sky130_fd_sc_hd__xor2_4
X_88366_ _86982_/CLK _40614_/Y _68498_/B sky130_fd_sc_hd__dfxtp_4
X_42772_ _42739_/X _42740_/X _41316_/X _87725_/Q _42750_/X _42773_/A
+ sky130_fd_sc_hd__o32ai_4
X_54758_ _54758_/A _54758_/X sky130_fd_sc_hd__buf_2
X_85578_ _85859_/CLK _85578_/D _85578_/Q sky130_fd_sc_hd__dfxtp_4
X_73592_ _73582_/Y _73591_/X _73592_/Y sky130_fd_sc_hd__xnor2_4
X_44511_ _40686_/A _44512_/A sky130_fd_sc_hd__buf_2
X_87317_ _83153_/CLK _87317_/D _87317_/Q sky130_fd_sc_hd__dfxtp_4
X_75331_ _80692_/Q _80948_/D _75331_/Y sky130_fd_sc_hd__nor2_4
X_41723_ _41814_/A _41723_/X sky130_fd_sc_hd__buf_2
X_53709_ _53713_/A _48559_/Y _53709_/Y sky130_fd_sc_hd__nand2_4
X_72543_ _72543_/A _72573_/A sky130_fd_sc_hd__buf_2
X_84529_ _84529_/CLK _84529_/D _76977_/A sky130_fd_sc_hd__dfxtp_4
X_45491_ _45488_/Y _45489_/X _45443_/X _45490_/Y _45491_/X sky130_fd_sc_hd__a211o_4
X_57477_ _57372_/X _57474_/Y _57476_/X _57478_/A sky130_fd_sc_hd__o21ai_4
X_88297_ _87022_/CLK _88297_/D _69279_/B sky130_fd_sc_hd__dfxtp_4
X_54689_ _54674_/A _54707_/B _54674_/C _47348_/A _54689_/X sky130_fd_sc_hd__and4_4
X_47230_ _47230_/A _54097_/B sky130_fd_sc_hd__inv_2
X_59216_ _84759_/Q _59216_/Y sky130_fd_sc_hd__inv_2
X_78050_ _84555_/Q _78050_/B _81859_/D sky130_fd_sc_hd__xor2_4
X_44442_ _44441_/Y _87106_/D sky130_fd_sc_hd__inv_2
X_56428_ _56109_/X _56426_/X _56427_/Y _85198_/D sky130_fd_sc_hd__o21ai_4
X_75262_ _75237_/X _75240_/X _75262_/X sky130_fd_sc_hd__xor2_4
X_41654_ _82908_/Q _41653_/X _41654_/X sky130_fd_sc_hd__or2_4
X_87248_ _87766_/CLK _43827_/X _87248_/Q sky130_fd_sc_hd__dfxtp_4
X_72474_ _72465_/Y _72358_/X _72470_/X _72473_/X _72474_/Y sky130_fd_sc_hd__a22oi_4
Xclkbuf_8_12_0_CLK clkbuf_7_6_0_CLK/X clkbuf_9_25_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_77001_ _84553_/Q _84425_/Q _77001_/X sky130_fd_sc_hd__xor2_4
X_74213_ _45931_/X _86213_/Q _72985_/X _74212_/X _74213_/X sky130_fd_sc_hd__a211o_4
X_40605_ _40604_/X _40605_/X sky130_fd_sc_hd__buf_2
X_47161_ _82376_/Q _54580_/D sky130_fd_sc_hd__inv_2
X_71425_ _71420_/X _83504_/Q _71424_/X _71425_/X sky130_fd_sc_hd__a21o_4
X_59147_ _58934_/X _85653_/Q _59081_/X _59147_/X sky130_fd_sc_hd__o21a_4
X_44373_ _41768_/X _44364_/X _87141_/Q _44365_/X _87141_/D sky130_fd_sc_hd__a2bb2o_4
X_56359_ _56153_/X _56350_/X _56358_/Y _85222_/D sky130_fd_sc_hd__o21ai_4
X_87179_ _87178_/CLK _87179_/D _44232_/B sky130_fd_sc_hd__dfxtp_4
X_75193_ _75182_/A _75162_/B _75162_/A _75193_/Y sky130_fd_sc_hd__nand3_4
X_41585_ _41548_/X _82313_/Q _41584_/X _41585_/Y sky130_fd_sc_hd__o21ai_4
X_46112_ _46112_/A _46111_/X _46138_/A sky130_fd_sc_hd__nor2_4
X_43324_ _41264_/X _43300_/X _87480_/Q _43302_/X _87480_/D sky130_fd_sc_hd__a2bb2o_4
X_74144_ _41963_/Y _56273_/X _72725_/A _74143_/Y _74144_/X sky130_fd_sc_hd__a211o_4
X_40536_ _40937_/A _40536_/B _40536_/X sky130_fd_sc_hd__or2_4
X_47092_ _47092_/A _47093_/A sky130_fd_sc_hd__inv_2
X_59078_ _84770_/Q _59078_/Y sky130_fd_sc_hd__inv_2
X_71356_ DATA_TO_HASH[5] _71427_/C sky130_fd_sc_hd__buf_2
X_46043_ _43585_/X _46043_/X sky130_fd_sc_hd__buf_2
X_58029_ _58010_/X _58026_/Y _58027_/Y _58028_/X _58015_/X _58029_/X
+ sky130_fd_sc_hd__o32a_4
X_70307_ _70303_/X _74748_/A _70306_/X _70307_/X sky130_fd_sc_hd__a21o_4
X_43255_ _41070_/X _43247_/X _87515_/Q _43248_/X _87515_/D sky130_fd_sc_hd__a2bb2o_4
X_78952_ _78952_/A _78951_/X _78956_/A sky130_fd_sc_hd__nand2_4
X_74075_ _43087_/Y _72895_/X _73486_/X _74074_/Y _74075_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_8_27_0_CLK clkbuf_8_27_0_CLK/A clkbuf_9_55_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_40467_ _82321_/Q _40467_/B _40467_/X sky130_fd_sc_hd__or2_4
X_71287_ _71136_/A _70696_/B _71287_/C _70578_/A _71287_/Y sky130_fd_sc_hd__nand4_4
X_42206_ _42205_/X _42200_/X _41321_/X _87980_/Q _42201_/X _42206_/Y
+ sky130_fd_sc_hd__o32ai_4
X_61040_ _60995_/Y _61008_/Y _60989_/X _84531_/Q _59509_/X _84531_/D
+ sky130_fd_sc_hd__o32a_4
X_77903_ _77891_/A _77890_/Y _77902_/X _77903_/Y sky130_fd_sc_hd__o21ai_4
X_73026_ _73530_/B _73026_/X sky130_fd_sc_hd__buf_2
X_70238_ _70238_/A _70238_/X sky130_fd_sc_hd__buf_2
X_43186_ _40890_/X _43180_/X _73341_/A _43185_/X _43186_/X sky130_fd_sc_hd__a2bb2o_4
X_78883_ _82635_/Q _78885_/A sky130_fd_sc_hd__inv_2
X_40398_ _82331_/Q _40385_/B _40398_/X sky130_fd_sc_hd__or2_4
X_49802_ _49807_/A _49802_/B _49795_/X _53015_/D _49802_/X sky130_fd_sc_hd__and4_4
X_42137_ _42137_/A _42137_/X sky130_fd_sc_hd__buf_2
X_77834_ _77847_/A _77833_/Y _77842_/A sky130_fd_sc_hd__xor2_4
X_70169_ _70209_/A _70169_/X sky130_fd_sc_hd__buf_2
X_47994_ _47872_/A _52573_/B sky130_fd_sc_hd__buf_2
X_49733_ _49678_/X _49751_/A sky130_fd_sc_hd__buf_2
X_46945_ _46939_/Y _46940_/X _46944_/X _46945_/Y sky130_fd_sc_hd__a21oi_4
X_42068_ _42067_/Y _88049_/D sky130_fd_sc_hd__inv_2
X_77765_ _77764_/B _77756_/Y _77765_/Y sky130_fd_sc_hd__nor2_4
X_62991_ _60259_/A _61694_/B _62926_/B _60281_/A _62186_/X _62991_/X
+ sky130_fd_sc_hd__a32o_4
X_74977_ _74987_/A _74988_/A _74978_/B sky130_fd_sc_hd__xor2_4
X_79504_ _79500_/Y _79504_/B _79510_/B sky130_fd_sc_hd__xor2_4
X_41019_ _82290_/Q _41019_/B _41019_/X sky130_fd_sc_hd__or2_4
X_64730_ _64720_/X _64727_/X _64729_/X _64730_/X sky130_fd_sc_hd__a21o_4
X_76716_ _76714_/Y _76715_/Y _76725_/A sky130_fd_sc_hd__xor2_4
X_49664_ _49651_/X _49642_/B _49669_/C _52879_/D _49664_/X sky130_fd_sc_hd__and4_4
X_61942_ _61929_/X _61932_/X _61941_/Y _84740_/Q _61895_/X _61942_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73928_ _72744_/X _85618_/Q _72857_/X _73927_/X _73928_/X sky130_fd_sc_hd__a211o_4
X_46876_ _46868_/A _46845_/X _46868_/C _52724_/D _46876_/X sky130_fd_sc_hd__and4_4
X_77696_ _77693_/C _77693_/D _77680_/X _77703_/B sky130_fd_sc_hd__a21bo_4
X_48615_ _48615_/A _52216_/B sky130_fd_sc_hd__buf_2
X_79435_ _58653_/A _79435_/B _79444_/A sky130_fd_sc_hd__xor2_4
X_45827_ _85029_/Q _45827_/B _45827_/Y sky130_fd_sc_hd__nor2_4
X_64661_ _64561_/X _64649_/Y _64660_/Y _64661_/Y sky130_fd_sc_hd__o21ai_4
X_76647_ _81682_/Q _81394_/Q _76965_/A sky130_fd_sc_hd__xnor2_4
X_61873_ _61736_/A _61879_/A sky130_fd_sc_hd__buf_2
X_49595_ _86358_/Q _49579_/X _49594_/Y _49595_/Y sky130_fd_sc_hd__o21ai_4
X_73859_ _73614_/A _73859_/X sky130_fd_sc_hd__buf_2
X_66400_ _66262_/A _66402_/B sky130_fd_sc_hd__buf_2
X_63612_ _61568_/B _63609_/X _63610_/X _63611_/Y _63612_/X sky130_fd_sc_hd__a211o_4
X_48546_ _52182_/A _48500_/X _48610_/C _48546_/X sky130_fd_sc_hd__and3_4
X_60824_ _60823_/Y _60824_/Y sky130_fd_sc_hd__inv_2
X_67380_ _67144_/A _67381_/A sky130_fd_sc_hd__buf_2
X_79366_ _79350_/X _79353_/Y _79366_/X sky130_fd_sc_hd__or2_4
X_45758_ _45754_/X _45756_/Y _45757_/X _45758_/X sky130_fd_sc_hd__a21o_4
X_64592_ _64803_/A _64593_/A sky130_fd_sc_hd__buf_2
X_76578_ _76550_/Y _76554_/B _76552_/Y _76578_/X sky130_fd_sc_hd__o21a_4
X_66331_ _84140_/Q _66332_/C sky130_fd_sc_hd__inv_2
X_78317_ _78318_/A _78335_/B _78318_/B _78317_/X sky130_fd_sc_hd__a21o_4
X_44709_ _44709_/A _44709_/Y sky130_fd_sc_hd__inv_2
X_63543_ _63554_/A _63554_/B _80475_/B _63543_/Y sky130_fd_sc_hd__nor3_4
X_75529_ _75528_/B _75530_/A sky130_fd_sc_hd__inv_2
X_48477_ _48470_/Y _48459_/X _48476_/X _48477_/Y sky130_fd_sc_hd__a21oi_4
X_60755_ _60761_/A _60752_/B _60755_/C _60755_/Y sky130_fd_sc_hd__nor3_4
X_79297_ _79297_/A _79296_/Y _82828_/D sky130_fd_sc_hd__xor2_4
X_45689_ _85070_/Q _45801_/A _45689_/Y sky130_fd_sc_hd__nor2_4
X_69050_ _69047_/X _69049_/X _69050_/Y sky130_fd_sc_hd__nand2_4
X_47428_ _47423_/Y _47414_/X _47427_/X _86636_/D sky130_fd_sc_hd__a21oi_4
X_66262_ _66262_/A _66389_/B sky130_fd_sc_hd__buf_2
X_78248_ _78248_/A _78248_/B _78251_/A sky130_fd_sc_hd__nor2_4
X_63474_ _63488_/A _61876_/X _63474_/X sky130_fd_sc_hd__and2_4
X_60686_ _60646_/Y _60677_/A _60713_/A _60686_/X sky130_fd_sc_hd__a21o_4
X_68001_ _87447_/Q _67953_/X _67954_/X _68000_/X _68001_/X sky130_fd_sc_hd__a211o_4
X_65213_ _65159_/A _86026_/Q _65213_/X sky130_fd_sc_hd__and2_4
X_62425_ _62416_/X _62421_/Y _62424_/X _84739_/Q _62367_/X _62425_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47359_ _47359_/A _47360_/A sky130_fd_sc_hd__inv_2
X_66193_ _66177_/A _66164_/B _66193_/C _66193_/Y sky130_fd_sc_hd__nor3_4
X_78179_ _78170_/Y _78177_/Y _78178_/Y _78179_/X sky130_fd_sc_hd__o21a_4
X_80210_ _80197_/Y _80201_/Y _80209_/X _80210_/Y sky130_fd_sc_hd__o21ai_4
X_65144_ _64946_/A _65144_/B _65144_/X sky130_fd_sc_hd__and2_4
X_50370_ _50383_/A _50370_/B _50370_/Y sky130_fd_sc_hd__nand2_4
X_62356_ _62344_/X _57660_/X _62315_/C _62355_/X _62356_/X sky130_fd_sc_hd__and4_4
X_81190_ _81190_/CLK _74927_/X _49161_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_371_0_CLK clkbuf_9_185_0_CLK/X _83049_/CLK sky130_fd_sc_hd__clkbuf_1
X_49029_ _49029_/A _49029_/B _49029_/Y sky130_fd_sc_hd__nor2_4
X_61307_ _61295_/A _72540_/B _72503_/A _61308_/A sky130_fd_sc_hd__o21a_4
X_80141_ _80132_/X _80141_/B _80141_/Y sky130_fd_sc_hd__nand2_4
X_69952_ _69535_/X _69537_/X _69939_/X _69952_/Y sky130_fd_sc_hd__a21oi_4
X_65075_ _64971_/X _86127_/Q _64972_/X _65074_/X _65075_/X sky130_fd_sc_hd__a211o_4
X_62287_ _62304_/A _58237_/X _62244_/C _62286_/X _62287_/X sky130_fd_sc_hd__and4_4
X_52040_ _52037_/Y _51987_/X _52039_/X _85901_/D sky130_fd_sc_hd__a21oi_4
X_68903_ _87082_/Q _68832_/X _68875_/X _68902_/X _68903_/X sky130_fd_sc_hd__a211o_4
X_64026_ _64026_/A _64091_/B sky130_fd_sc_hd__buf_2
X_61238_ _61086_/X _61238_/B _61238_/C _64454_/B _61238_/Y sky130_fd_sc_hd__nand4_4
X_80072_ _80071_/X _80072_/Y sky130_fd_sc_hd__inv_2
X_69883_ _69791_/A _69883_/B _69883_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_9_492_0_CLK clkbuf_9_493_0_CLK/A clkbuf_9_492_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_83900_ _82116_/CLK _83900_/D _83900_/Q sky130_fd_sc_hd__dfxtp_4
X_68834_ _73985_/A _68832_/X _68762_/X _68833_/X _68834_/X sky130_fd_sc_hd__a211o_4
X_61169_ _64225_/B _61169_/X sky130_fd_sc_hd__buf_2
X_84880_ _84849_/CLK _84880_/D _84880_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_386_0_CLK clkbuf_9_193_0_CLK/X _84333_/CLK sky130_fd_sc_hd__clkbuf_1
X_83831_ _83188_/CLK _83831_/D _83831_/Q sky130_fd_sc_hd__dfxtp_4
X_68765_ _68761_/X _68764_/X _68661_/X _68765_/Y sky130_fd_sc_hd__a21oi_4
X_53991_ _53991_/A _46367_/Y _53991_/Y sky130_fd_sc_hd__nand2_4
X_65977_ _65878_/A _65977_/B _65977_/X sky130_fd_sc_hd__and2_4
X_55730_ _55235_/A _55730_/B _55730_/X sky130_fd_sc_hd__and2_4
X_67716_ _68057_/A _68640_/A sky130_fd_sc_hd__buf_2
X_86550_ _85915_/CLK _86550_/D _73833_/B sky130_fd_sc_hd__dfxtp_4
X_52942_ _52922_/A _52954_/B _52926_/X _52942_/D _52942_/X sky130_fd_sc_hd__and4_4
X_64928_ _64777_/A _64929_/A sky130_fd_sc_hd__buf_2
X_83762_ _83476_/CLK _83762_/D _58372_/A sky130_fd_sc_hd__dfxtp_4
X_80974_ _81059_/CLK _75686_/X _75079_/B sky130_fd_sc_hd__dfxtp_4
X_68696_ _73873_/A _68640_/X _68070_/X _68695_/Y _68696_/X sky130_fd_sc_hd__a211o_4
X_85501_ _85499_/CLK _85501_/D _85501_/Q sky130_fd_sc_hd__dfxtp_4
X_82713_ _82803_/CLK _82713_/D _82669_/D sky130_fd_sc_hd__dfxtp_4
X_67647_ _67696_/A _67647_/B _67647_/X sky130_fd_sc_hd__and2_4
X_55661_ _55652_/Y _55654_/X _55660_/Y _55661_/X sky130_fd_sc_hd__o21a_4
X_86481_ _86191_/CLK _86481_/D _86481_/Q sky130_fd_sc_hd__dfxtp_4
X_52873_ _52870_/Y _52865_/X _52872_/X _52873_/Y sky130_fd_sc_hd__a21oi_4
X_64859_ _64679_/A _64859_/X sky130_fd_sc_hd__buf_2
X_83693_ _82381_/CLK _83693_/D _47183_/A sky130_fd_sc_hd__dfxtp_4
X_57400_ _44308_/X _57400_/X sky130_fd_sc_hd__buf_2
X_88220_ _88220_/CLK _41410_/Y _88220_/Q sky130_fd_sc_hd__dfxtp_4
X_54612_ _54589_/X _54607_/B _54591_/C _54612_/D _54612_/X sky130_fd_sc_hd__and4_4
X_85432_ _85431_/CLK _85432_/D _85432_/Q sky130_fd_sc_hd__dfxtp_4
X_51824_ _51805_/A _51815_/B _51810_/C _46744_/X _51824_/X sky130_fd_sc_hd__and4_4
X_58380_ _58380_/A _58369_/X _58380_/Y sky130_fd_sc_hd__nand2_4
X_82644_ _82642_/CLK _82644_/D _78966_/A sky130_fd_sc_hd__dfxtp_4
X_55592_ _55592_/A _55592_/B _55592_/X sky130_fd_sc_hd__and2_4
X_67578_ _67222_/A _67675_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_430_0_CLK clkbuf_9_430_0_CLK/A clkbuf_9_430_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_57331_ _57331_/A _57331_/B _57331_/C _57331_/Y sky130_fd_sc_hd__nand3_4
X_69317_ _88038_/Q _69315_/X _69245_/X _69316_/X _69317_/X sky130_fd_sc_hd__a211o_4
X_88151_ _88215_/CLK _88151_/D _88151_/Q sky130_fd_sc_hd__dfxtp_4
X_54543_ _85423_/Q _54540_/X _54542_/Y _54543_/Y sky130_fd_sc_hd__o21ai_4
X_66529_ _69315_/A _66529_/X sky130_fd_sc_hd__buf_2
X_85363_ _83630_/CLK _54870_/Y _85363_/Q sky130_fd_sc_hd__dfxtp_4
X_51755_ _51781_/A _51755_/X sky130_fd_sc_hd__buf_2
X_82575_ _82575_/CLK _82607_/Q _78177_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_324_0_CLK clkbuf_9_162_0_CLK/X _83690_/CLK sky130_fd_sc_hd__clkbuf_1
X_87102_ _88272_/CLK _44455_/X _87102_/Q sky130_fd_sc_hd__dfxtp_4
X_84314_ _84314_/CLK _63555_/Y _63554_/C sky130_fd_sc_hd__dfxtp_4
X_50706_ _50742_/A _50706_/X sky130_fd_sc_hd__buf_2
X_57262_ _57261_/X _56639_/X _45600_/A _57236_/X _57262_/X sky130_fd_sc_hd__a2bb2o_4
X_81526_ _84079_/CLK _81526_/D _81526_/Q sky130_fd_sc_hd__dfxtp_4
X_69248_ _68517_/A _69248_/X sky130_fd_sc_hd__buf_2
X_88082_ _88081_/CLK _41985_/Y _88082_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_954_0_CLK clkbuf_9_477_0_CLK/X _87820_/CLK sky130_fd_sc_hd__clkbuf_1
X_54474_ _85435_/Q _54457_/X _54473_/Y _54474_/Y sky130_fd_sc_hd__o21ai_4
X_85294_ _85192_/CLK _56111_/Y _55817_/B sky130_fd_sc_hd__dfxtp_4
X_51686_ _51697_/A _53209_/B _51686_/Y sky130_fd_sc_hd__nand2_4
X_59001_ _59061_/A _59001_/X sky130_fd_sc_hd__buf_2
X_56213_ _56252_/A _56214_/A sky130_fd_sc_hd__buf_2
X_87033_ _88301_/CLK _44612_/X _87033_/Q sky130_fd_sc_hd__dfxtp_4
X_53425_ _53423_/Y _53408_/X _53424_/X _53425_/Y sky130_fd_sc_hd__a21oi_4
X_84245_ _82436_/CLK _64453_/X _84245_/Q sky130_fd_sc_hd__dfxtp_4
X_50637_ _86162_/Q _50626_/X _50636_/Y _50637_/Y sky130_fd_sc_hd__o21ai_4
X_57193_ _56761_/X _56659_/Y _56894_/Y _57193_/D _57193_/Y sky130_fd_sc_hd__nand4_4
X_81457_ _81333_/CLK _76790_/B _81425_/D sky130_fd_sc_hd__dfxtp_4
X_69179_ _69179_/A _69179_/B _69179_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_445_0_CLK clkbuf_9_444_0_CLK/A clkbuf_9_445_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
Xpsn_inst_psn_buff_3 _44267_/A _44266_/C sky130_fd_sc_hd__buf_2
X_71210_ _71225_/A _71219_/C sky130_fd_sc_hd__buf_2
X_56144_ _56144_/A _56144_/X sky130_fd_sc_hd__buf_2
X_80408_ _80386_/Y _80404_/X _80407_/Y _80408_/Y sky130_fd_sc_hd__a21oi_4
X_53356_ _53221_/A _53357_/A sky130_fd_sc_hd__buf_2
X_41370_ _41324_/X _82897_/Q _41369_/X _41370_/Y sky130_fd_sc_hd__o21ai_4
X_72190_ _72172_/X _72187_/Y _72188_/Y _72189_/X _72176_/X _72190_/X
+ sky130_fd_sc_hd__o32a_4
X_84176_ _84175_/CLK _84176_/D _65817_/C sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_339_0_CLK clkbuf_9_169_0_CLK/X _83699_/CLK sky130_fd_sc_hd__clkbuf_1
X_50568_ _48894_/A _50560_/X _50568_/C _50568_/X sky130_fd_sc_hd__and3_4
X_81388_ _81482_/CLK _81388_/D _76884_/B sky130_fd_sc_hd__dfxtp_4
X_52307_ _52299_/A _52307_/B _52307_/Y sky130_fd_sc_hd__nand2_4
X_40321_ _40321_/A _46526_/A sky130_fd_sc_hd__buf_2
X_71141_ _71168_/A _71141_/B _71152_/C _70875_/X _71141_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_10_969_0_CLK clkbuf_9_484_0_CLK/X _86222_/CLK sky130_fd_sc_hd__clkbuf_1
X_83127_ _83145_/CLK _74004_/Y _83127_/Q sky130_fd_sc_hd__dfxtp_4
X_80339_ _80337_/Y _80338_/Y _80339_/X sky130_fd_sc_hd__xor2_4
X_56075_ _56104_/A _56100_/A sky130_fd_sc_hd__buf_2
X_53287_ _85661_/Q _53268_/X _53286_/Y _53287_/Y sky130_fd_sc_hd__o21ai_4
X_50499_ _50594_/A _50499_/X sky130_fd_sc_hd__buf_2
X_43040_ _43040_/A _87598_/D sky130_fd_sc_hd__inv_2
X_55026_ _55017_/X _55026_/B _55026_/C _55026_/D _55026_/X sky130_fd_sc_hd__and4_4
X_59903_ _59903_/A _59904_/B sky130_fd_sc_hd__inv_2
X_52238_ _52236_/Y _52232_/X _52237_/X _85862_/D sky130_fd_sc_hd__a21oi_4
X_71072_ _71072_/A _71078_/C sky130_fd_sc_hd__buf_2
X_83058_ _85571_/CLK _74479_/Y _83058_/Q sky130_fd_sc_hd__dfxtp_4
X_87935_ _88386_/CLK _42295_/Y _87935_/Q sky130_fd_sc_hd__dfxtp_4
X_74900_ _74900_/A _74900_/Y sky130_fd_sc_hd__inv_2
X_70023_ _69712_/X _69714_/X _70001_/X _70023_/Y sky130_fd_sc_hd__a21oi_4
X_82009_ _82009_/CLK _82041_/Q _77163_/A sky130_fd_sc_hd__dfxtp_4
X_59834_ _59834_/A _59833_/X _80400_/A _59834_/X sky130_fd_sc_hd__or3_4
X_52169_ _85875_/Q _52152_/X _52168_/Y _52169_/Y sky130_fd_sc_hd__o21ai_4
X_75880_ _75880_/A _75880_/B _75880_/Y sky130_fd_sc_hd__nand2_4
X_87866_ _82899_/CLK _87866_/D _87866_/Q sky130_fd_sc_hd__dfxtp_4
X_86817_ _86784_/CLK _86817_/D _67071_/B sky130_fd_sc_hd__dfxtp_4
X_74831_ _74831_/A _74844_/A sky130_fd_sc_hd__buf_2
X_59765_ _59765_/A _61770_/B sky130_fd_sc_hd__buf_2
X_44991_ _44988_/X _44990_/Y _44973_/X _44991_/Y sky130_fd_sc_hd__a21oi_4
X_56977_ _56976_/X _56685_/X _56977_/Y sky130_fd_sc_hd__nor2_4
X_87797_ _87285_/CLK _87797_/D _73507_/A sky130_fd_sc_hd__dfxtp_4
X_46730_ _46724_/Y _46704_/X _46729_/X _86710_/D sky130_fd_sc_hd__a21oi_4
X_58716_ _58847_/A _58716_/X sky130_fd_sc_hd__buf_2
X_77550_ _77551_/A _82116_/Q _77553_/B sky130_fd_sc_hd__nor2_4
X_43942_ _41454_/X _43939_/X _68071_/B _43941_/X _43942_/X sky130_fd_sc_hd__a2bb2o_4
X_55928_ _55928_/A _55928_/B _55928_/C _55927_/X _55956_/A sky130_fd_sc_hd__and4_4
X_74762_ _74762_/A _71507_/B _74762_/Y sky130_fd_sc_hd__nor2_4
X_86748_ _86246_/CLK _46323_/Y _86748_/Q sky130_fd_sc_hd__dfxtp_4
X_71974_ _71970_/A _71974_/B _71974_/Y sky130_fd_sc_hd__nand2_4
X_59696_ _59696_/A _66514_/B _80605_/A _59696_/Y sky130_fd_sc_hd__nor3_4
X_76501_ _81658_/Q _76501_/Y sky130_fd_sc_hd__inv_2
X_73713_ _73708_/X _73712_/X _73612_/X _73716_/A sky130_fd_sc_hd__a21o_4
Xclkbuf_10_907_0_CLK clkbuf_9_453_0_CLK/X _88111_/CLK sky130_fd_sc_hd__clkbuf_1
X_70925_ _70925_/A _70925_/X sky130_fd_sc_hd__buf_2
X_46661_ _83684_/Q _46662_/A sky130_fd_sc_hd__inv_2
X_58647_ _58643_/Y _58645_/Y _58646_/X _58647_/X sky130_fd_sc_hd__a21o_4
X_77481_ _77478_/X _77480_/Y _77481_/Y sky130_fd_sc_hd__nand2_4
X_43873_ _41264_/X _43868_/X _69033_/B _43870_/X _43873_/X sky130_fd_sc_hd__a2bb2o_4
X_55859_ _55856_/X _55858_/X _55516_/X _55859_/X sky130_fd_sc_hd__a21o_4
X_86679_ _86359_/CLK _47022_/Y _59118_/A sky130_fd_sc_hd__dfxtp_4
X_74693_ _74693_/A _74693_/Y sky130_fd_sc_hd__inv_2
X_48400_ _74383_/B _48401_/B sky130_fd_sc_hd__buf_2
X_79220_ _79203_/A _79201_/Y _79219_/Y _79220_/Y sky130_fd_sc_hd__a21oi_4
X_45612_ _45612_/A _45793_/B sky130_fd_sc_hd__buf_2
X_76432_ _76430_/X _76431_/Y _76432_/X sky130_fd_sc_hd__and2_4
X_42824_ _41454_/X _42821_/X _68067_/B _42822_/X _42824_/X sky130_fd_sc_hd__a2bb2o_4
X_49380_ _49397_/A _49369_/X _49380_/C _51768_/D _49380_/X sky130_fd_sc_hd__and4_4
X_73644_ _47863_/Y _73644_/B _73644_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_5_24_0_CLK clkbuf_4_12_1_CLK/X clkbuf_6_49_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_46592_ _57497_/A _54087_/B _46592_/Y sky130_fd_sc_hd__nand2_4
X_58578_ _58079_/X _58576_/Y _58577_/Y _58098_/X _58083_/X _58578_/X
+ sky130_fd_sc_hd__o32a_4
X_70856_ _70854_/A _71068_/B sky130_fd_sc_hd__inv_2
X_48331_ _48328_/Y _48322_/X _48330_/Y _86534_/D sky130_fd_sc_hd__a21boi_4
X_79151_ _79151_/A _79151_/B _79151_/X sky130_fd_sc_hd__xor2_4
X_45543_ _45541_/Y _45542_/Y _44939_/B _45543_/X sky130_fd_sc_hd__o21a_4
X_57529_ _57528_/X _73765_/A _57529_/Y sky130_fd_sc_hd__nand2_4
X_76363_ _81360_/Q _76363_/B _76363_/X sky130_fd_sc_hd__xor2_4
X_88349_ _82538_/CLK _40713_/X _88349_/Q sky130_fd_sc_hd__dfxtp_4
X_42755_ _41264_/X _42745_/X _69031_/B _42746_/X _87736_/D sky130_fd_sc_hd__a2bb2o_4
X_73575_ _88114_/Q _74095_/B _73575_/Y sky130_fd_sc_hd__nor2_4
X_70787_ _70873_/A _70791_/B _70791_/C _70791_/D _70787_/Y sky130_fd_sc_hd__nand4_4
X_78102_ _82566_/Q _78102_/B _78130_/A sky130_fd_sc_hd__xor2_4
X_75314_ _80691_/Q _80991_/Q _75314_/Y sky130_fd_sc_hd__nor2_4
X_41706_ _41672_/X _41673_/X _41705_/X _67683_/B _41668_/X _41707_/A
+ sky130_fd_sc_hd__o32ai_4
X_48262_ _48260_/Y _48233_/X _48261_/X _86546_/D sky130_fd_sc_hd__a21oi_4
X_60540_ _60482_/Y _60541_/C sky130_fd_sc_hd__buf_2
X_72526_ _72522_/Y _72525_/Y _59980_/X _72533_/A sky130_fd_sc_hd__a21o_4
X_79082_ _82623_/D _79082_/B _79084_/A sky130_fd_sc_hd__nand2_4
X_45474_ _85020_/Q _45474_/Y sky130_fd_sc_hd__inv_2
X_76294_ _76283_/A _76267_/B _76293_/A _76294_/Y sky130_fd_sc_hd__a21oi_4
X_42686_ _42685_/Y _87770_/D sky130_fd_sc_hd__inv_2
X_47213_ _47212_/Y _52918_/B sky130_fd_sc_hd__buf_2
X_78033_ _78033_/A _78033_/B _78033_/Y sky130_fd_sc_hd__nand2_4
X_44425_ _44381_/A _44425_/X sky130_fd_sc_hd__buf_2
X_75245_ _75245_/A _75244_/Y _75245_/Y sky130_fd_sc_hd__nand2_4
X_41637_ _40717_/X _41799_/A sky130_fd_sc_hd__buf_2
X_48193_ _48934_/A _48193_/X sky130_fd_sc_hd__buf_2
X_60471_ _63347_/C _60476_/C _60570_/B _60476_/A _60435_/C _60471_/X
+ sky130_fd_sc_hd__o41a_4
X_72457_ _57709_/X _85348_/Q _72456_/X _72457_/Y sky130_fd_sc_hd__o21ai_4
X_62210_ _60084_/A _62211_/D sky130_fd_sc_hd__buf_2
X_47144_ _47138_/Y _47128_/X _47143_/X _86666_/D sky130_fd_sc_hd__a21oi_4
X_71408_ _71191_/A _71411_/B sky130_fd_sc_hd__buf_2
X_44356_ _41715_/X _44345_/X _87151_/Q _44346_/X _87151_/D sky130_fd_sc_hd__a2bb2o_4
X_75176_ _75154_/Y _75151_/Y _75153_/A _75178_/C sky130_fd_sc_hd__o21ai_4
X_63190_ _63010_/A _63190_/X sky130_fd_sc_hd__buf_2
X_41568_ _81164_/Q _41584_/B _41568_/X sky130_fd_sc_hd__or2_4
X_72388_ _72305_/X _85355_/Q _72387_/X _72388_/Y sky130_fd_sc_hd__o21ai_4
X_43307_ _43306_/Y _87489_/D sky130_fd_sc_hd__inv_2
X_74127_ _73583_/A _74127_/B _74127_/X sky130_fd_sc_hd__and2_4
X_62141_ _62140_/X _62175_/B _62046_/C _62046_/D _62141_/Y sky130_fd_sc_hd__nand4_4
X_40519_ _40504_/X _82312_/Q _40518_/X _40519_/Y sky130_fd_sc_hd__o21ai_4
X_47075_ _47067_/A _47039_/B _47048_/C _52841_/D _47075_/X sky130_fd_sc_hd__and4_4
X_71339_ _50389_/B _71320_/A _71338_/Y _71339_/Y sky130_fd_sc_hd__o21ai_4
X_44287_ _44286_/Y _44287_/X sky130_fd_sc_hd__buf_2
X_79984_ _84656_/Q _64130_/C _79985_/B sky130_fd_sc_hd__xor2_4
X_41499_ _41489_/X _41490_/X _41498_/X _66752_/B _41474_/X _41500_/A
+ sky130_fd_sc_hd__o32ai_4
X_46026_ _40547_/Y _46022_/X _86807_/Q _46023_/X _46026_/X sky130_fd_sc_hd__a2bb2o_4
X_43238_ _43237_/Y _43238_/Y sky130_fd_sc_hd__inv_2
X_62072_ _63630_/A _59825_/B _61597_/A _59807_/A _62072_/X sky130_fd_sc_hd__a2bb2o_4
X_74058_ _74038_/A _66209_/B _74058_/X sky130_fd_sc_hd__and2_4
X_78935_ _78921_/Y _78923_/B _82638_/Q _82510_/D _78935_/X sky130_fd_sc_hd__a2bb2o_4
X_65900_ _65969_/A _65916_/A sky130_fd_sc_hd__buf_2
X_61023_ _61022_/Y _60994_/A _61012_/C _76985_/A _59829_/X _84537_/D
+ sky130_fd_sc_hd__a32o_4
X_73009_ _44539_/Y _73006_/X _73008_/Y _73021_/C sky130_fd_sc_hd__a21o_4
X_43169_ _43169_/A _87551_/D sky130_fd_sc_hd__inv_2
X_66880_ _66785_/A _86793_/Q _66880_/X sky130_fd_sc_hd__and2_4
X_78866_ _78866_/A _78860_/Y _78867_/B sky130_fd_sc_hd__nor2_4
X_65831_ _65855_/A _65916_/B _84175_/Q _65831_/X sky130_fd_sc_hd__and3_4
X_77817_ _77817_/A _77816_/X _77822_/A sky130_fd_sc_hd__nand2_4
X_47977_ _83771_/Q _47978_/A sky130_fd_sc_hd__inv_2
X_78797_ _78797_/A _78797_/B _82785_/D sky130_fd_sc_hd__nand2_4
X_49716_ _49688_/X _49716_/X sky130_fd_sc_hd__buf_2
X_68550_ _87096_/Q _68353_/X _68354_/X _68549_/X _68551_/B sky130_fd_sc_hd__a211o_4
X_46928_ _46928_/A _54446_/B sky130_fd_sc_hd__inv_2
X_65762_ _64903_/A _65763_/A sky130_fd_sc_hd__buf_2
X_77748_ _77747_/B _82260_/Q _77751_/C sky130_fd_sc_hd__nand2_4
X_62974_ _61675_/B _62936_/X _62982_/C _62908_/X _62974_/Y sky130_fd_sc_hd__nand4_4
X_67501_ _87404_/Q _67476_/X _67477_/X _67500_/X _67501_/X sky130_fd_sc_hd__a211o_4
X_64713_ _64713_/A _64752_/A sky130_fd_sc_hd__buf_2
X_49647_ _49645_/Y _49623_/X _49646_/X _49647_/Y sky130_fd_sc_hd__a21oi_4
X_61925_ _61879_/A _61919_/Y _61921_/Y _61924_/Y _61925_/Y sky130_fd_sc_hd__nand4_4
X_68481_ _88015_/Q _68402_/X _68359_/X _68480_/X _68481_/X sky130_fd_sc_hd__a211o_4
X_46859_ _46767_/A _46859_/X sky130_fd_sc_hd__buf_2
X_65693_ _65596_/X _83064_/Q _65540_/X _65692_/X _65694_/B sky130_fd_sc_hd__a211o_4
X_77679_ _77678_/X _77679_/Y sky130_fd_sc_hd__inv_2
X_67432_ _66953_/X _67432_/X sky130_fd_sc_hd__buf_2
X_79418_ _79418_/A _79418_/B _79418_/X sky130_fd_sc_hd__and2_4
X_64644_ _64615_/X _85535_/Q _64642_/X _64643_/X _64644_/X sky130_fd_sc_hd__a211o_4
X_49578_ _49575_/Y _49570_/X _49577_/X _49578_/Y sky130_fd_sc_hd__a21oi_4
X_61856_ _61856_/A _61874_/D sky130_fd_sc_hd__buf_2
X_80690_ _80696_/CLK _80690_/D _80690_/Q sky130_fd_sc_hd__dfxtp_4
X_60807_ _60792_/A _60810_/B _84562_/Q _60807_/Y sky130_fd_sc_hd__nor3_4
X_48529_ _81778_/Q _48529_/Y sky130_fd_sc_hd__inv_2
X_67363_ _67357_/X _67362_/X _67264_/X _67367_/A sky130_fd_sc_hd__a21o_4
X_79349_ _79342_/X _79344_/B _79349_/Y sky130_fd_sc_hd__nand2_4
X_64575_ _64570_/X _64573_/X _64574_/X _64582_/A sky130_fd_sc_hd__a21o_4
X_61787_ _61755_/A _61787_/X sky130_fd_sc_hd__buf_2
X_69102_ _69097_/X _69101_/X _69035_/X _69102_/X sky130_fd_sc_hd__a21o_4
X_66314_ _66117_/X _84965_/Q _66118_/X _66313_/X _66314_/X sky130_fd_sc_hd__a211o_4
X_51540_ _51622_/A _51545_/A sky130_fd_sc_hd__buf_2
X_63526_ _59411_/A _63491_/B _63514_/C _63491_/D _63526_/Y sky130_fd_sc_hd__nand4_4
X_82360_ _82570_/CLK _77214_/X _82360_/Q sky130_fd_sc_hd__dfxtp_4
X_60738_ _60624_/A _60687_/A _60632_/X _60738_/Y sky130_fd_sc_hd__nand3_4
X_67294_ _67248_/A _67294_/B _67294_/X sky130_fd_sc_hd__and2_4
X_81311_ _81279_/CLK _76999_/X _81311_/Q sky130_fd_sc_hd__dfxtp_4
X_69033_ _69011_/A _69033_/B _69033_/X sky130_fd_sc_hd__and2_4
X_66245_ _65781_/X _66135_/B _65784_/X _66245_/Y sky130_fd_sc_hd__nand3_4
X_51471_ _51033_/A _51552_/A sky130_fd_sc_hd__buf_2
X_63457_ _63454_/Y _63455_/X _63456_/Y _84322_/D sky130_fd_sc_hd__a21oi_4
X_82291_ _82103_/CLK _77127_/B _41014_/A sky130_fd_sc_hd__dfxtp_4
X_60669_ _60770_/A _63398_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_122_0_CLK clkbuf_6_61_0_CLK/X clkbuf_8_245_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_53210_ _85676_/Q _53198_/X _53209_/Y _53210_/Y sky130_fd_sc_hd__o21ai_4
X_84030_ _81154_/CLK _68136_/X _82070_/D sky130_fd_sc_hd__dfxtp_4
X_50422_ _50420_/Y _50380_/X _50421_/Y _50422_/Y sky130_fd_sc_hd__a21boi_4
X_62408_ _62337_/A _61939_/X _62364_/X _62392_/D _62408_/X sky130_fd_sc_hd__and4_4
X_81242_ _85338_/CLK _81050_/Q _81242_/Q sky130_fd_sc_hd__dfxtp_4
X_54190_ _54217_/A _54191_/B sky130_fd_sc_hd__buf_2
X_66176_ _84151_/Q _66177_/C sky130_fd_sc_hd__inv_2
X_63388_ _61354_/B _60834_/X _63386_/X _63387_/X _63388_/X sky130_fd_sc_hd__a211o_4
X_53141_ _53121_/X _53141_/B _53141_/Y sky130_fd_sc_hd__nand2_4
X_65127_ _64776_/A _65127_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_92_0_CLK clkbuf_9_46_0_CLK/X _84414_/CLK sky130_fd_sc_hd__clkbuf_1
X_50353_ _50350_/Y _50351_/X _50352_/Y _50353_/Y sky130_fd_sc_hd__a21boi_4
X_62339_ _62330_/X _62335_/Y _62338_/X _84745_/Q _62300_/X _62339_/Y
+ sky130_fd_sc_hd__o32ai_4
X_81173_ _82335_/CLK _74985_/B _81173_/Q sky130_fd_sc_hd__dfxtp_4
Xpsn_inst_psn_buff_10 _44196_/D _56278_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_21 _53441_/A _43019_/B1 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_32 _47002_/A _40352_/A sky130_fd_sc_hd__buf_2
X_80124_ _84669_/Q _63944_/C _80124_/X sky130_fd_sc_hd__xor2_4
X_53072_ _53080_/A _53072_/B _53072_/Y sky130_fd_sc_hd__nand2_4
X_65058_ _65009_/X _86160_/Q _64902_/X _65057_/X _65058_/X sky130_fd_sc_hd__a211o_4
X_69935_ _69900_/A _69935_/B _69935_/X sky130_fd_sc_hd__and2_4
X_50284_ _50500_/A _50285_/A sky130_fd_sc_hd__buf_2
X_85981_ _85981_/CLK _85981_/D _85981_/Q sky130_fd_sc_hd__dfxtp_4
X_56900_ _56866_/A _56899_/Y _56900_/X sky130_fd_sc_hd__and2_4
X_52023_ _52274_/A _52431_/A sky130_fd_sc_hd__buf_2
X_64009_ _64074_/A _64074_/B _80082_/B _64009_/Y sky130_fd_sc_hd__nor3_4
X_87720_ _87720_/CLK _87720_/D _87720_/Q sky130_fd_sc_hd__dfxtp_4
X_84932_ _84930_/CLK _84932_/D _84932_/Q sky130_fd_sc_hd__dfxtp_4
X_80055_ _80052_/Y _80035_/Y _80054_/X _80056_/B sky130_fd_sc_hd__o21ai_4
X_57880_ _57838_/X _86007_/Q _57879_/X _57880_/Y sky130_fd_sc_hd__o21ai_4
X_69866_ _87049_/Q _66608_/X _58827_/A _69865_/X _69866_/X sky130_fd_sc_hd__a211o_4
X_56831_ _55264_/A _55264_/C _56831_/X sky130_fd_sc_hd__and2_4
X_68817_ _68814_/X _68816_/X _68773_/X _68817_/X sky130_fd_sc_hd__a21o_4
X_87651_ _87394_/CLK _87651_/D _67714_/B sky130_fd_sc_hd__dfxtp_4
X_84863_ _84344_/CLK _84863_/D _58382_/A sky130_fd_sc_hd__dfxtp_4
X_69797_ _69797_/A _69797_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_253_0_CLK clkbuf_8_253_0_CLK/A clkbuf_9_506_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_86602_ _85961_/CLK _86602_/D _86602_/Q sky130_fd_sc_hd__dfxtp_4
X_59550_ _59564_/A _59516_/A _59581_/C _59551_/A sky130_fd_sc_hd__nand3_4
X_83814_ _83842_/CLK _70276_/X _74781_/A sky130_fd_sc_hd__dfxtp_4
X_56762_ _56733_/X _57003_/B sky130_fd_sc_hd__buf_2
X_68748_ _69678_/A _68748_/X sky130_fd_sc_hd__buf_2
X_87582_ _88327_/CLK _87582_/D _74053_/A sky130_fd_sc_hd__dfxtp_4
X_53974_ _53978_/A _52454_/B _53974_/Y sky130_fd_sc_hd__nand2_4
X_84794_ _86701_/CLK _84794_/D _84794_/Q sky130_fd_sc_hd__dfxtp_4
X_58501_ _64307_/C _63459_/B sky130_fd_sc_hd__buf_2
X_55713_ _55235_/A _55713_/B _55713_/X sky130_fd_sc_hd__and2_4
X_86533_ _86203_/CLK _48339_/Y _86533_/Q sky130_fd_sc_hd__dfxtp_4
X_52925_ _85729_/Q _52902_/X _52924_/Y _52925_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_30_0_CLK clkbuf_9_15_0_CLK/X _82979_/CLK sky130_fd_sc_hd__clkbuf_1
X_59481_ _64225_/C _63369_/B sky130_fd_sc_hd__buf_2
X_83745_ _83745_/CLK _83745_/D _47297_/A sky130_fd_sc_hd__dfxtp_4
X_56693_ _72765_/A _56672_/Y _56693_/C _56694_/C sky130_fd_sc_hd__nand3_4
X_68679_ _68599_/A _87751_/Q _68679_/X sky130_fd_sc_hd__and2_4
X_80957_ _81197_/CLK _75475_/B _75045_/A sky130_fd_sc_hd__dfxtp_4
X_70710_ _70710_/A _70703_/X _70710_/C _70710_/D _70710_/Y sky130_fd_sc_hd__nand4_4
X_58432_ _84849_/Q _63198_/A sky130_fd_sc_hd__inv_2
X_55644_ _55644_/A _56564_/D sky130_fd_sc_hd__buf_2
X_86464_ _83311_/CLK _48895_/Y _86464_/Q sky130_fd_sc_hd__dfxtp_4
X_52856_ _85742_/Q _52848_/X _52855_/Y _52856_/Y sky130_fd_sc_hd__o21ai_4
X_40870_ _40835_/A _40870_/X sky130_fd_sc_hd__buf_2
X_71690_ _71690_/A _71319_/B _71690_/Y sky130_fd_sc_hd__nor2_4
X_83676_ _83676_/CLK _70874_/Y _83676_/Q sky130_fd_sc_hd__dfxtp_4
X_80888_ _80991_/CLK _80888_/D _80888_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_263_0_CLK clkbuf_9_131_0_CLK/X _83763_/CLK sky130_fd_sc_hd__clkbuf_1
X_88203_ _87126_/CLK _88203_/D _88203_/Q sky130_fd_sc_hd__dfxtp_4
X_85415_ _85735_/CLK _54586_/Y _85415_/Q sky130_fd_sc_hd__dfxtp_4
X_51807_ _51796_/A _51807_/B _51807_/Y sky130_fd_sc_hd__nand2_4
X_70641_ _70773_/A _70925_/A sky130_fd_sc_hd__buf_2
X_82627_ _87421_/CLK _83979_/Q _82627_/Q sky130_fd_sc_hd__dfxtp_4
X_58363_ _63335_/A _58364_/A sky130_fd_sc_hd__buf_2
X_55575_ _44064_/X _45474_/Y _55575_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_893_0_CLK clkbuf_9_446_0_CLK/X _85822_/CLK sky130_fd_sc_hd__clkbuf_1
X_86395_ _86393_/CLK _86395_/D _86395_/Q sky130_fd_sc_hd__dfxtp_4
X_52787_ _52773_/A _52787_/B _52787_/Y sky130_fd_sc_hd__nand2_4
X_57314_ _56797_/A _57327_/B _56796_/Y _57315_/A sky130_fd_sc_hd__nand3_4
Xclkbuf_10_45_0_CLK clkbuf_9_22_0_CLK/X _85013_/CLK sky130_fd_sc_hd__clkbuf_1
X_88134_ _88133_/CLK _88134_/D _66892_/B sky130_fd_sc_hd__dfxtp_4
X_42540_ _42612_/A _42540_/X sky130_fd_sc_hd__buf_2
X_54526_ _54509_/A _54526_/B _54509_/C _54526_/D _54526_/X sky130_fd_sc_hd__and4_4
X_73360_ _73407_/A _86506_/Q _73360_/X sky130_fd_sc_hd__and2_4
X_85346_ _85346_/CLK _85346_/D _85346_/Q sky130_fd_sc_hd__dfxtp_4
X_51738_ _85954_/Q _50220_/X _51737_/Y _51738_/Y sky130_fd_sc_hd__o21ai_4
X_58294_ _83405_/Q _58294_/Y sky130_fd_sc_hd__inv_2
X_70572_ _71012_/A _70573_/B sky130_fd_sc_hd__buf_2
X_82558_ _82558_/CLK _82558_/D _82558_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_384_0_CLK clkbuf_8_192_0_CLK/X clkbuf_9_384_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_72311_ _72307_/Y _72310_/Y _72201_/X _72311_/X sky130_fd_sc_hd__a21o_4
X_57245_ _57244_/X _57245_/X sky130_fd_sc_hd__buf_2
X_81509_ _84087_/CLK _81553_/Q _81509_/Q sky130_fd_sc_hd__dfxtp_4
X_88065_ _87553_/CLK _88065_/D _73225_/A sky130_fd_sc_hd__dfxtp_4
X_54457_ _54376_/A _54457_/X sky130_fd_sc_hd__buf_2
X_42471_ _42470_/Y _87854_/D sky130_fd_sc_hd__inv_2
X_73291_ _48582_/A _73290_/Y _73291_/X sky130_fd_sc_hd__xor2_4
X_85277_ _85277_/CLK _85277_/D _56203_/C sky130_fd_sc_hd__dfxtp_4
X_51669_ _51657_/X _51684_/B _51684_/C _53191_/D _51669_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_278_0_CLK clkbuf_9_139_0_CLK/X _85404_/CLK sky130_fd_sc_hd__clkbuf_1
X_82489_ _82711_/CLK _82489_/D _82489_/Q sky130_fd_sc_hd__dfxtp_4
X_44210_ _44158_/Y _44210_/X sky130_fd_sc_hd__buf_2
X_75030_ _75030_/A _75023_/A _75047_/B sky130_fd_sc_hd__and2_4
X_87016_ _87011_/CLK _44652_/X _87016_/Q sky130_fd_sc_hd__dfxtp_4
X_41422_ _41422_/A _41379_/X _41422_/X sky130_fd_sc_hd__or2_4
X_53408_ _53355_/A _53408_/X sky130_fd_sc_hd__buf_2
X_72242_ _72240_/X _85687_/Q _72241_/X _72242_/X sky130_fd_sc_hd__o21a_4
X_84228_ _84228_/CLK _84228_/D _84228_/Q sky130_fd_sc_hd__dfxtp_4
X_45190_ _55814_/B _45134_/X _45189_/X _45190_/X sky130_fd_sc_hd__o21a_4
X_57176_ _57175_/Y _85068_/D sky130_fd_sc_hd__inv_2
X_54388_ _54378_/A _52696_/B _54388_/Y sky130_fd_sc_hd__nand2_4
X_44141_ _44140_/X _44141_/X sky130_fd_sc_hd__buf_2
X_56127_ _56147_/A _56127_/B _56127_/C _56143_/B sky130_fd_sc_hd__nor3_4
X_41353_ _41352_/X _41307_/X _88231_/Q _41308_/X _41353_/X sky130_fd_sc_hd__a2bb2o_4
X_53339_ _53339_/A _53330_/B _53330_/C _52827_/D _53339_/X sky130_fd_sc_hd__and4_4
X_72173_ _59238_/A _72220_/A sky130_fd_sc_hd__buf_2
X_84159_ _84166_/CLK _66067_/X _84159_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_399_0_CLK clkbuf_9_398_0_CLK/A clkbuf_9_399_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_8_206_0_CLK clkbuf_8_207_0_CLK/A clkbuf_9_413_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_201_0_CLK clkbuf_9_100_0_CLK/X _81048_/CLK sky130_fd_sc_hd__clkbuf_1
X_71124_ _49144_/X _71117_/X _71123_/Y _83599_/D sky130_fd_sc_hd__o21ai_4
X_44072_ _44072_/A _44072_/Y sky130_fd_sc_hd__inv_2
X_56058_ _56142_/A _56058_/X sky130_fd_sc_hd__buf_2
X_41284_ _41253_/A _41284_/X sky130_fd_sc_hd__buf_2
X_76981_ _76981_/A _76981_/B _76981_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_10_831_0_CLK clkbuf_9_415_0_CLK/X _86578_/CLK sky130_fd_sc_hd__clkbuf_1
X_47900_ _73717_/A _50264_/B sky130_fd_sc_hd__buf_2
X_43023_ _43023_/A _87603_/D sky130_fd_sc_hd__inv_2
X_55009_ _55013_/A _55026_/B _55013_/C _47616_/A _55009_/X sky130_fd_sc_hd__and4_4
X_78720_ _78720_/A _78721_/B sky130_fd_sc_hd__inv_2
X_71055_ _71055_/A _71055_/B _71055_/C _71055_/Y sky130_fd_sc_hd__nand3_4
X_75932_ _75932_/A _75933_/B sky130_fd_sc_hd__inv_2
X_87918_ _88171_/CLK _87918_/D _87918_/Q sky130_fd_sc_hd__dfxtp_4
X_48880_ _48651_/A _48880_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_322_0_CLK clkbuf_9_323_0_CLK/A clkbuf_9_322_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_70006_ _68559_/X _68561_/X _70005_/X _70006_/Y sky130_fd_sc_hd__a21oi_4
X_47831_ _47830_/Y _57489_/B sky130_fd_sc_hd__buf_2
X_59817_ _59754_/C _59631_/B _61202_/A _62183_/A _59840_/A _59817_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_78651_ _78628_/Y _78632_/B _78630_/Y _78651_/X sky130_fd_sc_hd__o21a_4
X_75863_ _75864_/A _75862_/Y _81024_/Q _75863_/Y sky130_fd_sc_hd__a21oi_4
X_87849_ _87851_/CLK _87849_/D _73795_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_216_0_CLK clkbuf_9_108_0_CLK/X _84520_/CLK sky130_fd_sc_hd__clkbuf_1
X_77602_ _77601_/Y _77603_/C sky130_fd_sc_hd__inv_2
X_74814_ _46220_/A _80668_/D sky130_fd_sc_hd__inv_2
X_47762_ _83472_/Q _47762_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_846_0_CLK clkbuf_9_423_0_CLK/X _86118_/CLK sky130_fd_sc_hd__clkbuf_1
X_59748_ _59742_/Y _59744_/Y _59745_/X _59746_/Y _59747_/Y _59748_/Y
+ sky130_fd_sc_hd__a41oi_4
X_78582_ _78582_/A _82772_/D _82484_/D sky130_fd_sc_hd__xor2_4
X_44974_ _44965_/X _44970_/Y _44973_/X _44974_/Y sky130_fd_sc_hd__a21oi_4
X_75794_ _81018_/Q _80890_/D _80986_/D sky130_fd_sc_hd__xor2_4
X_49501_ _49499_/Y _49487_/X _49500_/X _86376_/D sky130_fd_sc_hd__a21oi_4
X_46713_ _58688_/A _46672_/X _46712_/Y _46713_/Y sky130_fd_sc_hd__o21ai_4
X_77533_ _77532_/A _82103_/D _77533_/Y sky130_fd_sc_hd__nand2_4
X_43925_ _43916_/X _43924_/X _41408_/X _67891_/B _43917_/X _43926_/A
+ sky130_fd_sc_hd__o32ai_4
X_74745_ _74745_/A _74804_/C _74744_/X _74745_/D _74745_/Y sky130_fd_sc_hd__nand4_4
X_47693_ _47689_/Y _47651_/X _47692_/X _86608_/D sky130_fd_sc_hd__a21oi_4
X_71957_ _71957_/A _48876_/Y _71957_/Y sky130_fd_sc_hd__nand2_4
X_59679_ _59679_/A _59687_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_337_0_CLK clkbuf_8_168_0_CLK/X clkbuf_9_337_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_49432_ _86388_/Q _49415_/X _49431_/Y _49432_/Y sky130_fd_sc_hd__o21ai_4
X_61710_ _84729_/Q _59761_/A _62187_/C _59761_/B _61710_/Y sky130_fd_sc_hd__nand4_4
X_46644_ _58601_/A _46622_/X _46643_/Y _46644_/Y sky130_fd_sc_hd__o21ai_4
X_70908_ _70908_/A _70698_/A _70909_/A sky130_fd_sc_hd__nor2_4
X_77464_ _77460_/Y _77439_/Y _77463_/X _77465_/B sky130_fd_sc_hd__o21ai_4
X_43856_ _43855_/Y _43856_/Y sky130_fd_sc_hd__inv_2
X_74676_ _74679_/A _45728_/A _74676_/Y sky130_fd_sc_hd__nand2_4
X_62690_ _62658_/A _64248_/C _62676_/C _62657_/X _62690_/X sky130_fd_sc_hd__and4_4
X_71888_ _71870_/Y _83339_/Q _71887_/Y _83339_/D sky130_fd_sc_hd__a21o_4
X_79203_ _79203_/A _79201_/Y _79202_/Y _79205_/B sky130_fd_sc_hd__nand3_4
X_76415_ _76415_/A _76415_/Y sky130_fd_sc_hd__inv_2
X_42807_ _42806_/Y _87709_/D sky130_fd_sc_hd__inv_2
X_49363_ _86401_/Q _49360_/X _49362_/Y _49363_/Y sky130_fd_sc_hd__o21ai_4
X_61641_ _84871_/Q _61321_/Y _61642_/A sky130_fd_sc_hd__or2_4
X_73627_ _72892_/B _73627_/X sky130_fd_sc_hd__buf_2
X_46575_ _86724_/Q _46543_/X _46574_/Y _46575_/Y sky130_fd_sc_hd__o21ai_4
X_70839_ _70867_/A _70846_/B _70849_/C _70841_/D _70839_/Y sky130_fd_sc_hd__nand4_4
X_77395_ _77417_/A _77417_/B _77434_/B sky130_fd_sc_hd__xnor2_4
X_43787_ _43787_/A _87268_/D sky130_fd_sc_hd__inv_2
X_40999_ _40999_/A _40999_/X sky130_fd_sc_hd__buf_2
X_48314_ _48311_/Y _48273_/X _48313_/Y _48314_/Y sky130_fd_sc_hd__a21boi_4
X_79134_ _79134_/A _79134_/B _79134_/X sky130_fd_sc_hd__xor2_4
X_45526_ _45526_/A _45527_/A sky130_fd_sc_hd__inv_2
X_64360_ _59411_/A _64316_/B _64360_/Y sky130_fd_sc_hd__nor2_4
X_76346_ _76345_/A _81564_/Q _76347_/A sky130_fd_sc_hd__nand2_4
X_42738_ _42737_/Y _87743_/D sky130_fd_sc_hd__inv_2
X_49294_ _49292_/Y _49281_/X _49293_/X _86416_/D sky130_fd_sc_hd__a21oi_4
X_61572_ _61572_/A _61542_/B _61542_/C _61572_/D _61572_/Y sky130_fd_sc_hd__nand4_4
X_73558_ _87007_/Q _57092_/X _73557_/X _73558_/Y sky130_fd_sc_hd__o21ai_4
X_63311_ _59433_/Y _63259_/X _63234_/X _58978_/Y _63235_/X _63311_/Y
+ sky130_fd_sc_hd__o32ai_4
X_60523_ _60523_/A _60523_/X sky130_fd_sc_hd__buf_2
X_48245_ _66087_/B _48241_/X _48244_/Y _48245_/Y sky130_fd_sc_hd__o21ai_4
X_72509_ _72503_/A _72510_/C sky130_fd_sc_hd__buf_2
X_79065_ _79065_/A _79065_/Y sky130_fd_sc_hd__inv_2
X_45457_ _85117_/Q _45456_/X _45457_/Y sky130_fd_sc_hd__nor2_4
X_64291_ _79817_/B _64255_/X _64290_/X _64291_/X sky130_fd_sc_hd__a21o_4
X_76277_ _76276_/B _81643_/Q _76282_/C sky130_fd_sc_hd__nand2_4
X_42669_ _41028_/X _42652_/X _69354_/B _42653_/X _87779_/D sky130_fd_sc_hd__a2bb2o_4
X_73489_ _72861_/X _73489_/X sky130_fd_sc_hd__buf_2
X_66030_ _66030_/A _66029_/X _66030_/Y sky130_fd_sc_hd__nand2_4
X_78016_ _78011_/Y _77993_/B _78015_/Y _78018_/B sky130_fd_sc_hd__o21ai_4
X_44408_ _44407_/Y _87124_/D sky130_fd_sc_hd__inv_2
X_63242_ _63018_/X _63242_/X sky130_fd_sc_hd__buf_2
X_75228_ _75224_/Y _75225_/Y _75227_/Y _75228_/X sky130_fd_sc_hd__or3_4
X_48176_ _48903_/A _49173_/A sky130_fd_sc_hd__buf_2
X_60454_ _60454_/A _60562_/B sky130_fd_sc_hd__buf_2
X_45388_ _45596_/A _45388_/X sky130_fd_sc_hd__buf_2
X_47127_ _46653_/A _47128_/A sky130_fd_sc_hd__buf_2
X_44339_ _44339_/A _87159_/D sky130_fd_sc_hd__inv_2
X_63173_ _63169_/Y _63171_/X _63172_/X _63173_/Y sky130_fd_sc_hd__a21oi_4
X_75159_ _75158_/Y _75138_/Y _75140_/Y _75159_/Y sky130_fd_sc_hd__o21ai_4
X_60385_ _60385_/A _60182_/A _60386_/A sky130_fd_sc_hd__nor2_4
X_62124_ _61948_/A _62124_/B _61755_/X _61728_/A _62124_/X sky130_fd_sc_hd__and4_4
X_47058_ _54522_/D _52831_/D sky130_fd_sc_hd__buf_2
X_67981_ _67978_/X _67981_/B _67981_/Y sky130_fd_sc_hd__nand2_4
X_79967_ _79966_/X _79967_/Y sky130_fd_sc_hd__inv_2
X_46009_ _40496_/Y _46007_/X _67071_/B _46008_/X _86817_/D sky130_fd_sc_hd__a2bb2o_4
X_69720_ _73081_/A _68636_/X _68691_/X _69719_/Y _69720_/X sky130_fd_sc_hd__a211o_4
X_66932_ _66956_/A _66932_/B _66932_/X sky130_fd_sc_hd__and2_4
X_62055_ _62055_/A _62055_/B _59628_/A _59649_/A _62055_/X sky130_fd_sc_hd__and4_4
X_78918_ _78914_/Y _78918_/B _78918_/Y sky130_fd_sc_hd__nand2_4
X_79898_ _60153_/C _64200_/C _79898_/Y sky130_fd_sc_hd__nand2_4
X_61006_ _63734_/A _63765_/A sky130_fd_sc_hd__buf_2
X_69651_ _69651_/A _69680_/A sky130_fd_sc_hd__buf_2
X_66863_ _66628_/X _66863_/X sky130_fd_sc_hd__buf_2
X_78849_ _78874_/A _78854_/B _78856_/A _78849_/Y sky130_fd_sc_hd__o21ai_4
X_68602_ _44020_/A _69357_/A sky130_fd_sc_hd__buf_2
X_65814_ _65810_/X _65725_/B _65813_/X _65814_/Y sky130_fd_sc_hd__nand3_4
X_81860_ _81859_/CLK _78051_/X _81828_/D sky130_fd_sc_hd__dfxtp_4
X_69582_ _69582_/A _69582_/X sky130_fd_sc_hd__buf_2
X_66794_ _66794_/A _66794_/X sky130_fd_sc_hd__buf_2
X_80811_ _83957_/CLK _83955_/Q _75796_/B sky130_fd_sc_hd__dfxtp_4
X_68533_ _64584_/X _69014_/A sky130_fd_sc_hd__buf_2
X_65745_ _65888_/A _65802_/B _65745_/C _65745_/Y sky130_fd_sc_hd__nor3_4
X_50971_ _50971_/A _50971_/B _50971_/Y sky130_fd_sc_hd__nand2_4
X_62957_ _62965_/A _62664_/B _62140_/X _62957_/Y sky130_fd_sc_hd__nand3_4
X_81791_ _86807_/CLK _75950_/X _48384_/A sky130_fd_sc_hd__dfxtp_4
X_52710_ _52707_/Y _52702_/X _52709_/X _52710_/Y sky130_fd_sc_hd__a21oi_4
X_83530_ _86210_/CLK _71339_/Y _48152_/A sky130_fd_sc_hd__dfxtp_4
X_61908_ _61460_/B _61843_/B _61860_/C _61860_/D _61908_/Y sky130_fd_sc_hd__nand4_4
X_80742_ _81996_/CLK _80742_/D _81150_/D sky130_fd_sc_hd__dfxtp_4
X_68464_ _87855_/Q _68465_/B sky130_fd_sc_hd__inv_2
X_53690_ _85587_/Q _53687_/X _53689_/Y _53690_/Y sky130_fd_sc_hd__o21ai_4
X_65676_ _65676_/A _65675_/X _65676_/Y sky130_fd_sc_hd__nand2_4
X_62888_ _62965_/A _62935_/B _63610_/B _62888_/Y sky130_fd_sc_hd__nand3_4
X_67415_ _67342_/A _67415_/B _67415_/X sky130_fd_sc_hd__and2_4
X_52641_ _52637_/A _54332_/B _52641_/Y sky130_fd_sc_hd__nand2_4
X_64627_ _64680_/A _64627_/B _64627_/X sky130_fd_sc_hd__and2_4
X_83461_ _83464_/CLK _83461_/D _83461_/Q sky130_fd_sc_hd__dfxtp_4
X_61839_ _61839_/A _61839_/B _61839_/C _63089_/B _61839_/X sky130_fd_sc_hd__and4_4
X_80673_ _81807_/CLK _70157_/X _80673_/Q sky130_fd_sc_hd__dfxtp_4
X_68395_ _64584_/X _69651_/A sky130_fd_sc_hd__buf_2
X_85200_ _85297_/CLK _85200_/D _56420_/C sky130_fd_sc_hd__dfxtp_4
X_82412_ _82248_/CLK _82444_/Q _78455_/A sky130_fd_sc_hd__dfxtp_4
X_55360_ _55360_/A _55360_/X sky130_fd_sc_hd__buf_2
X_67346_ _87411_/Q _67274_/X _67344_/X _67345_/X _67346_/X sky130_fd_sc_hd__a211o_4
X_86180_ _85859_/CLK _86180_/D _86180_/Q sky130_fd_sc_hd__dfxtp_4
X_52572_ _65411_/B _52516_/X _52571_/Y _52572_/Y sky130_fd_sc_hd__o21ai_4
X_64558_ _64552_/Y _64555_/Y _64557_/Y _84866_/Q _64521_/X _64558_/Y
+ sky130_fd_sc_hd__o32ai_4
X_83392_ _85505_/CLK _83392_/D _47230_/A sky130_fd_sc_hd__dfxtp_4
XPHY_507 sky130_fd_sc_hd__decap_3
XPHY_518 sky130_fd_sc_hd__decap_3
X_54311_ _54366_/A _54311_/X sky130_fd_sc_hd__buf_2
XPHY_529 sky130_fd_sc_hd__decap_3
X_85131_ _85071_/CLK _85131_/D _85131_/Q sky130_fd_sc_hd__dfxtp_4
X_51523_ _51519_/Y _51503_/X _51522_/X _51523_/Y sky130_fd_sc_hd__a21oi_4
X_63509_ _63496_/A _58520_/A _63458_/X _63496_/D _63509_/X sky130_fd_sc_hd__and4_4
X_82343_ _82343_/CLK _77089_/X _48110_/A sky130_fd_sc_hd__dfxtp_4
X_55291_ _55263_/X _55290_/Y _55264_/Y _55291_/Y sky130_fd_sc_hd__a21boi_4
X_67277_ _67273_/X _67276_/X _67204_/X _67277_/X sky130_fd_sc_hd__a21o_4
X_64489_ _64483_/X _64486_/Y _64488_/Y _84873_/Q _64213_/X _64489_/Y
+ sky130_fd_sc_hd__o32ai_4
X_57030_ _56930_/X _57028_/Y _57029_/Y _57031_/A sky130_fd_sc_hd__o21ai_4
X_69016_ _87077_/Q _68948_/X _68993_/X _69015_/X _69016_/X sky130_fd_sc_hd__a211o_4
X_54242_ _54240_/Y _54226_/X _54241_/X _85478_/D sky130_fd_sc_hd__a21oi_4
X_66228_ _66224_/X _66227_/X _66228_/Y sky130_fd_sc_hd__nand2_4
X_85062_ _84998_/CLK _85062_/D _57210_/B sky130_fd_sc_hd__dfxtp_4
X_51454_ _51430_/X _52979_/B _51454_/Y sky130_fd_sc_hd__nand2_4
X_82274_ _82103_/CLK _82274_/D _82274_/Q sky130_fd_sc_hd__dfxtp_4
X_84013_ _84074_/CLK _68203_/X _82053_/D sky130_fd_sc_hd__dfxtp_4
X_50405_ _50432_/A _48380_/X _50405_/Y sky130_fd_sc_hd__nand2_4
X_81225_ _81224_/CLK _81033_/Q _81225_/Q sky130_fd_sc_hd__dfxtp_4
X_54173_ _54160_/A _54186_/B _54191_/C _53003_/D _54173_/X sky130_fd_sc_hd__and4_4
X_66159_ _57770_/A _66159_/B _66159_/X sky130_fd_sc_hd__and2_4
X_51385_ _51383_/Y _51366_/X _51384_/X _86020_/D sky130_fd_sc_hd__a21oi_4
X_53124_ _53097_/X _53133_/B sky130_fd_sc_hd__buf_2
X_50336_ _86221_/Q _50333_/X _50335_/Y _50336_/Y sky130_fd_sc_hd__o21ai_4
X_81156_ _81179_/CLK _81156_/D _40536_/B sky130_fd_sc_hd__dfxtp_4
X_58981_ _58981_/A _58982_/A sky130_fd_sc_hd__buf_2
X_80107_ _80107_/A _80106_/Y _81683_/D sky130_fd_sc_hd__xnor2_4
X_53055_ _85705_/Q _53038_/X _53054_/Y _53055_/Y sky130_fd_sc_hd__o21ai_4
X_57932_ _57781_/X _57930_/Y _57931_/Y _57893_/X _57795_/X _57932_/X
+ sky130_fd_sc_hd__o32a_4
X_69918_ _64615_/A _69918_/B _69918_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_7_52_0_CLK clkbuf_6_26_0_CLK/X clkbuf_7_52_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_50267_ _50265_/Y _50227_/X _50266_/Y _86235_/D sky130_fd_sc_hd__a21boi_4
X_85964_ _85962_/CLK _85964_/D _85964_/Q sky130_fd_sc_hd__dfxtp_4
X_81087_ _81087_/CLK _75688_/A _81087_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_192_0_CLK clkbuf_7_96_0_CLK/X clkbuf_8_192_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_52006_ _73901_/B _51994_/X _52005_/Y _52006_/Y sky130_fd_sc_hd__o21ai_4
X_87703_ _87221_/CLK _87703_/D _87703_/Q sky130_fd_sc_hd__dfxtp_4
X_80038_ _80026_/X _80027_/X _80037_/Y _80042_/A sky130_fd_sc_hd__a21boi_4
X_84915_ _84915_/CLK _84915_/D _84915_/Q sky130_fd_sc_hd__dfxtp_4
X_57863_ _57838_/X _86008_/Q _57862_/X _57863_/Y sky130_fd_sc_hd__o21ai_4
X_69849_ _43170_/A _66529_/X _68436_/X _69848_/X _69849_/X sky130_fd_sc_hd__a211o_4
X_50198_ _50196_/Y _50191_/X _50197_/X _50198_/Y sky130_fd_sc_hd__a21oi_4
X_85895_ _85895_/CLK _85895_/D _66283_/B sky130_fd_sc_hd__dfxtp_4
X_59602_ _59602_/A _59639_/A _59602_/C _59603_/A sky130_fd_sc_hd__and3_4
X_56814_ _56814_/A _56798_/B _56814_/Y sky130_fd_sc_hd__nand2_4
X_87634_ _87995_/CLK _42953_/X _66598_/B sky130_fd_sc_hd__dfxtp_4
X_72860_ _69622_/B _44128_/X _72858_/X _72859_/Y _72860_/X sky130_fd_sc_hd__a211o_4
X_84846_ _83457_/CLK _58447_/X _84846_/Q sky130_fd_sc_hd__dfxtp_4
X_57794_ _58635_/A _72417_/A sky130_fd_sc_hd__buf_2
X_71811_ _71813_/A _71427_/C _70852_/C _71811_/X sky130_fd_sc_hd__and3_4
Xclkbuf_7_67_0_CLK clkbuf_7_67_0_CLK/A clkbuf_7_67_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_59533_ _59899_/B _59899_/D _43969_/A _43969_/B _59546_/A sky130_fd_sc_hd__a22oi_4
X_56745_ _56742_/Y _56744_/Y _56696_/B _56745_/X sky130_fd_sc_hd__a21o_4
X_87565_ _83158_/CLK _43132_/Y _87565_/Q sky130_fd_sc_hd__dfxtp_4
X_53957_ _53956_/X _52440_/B _53957_/Y sky130_fd_sc_hd__nand2_4
X_41971_ _41960_/X _41951_/X _40743_/X _74204_/A _41953_/X _41972_/A
+ sky130_fd_sc_hd__o32ai_4
X_72791_ _72789_/X _72774_/X _72791_/C _72791_/Y sky130_fd_sc_hd__nand3_4
X_84777_ _86372_/CLK _84777_/D _84777_/Q sky130_fd_sc_hd__dfxtp_4
X_81989_ _81989_/CLK _81989_/D _77018_/A sky130_fd_sc_hd__dfxtp_4
X_43710_ _87299_/Q _69780_/B sky130_fd_sc_hd__inv_2
X_74530_ _51130_/B _74516_/X _74529_/Y _74530_/Y sky130_fd_sc_hd__o21ai_4
X_86516_ _86516_/CLK _86516_/D _86516_/Q sky130_fd_sc_hd__dfxtp_4
X_40922_ _40921_/X _40904_/X _88310_/Q _40905_/X _88310_/D sky130_fd_sc_hd__a2bb2o_4
X_52908_ _52895_/A _52916_/B _52900_/C _51214_/D _52908_/X sky130_fd_sc_hd__and4_4
X_71742_ _52924_/B _71737_/X _71741_/Y _71742_/Y sky130_fd_sc_hd__o21ai_4
X_83728_ _85484_/CLK _70674_/X _47458_/A sky130_fd_sc_hd__dfxtp_4
X_59464_ _59398_/A _59478_/B sky130_fd_sc_hd__buf_2
X_44690_ _44686_/X _44687_/X _40625_/Y _44688_/Y _44689_/X _87000_/D
+ sky130_fd_sc_hd__o32ai_4
X_56676_ _83333_/Q _56675_/X _56676_/Y sky130_fd_sc_hd__nand2_4
X_87496_ _87749_/CLK _87496_/D _87496_/Q sky130_fd_sc_hd__dfxtp_4
X_53888_ _52370_/A _53875_/B _53888_/C _53888_/X sky130_fd_sc_hd__and3_4
X_58415_ _58415_/A _58415_/B _58415_/Y sky130_fd_sc_hd__nand2_4
X_43641_ _87330_/Q _43641_/Y sky130_fd_sc_hd__inv_2
X_55627_ _55610_/A _55627_/X sky130_fd_sc_hd__buf_2
X_74461_ _74442_/X _48582_/A _74461_/Y sky130_fd_sc_hd__nand2_4
X_86447_ _85557_/CLK _86447_/D _65087_/B sky130_fd_sc_hd__dfxtp_4
X_40853_ _40324_/X _82864_/Q _40852_/X _40853_/X sky130_fd_sc_hd__o21a_4
X_52839_ _52783_/A _52839_/X sky130_fd_sc_hd__buf_2
X_71673_ _58468_/Y _71669_/X _71672_/Y _71673_/Y sky130_fd_sc_hd__o21ai_4
X_59395_ _84743_/Q _63127_/A sky130_fd_sc_hd__inv_2
X_83659_ _85444_/CLK _70929_/Y _46898_/A sky130_fd_sc_hd__dfxtp_4
X_76200_ _76200_/A _76200_/B _76200_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_130_0_CLK clkbuf_7_65_0_CLK/X clkbuf_8_130_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_73412_ _73410_/X _73412_/B _73412_/C _73412_/Y sky130_fd_sc_hd__nand3_4
X_70624_ _53005_/B _70583_/X _70623_/Y _83738_/D sky130_fd_sc_hd__o21ai_4
X_46360_ _46348_/X _81208_/Q _46359_/X _46361_/A sky130_fd_sc_hd__o21ai_4
X_58346_ _84872_/Q _63295_/A sky130_fd_sc_hd__inv_2
X_77180_ _77172_/A _77177_/B _77171_/A _77181_/B sky130_fd_sc_hd__o21ai_4
X_55558_ _55524_/A _45485_/Y _55558_/Y sky130_fd_sc_hd__nor2_4
X_43572_ _40520_/X _43560_/X _87354_/Q _43561_/X _87354_/D sky130_fd_sc_hd__a2bb2o_4
X_74392_ _74390_/Y _72107_/X _74391_/Y _74392_/Y sky130_fd_sc_hd__a21boi_4
X_86378_ _83666_/CLK _49490_/Y _86378_/Q sky130_fd_sc_hd__dfxtp_4
X_40784_ _40784_/A _40847_/B sky130_fd_sc_hd__buf_2
X_45311_ _80671_/Q _45311_/X sky130_fd_sc_hd__buf_2
X_76131_ _81727_/D _76139_/B _76135_/A sky130_fd_sc_hd__xnor2_4
X_88117_ _88121_/CLK _88117_/D _67290_/B sky130_fd_sc_hd__dfxtp_4
X_42523_ _42521_/X _42522_/X _40724_/X _68955_/A _42506_/X _42524_/A
+ sky130_fd_sc_hd__o32ai_4
X_54509_ _54509_/A _54503_/B _54509_/C _54509_/D _54509_/X sky130_fd_sc_hd__and4_4
X_85329_ _83550_/CLK _55045_/Y _85329_/Q sky130_fd_sc_hd__dfxtp_4
X_73343_ _45930_/X _73343_/X sky130_fd_sc_hd__buf_2
X_46291_ _72052_/A _46719_/A sky130_fd_sc_hd__buf_2
X_70555_ _71859_/A _70549_/X _70568_/C _70550_/D _70555_/Y sky130_fd_sc_hd__nor4_4
X_58277_ _58277_/A _58280_/B _58277_/Y sky130_fd_sc_hd__nand2_4
X_55489_ _55489_/A _55489_/B _55489_/Y sky130_fd_sc_hd__nor2_4
X_48030_ _83542_/Q _53552_/B sky130_fd_sc_hd__inv_2
X_45242_ _45239_/Y _45241_/Y _45212_/X _45242_/X sky130_fd_sc_hd__a21o_4
X_57228_ _57227_/Y _85059_/D sky130_fd_sc_hd__inv_2
X_76062_ _81718_/D _76062_/B _76068_/A sky130_fd_sc_hd__xor2_4
X_88048_ _88087_/CLK _88048_/D _88048_/Q sky130_fd_sc_hd__dfxtp_4
X_42454_ _51238_/B _42430_/X _40560_/X _68361_/A _42453_/X _42454_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73274_ _69835_/B _73224_/X _73194_/X _73273_/Y _73274_/X sky130_fd_sc_hd__a211o_4
X_70486_ _71337_/A _70483_/B _71777_/B _70486_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_145_0_CLK clkbuf_7_72_0_CLK/X clkbuf_9_291_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_75013_ _75010_/Y _75013_/B _75014_/B sky130_fd_sc_hd__xor2_4
X_41405_ _41405_/A _41405_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_140_0_CLK clkbuf_9_70_0_CLK/X _81620_/CLK sky130_fd_sc_hd__clkbuf_1
X_72225_ _59081_/A _72225_/X sky130_fd_sc_hd__buf_2
X_45173_ _45166_/X _45170_/Y _45172_/Y _45173_/Y sky130_fd_sc_hd__a21oi_4
X_57159_ _57427_/A _56750_/Y _57096_/Y _57159_/Y sky130_fd_sc_hd__a21oi_4
X_42385_ _42378_/X _42369_/X _40371_/X _87889_/Q _42370_/X _42386_/A
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_10_770_0_CLK clkbuf_9_385_0_CLK/X _82124_/CLK sky130_fd_sc_hd__clkbuf_1
X_44124_ _44124_/A _72814_/A sky130_fd_sc_hd__buf_2
X_79821_ _79812_/Y _79829_/A _79820_/Y _79822_/B sky130_fd_sc_hd__a21oi_4
X_41336_ _40686_/A _41336_/X sky130_fd_sc_hd__buf_2
X_60170_ _60170_/A _60344_/A sky130_fd_sc_hd__buf_2
X_72156_ _58847_/A _72156_/X sky130_fd_sc_hd__buf_2
X_49981_ _49981_/A _53193_/B _49981_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_261_0_CLK clkbuf_8_130_0_CLK/X clkbuf_9_261_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_71107_ _50153_/B _71095_/X _71106_/Y _71107_/Y sky130_fd_sc_hd__o21ai_4
X_48932_ _48901_/A _52287_/B _48932_/Y sky130_fd_sc_hd__nand2_4
X_44055_ _86755_/Q _55125_/A sky130_fd_sc_hd__buf_2
X_79752_ _84220_/Q _83268_/Q _79752_/Y sky130_fd_sc_hd__nand2_4
X_41267_ _41255_/X _40741_/A _41266_/X _41267_/Y sky130_fd_sc_hd__o21ai_4
X_72087_ _83287_/Q _72051_/X _72086_/Y _72087_/Y sky130_fd_sc_hd__o21ai_4
X_76964_ _76895_/Y _81373_/D sky130_fd_sc_hd__inv_2
Xclkbuf_10_155_0_CLK clkbuf_9_77_0_CLK/X _81660_/CLK sky130_fd_sc_hd__clkbuf_1
X_43006_ _43005_/X _42477_/A _40532_/X _87607_/Q _42463_/A _43006_/Y
+ sky130_fd_sc_hd__o32ai_4
X_78703_ _78685_/A _78702_/Y _78669_/B _78703_/Y sky130_fd_sc_hd__o21ai_4
X_71038_ _71005_/A _71183_/A sky130_fd_sc_hd__buf_2
X_75915_ _84513_/Q _75915_/B _75915_/X sky130_fd_sc_hd__xor2_4
X_48863_ _50056_/A _48684_/B _48863_/Y sky130_fd_sc_hd__nand2_4
X_79683_ _79660_/X _79673_/X _79683_/Y sky130_fd_sc_hd__nand2_4
X_41198_ _41184_/X _40676_/A _41197_/X _41198_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_785_0_CLK clkbuf_9_392_0_CLK/X _82529_/CLK sky130_fd_sc_hd__clkbuf_1
X_76895_ _81677_/Q _76895_/B _76895_/Y sky130_fd_sc_hd__xnor2_4
X_47814_ _47814_/A _53257_/D sky130_fd_sc_hd__buf_2
X_78634_ _78614_/Y _78616_/A _78613_/A _78634_/X sky130_fd_sc_hd__o21a_4
X_63860_ _61844_/X _63860_/B _63860_/C _63860_/D _63860_/Y sky130_fd_sc_hd__nand4_4
X_75846_ _75846_/A _80895_/D sky130_fd_sc_hd__inv_2
X_48794_ _86481_/Q _48781_/X _48793_/Y _48794_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_276_0_CLK clkbuf_9_277_0_CLK/A clkbuf_9_276_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_62811_ _60273_/A _62812_/B sky130_fd_sc_hd__buf_2
X_47745_ _47745_/A _47745_/X sky130_fd_sc_hd__buf_2
X_78565_ _82804_/Q _78569_/A sky130_fd_sc_hd__inv_2
X_44957_ _56203_/C _44911_/X _44956_/X _44957_/Y sky130_fd_sc_hd__o21ai_4
X_75777_ _81016_/Q _80888_/D _80984_/D sky130_fd_sc_hd__xor2_4
X_63791_ _61364_/B _63790_/X _63757_/C _63776_/X _63791_/Y sky130_fd_sc_hd__nand4_4
X_72989_ _73183_/A _65551_/B _72989_/X sky130_fd_sc_hd__and2_4
X_65530_ _64967_/X _65559_/A sky130_fd_sc_hd__buf_2
X_77516_ _77505_/Y _77509_/B _77508_/A _77516_/X sky130_fd_sc_hd__o21a_4
X_43908_ _43869_/X _43908_/X sky130_fd_sc_hd__buf_2
X_62742_ _62681_/X _62742_/X sky130_fd_sc_hd__buf_2
X_74728_ _70637_/A _74796_/B sky130_fd_sc_hd__buf_2
X_47676_ _47692_/A _47692_/B _47692_/C _53181_/D _47676_/X sky130_fd_sc_hd__and4_4
X_78496_ _78474_/A _78473_/X _78496_/X sky130_fd_sc_hd__xor2_4
X_44888_ _44887_/X _44889_/A sky130_fd_sc_hd__buf_2
X_49415_ _49415_/A _49415_/X sky130_fd_sc_hd__buf_2
X_46627_ _58577_/A _46622_/X _46626_/Y _46627_/Y sky130_fd_sc_hd__o21ai_4
X_65461_ _65458_/X _65461_/B _65461_/Y sky130_fd_sc_hd__nand2_4
X_77447_ _77447_/A _77444_/Y _77446_/Y _77447_/X sky130_fd_sc_hd__or3_4
X_43839_ _43810_/X _43824_/X _41174_/X _68681_/B _43811_/X _43840_/A
+ sky130_fd_sc_hd__o32ai_4
X_62673_ _62673_/A _62673_/B _84392_/Q _62673_/Y sky130_fd_sc_hd__nor3_4
X_74659_ _74659_/A _74659_/Y sky130_fd_sc_hd__inv_2
X_67200_ _67082_/A _67250_/A sky130_fd_sc_hd__buf_2
X_64412_ _64402_/X _64379_/B _64412_/C _64412_/X sky130_fd_sc_hd__and3_4
X_61624_ _61634_/A _61634_/B _79133_/B _61624_/Y sky130_fd_sc_hd__nor3_4
X_49346_ _49327_/X _54079_/B _49346_/Y sky130_fd_sc_hd__nand2_4
X_68180_ _68160_/A _68180_/X sky130_fd_sc_hd__buf_2
X_46558_ _82918_/Q _46527_/X _46558_/X sky130_fd_sc_hd__or2_4
X_65392_ _65289_/A _65392_/B _65392_/X sky130_fd_sc_hd__and2_4
X_77378_ _82221_/Q _77382_/A sky130_fd_sc_hd__inv_2
Xclkbuf_10_723_0_CLK clkbuf_9_361_0_CLK/X _87022_/CLK sky130_fd_sc_hd__clkbuf_1
X_67131_ _67131_/A _87612_/Q _67131_/X sky130_fd_sc_hd__and2_4
X_79117_ _78998_/B _79117_/Y sky130_fd_sc_hd__inv_2
X_45509_ _83002_/Q _45401_/X _45508_/X _45510_/A sky130_fd_sc_hd__o21ai_4
X_64343_ _64319_/X _64343_/B _64333_/X _64343_/X sky130_fd_sc_hd__and3_4
X_76329_ _76316_/A _76327_/Y _76328_/Y _76338_/A sky130_fd_sc_hd__o21a_4
X_49277_ _49273_/A _46417_/B _49277_/Y sky130_fd_sc_hd__nand2_4
X_61555_ _61546_/A _61546_/B _84471_/Q _61555_/Y sky130_fd_sc_hd__nor3_4
X_46489_ _83636_/Q _52526_/B sky130_fd_sc_hd__inv_2
Xclkbuf_9_214_0_CLK clkbuf_9_214_0_CLK/A clkbuf_9_214_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_48228_ _47937_/B _53504_/B sky130_fd_sc_hd__buf_2
X_60506_ _60500_/Y _60501_/Y _60482_/A _63247_/A sky130_fd_sc_hd__o21a_4
X_67062_ _45915_/X _67062_/X sky130_fd_sc_hd__buf_2
X_79048_ _82524_/D _79048_/B _79049_/A sky130_fd_sc_hd__and2_4
X_64274_ _64274_/A _64274_/X sky130_fd_sc_hd__buf_2
X_61486_ _61479_/Y _61482_/Y _61464_/X _61483_/Y _61485_/Y _61486_/X
+ sky130_fd_sc_hd__a41o_4
Xclkbuf_10_108_0_CLK clkbuf_9_54_0_CLK/X _84531_/CLK sky130_fd_sc_hd__clkbuf_1
X_66013_ _65924_/X _84986_/Q _65950_/X _66012_/X _66013_/X sky130_fd_sc_hd__a211o_4
X_63225_ _63288_/A _64434_/B _63312_/C _63192_/D _63225_/X sky130_fd_sc_hd__and4_4
X_48159_ _52093_/A _50391_/A sky130_fd_sc_hd__buf_2
X_60437_ _60436_/Y _84616_/D sky130_fd_sc_hd__inv_2
Xclkbuf_10_738_0_CLK clkbuf_9_369_0_CLK/X _86834_/CLK sky130_fd_sc_hd__clkbuf_1
X_81010_ _84197_/CLK _84218_/Q _81010_/Q sky130_fd_sc_hd__dfxtp_4
X_51170_ _51170_/A _51192_/C sky130_fd_sc_hd__buf_2
X_63156_ _63144_/X _84828_/Q _63146_/C _63135_/D _63156_/X sky130_fd_sc_hd__and4_4
X_60368_ _79566_/B _60323_/X _60305_/Y _60367_/Y _60368_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_9_229_0_CLK clkbuf_8_114_0_CLK/X clkbuf_9_229_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_50121_ _64948_/B _50113_/X _50120_/Y _50121_/Y sky130_fd_sc_hd__o21ai_4
X_62107_ _59605_/Y _62158_/C sky130_fd_sc_hd__buf_2
X_67964_ _67914_/X _67964_/B _67964_/X sky130_fd_sc_hd__and2_4
X_63087_ _60606_/X _63087_/X sky130_fd_sc_hd__buf_2
X_60299_ _60299_/A _60296_/X _60299_/C _60299_/Y sky130_fd_sc_hd__nand3_4
X_69703_ _69865_/A _88329_/Q _69703_/X sky130_fd_sc_hd__and2_4
X_50052_ _50056_/A _48878_/B _50052_/Y sky130_fd_sc_hd__nand2_4
X_66915_ _66915_/A _66915_/X sky130_fd_sc_hd__buf_2
X_62038_ _62037_/X _62021_/B _58487_/A _62020_/X _62038_/X sky130_fd_sc_hd__and4_4
X_82961_ _82961_/CLK _82769_/Q _82961_/Q sky130_fd_sc_hd__dfxtp_4
X_67895_ _67992_/A _88220_/Q _67895_/X sky130_fd_sc_hd__and2_4
X_84700_ _84329_/CLK _84700_/D _80484_/A sky130_fd_sc_hd__dfxtp_4
X_81912_ _82103_/CLK _81912_/D _82288_/D sky130_fd_sc_hd__dfxtp_4
X_69634_ _43126_/A _69506_/X _68436_/X _69633_/X _69634_/X sky130_fd_sc_hd__a211o_4
X_54860_ _85364_/Q _54839_/X _54859_/Y _54860_/Y sky130_fd_sc_hd__o21ai_4
X_66846_ _88392_/Q _66751_/X _66801_/X _66845_/X _66846_/X sky130_fd_sc_hd__a211o_4
X_85680_ _84797_/CLK _53192_/Y _85680_/Q sky130_fd_sc_hd__dfxtp_4
X_82892_ _86935_/CLK _78153_/B _82892_/Q sky130_fd_sc_hd__dfxtp_4
X_53811_ _53809_/Y _53773_/X _53810_/X _53811_/Y sky130_fd_sc_hd__a21oi_4
X_84631_ _84649_/CLK _60328_/X _79691_/A sky130_fd_sc_hd__dfxtp_4
X_81843_ _81857_/CLK _81875_/Q _77471_/A sky130_fd_sc_hd__dfxtp_4
X_69565_ _69580_/A _87315_/Q _69565_/X sky130_fd_sc_hd__and2_4
X_54791_ _85377_/Q _54784_/X _54790_/Y _54791_/Y sky130_fd_sc_hd__o21ai_4
X_66777_ _66728_/A _88139_/Q _66777_/X sky130_fd_sc_hd__and2_4
X_63989_ _63761_/A _64052_/D sky130_fd_sc_hd__buf_2
X_56530_ _56139_/X _56528_/X _56529_/Y _85161_/D sky130_fd_sc_hd__o21ai_4
X_68516_ _68300_/X _68516_/X sky130_fd_sc_hd__buf_2
X_87350_ _82899_/CLK _43578_/X _87350_/Q sky130_fd_sc_hd__dfxtp_4
X_53742_ _85577_/Q _53729_/X _53741_/Y _53742_/Y sky130_fd_sc_hd__o21ai_4
X_65728_ _65634_/A _65802_/B _65728_/C _65728_/Y sky130_fd_sc_hd__nor3_4
X_84562_ _84562_/CLK _84562_/D _84562_/Q sky130_fd_sc_hd__dfxtp_4
X_50954_ _50951_/Y _50928_/X _50953_/X _86101_/D sky130_fd_sc_hd__a21oi_4
X_81774_ _82053_/CLK _76061_/X _81774_/Q sky130_fd_sc_hd__dfxtp_4
X_69496_ _69493_/X _69495_/X _69399_/X _69496_/X sky130_fd_sc_hd__a21o_4
X_86301_ _86301_/CLK _49911_/Y _72174_/B sky130_fd_sc_hd__dfxtp_4
X_83513_ _83507_/CLK _71400_/X _83513_/Q sky130_fd_sc_hd__dfxtp_4
X_56461_ _56463_/A _56528_/A sky130_fd_sc_hd__buf_2
X_68447_ _68447_/A _68447_/X sky130_fd_sc_hd__buf_2
X_80725_ _84269_/CLK _80725_/D _80725_/Q sky130_fd_sc_hd__dfxtp_4
X_87281_ _88097_/CLK _87281_/D _69165_/B sky130_fd_sc_hd__dfxtp_4
X_53673_ _53670_/Y _53653_/X _53672_/X _85591_/D sky130_fd_sc_hd__a21oi_4
X_65659_ _65656_/X _65658_/X _65614_/X _65659_/X sky130_fd_sc_hd__a21o_4
X_84493_ _84493_/CLK _61269_/Y _84493_/Q sky130_fd_sc_hd__dfxtp_4
X_50885_ _86113_/Q _50882_/X _50884_/Y _50885_/Y sky130_fd_sc_hd__o21ai_4
X_58200_ _83373_/Q _58200_/Y sky130_fd_sc_hd__inv_2
X_55412_ _55200_/C _55412_/Y sky130_fd_sc_hd__inv_2
X_86232_ _86235_/CLK _86232_/D _86232_/Q sky130_fd_sc_hd__dfxtp_4
X_52624_ _52624_/A _54314_/B _52624_/Y sky130_fd_sc_hd__nand2_4
X_59180_ _59176_/Y _59179_/Y _59140_/X _59180_/X sky130_fd_sc_hd__a21o_4
X_83444_ _83763_/CLK _83444_/D _83444_/Q sky130_fd_sc_hd__dfxtp_4
X_56392_ _56383_/X _56386_/B _56392_/C _56392_/Y sky130_fd_sc_hd__nand3_4
X_80656_ _86772_/CLK _74835_/Y _80656_/Q sky130_fd_sc_hd__dfxtp_4
X_68378_ _66673_/X _69088_/A sky130_fd_sc_hd__buf_2
XPHY_304 sky130_fd_sc_hd__decap_3
X_58131_ _58721_/A _58649_/B sky130_fd_sc_hd__buf_2
XPHY_315 sky130_fd_sc_hd__decap_3
X_55343_ _55317_/A _57137_/A _55343_/X sky130_fd_sc_hd__and2_4
X_67329_ _63055_/A _68461_/A sky130_fd_sc_hd__buf_2
X_86163_ _85557_/CLK _86163_/D _86163_/Q sky130_fd_sc_hd__dfxtp_4
X_52555_ _52567_/A _54073_/B _52555_/Y sky130_fd_sc_hd__nand2_4
XPHY_326 sky130_fd_sc_hd__decap_3
X_83375_ _83372_/CLK _71791_/Y _83375_/Q sky130_fd_sc_hd__dfxtp_4
X_80587_ _84774_/Q _84166_/Q _80587_/X sky130_fd_sc_hd__xor2_4
XPHY_337 sky130_fd_sc_hd__decap_3
XPHY_348 sky130_fd_sc_hd__decap_3
XPHY_359 sky130_fd_sc_hd__decap_3
X_85114_ _85114_/CLK _85114_/D _45501_/A sky130_fd_sc_hd__dfxtp_4
X_51506_ _51502_/Y _51503_/X _51505_/X _85998_/D sky130_fd_sc_hd__a21oi_4
X_58062_ _58679_/A _58062_/X sky130_fd_sc_hd__buf_2
X_70340_ _70338_/A _70333_/B _83087_/Q _70332_/X _70340_/X sky130_fd_sc_hd__and4_4
X_82326_ _86758_/CLK _77147_/B _82326_/Q sky130_fd_sc_hd__dfxtp_4
X_55274_ _82982_/Q _55272_/X _55140_/X _55273_/X _55274_/X sky130_fd_sc_hd__a211o_4
X_86094_ _85778_/CLK _50990_/Y _86094_/Q sky130_fd_sc_hd__dfxtp_4
X_52486_ _52486_/A _52486_/X sky130_fd_sc_hd__buf_2
X_57013_ _57009_/Y _57012_/Y _44039_/X _57013_/X sky130_fd_sc_hd__o21a_4
X_54225_ _51822_/A _54253_/A sky130_fd_sc_hd__buf_2
X_85045_ _85042_/CLK _57260_/X _45585_/A sky130_fd_sc_hd__dfxtp_4
X_51437_ _51218_/X _51456_/A sky130_fd_sc_hd__buf_2
X_70271_ _70269_/X _74801_/B _70270_/X _83816_/D sky130_fd_sc_hd__a21o_4
X_82257_ _85381_/CLK _82257_/D _82257_/Q sky130_fd_sc_hd__dfxtp_4
X_72010_ _71993_/X _53834_/B _72010_/Y sky130_fd_sc_hd__nand2_4
X_81208_ _82933_/CLK _75060_/X _81208_/Q sky130_fd_sc_hd__dfxtp_4
X_42170_ _42096_/A _42170_/X sky130_fd_sc_hd__buf_2
X_54156_ _54160_/A _54160_/B _54146_/X _52989_/D _54156_/X sky130_fd_sc_hd__and4_4
X_51368_ _51367_/X _46539_/A _51368_/X sky130_fd_sc_hd__and2_4
X_82188_ _85404_/CLK _82188_/D _82188_/Q sky130_fd_sc_hd__dfxtp_4
X_53107_ _53107_/A _53113_/B _53107_/C _53107_/D _53107_/X sky130_fd_sc_hd__and4_4
X_41121_ _41121_/A _41121_/X sky130_fd_sc_hd__buf_2
X_50319_ _86224_/Q _50316_/X _50318_/Y _50319_/Y sky130_fd_sc_hd__o21ai_4
X_81139_ _80854_/CLK _80763_/Q _81139_/Q sky130_fd_sc_hd__dfxtp_4
X_58964_ _58904_/X _85762_/Q _58928_/X _58964_/X sky130_fd_sc_hd__o21a_4
X_54087_ _53801_/B _54087_/B _54087_/Y sky130_fd_sc_hd__nand2_4
X_51299_ _51297_/Y _51289_/X _51298_/X _51299_/Y sky130_fd_sc_hd__a21oi_4
X_86996_ _88363_/CLK _44698_/Y _44697_/A sky130_fd_sc_hd__dfxtp_4
X_41052_ _40879_/B _41019_/B _41052_/X sky130_fd_sc_hd__or2_4
X_53038_ _53065_/A _53038_/X sky130_fd_sc_hd__buf_2
X_57915_ _57773_/X _85716_/Q _44177_/X _57915_/X sky130_fd_sc_hd__o21a_4
X_73961_ _70117_/C _73939_/X _73960_/X _83129_/D sky130_fd_sc_hd__o21ai_4
X_85947_ _82206_/CLK _85947_/D _85947_/Q sky130_fd_sc_hd__dfxtp_4
X_58895_ _84792_/Q _58871_/X _58888_/X _58894_/X _58895_/Y sky130_fd_sc_hd__a2bb2oi_4
X_75700_ _75677_/Y _80782_/D sky130_fd_sc_hd__inv_2
X_72912_ _72908_/X _85596_/Q _72909_/X _72911_/X _72912_/X sky130_fd_sc_hd__a211o_4
X_57846_ _57846_/A _57845_/X _57846_/Y sky130_fd_sc_hd__nor2_4
X_45860_ _56920_/B _45798_/X _44889_/A _45860_/X sky130_fd_sc_hd__o21a_4
X_76680_ _76679_/Y _76666_/Y _76673_/A _76680_/Y sky130_fd_sc_hd__o21ai_4
X_73892_ _73892_/A _73869_/X _73892_/Y sky130_fd_sc_hd__nor2_4
X_85878_ _86196_/CLK _52157_/Y _85878_/Q sky130_fd_sc_hd__dfxtp_4
X_44811_ _41635_/Y _43939_/X _67361_/B _43941_/X _86942_/D sky130_fd_sc_hd__a2bb2o_4
X_75631_ _80776_/D _75619_/A _75631_/X sky130_fd_sc_hd__and2_4
X_87617_ _88387_/CLK _87617_/D _66995_/B sky130_fd_sc_hd__dfxtp_4
X_72843_ _72816_/X _72843_/B _72843_/X sky130_fd_sc_hd__and2_4
X_84829_ _84829_/CLK _58521_/Y _84829_/Q sky130_fd_sc_hd__dfxtp_4
X_45791_ _45784_/X _45788_/Y _45790_/Y _86854_/D sky130_fd_sc_hd__a21oi_4
X_57777_ _69768_/A _58002_/A sky130_fd_sc_hd__buf_2
X_54989_ _54985_/A _47582_/A _54989_/Y sky130_fd_sc_hd__nand2_4
X_47530_ _47530_/A _47530_/X sky130_fd_sc_hd__buf_2
X_59516_ _59516_/A _59562_/B sky130_fd_sc_hd__buf_2
X_78350_ _78350_/A _78345_/X _78346_/Y _78353_/B sky130_fd_sc_hd__nand3_4
X_44742_ _44532_/A _44742_/X sky130_fd_sc_hd__buf_2
X_56728_ _56842_/A _56700_/C _56676_/Y _57140_/A sky130_fd_sc_hd__nor3_4
X_75562_ _75562_/A _75552_/X _75559_/X _75563_/B sky130_fd_sc_hd__nand3_4
X_87548_ _88087_/CLK _43186_/X _73341_/A sky130_fd_sc_hd__dfxtp_4
X_41954_ _41932_/X _41951_/X _40707_/X _74051_/A _41953_/X _41955_/A
+ sky130_fd_sc_hd__o32ai_4
X_72774_ _72770_/X _72773_/X _72737_/X _72774_/X sky130_fd_sc_hd__a21o_4
X_77301_ _77301_/A _77301_/B _77318_/B sky130_fd_sc_hd__nor2_4
X_74513_ _46347_/A _50556_/B _74513_/Y sky130_fd_sc_hd__nand2_4
X_40905_ _40756_/A _40905_/X sky130_fd_sc_hd__buf_2
X_47461_ _86632_/Q _47429_/X _47460_/Y _47461_/Y sky130_fd_sc_hd__o21ai_4
X_71725_ _71729_/A _71302_/X _71724_/X _71725_/Y sky130_fd_sc_hd__nand3_4
X_59447_ _84730_/Q _59448_/A sky130_fd_sc_hd__inv_2
X_78281_ _78262_/X _78274_/A _78284_/B _78281_/Y sky130_fd_sc_hd__nand3_4
X_44673_ _44658_/X _44659_/X _40581_/X _87005_/Q _44660_/X _44674_/A
+ sky130_fd_sc_hd__o32ai_4
X_56659_ _56700_/C _56659_/Y sky130_fd_sc_hd__inv_2
X_75493_ _75493_/A _75492_/Y _75493_/Y sky130_fd_sc_hd__nor2_4
X_87479_ _87749_/CLK _87479_/D _87479_/Q sky130_fd_sc_hd__dfxtp_4
X_41885_ _42081_/A _42059_/A sky130_fd_sc_hd__buf_2
X_49200_ _40380_/X _81762_/Q _49199_/Y _72113_/A sky130_fd_sc_hd__o21ai_4
X_46412_ _46387_/A _46412_/B _46412_/Y sky130_fd_sc_hd__nand2_4
X_77232_ _77229_/Y _77231_/Y _77232_/Y sky130_fd_sc_hd__nor2_4
X_43624_ _55102_/A _43624_/X sky130_fd_sc_hd__buf_2
X_74444_ _83065_/Q _74441_/X _74443_/Y _74444_/Y sky130_fd_sc_hd__o21ai_4
X_40836_ _40836_/A _40836_/X sky130_fd_sc_hd__buf_2
X_47392_ _47418_/A _47408_/B _47377_/X _53019_/D _47392_/X sky130_fd_sc_hd__and4_4
X_59378_ _59325_/X _59376_/Y _59377_/Y _59342_/X _59329_/X _59378_/X
+ sky130_fd_sc_hd__o32a_4
X_71656_ _71660_/A _71223_/B _71660_/C _71656_/Y sky130_fd_sc_hd__nand3_4
X_49131_ _52385_/B _72079_/B sky130_fd_sc_hd__buf_2
X_46343_ _53980_/B _49245_/B sky130_fd_sc_hd__buf_2
X_70607_ _52986_/B _70584_/X _70606_/Y _70607_/Y sky130_fd_sc_hd__o21ai_4
X_58329_ _58329_/A _58331_/A sky130_fd_sc_hd__inv_2
X_77163_ _77163_/A _81921_/Q _77173_/C sky130_fd_sc_hd__nand2_4
X_43555_ _43542_/X _43546_/X _40474_/X _87362_/Q _43549_/X _43555_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74375_ _74375_/A _72113_/B _74366_/C _74375_/X sky130_fd_sc_hd__and3_4
X_40767_ _40767_/A _40767_/X sky130_fd_sc_hd__buf_2
X_71587_ _71581_/X _83448_/Q _71586_/Y _83448_/D sky130_fd_sc_hd__a21o_4
X_76114_ _81725_/D _76116_/B _76114_/X sky130_fd_sc_hd__or2_4
X_42506_ _42612_/A _42506_/X sky130_fd_sc_hd__buf_2
X_61340_ _61340_/A _61368_/B sky130_fd_sc_hd__buf_2
X_49062_ _49057_/Y _49038_/X _49061_/X _49062_/Y sky130_fd_sc_hd__a21oi_4
X_73326_ _69865_/B _72865_/X _72866_/X _73326_/X sky130_fd_sc_hd__o21a_4
X_70538_ _70554_/A _70538_/X sky130_fd_sc_hd__buf_2
X_46274_ _46274_/A _46328_/B _46274_/X sky130_fd_sc_hd__or2_4
X_77094_ _82095_/Q _77094_/B _77094_/X sky130_fd_sc_hd__xor2_4
X_43486_ _41701_/X _43484_/X _87398_/Q _43485_/X _87398_/D sky130_fd_sc_hd__a2bb2o_4
X_40698_ _49048_/A _40698_/X sky130_fd_sc_hd__buf_2
X_48013_ _48005_/Y _48007_/X _48012_/X _86577_/D sky130_fd_sc_hd__a21oi_4
X_45225_ _85164_/Q _45209_/X _45189_/X _45225_/X sky130_fd_sc_hd__o21a_4
X_76045_ _81523_/Q _81747_/D _81772_/D sky130_fd_sc_hd__xor2_4
X_42437_ _40528_/X _42434_/X _87864_/Q _42435_/X _87864_/D sky130_fd_sc_hd__a2bb2o_4
X_61271_ _61271_/A _61096_/X _61153_/C _61103_/X _61271_/Y sky130_fd_sc_hd__nand4_4
X_73257_ _73257_/A _73257_/X sky130_fd_sc_hd__buf_2
X_70469_ DATA_TO_HASH[6] _71424_/C sky130_fd_sc_hd__buf_2
X_63010_ _63010_/A _63010_/X sky130_fd_sc_hd__buf_2
X_60222_ _59640_/A _59615_/A _60222_/C _60222_/X sky130_fd_sc_hd__and3_4
X_72208_ _72143_/X _85370_/Q _72207_/X _72208_/Y sky130_fd_sc_hd__o21ai_4
X_45156_ _45156_/A _45182_/B _45156_/Y sky130_fd_sc_hd__nand2_4
X_42368_ _41768_/X _42356_/X _87897_/Q _42357_/X _87897_/D sky130_fd_sc_hd__a2bb2o_4
X_73188_ _73188_/A _73188_/B _73188_/Y sky130_fd_sc_hd__nand2_4
X_44107_ _43990_/Y _45938_/A _44107_/C _44107_/X sky130_fd_sc_hd__or3_4
X_79804_ _64841_/Y _72214_/Y _79803_/Y _79804_/X sky130_fd_sc_hd__o21a_4
X_41319_ _41513_/A _41319_/B _41319_/X sky130_fd_sc_hd__or2_4
X_72139_ _72277_/A _72139_/B _72139_/Y sky130_fd_sc_hd__nor2_4
X_60153_ _60151_/X _64638_/B _60153_/C _60153_/Y sky130_fd_sc_hd__nand3_4
X_49964_ _49973_/A _49943_/B _49973_/C _53177_/D _49964_/X sky130_fd_sc_hd__and4_4
X_45087_ _45237_/A _45087_/X sky130_fd_sc_hd__buf_2
X_42299_ _42279_/X _42297_/X _41574_/X _87933_/Q _42298_/X _42300_/A
+ sky130_fd_sc_hd__o32ai_4
X_77996_ _82255_/Q _81967_/Q _78012_/A sky130_fd_sc_hd__xnor2_4
X_48915_ _48915_/A _48959_/B _50578_/B sky130_fd_sc_hd__nor2_4
X_44038_ _44037_/X _44038_/X sky130_fd_sc_hd__buf_2
X_79735_ _79731_/Y _79734_/Y _79735_/X sky130_fd_sc_hd__xor2_4
X_64961_ _64961_/A _65984_/A sky130_fd_sc_hd__buf_2
X_60084_ _60084_/A _62198_/B _59976_/A _59985_/X _60085_/A sky130_fd_sc_hd__and4_4
X_76947_ _76946_/X _76953_/B sky130_fd_sc_hd__inv_2
X_49895_ _49901_/A _53109_/B _49895_/Y sky130_fd_sc_hd__nand2_4
X_66700_ _66602_/A _66700_/B _66700_/X sky130_fd_sc_hd__and2_4
X_63912_ _64328_/A _63912_/X sky130_fd_sc_hd__buf_2
X_48846_ _48844_/Y _48840_/X _48845_/X _86472_/D sky130_fd_sc_hd__a21oi_4
X_67680_ _87397_/Q _67628_/X _67581_/X _67679_/X _67680_/X sky130_fd_sc_hd__a211o_4
X_79666_ _79645_/B _79662_/X _79665_/Y _79666_/Y sky130_fd_sc_hd__a21oi_4
X_64892_ _64889_/Y _64814_/X _64891_/Y _84223_/D sky130_fd_sc_hd__a21o_4
X_76878_ _76910_/C _76877_/Y _76879_/B sky130_fd_sc_hd__xnor2_4
X_78617_ _78616_/Y _78617_/B _78617_/Y sky130_fd_sc_hd__nand2_4
X_66631_ _87441_/Q _66571_/X _66629_/X _66630_/X _66631_/X sky130_fd_sc_hd__a211o_4
X_63843_ _61831_/X _63860_/B _63860_/C _63860_/D _63843_/Y sky130_fd_sc_hd__nand4_4
X_75829_ _81102_/Q _75829_/B _75830_/B sky130_fd_sc_hd__xnor2_4
X_48777_ _48777_/A _52163_/B _48777_/Y sky130_fd_sc_hd__nand2_4
X_79597_ _79597_/A _79596_/Y _79598_/A sky130_fd_sc_hd__xor2_4
X_45989_ _45989_/A _45989_/Y sky130_fd_sc_hd__inv_2
X_69350_ _69347_/X _69349_/X _69171_/X _69350_/Y sky130_fd_sc_hd__a21oi_4
X_47728_ _72378_/A _47714_/X _47727_/Y _47728_/Y sky130_fd_sc_hd__o21ai_4
X_66562_ _69582_/A _66562_/X sky130_fd_sc_hd__buf_2
X_78548_ _78534_/Y _78546_/Y _78547_/Y _78548_/X sky130_fd_sc_hd__o21a_4
X_63774_ _64026_/A _63820_/B sky130_fd_sc_hd__buf_2
X_60986_ _84545_/Q _60979_/X _60980_/Y _60985_/Y _60986_/Y sky130_fd_sc_hd__a2bb2oi_4
X_68301_ _68300_/X _68301_/X sky130_fd_sc_hd__buf_2
X_65513_ _65449_/A _65546_/B _84196_/Q _65513_/X sky130_fd_sc_hd__and3_4
X_62725_ _62711_/A _64286_/C _62676_/C _62738_/D _62725_/X sky130_fd_sc_hd__and4_4
X_69281_ _69276_/X _69280_/X _69281_/Y sky130_fd_sc_hd__nand2_4
X_47659_ _47649_/A _53174_/B _47659_/Y sky130_fd_sc_hd__nand2_4
X_66493_ _65262_/X _66521_/B _65265_/X _66493_/Y sky130_fd_sc_hd__nand3_4
X_78479_ _78463_/B _78463_/A _78465_/A _78479_/Y sky130_fd_sc_hd__a21boi_4
Xclkbuf_10_662_0_CLK clkbuf_9_331_0_CLK/X _87686_/CLK sky130_fd_sc_hd__clkbuf_1
X_80510_ _80482_/Y _80485_/Y _80495_/X _80498_/Y _80510_/X sky130_fd_sc_hd__o22a_4
X_68232_ _67443_/X _67445_/X _68209_/X _68232_/Y sky130_fd_sc_hd__a21oi_4
X_65444_ _65753_/A _65444_/B _65444_/X sky130_fd_sc_hd__and2_4
X_50670_ _50657_/A _52367_/B _50670_/Y sky130_fd_sc_hd__nand2_4
X_62656_ _62655_/Y _62658_/A sky130_fd_sc_hd__buf_2
X_81490_ _81265_/CLK _81490_/D _81490_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_153_0_CLK clkbuf_8_76_0_CLK/X clkbuf_9_153_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_49329_ _49325_/Y _49326_/X _49328_/Y _49329_/Y sky130_fd_sc_hd__a21boi_4
X_61607_ _61558_/A _61607_/B _61590_/C _61607_/Y sky130_fd_sc_hd__nand3_4
X_80441_ _80441_/A _84152_/Q _80452_/A sky130_fd_sc_hd__xor2_4
X_68163_ _84023_/Q _68160_/X _68162_/X _68163_/X sky130_fd_sc_hd__a21bo_4
Xclkbuf_9_80_0_CLK clkbuf_8_40_0_CLK/X clkbuf_9_80_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_65375_ _65074_/A _65375_/B _65375_/X sky130_fd_sc_hd__and2_4
X_62587_ _62620_/A _63672_/B _62532_/X _62587_/Y sky130_fd_sc_hd__nand3_4
X_67114_ _67109_/X _67112_/X _67113_/X _67114_/Y sky130_fd_sc_hd__a21oi_4
X_52340_ _52262_/A _52340_/X sky130_fd_sc_hd__buf_2
X_64326_ _64267_/A _64326_/X sky130_fd_sc_hd__buf_2
X_83160_ _85895_/CLK _73223_/X _83160_/Q sky130_fd_sc_hd__dfxtp_4
X_61538_ _61499_/A _61538_/B _61538_/C _61538_/Y sky130_fd_sc_hd__nand3_4
X_80372_ _80370_/X _80372_/B _80372_/X sky130_fd_sc_hd__xor2_4
X_68094_ _68088_/X _66597_/Y _68089_/X _68093_/Y _68094_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_677_0_CLK clkbuf_9_338_0_CLK/X _87141_/CLK sky130_fd_sc_hd__clkbuf_1
X_82111_ _82860_/CLK _82123_/Q _82111_/Q sky130_fd_sc_hd__dfxtp_4
X_67045_ _80910_/D _66971_/X _67044_/X _67045_/X sky130_fd_sc_hd__a21bo_4
X_52271_ _52271_/A _52293_/A sky130_fd_sc_hd__buf_2
X_64257_ _64257_/A _64301_/B _64257_/Y sky130_fd_sc_hd__nor2_4
X_83091_ _81627_/CLK _83091_/D _70328_/C sky130_fd_sc_hd__dfxtp_4
X_61469_ _61686_/A _61484_/B sky130_fd_sc_hd__buf_2
Xclkbuf_9_168_0_CLK clkbuf_8_84_0_CLK/X clkbuf_9_168_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_54010_ _85523_/Q _53989_/X _54009_/Y _54010_/Y sky130_fd_sc_hd__o21ai_4
X_51222_ _51212_/A _51222_/B _51222_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_95_0_CLK clkbuf_9_94_0_CLK/A clkbuf_9_95_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_63208_ _63247_/A _63267_/D sky130_fd_sc_hd__buf_2
X_82042_ _82139_/CLK _77951_/B _82042_/Q sky130_fd_sc_hd__dfxtp_4
X_64188_ _64185_/X _64186_/X _64187_/Y _64188_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_600_0_CLK clkbuf_9_300_0_CLK/X _80962_/CLK sky130_fd_sc_hd__clkbuf_1
X_51153_ _86064_/Q _51128_/X _51152_/Y _51153_/Y sky130_fd_sc_hd__o21ai_4
X_63139_ _63139_/A _63113_/B _63103_/C _63092_/D _63139_/X sky130_fd_sc_hd__or4_4
X_86850_ _86882_/CLK _45852_/Y _63333_/B sky130_fd_sc_hd__dfxtp_4
X_68996_ _68992_/X _68995_/X _68737_/X _68996_/Y sky130_fd_sc_hd__a21oi_4
X_50104_ _86263_/Q _50088_/X _50103_/Y _50104_/Y sky130_fd_sc_hd__o21ai_4
X_85801_ _85514_/CLK _52544_/Y _65234_/B sky130_fd_sc_hd__dfxtp_4
X_51084_ _51084_/A _51071_/B _51071_/C _52775_/D _51084_/X sky130_fd_sc_hd__and4_4
X_55961_ _56386_/C _55689_/A _55611_/X _55960_/X _55961_/X sky130_fd_sc_hd__a211o_4
X_67947_ _84048_/Q _67925_/X _67946_/X _67947_/X sky130_fd_sc_hd__a21bo_4
X_86781_ _82317_/CLK _46073_/X _86781_/Q sky130_fd_sc_hd__dfxtp_4
X_83993_ _82896_/CLK _83993_/D _83993_/Q sky130_fd_sc_hd__dfxtp_4
X_57700_ _58098_/A _57700_/X sky130_fd_sc_hd__buf_2
X_54912_ _54893_/X _47741_/Y _54912_/Y sky130_fd_sc_hd__nand2_4
X_50035_ _49930_/X _51750_/C sky130_fd_sc_hd__buf_2
X_85732_ _86342_/CLK _52913_/Y _85732_/Q sky130_fd_sc_hd__dfxtp_4
X_58680_ _58605_/X _85944_/Q _58679_/X _58680_/X sky130_fd_sc_hd__o21a_4
X_82944_ _82368_/CLK _78112_/X _46265_/A sky130_fd_sc_hd__dfxtp_4
X_55892_ _55864_/X _56073_/A _74317_/C _55891_/X _55892_/X sky130_fd_sc_hd__and4_4
X_67878_ _81483_/D _67806_/X _67877_/X _84051_/D sky130_fd_sc_hd__a21bo_4
Xclkbuf_10_615_0_CLK clkbuf_9_307_0_CLK/X _80740_/CLK sky130_fd_sc_hd__clkbuf_1
X_57631_ _84965_/Q _57603_/X _57630_/Y _57631_/Y sky130_fd_sc_hd__o21ai_4
X_69617_ _69567_/A _69617_/X sky130_fd_sc_hd__buf_2
X_54843_ _54857_/A _54843_/B _54857_/C _53151_/D _54843_/X sky130_fd_sc_hd__and4_4
X_66829_ _87944_/Q _66759_/X _66807_/X _66828_/X _66829_/X sky130_fd_sc_hd__a211o_4
X_85663_ _85439_/CLK _53279_/Y _85663_/Q sky130_fd_sc_hd__dfxtp_4
X_82875_ _82596_/CLK _82467_/Q _82875_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_106_0_CLK clkbuf_8_53_0_CLK/X clkbuf_9_106_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_87402_ _86932_/CLK _87402_/D _87402_/Q sky130_fd_sc_hd__dfxtp_4
X_84614_ _84477_/CLK _84614_/D _79154_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_33_0_CLK clkbuf_9_33_0_CLK/A clkbuf_9_33_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_57562_ _47714_/A _57562_/X sky130_fd_sc_hd__buf_2
X_69548_ _87009_/Q _69414_/X _69430_/X _69547_/X _69548_/X sky130_fd_sc_hd__a211o_4
X_81826_ _84441_/CLK _81858_/Q _77233_/A sky130_fd_sc_hd__dfxtp_4
X_88382_ _88128_/CLK _40498_/X _88382_/Q sky130_fd_sc_hd__dfxtp_4
X_54774_ _54693_/X _54774_/X sky130_fd_sc_hd__buf_2
X_85594_ _85590_/CLK _85594_/D _85594_/Q sky130_fd_sc_hd__dfxtp_4
X_51986_ _85911_/Q _51945_/X _51985_/Y _51986_/Y sky130_fd_sc_hd__o21ai_4
X_59301_ _58766_/A _59301_/X sky130_fd_sc_hd__buf_2
X_56513_ _56523_/A _56520_/B _55823_/B _56513_/Y sky130_fd_sc_hd__nand3_4
X_87333_ _87333_/CLK _87333_/D _87333_/Q sky130_fd_sc_hd__dfxtp_4
X_53725_ _85580_/Q _53722_/X _53724_/Y _53725_/Y sky130_fd_sc_hd__o21ai_4
X_84545_ _84280_/CLK _60986_/Y _84545_/Q sky130_fd_sc_hd__dfxtp_4
X_50937_ _51074_/A _51021_/A sky130_fd_sc_hd__buf_2
X_57493_ _46542_/X _57493_/X sky130_fd_sc_hd__buf_2
X_81757_ _81783_/CLK _76121_/B _41304_/A sky130_fd_sc_hd__dfxtp_4
X_69479_ _69233_/A _69605_/A sky130_fd_sc_hd__buf_2
X_59232_ _59160_/X _85646_/Q _59205_/X _59232_/X sky130_fd_sc_hd__o21a_4
X_71510_ _71512_/A _70585_/X _71510_/Y sky130_fd_sc_hd__nand2_4
X_56444_ _56446_/A _56446_/B _56444_/C _56444_/Y sky130_fd_sc_hd__nand3_4
X_80708_ _80708_/CLK _80708_/D _80676_/D sky130_fd_sc_hd__dfxtp_4
X_41670_ _41670_/A _41670_/Y sky130_fd_sc_hd__inv_2
X_87264_ _88036_/CLK _43795_/Y _69397_/B sky130_fd_sc_hd__dfxtp_4
X_53656_ _53656_/A _74403_/B _53656_/Y sky130_fd_sc_hd__nand2_4
X_72490_ _63586_/A _72488_/B _72490_/Y sky130_fd_sc_hd__nand2_4
X_84476_ _84477_/CLK _61497_/Y _84476_/Q sky130_fd_sc_hd__dfxtp_4
X_50868_ _50228_/X _54079_/B _50868_/Y sky130_fd_sc_hd__nand2_4
X_81688_ _85003_/CLK _80162_/X _81688_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_48_0_CLK clkbuf_9_49_0_CLK/A clkbuf_9_48_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_86215_ _86213_/CLK _50369_/Y _86215_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_101 sky130_fd_sc_hd__decap_3
X_52607_ _52604_/Y _52592_/X _52606_/X _85788_/D sky130_fd_sc_hd__a21oi_4
X_40621_ _40620_/X _40621_/X sky130_fd_sc_hd__buf_2
X_59163_ _59105_/X _85748_/Q _59106_/X _59163_/X sky130_fd_sc_hd__o21a_4
X_71441_ _71238_/B _71485_/B _71444_/A sky130_fd_sc_hd__nor2_4
X_83427_ _82386_/CLK _71645_/Y _59500_/A sky130_fd_sc_hd__dfxtp_4
XPHY_112 sky130_fd_sc_hd__decap_3
X_56375_ _56458_/A _56363_/B _85217_/Q _56375_/Y sky130_fd_sc_hd__nand3_4
X_80639_ THREAD_COUNT[1] _80639_/LO sky130_fd_sc_hd__conb_1
X_87195_ _87195_/CLK _87195_/D _87195_/Q sky130_fd_sc_hd__dfxtp_4
X_53587_ _53723_/A _53601_/A sky130_fd_sc_hd__buf_2
XPHY_123 sky130_fd_sc_hd__decap_3
X_50799_ _50799_/A _50799_/B _50799_/Y sky130_fd_sc_hd__nand2_4
XPHY_134 sky130_fd_sc_hd__decap_3
X_58114_ _58112_/X _85988_/Q _58113_/X _58114_/Y sky130_fd_sc_hd__o21ai_4
XPHY_145 sky130_fd_sc_hd__decap_3
X_43340_ _41306_/X _43336_/X _87471_/Q _43337_/X _43340_/X sky130_fd_sc_hd__a2bb2o_4
X_55326_ _55310_/X _83751_/Q _55315_/X _55328_/C sky130_fd_sc_hd__nand3_4
X_86146_ _85554_/CLK _50726_/Y _86146_/Q sky130_fd_sc_hd__dfxtp_4
X_74160_ _57617_/B _74160_/B _74161_/B sky130_fd_sc_hd__xor2_4
XPHY_156 sky130_fd_sc_hd__decap_3
X_40552_ _40326_/A _86757_/Q _40591_/C _42446_/A sky130_fd_sc_hd__o21a_4
X_52538_ _52536_/Y _52486_/X _52537_/Y _85802_/D sky130_fd_sc_hd__a21boi_4
X_59094_ _59094_/A _59068_/B _59094_/Y sky130_fd_sc_hd__nor2_4
X_71372_ _71372_/A _71372_/Y sky130_fd_sc_hd__inv_2
X_83358_ _83756_/CLK _83358_/D _58548_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_3_6_0_CLK clkbuf_3_6_0_CLK/A clkbuf_3_6_1_CLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_167 sky130_fd_sc_hd__decap_3
XPHY_178 sky130_fd_sc_hd__decap_3
XPHY_189 sky130_fd_sc_hd__decap_3
X_73111_ _73104_/Y _73105_/Y _73110_/X _73121_/A sky130_fd_sc_hd__o21ai_4
X_58045_ _58043_/X _85994_/Q _58044_/X _58045_/Y sky130_fd_sc_hd__o21ai_4
X_70323_ _70328_/A _70328_/B _70323_/C _70328_/D _70323_/X sky130_fd_sc_hd__and4_4
X_82309_ _81195_/CLK _77022_/B _82309_/Q sky130_fd_sc_hd__dfxtp_4
X_43271_ _43270_/Y _43271_/Y sky130_fd_sc_hd__inv_2
X_55257_ _85033_/Q _55126_/X _55128_/X _55256_/X _55257_/X sky130_fd_sc_hd__a211o_4
X_74091_ _53567_/B _74090_/Y _74092_/B sky130_fd_sc_hd__xor2_4
X_86077_ _85757_/CLK _86077_/D _86077_/Q sky130_fd_sc_hd__dfxtp_4
X_52469_ _52467_/Y _52462_/X _52468_/Y _52469_/Y sky130_fd_sc_hd__a21boi_4
X_40483_ _40416_/A _81166_/Q _40483_/X sky130_fd_sc_hd__or2_4
X_83289_ _85536_/CLK _83289_/D _83289_/Q sky130_fd_sc_hd__dfxtp_4
X_45010_ _44975_/X _61398_/B _44995_/X _45010_/Y sky130_fd_sc_hd__o21ai_4
X_54208_ _54316_/A _54208_/X sky130_fd_sc_hd__buf_2
X_42222_ _42258_/A _42222_/X sky130_fd_sc_hd__buf_2
X_73042_ _73381_/A _73042_/B _73042_/X sky130_fd_sc_hd__and2_4
X_85028_ _85034_/CLK _85028_/D _85028_/Q sky130_fd_sc_hd__dfxtp_4
X_70254_ _70238_/X _74778_/B _70253_/X _83822_/D sky130_fd_sc_hd__a21o_4
X_55188_ _55185_/X _55187_/X _44109_/X _55188_/X sky130_fd_sc_hd__a21o_4
X_42153_ _41169_/X _42148_/X _88008_/Q _42150_/X _42153_/X sky130_fd_sc_hd__a2bb2o_4
X_54139_ _48755_/A _54249_/A sky130_fd_sc_hd__buf_2
X_77850_ _82159_/Q _77850_/B _77850_/X sky130_fd_sc_hd__xor2_4
X_70185_ _70231_/A _70200_/A sky130_fd_sc_hd__buf_2
X_59996_ _59950_/C _60091_/B sky130_fd_sc_hd__buf_2
X_41104_ _41104_/A _41104_/X sky130_fd_sc_hd__buf_2
X_76801_ _76801_/A _76801_/B _76802_/B sky130_fd_sc_hd__xor2_4
X_58947_ _58934_/X _85923_/Q _58793_/X _58947_/X sky130_fd_sc_hd__o21a_4
X_46961_ _46725_/A _46961_/X sky130_fd_sc_hd__buf_2
X_42084_ _42083_/X _42077_/X _40977_/X _88043_/Q _42078_/X _42084_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77781_ _77778_/X _77779_/Y _77780_/X _77782_/A sky130_fd_sc_hd__a21oi_4
X_74993_ _74993_/A _74993_/B _81199_/D sky130_fd_sc_hd__xor2_4
X_86979_ _87333_/CLK _44744_/Y _86979_/Q sky130_fd_sc_hd__dfxtp_4
X_48700_ _48652_/X _48146_/A _48699_/Y _74509_/A sky130_fd_sc_hd__o21ai_4
X_79520_ _79520_/A _79520_/B _79522_/A sky130_fd_sc_hd__nand2_4
X_45912_ _57673_/A _59498_/A sky130_fd_sc_hd__buf_2
X_41035_ _40991_/X _41207_/A _41034_/X _41035_/X sky130_fd_sc_hd__o21a_4
X_76732_ _76732_/A _76731_/Y _76733_/B sky130_fd_sc_hd__xnor2_4
X_49680_ _49685_/A _49669_/B _49669_/C _52895_/D _49680_/X sky130_fd_sc_hd__and4_4
X_73944_ _56548_/X _73944_/X sky130_fd_sc_hd__buf_2
X_46892_ _46892_/A _46941_/A sky130_fd_sc_hd__buf_2
X_58878_ _58877_/X _85929_/Q _58810_/X _58878_/X sky130_fd_sc_hd__o21a_4
X_48631_ _48631_/A _48632_/B sky130_fd_sc_hd__buf_2
X_79451_ _79442_/Y _79459_/A _79450_/Y _79451_/Y sky130_fd_sc_hd__a21oi_4
X_45843_ _85060_/Q _45740_/B _45843_/Y sky130_fd_sc_hd__nor2_4
X_57829_ _57718_/A _57829_/X sky130_fd_sc_hd__buf_2
X_76663_ _76663_/A _76662_/Y _76663_/Y sky130_fd_sc_hd__nand2_4
X_73875_ _73871_/X _73874_/X _73799_/X _73888_/B sky130_fd_sc_hd__a21o_4
X_78402_ _78403_/A _82709_/Q _78402_/Y sky130_fd_sc_hd__nor2_4
X_75614_ _80774_/D _75606_/A _75622_/A sky130_fd_sc_hd__nand2_4
X_60840_ _60671_/C _60675_/Y _60820_/B _60820_/A _60839_/Y _84554_/D
+ sky130_fd_sc_hd__a41oi_4
X_48562_ _86511_/Q _48536_/X _48561_/Y _48562_/Y sky130_fd_sc_hd__o21ai_4
X_72826_ _41988_/Y _72723_/X _72725_/X _72825_/Y _72826_/X sky130_fd_sc_hd__a211o_4
X_79382_ _84804_/Q _66433_/C _79382_/Y sky130_fd_sc_hd__nand2_4
X_45774_ _85129_/Q _45507_/X _45153_/A _45774_/X sky130_fd_sc_hd__o21a_4
X_76594_ _76595_/A _76595_/B _76597_/B sky130_fd_sc_hd__nor2_4
X_42986_ _42984_/X _42985_/X _40474_/X _87618_/Q _42976_/X _42986_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47513_ _47513_/A _47549_/B _47513_/C _53090_/D _47513_/X sky130_fd_sc_hd__and4_4
X_78333_ _78331_/B _78333_/Y sky130_fd_sc_hd__inv_2
X_44725_ _44725_/A _44725_/Y sky130_fd_sc_hd__inv_2
X_75545_ _75544_/X _75546_/C sky130_fd_sc_hd__inv_2
X_41937_ _41998_/A _41937_/X sky130_fd_sc_hd__buf_2
X_48493_ _48515_/A _52158_/B _48493_/Y sky130_fd_sc_hd__nand2_4
X_60771_ _63696_/A _63374_/A sky130_fd_sc_hd__buf_2
X_72757_ _72757_/A _73638_/A sky130_fd_sc_hd__buf_2
X_62510_ _61568_/B _62462_/X _62507_/X _62478_/X _62509_/X _62510_/X
+ sky130_fd_sc_hd__a41o_4
X_47444_ _47444_/A _53050_/B _47444_/Y sky130_fd_sc_hd__nand2_4
X_71708_ _71576_/X _71690_/A _71874_/D _71708_/Y sky130_fd_sc_hd__nor3_4
X_78264_ _78280_/B _78264_/Y sky130_fd_sc_hd__inv_2
X_44656_ _44638_/X _44639_/X _41081_/X _87013_/Q _44640_/X _44657_/A
+ sky130_fd_sc_hd__o32ai_4
X_63490_ _61447_/B _63487_/X _63488_/X _63489_/X _63490_/X sky130_fd_sc_hd__a211o_4
X_75476_ _75475_/Y _75477_/C sky130_fd_sc_hd__inv_2
X_41868_ _41992_/A _50731_/A sky130_fd_sc_hd__buf_2
X_72688_ _72688_/A _72697_/B sky130_fd_sc_hd__buf_2
XPHY_3 sky130_fd_sc_hd__decap_3
X_77215_ _77222_/A _77222_/B _77219_/A sky130_fd_sc_hd__xor2_4
X_62441_ _62429_/X _62435_/Y _62439_/X _84738_/Q _62440_/X _62441_/Y
+ sky130_fd_sc_hd__o32ai_4
X_43607_ _43607_/A _43607_/X sky130_fd_sc_hd__buf_2
X_74427_ _74424_/Y _74405_/X _74426_/X _74427_/Y sky130_fd_sc_hd__a21oi_4
X_40819_ _40817_/X _82294_/Q _40818_/X _40820_/A sky130_fd_sc_hd__o21ai_4
X_47375_ _86641_/Q _47332_/X _47374_/Y _47375_/Y sky130_fd_sc_hd__o21ai_4
X_71639_ _71637_/A _71228_/B _71637_/C _71639_/Y sky130_fd_sc_hd__nand3_4
X_78195_ _78192_/Y _78194_/X _78205_/A sky130_fd_sc_hd__nand2_4
X_44587_ _44587_/A _44679_/A sky130_fd_sc_hd__buf_2
X_41799_ _41799_/A _41799_/X sky130_fd_sc_hd__buf_2
X_49114_ _49109_/Y _49086_/X _49113_/X _86443_/D sky130_fd_sc_hd__a21oi_4
X_46326_ _46326_/A _50757_/B _46326_/Y sky130_fd_sc_hd__nand2_4
X_65160_ _65035_/X _85548_/Q _65036_/X _65159_/X _65160_/X sky130_fd_sc_hd__a211o_4
X_77146_ _77154_/A _77146_/B _77147_/B sky130_fd_sc_hd__xor2_4
X_43538_ _43518_/X _43523_/X _40426_/X _87369_/Q _43528_/X _43538_/Y
+ sky130_fd_sc_hd__o32ai_4
X_62372_ _62198_/Y _62406_/A sky130_fd_sc_hd__buf_2
X_74358_ _70346_/C _72699_/X _74357_/Y _83084_/D sky130_fd_sc_hd__a21bo_4
X_64111_ _59423_/Y _61003_/Y _62097_/X _60963_/X _64111_/X sky130_fd_sc_hd__a2bb2o_4
X_49045_ _53860_/B _50133_/B sky130_fd_sc_hd__buf_2
X_61323_ _61323_/A _61323_/B _61323_/X sky130_fd_sc_hd__or2_4
X_73309_ _73305_/X _73308_/X _73262_/X _73312_/A sky130_fd_sc_hd__a21o_4
X_46257_ _86752_/Q _46250_/X _46256_/Y _46257_/Y sky130_fd_sc_hd__o21ai_4
X_65091_ _64789_/A _65268_/B sky130_fd_sc_hd__buf_2
XPHY_690 sky130_fd_sc_hd__decap_3
X_77077_ _77077_/A _77086_/B _77080_/A sky130_fd_sc_hd__nand2_4
X_43469_ _43449_/X _43452_/X _41656_/X _87406_/Q _43456_/X _43470_/A
+ sky130_fd_sc_hd__o32ai_4
X_74289_ _72704_/A _74297_/A sky130_fd_sc_hd__buf_2
X_45208_ _56246_/C _45147_/X _45207_/X _45208_/Y sky130_fd_sc_hd__o21ai_4
X_76028_ _76028_/A _76028_/B _76031_/A sky130_fd_sc_hd__nand2_4
X_64042_ _84838_/Q _64091_/B _64091_/C _64091_/D _64042_/Y sky130_fd_sc_hd__nand4_4
X_61254_ _60267_/X _61254_/B _61254_/C _61254_/D _61254_/Y sky130_fd_sc_hd__nand4_4
X_46188_ _46188_/A _46114_/A _46217_/B sky130_fd_sc_hd__nor2_4
X_60205_ _60288_/C _60205_/X sky130_fd_sc_hd__buf_2
X_45139_ _55851_/B _45120_/X _45079_/X _45139_/X sky130_fd_sc_hd__o21a_4
X_68850_ _68759_/A _87232_/Q _68850_/X sky130_fd_sc_hd__and2_4
X_61185_ _61165_/A _61165_/B _61185_/C _61185_/Y sky130_fd_sc_hd__nor3_4
X_67801_ _67873_/A _67801_/B _67801_/X sky130_fd_sc_hd__and2_4
X_60136_ _60125_/A _60214_/B _60136_/C _60136_/Y sky130_fd_sc_hd__nor3_4
X_49947_ _49925_/X _49943_/B _49953_/C _53159_/D _49947_/X sky130_fd_sc_hd__and4_4
X_68781_ _68366_/X _42502_/Y _68781_/Y sky130_fd_sc_hd__nor2_4
X_65993_ _65990_/X _86235_/Q _65701_/X _65992_/X _65993_/X sky130_fd_sc_hd__a211o_4
X_77979_ _77980_/A _77972_/Y _77980_/C _77983_/A sky130_fd_sc_hd__a21o_4
X_79718_ _79715_/X _79717_/Y _79718_/X sky130_fd_sc_hd__xor2_4
X_67732_ _67658_/X _67732_/B _67732_/X sky130_fd_sc_hd__and2_4
X_64944_ _64666_/A _64944_/X sky130_fd_sc_hd__buf_2
X_60067_ _60081_/A _60081_/B _60067_/C _60067_/Y sky130_fd_sc_hd__nor3_4
X_49878_ _49875_/Y _49870_/X _49877_/X _86307_/D sky130_fd_sc_hd__a21oi_4
X_80990_ _80813_/CLK _80990_/D _80990_/Q sky130_fd_sc_hd__dfxtp_4
X_48829_ _50511_/A _48829_/B _48849_/C _48829_/X sky130_fd_sc_hd__and3_4
X_67663_ _81492_/D _67568_/X _67662_/X _67663_/X sky130_fd_sc_hd__a21bo_4
X_79649_ _79649_/A _79649_/B _79650_/B sky130_fd_sc_hd__xor2_4
X_64875_ _64858_/X _85527_/Q _64859_/X _64874_/X _64875_/X sky130_fd_sc_hd__a211o_4
X_69402_ _87020_/Q _69277_/X _69278_/X _69401_/X _69402_/X sky130_fd_sc_hd__a211o_4
X_66614_ _59802_/X _66614_/X sky130_fd_sc_hd__buf_2
X_51840_ _51820_/A _50976_/B _51840_/Y sky130_fd_sc_hd__nand2_4
X_63826_ _64172_/B _63877_/B sky130_fd_sc_hd__buf_2
X_82660_ _82596_/CLK _78330_/B _82660_/Q sky130_fd_sc_hd__dfxtp_4
X_67594_ _67120_/X _67594_/X sky130_fd_sc_hd__buf_2
X_81611_ _81632_/CLK _81611_/D _81803_/D sky130_fd_sc_hd__dfxtp_4
X_69333_ _87525_/Q _69098_/X _69124_/X _69332_/X _69333_/X sky130_fd_sc_hd__a211o_4
X_66545_ _87443_/Q _66538_/X _66540_/X _66544_/X _66545_/X sky130_fd_sc_hd__a211o_4
X_51771_ _85949_/Q _51763_/X _51770_/Y _51771_/Y sky130_fd_sc_hd__o21ai_4
X_63757_ _64223_/B _64192_/B _63757_/C _64192_/D _63757_/Y sky130_fd_sc_hd__nand4_4
X_82591_ _82671_/CLK _82623_/Q _78296_/A sky130_fd_sc_hd__dfxtp_4
X_60969_ _59831_/X _60969_/X sky130_fd_sc_hd__buf_2
X_53510_ _85623_/Q _53506_/X _53509_/Y _53510_/Y sky130_fd_sc_hd__o21ai_4
X_84330_ _84350_/CLK _63353_/Y _79158_/B sky130_fd_sc_hd__dfxtp_4
X_50722_ _86146_/Q _50654_/X _50721_/Y _50722_/Y sky130_fd_sc_hd__o21ai_4
X_62708_ _60309_/D _62708_/X sky130_fd_sc_hd__buf_2
X_81542_ _82053_/CLK _76689_/X _81542_/Q sky130_fd_sc_hd__dfxtp_4
X_69264_ _69260_/X _69263_/X _69251_/X _69264_/X sky130_fd_sc_hd__a21o_4
X_54490_ _54488_/Y _54475_/X _54489_/X _54490_/Y sky130_fd_sc_hd__a21oi_4
X_66476_ _65177_/X _66476_/B _65180_/X _66476_/Y sky130_fd_sc_hd__nand3_4
X_63688_ _63624_/X _63682_/X _63683_/X _63686_/X _63687_/Y _63688_/Y
+ sky130_fd_sc_hd__o41ai_4
X_68215_ _82050_/D _68200_/X _68214_/X _68215_/X sky130_fd_sc_hd__a21bo_4
X_53441_ _53441_/A _53817_/A sky130_fd_sc_hd__buf_2
X_65427_ _65424_/X _65426_/X _65277_/X _65427_/X sky130_fd_sc_hd__a21o_4
X_84261_ _84314_/CLK _64271_/X _79837_/B sky130_fd_sc_hd__dfxtp_4
X_50653_ _50650_/Y _50609_/X _50652_/X _50653_/Y sky130_fd_sc_hd__a21oi_4
X_62639_ _60271_/X _62910_/A sky130_fd_sc_hd__inv_2
X_81473_ _81473_/CLK _76956_/A _81473_/Q sky130_fd_sc_hd__dfxtp_4
X_69195_ _69192_/X _69194_/X _69025_/X _69195_/X sky130_fd_sc_hd__a21o_4
X_86000_ _85712_/CLK _86000_/D _86000_/Q sky130_fd_sc_hd__dfxtp_4
X_83212_ _82272_/CLK _83212_/D _79184_/B sky130_fd_sc_hd__dfxtp_4
X_56160_ _56169_/A _56150_/B _85285_/Q _56160_/Y sky130_fd_sc_hd__nand3_4
X_80424_ _80436_/A _80436_/B _80446_/B sky130_fd_sc_hd__xor2_4
X_68146_ _68144_/X _66909_/Y _68128_/X _68145_/Y _68146_/X sky130_fd_sc_hd__a211o_4
X_53372_ _53370_/Y _53355_/X _53371_/X _85646_/D sky130_fd_sc_hd__a21oi_4
X_65358_ _65252_/X _83284_/Q _65230_/X _65357_/X _65358_/X sky130_fd_sc_hd__a211o_4
X_84192_ _84192_/CLK _84192_/D _84192_/Q sky130_fd_sc_hd__dfxtp_4
X_50584_ _48928_/A _50560_/X _50568_/C _50584_/X sky130_fd_sc_hd__and3_4
X_55111_ _85316_/Q _55098_/X _55110_/Y _55111_/Y sky130_fd_sc_hd__o21ai_4
X_52323_ _52515_/A _52324_/A sky130_fd_sc_hd__buf_2
X_64309_ _64287_/A _58535_/A _64287_/C _64309_/Y sky130_fd_sc_hd__nand3_4
X_83143_ _83115_/CLK _83143_/D _70121_/A sky130_fd_sc_hd__dfxtp_4
X_80355_ _80353_/Y _80354_/Y _80355_/X sky130_fd_sc_hd__xor2_4
X_68077_ _68077_/A _68077_/B _68077_/Y sky130_fd_sc_hd__nand2_4
X_56091_ _55993_/Y _55994_/X _56098_/A _56091_/X sky130_fd_sc_hd__and3_4
X_65289_ _65289_/A _65289_/B _65289_/X sky130_fd_sc_hd__and2_4
X_55042_ _85329_/Q _55020_/X _55041_/Y _55042_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_6_30_0_CLK clkbuf_6_31_0_CLK/A clkbuf_7_61_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_67028_ _67028_/A _67028_/B _67028_/X sky130_fd_sc_hd__and2_4
X_52254_ _52251_/Y _52232_/X _52253_/X _85859_/D sky130_fd_sc_hd__a21oi_4
X_83074_ _85593_/CLK _74402_/Y _83074_/Q sky130_fd_sc_hd__dfxtp_4
X_87951_ _87950_/CLK _42264_/X _87951_/Q sky130_fd_sc_hd__dfxtp_4
X_80286_ _80280_/Y _80286_/B _80288_/B sky130_fd_sc_hd__nand2_4
X_51205_ _51184_/X _47174_/X _51205_/Y sky130_fd_sc_hd__nand2_4
X_86902_ _83022_/CLK _45055_/Y _64320_/B sky130_fd_sc_hd__dfxtp_4
X_82025_ _81989_/CLK _77792_/B _81993_/D sky130_fd_sc_hd__dfxtp_4
X_59850_ _59687_/A _59683_/A _59666_/A _59850_/Y sky130_fd_sc_hd__a21oi_4
X_52185_ _52185_/A _52185_/X sky130_fd_sc_hd__buf_2
X_87882_ _87883_/CLK _87882_/D _87882_/Q sky130_fd_sc_hd__dfxtp_4
X_58801_ _86703_/Q _58764_/B _58801_/Y sky130_fd_sc_hd__nor2_4
X_51136_ _51191_/A _51160_/A sky130_fd_sc_hd__buf_2
X_86833_ _88398_/CLK _86833_/D _66700_/B sky130_fd_sc_hd__dfxtp_4
X_59781_ _69814_/A _70056_/A sky130_fd_sc_hd__buf_2
X_56993_ _56737_/X _57149_/C _56735_/X _56994_/D _56726_/X _56993_/X
+ sky130_fd_sc_hd__a41o_4
X_68979_ _68517_/A _68979_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_554_0_CLK clkbuf_9_277_0_CLK/X _87472_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_45_0_CLK clkbuf_6_45_0_CLK/A clkbuf_7_91_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_58732_ _58703_/X _85460_/Q _58731_/X _58732_/Y sky130_fd_sc_hd__o21ai_4
X_51067_ _51056_/A _51071_/B _51071_/C _52758_/D _51067_/X sky130_fd_sc_hd__and4_4
X_55944_ _44989_/A _55619_/A _44102_/A _55943_/X _55945_/B sky130_fd_sc_hd__a211o_4
X_86764_ _80657_/CLK _46185_/X _86764_/Q sky130_fd_sc_hd__dfxtp_4
X_71990_ _71988_/Y _71969_/X _71989_/Y _71990_/Y sky130_fd_sc_hd__a21boi_4
X_83976_ _80961_/CLK _68413_/X _83976_/Q sky130_fd_sc_hd__dfxtp_4
X_50018_ _50027_/A _53232_/B _50018_/Y sky130_fd_sc_hd__nand2_4
X_85715_ _84766_/CLK _53004_/Y _85715_/Q sky130_fd_sc_hd__dfxtp_4
X_70941_ _51235_/B _70937_/X _70940_/Y _83657_/D sky130_fd_sc_hd__o21ai_4
X_58663_ _84809_/Q _58663_/Y sky130_fd_sc_hd__inv_2
X_82927_ _82933_/CLK _78226_/X _46459_/A sky130_fd_sc_hd__dfxtp_4
X_55875_ _56223_/C _44064_/X _44049_/X _55874_/X _55875_/X sky130_fd_sc_hd__a211o_4
X_86695_ _86695_/CLK _86695_/D _86695_/Q sky130_fd_sc_hd__dfxtp_4
X_57614_ _57612_/Y _57581_/X _57613_/Y _57614_/Y sky130_fd_sc_hd__a21boi_4
X_42840_ _42839_/Y _87692_/D sky130_fd_sc_hd__inv_2
X_54826_ _54824_/Y _54802_/X _54825_/X _54826_/Y sky130_fd_sc_hd__a21oi_4
X_85646_ _85648_/CLK _85646_/D _85646_/Q sky130_fd_sc_hd__dfxtp_4
X_73660_ _73605_/X _86237_/Q _44194_/X _73659_/X _73660_/X sky130_fd_sc_hd__a211o_4
X_58594_ _58928_/A _58594_/X sky130_fd_sc_hd__buf_2
X_70872_ _51812_/B _70855_/X _70871_/Y _70872_/Y sky130_fd_sc_hd__o21ai_4
X_82858_ _82855_/CLK _82858_/D _40888_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_569_0_CLK clkbuf_9_284_0_CLK/X _88376_/CLK sky130_fd_sc_hd__clkbuf_1
X_72611_ _83217_/Q _72590_/X _72585_/A _72610_/X _72611_/X sky130_fd_sc_hd__o22a_4
X_57545_ _57542_/Y _57543_/X _57544_/Y _57545_/Y sky130_fd_sc_hd__a21boi_4
X_81809_ _81260_/CLK _81809_/D _47378_/A sky130_fd_sc_hd__dfxtp_4
X_42771_ _41312_/X _42767_/X _67451_/B _42768_/X _42771_/X sky130_fd_sc_hd__a2bb2o_4
X_88365_ _83139_/CLK _40618_/X _88365_/Q sky130_fd_sc_hd__dfxtp_4
X_54757_ _54729_/A _54757_/X sky130_fd_sc_hd__buf_2
X_73591_ _73591_/A _73591_/B _73591_/X sky130_fd_sc_hd__xor2_4
X_85577_ _83564_/CLK _53744_/Y _85577_/Q sky130_fd_sc_hd__dfxtp_4
X_51969_ _51967_/Y _51934_/X _51968_/Y _85915_/D sky130_fd_sc_hd__a21boi_4
X_82789_ _82792_/CLK _82821_/Q _82789_/Q sky130_fd_sc_hd__dfxtp_4
X_44510_ _41281_/Y _44502_/X _87072_/Q _44503_/X _87072_/D sky130_fd_sc_hd__a2bb2o_4
X_75330_ _81076_/Q _75330_/Y sky130_fd_sc_hd__inv_2
X_87316_ _88084_/CLK _43677_/Y _87316_/Q sky130_fd_sc_hd__dfxtp_4
X_53708_ _53706_/Y _53696_/X _53707_/Y _85584_/D sky130_fd_sc_hd__a21boi_4
X_41722_ _41799_/A _41722_/X sky130_fd_sc_hd__buf_2
X_72542_ _72579_/B _72516_/C _72506_/C _72584_/A sky130_fd_sc_hd__nand3_4
X_84528_ _84400_/CLK _61050_/X _76976_/A sky130_fd_sc_hd__dfxtp_4
X_45490_ _85051_/Q _45490_/B _45490_/Y sky130_fd_sc_hd__nor2_4
X_57476_ _74139_/A _57067_/Y _57465_/A _56892_/B _57476_/X sky130_fd_sc_hd__a211o_4
X_88296_ _87790_/CLK _40997_/Y _88296_/Q sky130_fd_sc_hd__dfxtp_4
X_54688_ _85396_/Q _54676_/X _54687_/Y _54688_/Y sky130_fd_sc_hd__o21ai_4
X_59215_ _59204_/Y _59145_/X _59211_/X _59214_/X _84760_/D sky130_fd_sc_hd__a22oi_4
X_44441_ _44425_/X _44427_/X _41616_/X _87106_/Q _44428_/X _44441_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56427_ _56431_/A _56433_/B _85198_/Q _56427_/Y sky130_fd_sc_hd__nand3_4
X_75261_ _75261_/A _75261_/B _75279_/B sky130_fd_sc_hd__xor2_4
X_41653_ _40586_/A _41653_/X sky130_fd_sc_hd__buf_2
X_87247_ _87766_/CLK _43828_/X _87247_/Q sky130_fd_sc_hd__dfxtp_4
X_53639_ _85597_/Q _53610_/X _53638_/Y _53639_/Y sky130_fd_sc_hd__o21ai_4
X_72473_ _57800_/X _72471_/Y _72472_/Y _64761_/B _59833_/X _72473_/X
+ sky130_fd_sc_hd__o32a_4
X_84459_ _84469_/CLK _84459_/D _61690_/C sky130_fd_sc_hd__dfxtp_4
X_77000_ _84552_/Q _84424_/Q _77000_/X sky130_fd_sc_hd__xor2_4
X_74212_ _74232_/A _85893_/Q _74212_/X sky130_fd_sc_hd__and2_4
X_40604_ _40601_/X _81149_/Q _40603_/X _40604_/X sky130_fd_sc_hd__o21a_4
X_47160_ _86664_/Q _47145_/X _47159_/Y _47160_/Y sky130_fd_sc_hd__o21ai_4
X_59146_ _58858_/A _59146_/X sky130_fd_sc_hd__buf_2
X_71424_ _70407_/C _71432_/B _71424_/C _71365_/X _71424_/X sky130_fd_sc_hd__and4_4
X_44372_ _44372_/A _44372_/Y sky130_fd_sc_hd__inv_2
X_56358_ _56358_/A _56358_/B _55702_/B _56358_/Y sky130_fd_sc_hd__nand3_4
X_75192_ _75133_/Y _75147_/Y _75163_/X _75182_/A _75192_/Y sky130_fd_sc_hd__nand4_4
X_87178_ _87178_/CLK _87178_/D _87178_/Q sky130_fd_sc_hd__dfxtp_4
X_41584_ _41584_/A _41584_/B _41584_/X sky130_fd_sc_hd__or2_4
X_46111_ _46111_/A _46111_/B _46099_/X _46094_/X _46111_/X sky130_fd_sc_hd__or4_4
X_55309_ _44110_/X _55309_/X sky130_fd_sc_hd__buf_2
X_43323_ _41259_/X _43300_/X _87481_/Q _43302_/X _87481_/D sky130_fd_sc_hd__a2bb2o_4
X_74143_ _74143_/A _72795_/A _74143_/Y sky130_fd_sc_hd__nor2_4
X_86129_ _85527_/CLK _50809_/Y _86129_/Q sky130_fd_sc_hd__dfxtp_4
X_40535_ _40414_/X _40937_/A sky130_fd_sc_hd__buf_2
X_47091_ _46903_/A _47091_/X sky130_fd_sc_hd__buf_2
X_59077_ _84771_/Q _59043_/X _59069_/X _59076_/X _84771_/D sky130_fd_sc_hd__a2bb2oi_4
X_71355_ _71344_/X _83528_/Q _71354_/X _83528_/D sky130_fd_sc_hd__a21o_4
X_56289_ _56282_/Y _56360_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_507_0_CLK clkbuf_9_253_0_CLK/X _85786_/CLK sky130_fd_sc_hd__clkbuf_1
X_46042_ _41506_/Y _46029_/X _66785_/B _46030_/X _86797_/D sky130_fd_sc_hd__a2bb2o_4
X_58028_ _58098_/A _58028_/X sky130_fd_sc_hd__buf_2
X_70306_ _70296_/X _70297_/X _70306_/C _70301_/D _70306_/X sky130_fd_sc_hd__and4_4
X_43254_ _41064_/X _43247_/X _87516_/Q _43248_/X _87516_/D sky130_fd_sc_hd__a2bb2o_4
X_78951_ _78938_/A _78946_/A _78951_/X sky130_fd_sc_hd__and2_4
X_74074_ _87325_/Q _74073_/X _74074_/Y sky130_fd_sc_hd__nor2_4
X_40466_ _40932_/A _40467_/B sky130_fd_sc_hd__buf_2
X_71286_ _53219_/B _71264_/X _71285_/Y _71286_/Y sky130_fd_sc_hd__o21ai_4
X_42205_ _42204_/X _42205_/X sky130_fd_sc_hd__buf_2
X_77902_ _77902_/A _77902_/B _77902_/X sky130_fd_sc_hd__or2_4
X_73025_ _72771_/A _73530_/B sky130_fd_sc_hd__buf_2
X_70237_ _70224_/X _74755_/B _70236_/X _83827_/D sky130_fd_sc_hd__a21o_4
X_43185_ _43185_/A _43185_/X sky130_fd_sc_hd__buf_2
X_78882_ _82730_/Q _78882_/B _82698_/D sky130_fd_sc_hd__xor2_4
X_40397_ _40396_/Y _40397_/Y sky130_fd_sc_hd__inv_2
X_49801_ _57952_/B _49798_/X _49800_/Y _49801_/Y sky130_fd_sc_hd__o21ai_4
X_42136_ _51584_/A _42137_/A sky130_fd_sc_hd__buf_2
X_77833_ _82270_/Q _77833_/B _77833_/Y sky130_fd_sc_hd__xnor2_4
X_70168_ _70337_/A _70209_/A sky130_fd_sc_hd__buf_2
X_47993_ _57567_/A _50308_/A sky130_fd_sc_hd__buf_2
X_59979_ _59978_/Y _59979_/Y sky130_fd_sc_hd__inv_2
X_49732_ _49787_/A _49732_/X sky130_fd_sc_hd__buf_2
X_46944_ _46915_/X _46944_/B _46926_/C _52763_/D _46944_/X sky130_fd_sc_hd__and4_4
X_42067_ _42052_/X _42043_/X _40950_/X _88049_/Q _42044_/X _42067_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77764_ _77756_/Y _77764_/B _77764_/Y sky130_fd_sc_hd__nand2_4
X_62990_ _63713_/A _60159_/A _60212_/A _63348_/A _60304_/A _62990_/Y
+ sky130_fd_sc_hd__o32ai_4
X_70099_ _83134_/Q _70099_/Y sky130_fd_sc_hd__inv_2
X_74976_ _74972_/Y _74975_/X _74988_/A sky130_fd_sc_hd__nand2_4
X_79503_ _79503_/A _79503_/B _79504_/B sky130_fd_sc_hd__xnor2_4
X_41018_ _41018_/A _41018_/Y sky130_fd_sc_hd__inv_2
X_76715_ _81690_/Q _76715_/B _76715_/Y sky130_fd_sc_hd__xnor2_4
X_61941_ _61879_/A _61935_/Y _61938_/Y _61940_/Y _61941_/Y sky130_fd_sc_hd__nand4_4
X_49663_ _86346_/Q _49660_/X _49662_/Y _49663_/Y sky130_fd_sc_hd__o21ai_4
X_73927_ _44126_/X _73927_/B _73927_/X sky130_fd_sc_hd__and2_4
X_46875_ _54417_/D _52724_/D sky130_fd_sc_hd__buf_2
X_77695_ _77695_/A _77695_/B _77703_/A sky130_fd_sc_hd__or2_4
X_48614_ _48614_/A _48615_/A sky130_fd_sc_hd__inv_2
X_79434_ _58663_/Y _66407_/C _79433_/Y _79438_/A sky130_fd_sc_hd__o21a_4
X_45826_ _57473_/B _45826_/Y sky130_fd_sc_hd__inv_2
X_64660_ _64655_/X _64633_/B _64659_/X _64660_/Y sky130_fd_sc_hd__nand3_4
X_76646_ _81474_/Q _76648_/A sky130_fd_sc_hd__inv_2
X_49594_ _49580_/X _52807_/B _49594_/Y sky130_fd_sc_hd__nand2_4
X_61872_ _57656_/X _61824_/X _61838_/X _61870_/X _61871_/X _61872_/X
+ sky130_fd_sc_hd__a41o_4
X_73858_ _73853_/X _73856_/X _73857_/X _73863_/A sky130_fd_sc_hd__a21o_4
X_63611_ _63611_/A _63630_/B _63630_/C _63611_/Y sky130_fd_sc_hd__nor3_4
X_48545_ _48545_/A _48610_/C sky130_fd_sc_hd__buf_2
X_60823_ _61202_/A _63374_/A _61277_/B _60820_/Y _60822_/X _60823_/Y
+ sky130_fd_sc_hd__o41ai_4
X_72809_ _73535_/A _65455_/B _72809_/X sky130_fd_sc_hd__and2_4
X_79365_ _79361_/X _79364_/Y _79365_/X sky130_fd_sc_hd__xor2_4
X_45757_ _45757_/A _45757_/X sky130_fd_sc_hd__buf_2
X_64591_ _64829_/A _64591_/X sky130_fd_sc_hd__buf_2
X_76577_ _76576_/B _76575_/Y _76572_/Y _76577_/Y sky130_fd_sc_hd__o21ai_4
X_42969_ _40554_/X _43774_/A sky130_fd_sc_hd__buf_2
X_73789_ _73789_/A _73789_/B _73789_/Y sky130_fd_sc_hd__nand2_4
X_66330_ _66294_/X _66328_/Y _66329_/Y _66330_/Y sky130_fd_sc_hd__o21ai_4
X_78316_ _78316_/A _82659_/D _78335_/B sky130_fd_sc_hd__nand2_4
X_44708_ _43047_/A _44708_/X sky130_fd_sc_hd__buf_2
X_75528_ _75528_/A _75528_/B _75528_/X sky130_fd_sc_hd__xor2_4
X_63542_ _63495_/X _63533_/X _63534_/X _63538_/X _63541_/Y _63542_/Y
+ sky130_fd_sc_hd__o41ai_4
X_48476_ _50447_/A _48489_/B _48476_/C _48476_/X sky130_fd_sc_hd__and3_4
X_60754_ _60820_/A _60702_/Y _60754_/X sky130_fd_sc_hd__and2_4
X_79296_ _79275_/B _79292_/X _79295_/Y _79296_/Y sky130_fd_sc_hd__a21oi_4
X_45688_ _85102_/Q _45688_/Y sky130_fd_sc_hd__inv_2
X_47427_ _47418_/A _47415_/X _47466_/C _53044_/D _47427_/X sky130_fd_sc_hd__and4_4
X_66261_ _66179_/X _66258_/Y _66260_/Y _66261_/Y sky130_fd_sc_hd__o21ai_4
X_78247_ _78247_/A _78247_/B _78247_/X sky130_fd_sc_hd__xor2_4
X_44639_ _44567_/A _44639_/X sky130_fd_sc_hd__buf_2
X_63473_ _58541_/A _63436_/X _61440_/A _63437_/X _63473_/X sky130_fd_sc_hd__a2bb2o_4
X_75459_ _75457_/B _75457_/C _75457_/A _75509_/C sky130_fd_sc_hd__o21ai_4
X_60685_ _84584_/Q _60673_/X _60675_/Y _60684_/X _60685_/Y sky130_fd_sc_hd__a2bb2oi_4
X_68000_ _68044_/A _68000_/B _68000_/X sky130_fd_sc_hd__and2_4
X_65212_ _65718_/A _65212_/X sky130_fd_sc_hd__buf_2
X_62424_ _61499_/B _62390_/X _62363_/X _62407_/X _62423_/X _62424_/X
+ sky130_fd_sc_hd__a41o_4
X_47358_ _47354_/Y _47317_/X _47357_/X _86643_/D sky130_fd_sc_hd__a21oi_4
X_66192_ _84150_/Q _66193_/C sky130_fd_sc_hd__inv_2
X_78178_ _78177_/A _78177_/B _78178_/Y sky130_fd_sc_hd__nand2_4
X_46309_ _46450_/A _53511_/A sky130_fd_sc_hd__buf_2
X_65143_ _65140_/Y _65070_/X _65142_/Y _65143_/X sky130_fd_sc_hd__a21o_4
X_77129_ _77120_/Y _77127_/Y _77128_/Y _77129_/X sky130_fd_sc_hd__o21a_4
X_62355_ _62193_/A _62355_/X sky130_fd_sc_hd__buf_2
X_47289_ _54130_/B _52965_/B sky130_fd_sc_hd__buf_2
X_49028_ _46349_/A _49029_/B sky130_fd_sc_hd__buf_2
X_61306_ _61306_/A _72503_/A sky130_fd_sc_hd__buf_2
X_80140_ _80135_/X _80139_/Y _81686_/D sky130_fd_sc_hd__xor2_4
X_65074_ _65074_/A _65074_/B _65074_/X sky130_fd_sc_hd__and2_4
X_69951_ _69948_/X _69950_/X _69951_/Y sky130_fd_sc_hd__nand2_4
X_62286_ _62285_/X _62286_/X sky130_fd_sc_hd__buf_2
X_68902_ _68994_/A _88254_/Q _68902_/X sky130_fd_sc_hd__and2_4
X_64025_ _63217_/B _64118_/B _64040_/C _64025_/D _64025_/Y sky130_fd_sc_hd__nand4_4
X_61237_ _60296_/X _61188_/B _61188_/C _61237_/D _61237_/Y sky130_fd_sc_hd__nand4_4
X_80071_ _80071_/A _80070_/Y _80071_/X sky130_fd_sc_hd__xor2_4
X_69882_ _69882_/A _69883_/B sky130_fd_sc_hd__inv_2
X_68833_ _68785_/A _88353_/Q _68833_/X sky130_fd_sc_hd__and2_4
X_61168_ _72527_/A _72527_/B _84515_/Q _61167_/Y _61117_/X _84515_/D
+ sky130_fd_sc_hd__a32o_4
X_60119_ _60118_/X _60119_/Y sky130_fd_sc_hd__inv_2
X_83830_ _83191_/CLK _83830_/D _83830_/Q sky130_fd_sc_hd__dfxtp_4
X_68764_ _87088_/Q _68707_/X _68762_/X _68763_/X _68764_/X sky130_fd_sc_hd__a211o_4
X_53990_ _53990_/A _53991_/A sky130_fd_sc_hd__buf_2
X_65976_ _65976_/A _65976_/X sky130_fd_sc_hd__buf_2
X_61099_ _61172_/A _61230_/C sky130_fd_sc_hd__buf_2
X_67715_ _87907_/Q _67713_/X _67641_/X _67714_/X _67715_/X sky130_fd_sc_hd__a211o_4
X_52941_ _85726_/Q _52929_/X _52940_/Y _52941_/Y sky130_fd_sc_hd__o21ai_4
X_64927_ _64776_/A _64927_/X sky130_fd_sc_hd__buf_2
X_83761_ _83761_/CLK _83761_/D _83761_/Q sky130_fd_sc_hd__dfxtp_4
X_80973_ _81065_/CLK _75675_/X _80961_/D sky130_fd_sc_hd__dfxtp_4
X_68695_ _69661_/A _68695_/B _68695_/Y sky130_fd_sc_hd__nor2_4
X_85500_ _85499_/CLK _85500_/D _85500_/Q sky130_fd_sc_hd__dfxtp_4
X_82712_ _82803_/CLK _79011_/X _82668_/D sky130_fd_sc_hd__dfxtp_4
X_55660_ _55652_/Y _55654_/X _55659_/Y _55660_/Y sky130_fd_sc_hd__a21oi_4
X_67646_ _67643_/X _67645_/X _67619_/X _67649_/A sky130_fd_sc_hd__a21o_4
X_86480_ _86191_/CLK _48802_/Y _86480_/Q sky130_fd_sc_hd__dfxtp_4
X_52872_ _52867_/A _52853_/B _52872_/C _52872_/D _52872_/X sky130_fd_sc_hd__and4_4
X_64858_ _64678_/A _64858_/X sky130_fd_sc_hd__buf_2
X_83692_ _85635_/CLK _83692_/D _47194_/A sky130_fd_sc_hd__dfxtp_4
X_54611_ _54558_/A _54611_/X sky130_fd_sc_hd__buf_2
X_85431_ _85431_/CLK _54499_/Y _85431_/Q sky130_fd_sc_hd__dfxtp_4
X_51823_ _51823_/A _51823_/X sky130_fd_sc_hd__buf_2
X_63809_ _63809_/A _63804_/Y _63805_/Y _63809_/D _63809_/X sky130_fd_sc_hd__and4_4
X_82643_ _84003_/CLK _82643_/D _82643_/Q sky130_fd_sc_hd__dfxtp_4
X_67577_ _67577_/A _67577_/B _67577_/Y sky130_fd_sc_hd__nand2_4
X_55591_ _83005_/Q _55617_/A _44099_/X _55590_/X _55592_/B sky130_fd_sc_hd__a211o_4
X_64789_ _64789_/A _64913_/B sky130_fd_sc_hd__buf_2
X_57330_ _57330_/A _57330_/Y sky130_fd_sc_hd__inv_2
X_69316_ _69286_/A _87782_/Q _69316_/X sky130_fd_sc_hd__and2_4
X_88150_ _87436_/CLK _88150_/D _88150_/Q sky130_fd_sc_hd__dfxtp_4
X_54542_ _54546_/A _53364_/B _54542_/Y sky130_fd_sc_hd__nand2_4
X_66528_ _68386_/A _69315_/A sky130_fd_sc_hd__buf_2
X_85362_ _86289_/CLK _54875_/Y _85362_/Q sky130_fd_sc_hd__dfxtp_4
X_51754_ _52679_/A _51781_/A sky130_fd_sc_hd__buf_2
X_82574_ _82575_/CLK _82606_/Q _78161_/A sky130_fd_sc_hd__dfxtp_4
X_87101_ _88288_/CLK _44457_/Y _87101_/Q sky130_fd_sc_hd__dfxtp_4
X_84313_ _84314_/CLK _84313_/D _80455_/B sky130_fd_sc_hd__dfxtp_4
X_50705_ _50703_/Y _50699_/X _50704_/Y _50705_/Y sky130_fd_sc_hd__a21boi_4
X_57261_ _44287_/X _57261_/X sky130_fd_sc_hd__buf_2
X_81525_ _82053_/CLK _81525_/D _81525_/Q sky130_fd_sc_hd__dfxtp_4
X_69247_ _88043_/Q _69217_/X _69245_/X _69246_/X _69247_/X sky130_fd_sc_hd__a211o_4
X_88081_ _88081_/CLK _41987_/Y _88081_/Q sky130_fd_sc_hd__dfxtp_4
X_54473_ _54478_/A _54473_/B _54473_/Y sky130_fd_sc_hd__nand2_4
X_66459_ _65078_/X _66518_/B _65080_/X _66459_/Y sky130_fd_sc_hd__nand3_4
X_85293_ _85257_/CLK _85293_/D _85293_/Q sky130_fd_sc_hd__dfxtp_4
X_51685_ _51682_/Y _51667_/X _51684_/X _51685_/Y sky130_fd_sc_hd__a21oi_4
X_59000_ _58925_/X _85441_/Q _58999_/X _59000_/Y sky130_fd_sc_hd__o21ai_4
X_56212_ _56040_/X _56210_/X _56211_/Y _56212_/Y sky130_fd_sc_hd__o21ai_4
X_87032_ _87032_/CLK _87032_/D _87032_/Q sky130_fd_sc_hd__dfxtp_4
X_53424_ _53420_/A _53402_/B _53410_/C _51220_/D _53424_/X sky130_fd_sc_hd__and4_4
X_84244_ _84241_/CLK _64463_/Y _79658_/B sky130_fd_sc_hd__dfxtp_4
X_50636_ _50627_/X _52338_/B _50636_/Y sky130_fd_sc_hd__nand2_4
X_81456_ _81492_/CLK _76783_/B _81456_/Q sky130_fd_sc_hd__dfxtp_4
X_57192_ _57192_/A _85065_/Q _57195_/B sky130_fd_sc_hd__nand2_4
X_69178_ _69178_/A _69179_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_4 _44267_/A _44284_/C sky130_fd_sc_hd__buf_2
X_80407_ _80394_/X _80405_/X _80406_/X _80407_/Y sky130_fd_sc_hd__a21oi_4
X_56143_ _56117_/B _56143_/B _56144_/A sky130_fd_sc_hd__xnor2_4
X_68129_ _68129_/A _68129_/X sky130_fd_sc_hd__buf_2
X_53355_ _53355_/A _53355_/X sky130_fd_sc_hd__buf_2
X_84175_ _84175_/CLK _65832_/X _84175_/Q sky130_fd_sc_hd__dfxtp_4
X_50567_ _50538_/A _50568_/C sky130_fd_sc_hd__buf_2
X_81387_ _81322_/CLK _83923_/Q _76874_/B sky130_fd_sc_hd__dfxtp_4
X_40320_ _40326_/A _40321_/A sky130_fd_sc_hd__inv_2
X_52306_ _52304_/Y _52289_/X _52305_/X _85849_/D sky130_fd_sc_hd__a21oi_4
X_71140_ _70716_/A _71152_/C sky130_fd_sc_hd__buf_2
X_83126_ _83145_/CLK _83126_/D _83126_/Q sky130_fd_sc_hd__dfxtp_4
X_56074_ _56073_/Y _56074_/X sky130_fd_sc_hd__buf_2
X_80338_ _80320_/Y _80322_/B _80320_/A _80338_/Y sky130_fd_sc_hd__o21ai_4
X_53286_ _53276_/A _54464_/B _53286_/Y sky130_fd_sc_hd__nand2_4
X_50498_ _50495_/Y _50491_/X _50497_/X _86189_/D sky130_fd_sc_hd__a21oi_4
X_59902_ _60122_/A _59901_/Y _60122_/C _59903_/A sky130_fd_sc_hd__nand3_4
X_55025_ _54973_/A _55026_/C sky130_fd_sc_hd__buf_2
X_52237_ _48667_/A _52248_/B _52223_/C _52237_/X sky130_fd_sc_hd__and3_4
X_71071_ _71071_/A _71078_/A sky130_fd_sc_hd__buf_2
X_83057_ _85566_/CLK _83057_/D _83057_/Q sky130_fd_sc_hd__dfxtp_4
X_87934_ _82886_/CLK _87934_/D _87934_/Q sky130_fd_sc_hd__dfxtp_4
X_80269_ _80266_/Y _80268_/Y _80636_/A sky130_fd_sc_hd__nand2_4
Xclkbuf_10_493_0_CLK clkbuf_9_246_0_CLK/X _86398_/CLK sky130_fd_sc_hd__clkbuf_1
X_70022_ _83871_/Q _70010_/X _70021_/Y _70022_/X sky130_fd_sc_hd__a21bo_4
X_82008_ _82008_/CLK _82040_/Q _77174_/B sky130_fd_sc_hd__dfxtp_4
X_59833_ _65044_/A _59833_/X sky130_fd_sc_hd__buf_2
X_52168_ _52168_/A _50466_/B _52168_/Y sky130_fd_sc_hd__nand2_4
X_87865_ _87865_/CLK _87865_/D _87865_/Q sky130_fd_sc_hd__dfxtp_4
X_51119_ _51039_/A _51119_/X sky130_fd_sc_hd__buf_2
X_74830_ _74829_/Y _80658_/D sky130_fd_sc_hd__inv_2
X_86816_ _86784_/CLK _46011_/Y _67107_/B sky130_fd_sc_hd__dfxtp_4
X_59764_ _59722_/A _59765_/A sky130_fd_sc_hd__buf_2
X_44990_ _44990_/A _45033_/B _44990_/Y sky130_fd_sc_hd__nand2_4
X_52099_ _52096_/Y _52049_/X _52098_/X _85889_/D sky130_fd_sc_hd__a21oi_4
X_56976_ _56985_/D _56976_/X sky130_fd_sc_hd__buf_2
X_87796_ _88085_/CLK _42625_/Y _73527_/A sky130_fd_sc_hd__dfxtp_4
X_58715_ _64679_/A _58847_/A sky130_fd_sc_hd__buf_2
X_43941_ _45964_/A _43941_/X sky130_fd_sc_hd__buf_2
X_55927_ _55926_/X _55927_/X sky130_fd_sc_hd__buf_2
X_74761_ _70325_/Y _71012_/B _74760_/Y _74761_/Y sky130_fd_sc_hd__o21ai_4
X_86747_ _85822_/CLK _46332_/Y _86747_/Q sky130_fd_sc_hd__dfxtp_4
X_71973_ _83310_/Q _57635_/X _71972_/Y _71973_/Y sky130_fd_sc_hd__o21ai_4
X_59695_ _59691_/X _62183_/A _59631_/Y _59695_/Y sky130_fd_sc_hd__o21ai_4
X_83959_ _80991_/CLK _68837_/X _83959_/Q sky130_fd_sc_hd__dfxtp_4
X_76500_ _76500_/A _76499_/X _76500_/X sky130_fd_sc_hd__xor2_4
X_73712_ _73609_/X _85627_/Q _73661_/X _73711_/X _73712_/X sky130_fd_sc_hd__a211o_4
X_46660_ _46652_/Y _46654_/X _46659_/X _86717_/D sky130_fd_sc_hd__a21oi_4
X_58646_ _58939_/A _58646_/X sky130_fd_sc_hd__buf_2
X_70924_ _51037_/B _70909_/X _70923_/Y _83661_/D sky130_fd_sc_hd__o21ai_4
X_77480_ _77479_/X _77480_/Y sky130_fd_sc_hd__inv_2
X_43872_ _41259_/X _43868_/X _69011_/B _43870_/X _87225_/D sky130_fd_sc_hd__a2bb2o_4
X_55858_ _56414_/C _55489_/A _55512_/X _55857_/X _55858_/X sky130_fd_sc_hd__a211o_4
X_74692_ _74675_/X _56873_/X _74691_/Y _74693_/A sky130_fd_sc_hd__o21ai_4
X_86678_ _86359_/CLK _86678_/D _59131_/A sky130_fd_sc_hd__dfxtp_4
X_45611_ _45611_/A _55470_/B sky130_fd_sc_hd__inv_2
X_76431_ _76430_/B _76430_/C _76430_/A _76431_/Y sky130_fd_sc_hd__o21ai_4
X_54809_ _54889_/A _54831_/C sky130_fd_sc_hd__buf_2
X_42823_ _41447_/X _42821_/X _87701_/Q _42822_/X _42823_/X sky130_fd_sc_hd__a2bb2o_4
X_73643_ _73643_/A _73642_/X _73644_/B sky130_fd_sc_hd__nand2_4
X_85629_ _86237_/CLK _85629_/D _85629_/Q sky130_fd_sc_hd__dfxtp_4
X_70855_ _70855_/A _70855_/X sky130_fd_sc_hd__buf_2
X_46591_ _46591_/A _54087_/B sky130_fd_sc_hd__buf_2
X_58577_ _58577_/A _58614_/B _58577_/Y sky130_fd_sc_hd__nor2_4
X_55789_ _45244_/A _55306_/X _55172_/X _55788_/X _55790_/B sky130_fd_sc_hd__a211o_4
X_48330_ _48348_/A _50372_/B _48330_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_431_0_CLK clkbuf_9_215_0_CLK/X _84177_/CLK sky130_fd_sc_hd__clkbuf_1
X_79150_ _79150_/A _79150_/B _82458_/D sky130_fd_sc_hd__xor2_4
X_45542_ _85144_/Q _45464_/X _44964_/X _45542_/Y sky130_fd_sc_hd__o21ai_4
X_57528_ _46366_/A _57528_/X sky130_fd_sc_hd__buf_2
X_76362_ _76355_/Y _76361_/Y _76363_/B sky130_fd_sc_hd__xor2_4
X_42754_ _41259_/X _42745_/X _69008_/B _42746_/X _42754_/X sky130_fd_sc_hd__a2bb2o_4
X_88348_ _87851_/CLK _40721_/X _88348_/Q sky130_fd_sc_hd__dfxtp_4
X_73574_ _83145_/Q _73549_/X _73573_/Y _83145_/D sky130_fd_sc_hd__a21o_4
X_70786_ _70786_/A _70873_/A sky130_fd_sc_hd__buf_2
X_78101_ _82661_/Q _78101_/B _78101_/X sky130_fd_sc_hd__xor2_4
X_75313_ _75299_/Y _75311_/Y _75312_/Y _75322_/A sky130_fd_sc_hd__o21a_4
X_41705_ _41704_/X _41705_/X sky130_fd_sc_hd__buf_2
X_48261_ _50308_/A _48201_/B _48195_/X _48261_/X sky130_fd_sc_hd__and3_4
X_72525_ _72525_/A _72525_/Y sky130_fd_sc_hd__inv_2
X_79081_ _82751_/Q _79082_/B sky130_fd_sc_hd__inv_2
X_45473_ _45470_/Y _45439_/X _45471_/X _45472_/Y _45473_/X sky130_fd_sc_hd__a211o_4
X_57459_ _57441_/X _56761_/X _57458_/X _57459_/X sky130_fd_sc_hd__o21a_4
X_76293_ _76293_/A _76283_/Y _76273_/A _76293_/Y sky130_fd_sc_hd__nor3_4
X_88279_ _87011_/CLK _41094_/X _69526_/B sky130_fd_sc_hd__dfxtp_4
X_42685_ _42665_/X _42666_/X _41076_/X _69480_/B _42673_/X _42685_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47212_ _47212_/A _47212_/Y sky130_fd_sc_hd__inv_2
X_78032_ _78021_/C _78027_/B _78030_/A _78033_/B sky130_fd_sc_hd__nand3_4
X_44424_ _41570_/X _44412_/X _87114_/Q _44413_/X _87114_/D sky130_fd_sc_hd__a2bb2o_4
X_75244_ _75223_/Y _75244_/Y sky130_fd_sc_hd__inv_2
X_41636_ _41635_/Y _41636_/X sky130_fd_sc_hd__buf_2
X_48192_ _48192_/A _48934_/A sky130_fd_sc_hd__buf_2
X_60470_ _60469_/X _60476_/A sky130_fd_sc_hd__buf_2
X_72456_ _57712_/X _85316_/Q _72324_/X _72456_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_10_446_0_CLK clkbuf_9_223_0_CLK/X _84192_/CLK sky130_fd_sc_hd__clkbuf_1
X_47143_ _47113_/A _47133_/B _47143_/C _52879_/D _47143_/X sky130_fd_sc_hd__and4_4
X_59129_ _59043_/A _59129_/X sky130_fd_sc_hd__buf_2
X_71407_ _71397_/X _83510_/Q _71406_/Y _71407_/X sky130_fd_sc_hd__a21o_4
X_44355_ _44355_/A _87152_/D sky130_fd_sc_hd__inv_2
X_75175_ _75175_/A _75175_/B _75175_/C _75178_/B sky130_fd_sc_hd__nand3_4
X_41567_ _41567_/A _41567_/Y sky130_fd_sc_hd__inv_2
X_72387_ _72339_/X _85323_/Q _72386_/X _72387_/X sky130_fd_sc_hd__o21a_4
X_43306_ _43296_/X _43305_/X _41209_/X _87489_/Q _43273_/X _43306_/Y
+ sky130_fd_sc_hd__o32ai_4
X_62140_ _84782_/Q _62140_/X sky130_fd_sc_hd__buf_2
X_74126_ _74119_/Y _74120_/Y _74125_/X _74126_/Y sky130_fd_sc_hd__o21ai_4
X_40518_ _40416_/A _40518_/B _40518_/X sky130_fd_sc_hd__or2_4
X_47074_ _47074_/A _52841_/D sky130_fd_sc_hd__buf_2
X_71338_ _71338_/A _70431_/C _71779_/B _71338_/Y sky130_fd_sc_hd__nand3_4
X_44286_ _44274_/X _44286_/Y sky130_fd_sc_hd__inv_2
X_79983_ _84928_/Q _65817_/C _79985_/A sky130_fd_sc_hd__xor2_4
X_41498_ _41497_/X _41498_/X sky130_fd_sc_hd__buf_2
X_46025_ _40541_/Y _46022_/X _67287_/B _46023_/X _86808_/D sky130_fd_sc_hd__a2bb2o_4
X_43237_ _43226_/X _43229_/X _41021_/X _87524_/Q _43232_/X _43237_/Y
+ sky130_fd_sc_hd__o32ai_4
X_62071_ _83243_/Q _63630_/A sky130_fd_sc_hd__inv_2
X_74057_ _86986_/Q _73916_/B _74056_/X _74057_/Y sky130_fd_sc_hd__o21ai_4
X_78934_ _78912_/B _82510_/D sky130_fd_sc_hd__inv_2
X_40449_ _40448_/Y _88390_/D sky130_fd_sc_hd__inv_2
X_71269_ _71168_/A _71276_/B _71276_/C _70656_/D _71269_/Y sky130_fd_sc_hd__nand4_4
X_61022_ _60998_/X _60992_/X _65296_/A _61022_/Y sky130_fd_sc_hd__a21oi_4
X_73008_ _88330_/Q _72803_/X _73007_/X _73008_/Y sky130_fd_sc_hd__o21ai_4
X_43168_ _43162_/X _43167_/X _40874_/X _73275_/A _43154_/X _43169_/A
+ sky130_fd_sc_hd__o32ai_4
X_78865_ _78852_/X _78865_/B _78865_/X sky130_fd_sc_hd__and2_4
X_65830_ _65757_/A _65830_/X sky130_fd_sc_hd__buf_2
X_42119_ _42118_/Y _42119_/Y sky130_fd_sc_hd__inv_2
X_77816_ _77795_/X _77808_/X _77816_/X sky130_fd_sc_hd__and2_4
X_47976_ _47970_/Y _47954_/X _47975_/X _47976_/Y sky130_fd_sc_hd__a21oi_4
X_43099_ _43085_/X _43086_/X _40739_/X _43098_/Y _43090_/X _87576_/D
+ sky130_fd_sc_hd__o32ai_4
X_78796_ _78782_/Y _78786_/X _78794_/A _78797_/B sky130_fd_sc_hd__nand3_4
X_49715_ _49632_/A _49715_/X sky130_fd_sc_hd__buf_2
X_46927_ _46923_/Y _46891_/X _46926_/X _46927_/Y sky130_fd_sc_hd__a21oi_4
X_65761_ _64902_/A _65761_/X sky130_fd_sc_hd__buf_2
X_77747_ _82260_/Q _77747_/B _77747_/X sky130_fd_sc_hd__or2_4
X_62973_ _62927_/A _62664_/B _62162_/X _62973_/Y sky130_fd_sc_hd__nand3_4
X_74959_ _74959_/A _74959_/B _74959_/Y sky130_fd_sc_hd__nand2_4
X_67500_ _67572_/A _86936_/Q _67500_/X sky130_fd_sc_hd__and2_4
X_64712_ _64702_/X _64712_/B _64711_/X _64737_/A sky130_fd_sc_hd__nand3_4
X_49646_ _49625_/A _49642_/B _49629_/X _52861_/D _49646_/X sky130_fd_sc_hd__and4_4
X_61924_ _61922_/X _61924_/B _61878_/C _61910_/D _61924_/Y sky130_fd_sc_hd__nand4_4
X_68480_ _68553_/A _68480_/B _68480_/X sky130_fd_sc_hd__and2_4
X_46858_ _46853_/Y _46844_/X _46857_/X _86696_/D sky130_fd_sc_hd__a21oi_4
X_65692_ _65825_/A _86512_/Q _65692_/X sky130_fd_sc_hd__and2_4
X_77678_ _77655_/A _77652_/Y _77653_/Y _77678_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_9_505_0_CLK clkbuf_9_505_0_CLK/A clkbuf_9_505_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_67431_ _67428_/X _67430_/X _67383_/X _67436_/A sky130_fd_sc_hd__a21o_4
X_79417_ _79439_/A _79417_/Y sky130_fd_sc_hd__inv_2
X_45809_ _57210_/B _45736_/B _45809_/Y sky130_fd_sc_hd__nor2_4
X_64643_ _64769_/A _64643_/B _64643_/X sky130_fd_sc_hd__and2_4
X_76629_ _81376_/Q _76628_/A _76629_/Y sky130_fd_sc_hd__xnor2_4
X_49577_ _49571_/X _49561_/B _49577_/C _52790_/D _49577_/X sky130_fd_sc_hd__and4_4
X_61855_ _62185_/B _61874_/B sky130_fd_sc_hd__buf_2
X_46789_ _86703_/Q _46767_/X _46788_/Y _46789_/Y sky130_fd_sc_hd__o21ai_4
X_48528_ _86514_/Q _48478_/X _48527_/Y _48528_/Y sky130_fd_sc_hd__o21ai_4
X_60806_ _60715_/X _60810_/B sky130_fd_sc_hd__buf_2
X_67362_ _87410_/Q _67358_/X _67360_/X _67361_/X _67362_/X sky130_fd_sc_hd__a211o_4
X_79348_ _79355_/B _79347_/Y _79348_/X sky130_fd_sc_hd__xor2_4
X_64574_ _64619_/A _64574_/X sky130_fd_sc_hd__buf_2
X_61786_ _59765_/A _61823_/B sky130_fd_sc_hd__buf_2
X_69101_ _87477_/Q _69098_/X _69010_/X _69100_/X _69101_/X sky130_fd_sc_hd__a211o_4
X_66313_ _66326_/A _86533_/Q _66313_/X sky130_fd_sc_hd__and2_4
X_63525_ _61489_/B _63487_/X _63523_/X _63524_/X _63525_/X sky130_fd_sc_hd__a211o_4
X_60737_ _60736_/X _60804_/C _60694_/C _60804_/B _59846_/X _60737_/Y
+ sky130_fd_sc_hd__a41oi_4
X_48459_ _48651_/A _48459_/X sky130_fd_sc_hd__buf_2
X_79279_ _84339_/Q _79279_/B _79285_/B sky130_fd_sc_hd__xor2_4
X_67293_ _67055_/X _67293_/X sky130_fd_sc_hd__buf_2
X_81310_ _81632_/CLK _76998_/X _81310_/Q sky130_fd_sc_hd__dfxtp_4
X_69032_ _87992_/Q _69007_/X _68916_/X _69031_/X _69032_/X sky130_fd_sc_hd__a211o_4
X_66244_ _66244_/A _66244_/B _66244_/Y sky130_fd_sc_hd__nand2_4
X_51470_ _86004_/Q _51458_/X _51469_/Y _51470_/Y sky130_fd_sc_hd__o21ai_4
X_63456_ _63456_/A _63456_/B _84322_/Q _63456_/Y sky130_fd_sc_hd__nor3_4
X_82290_ _82103_/CLK _82290_/D _82290_/Q sky130_fd_sc_hd__dfxtp_4
X_60668_ _60642_/C _60616_/Y _60644_/C _60667_/Y _60770_/A sky130_fd_sc_hd__and4_4
Xclkbuf_8_73_0_CLK clkbuf_8_73_0_CLK/A clkbuf_8_73_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_50421_ _50556_/A _52123_/B _50421_/Y sky130_fd_sc_hd__nand2_4
X_62407_ _62478_/A _62407_/X sky130_fd_sc_hd__buf_2
X_81241_ _85338_/CLK _81049_/Q _81241_/Q sky130_fd_sc_hd__dfxtp_4
X_66175_ _66046_/A _66177_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_5_0_CLK clkbuf_6_2_0_CLK/X clkbuf_7_5_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_63387_ _63400_/A _58225_/A _63400_/C _63387_/X sky130_fd_sc_hd__and3_4
X_60599_ _60599_/A _60403_/A _60403_/B _59508_/X _60599_/X sky130_fd_sc_hd__and4_4
X_65126_ _65126_/A _65125_/X _65126_/Y sky130_fd_sc_hd__nand2_4
X_53140_ _53136_/Y _53137_/X _53139_/X _85690_/D sky130_fd_sc_hd__a21oi_4
X_50352_ _50356_/A _57609_/B _50352_/Y sky130_fd_sc_hd__nand2_4
X_62338_ _61427_/B _62278_/X _60027_/A _62323_/X _62337_/X _62338_/X
+ sky130_fd_sc_hd__a41o_4
X_81172_ _82335_/CLK _74978_/B _41523_/A sky130_fd_sc_hd__dfxtp_4
Xpsn_inst_psn_buff_11 _44133_/Y _44134_/D sky130_fd_sc_hd__buf_8
Xpsn_inst_psn_buff_22 _53441_/A _43182_/B1 sky130_fd_sc_hd__buf_2
X_80123_ _84941_/Q _84189_/Q _80125_/A sky130_fd_sc_hd__xor2_4
X_53071_ _53068_/Y _53056_/X _53070_/X _85703_/D sky130_fd_sc_hd__a21oi_4
X_65057_ _64904_/A _85840_/Q _65057_/X sky130_fd_sc_hd__and2_4
X_69934_ _69931_/X _69933_/X _69624_/X _69937_/A sky130_fd_sc_hd__a21o_4
X_50283_ _50595_/A _50500_/A sky130_fd_sc_hd__buf_2
X_62269_ _62269_/A _62269_/X sky130_fd_sc_hd__buf_2
X_85980_ _85692_/CLK _85980_/D _85980_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_88_0_CLK clkbuf_8_89_0_CLK/A clkbuf_8_88_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_52022_ _52462_/A _52022_/X sky130_fd_sc_hd__buf_2
X_64008_ _63849_/A _64074_/B sky130_fd_sc_hd__buf_2
X_84931_ _86312_/CLK _84931_/D _84931_/Q sky130_fd_sc_hd__dfxtp_4
X_80054_ _80042_/A _80041_/Y _80053_/X _80054_/X sky130_fd_sc_hd__a21o_4
X_69865_ _69865_/A _69865_/B _69865_/X sky130_fd_sc_hd__and2_4
X_56830_ _56774_/A _85129_/Q _44135_/X _56830_/Y sky130_fd_sc_hd__nor3_4
X_68816_ _87489_/Q _68792_/X _68545_/X _68815_/X _68816_/X sky130_fd_sc_hd__a211o_4
X_87650_ _87394_/CLK _87650_/D _87650_/Q sky130_fd_sc_hd__dfxtp_4
X_84862_ _84344_/CLK _84862_/D _84862_/Q sky130_fd_sc_hd__dfxtp_4
X_69796_ _69796_/A _69796_/X sky130_fd_sc_hd__buf_2
X_86601_ _85961_/CLK _86601_/D _72405_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_11_0_CLK clkbuf_7_5_0_CLK/X clkbuf_9_23_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_83813_ _83813_/CLK _70278_/X _74775_/B sky130_fd_sc_hd__dfxtp_4
X_56761_ _56788_/A _56761_/X sky130_fd_sc_hd__buf_2
X_68747_ _41938_/A _68493_/X _68745_/X _68746_/Y _68747_/X sky130_fd_sc_hd__a211o_4
X_87581_ _87542_/CLK _43088_/Y _87581_/Q sky130_fd_sc_hd__dfxtp_4
X_53973_ _53929_/A _53978_/A sky130_fd_sc_hd__buf_2
X_65959_ _64694_/A _86589_/Q _65959_/X sky130_fd_sc_hd__and2_4
X_84793_ _86701_/CLK _58885_/Y _84793_/Q sky130_fd_sc_hd__dfxtp_4
X_58500_ _83425_/Q _58500_/Y sky130_fd_sc_hd__inv_2
X_55712_ _55711_/X _85283_/Q _55172_/A _55712_/Y sky130_fd_sc_hd__a21oi_4
X_86532_ _86490_/CLK _86532_/D _66326_/B sky130_fd_sc_hd__dfxtp_4
X_52924_ _52910_/A _52924_/B _52924_/Y sky130_fd_sc_hd__nand2_4
X_83744_ _86647_/CLK _83744_/D _47305_/A sky130_fd_sc_hd__dfxtp_4
X_59480_ _83432_/Q _59480_/Y sky130_fd_sc_hd__inv_2
X_56692_ _56663_/X _56693_/C sky130_fd_sc_hd__inv_2
X_80956_ _80991_/CLK _80956_/D _80956_/Q sky130_fd_sc_hd__dfxtp_4
X_68678_ _68674_/X _68677_/X _68477_/X _68678_/Y sky130_fd_sc_hd__a21oi_4
X_58431_ _58334_/X _58429_/Y _58430_/Y _84850_/D sky130_fd_sc_hd__a21oi_4
X_55643_ _55643_/A _55642_/X _55644_/A sky130_fd_sc_hd__and2_4
X_67629_ _67582_/A _67629_/B _67629_/X sky130_fd_sc_hd__and2_4
X_86463_ _83623_/CLK _86463_/D _64658_/B sky130_fd_sc_hd__dfxtp_4
X_52855_ _52850_/A _52855_/B _52855_/Y sky130_fd_sc_hd__nand2_4
X_83675_ _83676_/CLK _70877_/Y _83675_/Q sky130_fd_sc_hd__dfxtp_4
X_80887_ _80854_/CLK _80887_/D _80887_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_26_0_CLK clkbuf_8_27_0_CLK/A clkbuf_9_53_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_88202_ _87126_/CLK _41508_/X _88202_/Q sky130_fd_sc_hd__dfxtp_4
X_85414_ _86054_/CLK _85414_/D _85414_/Q sky130_fd_sc_hd__dfxtp_4
X_51806_ _51801_/Y _51793_/X _51805_/X _51806_/Y sky130_fd_sc_hd__a21oi_4
X_70640_ _53012_/B _70632_/X _70639_/Y _83737_/D sky130_fd_sc_hd__o21ai_4
X_58362_ _84868_/Q _63335_/A sky130_fd_sc_hd__inv_2
X_82626_ _81179_/CLK _82626_/D _82626_/Q sky130_fd_sc_hd__dfxtp_4
X_55574_ _85116_/Q _55571_/X _44049_/X _55573_/Y _55574_/X sky130_fd_sc_hd__a211o_4
X_86394_ _86393_/CLK _86394_/D _86394_/Q sky130_fd_sc_hd__dfxtp_4
X_52786_ _52782_/Y _52783_/X _52785_/X _52786_/Y sky130_fd_sc_hd__a21oi_4
X_57313_ _57049_/A _85036_/Q _57326_/C _57313_/Y sky130_fd_sc_hd__nor3_4
X_88133_ _88133_/CLK _41829_/Y _66920_/B sky130_fd_sc_hd__dfxtp_4
X_54525_ _85426_/Q _54512_/X _54524_/Y _54525_/Y sky130_fd_sc_hd__o21ai_4
X_85345_ _83711_/CLK _85345_/D _85345_/Q sky130_fd_sc_hd__dfxtp_4
X_51737_ _51737_/A _53259_/B _51737_/Y sky130_fd_sc_hd__nand2_4
X_70571_ _70570_/Y _71867_/A sky130_fd_sc_hd__buf_2
X_82557_ _82557_/CLK _82557_/D _78903_/B sky130_fd_sc_hd__dfxtp_4
X_58293_ _58282_/X _58290_/Y _58292_/Y _84886_/D sky130_fd_sc_hd__a21oi_4
X_72310_ _72209_/X _85970_/Q _72309_/X _72310_/Y sky130_fd_sc_hd__o21ai_4
X_57244_ _57235_/Y _57244_/X sky130_fd_sc_hd__buf_2
X_81508_ _83918_/CLK _76171_/B _81508_/Q sky130_fd_sc_hd__dfxtp_4
X_88064_ _87813_/CLK _88064_/D _73247_/A sky130_fd_sc_hd__dfxtp_4
X_42470_ _42466_/X _42467_/X _40610_/X _68490_/A _42453_/X _42470_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54456_ _54452_/Y _54448_/X _54455_/X _85439_/D sky130_fd_sc_hd__a21oi_4
X_73290_ _73290_/A _73290_/B _73290_/Y sky130_fd_sc_hd__nand2_4
X_85276_ _85277_/CLK _56207_/Y _56206_/C sky130_fd_sc_hd__dfxtp_4
X_51668_ _51694_/A _51684_/B sky130_fd_sc_hd__buf_2
X_82488_ _82518_/CLK _82488_/D _78174_/B sky130_fd_sc_hd__dfxtp_4
X_41421_ _41072_/X _41421_/X sky130_fd_sc_hd__buf_2
X_87015_ _88283_/CLK _44653_/X _87015_/Q sky130_fd_sc_hd__dfxtp_4
X_53407_ _85639_/Q _53404_/X _53406_/Y _53407_/Y sky130_fd_sc_hd__o21ai_4
X_72241_ _64591_/X _72241_/X sky130_fd_sc_hd__buf_2
X_84227_ _84231_/CLK _84227_/D _84227_/Q sky130_fd_sc_hd__dfxtp_4
X_50619_ _50577_/A _50619_/X sky130_fd_sc_hd__buf_2
X_57175_ _57175_/A _57175_/B _57175_/Y sky130_fd_sc_hd__nand2_4
X_81439_ _81532_/CLK _81471_/Q _76139_/B sky130_fd_sc_hd__dfxtp_4
X_54387_ _54383_/Y _54366_/X _54386_/X _85452_/D sky130_fd_sc_hd__a21oi_4
X_51599_ _51597_/Y _51585_/X _51598_/X _85981_/D sky130_fd_sc_hd__a21oi_4
X_44140_ _60665_/C _44003_/X _62975_/D _44140_/X sky130_fd_sc_hd__a21o_4
X_56126_ _56117_/C _56147_/A sky130_fd_sc_hd__inv_2
X_41352_ _41351_/Y _41352_/X sky130_fd_sc_hd__buf_2
X_53338_ _53311_/A _53339_/A sky130_fd_sc_hd__buf_2
X_72172_ _58864_/A _72172_/X sky130_fd_sc_hd__buf_2
X_84158_ _84166_/CLK _84158_/D _84158_/Q sky130_fd_sc_hd__dfxtp_4
X_71123_ _71112_/X _71055_/B _71119_/C _71123_/Y sky130_fd_sc_hd__nand3_4
X_83109_ _82998_/CLK _74296_/X _70277_/C sky130_fd_sc_hd__dfxtp_4
X_44071_ _44071_/A _44232_/B _87178_/Q _44071_/X sky130_fd_sc_hd__and3_4
X_56057_ _56029_/X _56055_/X _56056_/Y _56057_/Y sky130_fd_sc_hd__o21ai_4
X_41283_ _41181_/A _41283_/X sky130_fd_sc_hd__buf_2
X_53269_ _53269_/A _53276_/A sky130_fd_sc_hd__buf_2
X_76980_ _76980_/A _62527_/C _76980_/X sky130_fd_sc_hd__xor2_4
X_84089_ _81507_/CLK _84089_/D _80913_/D sky130_fd_sc_hd__dfxtp_4
X_43022_ _42439_/X _43017_/X _40560_/X _73554_/A _43021_/X _43023_/A
+ sky130_fd_sc_hd__o32ai_4
X_55008_ _85336_/Q _54994_/X _55007_/Y _55008_/Y sky130_fd_sc_hd__o21ai_4
X_71054_ _71054_/A _71055_/B sky130_fd_sc_hd__buf_2
X_75931_ _81700_/D _75930_/B _75932_/A sky130_fd_sc_hd__nand2_4
X_87917_ _86934_/CLK _87917_/D _87917_/Q sky130_fd_sc_hd__dfxtp_4
X_70005_ _69655_/A _70005_/X sky130_fd_sc_hd__buf_2
X_47830_ _83561_/Q _47830_/Y sky130_fd_sc_hd__inv_2
X_59816_ _59816_/A _61202_/A sky130_fd_sc_hd__buf_2
X_78650_ _78649_/B _78648_/Y _78645_/Y _78654_/C sky130_fd_sc_hd__o21ai_4
X_75862_ _75860_/B _75860_/A _75862_/Y sky130_fd_sc_hd__nand2_4
X_87848_ _87595_/CLK _42490_/Y _73820_/A sky130_fd_sc_hd__dfxtp_4
X_77601_ _77601_/A _82107_/D _77601_/Y sky130_fd_sc_hd__nand2_4
X_74813_ _46216_/A _74813_/Y sky130_fd_sc_hd__inv_2
X_47761_ _47620_/X _47799_/A sky130_fd_sc_hd__buf_2
X_59747_ _59737_/A _59711_/B _80539_/A _59747_/Y sky130_fd_sc_hd__nor3_4
X_78581_ _78600_/A _78581_/B _82772_/D sky130_fd_sc_hd__xor2_4
X_56959_ _56949_/X _56619_/X _45535_/A _56947_/X _85112_/D sky130_fd_sc_hd__a2bb2o_4
X_44973_ _44972_/X _44973_/X sky130_fd_sc_hd__buf_2
X_75793_ _75793_/A _75793_/B _80890_/D sky130_fd_sc_hd__xor2_4
X_87779_ _87533_/CLK _87779_/D _69354_/B sky130_fd_sc_hd__dfxtp_4
X_49500_ _49500_/A _49500_/B _49493_/X _52716_/D _49500_/X sky130_fd_sc_hd__and4_4
X_46712_ _46712_/A _51800_/B _46712_/Y sky130_fd_sc_hd__nand2_4
X_77532_ _77532_/A _82103_/D _77537_/A sky130_fd_sc_hd__nor2_4
X_43924_ _43854_/A _43924_/X sky130_fd_sc_hd__buf_2
X_74744_ _70732_/X _74744_/X sky130_fd_sc_hd__buf_2
X_47692_ _47692_/A _47692_/B _47692_/C _53191_/D _47692_/X sky130_fd_sc_hd__and4_4
X_71956_ _71942_/Y _83314_/Q _71955_/Y _71956_/X sky130_fd_sc_hd__a21o_4
X_59678_ _59621_/X _59619_/X _59753_/B _72569_/C _59600_/X _59680_/A
+ sky130_fd_sc_hd__a32oi_4
X_49431_ _49418_/A _46740_/X _49431_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_370_0_CLK clkbuf_9_185_0_CLK/X _86361_/CLK sky130_fd_sc_hd__clkbuf_1
X_46643_ _46651_/A _51765_/B _46643_/Y sky130_fd_sc_hd__nand2_4
X_58629_ _58112_/X _86108_/Q _58628_/X _58629_/Y sky130_fd_sc_hd__o21ai_4
X_70907_ _70358_/X _70907_/B _70495_/A _70908_/A sky130_fd_sc_hd__nand3_4
X_77463_ _77461_/X _77431_/Y _77462_/Y _77463_/X sky130_fd_sc_hd__a21o_4
X_43855_ _43846_/X _43854_/X _41214_/X _87232_/Q _43847_/X _43855_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74675_ _74675_/A _74675_/X sky130_fd_sc_hd__buf_2
X_71887_ _71887_/A _71783_/A _71783_/C _71883_/D _71887_/Y sky130_fd_sc_hd__nor4_4
X_79202_ _84789_/Q _66509_/C _79202_/Y sky130_fd_sc_hd__nand2_4
X_76414_ _76395_/Y _76392_/Y _76394_/A _76415_/A sky130_fd_sc_hd__o21a_4
X_42806_ _42795_/X _42796_/X _41403_/X _87709_/Q _42805_/X _42806_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49362_ _49382_/A _51744_/B _49362_/Y sky130_fd_sc_hd__nand2_4
X_61640_ _61640_/A _61611_/B _61611_/C _61639_/X _61640_/Y sky130_fd_sc_hd__nand4_4
X_73626_ _41889_/Y _73529_/X _73344_/X _73625_/Y _73626_/X sky130_fd_sc_hd__a211o_4
X_70838_ _70832_/A _70849_/C sky130_fd_sc_hd__buf_2
X_46574_ _46547_/A _50870_/B _46574_/Y sky130_fd_sc_hd__nand2_4
X_77394_ _77394_/A _77394_/B _77417_/B sky130_fd_sc_hd__xor2_4
X_43786_ _43774_/X _43781_/X _41021_/X _87268_/Q _43776_/X _43787_/A
+ sky130_fd_sc_hd__o32ai_4
X_40998_ _40686_/A _40999_/A sky130_fd_sc_hd__buf_2
X_48313_ _48275_/X _50356_/B _48313_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_491_0_CLK clkbuf_9_491_0_CLK/A clkbuf_9_491_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_79133_ _79133_/A _79133_/B _79133_/X sky130_fd_sc_hd__xor2_4
X_45525_ _56614_/B _45343_/X _45378_/X _45525_/X sky130_fd_sc_hd__o21a_4
X_76345_ _76345_/A _81564_/Q _76348_/B sky130_fd_sc_hd__nor2_4
X_42737_ _42721_/X _42723_/X _41220_/X _68868_/B _42732_/X _42737_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49293_ _50812_/A _49283_/B _49234_/X _49293_/X sky130_fd_sc_hd__and3_4
X_61571_ _61342_/X _61572_/D sky130_fd_sc_hd__buf_2
X_73557_ _88371_/Q _72769_/B _72866_/X _73557_/X sky130_fd_sc_hd__o21a_4
X_70769_ _70863_/A _70779_/B _70766_/C _70769_/D _70769_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_10_385_0_CLK clkbuf_9_192_0_CLK/X _83216_/CLK sky130_fd_sc_hd__clkbuf_1
X_63310_ _72381_/A _63310_/X sky130_fd_sc_hd__buf_2
X_48244_ _48244_/A _50293_/B _48244_/Y sky130_fd_sc_hd__nand2_4
X_60522_ _60522_/A _60523_/A sky130_fd_sc_hd__buf_2
X_72508_ _72508_/A _72516_/A sky130_fd_sc_hd__buf_2
X_79064_ _79064_/A _79064_/B _79065_/A sky130_fd_sc_hd__xor2_4
X_45456_ _45612_/A _45456_/X sky130_fd_sc_hd__buf_2
X_64290_ _64282_/Y _64289_/X _64269_/X _64290_/X sky130_fd_sc_hd__o21a_4
X_76276_ _81643_/Q _76276_/B _76276_/X sky130_fd_sc_hd__or2_4
X_42668_ _42667_/Y _42668_/Y sky130_fd_sc_hd__inv_2
X_73488_ _43199_/Y _72895_/X _73486_/X _73487_/Y _73488_/X sky130_fd_sc_hd__a211o_4
X_78015_ _82079_/Q _78012_/Y _78014_/X _78015_/Y sky130_fd_sc_hd__o21ai_4
X_44407_ _44404_/X _44405_/X _41515_/X _87124_/Q _44406_/X _44407_/Y
+ sky130_fd_sc_hd__o32ai_4
X_63241_ _63216_/X _63241_/B _63241_/C _63240_/X _63241_/X sky130_fd_sc_hd__and4_4
X_75227_ _75226_/Y _75227_/Y sky130_fd_sc_hd__inv_2
X_41619_ _81155_/Q _41563_/B _41619_/X sky130_fd_sc_hd__or2_4
X_60453_ _60452_/X _60454_/A sky130_fd_sc_hd__buf_2
X_72439_ _64758_/X _85318_/Q _72386_/X _72439_/X sky130_fd_sc_hd__o21a_4
X_48175_ _48226_/A _48175_/X sky130_fd_sc_hd__buf_2
X_45387_ _45387_/A _45596_/A sky130_fd_sc_hd__buf_2
X_42599_ _42599_/A _42599_/Y sky130_fd_sc_hd__inv_2
X_47126_ _59270_/A _47096_/X _47125_/Y _47126_/Y sky130_fd_sc_hd__o21ai_4
X_44338_ _44330_/X _44331_/X _41676_/X _87159_/Q _44332_/X _44339_/A
+ sky130_fd_sc_hd__o32ai_4
X_63172_ _63231_/A _63172_/X sky130_fd_sc_hd__buf_2
X_75158_ _81063_/Q _75158_/Y sky130_fd_sc_hd__inv_2
X_60384_ _60392_/A _60392_/C _60404_/C sky130_fd_sc_hd__and2_4
X_62123_ _62118_/Y _62101_/X _62122_/Y _84432_/D sky130_fd_sc_hd__a21oi_4
X_74109_ _74152_/A _66238_/B _74109_/X sky130_fd_sc_hd__and2_4
X_47057_ _82387_/Q _54522_/D sky130_fd_sc_hd__inv_2
X_44269_ _44187_/A _72908_/A sky130_fd_sc_hd__buf_2
X_67980_ _86948_/Q _67906_/X _67908_/X _67979_/X _67981_/B sky130_fd_sc_hd__a211o_4
X_79966_ _79964_/Y _79965_/Y _79966_/X sky130_fd_sc_hd__xor2_4
X_75089_ _75087_/Y _81058_/Q _75088_/Y _75091_/B sky130_fd_sc_hd__a21bo_4
X_46008_ _45975_/X _46008_/X sky130_fd_sc_hd__buf_2
X_66931_ _66928_/X _66930_/X _66905_/X _66931_/X sky130_fd_sc_hd__a21o_4
X_62054_ _59588_/Y _62055_/A sky130_fd_sc_hd__buf_2
X_78917_ _82637_/Q _82509_/D _78916_/X _78918_/B sky130_fd_sc_hd__o21ai_4
X_79897_ _79896_/Y _60152_/A _79899_/A sky130_fd_sc_hd__nand2_4
X_61005_ _60854_/Y _60915_/A _60928_/X _63734_/A sky130_fd_sc_hd__a21boi_4
Xclkbuf_10_323_0_CLK clkbuf_9_161_0_CLK/X _85725_/CLK sky130_fd_sc_hd__clkbuf_1
X_69650_ _69647_/X _69649_/X _69385_/X _69650_/X sky130_fd_sc_hd__a21o_4
X_66862_ _87879_/Q _66816_/X _66794_/X _66861_/X _66862_/X sky130_fd_sc_hd__a211o_4
X_78848_ _78839_/X _78840_/A _78856_/A sky130_fd_sc_hd__nand2_4
Xclkbuf_10_953_0_CLK clkbuf_9_476_0_CLK/X _88081_/CLK sky130_fd_sc_hd__clkbuf_1
X_68601_ _68450_/A _68601_/X sky130_fd_sc_hd__buf_2
X_65813_ _65811_/X _83056_/Q _65768_/X _65812_/X _65813_/X sky130_fd_sc_hd__a211o_4
X_69581_ _43115_/A _69506_/X _66349_/X _69580_/X _69581_/X sky130_fd_sc_hd__a211o_4
X_47959_ _47959_/A _73864_/A sky130_fd_sc_hd__inv_2
X_78779_ _78778_/X _78779_/Y sky130_fd_sc_hd__inv_2
X_66793_ _66910_/A _66793_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_444_0_CLK clkbuf_9_444_0_CLK/A clkbuf_9_444_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_80810_ _80821_/CLK _83954_/Q _75786_/B sky130_fd_sc_hd__dfxtp_4
X_68532_ _68529_/X _68531_/X _68429_/X _68532_/X sky130_fd_sc_hd__a21o_4
X_65744_ _84181_/Q _65745_/C sky130_fd_sc_hd__inv_2
X_50970_ _50968_/Y _50957_/X _50969_/X _50970_/Y sky130_fd_sc_hd__a21oi_4
X_62956_ _58198_/A _62808_/X _62827_/X _62818_/X _62955_/X _62956_/Y
+ sky130_fd_sc_hd__a41oi_4
X_81790_ _83133_/CLK _81790_/D _48914_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_338_0_CLK clkbuf_9_169_0_CLK/X _82381_/CLK sky130_fd_sc_hd__clkbuf_1
X_49629_ _49548_/A _49629_/X sky130_fd_sc_hd__buf_2
X_61907_ _61461_/X _61874_/B _61907_/C _61874_/D _61907_/Y sky130_fd_sc_hd__nand4_4
X_80741_ _81994_/CLK _80741_/D _81149_/D sky130_fd_sc_hd__dfxtp_4
X_68463_ _69645_/A _68463_/X sky130_fd_sc_hd__buf_2
X_65675_ _65596_/X _83065_/Q _65540_/X _65674_/X _65675_/X sky130_fd_sc_hd__a211o_4
X_62887_ _60362_/A _62965_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_968_0_CLK clkbuf_9_484_0_CLK/X _86541_/CLK sky130_fd_sc_hd__clkbuf_1
X_67414_ _67055_/X _67414_/X sky130_fd_sc_hd__buf_2
X_52640_ _52638_/Y _52619_/X _52639_/X _52640_/Y sky130_fd_sc_hd__a21oi_4
X_64626_ _64803_/A _64680_/A sky130_fd_sc_hd__buf_2
X_83460_ _83495_/CLK _71549_/X _83460_/Q sky130_fd_sc_hd__dfxtp_4
X_61838_ _61755_/X _61838_/X sky130_fd_sc_hd__buf_2
X_80672_ _80672_/CLK _80672_/D _80672_/Q sky130_fd_sc_hd__dfxtp_4
X_68394_ _68394_/A _68394_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_459_0_CLK clkbuf_9_459_0_CLK/A clkbuf_9_459_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_82411_ _82443_/CLK _82411_/D _78432_/A sky130_fd_sc_hd__dfxtp_4
X_67345_ _67320_/A _86943_/Q _67345_/X sky130_fd_sc_hd__and2_4
X_52571_ _52518_/A _52571_/B _52571_/Y sky130_fd_sc_hd__nand2_4
X_64557_ _58993_/Y _61085_/X _64556_/Y _64557_/Y sky130_fd_sc_hd__o21ai_4
X_83391_ _85407_/CLK _83391_/D _47242_/A sky130_fd_sc_hd__dfxtp_4
X_61769_ _61767_/Y _61699_/X _61768_/Y _61769_/Y sky130_fd_sc_hd__a21oi_4
XPHY_508 sky130_fd_sc_hd__decap_3
X_54310_ _85465_/Q _54294_/X _54309_/Y _54310_/Y sky130_fd_sc_hd__o21ai_4
XPHY_519 sky130_fd_sc_hd__decap_3
X_85130_ _85067_/CLK _56827_/Y _85130_/Q sky130_fd_sc_hd__dfxtp_4
X_51522_ _51521_/X _51527_/B _51522_/C _53048_/D _51522_/X sky130_fd_sc_hd__and4_4
X_63508_ _63506_/Y _63455_/X _63507_/Y _84318_/D sky130_fd_sc_hd__a21oi_4
X_82342_ _82369_/CLK _77081_/X _82342_/Q sky130_fd_sc_hd__dfxtp_4
X_55290_ _55290_/A _55290_/Y sky130_fd_sc_hd__inv_2
X_67276_ _87414_/Q _67274_/X _67226_/X _67275_/X _67276_/X sky130_fd_sc_hd__a211o_4
X_64488_ _58970_/A _61085_/X _64487_/Y _64488_/Y sky130_fd_sc_hd__o21ai_4
X_69015_ _69059_/A _88249_/Q _69015_/X sky130_fd_sc_hd__and2_4
X_54241_ _54255_/A _54237_/B _54237_/C _53074_/D _54241_/X sky130_fd_sc_hd__and4_4
X_66227_ _66225_/X _84971_/Q _66186_/X _66226_/X _66227_/X sky130_fd_sc_hd__a211o_4
X_85061_ _85128_/CLK _85061_/D _57217_/B sky130_fd_sc_hd__dfxtp_4
X_51453_ _51446_/Y _51448_/X _51452_/X _86008_/D sky130_fd_sc_hd__a21oi_4
X_63439_ _63427_/A _61831_/X _63439_/X sky130_fd_sc_hd__and2_4
X_82273_ _83508_/CLK _80634_/Y _82273_/Q sky130_fd_sc_hd__dfxtp_4
X_84012_ _84074_/CLK _68206_/X _82052_/D sky130_fd_sc_hd__dfxtp_4
X_50404_ _50213_/X _50432_/A sky130_fd_sc_hd__buf_2
X_81224_ _81224_/CLK _81032_/Q _81224_/Q sky130_fd_sc_hd__dfxtp_4
X_54172_ _54254_/A _54191_/C sky130_fd_sc_hd__buf_2
X_66158_ _66391_/A _66385_/B sky130_fd_sc_hd__buf_2
X_51384_ _51367_/X _51384_/B _51384_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_906_0_CLK clkbuf_9_453_0_CLK/X _87850_/CLK sky130_fd_sc_hd__clkbuf_1
X_53123_ _85693_/Q _53120_/X _53122_/Y _53123_/Y sky130_fd_sc_hd__o21ai_4
X_65109_ _65005_/X _65109_/B _65109_/X sky130_fd_sc_hd__and2_4
X_50335_ _50398_/A _52036_/B _50335_/Y sky130_fd_sc_hd__nand2_4
X_81155_ _81179_/CLK _74853_/B _81155_/Q sky130_fd_sc_hd__dfxtp_4
X_66089_ _66426_/A _65741_/B _66426_/C _66089_/Y sky130_fd_sc_hd__nand3_4
X_58980_ _58559_/X _83438_/Q _58979_/Y _84782_/D sky130_fd_sc_hd__o21a_4
Xclkbuf_5_23_0_CLK clkbuf_5_23_0_CLK/A clkbuf_6_47_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_80106_ _80098_/B _80098_/A _80105_/X _80106_/Y sky130_fd_sc_hd__a21boi_4
X_53054_ _53040_/X _53054_/B _53054_/Y sky130_fd_sc_hd__nand2_4
X_57931_ _86643_/Q _57791_/X _57931_/Y sky130_fd_sc_hd__nor2_4
X_69917_ _69917_/A _69918_/B sky130_fd_sc_hd__inv_2
X_50266_ _50230_/A _53488_/B _50266_/Y sky130_fd_sc_hd__nand2_4
X_85963_ _85962_/CLK _85963_/D _85963_/Q sky130_fd_sc_hd__dfxtp_4
X_81086_ _81087_/CLK _81118_/Q _81086_/Q sky130_fd_sc_hd__dfxtp_4
X_52005_ _52027_/A _50302_/B _52005_/Y sky130_fd_sc_hd__nand2_4
X_87702_ _87221_/CLK _87702_/D _87702_/Q sky130_fd_sc_hd__dfxtp_4
X_80037_ _84932_/Q _84180_/Q _80037_/Y sky130_fd_sc_hd__nand2_4
X_84914_ _84914_/CLK _84914_/D _58177_/A sky130_fd_sc_hd__dfxtp_4
X_57862_ _57852_/X _85720_/Q _57814_/X _57862_/X sky130_fd_sc_hd__o21a_4
X_69848_ _69633_/A _73299_/A _69848_/X sky130_fd_sc_hd__and2_4
X_50197_ _51242_/A _50710_/B _50197_/X sky130_fd_sc_hd__and2_4
X_85894_ _86213_/CLK _85894_/D _66296_/B sky130_fd_sc_hd__dfxtp_4
X_59601_ _59751_/A _59752_/A _59639_/A sky130_fd_sc_hd__and2_4
X_56813_ _57029_/A _56812_/X _56814_/A sky130_fd_sc_hd__nand2_4
X_87633_ _88201_/CLK _87633_/D _66616_/B sky130_fd_sc_hd__dfxtp_4
X_84845_ _84877_/CLK _84845_/D _84845_/Q sky130_fd_sc_hd__dfxtp_4
X_57793_ _58007_/A _57793_/X sky130_fd_sc_hd__buf_2
X_69779_ _69779_/A _69779_/X sky130_fd_sc_hd__buf_2
X_71810_ _70502_/Y _71813_/A sky130_fd_sc_hd__buf_2
X_59532_ _59532_/A _59716_/B sky130_fd_sc_hd__buf_2
X_56744_ _57179_/A _85135_/Q _56744_/Y sky130_fd_sc_hd__nand2_4
X_41970_ _41965_/X _41956_/X _40739_/X _41969_/Y _41967_/X _41970_/Y
+ sky130_fd_sc_hd__o32ai_4
X_87564_ _87821_/CLK _87564_/D _43133_/A sky130_fd_sc_hd__dfxtp_4
X_53956_ _53956_/A _53956_/X sky130_fd_sc_hd__buf_2
X_72790_ _72774_/X _72791_/C _72789_/X _72790_/X sky130_fd_sc_hd__a21o_4
X_84776_ _86688_/CLK _84776_/D _84776_/Q sky130_fd_sc_hd__dfxtp_4
X_81988_ _82104_/CLK _81988_/D _77009_/A sky130_fd_sc_hd__dfxtp_4
X_86515_ _85581_/CLK _86515_/D _86515_/Q sky130_fd_sc_hd__dfxtp_4
X_40921_ _40921_/A _40921_/X sky130_fd_sc_hd__buf_2
X_52907_ _52852_/A _52916_/B sky130_fd_sc_hd__buf_2
X_71741_ _71168_/A _70656_/B _71279_/C _71744_/D _71741_/Y sky130_fd_sc_hd__nand4_4
X_59463_ _59463_/A _59463_/Y sky130_fd_sc_hd__inv_2
X_83727_ _85381_/CLK _83727_/D _47468_/A sky130_fd_sc_hd__dfxtp_4
X_56675_ _83332_/Q _56675_/X sky130_fd_sc_hd__buf_2
X_80939_ _80804_/CLK _80983_/Q _80939_/Q sky130_fd_sc_hd__dfxtp_4
X_87495_ _87758_/CLK _87495_/D _87495_/Q sky130_fd_sc_hd__dfxtp_4
X_53887_ _85548_/Q _53869_/X _53886_/Y _53887_/Y sky130_fd_sc_hd__o21ai_4
X_58414_ _84854_/Q _58415_/A sky130_fd_sc_hd__inv_2
X_43640_ _40678_/X _43624_/X _87331_/Q _43625_/X _43640_/X sky130_fd_sc_hd__a2bb2o_4
X_74460_ _74457_/Y _74430_/X _74459_/X _74460_/Y sky130_fd_sc_hd__a21oi_4
X_55626_ _45409_/A _55617_/X _44052_/A _55625_/Y _55626_/X sky130_fd_sc_hd__a211o_4
X_86446_ _85557_/CLK _86446_/D _65100_/B sky130_fd_sc_hd__dfxtp_4
X_40852_ _40829_/A _40852_/B _40852_/X sky130_fd_sc_hd__or2_4
X_52838_ _85745_/Q _52821_/X _52837_/Y _52838_/Y sky130_fd_sc_hd__o21ai_4
X_83658_ _83660_/CLK _70931_/Y _46911_/A sky130_fd_sc_hd__dfxtp_4
X_71672_ _71680_/A _71671_/X _71672_/C _71672_/Y sky130_fd_sc_hd__nand3_4
X_59394_ _58982_/A _59394_/X sky130_fd_sc_hd__buf_2
X_73411_ _73412_/B _73412_/C _73410_/X _73411_/X sky130_fd_sc_hd__a21o_4
X_70623_ _70727_/A _70620_/B _70620_/C _70620_/D _70623_/Y sky130_fd_sc_hd__nand4_4
X_58345_ _58341_/X _58342_/Y _58344_/Y _84873_/D sky130_fd_sc_hd__a21oi_4
X_82609_ _82702_/CLK _78947_/B _82609_/Q sky130_fd_sc_hd__dfxtp_4
X_43571_ _43570_/Y _87355_/D sky130_fd_sc_hd__inv_2
X_55557_ _55554_/X _55556_/X _44113_/X _56595_/A sky130_fd_sc_hd__a21o_4
X_74391_ _74391_/A _52123_/B _74391_/Y sky130_fd_sc_hd__nand2_4
X_86377_ _83666_/CLK _86377_/D _86377_/Q sky130_fd_sc_hd__dfxtp_4
X_40783_ _40783_/A _40783_/X sky130_fd_sc_hd__buf_2
X_52769_ _85758_/Q _52765_/X _52768_/Y _52769_/Y sky130_fd_sc_hd__o21ai_4
X_83589_ _83589_/CLK _71153_/Y _83589_/Q sky130_fd_sc_hd__dfxtp_4
X_45310_ _45302_/X _45307_/Y _45309_/Y _45310_/Y sky130_fd_sc_hd__a21oi_4
X_76130_ _76130_/A _76130_/B _76130_/X sky130_fd_sc_hd__xor2_4
X_88116_ _88116_/CLK _88116_/D _88116_/Q sky130_fd_sc_hd__dfxtp_4
X_42522_ _42574_/A _42522_/X sky130_fd_sc_hd__buf_2
X_54508_ _54401_/A _54509_/C sky130_fd_sc_hd__buf_2
X_73342_ _69873_/Y _73224_/X _56935_/X _73341_/Y _73342_/X sky130_fd_sc_hd__a211o_4
X_85328_ _83550_/CLK _85328_/D _85328_/Q sky130_fd_sc_hd__dfxtp_4
X_46290_ _46290_/A _72052_/A sky130_fd_sc_hd__buf_2
X_70554_ _70554_/A _70568_/C sky130_fd_sc_hd__buf_2
X_58276_ _84890_/Q _58277_/A sky130_fd_sc_hd__inv_2
X_55488_ _85138_/Q _55489_/B sky130_fd_sc_hd__inv_2
X_45241_ _85195_/Q _45176_/X _45240_/X _45241_/Y sky130_fd_sc_hd__o21ai_4
X_57227_ _57121_/X _56917_/A _57226_/X _57227_/Y sky130_fd_sc_hd__o21ai_4
X_76061_ _81525_/Q _76061_/B _76061_/X sky130_fd_sc_hd__xor2_4
X_88047_ _87544_/CLK _42071_/Y _88047_/Q sky130_fd_sc_hd__dfxtp_4
X_42453_ _42612_/A _42453_/X sky130_fd_sc_hd__buf_2
X_54439_ _54385_/A _54440_/B sky130_fd_sc_hd__buf_2
X_85259_ _85192_/CLK _85259_/D _56250_/C sky130_fd_sc_hd__dfxtp_4
X_73273_ _73273_/A _73196_/B _73273_/Y sky130_fd_sc_hd__nor2_4
X_70485_ _70400_/A _71777_/B sky130_fd_sc_hd__buf_2
X_75012_ _80768_/Q _75020_/C _75011_/Y _75013_/B sky130_fd_sc_hd__a21oi_4
X_41404_ _41399_/X _41400_/X _41403_/X _67860_/B _41388_/X _41405_/A
+ sky130_fd_sc_hd__o32ai_4
X_72224_ _72224_/A _72224_/Y sky130_fd_sc_hd__inv_2
X_45172_ _45127_/X _61538_/B _45144_/X _45172_/Y sky130_fd_sc_hd__o21ai_4
X_57158_ _57158_/A _57158_/B _57158_/C _57158_/Y sky130_fd_sc_hd__nor3_4
X_42384_ _40331_/X _42374_/X _87890_/Q _42375_/X _42384_/X sky130_fd_sc_hd__a2bb2o_4
X_44123_ _44187_/A _44124_/A sky130_fd_sc_hd__inv_2
X_56109_ _56109_/A _56109_/X sky130_fd_sc_hd__buf_2
X_79820_ _79804_/X _79820_/B _79820_/Y sky130_fd_sc_hd__nor2_4
X_41335_ _41334_/Y _88234_/D sky130_fd_sc_hd__inv_2
X_72155_ _72155_/A _72155_/X sky130_fd_sc_hd__buf_2
X_49980_ _49976_/Y _49977_/X _49979_/X _86288_/D sky130_fd_sc_hd__a21oi_4
X_57089_ _73183_/A _73186_/A sky130_fd_sc_hd__buf_2
X_71106_ _71101_/X _71082_/B _71099_/C _71106_/Y sky130_fd_sc_hd__nand3_4
X_48931_ _48931_/A _52287_/B sky130_fd_sc_hd__buf_2
X_44054_ _87180_/Q _44054_/Y sky130_fd_sc_hd__inv_2
X_79751_ _79745_/Y _79750_/Y _79751_/X sky130_fd_sc_hd__xor2_4
X_41266_ _41266_/A _41280_/B _41266_/X sky130_fd_sc_hd__or2_4
X_72086_ _72053_/A _49144_/A _72086_/Y sky130_fd_sc_hd__nand2_4
X_76963_ _76874_/Y _76963_/Y sky130_fd_sc_hd__inv_2
X_43005_ _43774_/A _43005_/X sky130_fd_sc_hd__buf_2
X_78702_ _78684_/X _78702_/Y sky130_fd_sc_hd__inv_2
X_71037_ _53167_/B _71013_/A _71036_/Y _83628_/D sky130_fd_sc_hd__o21ai_4
X_75914_ _61185_/C _62766_/C _75914_/X sky130_fd_sc_hd__xor2_4
X_48862_ _48837_/A _50056_/A sky130_fd_sc_hd__buf_2
X_79682_ _79678_/X _79682_/B _79704_/B sky130_fd_sc_hd__xor2_4
X_41197_ _81713_/Q _41197_/B _41197_/X sky130_fd_sc_hd__or2_4
X_76894_ _76894_/A _76894_/Y sky130_fd_sc_hd__inv_2
X_47813_ _81219_/Q _47814_/A sky130_fd_sc_hd__inv_2
X_78633_ _78632_/B _78632_/C _78628_/Y _78637_/C sky130_fd_sc_hd__o21ai_4
X_75845_ _75841_/Y _75844_/Y _75846_/A sky130_fd_sc_hd__xor2_4
X_48793_ _48793_/A _48540_/B _48793_/Y sky130_fd_sc_hd__nand2_4
X_62810_ _57672_/X _62808_/X _62768_/X _62759_/X _62809_/X _62810_/Y
+ sky130_fd_sc_hd__a41oi_4
X_47744_ _86602_/Q _47714_/X _47743_/Y _47744_/Y sky130_fd_sc_hd__o21ai_4
X_78564_ _82515_/Q _82771_/D _78564_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_7_121_0_CLK clkbuf_6_60_0_CLK/X clkbuf_8_243_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_44956_ _85245_/Q _44874_/X _44926_/X _44956_/X sky130_fd_sc_hd__o21a_4
X_63790_ _61003_/A _63790_/X sky130_fd_sc_hd__buf_2
X_75776_ _75771_/Y _75775_/Y _80888_/D sky130_fd_sc_hd__xor2_4
X_72988_ _72720_/A _72988_/X sky130_fd_sc_hd__buf_2
X_77515_ _81941_/Q _82197_/D _81909_/D sky130_fd_sc_hd__xor2_4
X_43907_ _43842_/A _43907_/X sky130_fd_sc_hd__buf_2
X_62741_ _62679_/X _62743_/B sky130_fd_sc_hd__buf_2
X_74727_ _74727_/A _74796_/C _71738_/X _71016_/A _74730_/C sky130_fd_sc_hd__nand4_4
X_47675_ _47675_/A _53181_/D sky130_fd_sc_hd__buf_2
X_71939_ _71938_/Y _71939_/X sky130_fd_sc_hd__buf_2
X_78495_ _78486_/Y _78515_/A _78499_/A sky130_fd_sc_hd__xor2_4
X_44887_ _80672_/Q _44887_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_91_0_CLK clkbuf_9_45_0_CLK/X _84421_/CLK sky130_fd_sc_hd__clkbuf_1
X_49414_ _49411_/Y _49405_/X _49413_/X _49414_/Y sky130_fd_sc_hd__a21oi_4
X_46626_ _46651_/A _46625_/X _46626_/Y sky130_fd_sc_hd__nand2_4
X_65460_ _65428_/X _83079_/Q _65407_/X _65459_/X _65461_/B sky130_fd_sc_hd__a211o_4
X_77446_ _77446_/A _77446_/Y sky130_fd_sc_hd__inv_2
X_43838_ _41169_/X _43832_/X _87240_/Q _43833_/X _43838_/X sky130_fd_sc_hd__a2bb2o_4
X_62672_ _62672_/A _62673_/B sky130_fd_sc_hd__buf_2
X_74658_ _56666_/Y _74656_/X _74657_/Y _74659_/A sky130_fd_sc_hd__a21bo_4
X_64411_ _64377_/X _64411_/B _64391_/X _64411_/X sky130_fd_sc_hd__and3_4
X_49345_ _65343_/B _49334_/X _49344_/Y _49345_/Y sky130_fd_sc_hd__o21ai_4
X_61623_ _61617_/Y _61619_/Y _61583_/Y _61620_/Y _61622_/Y _61623_/X
+ sky130_fd_sc_hd__a41o_4
X_73609_ _74012_/A _73609_/X sky130_fd_sc_hd__buf_2
X_46557_ _86726_/Q _46543_/X _46556_/Y _46557_/Y sky130_fd_sc_hd__o21ai_4
X_65391_ _64991_/A _65391_/X sky130_fd_sc_hd__buf_2
X_77377_ _77367_/X _82220_/Q _77376_/Y _77386_/A sky130_fd_sc_hd__a21boi_4
X_43769_ _40982_/X _43752_/X _69262_/B _43753_/X _43769_/X sky130_fd_sc_hd__a2bb2o_4
X_74589_ _74575_/X _74583_/X _56099_/A _74584_/X _74589_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_opt_8_CLK clkbuf_opt_9_CLK/A _84888_/CLK sky130_fd_sc_hd__clkbuf_16
X_67130_ _67130_/A _67129_/X _67130_/Y sky130_fd_sc_hd__nand2_4
X_79116_ _78960_/Y _82515_/D sky130_fd_sc_hd__inv_2
X_45508_ _85146_/Q _45507_/X _45429_/X _45508_/X sky130_fd_sc_hd__o21a_4
X_64342_ _64304_/A _64303_/X _57664_/A _64318_/D _64342_/X sky130_fd_sc_hd__and4_4
X_76328_ _76328_/A _81518_/D _76328_/Y sky130_fd_sc_hd__nand2_4
X_49276_ _86419_/Q _49255_/X _49275_/Y _49276_/Y sky130_fd_sc_hd__o21ai_4
X_61554_ _61548_/Y _61550_/Y _61525_/X _61551_/Y _61553_/Y _61554_/X
+ sky130_fd_sc_hd__a41o_4
X_46488_ _46479_/Y _46445_/X _46487_/X _46488_/Y sky130_fd_sc_hd__a21oi_4
X_48227_ _49173_/A _48229_/A sky130_fd_sc_hd__buf_2
X_60505_ _60566_/A _60595_/C _59512_/A _60586_/D sky130_fd_sc_hd__a21oi_4
X_67061_ _67058_/X _67060_/X _66964_/X _67061_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_8_252_0_CLK clkbuf_8_253_0_CLK/A clkbuf_9_505_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_79047_ _82748_/Q _79047_/B _82716_/D sky130_fd_sc_hd__xor2_4
X_45439_ _45596_/A _45439_/X sky130_fd_sc_hd__buf_2
X_64273_ _64273_/A _64273_/B _84900_/Q _64304_/D _64273_/X sky130_fd_sc_hd__and4_4
X_76259_ _81353_/Q _76258_/Y _81321_/D sky130_fd_sc_hd__xor2_4
X_61485_ _61485_/A _61485_/Y sky130_fd_sc_hd__inv_2
X_66012_ _66011_/X _86554_/Q _66012_/X sky130_fd_sc_hd__and2_4
X_63224_ _60466_/X _63312_/C sky130_fd_sc_hd__buf_2
X_48158_ _46301_/X _82338_/Q _48157_/X _52093_/A sky130_fd_sc_hd__o21ai_4
X_60436_ _79156_/A _60074_/X _60435_/Y _60436_/Y sky130_fd_sc_hd__o21ai_4
X_47109_ _47109_/A _52859_/B _47109_/Y sky130_fd_sc_hd__nand2_4
X_63155_ _63154_/X _64364_/B _63108_/C _63121_/D _63155_/X sky130_fd_sc_hd__and4_4
X_48089_ _48084_/Y _48055_/X _48088_/X _48089_/Y sky130_fd_sc_hd__a21oi_4
X_60367_ _60267_/X _60367_/B _60367_/C _60367_/D _60367_/Y sky130_fd_sc_hd__nand4_4
X_50120_ _50120_/A _49015_/X _50120_/Y sky130_fd_sc_hd__nand2_4
X_62106_ _59684_/X _62170_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_262_0_CLK clkbuf_9_131_0_CLK/X _83451_/CLK sky130_fd_sc_hd__clkbuf_1
X_67963_ _87897_/Q _67888_/X _67865_/X _67962_/X _67963_/X sky130_fd_sc_hd__a211o_4
X_63086_ _60503_/X _63088_/A sky130_fd_sc_hd__buf_2
X_79949_ _79947_/Y _79948_/Y _79949_/X sky130_fd_sc_hd__xor2_4
X_60298_ _60402_/A _60406_/B _60298_/C _60299_/C sky130_fd_sc_hd__and3_4
Xclkbuf_10_892_0_CLK clkbuf_9_446_0_CLK/X _86139_/CLK sky130_fd_sc_hd__clkbuf_1
X_69702_ _69699_/X _69701_/X _66579_/X _69702_/X sky130_fd_sc_hd__a21o_4
X_50051_ _50049_/Y _50029_/X _50050_/X _86274_/D sky130_fd_sc_hd__a21oi_4
X_66914_ _68392_/A _66915_/A sky130_fd_sc_hd__buf_2
X_62037_ _62094_/B _62037_/X sky130_fd_sc_hd__buf_2
X_82960_ _82769_/CLK _82960_/D _82960_/Q sky130_fd_sc_hd__dfxtp_4
X_67894_ _67657_/X _67992_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_44_0_CLK clkbuf_9_22_0_CLK/X _85049_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_9_383_0_CLK clkbuf_9_382_0_CLK/A clkbuf_9_383_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_81911_ _82005_/CLK _81911_/D _82287_/D sky130_fd_sc_hd__dfxtp_4
X_69633_ _69633_/A _87310_/Q _69633_/X sky130_fd_sc_hd__and2_4
X_66845_ _66823_/A _66845_/B _66845_/X sky130_fd_sc_hd__and2_4
X_82891_ _87926_/CLK _78144_/B _82891_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_277_0_CLK clkbuf_9_138_0_CLK/X _85505_/CLK sky130_fd_sc_hd__clkbuf_1
X_53810_ _52291_/A _53806_/B _53806_/C _53810_/X sky130_fd_sc_hd__and3_4
X_84630_ _84645_/CLK _60333_/Y _79680_/A sky130_fd_sc_hd__dfxtp_4
X_69564_ _69696_/A _69564_/X sky130_fd_sc_hd__buf_2
X_81842_ _81857_/CLK _81842_/D _77468_/A sky130_fd_sc_hd__dfxtp_4
X_54790_ _54790_/A _47526_/Y _54790_/Y sky130_fd_sc_hd__nand2_4
X_66776_ _66773_/X _66775_/X _66726_/X _66776_/X sky130_fd_sc_hd__a21o_4
X_63988_ _64067_/A _64052_/B sky130_fd_sc_hd__buf_2
X_68515_ _83972_/Q _68462_/X _68514_/X _68515_/X sky130_fd_sc_hd__a21bo_4
X_53741_ _53750_/A _48627_/A _53741_/Y sky130_fd_sc_hd__nand2_4
X_65727_ _84182_/Q _65728_/C sky130_fd_sc_hd__inv_2
X_84561_ _84562_/CLK _84561_/D _60810_/C sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_59_0_CLK clkbuf_9_29_0_CLK/X _85037_/CLK sky130_fd_sc_hd__clkbuf_1
X_50953_ _50963_/A _50941_/B _50963_/C _46736_/X _50953_/X sky130_fd_sc_hd__and4_4
X_62939_ _60360_/X _62939_/X sky130_fd_sc_hd__buf_2
X_81773_ _81575_/CLK _76054_/X _81773_/Q sky130_fd_sc_hd__dfxtp_4
X_69495_ _87513_/Q _69442_/X _69396_/X _69494_/X _69495_/X sky130_fd_sc_hd__a211o_4
X_86300_ _86301_/CLK _49917_/Y _72187_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_398_0_CLK clkbuf_9_398_0_CLK/A clkbuf_9_398_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_83512_ _83507_/CLK _83512_/D _83512_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_205_0_CLK clkbuf_8_205_0_CLK/A clkbuf_9_411_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_56460_ _73024_/B _56460_/B _56370_/C _56460_/D _56463_/A sky130_fd_sc_hd__nand4_4
X_80724_ _80676_/CLK _75910_/X _80692_/D sky130_fd_sc_hd__dfxtp_4
X_68446_ _68446_/A _68445_/X _68446_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_200_0_CLK clkbuf_9_100_0_CLK/X _81082_/CLK sky130_fd_sc_hd__clkbuf_1
X_87280_ _88087_/CLK _87280_/D _69179_/B sky130_fd_sc_hd__dfxtp_4
X_53672_ _50447_/A _53666_/X _53692_/C _53672_/X sky130_fd_sc_hd__and3_4
X_65658_ _65503_/X _85586_/Q _65504_/X _65657_/X _65658_/X sky130_fd_sc_hd__a211o_4
X_84492_ _84520_/CLK _84492_/D _84492_/Q sky130_fd_sc_hd__dfxtp_4
X_50884_ _50906_/A _51744_/B _50884_/Y sky130_fd_sc_hd__nand2_4
X_55411_ _55410_/Y _55200_/C _55411_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_830_0_CLK clkbuf_9_415_0_CLK/X _86753_/CLK sky130_fd_sc_hd__clkbuf_1
X_86231_ _86235_/CLK _86231_/D _86231_/Q sky130_fd_sc_hd__dfxtp_4
X_52623_ _52617_/Y _52619_/X _52622_/X _85785_/D sky130_fd_sc_hd__a21oi_4
X_64609_ _66195_/B _64638_/B _84233_/Q _64609_/X sky130_fd_sc_hd__and3_4
X_83443_ _83763_/CLK _83443_/D _83443_/Q sky130_fd_sc_hd__dfxtp_4
X_56391_ _56031_/X _56378_/X _56390_/Y _85212_/D sky130_fd_sc_hd__o21ai_4
X_80655_ _86896_/CLK _80655_/D _80655_/Q sky130_fd_sc_hd__dfxtp_4
X_68377_ _68377_/A _68377_/X sky130_fd_sc_hd__buf_2
X_65589_ _65587_/Y _65529_/X _65588_/X _84191_/D sky130_fd_sc_hd__a21o_4
X_58130_ _57991_/A _58130_/B _58130_/Y sky130_fd_sc_hd__nor2_4
XPHY_305 sky130_fd_sc_hd__decap_3
X_55342_ _44059_/X _55342_/X sky130_fd_sc_hd__buf_2
X_67328_ _84074_/Q _67211_/X _67327_/X _84074_/D sky130_fd_sc_hd__a21bo_4
X_86162_ _83303_/CLK _50641_/Y _86162_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_321_0_CLK clkbuf_8_160_0_CLK/X clkbuf_9_321_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_316 sky130_fd_sc_hd__decap_3
X_52554_ _52552_/Y _52541_/X _52553_/Y _52554_/Y sky130_fd_sc_hd__a21boi_4
X_83374_ _83372_/CLK _71793_/Y _58196_/A sky130_fd_sc_hd__dfxtp_4
XPHY_327 sky130_fd_sc_hd__decap_3
X_80586_ _80580_/A _80580_/B _80585_/Y _80608_/A sky130_fd_sc_hd__a21boi_4
XPHY_338 sky130_fd_sc_hd__decap_3
X_85113_ _85057_/CLK _85113_/D _85113_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_349 sky130_fd_sc_hd__decap_3
X_51505_ _51509_/A _51527_/B _51522_/C _53031_/D _51505_/X sky130_fd_sc_hd__and4_4
X_58061_ _58010_/X _58058_/Y _58060_/Y _58028_/X _58015_/X _58061_/X
+ sky130_fd_sc_hd__o32a_4
Xclkbuf_10_215_0_CLK clkbuf_9_107_0_CLK/X _84620_/CLK sky130_fd_sc_hd__clkbuf_1
X_82325_ _82327_/CLK _77139_/B _82325_/Q sky130_fd_sc_hd__dfxtp_4
X_55273_ _55252_/A _56887_/B _55273_/X sky130_fd_sc_hd__and2_4
X_67259_ _67259_/A _67259_/B _67259_/X sky130_fd_sc_hd__and2_4
X_86093_ _85773_/CLK _86093_/D _86093_/Q sky130_fd_sc_hd__dfxtp_4
X_52485_ _85812_/Q _52470_/X _52484_/Y _52485_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_845_0_CLK clkbuf_9_422_0_CLK/X _82975_/CLK sky130_fd_sc_hd__clkbuf_1
X_57012_ _57010_/Y _57011_/Y _57012_/Y sky130_fd_sc_hd__nor2_4
X_54224_ _85481_/Q _54220_/X _54223_/Y _54224_/Y sky130_fd_sc_hd__o21ai_4
X_85044_ _85075_/CLK _57262_/X _45600_/A sky130_fd_sc_hd__dfxtp_4
X_51436_ _86010_/Q _51429_/X _51435_/Y _51436_/Y sky130_fd_sc_hd__o21ai_4
X_70270_ _70267_/A _70267_/B _83112_/Q _70264_/X _70270_/X sky130_fd_sc_hd__and4_4
X_82256_ _85381_/CLK _82256_/D _82256_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_336_0_CLK clkbuf_8_168_0_CLK/X clkbuf_9_336_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_81207_ _81211_/CLK _75054_/X _48986_/A sky130_fd_sc_hd__dfxtp_4
X_54155_ _53418_/X _54160_/A sky130_fd_sc_hd__buf_2
X_51367_ _51282_/A _51367_/X sky130_fd_sc_hd__buf_2
X_82187_ _84951_/CLK _82187_/D _82187_/Q sky130_fd_sc_hd__dfxtp_4
X_41120_ _41100_/X _40571_/A _41119_/X _41121_/A sky130_fd_sc_hd__o21ai_4
X_53106_ _85696_/Q _53093_/X _53105_/Y _53106_/Y sky130_fd_sc_hd__o21ai_4
X_50318_ _50317_/X _48016_/B _50318_/Y sky130_fd_sc_hd__nand2_4
X_81138_ _82327_/CLK _80762_/Q _40671_/A sky130_fd_sc_hd__dfxtp_4
X_58963_ _58925_/X _85442_/Q _58962_/X _58963_/Y sky130_fd_sc_hd__o21ai_4
X_54086_ _85507_/Q _54067_/X _54085_/Y _54086_/Y sky130_fd_sc_hd__o21ai_4
X_51298_ _51298_/A _46391_/A _51298_/X sky130_fd_sc_hd__and2_4
X_86995_ _86998_/CLK _44700_/Y _86995_/Q sky130_fd_sc_hd__dfxtp_4
X_53037_ _53034_/Y _53028_/X _53036_/X _85709_/D sky130_fd_sc_hd__a21oi_4
X_57914_ _57760_/X _85396_/Q _57913_/X _57914_/Y sky130_fd_sc_hd__o21ai_4
X_41051_ _41050_/X _40987_/X _69415_/B _40989_/X _88287_/D sky130_fd_sc_hd__a2bb2o_4
X_50249_ _50241_/Y _50243_/X _50248_/X _86238_/D sky130_fd_sc_hd__a21oi_4
X_73960_ _73958_/X _73959_/Y _73839_/X _73960_/X sky130_fd_sc_hd__a21o_4
X_85946_ _82206_/CLK _85946_/D _85946_/Q sky130_fd_sc_hd__dfxtp_4
X_81069_ _80817_/CLK _75817_/A _75224_/A sky130_fd_sc_hd__dfxtp_4
X_58894_ _58890_/Y _58893_/Y _58883_/X _58894_/X sky130_fd_sc_hd__a21o_4
X_72911_ _73381_/A _72911_/B _72911_/X sky130_fd_sc_hd__and2_4
X_57845_ _58676_/A _57845_/X sky130_fd_sc_hd__buf_2
X_73891_ _73250_/A _73891_/X sky130_fd_sc_hd__buf_2
X_85877_ _86193_/CLK _85877_/D _85877_/Q sky130_fd_sc_hd__dfxtp_4
X_44810_ _44810_/A _86943_/D sky130_fd_sc_hd__inv_2
X_75630_ _75630_/A _75629_/X _75639_/B sky130_fd_sc_hd__xnor2_4
X_87616_ _88387_/CLK _87616_/D _87616_/Q sky130_fd_sc_hd__dfxtp_4
X_72842_ _72837_/X _72841_/X _72812_/X _72845_/A sky130_fd_sc_hd__a21o_4
X_84828_ _84829_/CLK _84828_/D _84828_/Q sky130_fd_sc_hd__dfxtp_4
X_45790_ _45748_/X _61630_/A _45765_/X _45790_/Y sky130_fd_sc_hd__o21ai_4
X_57776_ _57776_/A _69768_/A sky130_fd_sc_hd__buf_2
X_54988_ _54986_/Y _54971_/X _54987_/X _54988_/Y sky130_fd_sc_hd__a21oi_4
X_59515_ _59876_/B _59521_/A _59557_/A sky130_fd_sc_hd__nor2_4
X_44741_ _41936_/A _44741_/X sky130_fd_sc_hd__buf_2
X_56727_ _56726_/X _56727_/X sky130_fd_sc_hd__buf_2
X_75561_ _75553_/Y _75561_/B _75561_/Y sky130_fd_sc_hd__nand2_4
X_87547_ _87814_/CLK _87547_/D _73374_/A sky130_fd_sc_hd__dfxtp_4
X_41953_ _42025_/A _41953_/X sky130_fd_sc_hd__buf_2
X_53939_ _53937_/Y _53892_/X _53938_/X _85538_/D sky130_fd_sc_hd__a21oi_4
X_84759_ _85485_/CLK _84759_/D _84759_/Q sky130_fd_sc_hd__dfxtp_4
X_72773_ _43115_/Y _72731_/X _56935_/X _72772_/Y _72773_/X sky130_fd_sc_hd__a211o_4
X_77300_ _77300_/A _77301_/B sky130_fd_sc_hd__inv_2
X_74512_ _83050_/Q _74387_/X _74511_/Y _74512_/Y sky130_fd_sc_hd__o21ai_4
X_40904_ _40793_/A _40904_/X sky130_fd_sc_hd__buf_2
X_47460_ _47444_/A _53060_/B _47460_/Y sky130_fd_sc_hd__nand2_4
X_71724_ _70939_/A _71724_/X sky130_fd_sc_hd__buf_2
X_59446_ _59442_/X _83339_/Q _59445_/Y _84731_/D sky130_fd_sc_hd__o21a_4
X_78280_ _78262_/X _78280_/B _78274_/A _78284_/B _78280_/Y sky130_fd_sc_hd__nand4_4
X_44672_ _44672_/A _44672_/Y sky130_fd_sc_hd__inv_2
X_56658_ _83335_/Q _83334_/Q _56700_/C sky130_fd_sc_hd__nand2_4
X_75492_ _75492_/A _75492_/Y sky130_fd_sc_hd__inv_2
X_87478_ _87990_/CLK _43328_/X _87478_/Q sky130_fd_sc_hd__dfxtp_4
X_41884_ _41884_/A _41884_/Y sky130_fd_sc_hd__inv_2
X_46411_ _46411_/A _46412_/B sky130_fd_sc_hd__buf_2
X_77231_ _77230_/Y _77231_/Y sky130_fd_sc_hd__inv_2
X_43623_ _40646_/X _43604_/X _73797_/A _43607_/X _87337_/D sky130_fd_sc_hd__a2bb2o_4
X_55609_ _44116_/B _55641_/A sky130_fd_sc_hd__buf_2
X_74443_ _74442_/X _48538_/Y _74443_/Y sky130_fd_sc_hd__nand2_4
X_86429_ _86246_/CLK _86429_/D _64710_/B sky130_fd_sc_hd__dfxtp_4
X_40835_ _40835_/A _40835_/X sky130_fd_sc_hd__buf_2
X_47391_ _47391_/A _53019_/D sky130_fd_sc_hd__buf_2
X_71655_ _71655_/A _71660_/C sky130_fd_sc_hd__buf_2
X_59377_ _59377_/A _59306_/B _59377_/Y sky130_fd_sc_hd__nor2_4
X_56589_ _56589_/A _56589_/X sky130_fd_sc_hd__buf_2
X_49130_ _49128_/X _48632_/A _49129_/Y _52385_/B sky130_fd_sc_hd__a21o_4
X_46342_ _83649_/Q _53980_/B sky130_fd_sc_hd__inv_2
X_70606_ _70717_/A _70613_/B _74533_/D _70594_/X _70606_/Y sky130_fd_sc_hd__nand4_4
X_58328_ _58328_/A _58328_/X sky130_fd_sc_hd__buf_2
X_77162_ _77163_/A _81921_/Q _77173_/B sky130_fd_sc_hd__or2_4
X_43554_ _40469_/X _43532_/X _87363_/Q _43533_/X _87363_/D sky130_fd_sc_hd__a2bb2o_4
X_74374_ _83079_/Q _72066_/X _74373_/Y _74374_/Y sky130_fd_sc_hd__o21ai_4
X_40766_ _40731_/X _82305_/Q _40765_/X _40767_/A sky130_fd_sc_hd__o21ai_4
X_71586_ _71586_/A _71590_/B _71582_/X _71586_/Y sky130_fd_sc_hd__nor3_4
X_76113_ _76113_/A _76113_/B _76113_/X sky130_fd_sc_hd__xor2_4
X_42505_ _42505_/A _87842_/D sky130_fd_sc_hd__inv_2
X_49061_ _50142_/A _48940_/B _48928_/C _49061_/X sky130_fd_sc_hd__and3_4
X_73325_ _73321_/X _73324_/X _72862_/X _73325_/X sky130_fd_sc_hd__a21o_4
X_46273_ _86751_/Q _46250_/X _46272_/Y _46273_/Y sky130_fd_sc_hd__o21ai_4
X_70537_ _70530_/Y _70554_/A sky130_fd_sc_hd__buf_2
X_58259_ _58259_/A _58268_/B _58259_/Y sky130_fd_sc_hd__nand2_4
X_77093_ _77096_/B _77093_/B _77094_/B sky130_fd_sc_hd__xnor2_4
X_43485_ _43466_/X _43485_/X sky130_fd_sc_hd__buf_2
X_40697_ _40696_/X _40651_/X _88352_/Q _40652_/X _40697_/X sky130_fd_sc_hd__a2bb2o_4
X_48012_ _50314_/A _48069_/B _47919_/X _48012_/X sky130_fd_sc_hd__and3_4
X_45224_ _85260_/Q _45222_/X _45223_/X _45224_/Y sky130_fd_sc_hd__o21ai_4
X_76044_ _76047_/B _76043_/Y _81747_/D sky130_fd_sc_hd__xnor2_4
X_42436_ _40524_/X _42434_/X _87865_/Q _42435_/X _87865_/D sky130_fd_sc_hd__a2bb2o_4
X_61270_ _84492_/Q _60979_/X _61097_/X _61170_/Y _84492_/D sky130_fd_sc_hd__a2bb2oi_4
X_73256_ _87052_/Q _73129_/X _73255_/X _73270_/C sky130_fd_sc_hd__o21ai_4
X_70468_ _71483_/B _71366_/A sky130_fd_sc_hd__buf_2
X_60221_ _60221_/A _60344_/A _60344_/B _60344_/C _60299_/A sky130_fd_sc_hd__nand4_4
X_72207_ _72196_/X _85338_/Q _72120_/X _72207_/X sky130_fd_sc_hd__o21a_4
X_45155_ _83025_/Q _45156_/A sky130_fd_sc_hd__inv_2
X_42367_ _42367_/A _42367_/Y sky130_fd_sc_hd__inv_2
X_73187_ _44189_/X _83065_/Q _73238_/A _73186_/X _73188_/B sky130_fd_sc_hd__a211o_4
X_70399_ DATA_TO_HASH[1] _70400_/A sky130_fd_sc_hd__buf_2
X_44106_ _44104_/Y _86840_/Q _44106_/C _44107_/C sky130_fd_sc_hd__nand3_4
X_79803_ _79796_/X _79798_/B _79803_/Y sky130_fd_sc_hd__nand2_4
X_41318_ _41317_/Y _88237_/D sky130_fd_sc_hd__inv_2
X_60152_ _60152_/A _60153_/C sky130_fd_sc_hd__inv_2
X_72138_ _59255_/A _72277_/A sky130_fd_sc_hd__buf_2
X_49963_ _72294_/B _49960_/X _49962_/Y _49963_/Y sky130_fd_sc_hd__o21ai_4
X_45086_ _45078_/X _45083_/Y _45085_/Y _45086_/Y sky130_fd_sc_hd__a21oi_4
X_42298_ _42276_/A _42298_/X sky130_fd_sc_hd__buf_2
X_77995_ _82079_/Q _77997_/A sky130_fd_sc_hd__inv_2
X_48914_ _48914_/A _48914_/B _50578_/A sky130_fd_sc_hd__nor2_4
X_44037_ _44036_/Y _44037_/X sky130_fd_sc_hd__buf_2
X_79734_ _79732_/X _79739_/B _79734_/Y sky130_fd_sc_hd__xnor2_4
X_41249_ _41184_/X _40727_/A _41248_/X _41249_/Y sky130_fd_sc_hd__o21ai_4
X_64960_ _64955_/X _64958_/X _64959_/X _64960_/X sky130_fd_sc_hd__a21o_4
X_60083_ _62463_/A _60084_/A sky130_fd_sc_hd__buf_2
X_72069_ _83291_/Q _72066_/X _72068_/Y _72069_/Y sky130_fd_sc_hd__o21ai_4
X_76946_ _81376_/D _76946_/B _76946_/X sky130_fd_sc_hd__and2_4
X_49894_ _49892_/Y _49870_/X _49893_/X _49894_/Y sky130_fd_sc_hd__a21oi_4
X_63911_ _63903_/X _63890_/X _63905_/Y _63908_/Y _63910_/X _63911_/X
+ sky130_fd_sc_hd__a41o_4
X_48845_ _48845_/A _48849_/B _48849_/C _48845_/X sky130_fd_sc_hd__and3_4
X_79665_ _79652_/X _79663_/X _79664_/X _79665_/Y sky130_fd_sc_hd__a21oi_4
X_64891_ _64870_/A _64870_/B _64891_/C _64891_/Y sky130_fd_sc_hd__nor3_4
X_76877_ _81498_/Q _81370_/D _76876_/X _76877_/Y sky130_fd_sc_hd__a21oi_4
X_66630_ _66602_/A _86804_/Q _66630_/X sky130_fd_sc_hd__and2_4
X_78616_ _78616_/A _78616_/B _78616_/Y sky130_fd_sc_hd__nor2_4
X_63842_ _63836_/Y _63838_/Y _63840_/Y _63841_/Y _63842_/X sky130_fd_sc_hd__and4_4
X_75828_ _80926_/Q _75830_/A sky130_fd_sc_hd__inv_2
X_48776_ _48774_/Y _48760_/X _48775_/X _86485_/D sky130_fd_sc_hd__a21oi_4
X_79596_ _79580_/A _79580_/B _79575_/Y _79596_/Y sky130_fd_sc_hd__o21ai_4
X_45988_ _45980_/X _45987_/X _40439_/X _86826_/Q _45982_/X _45989_/A
+ sky130_fd_sc_hd__o32ai_4
X_47727_ _47715_/X _53209_/B _47727_/Y sky130_fd_sc_hd__nand2_4
X_66561_ _66560_/X _69582_/A sky130_fd_sc_hd__buf_2
X_78547_ _78547_/A _82674_/D _78547_/Y sky130_fd_sc_hd__nand2_4
X_44939_ _44937_/Y _44939_/B _44939_/X sky130_fd_sc_hd__and2_4
X_63773_ _60867_/Y _64026_/A sky130_fd_sc_hd__buf_2
X_75759_ _75759_/A _75759_/B _75760_/B sky130_fd_sc_hd__xor2_4
X_60985_ _60911_/X _60921_/X _63738_/B _63738_/D _60985_/Y sky130_fd_sc_hd__a22oi_4
X_68300_ _64731_/A _68300_/X sky130_fd_sc_hd__buf_2
X_65512_ _65512_/A _65511_/Y _65512_/Y sky130_fd_sc_hd__nand2_4
X_62724_ _60199_/X _62738_/D sky130_fd_sc_hd__buf_2
X_69280_ _87029_/Q _69277_/X _69278_/X _69279_/X _69280_/X sky130_fd_sc_hd__a211o_4
X_47658_ _54867_/B _53174_/B sky130_fd_sc_hd__buf_2
X_66492_ _66391_/A _66521_/B sky130_fd_sc_hd__buf_2
X_78478_ _78464_/X _78478_/B _78478_/Y sky130_fd_sc_hd__nand2_4
X_68231_ _84006_/Q _68220_/X _68230_/X _84006_/D sky130_fd_sc_hd__a21bo_4
X_46609_ _86721_/Q _46474_/X _46608_/Y _46609_/Y sky130_fd_sc_hd__o21ai_4
X_65443_ _65440_/X _65442_/X _65389_/X _65446_/A sky130_fd_sc_hd__a21o_4
X_77429_ _77428_/X _77431_/B sky130_fd_sc_hd__inv_2
X_62655_ _60204_/A _60156_/Y _62655_/Y sky130_fd_sc_hd__nor2_4
X_47589_ _83706_/Q _47589_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_51_0_CLK clkbuf_7_50_0_CLK/A clkbuf_7_51_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_49328_ _49327_/X _50850_/B _49328_/Y sky130_fd_sc_hd__nand2_4
X_61606_ _61602_/X _61576_/X _61605_/Y _84467_/D sky130_fd_sc_hd__a21oi_4
X_80440_ _59216_/Y _66177_/C _80439_/Y _80458_/A sky130_fd_sc_hd__o21a_4
X_68162_ _68155_/X _67005_/Y _68148_/X _68161_/Y _68162_/X sky130_fd_sc_hd__a211o_4
X_65374_ _65370_/Y _65347_/X _65373_/Y _84204_/D sky130_fd_sc_hd__a21o_4
Xclkbuf_8_191_0_CLK clkbuf_7_95_0_CLK/X clkbuf_9_382_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_62586_ _61655_/A _62566_/B _62501_/X _62597_/D _62586_/Y sky130_fd_sc_hd__nand4_4
X_67113_ _66410_/A _67113_/X sky130_fd_sc_hd__buf_2
X_64325_ _58317_/A _64308_/X _64324_/Y _64325_/Y sky130_fd_sc_hd__o21ai_4
X_49259_ _49263_/A _53993_/B _49259_/Y sky130_fd_sc_hd__nand2_4
X_61537_ _61533_/X _61517_/X _61536_/Y _61537_/Y sky130_fd_sc_hd__a21oi_4
X_80371_ _80371_/A _80371_/B _80372_/B sky130_fd_sc_hd__xor2_4
X_68093_ _66607_/X _66610_/X _67897_/X _68093_/Y sky130_fd_sc_hd__a21oi_4
X_82110_ _82860_/CLK _82110_/D _77208_/A sky130_fd_sc_hd__dfxtp_4
X_67044_ _66947_/X _67030_/Y _67031_/X _67043_/Y _67044_/X sky130_fd_sc_hd__a211o_4
X_52270_ _52126_/A _52271_/A sky130_fd_sc_hd__buf_2
X_64256_ _64315_/A _64301_/B sky130_fd_sc_hd__buf_2
X_83090_ _81627_/CLK _83090_/D _83090_/Q sky130_fd_sc_hd__dfxtp_4
X_61468_ _61468_/A _61468_/B _61467_/X _61451_/D _61468_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_7_66_0_CLK clkbuf_7_67_0_CLK/A clkbuf_7_66_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_51221_ _51217_/Y _51201_/X _51220_/X _51221_/Y sky130_fd_sc_hd__a21oi_4
X_63207_ _63201_/Y _63202_/X _63205_/X _63206_/X _63183_/X _63207_/Y
+ sky130_fd_sc_hd__o41ai_4
X_82041_ _82009_/CLK _77942_/B _82041_/Q sky130_fd_sc_hd__dfxtp_4
X_60419_ _60502_/A _60420_/A sky130_fd_sc_hd__buf_2
X_64187_ _64187_/A _64187_/B _79908_/B _64187_/Y sky130_fd_sc_hd__nor3_4
X_61399_ _84851_/Q _61399_/X sky130_fd_sc_hd__buf_2
X_51152_ _51130_/A _52843_/B _51152_/Y sky130_fd_sc_hd__nand2_4
X_63138_ _63132_/Y _63133_/X _63135_/X _63137_/X _63125_/X _63138_/Y
+ sky130_fd_sc_hd__o41ai_4
X_68995_ _86982_/Q _68948_/X _68993_/X _68994_/X _68995_/X sky130_fd_sc_hd__a211o_4
X_50103_ _50103_/A _48982_/X _50103_/Y sky130_fd_sc_hd__nand2_4
X_85800_ _85800_/CLK _85800_/D _85800_/Q sky130_fd_sc_hd__dfxtp_4
X_51083_ _51191_/A _51084_/A sky130_fd_sc_hd__buf_2
X_55960_ _55691_/A _55960_/B _55960_/X sky130_fd_sc_hd__and2_4
X_67946_ _67782_/X _67934_/Y _67863_/X _67945_/Y _67946_/X sky130_fd_sc_hd__a211o_4
X_63069_ _63069_/A _63081_/B _63081_/C _63033_/D _63069_/X sky130_fd_sc_hd__or4_4
X_86780_ _86814_/CLK _46075_/Y _86780_/Q sky130_fd_sc_hd__dfxtp_4
X_83992_ _82896_/CLK _83992_/D _82640_/D sky130_fd_sc_hd__dfxtp_4
X_50034_ _86277_/Q _50012_/X _50033_/Y _50034_/Y sky130_fd_sc_hd__o21ai_4
X_54911_ _54908_/Y _54909_/X _54910_/X _85355_/D sky130_fd_sc_hd__a21oi_4
X_85731_ _85635_/CLK _52917_/Y _85731_/Q sky130_fd_sc_hd__dfxtp_4
X_82943_ _82925_/CLK _78107_/X _46274_/A sky130_fd_sc_hd__dfxtp_4
X_55891_ _55891_/A _55890_/X _55891_/X sky130_fd_sc_hd__and2_4
X_67877_ _67664_/X _67862_/Y _67863_/X _67876_/Y _67877_/X sky130_fd_sc_hd__a211o_4
X_57630_ _57630_/A _48122_/Y _57630_/Y sky130_fd_sc_hd__nand2_4
X_69616_ _83910_/Q _69564_/X _69615_/X _69616_/X sky130_fd_sc_hd__a21bo_4
X_54842_ _85368_/Q _54839_/X _54841_/Y _54842_/Y sky130_fd_sc_hd__o21ai_4
X_66828_ _66760_/A _66828_/B _66828_/X sky130_fd_sc_hd__and2_4
X_85662_ _85439_/CLK _53285_/Y _85662_/Q sky130_fd_sc_hd__dfxtp_4
X_82874_ _82855_/CLK _78248_/B _82874_/Q sky130_fd_sc_hd__dfxtp_4
X_87401_ _87397_/CLK _87401_/D _87401_/Q sky130_fd_sc_hd__dfxtp_4
X_84613_ _84606_/CLK _60478_/Y _79153_/A sky130_fd_sc_hd__dfxtp_4
X_57561_ _57559_/Y _57543_/X _57560_/Y _84979_/D sky130_fd_sc_hd__a21boi_4
X_81825_ _81695_/CLK _81825_/D _47226_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_144_0_CLK clkbuf_7_72_0_CLK/X clkbuf_8_144_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_69547_ _44022_/X _69547_/B _69547_/X sky130_fd_sc_hd__and2_4
X_88381_ _87116_/CLK _40503_/Y _88381_/Q sky130_fd_sc_hd__dfxtp_4
X_54773_ _85380_/Q _54757_/X _54772_/Y _54773_/Y sky130_fd_sc_hd__o21ai_4
X_66759_ _66758_/X _66759_/X sky130_fd_sc_hd__buf_2
X_85593_ _85593_/CLK _85593_/D _85593_/Q sky130_fd_sc_hd__dfxtp_4
X_51985_ _51947_/A _48231_/B _51985_/Y sky130_fd_sc_hd__nand2_4
X_59300_ _86665_/Q _59226_/B _59300_/Y sky130_fd_sc_hd__nor2_4
X_56512_ _56525_/A _56523_/A sky130_fd_sc_hd__buf_2
X_87332_ _87045_/CLK _87332_/D _73921_/A sky130_fd_sc_hd__dfxtp_4
X_53724_ _53791_/A _48593_/A _53724_/Y sky130_fd_sc_hd__nand2_4
X_84544_ _84549_/CLK _84544_/D _84544_/Q sky130_fd_sc_hd__dfxtp_4
X_50936_ _50819_/X _50936_/X sky130_fd_sc_hd__buf_2
X_57492_ _57490_/Y _47791_/X _57491_/Y _57492_/Y sky130_fd_sc_hd__a21oi_4
X_81756_ _81756_/CLK _76113_/B _41310_/A sky130_fd_sc_hd__dfxtp_4
X_69478_ _69478_/A _69478_/X sky130_fd_sc_hd__buf_2
X_59231_ _57708_/X _59231_/X sky130_fd_sc_hd__buf_2
X_56443_ _56144_/X _56439_/X _56442_/Y _85192_/D sky130_fd_sc_hd__o21ai_4
X_68429_ _68429_/A _68429_/X sky130_fd_sc_hd__buf_2
X_80707_ _81834_/CLK _75893_/X _80675_/D sky130_fd_sc_hd__dfxtp_4
X_87263_ _87273_/CLK _87263_/D _69411_/B sky130_fd_sc_hd__dfxtp_4
X_53655_ _53652_/Y _53653_/X _53654_/X _85594_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_260_0_CLK clkbuf_8_130_0_CLK/X clkbuf_9_260_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_7_19_0_CLK clkbuf_6_9_0_CLK/X clkbuf_8_39_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_84475_ _84477_/CLK _84475_/D _84475_/Q sky130_fd_sc_hd__dfxtp_4
X_50867_ _86117_/Q _50856_/X _50866_/Y _50867_/Y sky130_fd_sc_hd__o21ai_4
X_81687_ _81801_/CLK _81687_/D _81687_/Q sky130_fd_sc_hd__dfxtp_4
X_86214_ _86213_/CLK _50373_/Y _86214_/Q sky130_fd_sc_hd__dfxtp_4
X_40620_ _48461_/A _40620_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_159_0_CLK clkbuf_7_79_0_CLK/X clkbuf_9_318_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_52606_ _52614_/A _52605_/X _52622_/C _51777_/D _52606_/X sky130_fd_sc_hd__and4_4
X_59162_ _59146_/X _85428_/Q _59161_/X _59162_/Y sky130_fd_sc_hd__o21ai_4
X_71440_ _71419_/Y _83498_/Q _71439_/X _71440_/X sky130_fd_sc_hd__a21o_4
X_83426_ _82386_/CLK _71647_/Y _59504_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_154_0_CLK clkbuf_9_77_0_CLK/X _81330_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_102 sky130_fd_sc_hd__decap_3
X_56374_ _56435_/A _56458_/A sky130_fd_sc_hd__buf_2
X_80638_ _41796_/Y _46258_/A _88403_/Q _40354_/X _88403_/D sky130_fd_sc_hd__a2bb2o_4
X_87194_ _87446_/CLK _43932_/Y _67939_/B sky130_fd_sc_hd__dfxtp_4
X_53586_ _53846_/A _53586_/X sky130_fd_sc_hd__buf_2
XPHY_113 sky130_fd_sc_hd__decap_3
X_50798_ _50796_/Y _50792_/X _50797_/Y _50798_/Y sky130_fd_sc_hd__a21boi_4
XPHY_124 sky130_fd_sc_hd__decap_3
X_58113_ _57947_/X _85700_/Q _57948_/X _58113_/X sky130_fd_sc_hd__o21a_4
XPHY_135 sky130_fd_sc_hd__decap_3
Xclkbuf_10_784_0_CLK clkbuf_9_392_0_CLK/X _82803_/CLK sky130_fd_sc_hd__clkbuf_1
X_55325_ _55322_/X _55324_/X _83750_/Q _55325_/X sky130_fd_sc_hd__a21o_4
X_86145_ _86145_/CLK _86145_/D _86145_/Q sky130_fd_sc_hd__dfxtp_4
X_52537_ _52487_/X _49322_/B _52537_/Y sky130_fd_sc_hd__nand2_4
XPHY_146 sky130_fd_sc_hd__decap_3
X_40551_ _43175_/B _40591_/C sky130_fd_sc_hd__inv_2
X_71371_ _71163_/A _71342_/B _71372_/A sky130_fd_sc_hd__nor2_4
X_59093_ _59029_/A _86361_/Q _59093_/Y sky130_fd_sc_hd__nor2_4
X_83357_ _83421_/CLK _83357_/D _83357_/Q sky130_fd_sc_hd__dfxtp_4
X_80569_ _80567_/X _80569_/B _80570_/B sky130_fd_sc_hd__xnor2_4
XPHY_157 sky130_fd_sc_hd__decap_3
XPHY_168 sky130_fd_sc_hd__decap_3
X_73110_ _73107_/X _73109_/X _72982_/X _73110_/X sky130_fd_sc_hd__a21o_4
XPHY_179 sky130_fd_sc_hd__decap_3
X_58044_ _57966_/X _85706_/Q _58020_/X _58044_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_9_275_0_CLK clkbuf_9_274_0_CLK/A clkbuf_9_275_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_70322_ _70320_/X _74782_/B _70321_/X _83798_/D sky130_fd_sc_hd__a21o_4
X_82308_ _81179_/CLK _77016_/Y _82308_/Q sky130_fd_sc_hd__dfxtp_4
X_43270_ _43260_/X _43269_/X _41116_/X _87507_/Q _43250_/X _43270_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55256_ _55135_/A _85001_/Q _55256_/X sky130_fd_sc_hd__and2_4
X_74090_ _74090_/A _74090_/B _74090_/Y sky130_fd_sc_hd__nand2_4
X_86076_ _85757_/CLK _86076_/D _86076_/Q sky130_fd_sc_hd__dfxtp_4
X_40482_ _40481_/Y _88385_/D sky130_fd_sc_hd__inv_2
X_52468_ _52468_/A _52468_/B _52468_/Y sky130_fd_sc_hd__nand2_4
X_83288_ _85542_/CLK _83288_/D _83288_/Q sky130_fd_sc_hd__dfxtp_4
X_42221_ _41367_/X _42209_/X _87972_/Q _42210_/X _42221_/X sky130_fd_sc_hd__a2bb2o_4
X_54207_ _53282_/A _54316_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_169_0_CLK clkbuf_9_84_0_CLK/X _81582_/CLK sky130_fd_sc_hd__clkbuf_1
X_73041_ _72870_/X _86199_/Q _72905_/X _73040_/X _73041_/X sky130_fd_sc_hd__a211o_4
X_85027_ _85031_/CLK _85027_/D _85027_/Q sky130_fd_sc_hd__dfxtp_4
X_51419_ _86013_/Q _51402_/X _51418_/Y _51419_/Y sky130_fd_sc_hd__o21ai_4
X_70253_ _70260_/A _70260_/B _83182_/Q _70260_/D _70253_/X sky130_fd_sc_hd__and4_4
X_82239_ _82531_/CLK _82271_/Q _82239_/Q sky130_fd_sc_hd__dfxtp_4
X_55187_ _85101_/Q _55145_/A _44044_/X _55186_/Y _55187_/X sky130_fd_sc_hd__a211o_4
X_52399_ _52630_/A _52602_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_799_0_CLK clkbuf_9_399_0_CLK/X _84111_/CLK sky130_fd_sc_hd__clkbuf_1
X_42152_ _41165_/X _42148_/X _88009_/Q _42150_/X _88009_/D sky130_fd_sc_hd__a2bb2o_4
X_54138_ _54135_/Y _54117_/X _54137_/X _54138_/Y sky130_fd_sc_hd__a21oi_4
X_70184_ _70169_/X _83845_/Q _70183_/X _83845_/D sky130_fd_sc_hd__a21o_4
X_59995_ _59995_/A _59995_/X sky130_fd_sc_hd__buf_2
X_41103_ _41100_/X _81699_/Q _41102_/X _41104_/A sky130_fd_sc_hd__o21ai_4
X_76800_ _76795_/Y _76800_/B _76801_/B sky130_fd_sc_hd__nand2_4
X_46960_ _86685_/Q _46955_/X _46959_/Y _46960_/Y sky130_fd_sc_hd__o21ai_4
X_42083_ _42083_/A _42083_/X sky130_fd_sc_hd__buf_2
X_58946_ _84787_/Q _58946_/Y sky130_fd_sc_hd__inv_2
X_54069_ _54068_/X _54069_/B _54069_/Y sky130_fd_sc_hd__nand2_4
X_77780_ _81927_/D _77780_/B _77780_/X sky130_fd_sc_hd__and2_4
X_74992_ _74986_/X _75001_/A _74993_/B sky130_fd_sc_hd__xor2_4
X_86978_ _82538_/CLK _86978_/D _44745_/A sky130_fd_sc_hd__dfxtp_4
X_45911_ _44184_/X _57673_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_722_0_CLK clkbuf_9_361_0_CLK/X _87011_/CLK sky130_fd_sc_hd__clkbuf_1
X_41034_ _41034_/A _41019_/B _41034_/X sky130_fd_sc_hd__or2_4
X_76731_ _76724_/Y _76725_/A _76730_/Y _76731_/Y sky130_fd_sc_hd__a21oi_4
X_73943_ _43070_/Y _72900_/X _73894_/X _73942_/Y _73943_/X sky130_fd_sc_hd__a211o_4
X_85929_ _86089_/CLK _51883_/Y _85929_/Q sky130_fd_sc_hd__dfxtp_4
X_46891_ _47081_/A _46891_/X sky130_fd_sc_hd__buf_2
X_58877_ _58877_/A _58877_/X sky130_fd_sc_hd__buf_2
X_48630_ _81769_/Q _48632_/A sky130_fd_sc_hd__inv_2
X_79450_ _79438_/A _79438_/B _79450_/Y sky130_fd_sc_hd__nor2_4
X_45842_ _85092_/Q _45842_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_9_213_0_CLK clkbuf_8_106_0_CLK/X clkbuf_9_213_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_57828_ _57726_/X _86011_/Q _57827_/X _57828_/Y sky130_fd_sc_hd__o21ai_4
X_76662_ _76662_/A _76658_/Y _76662_/C _76662_/Y sky130_fd_sc_hd__nand3_4
X_73874_ _68695_/B _73872_/X _73772_/X _73873_/Y _73874_/X sky130_fd_sc_hd__a211o_4
X_78401_ _82504_/Q _82760_/D _78401_/X sky130_fd_sc_hd__xor2_4
X_75613_ _75621_/A _80775_/D _75616_/A sky130_fd_sc_hd__xnor2_4
Xclkbuf_10_107_0_CLK clkbuf_9_53_0_CLK/X _87178_/CLK sky130_fd_sc_hd__clkbuf_1
X_48561_ _48604_/A _48561_/B _48561_/Y sky130_fd_sc_hd__nand2_4
X_72825_ _42550_/A _73000_/B _72825_/Y sky130_fd_sc_hd__nor2_4
X_79381_ _79375_/Y _79381_/B _82836_/D sky130_fd_sc_hd__xor2_4
X_45773_ _45770_/X _45772_/Y _45757_/X _45773_/X sky130_fd_sc_hd__a21o_4
X_57759_ _57837_/A _57759_/X sky130_fd_sc_hd__buf_2
X_76593_ _76593_/A _76593_/Y sky130_fd_sc_hd__inv_2
X_42985_ _41992_/A _42985_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_737_0_CLK clkbuf_9_368_0_CLK/X _87990_/CLK sky130_fd_sc_hd__clkbuf_1
X_47512_ _47511_/Y _53090_/D sky130_fd_sc_hd__buf_2
X_78332_ _78332_/A _78332_/Y sky130_fd_sc_hd__inv_2
X_44724_ _44723_/Y _44724_/Y sky130_fd_sc_hd__inv_2
X_75544_ _75540_/X _75543_/X _75544_/X sky130_fd_sc_hd__xor2_4
X_41936_ _41936_/A _41998_/A sky130_fd_sc_hd__buf_2
X_48492_ _53678_/B _52158_/B sky130_fd_sc_hd__buf_2
X_72756_ _44124_/A _72757_/A sky130_fd_sc_hd__buf_2
X_60770_ _60770_/A _63696_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_228_0_CLK clkbuf_8_114_0_CLK/X clkbuf_9_228_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_47443_ _47442_/Y _53050_/B sky130_fd_sc_hd__buf_2
X_71707_ _58303_/Y _71695_/X _71706_/Y _83403_/D sky130_fd_sc_hd__o21ai_4
X_59429_ _59426_/X _59427_/Y _59428_/Y _84736_/D sky130_fd_sc_hd__a21oi_4
X_78263_ _78263_/A _78263_/B _78280_/B sky130_fd_sc_hd__and2_4
X_44655_ _44655_/A _44655_/Y sky130_fd_sc_hd__inv_2
X_75475_ _75475_/A _75475_/B _75475_/Y sky130_fd_sc_hd__nand2_4
X_41867_ _42429_/A _41992_/A sky130_fd_sc_hd__buf_2
X_72687_ _72687_/A _72697_/A sky130_fd_sc_hd__buf_2
X_77214_ _82111_/Q _77214_/B _77214_/X sky130_fd_sc_hd__xor2_4
X_43606_ _43606_/A _43607_/A sky130_fd_sc_hd__buf_2
XPHY_4 sky130_fd_sc_hd__decap_3
X_62440_ _62214_/A _62440_/X sky130_fd_sc_hd__buf_2
X_74426_ _48498_/A _74420_/X _74425_/X _74426_/X sky130_fd_sc_hd__and3_4
X_40818_ _82870_/Q _40779_/B _40818_/X sky130_fd_sc_hd__or2_4
X_47374_ _47333_/X _53012_/B _47374_/Y sky130_fd_sc_hd__nand2_4
X_71638_ _59488_/Y _71628_/X _71637_/Y _71638_/Y sky130_fd_sc_hd__o21ai_4
X_78194_ _78193_/Y _78191_/C _78194_/X sky130_fd_sc_hd__and2_4
X_44586_ _44586_/A _87044_/D sky130_fd_sc_hd__inv_2
X_41798_ _41797_/X _41750_/X _66583_/B _41751_/X _88147_/D sky130_fd_sc_hd__a2bb2o_4
X_49113_ _50677_/A _49113_/B _49091_/C _49113_/X sky130_fd_sc_hd__and3_4
X_46325_ _53971_/B _50757_/B sky130_fd_sc_hd__buf_2
X_77145_ _77142_/Y _77144_/X _77146_/B sky130_fd_sc_hd__nand2_4
X_43537_ _40418_/X _43532_/X _87370_/Q _43533_/X _87370_/D sky130_fd_sc_hd__a2bb2o_4
X_74357_ _45954_/X _58334_/A _56163_/A _74357_/Y sky130_fd_sc_hd__nand3_4
X_62371_ _62344_/X _57664_/X _62315_/C _62355_/X _62371_/X sky130_fd_sc_hd__and4_4
X_40749_ _40748_/Y _40749_/X sky130_fd_sc_hd__buf_2
X_71569_ _71557_/X _83453_/Q _71568_/Y _71569_/X sky130_fd_sc_hd__a21o_4
X_64110_ _58970_/A _64102_/B _64110_/Y sky130_fd_sc_hd__nor2_4
X_49044_ _49044_/A _53860_/B sky130_fd_sc_hd__inv_2
X_61322_ _61321_/Y _61323_/B sky130_fd_sc_hd__buf_2
X_73308_ _73210_/X _85580_/Q _73284_/X _73307_/X _73308_/X sky130_fd_sc_hd__a211o_4
X_46256_ _46272_/A _49212_/B _46256_/Y sky130_fd_sc_hd__nand2_4
XPHY_680 sky130_fd_sc_hd__decap_3
X_65090_ _65090_/A _65089_/Y _65090_/Y sky130_fd_sc_hd__nand2_4
X_77076_ _81997_/Q _82285_/D _77086_/B sky130_fd_sc_hd__nand2_4
X_43468_ _41651_/X _43465_/X _87407_/Q _43467_/X _87407_/D sky130_fd_sc_hd__a2bb2o_4
X_74288_ _72686_/A _74288_/X sky130_fd_sc_hd__buf_2
XPHY_691 sky130_fd_sc_hd__decap_3
X_45207_ _56341_/C _45206_/X _45161_/X _45207_/X sky130_fd_sc_hd__o21a_4
X_64041_ _60930_/C _64091_/D sky130_fd_sc_hd__buf_2
X_76027_ _81713_/D _76027_/B _76028_/B sky130_fd_sc_hd__nand2_4
X_42419_ _42419_/A _42419_/Y sky130_fd_sc_hd__inv_2
X_61253_ _61153_/C _61271_/A _61202_/B _61254_/D sky130_fd_sc_hd__o21ai_4
X_73239_ _73239_/A _86511_/Q _73239_/X sky130_fd_sc_hd__and2_4
X_46187_ _46187_/A _74842_/B sky130_fd_sc_hd__buf_2
X_43399_ _43296_/A _43399_/X sky130_fd_sc_hd__buf_2
X_60204_ _60204_/A _60288_/C sky130_fd_sc_hd__buf_2
X_45138_ _45133_/Y _45136_/Y _45137_/X _45138_/X sky130_fd_sc_hd__a21o_4
X_61184_ _84513_/Q _60979_/X _61176_/Y _61183_/Y _84513_/D sky130_fd_sc_hd__a2bb2oi_4
X_67800_ _67794_/X _67797_/X _67799_/X _67800_/X sky130_fd_sc_hd__a21o_4
X_60135_ _60134_/X _84656_/D sky130_fd_sc_hd__inv_2
X_49946_ _72251_/B _49934_/X _49945_/Y _49946_/Y sky130_fd_sc_hd__o21ai_4
X_45069_ _64334_/B _61447_/B sky130_fd_sc_hd__buf_2
X_68780_ _43070_/A _68778_/X _68552_/X _68779_/X _68780_/X sky130_fd_sc_hd__a211o_4
X_65992_ _65992_/A _73707_/B _65992_/X sky130_fd_sc_hd__and2_4
X_77978_ _77975_/Y _77977_/Y _77980_/C sky130_fd_sc_hd__nor2_4
X_67731_ _67728_/X _67730_/X _67681_/X _67731_/X sky130_fd_sc_hd__a21o_4
X_79717_ _79703_/Y _79708_/Y _79716_/X _79717_/Y sky130_fd_sc_hd__o21ai_4
X_64943_ _64938_/Y _64939_/X _64942_/Y _84221_/D sky130_fd_sc_hd__a21o_4
X_60066_ _59842_/A _60081_/A sky130_fd_sc_hd__buf_2
X_76929_ _81680_/Q _76929_/B _76945_/A sky130_fd_sc_hd__xnor2_4
X_49877_ _49893_/A _49884_/B _49893_/C _53090_/D _49877_/X sky130_fd_sc_hd__and4_4
X_48828_ _48853_/A _48849_/C sky130_fd_sc_hd__buf_2
X_67662_ _67522_/X _67649_/Y _67624_/X _67661_/Y _67662_/X sky130_fd_sc_hd__a211o_4
X_79648_ _84211_/Q _83259_/Q _79648_/X sky130_fd_sc_hd__xor2_4
X_64874_ _64804_/A _64874_/B _64874_/X sky130_fd_sc_hd__and2_4
X_69401_ _69322_/A _69401_/B _69401_/X sky130_fd_sc_hd__and2_4
X_66613_ _84104_/Q _59803_/X _66612_/X _84104_/D sky130_fd_sc_hd__a21bo_4
X_63825_ _61811_/X _63860_/B _63860_/C _63860_/D _63825_/Y sky130_fd_sc_hd__nand4_4
X_48759_ _48759_/A _48840_/A sky130_fd_sc_hd__buf_2
X_67593_ _87976_/Q _67591_/X _67524_/X _67592_/X _67593_/X sky130_fd_sc_hd__a211o_4
X_79579_ _79547_/Y _79561_/Y _79559_/Y _79580_/B sky130_fd_sc_hd__a21oi_4
X_81610_ _83184_/CLK _81610_/D _81802_/D sky130_fd_sc_hd__dfxtp_4
X_69332_ _69236_/A _69332_/B _69332_/X sky130_fd_sc_hd__and2_4
X_66544_ _68999_/A _66544_/B _66544_/X sky130_fd_sc_hd__and2_4
X_51770_ _51779_/A _51770_/B _51770_/Y sky130_fd_sc_hd__nand2_4
X_63756_ _64045_/A _64192_/D sky130_fd_sc_hd__buf_2
X_82590_ _82671_/CLK _82622_/Q _82590_/Q sky130_fd_sc_hd__dfxtp_4
X_60968_ _60950_/Y _60993_/B _60967_/X _60968_/X sky130_fd_sc_hd__a21o_4
X_50721_ _50657_/A _50721_/B _50721_/Y sky130_fd_sc_hd__nand2_4
X_62707_ _62705_/X _62652_/X _62706_/Y _62707_/Y sky130_fd_sc_hd__a21oi_4
X_81541_ _81412_/CLK _76682_/X _81541_/Q sky130_fd_sc_hd__dfxtp_4
X_69263_ _87530_/Q _69261_/X _69248_/X _69262_/X _69263_/X sky130_fd_sc_hd__a211o_4
X_66475_ _66411_/A _66475_/X sky130_fd_sc_hd__buf_2
X_63687_ _58360_/A _63416_/A _63661_/C _63699_/D _63687_/Y sky130_fd_sc_hd__nand4_4
X_60899_ _60881_/Y _61036_/C _60897_/Y _84553_/Q _60898_/X _60899_/X
+ sky130_fd_sc_hd__o32a_4
X_68214_ _68196_/X _67316_/Y _68207_/X _68213_/Y _68214_/X sky130_fd_sc_hd__a211o_4
X_53440_ _53435_/Y _53437_/X _53439_/X _53440_/Y sky130_fd_sc_hd__a21oi_4
X_65426_ _65272_/X _85601_/Q _65326_/X _65425_/X _65426_/X sky130_fd_sc_hd__a211o_4
X_84260_ _84314_/CLK _84260_/D _84260_/Q sky130_fd_sc_hd__dfxtp_4
X_50652_ _50142_/A _50651_/X _50568_/C _50652_/X sky130_fd_sc_hd__and3_4
X_62638_ _59478_/A _60337_/C _62638_/Y sky130_fd_sc_hd__nor2_4
X_81472_ _81322_/CLK _76938_/X _81440_/D sky130_fd_sc_hd__dfxtp_4
X_69194_ _87535_/Q _69044_/X _68979_/X _69193_/X _69194_/X sky130_fd_sc_hd__a211o_4
X_83211_ _83216_/CLK _72627_/Y _79168_/A sky130_fd_sc_hd__dfxtp_4
X_80423_ _80423_/A _80423_/B _80436_/B sky130_fd_sc_hd__xnor2_4
X_68145_ _66918_/X _66921_/X _68133_/X _68145_/Y sky130_fd_sc_hd__a21oi_4
X_53371_ _53371_/A _53371_/B _53371_/C _52857_/D _53371_/X sky130_fd_sc_hd__and4_4
X_65357_ _65408_/A _65357_/B _65357_/X sky130_fd_sc_hd__and2_4
X_84191_ _84192_/CLK _84191_/D _84191_/Q sky130_fd_sc_hd__dfxtp_4
X_50583_ _86173_/Q _50563_/X _50582_/Y _50583_/Y sky130_fd_sc_hd__o21ai_4
X_62569_ _62622_/A _62569_/B _62569_/C _62569_/D _62569_/Y sky130_fd_sc_hd__nand4_4
X_55110_ _55118_/A _47798_/A _55110_/Y sky130_fd_sc_hd__nand2_4
X_52322_ _52322_/A _52515_/A sky130_fd_sc_hd__buf_2
X_64308_ _64249_/A _64308_/X sky130_fd_sc_hd__buf_2
X_83142_ _83115_/CLK _73648_/Y _83142_/Q sky130_fd_sc_hd__dfxtp_4
X_56090_ _56089_/X _56098_/A sky130_fd_sc_hd__buf_2
X_80354_ _80338_/Y _80334_/Y _80336_/Y _80354_/Y sky130_fd_sc_hd__a21boi_4
X_68076_ _86944_/Q _68023_/X _68024_/X _68075_/X _68077_/B sky130_fd_sc_hd__a211o_4
X_65288_ _65283_/X _65286_/X _65287_/X _65288_/X sky130_fd_sc_hd__a21o_4
X_55041_ _55037_/A _47679_/A _55041_/Y sky130_fd_sc_hd__nand2_4
X_67027_ _67020_/X _67024_/X _67026_/X _67027_/X sky130_fd_sc_hd__a21o_4
X_52253_ _48702_/A _52267_/B _52267_/C _52253_/X sky130_fd_sc_hd__and3_4
X_64239_ _64234_/X _64235_/X _64236_/X _64238_/Y _64229_/X _64239_/X
+ sky130_fd_sc_hd__o41a_4
X_83073_ _83584_/CLK _83073_/D _83073_/Q sky130_fd_sc_hd__dfxtp_4
X_87950_ _87950_/CLK _42265_/X _87950_/Q sky130_fd_sc_hd__dfxtp_4
X_80285_ _80283_/Y _80284_/Y _80286_/B sky130_fd_sc_hd__nand2_4
X_51204_ _51200_/Y _51201_/X _51203_/X _51204_/Y sky130_fd_sc_hd__a21oi_4
X_86901_ _85177_/CLK _45072_/Y _64334_/B sky130_fd_sc_hd__dfxtp_4
X_82024_ _81989_/CLK _77785_/B _81992_/D sky130_fd_sc_hd__dfxtp_4
X_52184_ _52438_/A _52184_/X sky130_fd_sc_hd__buf_2
X_87881_ _87625_/CLK _87881_/D _87881_/Q sky130_fd_sc_hd__dfxtp_4
X_58800_ _58763_/A _58800_/B _58800_/Y sky130_fd_sc_hd__nor2_4
X_51135_ _86067_/Q _51128_/X _51134_/Y _51135_/Y sky130_fd_sc_hd__o21ai_4
X_86832_ _87225_/CLK _86832_/D _86832_/Q sky130_fd_sc_hd__dfxtp_4
X_59780_ _59780_/A _59780_/Y sky130_fd_sc_hd__inv_2
X_56992_ _56991_/Y _56994_/D sky130_fd_sc_hd__buf_2
X_68978_ _87994_/Q _68975_/X _68976_/X _68977_/X _68978_/X sky130_fd_sc_hd__a211o_4
X_58731_ _58730_/X _85940_/Q _58679_/X _58731_/X sky130_fd_sc_hd__o21a_4
X_51066_ _51013_/A _51071_/B sky130_fd_sc_hd__buf_2
X_67929_ _67955_/A _67929_/B _67929_/X sky130_fd_sc_hd__and2_4
X_55943_ _44085_/C _55943_/B _55943_/X sky130_fd_sc_hd__and2_4
X_86763_ _80672_/CLK _86763_/D _46186_/A sky130_fd_sc_hd__dfxtp_4
X_83975_ _80961_/CLK _68435_/X _83975_/Q sky130_fd_sc_hd__dfxtp_4
X_50017_ _50015_/Y _50003_/X _50016_/X _86281_/D sky130_fd_sc_hd__a21oi_4
X_85714_ _84757_/CLK _53009_/Y _85714_/Q sky130_fd_sc_hd__dfxtp_4
X_70940_ _70942_/A _70940_/B _70947_/C _70940_/Y sky130_fd_sc_hd__nand3_4
X_58662_ _58653_/Y _58624_/X _58658_/X _58661_/X _84810_/D sky130_fd_sc_hd__a22oi_4
X_82926_ _81198_/CLK _78218_/X _82926_/Q sky130_fd_sc_hd__dfxtp_4
X_55874_ _55843_/A _55874_/B _55874_/X sky130_fd_sc_hd__and2_4
X_86694_ _86695_/CLK _86694_/D _86694_/Q sky130_fd_sc_hd__dfxtp_4
X_57613_ _57608_/X _50356_/B _57613_/Y sky130_fd_sc_hd__nand2_4
X_54825_ _54825_/A _54843_/B _54831_/C _53133_/D _54825_/X sky130_fd_sc_hd__and4_4
X_85645_ _85645_/CLK _85645_/D _85645_/Q sky130_fd_sc_hd__dfxtp_4
X_70871_ _70871_/A _70869_/B _70869_/C _70869_/D _70871_/Y sky130_fd_sc_hd__nand4_4
X_58593_ _58591_/X _85471_/Q _58592_/X _58593_/Y sky130_fd_sc_hd__o21ai_4
X_82857_ _82349_/CLK _78124_/B _82857_/Q sky130_fd_sc_hd__dfxtp_4
X_72610_ _72537_/B _72549_/B _61112_/X _72610_/X sky130_fd_sc_hd__a21bo_4
X_57544_ _57531_/A _53516_/B _57544_/Y sky130_fd_sc_hd__nand2_4
X_81808_ _81808_/CLK _81808_/D _81808_/Q sky130_fd_sc_hd__dfxtp_4
X_88364_ _88363_/CLK _88364_/D _88364_/Q sky130_fd_sc_hd__dfxtp_4
X_42770_ _41306_/X _42767_/X _67437_/B _42768_/X _42770_/X sky130_fd_sc_hd__a2bb2o_4
X_54756_ _54751_/Y _54747_/X _54755_/X _85384_/D sky130_fd_sc_hd__a21oi_4
X_73590_ _73590_/A _73589_/X _73591_/B sky130_fd_sc_hd__nand2_4
X_85576_ _86500_/CLK _53749_/Y _85576_/Q sky130_fd_sc_hd__dfxtp_4
X_51968_ _51941_/A _53488_/B _51968_/Y sky130_fd_sc_hd__nand2_4
X_82788_ _83238_/CLK _82820_/Q _78331_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_1009_0_CLK clkbuf_9_504_0_CLK/X _83307_/CLK sky130_fd_sc_hd__clkbuf_1
X_87315_ _83153_/CLK _43678_/X _87315_/Q sky130_fd_sc_hd__dfxtp_4
X_41721_ _41720_/Y _41721_/X sky130_fd_sc_hd__buf_2
X_53707_ _53778_/A _52188_/B _53707_/Y sky130_fd_sc_hd__nand2_4
X_72541_ _72540_/Y _72579_/B sky130_fd_sc_hd__inv_2
X_84527_ _84287_/CLK _84527_/D _76975_/A sky130_fd_sc_hd__dfxtp_4
X_50919_ _50941_/A _50919_/B _50897_/X _50919_/D _50919_/X sky130_fd_sc_hd__and4_4
X_57475_ _56649_/X _74139_/A sky130_fd_sc_hd__buf_2
X_81739_ _81783_/CLK _81739_/D _41743_/B sky130_fd_sc_hd__dfxtp_4
X_88295_ _87790_/CLK _41006_/Y _88295_/Q sky130_fd_sc_hd__dfxtp_4
X_54687_ _54682_/A _47344_/A _54687_/Y sky130_fd_sc_hd__nand2_4
X_51899_ _51896_/Y _51877_/X _51898_/X _51899_/Y sky130_fd_sc_hd__a21oi_4
X_59214_ _59152_/X _59212_/Y _59213_/Y _59169_/X _59156_/X _59214_/X
+ sky130_fd_sc_hd__o32a_4
X_56426_ _56439_/A _56426_/X sky130_fd_sc_hd__buf_2
X_44440_ _44439_/Y _87107_/D sky130_fd_sc_hd__inv_2
X_75260_ _75258_/X _75259_/Y _75261_/B sky130_fd_sc_hd__and2_4
X_87246_ _87249_/CLK _43830_/Y _87246_/Q sky130_fd_sc_hd__dfxtp_4
X_53638_ _53611_/X _74383_/B _53638_/Y sky130_fd_sc_hd__nand2_4
X_41652_ _41651_/X _41638_/X _67434_/B _41639_/X _88175_/D sky130_fd_sc_hd__a2bb2o_4
X_72472_ _86595_/Q _72401_/B _72472_/Y sky130_fd_sc_hd__nor2_4
X_84458_ _84458_/CLK _61701_/Y _84458_/Q sky130_fd_sc_hd__dfxtp_4
X_74211_ _74208_/X _74210_/Y _74211_/Y sky130_fd_sc_hd__nand2_4
X_40603_ _47943_/A _82877_/Q _40603_/X sky130_fd_sc_hd__or2_4
X_59145_ _72358_/A _59145_/X sky130_fd_sc_hd__buf_2
X_71423_ _71420_/X _83505_/Q _71422_/X _83505_/D sky130_fd_sc_hd__a21o_4
X_83409_ _83338_/CLK _83409_/D _83409_/Q sky130_fd_sc_hd__dfxtp_4
X_44371_ _44350_/X _44351_/X _41762_/X _87142_/Q _44353_/X _44372_/A
+ sky130_fd_sc_hd__o32ai_4
X_56357_ _56148_/X _56350_/X _56356_/Y _85223_/D sky130_fd_sc_hd__o21ai_4
X_75191_ _75189_/X _75190_/Y _75217_/A sky130_fd_sc_hd__nand2_4
X_41583_ _41580_/X _41581_/X _67128_/B _41582_/X _88188_/D sky130_fd_sc_hd__a2bb2o_4
X_87177_ _87174_/CLK _87177_/D _43971_/A sky130_fd_sc_hd__dfxtp_4
X_53569_ _53671_/A _53620_/C sky130_fd_sc_hd__buf_2
X_84389_ _84555_/CLK _62707_/Y _84389_/Q sky130_fd_sc_hd__dfxtp_4
X_46110_ _46092_/X _46162_/B sky130_fd_sc_hd__inv_2
X_43322_ _41250_/X _43300_/X _87482_/Q _43302_/X _87482_/D sky130_fd_sc_hd__a2bb2o_4
X_55308_ _45673_/A _55305_/X _44045_/X _55307_/Y _55308_/X sky130_fd_sc_hd__a211o_4
X_74142_ _88346_/Q _73633_/X _73028_/X _74142_/Y sky130_fd_sc_hd__o21ai_4
X_86128_ _86139_/CLK _50813_/Y _86128_/Q sky130_fd_sc_hd__dfxtp_4
X_40534_ _40534_/A _88375_/D sky130_fd_sc_hd__inv_2
X_59076_ _59072_/Y _59075_/Y _59053_/X _59076_/X sky130_fd_sc_hd__a21o_4
X_47090_ _59226_/A _47050_/X _47089_/Y _47090_/Y sky130_fd_sc_hd__o21ai_4
X_71354_ _71504_/C _71351_/X _71424_/C _71363_/D _71354_/X sky130_fd_sc_hd__and4_4
X_56288_ _56284_/X _55987_/X _56287_/Y _85249_/D sky130_fd_sc_hd__o21ai_4
X_58027_ _86635_/Q _58039_/B _58027_/Y sky130_fd_sc_hd__nor2_4
X_70305_ _70303_/X _83804_/Q _70304_/X _83804_/D sky130_fd_sc_hd__a21o_4
X_46041_ _41502_/Y _46029_/X _66765_/B _46030_/X _86798_/D sky130_fd_sc_hd__a2bb2o_4
X_43253_ _41059_/X _43247_/X _87517_/Q _43248_/X _87517_/D sky130_fd_sc_hd__a2bb2o_4
X_55239_ _55243_/B _55240_/B sky130_fd_sc_hd__inv_2
X_78950_ _78948_/Y _79115_/A _78957_/A sky130_fd_sc_hd__xor2_4
X_86059_ _85741_/CLK _51182_/Y _86059_/Q sky130_fd_sc_hd__dfxtp_4
X_74073_ _72978_/A _74073_/X sky130_fd_sc_hd__buf_2
X_40465_ _40784_/A _40932_/A sky130_fd_sc_hd__buf_2
X_71285_ _71041_/X _71268_/A _71279_/C _70638_/A _71285_/Y sky130_fd_sc_hd__nand4_4
X_42204_ _43161_/A _42204_/X sky130_fd_sc_hd__buf_2
X_77901_ _77899_/Y _77900_/Y _77904_/A sky130_fd_sc_hd__xor2_4
X_73024_ _73024_/A _73024_/B _73024_/Y sky130_fd_sc_hd__nor2_4
X_70236_ _70239_/A _70239_/B _70236_/C _70239_/D _70236_/X sky130_fd_sc_hd__and4_4
X_43184_ _43217_/A _43185_/A sky130_fd_sc_hd__buf_2
X_78881_ _78881_/A _78880_/Y _78882_/B sky130_fd_sc_hd__xor2_4
X_40396_ _57491_/A _40364_/X _40395_/X _88398_/Q _40375_/X _40396_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49800_ _49809_/A _53012_/B _49800_/Y sky130_fd_sc_hd__nand2_4
X_42135_ _42134_/Y _42135_/Y sky130_fd_sc_hd__inv_2
X_77832_ _77832_/A _77847_/A sky130_fd_sc_hd__inv_2
Xclkbuf_10_661_0_CLK clkbuf_9_330_0_CLK/X _82888_/CLK sky130_fd_sc_hd__clkbuf_1
X_70167_ _70157_/A _70337_/A sky130_fd_sc_hd__inv_2
X_47992_ _46493_/X _82354_/Q _47991_/Y _57567_/A sky130_fd_sc_hd__o21ai_4
X_59978_ _59974_/Y _59977_/Y _59978_/Y sky130_fd_sc_hd__nand2_4
X_49731_ _86333_/Q _49715_/X _49730_/Y _49731_/Y sky130_fd_sc_hd__o21ai_4
X_46943_ _46942_/Y _52763_/D sky130_fd_sc_hd__buf_2
X_42066_ _40939_/X _41907_/X _88050_/Q _41912_/X _88050_/D sky130_fd_sc_hd__a2bb2o_4
X_58929_ _58904_/X _85765_/Q _58928_/X _58929_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_9_152_0_CLK clkbuf_8_76_0_CLK/X clkbuf_9_152_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_77763_ _77771_/B _81926_/D _77763_/Y sky130_fd_sc_hd__xnor2_4
X_74975_ _74966_/Y _74973_/Y _74974_/Y _74975_/X sky130_fd_sc_hd__o21a_4
X_70098_ _83135_/Q _70102_/A sky130_fd_sc_hd__inv_2
X_79502_ _79502_/A _79502_/B _79503_/B sky130_fd_sc_hd__xor2_4
X_41017_ _40999_/X _41000_/X _41016_/X _88293_/Q _40995_/X _41018_/A
+ sky130_fd_sc_hd__o32ai_4
X_76714_ _76714_/A _76714_/Y sky130_fd_sc_hd__inv_2
X_49662_ _49661_/X _52876_/B _49662_/Y sky130_fd_sc_hd__nand2_4
X_61940_ _61939_/X _61924_/B _61878_/C _61910_/D _61940_/Y sky130_fd_sc_hd__nand4_4
X_73926_ _72894_/X _86226_/Q _45896_/X _73925_/X _73926_/X sky130_fd_sc_hd__a211o_4
X_46874_ _82950_/Q _54417_/D sky130_fd_sc_hd__inv_2
X_77694_ _77694_/A _77695_/A sky130_fd_sc_hd__inv_2
X_48613_ _48613_/A _48661_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_676_0_CLK clkbuf_9_338_0_CLK/X _87144_/CLK sky130_fd_sc_hd__clkbuf_1
X_79433_ _79433_/A _79433_/B _79433_/Y sky130_fd_sc_hd__nand2_4
X_45825_ _45823_/Y _45394_/X _45571_/X _45824_/Y _45825_/X sky130_fd_sc_hd__a211o_4
X_76645_ _76645_/A _76644_/Y _76645_/Y sky130_fd_sc_hd__nand2_4
X_49593_ _49591_/Y _49570_/X _49592_/X _86359_/D sky130_fd_sc_hd__a21oi_4
X_73857_ _73262_/A _73857_/X sky130_fd_sc_hd__buf_2
X_61871_ _61871_/A _61839_/B _61839_/C _63110_/B _61871_/X sky130_fd_sc_hd__and4_4
X_63610_ _63657_/A _63610_/B _63610_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_167_0_CLK clkbuf_8_83_0_CLK/X clkbuf_9_167_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_48544_ _48544_/A _52182_/A sky130_fd_sc_hd__buf_2
X_60822_ _64561_/A _57872_/A _60822_/C _60822_/X sky130_fd_sc_hd__or3_4
X_72808_ _72806_/X _86207_/Q _72746_/X _72807_/X _72808_/X sky130_fd_sc_hd__a211o_4
X_79364_ _79362_/X _79369_/B _79364_/Y sky130_fd_sc_hd__xnor2_4
X_45756_ _57326_/B _45675_/X _45755_/X _45756_/Y sky130_fd_sc_hd__o21ai_4
X_64590_ _44175_/A _64829_/A sky130_fd_sc_hd__buf_2
X_76576_ _76572_/Y _76576_/B _76575_/Y _76576_/X sky130_fd_sc_hd__or3_4
X_42968_ _42968_/A _42968_/Y sky130_fd_sc_hd__inv_2
X_73788_ _73786_/X _84984_/Q _73740_/X _73787_/X _73789_/B sky130_fd_sc_hd__a211o_4
Xclkbuf_9_94_0_CLK clkbuf_9_94_0_CLK/A clkbuf_9_94_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_78315_ _78316_/A _82659_/D _78318_/A sky130_fd_sc_hd__or2_4
X_44707_ _44529_/A _44707_/X sky130_fd_sc_hd__buf_2
X_63541_ _59415_/A _63541_/B _63514_/C _63541_/D _63541_/Y sky130_fd_sc_hd__nand4_4
X_75527_ _75505_/Y _75538_/B _75503_/Y _75528_/B sky130_fd_sc_hd__o21a_4
X_41919_ _42477_/A _41919_/X sky130_fd_sc_hd__buf_2
X_48475_ _74416_/A _50447_/A sky130_fd_sc_hd__buf_2
X_60753_ _60748_/X _60750_/X _60684_/X _60726_/Y _60752_/Y _60753_/Y
+ sky130_fd_sc_hd__a41oi_4
X_72739_ _72739_/A _72739_/X sky130_fd_sc_hd__buf_2
X_79295_ _79282_/X _79293_/X _79294_/X _79295_/Y sky130_fd_sc_hd__a21oi_4
X_45687_ _45679_/X _45683_/Y _45686_/Y _45687_/Y sky130_fd_sc_hd__a21oi_4
X_42899_ _51949_/A _42962_/A sky130_fd_sc_hd__buf_2
X_47426_ _47426_/A _53044_/D sky130_fd_sc_hd__buf_2
X_66260_ _65796_/X _66276_/B _65798_/X _66260_/Y sky130_fd_sc_hd__nand3_4
X_78246_ _78246_/A _78245_/Y _78247_/B sky130_fd_sc_hd__xor2_4
X_44638_ _44679_/A _44638_/X sky130_fd_sc_hd__buf_2
X_75458_ _75458_/A _75458_/X sky130_fd_sc_hd__buf_2
X_63472_ _63448_/A _58506_/A _63458_/X _63496_/D _63472_/X sky130_fd_sc_hd__and4_4
X_60684_ _63416_/A _60732_/C _60804_/C _63699_/D _60684_/X sky130_fd_sc_hd__a211o_4
X_65211_ _65859_/A _65211_/X sky130_fd_sc_hd__buf_2
X_62423_ _62479_/A _61954_/X _62364_/X _62392_/D _62423_/X sky130_fd_sc_hd__and4_4
X_74409_ _83072_/Q _74377_/X _74408_/Y _74409_/Y sky130_fd_sc_hd__o21ai_4
X_47357_ _47380_/A _47349_/B _47370_/C _53003_/D _47357_/X sky130_fd_sc_hd__and4_4
X_66191_ _66179_/X _66189_/Y _66190_/Y _66191_/Y sky130_fd_sc_hd__o21ai_4
X_78177_ _78177_/A _78177_/B _78177_/Y sky130_fd_sc_hd__nor2_4
X_44569_ _44565_/X _44567_/X _40866_/X _87052_/Q _44568_/X _44570_/A
+ sky130_fd_sc_hd__o32ai_4
X_75389_ _75369_/Y _75404_/B _75404_/A _75390_/B sky130_fd_sc_hd__a21boi_4
X_46308_ _46308_/A _46428_/B sky130_fd_sc_hd__buf_2
X_65142_ _65047_/A _65047_/B _65142_/C _65142_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_10_614_0_CLK clkbuf_9_307_0_CLK/X _80854_/CLK sky130_fd_sc_hd__clkbuf_1
X_77128_ _77127_/A _77127_/B _77128_/Y sky130_fd_sc_hd__nand2_4
X_62354_ _62352_/Y _62327_/X _62353_/Y _84416_/D sky130_fd_sc_hd__a21oi_4
X_47288_ _83386_/Q _54130_/B sky130_fd_sc_hd__inv_2
X_61305_ _61305_/A _61301_/X _72583_/C _61305_/Y sky130_fd_sc_hd__nand3_4
X_49027_ _64992_/B _49003_/X _49026_/Y _49027_/Y sky130_fd_sc_hd__o21ai_4
X_46239_ _46239_/A _48882_/A sky130_fd_sc_hd__inv_2
X_65073_ _65069_/Y _65070_/X _65072_/Y _84216_/D sky130_fd_sc_hd__a21o_4
Xclkbuf_9_105_0_CLK clkbuf_8_52_0_CLK/X clkbuf_9_105_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_69950_ _87042_/Q _44225_/B _57800_/A _69949_/X _69950_/X sky130_fd_sc_hd__a211o_4
X_77059_ _77067_/A _77068_/A _77060_/B sky130_fd_sc_hd__xor2_4
X_62285_ _62276_/X _62285_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_32_0_CLK clkbuf_9_33_0_CLK/A clkbuf_9_32_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_64024_ _63749_/A _64118_/B sky130_fd_sc_hd__buf_2
X_68901_ _69014_/A _68994_/A sky130_fd_sc_hd__buf_2
X_61236_ _61198_/X _64203_/B _61237_/D sky130_fd_sc_hd__nand2_4
X_80070_ _80068_/X _80069_/X _80070_/Y sky130_fd_sc_hd__xnor2_4
X_69881_ _81962_/D _69831_/X _69880_/X _83890_/D sky130_fd_sc_hd__a21bo_4
Xclkbuf_10_629_0_CLK clkbuf_9_314_0_CLK/X _81970_/CLK sky130_fd_sc_hd__clkbuf_1
X_68832_ _68059_/A _68832_/X sky130_fd_sc_hd__buf_2
X_61167_ _61097_/X _61103_/X _59980_/X _61167_/Y sky130_fd_sc_hd__a21oi_4
X_60118_ _62244_/D _59950_/B _59977_/B _60118_/X sky130_fd_sc_hd__and3_4
X_49929_ _72220_/B _49906_/X _49928_/Y _49929_/Y sky130_fd_sc_hd__o21ai_4
X_68763_ _68735_/A _68763_/B _68763_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_47_0_CLK clkbuf_9_47_0_CLK/A clkbuf_9_47_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_65975_ _68347_/A _65976_/A sky130_fd_sc_hd__buf_2
X_61098_ _61083_/C _61172_/A sky130_fd_sc_hd__buf_2
X_67714_ _67690_/X _67714_/B _67714_/X sky130_fd_sc_hd__and2_4
X_52940_ _52944_/A _52940_/B _52940_/Y sky130_fd_sc_hd__nand2_4
X_64926_ _64926_/A _64926_/B _64926_/Y sky130_fd_sc_hd__nand2_4
X_60049_ _60049_/A _60049_/Y sky130_fd_sc_hd__inv_2
X_83760_ _83421_/CLK _83760_/D _57655_/A sky130_fd_sc_hd__dfxtp_4
X_80972_ _80931_/CLK _75667_/X _75554_/B sky130_fd_sc_hd__dfxtp_4
X_68694_ _88102_/Q _68636_/X _68691_/X _68693_/Y _68694_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_3_5_0_CLK clkbuf_2_2_2_CLK/X clkbuf_3_5_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_82711_ _82711_/CLK _82711_/D _82667_/D sky130_fd_sc_hd__dfxtp_4
X_67645_ _87462_/Q _67594_/X _67595_/X _67644_/X _67645_/X sky130_fd_sc_hd__a211o_4
X_52871_ _52845_/A _52872_/C sky130_fd_sc_hd__buf_2
X_64857_ _64817_/X _86136_/Q _64776_/X _64856_/X _64857_/X sky130_fd_sc_hd__a211o_4
X_83691_ _85635_/CLK _83691_/D _47204_/A sky130_fd_sc_hd__dfxtp_4
X_54610_ _85410_/Q _54593_/X _54609_/Y _54610_/Y sky130_fd_sc_hd__o21ai_4
X_85430_ _85431_/CLK _54504_/Y _85430_/Q sky130_fd_sc_hd__dfxtp_4
X_51822_ _51822_/A _51823_/A sky130_fd_sc_hd__buf_2
X_63808_ _58232_/X _63858_/B _63858_/C _63793_/D _63809_/D sky130_fd_sc_hd__nand4_4
X_82642_ _82642_/CLK _83994_/Q _78948_/A sky130_fd_sc_hd__dfxtp_4
X_55590_ _55908_/A _55590_/B _55590_/X sky130_fd_sc_hd__and2_4
X_67576_ _87157_/Q _67551_/X _67552_/X _67575_/X _67577_/B sky130_fd_sc_hd__a211o_4
X_64788_ _66002_/A _64789_/A sky130_fd_sc_hd__buf_2
X_69315_ _69315_/A _69315_/X sky130_fd_sc_hd__buf_2
X_54541_ _54486_/A _54546_/A sky130_fd_sc_hd__buf_2
X_66527_ _44147_/A _68386_/A sky130_fd_sc_hd__buf_2
X_85361_ _86289_/CLK _85361_/D _85361_/Q sky130_fd_sc_hd__dfxtp_4
X_51753_ _85952_/Q _51387_/X _51752_/Y _51753_/Y sky130_fd_sc_hd__o21ai_4
X_63739_ _84905_/Q _60921_/X _60895_/X _63739_/Y sky130_fd_sc_hd__o21ai_4
X_82573_ _82604_/CLK _82605_/Q _78154_/A sky130_fd_sc_hd__dfxtp_4
X_87100_ _88272_/CLK _87100_/D _87100_/Q sky130_fd_sc_hd__dfxtp_4
X_84312_ _84314_/CLK _63580_/Y _80442_/B sky130_fd_sc_hd__dfxtp_4
X_50704_ _50695_/A _53919_/B _50704_/Y sky130_fd_sc_hd__nand2_4
X_57260_ _57243_/X _56634_/X _45585_/A _57245_/X _57260_/X sky130_fd_sc_hd__a2bb2o_4
X_81524_ _81532_/CLK _81568_/Q _76054_/A sky130_fd_sc_hd__dfxtp_4
X_69246_ _69191_/A _87787_/Q _69246_/X sky130_fd_sc_hd__and2_4
X_88080_ _87824_/CLK _88080_/D _88080_/Q sky130_fd_sc_hd__dfxtp_4
X_54472_ _54470_/Y _54448_/X _54471_/X _85436_/D sky130_fd_sc_hd__a21oi_4
X_66458_ _66173_/A _66517_/B _66173_/C _66458_/Y sky130_fd_sc_hd__nand3_4
X_85292_ _80671_/CLK _56125_/Y _56124_/C sky130_fd_sc_hd__dfxtp_4
X_51684_ _51695_/A _51684_/B _51684_/C _53207_/D _51684_/X sky130_fd_sc_hd__and4_4
X_56211_ _56200_/X _56205_/X _56211_/C _56211_/Y sky130_fd_sc_hd__nand3_4
X_87031_ _87333_/CLK _87031_/D _87031_/Q sky130_fd_sc_hd__dfxtp_4
X_53423_ _85636_/Q _53404_/X _53422_/Y _53423_/Y sky130_fd_sc_hd__o21ai_4
X_65409_ _65252_/X _83282_/Q _65407_/X _65408_/X _65409_/X sky130_fd_sc_hd__a211o_4
X_84243_ _84458_/CLK _64472_/X _79649_/B sky130_fd_sc_hd__dfxtp_4
X_50635_ _50633_/Y _50619_/X _50634_/Y _86163_/D sky130_fd_sc_hd__a21boi_4
X_57191_ _57331_/A _57331_/C _57121_/X _57195_/A sky130_fd_sc_hd__a21o_4
X_81455_ _81333_/CLK _76771_/B _81423_/D sky130_fd_sc_hd__dfxtp_4
X_69177_ _88048_/Q _68975_/X _68976_/X _69176_/X _69177_/X sky130_fd_sc_hd__a211o_4
X_66389_ _66389_/A _66389_/B _66389_/C _66389_/Y sky130_fd_sc_hd__nor3_4
X_56142_ _56142_/A _56142_/X sky130_fd_sc_hd__buf_2
X_80406_ _80406_/A _80406_/B _80406_/X sky130_fd_sc_hd__and2_4
X_68128_ _68089_/A _68128_/X sky130_fd_sc_hd__buf_2
X_53354_ _85649_/Q _53351_/X _53353_/Y _53354_/Y sky130_fd_sc_hd__o21ai_4
Xpsn_inst_psn_buff_5 _71215_/Y _71216_/A sky130_fd_sc_hd__buf_8
X_84174_ _85346_/CLK _84174_/D _84174_/Q sky130_fd_sc_hd__dfxtp_4
X_50566_ _86176_/Q _50563_/X _50565_/Y _50566_/Y sky130_fd_sc_hd__o21ai_4
X_81386_ _81352_/CLK _83922_/Q _76864_/B sky130_fd_sc_hd__dfxtp_4
X_52305_ _52295_/A _48969_/A _52305_/X sky130_fd_sc_hd__and2_4
X_83125_ _83145_/CLK _74050_/Y _70110_/A sky130_fd_sc_hd__dfxtp_4
X_56073_ _56073_/A _55864_/X _56073_/Y sky130_fd_sc_hd__xnor2_4
X_80337_ _80334_/Y _80336_/Y _80337_/Y sky130_fd_sc_hd__nand2_4
X_68059_ _68059_/A _68059_/X sky130_fd_sc_hd__buf_2
X_53285_ _53281_/Y _53272_/X _53284_/X _53285_/Y sky130_fd_sc_hd__a21oi_4
X_50497_ _52204_/A _50526_/B _50497_/C _50497_/X sky130_fd_sc_hd__and3_4
X_55024_ _54253_/A _55024_/X sky130_fd_sc_hd__buf_2
X_59901_ _59901_/A _59705_/X _59901_/C _59901_/Y sky130_fd_sc_hd__nand3_4
X_52236_ _85862_/Q _52214_/X _52235_/Y _52236_/Y sky130_fd_sc_hd__o21ai_4
X_71070_ _71070_/A _71070_/X sky130_fd_sc_hd__buf_2
X_83056_ _85571_/CLK _83056_/D _83056_/Q sky130_fd_sc_hd__dfxtp_4
X_87933_ _87421_/CLK _42300_/Y _87933_/Q sky130_fd_sc_hd__dfxtp_4
X_80268_ _80267_/Y _80268_/B _80268_/Y sky130_fd_sc_hd__nand2_4
X_70021_ _70021_/A _70020_/X _70021_/C _70021_/Y sky130_fd_sc_hd__nand3_4
X_82007_ _82008_/CLK _82007_/D _77157_/A sky130_fd_sc_hd__dfxtp_4
X_59832_ _59831_/X _59834_/A sky130_fd_sc_hd__buf_2
X_52167_ _52164_/Y _52145_/X _52166_/X _85876_/D sky130_fd_sc_hd__a21oi_4
X_87864_ _87865_/CLK _87864_/D _87864_/Q sky130_fd_sc_hd__dfxtp_4
X_80199_ _80173_/Y _80176_/Y _80184_/Y _80187_/Y _80199_/X sky130_fd_sc_hd__o22a_4
X_51118_ _86070_/Q _51101_/X _51117_/Y _51118_/Y sky130_fd_sc_hd__o21ai_4
X_86815_ _81182_/CLK _86815_/D _67133_/B sky130_fd_sc_hd__dfxtp_4
X_59763_ _59763_/A _59716_/A _59716_/B _59763_/X sky130_fd_sc_hd__and3_4
X_52098_ _53620_/A _52098_/B _52097_/X _52098_/X sky130_fd_sc_hd__and3_4
X_56975_ _57193_/D _56922_/X _83329_/Q _56975_/Y sky130_fd_sc_hd__nor3_4
X_87795_ _88084_/CLK _42635_/X _87795_/Q sky130_fd_sc_hd__dfxtp_4
X_58714_ _58846_/A _58714_/X sky130_fd_sc_hd__buf_2
X_51049_ _51058_/A _46899_/X _51049_/Y sky130_fd_sc_hd__nand2_4
X_55926_ _55926_/A _55926_/B _55926_/X sky130_fd_sc_hd__and2_4
X_43940_ _43605_/A _45964_/A sky130_fd_sc_hd__buf_2
X_74760_ _74760_/A _74720_/C _74804_/D _74780_/D _74760_/Y sky130_fd_sc_hd__nand4_4
X_86746_ _85818_/CLK _86746_/D _86746_/Q sky130_fd_sc_hd__dfxtp_4
X_71972_ _71972_/A _71972_/B _71972_/Y sky130_fd_sc_hd__nand2_4
X_83958_ _80821_/CLK _68857_/X _83958_/Q sky130_fd_sc_hd__dfxtp_4
X_59694_ _62185_/B _62183_/A sky130_fd_sc_hd__buf_2
X_73711_ _73711_/A _73711_/B _73711_/X sky130_fd_sc_hd__and2_4
X_58645_ _58112_/X _86107_/Q _58644_/X _58645_/Y sky130_fd_sc_hd__o21ai_4
X_70923_ _70871_/A _70914_/B _70914_/C _70919_/D _70923_/Y sky130_fd_sc_hd__nand4_4
X_82909_ _87416_/CLK _78278_/B _82909_/Q sky130_fd_sc_hd__dfxtp_4
X_43871_ _41250_/X _43868_/X _68980_/B _43870_/X _43871_/X sky130_fd_sc_hd__a2bb2o_4
X_55857_ _44079_/X _55857_/B _55857_/X sky130_fd_sc_hd__and2_4
X_74691_ _74691_/A _74691_/B _74691_/Y sky130_fd_sc_hd__nand2_4
X_86677_ _86359_/CLK _86677_/D _86677_/Q sky130_fd_sc_hd__dfxtp_4
X_83889_ _82339_/CLK _83889_/D _83889_/Q sky130_fd_sc_hd__dfxtp_4
X_45610_ _45603_/X _45606_/X _45609_/Y _86866_/D sky130_fd_sc_hd__a21oi_4
X_76430_ _76430_/A _76430_/B _76430_/C _76430_/X sky130_fd_sc_hd__or3_4
X_42822_ _42822_/A _42822_/X sky130_fd_sc_hd__buf_2
X_54808_ _54400_/A _54889_/A sky130_fd_sc_hd__buf_2
X_73642_ _72829_/X _84990_/Q _73614_/X _73641_/X _73642_/X sky130_fd_sc_hd__a211o_4
X_85628_ _86237_/CLK _53485_/Y _85628_/Q sky130_fd_sc_hd__dfxtp_4
X_46590_ _46578_/X _49190_/A _46589_/X _46591_/A sky130_fd_sc_hd__o21ai_4
X_58576_ _58576_/A _58576_/B _58576_/Y sky130_fd_sc_hd__nor2_4
X_70854_ _70854_/A _70698_/A _70855_/A sky130_fd_sc_hd__nor2_4
X_55788_ _55761_/A _85291_/Q _55788_/X sky130_fd_sc_hd__and2_4
X_57527_ _46542_/X _57527_/X sky130_fd_sc_hd__buf_2
X_45541_ _83000_/Q _45604_/B _45541_/Y sky130_fd_sc_hd__nor2_4
X_76361_ _76324_/Y _76356_/Y _76360_/Y _76361_/Y sky130_fd_sc_hd__a21oi_4
X_88347_ _87859_/CLK _40726_/Y _88347_/Q sky130_fd_sc_hd__dfxtp_4
X_42753_ _41250_/X _42745_/X _68977_/B _42746_/X _42753_/X sky130_fd_sc_hd__a2bb2o_4
X_54739_ _54748_/A _54755_/B _54748_/C _54739_/D _54739_/X sky130_fd_sc_hd__and4_4
X_73573_ _74117_/A _73572_/Y _73573_/Y sky130_fd_sc_hd__nor2_4
X_85559_ _83305_/CLK _53835_/Y _85559_/Q sky130_fd_sc_hd__dfxtp_4
X_70785_ _52859_/B _70761_/X _70784_/Y _70785_/Y sky130_fd_sc_hd__o21ai_4
X_78100_ _78100_/A _78099_/Y _78101_/B sky130_fd_sc_hd__xor2_4
X_75312_ _80690_/Q _80990_/Q _75312_/Y sky130_fd_sc_hd__nand2_4
X_41704_ _41603_/X _82899_/Q _41703_/X _41704_/X sky130_fd_sc_hd__o21a_4
X_48260_ _86546_/Q _48188_/X _48259_/Y _48260_/Y sky130_fd_sc_hd__o21ai_4
X_72524_ _72602_/A _72525_/A sky130_fd_sc_hd__buf_2
X_79080_ _79080_/A _82623_/D sky130_fd_sc_hd__inv_2
X_45472_ _85116_/Q _45456_/X _45472_/Y sky130_fd_sc_hd__nor2_4
X_57458_ _55248_/B _57463_/B _57458_/X sky130_fd_sc_hd__or2_4
X_76292_ _76291_/X _76296_/A sky130_fd_sc_hd__inv_2
X_42684_ _41070_/X _42679_/X _69466_/B _42681_/X _42684_/X sky130_fd_sc_hd__a2bb2o_4
X_88278_ _82301_/CLK _88278_/D _69536_/B sky130_fd_sc_hd__dfxtp_4
X_47211_ _47207_/Y _47177_/X _47210_/X _47211_/Y sky130_fd_sc_hd__a21oi_4
X_78031_ _78031_/A _78031_/B _78033_/A sky130_fd_sc_hd__nand2_4
X_44423_ _44422_/Y _87115_/D sky130_fd_sc_hd__inv_2
X_56409_ _56439_/A _56409_/X sky130_fd_sc_hd__buf_2
X_75243_ _75243_/A _75243_/Y sky130_fd_sc_hd__inv_2
X_41635_ _41577_/X _82912_/Q _41634_/X _41635_/Y sky130_fd_sc_hd__o21ai_4
X_87229_ _87235_/CLK _43861_/X _68920_/B sky130_fd_sc_hd__dfxtp_4
X_48191_ _86558_/Q _48188_/X _48190_/Y _48191_/Y sky130_fd_sc_hd__o21ai_4
X_72455_ _83252_/Q _79549_/B sky130_fd_sc_hd__inv_2
X_57389_ _57384_/X _56584_/X _85021_/Q _57385_/X _57389_/X sky130_fd_sc_hd__a2bb2o_4
X_47142_ _54571_/D _52879_/D sky130_fd_sc_hd__buf_2
X_59128_ _84767_/Q _59043_/X _59120_/X _59127_/X _59128_/Y sky130_fd_sc_hd__a2bb2oi_4
X_71406_ _70679_/A _71404_/B _71411_/C _71406_/Y sky130_fd_sc_hd__nor3_4
X_44354_ _44350_/X _44351_/X _41710_/X _87152_/Q _44353_/X _44355_/A
+ sky130_fd_sc_hd__o32ai_4
X_75174_ _75169_/Y _75175_/A sky130_fd_sc_hd__inv_2
X_41566_ _41540_/X _41541_/X _41565_/X _67052_/B _41537_/X _41567_/A
+ sky130_fd_sc_hd__o32ai_4
X_72386_ _72255_/A _72386_/X sky130_fd_sc_hd__buf_2
X_43305_ _43305_/A _43305_/X sky130_fd_sc_hd__buf_2
X_74125_ _74122_/X _74124_/X _72737_/A _74125_/X sky130_fd_sc_hd__a21o_4
X_40517_ _40516_/Y _88379_/D sky130_fd_sc_hd__inv_2
X_47073_ _82385_/Q _47074_/A sky130_fd_sc_hd__inv_2
X_59059_ _59048_/X _85660_/Q _59010_/X _59059_/X sky130_fd_sc_hd__o21a_4
X_71337_ _71337_/A _71338_/A sky130_fd_sc_hd__buf_2
X_44285_ _45950_/A _44268_/A _44210_/X _44285_/Y sky130_fd_sc_hd__nor3_4
X_79982_ _79982_/A _79981_/Y _79982_/X sky130_fd_sc_hd__xor2_4
X_41497_ _41344_/X _40402_/B _41496_/X _41497_/X sky130_fd_sc_hd__o21a_4
X_46024_ _40537_/Y _46022_/X _86809_/Q _46023_/X _86809_/D sky130_fd_sc_hd__a2bb2o_4
X_43236_ _43236_/A _87525_/D sky130_fd_sc_hd__inv_2
X_62070_ _62037_/X _62021_/B _58495_/A _62020_/X _62070_/X sky130_fd_sc_hd__and4_4
X_74056_ _68892_/B _72899_/X _73898_/X _74056_/X sky130_fd_sc_hd__o21a_4
X_78933_ _78923_/B _82511_/D sky130_fd_sc_hd__inv_2
X_40448_ _40437_/X _40443_/X _40446_/X _88390_/Q _40447_/X _40448_/Y
+ sky130_fd_sc_hd__o32ai_4
X_71268_ _71268_/A _71276_/B sky130_fd_sc_hd__buf_2
X_73007_ _73007_/A _73007_/X sky130_fd_sc_hd__buf_2
X_61021_ _61018_/Y _60952_/X _61019_/X _76986_/A _61020_/X _84538_/D
+ sky130_fd_sc_hd__o32a_4
X_70219_ _70229_/A _70229_/B _70219_/C _70229_/D _70219_/X sky130_fd_sc_hd__and4_4
X_43167_ _43167_/A _43167_/X sky130_fd_sc_hd__buf_2
X_78864_ _78877_/B _78877_/A _78868_/A sky130_fd_sc_hd__xnor2_4
X_40379_ _47825_/A _40380_/A sky130_fd_sc_hd__buf_2
X_71199_ _71197_/A _71055_/B _71197_/C _71199_/Y sky130_fd_sc_hd__nand3_4
X_42118_ _42099_/X _42116_/X _41076_/X _88026_/Q _42117_/X _42118_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77815_ _77828_/A _77814_/Y _77835_/A sky130_fd_sc_hd__xor2_4
X_47975_ _47946_/A _47975_/B _47975_/X sky130_fd_sc_hd__and2_4
X_43098_ _43098_/A _43098_/Y sky130_fd_sc_hd__inv_2
X_78795_ _78795_/A _78795_/B _78797_/A sky130_fd_sc_hd__nand2_4
X_49714_ _49711_/Y _49706_/X _49713_/X _49714_/Y sky130_fd_sc_hd__a21oi_4
X_46926_ _46915_/X _46896_/B _46926_/C _52750_/D _46926_/X sky130_fd_sc_hd__and4_4
X_42049_ _41993_/A _42049_/X sky130_fd_sc_hd__buf_2
X_65760_ _65188_/X _65653_/B _65191_/X _65772_/A sky130_fd_sc_hd__nand3_4
X_77746_ _81972_/Q _77747_/B sky130_fd_sc_hd__inv_2
X_74958_ _74958_/A _74958_/B _74961_/B _74959_/B sky130_fd_sc_hd__and3_4
X_62972_ _58207_/A _62924_/C _62827_/X _62644_/X _62971_/X _62972_/Y
+ sky130_fd_sc_hd__a41oi_4
X_64711_ _64704_/X _86749_/Q _64707_/X _64710_/X _64711_/X sky130_fd_sc_hd__a211o_4
X_49645_ _59244_/B _49632_/X _49644_/Y _49645_/Y sky130_fd_sc_hd__o21ai_4
X_61923_ _61712_/X _61924_/B sky130_fd_sc_hd__buf_2
X_73909_ _73907_/X _84979_/Q _73859_/X _73908_/X _73910_/B sky130_fd_sc_hd__a211o_4
X_46857_ _46830_/A _46845_/X _46868_/C _52716_/D _46857_/X sky130_fd_sc_hd__and4_4
X_65691_ _65688_/X _65690_/X _65642_/X _65694_/A sky130_fd_sc_hd__a21o_4
X_77677_ _77673_/Y _77675_/Y _77676_/A _77677_/Y sky130_fd_sc_hd__o21ai_4
X_74889_ _74889_/A _74890_/B sky130_fd_sc_hd__buf_2
X_67430_ _87407_/Q _67358_/X _67360_/X _67429_/X _67430_/X sky130_fd_sc_hd__a211o_4
X_79416_ _79416_/A _79416_/B _79439_/A sky130_fd_sc_hd__xor2_4
X_45808_ _45808_/A _45808_/Y sky130_fd_sc_hd__inv_2
X_64642_ _64642_/A _64642_/X sky130_fd_sc_hd__buf_2
X_76628_ _76628_/A _76628_/Y sky130_fd_sc_hd__inv_2
X_61854_ _57652_/X _61824_/X _61838_/X _61790_/X _61853_/X _61854_/X
+ sky130_fd_sc_hd__a41o_4
X_49576_ _49548_/A _49577_/C sky130_fd_sc_hd__buf_2
X_46788_ _46806_/A _50981_/B _46788_/Y sky130_fd_sc_hd__nand2_4
X_60805_ _60804_/Y _60805_/Y sky130_fd_sc_hd__inv_2
X_48527_ _48515_/A _48788_/B _48527_/Y sky130_fd_sc_hd__nand2_4
X_79347_ _79333_/Y _79339_/B _79346_/X _79347_/Y sky130_fd_sc_hd__o21ai_4
X_67361_ _67308_/A _67361_/B _67361_/X sky130_fd_sc_hd__and2_4
X_45739_ _45193_/A _45740_/B sky130_fd_sc_hd__buf_2
X_64573_ _44149_/X _85537_/Q _64571_/X _64572_/X _64573_/X sky130_fd_sc_hd__a211o_4
X_76559_ _76559_/A _76559_/Y sky130_fd_sc_hd__inv_2
X_61785_ _61783_/Y _61699_/X _61784_/Y _61785_/Y sky130_fd_sc_hd__a21oi_4
X_69100_ _69236_/A _69100_/B _69100_/X sky130_fd_sc_hd__and2_4
X_66312_ _66309_/X _66311_/X _66240_/X _66312_/X sky130_fd_sc_hd__a21o_4
X_63524_ _63512_/A _63524_/B _63476_/C _63524_/X sky130_fd_sc_hd__and3_4
X_48458_ _48934_/A _48651_/A sky130_fd_sc_hd__buf_2
X_60736_ _63400_/C _60736_/X sky130_fd_sc_hd__buf_2
X_67292_ _67292_/A _67291_/X _67292_/Y sky130_fd_sc_hd__nand2_4
X_79278_ _84795_/Q _84115_/Q _79278_/X sky130_fd_sc_hd__xor2_4
X_69031_ _69134_/A _69031_/B _69031_/X sky130_fd_sc_hd__and2_4
X_47409_ _47405_/Y _47364_/X _47408_/X _47409_/Y sky130_fd_sc_hd__a21oi_4
X_66243_ _66225_/X _84970_/Q _66186_/X _66242_/X _66244_/B sky130_fd_sc_hd__a211o_4
X_78229_ _78234_/A _78225_/A _78228_/Y _78229_/Y sky130_fd_sc_hd__a21boi_4
X_63455_ _63516_/A _63455_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_553_0_CLK clkbuf_9_276_0_CLK/X _82896_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_44_0_CLK clkbuf_6_45_0_CLK/A clkbuf_7_89_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_48389_ _48382_/Y _48383_/X _48388_/X _48389_/Y sky130_fd_sc_hd__a21oi_4
X_60667_ _60667_/A _60667_/Y sky130_fd_sc_hd__inv_2
X_50420_ _86204_/Q _50387_/X _50419_/Y _50420_/Y sky130_fd_sc_hd__o21ai_4
X_81240_ _85334_/CLK _81048_/Q _81240_/Q sky130_fd_sc_hd__dfxtp_4
X_62406_ _62406_/A _62401_/Y _62406_/C _62405_/Y _62406_/Y sky130_fd_sc_hd__nand4_4
X_66174_ _66068_/X _65710_/Y _66173_/Y _66174_/Y sky130_fd_sc_hd__o21ai_4
X_63386_ _63374_/A _61762_/X _63386_/X sky130_fd_sc_hd__and2_4
X_60598_ _60533_/Y _60566_/A _60598_/Y sky130_fd_sc_hd__nand2_4
X_65125_ _65099_/X _86733_/Q _65028_/X _65124_/X _65125_/X sky130_fd_sc_hd__a211o_4
X_50351_ _50227_/A _50351_/X sky130_fd_sc_hd__buf_2
X_62337_ _62337_/A _61861_/X _62237_/X _62280_/D _62337_/X sky130_fd_sc_hd__and4_4
X_81171_ _81179_/CLK _74969_/B _81171_/Q sky130_fd_sc_hd__dfxtp_4
X_80122_ _57912_/Y _65634_/C _80121_/Y _80122_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_10_568_0_CLK clkbuf_9_284_0_CLK/X _87416_/CLK sky130_fd_sc_hd__clkbuf_1
Xpsn_inst_psn_buff_12 _44134_/D _55686_/C sky130_fd_sc_hd__buf_2
X_53070_ _53074_/A _53069_/X _53074_/C _53070_/D _53070_/X sky130_fd_sc_hd__and4_4
X_65056_ _65053_/X _65056_/B _65055_/X _65056_/Y sky130_fd_sc_hd__nand3_4
X_69933_ _73465_/A _69837_/X _68741_/X _69932_/Y _69933_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_6_59_0_CLK clkbuf_6_59_0_CLK/A clkbuf_6_59_0_CLK/X sky130_fd_sc_hd__clkbuf_1
Xpsn_inst_psn_buff_23 _53441_/A _53447_/A sky130_fd_sc_hd__buf_2
X_50282_ _50219_/X _50282_/X sky130_fd_sc_hd__buf_2
X_62268_ _62264_/Y _62253_/X _62267_/Y _84422_/D sky130_fd_sc_hd__a21oi_4
X_52021_ _52021_/A _52462_/A sky130_fd_sc_hd__buf_2
X_64007_ _60034_/X _64074_/A sky130_fd_sc_hd__buf_2
X_61219_ _61218_/Y _61125_/A _84505_/Q _59803_/X _84505_/D sky130_fd_sc_hd__a2bb2o_4
X_84930_ _84930_/CLK _84930_/D _84930_/Q sky130_fd_sc_hd__dfxtp_4
X_80053_ _80025_/Y _80043_/B _80042_/A _80041_/Y _80053_/X sky130_fd_sc_hd__o22a_4
X_69864_ _69861_/X _69863_/X _66579_/X _69864_/X sky130_fd_sc_hd__a21o_4
X_62199_ _62198_/Y _62572_/A sky130_fd_sc_hd__buf_2
X_68815_ _68770_/X _68815_/B _68815_/X sky130_fd_sc_hd__and2_4
X_84861_ _84250_/CLK _84861_/D _84861_/Q sky130_fd_sc_hd__dfxtp_4
X_69795_ _69792_/X _69794_/X _69768_/X _69795_/X sky130_fd_sc_hd__a21o_4
X_86600_ _86600_/CLK _86600_/D _86600_/Q sky130_fd_sc_hd__dfxtp_4
X_83812_ _83842_/CLK _83812_/D _83812_/Q sky130_fd_sc_hd__dfxtp_4
X_56760_ _56759_/X _56788_/A sky130_fd_sc_hd__buf_2
X_68746_ _68746_/A _68746_/B _68746_/Y sky130_fd_sc_hd__nor2_4
X_87580_ _87542_/CLK _87580_/D _87580_/Q sky130_fd_sc_hd__dfxtp_4
X_53972_ _85531_/Q _53955_/X _53971_/Y _53972_/Y sky130_fd_sc_hd__o21ai_4
X_65958_ _72123_/A _86237_/Q _45922_/X _65957_/X _65958_/X sky130_fd_sc_hd__a211o_4
X_84792_ _86697_/CLK _58895_/Y _84792_/Q sky130_fd_sc_hd__dfxtp_4
X_55711_ _55711_/A _55711_/X sky130_fd_sc_hd__buf_2
X_86531_ _86490_/CLK _86531_/D _86531_/Q sky130_fd_sc_hd__dfxtp_4
X_52923_ _52919_/Y _52920_/X _52922_/X _52923_/Y sky130_fd_sc_hd__a21oi_4
X_64909_ _64877_/X _86454_/Q _64909_/X sky130_fd_sc_hd__and2_4
X_83743_ _86322_/CLK _83743_/D _47313_/A sky130_fd_sc_hd__dfxtp_4
X_56691_ _56691_/A _72765_/A sky130_fd_sc_hd__buf_2
X_80955_ _80740_/CLK _80955_/D _80955_/Q sky130_fd_sc_hd__dfxtp_4
X_68677_ _86995_/Q _68394_/X _68421_/X _68676_/X _68677_/X sky130_fd_sc_hd__a211o_4
X_65889_ _65886_/Y _65830_/X _65888_/Y _84171_/D sky130_fd_sc_hd__a21o_4
X_58430_ _58151_/A _83362_/Q _58430_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_506_0_CLK clkbuf_9_253_0_CLK/X _84807_/CLK sky130_fd_sc_hd__clkbuf_1
X_55642_ _83009_/Q _55619_/A _44101_/A _55641_/Y _55642_/X sky130_fd_sc_hd__a211o_4
X_67628_ _67987_/A _67628_/X sky130_fd_sc_hd__buf_2
X_86462_ _83623_/CLK _48919_/Y _64684_/B sky130_fd_sc_hd__dfxtp_4
X_52854_ _52851_/Y _52839_/X _52853_/X _52854_/Y sky130_fd_sc_hd__a21oi_4
X_83674_ _83673_/CLK _70881_/Y _83674_/Q sky130_fd_sc_hd__dfxtp_4
X_80886_ _80740_/CLK _75760_/B _80854_/D sky130_fd_sc_hd__dfxtp_4
X_88201_ _88201_/CLK _41512_/X _88201_/Q sky130_fd_sc_hd__dfxtp_4
X_85413_ _83690_/CLK _85413_/D _85413_/Q sky130_fd_sc_hd__dfxtp_4
X_51805_ _51805_/A _51794_/B _51794_/C _46716_/X _51805_/X sky130_fd_sc_hd__and4_4
X_58361_ _58328_/X _83765_/Q _58360_/Y _84869_/D sky130_fd_sc_hd__o21a_4
X_82625_ _82743_/CLK _82625_/D _82625_/Q sky130_fd_sc_hd__dfxtp_4
X_55573_ _55572_/X _45470_/Y _55573_/Y sky130_fd_sc_hd__nor2_4
X_67559_ _67582_/A _67559_/B _67559_/X sky130_fd_sc_hd__and2_4
X_86393_ _86393_/CLK _86393_/D _86393_/Q sky130_fd_sc_hd__dfxtp_4
X_52785_ _52784_/X _52775_/B _52775_/C _52785_/D _52785_/X sky130_fd_sc_hd__and4_4
X_57312_ _57311_/X _57303_/Y _56704_/X _57312_/Y sky130_fd_sc_hd__a21oi_4
X_88132_ _88394_/CLK _41831_/Y _88132_/Q sky130_fd_sc_hd__dfxtp_4
X_54524_ _54518_/A _53345_/B _54524_/Y sky130_fd_sc_hd__nand2_4
X_85344_ _83711_/CLK _54965_/Y _85344_/Q sky130_fd_sc_hd__dfxtp_4
X_51736_ _51733_/Y _51719_/X _51735_/X _85955_/D sky130_fd_sc_hd__a21oi_4
X_70570_ DATA_TO_HASH[0] _70570_/Y sky130_fd_sc_hd__inv_2
X_58292_ _63672_/B _58248_/B _58292_/Y sky130_fd_sc_hd__nor2_4
X_82556_ _82557_/CLK _82556_/D _82556_/Q sky130_fd_sc_hd__dfxtp_4
X_69229_ _83939_/Q _69161_/X _69228_/X _69229_/X sky130_fd_sc_hd__a21bo_4
X_57243_ _44287_/X _57243_/X sky130_fd_sc_hd__buf_2
X_81507_ _81507_/CLK _76158_/B _75929_/A sky130_fd_sc_hd__dfxtp_4
X_88063_ _87814_/CLK _42034_/Y _73273_/A sky130_fd_sc_hd__dfxtp_4
X_54455_ _54453_/X _54440_/B _54471_/C _46942_/Y _54455_/X sky130_fd_sc_hd__and4_4
X_85275_ _85277_/CLK _85275_/D _56208_/C sky130_fd_sc_hd__dfxtp_4
X_51667_ _51639_/A _51667_/X sky130_fd_sc_hd__buf_2
X_82487_ _82580_/CLK _82487_/D _78177_/B sky130_fd_sc_hd__dfxtp_4
X_87014_ _88288_/CLK _44655_/Y _87014_/Q sky130_fd_sc_hd__dfxtp_4
X_41420_ _41416_/X _41418_/X _67909_/B _41419_/X _88219_/D sky130_fd_sc_hd__a2bb2o_4
X_53406_ _53405_/X _47165_/Y _53406_/Y sky130_fd_sc_hd__nand2_4
X_72240_ _72155_/A _72240_/X sky130_fd_sc_hd__buf_2
X_84226_ _85315_/CLK _84226_/D _84226_/Q sky130_fd_sc_hd__dfxtp_4
X_50618_ _86166_/Q _50594_/X _50617_/Y _50618_/Y sky130_fd_sc_hd__o21ai_4
X_57174_ _57172_/Y _57173_/Y _57121_/X _57175_/B sky130_fd_sc_hd__o21ai_4
X_81438_ _81532_/CLK _81470_/Q _76133_/B sky130_fd_sc_hd__dfxtp_4
X_54386_ _54395_/A _54395_/B _54395_/C _46820_/Y _54386_/X sky130_fd_sc_hd__and4_4
X_51598_ _51580_/A _51603_/B _51603_/C _53125_/D _51598_/X sky130_fd_sc_hd__and4_4
X_56125_ _56112_/X _56121_/X _56124_/Y _56125_/Y sky130_fd_sc_hd__o21ai_4
X_41351_ _41324_/X _82901_/Q _41350_/X _41351_/Y sky130_fd_sc_hd__o21ai_4
X_53337_ _85652_/Q _53324_/X _53336_/Y _53337_/Y sky130_fd_sc_hd__o21ai_4
X_72171_ _72168_/Y _72170_/Y _59297_/X _72171_/X sky130_fd_sc_hd__a21o_4
X_84157_ _84161_/CLK _66093_/X _84157_/Q sky130_fd_sc_hd__dfxtp_4
X_50549_ _50541_/A _48695_/B _50549_/Y sky130_fd_sc_hd__nand2_4
X_81369_ _81428_/CLK _76867_/Y _76500_/A sky130_fd_sc_hd__dfxtp_4
X_71122_ _49135_/X _71117_/X _71121_/Y _83600_/D sky130_fd_sc_hd__o21ai_4
X_83108_ _82998_/CLK _74298_/X _70280_/A sky130_fd_sc_hd__dfxtp_4
X_44070_ _87176_/Q _44070_/B _43972_/B _44071_/A sky130_fd_sc_hd__nor3_4
X_56056_ _56052_/A _56052_/B _55915_/B _56056_/Y sky130_fd_sc_hd__nand3_4
X_41282_ _41281_/Y _41282_/X sky130_fd_sc_hd__buf_2
X_53268_ _51900_/A _53268_/X sky130_fd_sc_hd__buf_2
X_84088_ _83918_/CLK _66993_/X _84088_/Q sky130_fd_sc_hd__dfxtp_4
X_43021_ _43024_/A _43021_/X sky130_fd_sc_hd__buf_2
X_55007_ _55011_/A _47610_/A _55007_/Y sky130_fd_sc_hd__nand2_4
X_52219_ _52217_/Y _52203_/X _52218_/X _85866_/D sky130_fd_sc_hd__a21oi_4
X_71053_ _48889_/B _71047_/X _71052_/Y _71053_/Y sky130_fd_sc_hd__o21ai_4
X_75930_ _81700_/D _75930_/B _75933_/A sky130_fd_sc_hd__nor2_4
X_83039_ _85311_/CLK _74546_/Y _74545_/C sky130_fd_sc_hd__dfxtp_4
X_87916_ _88171_/CLK _42335_/Y _87916_/Q sky130_fd_sc_hd__dfxtp_4
X_53199_ _53199_/A _53219_/A sky130_fd_sc_hd__buf_2
X_70004_ _82555_/D _69988_/X _70003_/X _70004_/X sky130_fd_sc_hd__a21bo_4
X_59815_ _59805_/Y _59840_/A _59812_/Y _80442_/A _59814_/X _84696_/D
+ sky130_fd_sc_hd__o32a_4
X_75861_ _75860_/A _75860_/B _75864_/A sky130_fd_sc_hd__or2_4
X_87847_ _87850_/CLK _87847_/D _68668_/A sky130_fd_sc_hd__dfxtp_4
X_77600_ _77601_/A _82107_/D _77600_/Y sky130_fd_sc_hd__nor2_4
X_74812_ _46168_/Y _46169_/Y _46171_/Y _80665_/D sky130_fd_sc_hd__a21oi_4
X_47760_ _47714_/A _47760_/X sky130_fd_sc_hd__buf_2
X_59746_ _59689_/A _59631_/B _59746_/Y sky130_fd_sc_hd__nand2_4
X_78580_ _78561_/A _78577_/X _78579_/Y _78581_/B sky130_fd_sc_hd__a21oi_4
X_44972_ _44972_/A _44972_/X sky130_fd_sc_hd__buf_2
X_56958_ _56613_/X _56952_/X _56957_/Y _85113_/D sky130_fd_sc_hd__a21oi_4
X_75792_ _75788_/Y _75775_/Y _75791_/Y _75793_/B sky130_fd_sc_hd__o21ai_4
X_87778_ _87533_/CLK _87778_/D _87778_/Q sky130_fd_sc_hd__dfxtp_4
X_46711_ _52632_/B _51800_/B sky130_fd_sc_hd__buf_2
X_77531_ _77519_/A _77529_/Y _77530_/Y _77540_/A sky130_fd_sc_hd__o21a_4
X_43923_ _43922_/Y _87197_/D sky130_fd_sc_hd__inv_2
X_55909_ _56216_/C _44106_/C _44051_/A _55908_/X _55909_/X sky130_fd_sc_hd__a211o_4
X_74743_ _70730_/X _74804_/C sky130_fd_sc_hd__buf_2
X_86729_ _86121_/CLK _46532_/Y _86729_/Q sky130_fd_sc_hd__dfxtp_4
X_47691_ _47691_/A _53191_/D sky130_fd_sc_hd__buf_2
X_71955_ _71867_/A _70538_/X _71404_/B _71955_/Y sky130_fd_sc_hd__nor3_4
X_59677_ _59655_/X _59687_/B _59651_/C _59763_/A _59676_/Y _59677_/Y
+ sky130_fd_sc_hd__a41oi_4
X_56889_ _55288_/A _56889_/B _56889_/X sky130_fd_sc_hd__and2_4
X_49430_ _49428_/Y _49405_/X _49429_/X _49430_/Y sky130_fd_sc_hd__a21oi_4
X_70906_ _51008_/B _70885_/A _70905_/Y _83666_/D sky130_fd_sc_hd__o21ai_4
X_58628_ _58125_/X _85788_/Q _58126_/X _58628_/X sky130_fd_sc_hd__o21a_4
X_46642_ _52590_/B _51765_/B sky130_fd_sc_hd__buf_2
X_77462_ _77447_/X _77448_/Y _77442_/X _77462_/Y sky130_fd_sc_hd__a21boi_4
X_43854_ _43854_/A _43854_/X sky130_fd_sc_hd__buf_2
X_74674_ _74630_/X _57007_/X _74673_/Y _74674_/X sky130_fd_sc_hd__o21a_4
X_71886_ _71870_/Y _83340_/Q _71885_/Y _71886_/X sky130_fd_sc_hd__a21o_4
X_79201_ _79201_/A _79201_/Y sky130_fd_sc_hd__inv_2
X_76413_ _76409_/Y _76411_/Y _76408_/Y _76417_/C sky130_fd_sc_hd__o21ai_4
X_42805_ _42700_/A _42805_/X sky130_fd_sc_hd__buf_2
X_49361_ _49205_/A _49382_/A sky130_fd_sc_hd__buf_2
X_73625_ _87856_/Q _73624_/X _73625_/Y sky130_fd_sc_hd__nor2_4
X_46573_ _52563_/B _50870_/B sky130_fd_sc_hd__buf_2
X_70837_ _46625_/X _70831_/X _70836_/Y _70837_/Y sky130_fd_sc_hd__o21ai_4
X_58559_ _58423_/A _58559_/X sky130_fd_sc_hd__buf_2
X_77393_ _77406_/A _82094_/D _77394_/B sky130_fd_sc_hd__xor2_4
X_43785_ _43784_/Y _87269_/D sky130_fd_sc_hd__inv_2
X_40997_ _40996_/Y _40997_/Y sky130_fd_sc_hd__inv_2
X_48312_ _48088_/B _50356_/B sky130_fd_sc_hd__buf_2
X_79132_ _79132_/A _79132_/B _79132_/X sky130_fd_sc_hd__xor2_4
X_45524_ _45518_/X _45522_/X _45523_/X _45524_/X sky130_fd_sc_hd__a21o_4
X_76344_ _81648_/Q _76344_/Y sky130_fd_sc_hd__inv_2
X_42736_ _42736_/A _87744_/D sky130_fd_sc_hd__inv_2
X_61570_ _61541_/A _61570_/B _61541_/C _61570_/Y sky130_fd_sc_hd__nand3_4
X_49292_ _65054_/B _49204_/X _49291_/Y _49292_/Y sky130_fd_sc_hd__o21ai_4
X_73556_ _73553_/X _73555_/X _73489_/X _73556_/X sky130_fd_sc_hd__a21o_4
X_70768_ _70768_/A _70863_/A sky130_fd_sc_hd__buf_2
X_48243_ _49223_/A _48244_/A sky130_fd_sc_hd__buf_2
X_60521_ _60400_/Y _60430_/Y _60482_/A _60522_/A sky130_fd_sc_hd__nand3_4
X_72507_ _72507_/A _72508_/A sky130_fd_sc_hd__inv_2
X_79063_ _82830_/Q _82542_/Q _79064_/B sky130_fd_sc_hd__xnor2_4
X_45455_ _45455_/A _45455_/Y sky130_fd_sc_hd__inv_2
X_76275_ _81259_/Q _81515_/D _76276_/B sky130_fd_sc_hd__xor2_4
X_42667_ _42665_/X _42666_/X _41021_/X _87780_/Q _42658_/X _42667_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73487_ _73487_/A _72896_/B _73487_/Y sky130_fd_sc_hd__nor2_4
X_70699_ _70699_/A _70699_/X sky130_fd_sc_hd__buf_2
X_78014_ _77997_/A _78012_/A _82078_/Q _78013_/Y _78014_/X sky130_fd_sc_hd__a2bb2o_4
X_44406_ _44352_/X _44406_/X sky130_fd_sc_hd__buf_2
X_63240_ _60482_/Y _63240_/X sky130_fd_sc_hd__buf_2
X_75226_ _75226_/A _80985_/Q _75226_/Y sky130_fd_sc_hd__nand2_4
X_41618_ _41617_/Y _88182_/D sky130_fd_sc_hd__inv_2
X_48174_ _73588_/B _48170_/X _48173_/Y _48174_/Y sky130_fd_sc_hd__o21ai_4
X_60452_ _60387_/X _60430_/Y _60452_/X sky130_fd_sc_hd__and2_4
X_72438_ _72413_/X _72436_/Y _72437_/Y _57793_/X _72417_/X _72438_/X
+ sky130_fd_sc_hd__o32a_4
X_45386_ _45386_/A _55635_/B sky130_fd_sc_hd__inv_2
X_42598_ _42590_/X _42592_/X _40874_/X _87807_/Q _42597_/X _42599_/A
+ sky130_fd_sc_hd__o32ai_4
X_47125_ _47109_/A _52869_/B _47125_/Y sky130_fd_sc_hd__nand2_4
X_44337_ _44336_/Y _87160_/D sky130_fd_sc_hd__inv_2
X_63171_ _59413_/Y _63170_/X _63161_/C _63149_/X _63171_/X sky130_fd_sc_hd__or4_4
X_75157_ _75156_/Y _75157_/B _75153_/A _75161_/B sky130_fd_sc_hd__nand3_4
X_41549_ _41482_/A _41584_/B sky130_fd_sc_hd__buf_2
X_72369_ _72270_/X _72366_/Y _72368_/Y _72296_/X _72274_/X _72369_/X
+ sky130_fd_sc_hd__o32a_4
X_60383_ _60383_/A _60515_/C sky130_fd_sc_hd__buf_2
X_74108_ _72910_/A _74152_/A sky130_fd_sc_hd__buf_2
X_62122_ _62144_/A _62121_/X _62122_/C _62122_/Y sky130_fd_sc_hd__nor3_4
X_47056_ _46961_/X _47067_/A sky130_fd_sc_hd__buf_2
X_44268_ _44268_/A _43986_/A _44242_/C _44268_/Y sky130_fd_sc_hd__nand3_4
X_75088_ _75086_/A _75079_/B _75088_/Y sky130_fd_sc_hd__nand2_4
X_79965_ _79947_/Y _79948_/Y _79944_/Y _79965_/Y sky130_fd_sc_hd__o21ai_4
X_46007_ _45962_/X _46007_/X sky130_fd_sc_hd__buf_2
X_43219_ _40968_/X _43216_/X _87533_/Q _43218_/X _43219_/X sky130_fd_sc_hd__a2bb2o_4
X_66930_ _87428_/Q _66878_/X _66879_/X _66929_/X _66930_/X sky130_fd_sc_hd__a211o_4
X_62053_ _62049_/Y _62033_/X _62052_/Y _62053_/Y sky130_fd_sc_hd__a21oi_4
X_74039_ _74012_/X _86221_/Q _73948_/X _74038_/X _74039_/X sky130_fd_sc_hd__a211o_4
X_78916_ _78902_/Y _78903_/Y _82636_/Q _82508_/D _78916_/X sky130_fd_sc_hd__a2bb2o_4
X_44199_ _57043_/B _44220_/B sky130_fd_sc_hd__buf_2
X_79896_ _64200_/C _79896_/Y sky130_fd_sc_hd__inv_2
X_61004_ _61003_/Y _61004_/Y sky130_fd_sc_hd__inv_2
X_66861_ _66912_/A _66861_/B _66861_/X sky130_fd_sc_hd__and2_4
X_78847_ _78857_/B _78857_/A _78874_/B sky130_fd_sc_hd__xnor2_4
X_68600_ _88010_/Q _68527_/X _68501_/X _68599_/X _68600_/X sky130_fd_sc_hd__a211o_4
X_65812_ _65812_/A _86504_/Q _65812_/X sky130_fd_sc_hd__and2_4
X_69580_ _69580_/A _87314_/Q _69580_/X sky130_fd_sc_hd__and2_4
X_47958_ _47953_/Y _47954_/X _47957_/X _86582_/D sky130_fd_sc_hd__a21oi_4
X_66792_ _59801_/A _66910_/A sky130_fd_sc_hd__buf_2
X_78778_ _78778_/A _78778_/B _78778_/X sky130_fd_sc_hd__xor2_4
X_68531_ _87501_/Q _68504_/X _68450_/X _68530_/X _68531_/X sky130_fd_sc_hd__a211o_4
X_46909_ _46249_/A _46909_/X sky130_fd_sc_hd__buf_2
X_65743_ _64739_/A _65888_/A sky130_fd_sc_hd__buf_2
X_77729_ _77732_/B _77730_/A sky130_fd_sc_hd__inv_2
X_62955_ _62971_/A _84886_/Q _60302_/X _62979_/D _62955_/X sky130_fd_sc_hd__and4_4
X_47889_ _83556_/Q _73692_/A sky130_fd_sc_hd__inv_2
X_61906_ _57664_/X _61902_/X _61838_/X _61870_/X _61905_/X _61906_/X
+ sky130_fd_sc_hd__a41o_4
X_49628_ _86352_/Q _49606_/X _49627_/Y _49628_/Y sky130_fd_sc_hd__o21ai_4
X_80740_ _80740_/CLK _75108_/X _75042_/A sky130_fd_sc_hd__dfxtp_4
X_68462_ _68586_/A _68462_/X sky130_fd_sc_hd__buf_2
X_65674_ _65825_/A _86513_/Q _65674_/X sky130_fd_sc_hd__and2_4
X_62886_ _62886_/A _62886_/X sky130_fd_sc_hd__buf_2
X_67413_ _67410_/X _67413_/B _67413_/Y sky130_fd_sc_hd__nand2_4
X_64625_ _59345_/X _86176_/Q _64583_/X _64624_/X _64625_/X sky130_fd_sc_hd__a211o_4
X_49559_ _59044_/B _49551_/X _49558_/Y _49559_/Y sky130_fd_sc_hd__o21ai_4
X_61837_ _61823_/A _61823_/B _63448_/B _61788_/X _61837_/X sky130_fd_sc_hd__and4_4
X_80671_ _80671_/CLK _80671_/D _80671_/Q sky130_fd_sc_hd__dfxtp_4
X_68393_ _69607_/A _68394_/A sky130_fd_sc_hd__buf_2
X_82410_ _82443_/CLK _82410_/D _78417_/A sky130_fd_sc_hd__dfxtp_4
X_67344_ _67226_/A _67344_/X sky130_fd_sc_hd__buf_2
X_52570_ _52568_/Y _51951_/X _52569_/Y _85795_/D sky130_fd_sc_hd__a21boi_4
X_64556_ _64455_/X _61694_/B _61102_/X _64556_/Y sky130_fd_sc_hd__nand3_4
X_83390_ _85407_/CLK _83390_/D _83390_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_492_0_CLK clkbuf_9_246_0_CLK/X _86400_/CLK sky130_fd_sc_hd__clkbuf_1
X_61768_ _61752_/A _61723_/X _78078_/B _61768_/Y sky130_fd_sc_hd__nor3_4
XPHY_509 sky130_fd_sc_hd__decap_3
X_51521_ _51629_/A _51521_/X sky130_fd_sc_hd__buf_2
X_63507_ _63517_/A _63517_/B _80506_/B _63507_/Y sky130_fd_sc_hd__nor3_4
X_82341_ _86753_/CLK _82341_/D _82341_/Q sky130_fd_sc_hd__dfxtp_4
X_60719_ _59756_/A _60719_/X sky130_fd_sc_hd__buf_2
X_67275_ _67250_/A _86777_/Q _67275_/X sky130_fd_sc_hd__and2_4
X_64487_ _61182_/X _61618_/X _64211_/C _64487_/Y sky130_fd_sc_hd__nand3_4
X_61699_ _61645_/A _61699_/X sky130_fd_sc_hd__buf_2
X_69014_ _69014_/A _69059_/A sky130_fd_sc_hd__buf_2
X_54240_ _85478_/Q _54220_/X _54239_/Y _54240_/Y sky130_fd_sc_hd__o21ai_4
X_66226_ _66226_/A _86539_/Q _66226_/X sky130_fd_sc_hd__and2_4
X_85060_ _85034_/CLK _85060_/D _85060_/Q sky130_fd_sc_hd__dfxtp_4
X_51452_ _51456_/A _51473_/B _51467_/C _52977_/D _51452_/X sky130_fd_sc_hd__and4_4
X_63438_ _58424_/Y _63436_/X _61406_/A _63437_/X _63438_/X sky130_fd_sc_hd__a2bb2o_4
X_82272_ _82272_/CLK _82272_/D _82272_/Q sky130_fd_sc_hd__dfxtp_4
X_84011_ _81475_/CLK _68212_/X _84011_/Q sky130_fd_sc_hd__dfxtp_4
X_50403_ _50464_/A _50403_/X sky130_fd_sc_hd__buf_2
X_81223_ _85351_/CLK _81031_/Q _81223_/Q sky130_fd_sc_hd__dfxtp_4
X_54171_ _53436_/X _54171_/X sky130_fd_sc_hd__buf_2
X_66157_ _66154_/X _66156_/X _65961_/X _66453_/A sky130_fd_sc_hd__a21o_4
X_51383_ _86020_/Q _51362_/X _51382_/Y _51383_/Y sky130_fd_sc_hd__o21ai_4
X_63369_ _63410_/A _63369_/B _63384_/C _63384_/D _63369_/X sky130_fd_sc_hd__and4_4
X_53122_ _53121_/X _53122_/B _53122_/Y sky130_fd_sc_hd__nand2_4
X_65108_ _64991_/A _65108_/X sky130_fd_sc_hd__buf_2
X_50334_ _50213_/X _50398_/A sky130_fd_sc_hd__buf_2
X_81154_ _81154_/CLK _74849_/B _41624_/A sky130_fd_sc_hd__dfxtp_4
X_66088_ _65924_/X _84981_/Q _65950_/X _66087_/X _66426_/C sky130_fd_sc_hd__a211o_4
X_80105_ _80089_/X _80105_/B _80105_/X sky130_fd_sc_hd__or2_4
X_53053_ _53051_/Y _53028_/X _53052_/X _53053_/Y sky130_fd_sc_hd__a21oi_4
X_57930_ _57952_/A _86323_/Q _57930_/Y sky130_fd_sc_hd__nor2_4
X_65039_ _65033_/X _65038_/X _64959_/X _65039_/X sky130_fd_sc_hd__a21o_4
X_69916_ _64834_/A _69916_/X sky130_fd_sc_hd__buf_2
X_50265_ _86235_/Q _50250_/X _50264_/Y _50265_/Y sky130_fd_sc_hd__o21ai_4
X_85962_ _85962_/CLK _85962_/D _85962_/Q sky130_fd_sc_hd__dfxtp_4
X_81085_ _81087_/CLK _75669_/A _75473_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_430_0_CLK clkbuf_9_215_0_CLK/X _82833_/CLK sky130_fd_sc_hd__clkbuf_1
X_52004_ _52002_/Y _51981_/X _52003_/Y _85908_/D sky130_fd_sc_hd__a21boi_4
X_87701_ _88201_/CLK _42823_/X _87701_/Q sky130_fd_sc_hd__dfxtp_4
X_80036_ _80030_/Y _80035_/Y _80036_/X sky130_fd_sc_hd__xor2_4
X_84913_ _84906_/CLK _58185_/Y _84913_/Q sky130_fd_sc_hd__dfxtp_4
X_57861_ _57811_/X _85400_/Q _57860_/X _57861_/Y sky130_fd_sc_hd__o21ai_4
X_69847_ _83893_/Q _69831_/X _69846_/X _83893_/D sky130_fd_sc_hd__a21bo_4
X_50196_ _65327_/B _50185_/X _50195_/Y _50196_/Y sky130_fd_sc_hd__o21ai_4
X_85893_ _86203_/CLK _52080_/Y _85893_/Q sky130_fd_sc_hd__dfxtp_4
X_59600_ _60392_/B _60174_/C _60636_/B _60407_/A _59600_/X sky130_fd_sc_hd__and4_4
X_56812_ _56808_/Y _56811_/Y _56794_/Y _56688_/X _56812_/X sky130_fd_sc_hd__a211o_4
X_87632_ _87888_/CLK _42957_/X _87632_/Q sky130_fd_sc_hd__dfxtp_4
X_84844_ _84299_/CLK _84844_/D _84844_/Q sky130_fd_sc_hd__dfxtp_4
X_57792_ _57792_/A _57791_/X _57792_/Y sky130_fd_sc_hd__nor2_4
X_69778_ _73175_/A _69747_/X _68691_/X _69777_/Y _69778_/X sky130_fd_sc_hd__a211o_4
X_59531_ _61183_/A _59532_/A sky130_fd_sc_hd__inv_2
X_56743_ _56852_/A _57179_/A sky130_fd_sc_hd__buf_2
X_68729_ _73892_/A _68650_/X _68651_/X _68728_/Y _68729_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_445_0_CLK clkbuf_9_222_0_CLK/X _85351_/CLK sky130_fd_sc_hd__clkbuf_1
X_87563_ _83158_/CLK _43136_/Y _87563_/Q sky130_fd_sc_hd__dfxtp_4
X_53955_ _53921_/A _53955_/X sky130_fd_sc_hd__buf_2
X_84775_ _86688_/CLK _84775_/D _84775_/Q sky130_fd_sc_hd__dfxtp_4
X_81987_ _82104_/CLK _81987_/D _77013_/A sky130_fd_sc_hd__dfxtp_4
X_86514_ _83572_/CLK _86514_/D _86514_/Q sky130_fd_sc_hd__dfxtp_4
X_40920_ _40877_/X _82852_/Q _40919_/X _40921_/A sky130_fd_sc_hd__o21ai_4
X_52906_ _85733_/Q _52902_/X _52905_/Y _52906_/Y sky130_fd_sc_hd__o21ai_4
X_71740_ _71753_/D _71744_/D sky130_fd_sc_hd__buf_2
X_83726_ _85381_/CLK _83726_/D _47480_/A sky130_fd_sc_hd__dfxtp_4
X_59462_ _58982_/A _59462_/X sky130_fd_sc_hd__buf_2
X_56674_ _56655_/A _56674_/X sky130_fd_sc_hd__buf_2
X_80938_ _80776_/CLK _80938_/D _74906_/A sky130_fd_sc_hd__dfxtp_4
X_87494_ _87749_/CLK _87494_/D _87494_/Q sky130_fd_sc_hd__dfxtp_4
X_53886_ _53871_/X _53886_/B _53886_/Y sky130_fd_sc_hd__nand2_4
X_58413_ _58406_/X _83367_/Q _58412_/Y _58413_/X sky130_fd_sc_hd__o21a_4
X_55625_ _44087_/B _55625_/B _55625_/Y sky130_fd_sc_hd__nor2_4
X_86445_ _86155_/CLK _86445_/D _86445_/Q sky130_fd_sc_hd__dfxtp_4
X_40851_ _40850_/Y _88323_/D sky130_fd_sc_hd__inv_2
X_52837_ _52843_/A _52837_/B _52837_/Y sky130_fd_sc_hd__nand2_4
X_71671_ _71641_/A _71671_/X sky130_fd_sc_hd__buf_2
X_59393_ _58982_/X _83488_/Q _59392_/Y _84744_/D sky130_fd_sc_hd__o21a_4
X_83657_ _85822_/CLK _83657_/D _46242_/A sky130_fd_sc_hd__dfxtp_4
X_80869_ _81125_/CLK _75604_/B _80837_/D sky130_fd_sc_hd__dfxtp_4
X_73410_ _48639_/A _73409_/Y _73410_/X sky130_fd_sc_hd__xor2_4
X_70622_ _70824_/A _70727_/A sky130_fd_sc_hd__buf_2
X_82608_ _82702_/CLK _78939_/B _82576_/D sky130_fd_sc_hd__dfxtp_4
X_58344_ _58344_/A _58344_/B _58344_/Y sky130_fd_sc_hd__nor2_4
X_43570_ _43557_/X _43563_/X _40515_/X _87355_/Q _43058_/A _43570_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55556_ _45504_/A _55522_/X _55513_/X _55555_/Y _55556_/X sky130_fd_sc_hd__a211o_4
X_86376_ _83666_/CLK _86376_/D _86376_/Q sky130_fd_sc_hd__dfxtp_4
X_74390_ _83076_/Q _74387_/X _74389_/Y _74390_/Y sky130_fd_sc_hd__o21ai_4
X_40782_ _40781_/X _40754_/X _69612_/B _40756_/X _88336_/D sky130_fd_sc_hd__a2bb2o_4
X_52768_ _52773_/A _52768_/B _52768_/Y sky130_fd_sc_hd__nand2_4
X_83588_ _86525_/CLK _71156_/Y _83588_/Q sky130_fd_sc_hd__dfxtp_4
X_88115_ _88108_/CLK _88115_/D _73552_/A sky130_fd_sc_hd__dfxtp_4
X_42521_ _42610_/A _42521_/X sky130_fd_sc_hd__buf_2
X_54507_ _54481_/A _54509_/A sky130_fd_sc_hd__buf_2
X_73341_ _73341_/A _73196_/B _73341_/Y sky130_fd_sc_hd__nor2_4
X_85327_ _83550_/CLK _85327_/D _85327_/Q sky130_fd_sc_hd__dfxtp_4
X_51719_ _51719_/A _51719_/X sky130_fd_sc_hd__buf_2
X_70553_ _70552_/Y _71859_/A sky130_fd_sc_hd__buf_2
X_58275_ _58271_/X _83443_/Q _58274_/Y _84891_/D sky130_fd_sc_hd__o21a_4
X_82539_ _82541_/CLK _83859_/Q _82539_/Q sky130_fd_sc_hd__dfxtp_4
X_55487_ _55453_/X _55489_/A sky130_fd_sc_hd__buf_2
X_52699_ _52697_/Y _52673_/X _52698_/X _52699_/Y sky130_fd_sc_hd__a21oi_4
X_45240_ _56523_/C _45209_/X _45189_/X _45240_/X sky130_fd_sc_hd__o21a_4
X_57226_ _45947_/B _85059_/Q _57225_/Y _57158_/C _57226_/X sky130_fd_sc_hd__a211o_4
X_76060_ _76057_/Y _76060_/B _76061_/B sky130_fd_sc_hd__xor2_4
X_88046_ _87789_/CLK _42074_/X _88046_/Q sky130_fd_sc_hd__dfxtp_4
X_54438_ _85442_/Q _54431_/X _54437_/Y _54438_/Y sky130_fd_sc_hd__o21ai_4
X_42452_ _42488_/A _42612_/A sky130_fd_sc_hd__buf_2
X_73272_ _83158_/Q _73193_/X _73271_/Y _73272_/X sky130_fd_sc_hd__a21o_4
X_85258_ _85257_/CLK _56254_/Y _56253_/C sky130_fd_sc_hd__dfxtp_4
X_70484_ _70466_/Y _83764_/Q _70483_/X _83764_/D sky130_fd_sc_hd__a21o_4
X_75011_ _75001_/Y _75004_/X _74999_/X _75011_/Y sky130_fd_sc_hd__a21boi_4
X_41403_ _41402_/X _41403_/X sky130_fd_sc_hd__buf_2
X_72223_ _72214_/Y _72152_/X _72219_/X _72222_/X _83273_/D sky130_fd_sc_hd__a22oi_4
X_84209_ _85315_/CLK _65246_/X _84209_/Q sky130_fd_sc_hd__dfxtp_4
X_45171_ _64411_/B _61538_/B sky130_fd_sc_hd__buf_2
X_57157_ _56801_/X _57170_/B _57155_/D _57156_/X _57003_/B _57158_/B
+ sky130_fd_sc_hd__a41oi_4
X_42383_ _41797_/X _42374_/X _87891_/Q _42375_/X _87891_/D sky130_fd_sc_hd__a2bb2o_4
X_54369_ _54355_/A _52677_/B _54369_/Y sky130_fd_sc_hd__nand2_4
X_85189_ _85156_/CLK _85189_/D _56450_/C sky130_fd_sc_hd__dfxtp_4
X_44122_ HASH_EN _44196_/B sky130_fd_sc_hd__buf_2
X_56108_ _56108_/A _56108_/B _56109_/A sky130_fd_sc_hd__xnor2_4
X_41334_ _41239_/X _41241_/X _41332_/X _67553_/B _41333_/X _41334_/Y
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_9_504_0_CLK clkbuf_9_505_0_CLK/A clkbuf_9_504_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_72154_ _59231_/X _85374_/Q _72153_/X _72154_/Y sky130_fd_sc_hd__o21ai_4
X_57088_ _72814_/A _73183_/A sky130_fd_sc_hd__buf_2
X_71105_ _49073_/X _71095_/X _71104_/Y _83606_/D sky130_fd_sc_hd__o21ai_4
X_48930_ _48930_/A _48931_/A sky130_fd_sc_hd__inv_2
X_56039_ _55927_/X _56001_/A _56039_/Y sky130_fd_sc_hd__xnor2_4
X_44053_ _44053_/A _44202_/A sky130_fd_sc_hd__inv_2
X_79750_ _79728_/Y _79746_/X _79749_/Y _79750_/Y sky130_fd_sc_hd__a21oi_4
X_41265_ _41264_/X _41251_/X _88248_/Q _41253_/X _41265_/X sky130_fd_sc_hd__a2bb2o_4
X_72085_ _72082_/Y _72083_/X _72084_/Y _83288_/D sky130_fd_sc_hd__a21boi_4
X_76962_ _76840_/Y _81367_/D sky130_fd_sc_hd__inv_2
X_43004_ _40528_/X _42994_/X _87608_/Q _42995_/X _43004_/X sky130_fd_sc_hd__a2bb2o_4
X_78701_ _78701_/A _78701_/B _78701_/X sky130_fd_sc_hd__and2_4
X_71036_ _71181_/A _71030_/B _71030_/C _71039_/D _71036_/Y sky130_fd_sc_hd__nand4_4
X_75913_ _84511_/Q _84383_/Q _75913_/X sky130_fd_sc_hd__xor2_4
X_48861_ _48836_/A _48861_/X sky130_fd_sc_hd__buf_2
X_79681_ _79679_/X _79681_/B _79682_/B sky130_fd_sc_hd__xnor2_4
X_41196_ _41196_/A _88260_/D sky130_fd_sc_hd__inv_2
X_76893_ _76893_/A _76893_/Y sky130_fd_sc_hd__inv_2
X_47812_ _49379_/A _49374_/A sky130_fd_sc_hd__buf_2
X_78632_ _78628_/Y _78632_/B _78632_/C _78632_/X sky130_fd_sc_hd__or3_4
X_75844_ _75836_/A _75836_/B _75843_/Y _75844_/Y sky130_fd_sc_hd__o21ai_4
X_48792_ _48789_/Y _48785_/X _48791_/X _48792_/Y sky130_fd_sc_hd__a21oi_4
X_47743_ _47715_/X _53219_/B _47743_/Y sky130_fd_sc_hd__nand2_4
X_59729_ _59635_/Y _59730_/A sky130_fd_sc_hd__buf_2
X_78563_ _78563_/A _78562_/X _82771_/D sky130_fd_sc_hd__xor2_4
X_44955_ _44948_/X _44952_/X _44954_/Y _44955_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_8_72_0_CLK clkbuf_8_73_0_CLK/A clkbuf_8_72_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_75775_ _75759_/B _75772_/X _75774_/Y _75775_/Y sky130_fd_sc_hd__a21oi_4
X_72987_ _72978_/A _86201_/Q _72985_/X _72986_/X _72987_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_7_4_0_CLK clkbuf_6_2_0_CLK/X clkbuf_8_9_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_77514_ _77514_/A _77514_/B _82197_/D sky130_fd_sc_hd__xnor2_4
X_43906_ _41356_/X _43886_/X _67644_/B _43887_/X _43906_/X sky130_fd_sc_hd__a2bb2o_4
X_62740_ _62727_/A _62727_/B _61844_/X _62740_/Y sky130_fd_sc_hd__nand3_4
X_74726_ _70730_/X _74796_/C sky130_fd_sc_hd__buf_2
X_47674_ _47674_/A _47675_/A sky130_fd_sc_hd__inv_2
X_71938_ _70554_/A _71411_/B _71938_/Y sky130_fd_sc_hd__nor2_4
X_78494_ _78494_/A _78515_/A sky130_fd_sc_hd__buf_2
X_44886_ _85217_/Q _44880_/X _44885_/X _44886_/Y sky130_fd_sc_hd__o21ai_4
X_49413_ _49420_/A _49420_/B _49420_/C _46707_/X _49413_/X sky130_fd_sc_hd__and4_4
X_46625_ _46624_/Y _46625_/X sky130_fd_sc_hd__buf_2
X_77445_ _77444_/A _77444_/B _77446_/A sky130_fd_sc_hd__nand2_4
X_43837_ _41165_/X _43832_/X _68627_/B _43833_/X _87241_/D sky130_fd_sc_hd__a2bb2o_4
X_62671_ _62671_/A _62673_/A sky130_fd_sc_hd__buf_2
X_74657_ _74694_/A _45638_/A _74657_/Y sky130_fd_sc_hd__nand2_4
X_71869_ _71823_/A _71713_/Y _70454_/Y _71870_/A sky130_fd_sc_hd__nor3_4
X_64410_ _63573_/A _61226_/X _64410_/Y sky130_fd_sc_hd__nor2_4
X_49344_ _49352_/A _51378_/B _49344_/Y sky130_fd_sc_hd__nand2_4
X_73608_ _73605_/X _86239_/Q _44194_/X _73607_/X _73608_/X sky130_fd_sc_hd__a211o_4
X_61622_ _61621_/X _61622_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_87_0_CLK clkbuf_8_87_0_CLK/A clkbuf_8_87_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_46556_ _46547_/A _50862_/B _46556_/Y sky130_fd_sc_hd__nand2_4
X_65390_ _65385_/X _65388_/X _65389_/X _65390_/X sky130_fd_sc_hd__a21o_4
X_77376_ _77376_/A _77376_/B _77376_/Y sky130_fd_sc_hd__nand2_4
X_43768_ _43767_/Y _43768_/Y sky130_fd_sc_hd__inv_2
X_74588_ _56094_/X _74625_/A _74587_/Y _83025_/D sky130_fd_sc_hd__a21boi_4
X_79115_ _79115_/A _79115_/Y sky130_fd_sc_hd__inv_2
X_45507_ _45705_/A _45507_/X sky130_fd_sc_hd__buf_2
X_64341_ _59403_/A _64316_/B _64341_/Y sky130_fd_sc_hd__nor2_4
X_76327_ _76328_/A _81518_/D _76327_/Y sky130_fd_sc_hd__nor2_4
X_42719_ _41169_/X _42717_/X _87752_/Q _42718_/X _87752_/D sky130_fd_sc_hd__a2bb2o_4
X_49275_ _49261_/A _46412_/B _49275_/Y sky130_fd_sc_hd__nand2_4
X_61553_ _61553_/A _61553_/Y sky130_fd_sc_hd__inv_2
X_73539_ _73536_/X _73538_/X _72949_/X _73542_/A sky130_fd_sc_hd__a21o_4
X_46487_ _52524_/A _46487_/B _46472_/C _46487_/X sky130_fd_sc_hd__and3_4
X_43699_ _87303_/Q _69722_/B sky130_fd_sc_hd__inv_2
X_48226_ _48226_/A _48226_/X sky130_fd_sc_hd__buf_2
X_60504_ _60503_/X _60595_/C sky130_fd_sc_hd__buf_2
X_67060_ _87359_/Q _67035_/X _66984_/X _67059_/X _67060_/X sky130_fd_sc_hd__a211o_4
X_79046_ _79045_/X _79047_/B sky130_fd_sc_hd__buf_2
X_45438_ _85086_/Q _45438_/Y sky130_fd_sc_hd__inv_2
X_64272_ _64272_/A _64301_/B _64272_/Y sky130_fd_sc_hd__nor2_4
X_76258_ _76268_/D _76257_/Y _76258_/Y sky130_fd_sc_hd__xnor2_4
X_61484_ _59407_/A _61484_/B _61484_/C _61452_/D _61485_/A sky130_fd_sc_hd__nand4_4
Xclkbuf_8_10_0_CLK clkbuf_7_5_0_CLK/X clkbuf_8_10_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_66011_ _64611_/A _66011_/X sky130_fd_sc_hd__buf_2
X_75209_ _75196_/Y _75189_/X _75190_/Y _75210_/B sky130_fd_sc_hd__a21boi_4
X_63223_ _58385_/Y _63190_/X _63175_/X _58261_/Y _63176_/X _63223_/Y
+ sky130_fd_sc_hd__o32ai_4
X_48157_ _47943_/A _48157_/B _48157_/X sky130_fd_sc_hd__or2_4
X_60435_ _60435_/A _72577_/B _60435_/C _60435_/Y sky130_fd_sc_hd__nand3_4
X_45369_ _45369_/A _45452_/A sky130_fd_sc_hd__buf_2
X_76189_ _76189_/A _76189_/B _76187_/Y _76193_/C sky130_fd_sc_hd__nand3_4
X_47108_ _53373_/B _52859_/B sky130_fd_sc_hd__buf_2
X_63154_ _60452_/X _63154_/X sky130_fd_sc_hd__buf_2
X_60366_ _60359_/X _60363_/Y _59892_/Y _60285_/A _60365_/Y _60366_/Y
+ sky130_fd_sc_hd__a41oi_4
X_48088_ _48138_/A _48088_/B _48088_/X sky130_fd_sc_hd__and2_4
X_62105_ _59668_/B _62105_/X sky130_fd_sc_hd__buf_2
X_47039_ _47029_/A _47039_/B _47029_/C _52818_/D _47039_/X sky130_fd_sc_hd__and4_4
Xclkbuf_8_25_0_CLK clkbuf_8_25_0_CLK/A clkbuf_9_51_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_67962_ _68028_/A _87641_/Q _67962_/X sky130_fd_sc_hd__and2_4
X_79948_ _79932_/A _79931_/B _79928_/Y _79948_/Y sky130_fd_sc_hd__a21oi_4
X_63085_ _63038_/A _64294_/B _63085_/C _63085_/D _63085_/X sky130_fd_sc_hd__and4_4
X_60297_ _57686_/A _59741_/A _59705_/X _62640_/C _60298_/C sky130_fd_sc_hd__nand4_4
X_69701_ _73036_/A _68377_/X _66574_/X _69700_/Y _69701_/X sky130_fd_sc_hd__a211o_4
X_50050_ _50050_/A _50045_/X _51750_/C _53261_/D _50050_/X sky130_fd_sc_hd__and4_4
X_66913_ _87877_/Q _66816_/X _66911_/X _66912_/X _66913_/X sky130_fd_sc_hd__a211o_4
X_62036_ _59721_/A _62094_/B sky130_fd_sc_hd__buf_2
X_67893_ _67890_/X _67892_/X _67799_/X _67893_/X sky130_fd_sc_hd__a21o_4
X_79879_ _79874_/X _79878_/Y _79879_/X sky130_fd_sc_hd__xor2_4
X_81910_ _82005_/CLK _81910_/D _81910_/Q sky130_fd_sc_hd__dfxtp_4
X_69632_ _69696_/A _69632_/X sky130_fd_sc_hd__buf_2
X_66844_ _66839_/X _66842_/X _66843_/X _66844_/X sky130_fd_sc_hd__a21o_4
X_82890_ _83987_/CLK _78139_/B _41747_/A sky130_fd_sc_hd__dfxtp_4
X_81841_ _81094_/CLK _81841_/D _77444_/A sky130_fd_sc_hd__dfxtp_4
X_69563_ _83914_/Q _69504_/X _69562_/X _83914_/D sky130_fd_sc_hd__a21bo_4
X_66775_ _87371_/Q _66678_/X _66747_/X _66774_/X _66775_/X sky130_fd_sc_hd__a211o_4
X_63987_ _61969_/X _63955_/X _64050_/C _64033_/D _63987_/Y sky130_fd_sc_hd__nand4_4
X_68514_ _68376_/X _66524_/B _68500_/Y _68513_/Y _68514_/X sky130_fd_sc_hd__a211o_4
X_53740_ _53737_/Y _53715_/X _53739_/X _85578_/D sky130_fd_sc_hd__a21oi_4
X_65726_ _65516_/X _65102_/Y _65725_/Y _65726_/Y sky130_fd_sc_hd__o21ai_4
X_84560_ _84562_/CLK _84560_/D _84560_/Q sky130_fd_sc_hd__dfxtp_4
X_50952_ _50952_/A _50963_/C sky130_fd_sc_hd__buf_2
X_62938_ _61629_/B _62936_/X _62982_/C _62908_/X _62938_/Y sky130_fd_sc_hd__nand4_4
X_69494_ _69454_/A _69494_/B _69494_/X sky130_fd_sc_hd__and2_4
X_81772_ _82368_/CLK _81772_/D _81772_/Q sky130_fd_sc_hd__dfxtp_4
X_83511_ _83507_/CLK _83511_/D _83511_/Q sky130_fd_sc_hd__dfxtp_4
X_80723_ _80676_/CLK _80723_/D _80691_/D sky130_fd_sc_hd__dfxtp_4
X_68445_ _44675_/A _68023_/X _68024_/X _68444_/X _68445_/X sky130_fd_sc_hd__a211o_4
X_65657_ _65735_/A _86482_/Q _65657_/X sky130_fd_sc_hd__and2_4
X_53671_ _53671_/A _53692_/C sky130_fd_sc_hd__buf_2
X_84491_ _84241_/CLK _61273_/X _84491_/Q sky130_fd_sc_hd__dfxtp_4
X_50883_ _50728_/A _50906_/A sky130_fd_sc_hd__buf_2
X_62869_ _62869_/A _62935_/B _63585_/B _62869_/Y sky130_fd_sc_hd__nand3_4
X_55410_ _55399_/X _55409_/Y _55410_/Y sky130_fd_sc_hd__nand2_4
X_86230_ _86235_/CLK _50292_/Y _86230_/Q sky130_fd_sc_hd__dfxtp_4
X_52622_ _52643_/A _52605_/X _52622_/C _52622_/D _52622_/X sky130_fd_sc_hd__and4_4
X_64608_ _64608_/A _66195_/B sky130_fd_sc_hd__buf_2
X_83442_ _83763_/CLK _71601_/X _83442_/Q sky130_fd_sc_hd__dfxtp_4
X_56390_ _56383_/X _56386_/B _56390_/C _56390_/Y sky130_fd_sc_hd__nand3_4
X_80654_ _86772_/CLK _80654_/D _74846_/B sky130_fd_sc_hd__dfxtp_4
X_68376_ _68376_/A _68376_/X sky130_fd_sc_hd__buf_2
X_65588_ _65559_/A _65559_/B _84191_/Q _65588_/X sky130_fd_sc_hd__and3_4
X_55341_ _55445_/B _55445_/D _55362_/A sky130_fd_sc_hd__and2_4
X_67327_ _67305_/X _67316_/Y _67269_/X _67326_/Y _67327_/X sky130_fd_sc_hd__a211o_4
X_86161_ _85557_/CLK _50648_/Y _86161_/Q sky130_fd_sc_hd__dfxtp_4
X_52553_ _52542_/X _54071_/B _52553_/Y sky130_fd_sc_hd__nand2_4
XPHY_306 sky130_fd_sc_hd__decap_3
X_64539_ _64534_/X _64535_/X _64536_/X _64538_/Y _64219_/B _64539_/X
+ sky130_fd_sc_hd__o41a_4
X_83373_ _83372_/CLK _71795_/Y _83373_/Q sky130_fd_sc_hd__dfxtp_4
X_80585_ _84773_/Q _65970_/C _80585_/Y sky130_fd_sc_hd__nand2_4
XPHY_317 sky130_fd_sc_hd__decap_3
XPHY_328 sky130_fd_sc_hd__decap_3
X_85112_ _85144_/CLK _85112_/D _45535_/A sky130_fd_sc_hd__dfxtp_4
XPHY_339 sky130_fd_sc_hd__decap_3
X_51504_ _51504_/A _51527_/B sky130_fd_sc_hd__buf_2
X_58060_ _86632_/Q _58136_/B _58060_/Y sky130_fd_sc_hd__nor2_4
X_82324_ _82327_/CLK _77132_/B _82324_/Q sky130_fd_sc_hd__dfxtp_4
X_55272_ _55272_/A _55272_/X sky130_fd_sc_hd__buf_2
X_67258_ _80901_/D _67211_/X _67257_/X _67258_/X sky130_fd_sc_hd__a21bo_4
X_86092_ _85773_/CLK _51002_/Y _86092_/Q sky130_fd_sc_hd__dfxtp_4
X_52484_ _52476_/A _52484_/B _52484_/Y sky130_fd_sc_hd__nand2_4
X_57011_ _56783_/X _56700_/Y _56768_/Y _57024_/D _57011_/Y sky130_fd_sc_hd__nand4_4
X_54223_ _54230_/A _53054_/B _54223_/Y sky130_fd_sc_hd__nand2_4
X_66209_ _65763_/A _66209_/B _66209_/X sky130_fd_sc_hd__and2_4
X_85043_ _85042_/CLK _85043_/D _45617_/A sky130_fd_sc_hd__dfxtp_4
X_51435_ _51430_/X _52965_/B _51435_/Y sky130_fd_sc_hd__nand2_4
X_82255_ _85381_/CLK _80438_/Y _82255_/Q sky130_fd_sc_hd__dfxtp_4
X_67189_ _87929_/Q _67117_/X _67167_/X _67188_/X _67189_/X sky130_fd_sc_hd__a211o_4
X_81206_ _81197_/CLK _75045_/X _48996_/A sky130_fd_sc_hd__dfxtp_4
X_54154_ _85494_/Q _54140_/X _54153_/Y _54154_/Y sky130_fd_sc_hd__o21ai_4
X_51366_ _51793_/A _51366_/X sky130_fd_sc_hd__buf_2
X_82186_ _84951_/CLK _82186_/D _82186_/Q sky130_fd_sc_hd__dfxtp_4
X_53105_ _53115_/A _53105_/B _53105_/Y sky130_fd_sc_hd__nand2_4
X_50317_ _50500_/A _50317_/X sky130_fd_sc_hd__buf_2
X_81137_ _80968_/CLK _81137_/D _40676_/A sky130_fd_sc_hd__dfxtp_4
X_58962_ _58961_/X _85922_/Q _58900_/X _58962_/X sky130_fd_sc_hd__o21a_4
X_54085_ _54068_/X _46585_/Y _54085_/Y sky130_fd_sc_hd__nand2_4
X_51297_ _64920_/B _51285_/X _51296_/Y _51297_/Y sky130_fd_sc_hd__o21ai_4
X_86994_ _86998_/CLK _44702_/Y _86994_/Q sky130_fd_sc_hd__dfxtp_4
X_41050_ _41050_/A _41050_/X sky130_fd_sc_hd__buf_2
X_53036_ _53048_/A _53036_/B _53058_/C _53036_/D _53036_/X sky130_fd_sc_hd__and4_4
X_57913_ _57884_/X _85492_/Q _57763_/X _57913_/X sky130_fd_sc_hd__o21a_4
X_50248_ _48196_/A _74509_/C _50247_/X _50248_/X sky130_fd_sc_hd__and3_4
X_85945_ _82774_/CLK _51795_/Y _85945_/Q sky130_fd_sc_hd__dfxtp_4
X_81068_ _80813_/CLK _81100_/Q _81068_/Q sky130_fd_sc_hd__dfxtp_4
X_58893_ _58891_/X _86088_/Q _58892_/X _58893_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_490_0_CLK clkbuf_9_491_0_CLK/A clkbuf_9_490_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_72910_ _72910_/A _73381_/A sky130_fd_sc_hd__buf_2
X_80019_ _80019_/A _80018_/X _80019_/Y sky130_fd_sc_hd__xnor2_4
X_57844_ _58805_/A _58676_/A sky130_fd_sc_hd__buf_2
X_50179_ _50693_/A _50693_/B _47848_/X _50179_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_10_384_0_CLK clkbuf_9_192_0_CLK/X _83218_/CLK sky130_fd_sc_hd__clkbuf_1
X_85876_ _86193_/CLK _85876_/D _85876_/Q sky130_fd_sc_hd__dfxtp_4
X_73890_ _70101_/Y _73818_/X _73889_/X _83132_/D sky130_fd_sc_hd__o21ai_4
X_87615_ _82888_/CLK _42992_/Y _87615_/Q sky130_fd_sc_hd__dfxtp_4
X_72841_ _72750_/X _85598_/Q _72839_/X _72840_/X _72841_/X sky130_fd_sc_hd__a211o_4
X_84827_ _84829_/CLK _84827_/D _64379_/C sky130_fd_sc_hd__dfxtp_4
X_57775_ _72476_/B _86013_/Q _57774_/X _57775_/Y sky130_fd_sc_hd__o21ai_4
X_54987_ _54964_/A _54978_/X _54974_/C _47578_/A _54987_/X sky130_fd_sc_hd__and4_4
X_59514_ _59538_/C _59521_/A sky130_fd_sc_hd__inv_2
X_44740_ _44528_/A _44740_/X sky130_fd_sc_hd__buf_2
X_56726_ _56684_/C _56726_/X sky130_fd_sc_hd__buf_2
X_75560_ _75559_/X _75561_/B sky130_fd_sc_hd__inv_2
X_87546_ _88062_/CLK _87546_/D _43190_/A sky130_fd_sc_hd__dfxtp_4
X_53938_ _50209_/A _53875_/B _53888_/C _53938_/X sky130_fd_sc_hd__and3_4
X_41952_ _41881_/A _42025_/A sky130_fd_sc_hd__buf_2
X_72772_ _87314_/Q _72924_/B _72772_/Y sky130_fd_sc_hd__nor2_4
X_84758_ _84760_/CLK _59243_/Y _59229_/A sky130_fd_sc_hd__dfxtp_4
X_74511_ _74466_/A _48704_/Y _74511_/Y sky130_fd_sc_hd__nand2_4
X_40903_ _40903_/A _40903_/X sky130_fd_sc_hd__buf_2
X_71723_ _70504_/A _71729_/A sky130_fd_sc_hd__buf_2
X_83709_ _83707_/CLK _70750_/Y _47561_/A sky130_fd_sc_hd__dfxtp_4
X_59445_ _59445_/A _59444_/X _59445_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_399_0_CLK clkbuf_9_199_0_CLK/X _84187_/CLK sky130_fd_sc_hd__clkbuf_1
X_44671_ _44658_/X _44659_/X _40573_/X _87006_/Q _44660_/X _44672_/A
+ sky130_fd_sc_hd__o32ai_4
X_56657_ _56912_/A _56645_/Y _56660_/A sky130_fd_sc_hd__nand2_4
X_87477_ _87952_/CLK _43332_/Y _87477_/Q sky130_fd_sc_hd__dfxtp_4
X_75491_ _75488_/Y _75491_/B _75491_/C _75492_/A sky130_fd_sc_hd__nand3_4
X_41883_ _57491_/B _41879_/X _40581_/X _73595_/A _41882_/X _41884_/A
+ sky130_fd_sc_hd__o32ai_4
X_53869_ _53729_/A _53869_/X sky130_fd_sc_hd__buf_2
X_84689_ _84358_/CLK _84689_/D _80371_/A sky130_fd_sc_hd__dfxtp_4
X_46410_ _46410_/A _46411_/A sky130_fd_sc_hd__inv_2
X_77230_ _77230_/A _77230_/B _77230_/C _77230_/Y sky130_fd_sc_hd__nand3_4
X_43622_ _43622_/A _43622_/Y sky130_fd_sc_hd__inv_2
X_55608_ _85119_/Q _55605_/X _44090_/B _55607_/Y _55608_/X sky130_fd_sc_hd__a211o_4
X_74442_ _46280_/A _74442_/X sky130_fd_sc_hd__buf_2
X_86428_ _86246_/CLK _49236_/Y _64749_/B sky130_fd_sc_hd__dfxtp_4
X_40834_ _40833_/Y _88326_/D sky130_fd_sc_hd__inv_2
X_47390_ _81808_/Q _47391_/A sky130_fd_sc_hd__inv_2
X_59376_ _59326_/X _59376_/B _59376_/Y sky130_fd_sc_hd__nor2_4
X_71654_ _70426_/A _71660_/A sky130_fd_sc_hd__buf_2
X_56588_ _72648_/C _55570_/X _56589_/A sky130_fd_sc_hd__xnor2_4
X_46341_ _46336_/Y _46258_/X _46340_/Y _86746_/D sky130_fd_sc_hd__a21boi_4
X_70605_ _70994_/A _70717_/A sky130_fd_sc_hd__buf_2
X_58327_ _58310_/X _83453_/Q _58326_/Y _84877_/D sky130_fd_sc_hd__o21a_4
X_77161_ _77161_/A _77161_/B _77161_/X sky130_fd_sc_hd__xor2_4
X_55539_ _55498_/X _55539_/B _55539_/Y sky130_fd_sc_hd__nor2_4
X_43553_ _43553_/A _87364_/D sky130_fd_sc_hd__inv_2
X_74373_ _72068_/A _74373_/B _74373_/Y sky130_fd_sc_hd__nand2_4
X_86359_ _86359_/CLK _86359_/D _86359_/Q sky130_fd_sc_hd__dfxtp_4
X_40765_ _82881_/Q _40765_/B _40765_/X sky130_fd_sc_hd__or2_4
X_71585_ _71585_/A _71590_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_322_0_CLK clkbuf_9_161_0_CLK/X _86651_/CLK sky130_fd_sc_hd__clkbuf_1
X_76112_ _76112_/A _76112_/B _76113_/B sky130_fd_sc_hd__xor2_4
X_42504_ _42495_/X _42496_/X _40682_/X _68801_/A _42480_/X _42505_/A
+ sky130_fd_sc_hd__o32ai_4
X_49060_ _49060_/A _50142_/A sky130_fd_sc_hd__buf_2
X_73324_ _69862_/B _44128_/X _72858_/X _73323_/Y _73324_/X sky130_fd_sc_hd__a211o_4
X_46272_ _46272_/A _50738_/B _46272_/Y sky130_fd_sc_hd__nand2_4
X_70536_ _71012_/A _70692_/B sky130_fd_sc_hd__buf_2
X_58258_ _58258_/A _58259_/A sky130_fd_sc_hd__inv_2
Xclkbuf_10_952_0_CLK clkbuf_9_476_0_CLK/X _87824_/CLK sky130_fd_sc_hd__clkbuf_1
X_77092_ _77097_/A _77096_/A _77091_/Y _77093_/B sky130_fd_sc_hd__a21boi_4
X_43484_ _43513_/A _43484_/X sky130_fd_sc_hd__buf_2
X_40696_ _40695_/Y _40696_/X sky130_fd_sc_hd__buf_2
X_48011_ _48011_/A _50314_/A sky130_fd_sc_hd__buf_2
X_45223_ _85228_/Q _45206_/X _45161_/X _45223_/X sky130_fd_sc_hd__o21a_4
X_57209_ _57208_/Y _57129_/A _56704_/X _57209_/Y sky130_fd_sc_hd__a21oi_4
X_76043_ _76039_/B _76047_/A _76042_/Y _76043_/Y sky130_fd_sc_hd__a21boi_4
X_42435_ _41911_/A _42435_/X sky130_fd_sc_hd__buf_2
X_88029_ _87767_/CLK _42113_/X _88029_/Q sky130_fd_sc_hd__dfxtp_4
X_73255_ _69826_/B _73086_/X _73202_/X _73255_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_9_443_0_CLK clkbuf_9_443_0_CLK/A clkbuf_9_443_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_70467_ _71337_/A _71706_/A sky130_fd_sc_hd__buf_2
X_58189_ _57677_/X _58186_/Y _58188_/Y _84912_/D sky130_fd_sc_hd__a21oi_4
X_60220_ _60220_/A _60344_/C sky130_fd_sc_hd__buf_2
X_72206_ _72137_/X _72204_/Y _72205_/Y _72194_/X _72141_/X _72206_/X
+ sky130_fd_sc_hd__o32a_4
X_45154_ _85297_/Q _45120_/X _45153_/X _45154_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_10_337_0_CLK clkbuf_9_168_0_CLK/X _85735_/CLK sky130_fd_sc_hd__clkbuf_1
X_42366_ _42350_/X _42346_/X _41762_/X _87898_/Q _42347_/X _42367_/A
+ sky130_fd_sc_hd__o32ai_4
X_73186_ _73186_/A _86513_/Q _73186_/X sky130_fd_sc_hd__and2_4
X_70398_ _50870_/B _70364_/A _70397_/Y _83780_/D sky130_fd_sc_hd__o21ai_4
X_44105_ _44086_/A _44106_/C sky130_fd_sc_hd__buf_2
X_79802_ _79799_/X _79801_/Y _79802_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_10_967_0_CLK clkbuf_9_483_0_CLK/X _85538_/CLK sky130_fd_sc_hd__clkbuf_1
X_41317_ _41239_/X _41241_/X _41316_/X _88237_/Q _41236_/X _41317_/Y
+ sky130_fd_sc_hd__o32ai_4
X_60151_ _65198_/A _60151_/X sky130_fd_sc_hd__buf_2
X_72137_ _59325_/A _72137_/X sky130_fd_sc_hd__buf_2
X_49962_ _49981_/A _53174_/B _49962_/Y sky130_fd_sc_hd__nand2_4
X_45085_ _45052_/X _61460_/B _45070_/X _45085_/Y sky130_fd_sc_hd__o21ai_4
X_42297_ _42199_/X _42297_/X sky130_fd_sc_hd__buf_2
X_77994_ _77994_/A _77994_/B _82142_/D sky130_fd_sc_hd__xor2_4
X_48913_ _64684_/B _48896_/X _48912_/Y _48913_/Y sky130_fd_sc_hd__o21ai_4
X_44036_ _44010_/A _44036_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_9_458_0_CLK clkbuf_9_459_0_CLK/A clkbuf_9_458_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_79733_ _79733_/A _79733_/B _79739_/B sky130_fd_sc_hd__xor2_4
X_41248_ _81704_/Q _41197_/B _41248_/X sky130_fd_sc_hd__or2_4
X_60082_ _60078_/X _60079_/Y _60403_/A _72625_/B _60081_/Y _60082_/Y
+ sky130_fd_sc_hd__a41oi_4
X_72068_ _72068_/A _49106_/Y _72068_/Y sky130_fd_sc_hd__nand2_4
X_76945_ _76945_/A _81376_/D sky130_fd_sc_hd__inv_2
X_49893_ _49893_/A _49893_/B _49893_/C _53107_/D _49893_/X sky130_fd_sc_hd__and4_4
X_63910_ _63942_/A _59399_/A _63862_/C _63910_/X sky130_fd_sc_hd__and3_4
X_71019_ _53141_/B _71013_/X _71018_/Y _83633_/D sky130_fd_sc_hd__o21ai_4
X_48844_ _86472_/Q _48836_/X _48843_/Y _48844_/Y sky130_fd_sc_hd__o21ai_4
X_79664_ _79664_/A _79647_/X _79664_/X sky130_fd_sc_hd__and2_4
X_41179_ _41178_/Y _41179_/X sky130_fd_sc_hd__buf_2
X_64890_ _84223_/Q _64891_/C sky130_fd_sc_hd__inv_2
X_76876_ _76870_/Y _76910_/A _76876_/X sky130_fd_sc_hd__and2_4
X_78615_ _78616_/A _78616_/B _78614_/Y _78615_/X sky130_fd_sc_hd__o21a_4
X_63841_ _58241_/X _63858_/B _63858_/C _63793_/D _63841_/Y sky130_fd_sc_hd__nand4_4
X_75827_ _75825_/X _75827_/B _80989_/D sky130_fd_sc_hd__nand2_4
X_48775_ _52161_/A _48770_/X _48786_/C _48775_/X sky130_fd_sc_hd__and3_4
X_79595_ _79592_/Y _79594_/Y _79597_/A sky130_fd_sc_hd__nand2_4
X_45987_ _46001_/A _45987_/X sky130_fd_sc_hd__buf_2
X_47726_ _54903_/B _53209_/B sky130_fd_sc_hd__buf_2
X_66560_ _44147_/A _66560_/X sky130_fd_sc_hd__buf_2
X_78546_ _78547_/A _82674_/D _78546_/Y sky130_fd_sc_hd__nor2_4
X_44938_ _45819_/A _44939_/B sky130_fd_sc_hd__buf_2
X_63772_ _61358_/A _63772_/B _63721_/C _61012_/A _63772_/Y sky130_fd_sc_hd__nand4_4
X_75758_ _75753_/Y _75740_/B _75757_/Y _75759_/B sky130_fd_sc_hd__o21ai_4
X_60984_ _60984_/A _63738_/D sky130_fd_sc_hd__buf_2
X_65511_ _65507_/X _65663_/B _65510_/X _65511_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_905_0_CLK clkbuf_9_452_0_CLK/X _86984_/CLK sky130_fd_sc_hd__clkbuf_1
X_74709_ _74711_/A _74709_/Y sky130_fd_sc_hd__inv_2
X_62723_ _62719_/X _62721_/X _62722_/Y _62723_/Y sky130_fd_sc_hd__a21oi_4
X_47657_ _47657_/A _54867_/B sky130_fd_sc_hd__inv_2
X_66491_ _66488_/Y _66483_/X _66490_/X _84113_/D sky130_fd_sc_hd__a21o_4
X_78477_ _78465_/A _78478_/B sky130_fd_sc_hd__inv_2
X_44869_ _45387_/A _45612_/A sky130_fd_sc_hd__buf_2
X_75689_ _75689_/A _75688_/Y _75692_/A sky130_fd_sc_hd__xor2_4
X_68230_ _68188_/X _67413_/Y _68228_/X _68229_/Y _68230_/X sky130_fd_sc_hd__a211o_4
X_46608_ _46491_/A _51744_/B _46608_/Y sky130_fd_sc_hd__nand2_4
X_65442_ _65059_/X _85600_/Q _65060_/X _65441_/X _65442_/X sky130_fd_sc_hd__a211o_4
X_77428_ _77412_/A _77412_/B _77410_/Y _77428_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_5_22_0_CLK clkbuf_5_23_0_CLK/A clkbuf_6_45_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_62654_ _62651_/Y _62652_/X _62653_/Y _62654_/Y sky130_fd_sc_hd__a21oi_4
X_47588_ _47584_/Y _47555_/X _47587_/X _86619_/D sky130_fd_sc_hd__a21oi_4
X_49327_ _48995_/A _49327_/X sky130_fd_sc_hd__buf_2
X_61605_ _61634_/A _61634_/B _79135_/B _61605_/Y sky130_fd_sc_hd__nor3_4
X_68161_ _67010_/X _67012_/X _68129_/X _68161_/Y sky130_fd_sc_hd__a21oi_4
X_46539_ _46539_/A _50854_/B sky130_fd_sc_hd__buf_2
X_65373_ _65397_/A _65397_/B _65373_/C _65373_/Y sky130_fd_sc_hd__nor3_4
X_77359_ _77359_/A _77360_/A sky130_fd_sc_hd__inv_2
X_62585_ _62487_/X _58198_/A _62618_/C _62608_/D _62585_/X sky130_fd_sc_hd__and4_4
X_67112_ _88381_/Q _67110_/X _67040_/X _67111_/X _67112_/X sky130_fd_sc_hd__a211o_4
X_64324_ _64336_/A _84824_/Q _64323_/X _64324_/Y sky130_fd_sc_hd__nand3_4
X_49258_ _86423_/Q _49255_/X _49257_/Y _49258_/Y sky130_fd_sc_hd__o21ai_4
X_61536_ _61546_/A _61546_/B _79141_/B _61536_/Y sky130_fd_sc_hd__nor3_4
X_80370_ _84753_/Q _84145_/Q _80370_/X sky130_fd_sc_hd__xor2_4
X_68092_ _82081_/D _68040_/X _68091_/X _68092_/X sky130_fd_sc_hd__a21bo_4
Xclkbuf_10_9_0_CLK clkbuf_9_4_0_CLK/X _85277_/CLK sky130_fd_sc_hd__clkbuf_1
X_48209_ _48206_/Y _48175_/X _48208_/Y _86556_/D sky130_fd_sc_hd__a21boi_4
X_67043_ _67038_/X _67042_/X _67015_/X _67043_/Y sky130_fd_sc_hd__a21oi_4
X_79029_ _82651_/Q _79029_/Y sky130_fd_sc_hd__inv_2
X_64255_ _64314_/A _64255_/X sky130_fd_sc_hd__buf_2
X_61467_ _72529_/C _61467_/X sky130_fd_sc_hd__buf_2
X_49189_ _49405_/A _49189_/X sky130_fd_sc_hd__buf_2
X_51220_ _51220_/A _51203_/B _51197_/C _51220_/D _51220_/X sky130_fd_sc_hd__and4_4
X_63206_ _63157_/X _63206_/B _63241_/C _63181_/X _63206_/X sky130_fd_sc_hd__and4_4
X_82040_ _82009_/CLK _77934_/B _82040_/Q sky130_fd_sc_hd__dfxtp_4
X_60418_ _60155_/C _60407_/A _60403_/B _60418_/D _60502_/A sky130_fd_sc_hd__and4_4
X_64186_ _63912_/X _64186_/X sky130_fd_sc_hd__buf_2
X_61398_ _61375_/A _61398_/B _61398_/C _61398_/Y sky130_fd_sc_hd__nand3_4
X_51151_ _51145_/Y _51147_/X _51150_/X _51151_/Y sky130_fd_sc_hd__a21oi_4
X_63137_ _63100_/A _63137_/B _63147_/C _63124_/D _63137_/X sky130_fd_sc_hd__and4_4
X_60349_ _64939_/A _60349_/X sky130_fd_sc_hd__buf_2
X_68994_ _68994_/A _88346_/Q _68994_/X sky130_fd_sc_hd__and2_4
X_50102_ _50100_/Y _50092_/X _50101_/X _50102_/Y sky130_fd_sc_hd__a21oi_4
X_51082_ _50946_/A _51191_/A sky130_fd_sc_hd__buf_2
X_67945_ _67941_/X _67944_/X _67897_/X _67945_/Y sky130_fd_sc_hd__a21oi_4
X_63068_ _63061_/Y _63063_/X _63064_/X _63066_/X _63067_/X _63068_/Y
+ sky130_fd_sc_hd__o41ai_4
X_83991_ _82896_/CLK _83991_/D _82639_/D sky130_fd_sc_hd__dfxtp_4
X_50033_ _50027_/A _53246_/B _50033_/Y sky130_fd_sc_hd__nand2_4
X_54910_ _54910_/A _54910_/B _54910_/C _53217_/D _54910_/X sky130_fd_sc_hd__and4_4
X_85730_ _83690_/CLK _52923_/Y _85730_/Q sky130_fd_sc_hd__dfxtp_4
X_62019_ _59765_/A _62021_/B sky130_fd_sc_hd__buf_2
X_82942_ _82942_/CLK _78101_/X _46285_/A sky130_fd_sc_hd__dfxtp_4
X_55890_ _45081_/A _55617_/A _44099_/X _55889_/X _55890_/X sky130_fd_sc_hd__a211o_4
X_67876_ _67871_/X _67874_/X _67875_/X _67876_/Y sky130_fd_sc_hd__a21oi_4
X_69615_ _69186_/Y _69603_/X _69604_/X _69614_/Y _69615_/X sky130_fd_sc_hd__a211o_4
X_54841_ _54850_/A _47610_/A _54841_/Y sky130_fd_sc_hd__nand2_4
X_66827_ _80919_/D _66734_/X _66826_/X _66827_/X sky130_fd_sc_hd__a21bo_4
X_85661_ _85436_/CLK _53289_/Y _85661_/Q sky130_fd_sc_hd__dfxtp_4
X_82873_ _82942_/CLK _78241_/B _82873_/Q sky130_fd_sc_hd__dfxtp_4
X_87400_ _87653_/CLK _43482_/X _87400_/Q sky130_fd_sc_hd__dfxtp_4
X_84612_ _84469_/CLK _84612_/D _79152_/A sky130_fd_sc_hd__dfxtp_4
X_81824_ _83761_/CLK _81632_/Q _81824_/Q sky130_fd_sc_hd__dfxtp_4
X_57560_ _57597_/A _48257_/B _57560_/Y sky130_fd_sc_hd__nand2_4
X_69546_ _69543_/X _69545_/X _64629_/A _69546_/X sky130_fd_sc_hd__a21o_4
X_88380_ _87865_/CLK _88380_/D _88380_/Q sky130_fd_sc_hd__dfxtp_4
X_54772_ _54758_/X _54772_/B _54772_/Y sky130_fd_sc_hd__nand2_4
X_85592_ _85590_/CLK _53668_/Y _85592_/Q sky130_fd_sc_hd__dfxtp_4
X_66758_ _68386_/A _66758_/X sky130_fd_sc_hd__buf_2
X_51984_ _51980_/Y _51981_/X _51983_/Y _51984_/Y sky130_fd_sc_hd__a21boi_4
X_56511_ _56099_/X _56499_/X _56510_/Y _85168_/D sky130_fd_sc_hd__o21ai_4
X_87331_ _87045_/CLK _43640_/X _87331_/Q sky130_fd_sc_hd__dfxtp_4
X_53723_ _53723_/A _53791_/A sky130_fd_sc_hd__buf_2
X_65709_ _65596_/X _83063_/Q _65707_/X _65708_/X _65710_/B sky130_fd_sc_hd__a211o_4
X_84543_ _84529_/CLK _84543_/D _84543_/Q sky130_fd_sc_hd__dfxtp_4
X_50935_ _50933_/Y _50928_/X _50934_/X _50935_/Y sky130_fd_sc_hd__a21oi_4
X_57491_ _57491_/A _57491_/B _57491_/C _57491_/Y sky130_fd_sc_hd__nor3_4
X_81755_ _81755_/CLK _76104_/B _41314_/A sky130_fd_sc_hd__dfxtp_4
X_69477_ _81385_/D _69439_/X _69476_/X _83921_/D sky130_fd_sc_hd__a21bo_4
X_66689_ _66689_/A _66689_/B _66689_/X sky130_fd_sc_hd__and2_4
X_59230_ _72358_/A _59230_/X sky130_fd_sc_hd__buf_2
X_56442_ _56446_/A _56446_/B _56442_/C _56442_/Y sky130_fd_sc_hd__nand3_4
X_68428_ _87505_/Q _68365_/X _68053_/X _68427_/X _68428_/X sky130_fd_sc_hd__a211o_4
X_80706_ _81104_/CLK _75892_/X _80674_/D sky130_fd_sc_hd__dfxtp_4
X_87262_ _87776_/CLK _43799_/Y _69427_/B sky130_fd_sc_hd__dfxtp_4
X_53654_ _52135_/A _53658_/B _53667_/C _53654_/X sky130_fd_sc_hd__and3_4
X_84474_ _82822_/CLK _61519_/Y _79142_/B sky130_fd_sc_hd__dfxtp_4
X_50866_ _50857_/X _51378_/B _50866_/Y sky130_fd_sc_hd__nand2_4
X_81686_ _81257_/CLK _81686_/D _81686_/Q sky130_fd_sc_hd__dfxtp_4
X_86213_ _86213_/CLK _50377_/Y _86213_/Q sky130_fd_sc_hd__dfxtp_4
X_52605_ _52605_/A _52605_/X sky130_fd_sc_hd__buf_2
X_59161_ _59160_/X _85652_/Q _59081_/X _59161_/X sky130_fd_sc_hd__o21a_4
X_83425_ _82386_/CLK _83425_/D _83425_/Q sky130_fd_sc_hd__dfxtp_4
X_56373_ _56370_/Y _56435_/A sky130_fd_sc_hd__buf_2
X_80637_ _46128_/D _46158_/B _80651_/D sky130_fd_sc_hd__nand2_4
X_68359_ _68651_/A _68359_/X sky130_fd_sc_hd__buf_2
X_87193_ _87189_/CLK _87193_/D _67955_/B sky130_fd_sc_hd__dfxtp_4
X_53585_ _53661_/A _53846_/A sky130_fd_sc_hd__buf_2
XPHY_103 sky130_fd_sc_hd__decap_3
X_50797_ _50787_/X _46417_/B _50797_/Y sky130_fd_sc_hd__nand2_4
XPHY_114 sky130_fd_sc_hd__decap_3
X_58112_ _58796_/A _58112_/X sky130_fd_sc_hd__buf_2
XPHY_125 sky130_fd_sc_hd__decap_3
X_55324_ _82990_/Q _55311_/X _55312_/X _55323_/X _55324_/X sky130_fd_sc_hd__a211o_4
X_86144_ _85535_/CLK _50737_/Y _86144_/Q sky130_fd_sc_hd__dfxtp_4
X_40550_ _44733_/A _40550_/X sky130_fd_sc_hd__buf_2
X_52536_ _65209_/B _52500_/X _52535_/Y _52536_/Y sky130_fd_sc_hd__o21ai_4
XPHY_136 sky130_fd_sc_hd__decap_3
X_59092_ _59078_/Y _58857_/X _59088_/X _59091_/X _59092_/Y sky130_fd_sc_hd__a22oi_4
X_71370_ _71344_/A _83522_/Q _71369_/X _71370_/X sky130_fd_sc_hd__a21o_4
X_83356_ _83414_/CLK _83356_/D _83356_/Q sky130_fd_sc_hd__dfxtp_4
X_80568_ _80568_/A _80568_/B _80569_/B sky130_fd_sc_hd__xor2_4
XPHY_147 sky130_fd_sc_hd__decap_3
XPHY_158 sky130_fd_sc_hd__decap_3
XPHY_169 sky130_fd_sc_hd__decap_3
X_58043_ _58618_/A _58043_/X sky130_fd_sc_hd__buf_2
X_70321_ _70328_/A _70328_/B _70321_/C _70328_/D _70321_/X sky130_fd_sc_hd__and4_4
X_82307_ _80835_/CLK _77006_/Y _82307_/Q sky130_fd_sc_hd__dfxtp_4
X_55255_ _55254_/A _55253_/X _83320_/Q _55678_/A sky130_fd_sc_hd__a21o_4
X_86075_ _85754_/CLK _86075_/D _86075_/Q sky130_fd_sc_hd__dfxtp_4
X_40481_ _40477_/X _40443_/X _40480_/X _88385_/Q _40447_/X _40481_/Y
+ sky130_fd_sc_hd__o32ai_4
X_52467_ _85816_/Q _52438_/X _52466_/Y _52467_/Y sky130_fd_sc_hd__o21ai_4
X_83287_ _85542_/CLK _83287_/D _83287_/Q sky130_fd_sc_hd__dfxtp_4
X_80499_ _80495_/X _80498_/Y _80502_/A sky130_fd_sc_hd__xor2_4
Xclkbuf_7_120_0_CLK clkbuf_6_60_0_CLK/X clkbuf_8_241_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_42220_ _41361_/X _42209_/X _87973_/Q _42210_/X _87973_/D sky130_fd_sc_hd__a2bb2o_4
X_54206_ _85484_/Q _54193_/X _54205_/Y _54206_/Y sky130_fd_sc_hd__o21ai_4
X_73040_ _73040_/A _73040_/B _73040_/X sky130_fd_sc_hd__and2_4
X_85026_ _85100_/CLK _57370_/X _85026_/Q sky130_fd_sc_hd__dfxtp_4
X_51418_ _51403_/X _52944_/B _51418_/Y sky130_fd_sc_hd__nand2_4
X_70252_ _70238_/X _74790_/B _70251_/X _70252_/X sky130_fd_sc_hd__a21o_4
X_82238_ _82515_/CLK _82270_/Q _82238_/Q sky130_fd_sc_hd__dfxtp_4
X_55186_ _55174_/X _55186_/B _55186_/Y sky130_fd_sc_hd__nor2_4
X_52398_ _52398_/A _52630_/A sky130_fd_sc_hd__buf_2
Xclkbuf_2_3_1_CLK clkbuf_2_3_0_CLK/X clkbuf_2_3_1_CLK/X sky130_fd_sc_hd__clkbuf_1
X_42151_ _41161_/X _42148_/X _88010_/Q _42150_/X _42151_/X sky130_fd_sc_hd__a2bb2o_4
X_54137_ _54127_/X _54160_/B _54118_/X _52971_/D _54137_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_90_0_CLK clkbuf_9_45_0_CLK/X _84403_/CLK sky130_fd_sc_hd__clkbuf_1
X_51349_ _51346_/Y _51339_/X _51348_/X _51349_/Y sky130_fd_sc_hd__a21oi_4
X_70183_ _70183_/A _70183_/B _70183_/C _70183_/D _70183_/X sky130_fd_sc_hd__and4_4
X_82169_ _82047_/CLK _84161_/Q _77942_/A sky130_fd_sc_hd__dfxtp_4
X_59994_ _66064_/A _60543_/B sky130_fd_sc_hd__buf_2
X_41102_ _82275_/Q _41102_/B _41102_/X sky130_fd_sc_hd__or2_4
X_42082_ _43161_/A _42083_/A sky130_fd_sc_hd__buf_2
X_58945_ _79180_/A _58857_/X _58940_/X _58944_/X _58945_/Y sky130_fd_sc_hd__a22oi_4
X_54068_ _53990_/A _54068_/X sky130_fd_sc_hd__buf_2
X_74991_ _74988_/Y _74990_/X _75001_/A sky130_fd_sc_hd__nand2_4
X_86977_ _88363_/CLK _86977_/D _44747_/A sky130_fd_sc_hd__dfxtp_4
X_45910_ _45893_/B _86770_/Q _45909_/X _86844_/D sky130_fd_sc_hd__a21o_4
X_41033_ _41032_/X _40987_/X _69376_/B _40989_/X _88290_/D sky130_fd_sc_hd__a2bb2o_4
X_53019_ _53019_/A _53036_/B _53019_/C _53019_/D _53019_/X sky130_fd_sc_hd__and4_4
X_76730_ _76714_/Y _76715_/Y _76730_/Y sky130_fd_sc_hd__nor2_4
X_73942_ _87331_/Q _74246_/B _73942_/Y sky130_fd_sc_hd__nor2_4
X_85928_ _86089_/CLK _51888_/Y _85928_/Q sky130_fd_sc_hd__dfxtp_4
X_46890_ _46653_/A _47081_/A sky130_fd_sc_hd__buf_2
X_58876_ _58876_/A _58877_/A sky130_fd_sc_hd__buf_2
X_45841_ _55231_/B _45394_/X _45396_/X _45840_/Y _45841_/X sky130_fd_sc_hd__a211o_4
X_57827_ _57739_/X _85723_/Q _57814_/X _57827_/X sky130_fd_sc_hd__o21a_4
X_76661_ _76661_/A _76663_/A sky130_fd_sc_hd__inv_2
X_73873_ _73873_/A _73873_/B _73873_/Y sky130_fd_sc_hd__nor2_4
X_85859_ _85859_/CLK _85859_/D _85859_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_251_0_CLK clkbuf_8_251_0_CLK/A clkbuf_9_502_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_78400_ _78400_/A _78400_/B _82760_/D sky130_fd_sc_hd__xor2_4
X_75612_ _81111_/Q _75612_/B _80775_/D sky130_fd_sc_hd__xor2_4
X_48560_ _48559_/Y _48561_/B sky130_fd_sc_hd__buf_2
X_72824_ _83175_/Q _72794_/X _72823_/Y _83175_/D sky130_fd_sc_hd__a21o_4
X_79380_ _79358_/Y _79376_/X _79379_/Y _79381_/B sky130_fd_sc_hd__a21oi_4
X_45772_ _85033_/Q _44933_/X _45771_/X _45772_/Y sky130_fd_sc_hd__o21ai_4
X_57758_ _58857_/A _57758_/X sky130_fd_sc_hd__buf_2
X_76592_ _81374_/Q _76591_/X _76592_/X sky130_fd_sc_hd__xor2_4
X_42984_ _43774_/A _42984_/X sky130_fd_sc_hd__buf_2
X_47511_ _81795_/Q _47511_/Y sky130_fd_sc_hd__inv_2
X_78331_ _78329_/Y _78331_/B _78332_/A _78337_/C sky130_fd_sc_hd__nand3_4
X_44723_ _44712_/X _44713_/X _40707_/X _86986_/Q _44714_/X _44723_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56709_ _57284_/A _57416_/A sky130_fd_sc_hd__buf_2
X_75543_ _75543_/A _75543_/B _75543_/X sky130_fd_sc_hd__xor2_4
X_41935_ _42081_/A _41936_/A sky130_fd_sc_hd__buf_2
X_87529_ _87533_/CLK _43225_/X _87529_/Q sky130_fd_sc_hd__dfxtp_4
X_48491_ _83581_/Q _53678_/B sky130_fd_sc_hd__inv_2
X_72755_ _73359_/A _72755_/X sky130_fd_sc_hd__buf_2
X_57689_ _57689_/A _58094_/A sky130_fd_sc_hd__buf_2
X_47442_ _83730_/Q _47442_/Y sky130_fd_sc_hd__inv_2
X_71706_ _71706_/A _71637_/C _71777_/B _71706_/Y sky130_fd_sc_hd__nand3_4
X_59428_ _58548_/A _83344_/Q _59428_/Y sky130_fd_sc_hd__nor2_4
X_78262_ _78262_/A _78262_/B _78262_/X sky130_fd_sc_hd__xor2_4
X_44654_ _44638_/X _44639_/X _41076_/A _87014_/Q _44640_/X _44655_/A
+ sky130_fd_sc_hd__o32ai_4
X_75474_ _75475_/A _75475_/B _75477_/B sky130_fd_sc_hd__nor2_4
X_41866_ _41877_/A _42429_/A sky130_fd_sc_hd__buf_2
X_72686_ _72686_/A _72686_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_261_0_CLK clkbuf_9_130_0_CLK/X _83480_/CLK sky130_fd_sc_hd__clkbuf_1
X_77213_ _77213_/A _77212_/Y _77214_/B sky130_fd_sc_hd__xor2_4
X_43605_ _43605_/A _43606_/A sky130_fd_sc_hd__buf_2
X_74425_ _74458_/A _74425_/X sky130_fd_sc_hd__buf_2
X_40817_ _40817_/A _40817_/X sky130_fd_sc_hd__buf_2
X_47373_ _47372_/Y _53012_/B sky130_fd_sc_hd__buf_2
X_59359_ _59356_/Y _59358_/Y _59297_/X _59359_/X sky130_fd_sc_hd__a21o_4
X_71637_ _71637_/A _71226_/B _71637_/C _71637_/Y sky130_fd_sc_hd__nand3_4
XPHY_5 sky130_fd_sc_hd__decap_3
X_78193_ _78191_/B _78193_/B _78174_/B _78193_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_891_0_CLK clkbuf_9_445_0_CLK/X _86145_/CLK sky130_fd_sc_hd__clkbuf_1
X_44585_ _44565_/X _44567_/X _40909_/X _87044_/Q _44568_/X _44586_/A
+ sky130_fd_sc_hd__o32ai_4
X_41797_ _41796_/Y _41797_/X sky130_fd_sc_hd__buf_2
X_49112_ _49112_/A _50677_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_43_0_CLK clkbuf_9_21_0_CLK/X _83843_/CLK sky130_fd_sc_hd__clkbuf_1
X_46324_ _83651_/Q _53971_/B sky130_fd_sc_hd__inv_2
X_77144_ _77143_/Y _77141_/C _77144_/X sky130_fd_sc_hd__and2_4
X_43536_ _40408_/X _43532_/X _87371_/Q _43533_/X _87371_/D sky130_fd_sc_hd__a2bb2o_4
X_62370_ _62368_/Y _62327_/X _62369_/Y _84415_/D sky130_fd_sc_hd__a21oi_4
X_74356_ _83085_/Q _72699_/X _74355_/Y _74356_/X sky130_fd_sc_hd__a21bo_4
X_40748_ _40628_/X _81124_/Q _40747_/X _40748_/Y sky130_fd_sc_hd__o21ai_4
X_71568_ _70558_/X _71583_/B _71558_/X _71568_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_9_382_0_CLK clkbuf_9_382_0_CLK/A clkbuf_9_382_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_61321_ _72507_/A _61317_/A _61313_/A _61321_/Y sky130_fd_sc_hd__nand3_4
X_49043_ _49037_/Y _49038_/X _49042_/X _86450_/D sky130_fd_sc_hd__a21oi_4
X_73307_ _73426_/A _86476_/Q _73307_/X sky130_fd_sc_hd__and2_4
X_46255_ _53946_/B _49212_/B sky130_fd_sc_hd__buf_2
X_70519_ _57668_/Y _70501_/X _70518_/Y _70519_/Y sky130_fd_sc_hd__o21ai_4
XPHY_670 sky130_fd_sc_hd__decap_3
X_77075_ _81997_/Q _82285_/D _77077_/A sky130_fd_sc_hd__or2_4
X_43467_ _43466_/X _43467_/X sky130_fd_sc_hd__buf_2
X_74287_ _83112_/Q _72702_/X _74286_/Y _83112_/D sky130_fd_sc_hd__a21bo_4
XPHY_681 sky130_fd_sc_hd__decap_3
Xclkbuf_10_276_0_CLK clkbuf_9_138_0_CLK/X _85407_/CLK sky130_fd_sc_hd__clkbuf_1
X_40679_ _40678_/X _40651_/X _88355_/Q _40652_/X _88355_/D sky130_fd_sc_hd__a2bb2o_4
X_71499_ _71487_/X _83477_/Q _71498_/X _83477_/D sky130_fd_sc_hd__a21o_4
XPHY_692 sky130_fd_sc_hd__decap_3
X_45206_ _45281_/A _45206_/X sky130_fd_sc_hd__buf_2
X_64040_ _63227_/B _64118_/B _64040_/C _64142_/D _64040_/Y sky130_fd_sc_hd__nand4_4
X_76026_ _81713_/D _76027_/B _76028_/A sky130_fd_sc_hd__or2_4
X_42418_ _42417_/X _42410_/X _40474_/X _87874_/Q _42411_/X _42419_/A
+ sky130_fd_sc_hd__o32ai_4
X_61252_ _72590_/A _61252_/X sky130_fd_sc_hd__buf_2
X_73238_ _73238_/A _73238_/X sky130_fd_sc_hd__buf_2
X_46186_ _46186_/A _46125_/A _46186_/X sky130_fd_sc_hd__or2_4
X_43398_ _41469_/X _43396_/X _87441_/Q _43397_/X _87441_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_10_58_0_CLK clkbuf_9_29_0_CLK/X _85040_/CLK sky130_fd_sc_hd__clkbuf_1
X_60203_ _62737_/A _60218_/A sky130_fd_sc_hd__buf_2
X_45137_ _45212_/A _45137_/X sky130_fd_sc_hd__buf_2
X_42349_ _42348_/Y _87909_/D sky130_fd_sc_hd__inv_2
X_61183_ _61183_/A _61177_/Y _61178_/Y _61182_/X _61183_/Y sky130_fd_sc_hd__nor4_4
X_73169_ _74437_/B _73169_/B _73169_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_9_397_0_CLK clkbuf_8_198_0_CLK/X clkbuf_9_397_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_8_204_0_CLK clkbuf_8_205_0_CLK/A clkbuf_9_409_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_60134_ _84656_/Q _60132_/X _60133_/Y _60015_/Y _60134_/X sky130_fd_sc_hd__a2bb2o_4
X_49945_ _49955_/A _53157_/B _49945_/Y sky130_fd_sc_hd__nand2_4
X_45068_ _45065_/X _45067_/Y _45049_/X _45068_/Y sky130_fd_sc_hd__a21oi_4
X_65991_ _65486_/A _65992_/A sky130_fd_sc_hd__buf_2
X_77977_ _77977_/A _77977_/Y sky130_fd_sc_hd__inv_2
X_44019_ _44019_/A _44020_/A sky130_fd_sc_hd__buf_2
X_67730_ _87459_/Q _67628_/X _67702_/X _67729_/X _67730_/X sky130_fd_sc_hd__a211o_4
X_79716_ _79702_/A _79701_/Y _79716_/X sky130_fd_sc_hd__or2_4
X_64942_ _65047_/A _64870_/B _64942_/C _64942_/Y sky130_fd_sc_hd__nor3_4
X_60065_ _59951_/D _60061_/Y _60063_/Y _60129_/B _60064_/Y _84668_/D
+ sky130_fd_sc_hd__a41oi_4
X_76928_ _76928_/A _76927_/Y _81567_/D sky130_fd_sc_hd__nand2_4
X_49876_ _49794_/X _49893_/C sky130_fd_sc_hd__buf_2
Xclkbuf_9_320_0_CLK clkbuf_8_160_0_CLK/X clkbuf_9_320_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_48827_ _47918_/A _48853_/A sky130_fd_sc_hd__buf_2
X_67661_ _67656_/X _67660_/X _67637_/X _67661_/Y sky130_fd_sc_hd__a21oi_4
X_79647_ _65221_/C _72394_/Y _79646_/Y _79647_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_8_219_0_CLK clkbuf_8_219_0_CLK/A clkbuf_9_438_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_64873_ _64817_/X _86135_/Q _64776_/X _64872_/X _64873_/X sky130_fd_sc_hd__a211o_4
X_76859_ _76847_/Y _81368_/D sky130_fd_sc_hd__inv_2
Xclkbuf_10_214_0_CLK clkbuf_9_107_0_CLK/X _84623_/CLK sky130_fd_sc_hd__clkbuf_1
X_69400_ _69395_/X _69398_/X _69399_/X _69400_/X sky130_fd_sc_hd__a21o_4
X_66612_ _66526_/X _66597_/Y _59782_/X _66611_/Y _66612_/X sky130_fd_sc_hd__a211o_4
X_63824_ _60882_/X _63860_/C sky130_fd_sc_hd__buf_2
Xclkbuf_10_844_0_CLK clkbuf_9_422_0_CLK/X _82748_/CLK sky130_fd_sc_hd__clkbuf_1
X_48758_ _73012_/B _48754_/X _48757_/Y _48758_/Y sky130_fd_sc_hd__o21ai_4
X_67592_ _67569_/X _87720_/Q _67592_/X sky130_fd_sc_hd__and2_4
X_79578_ _79575_/Y _79578_/B _79580_/A sky130_fd_sc_hd__nand2_4
X_69331_ _88037_/Q _69121_/X _69232_/X _69330_/X _69331_/X sky130_fd_sc_hd__a211o_4
X_47709_ _81230_/Q _47710_/A sky130_fd_sc_hd__inv_2
X_66543_ _68614_/A _68999_/A sky130_fd_sc_hd__buf_2
X_78529_ _78521_/X _78528_/X _78529_/Y sky130_fd_sc_hd__xnor2_4
X_63755_ _60879_/D _64045_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_335_0_CLK clkbuf_9_335_0_CLK/A clkbuf_9_335_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_60967_ _60967_/A _60967_/X sky130_fd_sc_hd__buf_2
X_48689_ _74505_/A _48691_/A sky130_fd_sc_hd__buf_2
X_50720_ _50717_/Y _50699_/X _50719_/Y _86147_/D sky130_fd_sc_hd__a21boi_4
X_62706_ _62673_/A _62673_/B _84389_/Q _62706_/Y sky130_fd_sc_hd__nor3_4
X_81540_ _83940_/CLK _81540_/D _81528_/D sky130_fd_sc_hd__dfxtp_4
X_69262_ _69179_/A _69262_/B _69262_/X sky130_fd_sc_hd__and2_4
X_66474_ _66472_/Y _66449_/X _66473_/X _84116_/D sky130_fd_sc_hd__a21o_4
Xclkbuf_10_229_0_CLK clkbuf_9_114_0_CLK/X _84438_/CLK sky130_fd_sc_hd__clkbuf_1
X_63686_ _61663_/B _63609_/X _63684_/X _63685_/X _63686_/X sky130_fd_sc_hd__a211o_4
X_60898_ _60341_/A _60898_/X sky130_fd_sc_hd__buf_2
X_68213_ _67323_/X _67325_/X _68209_/X _68213_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_859_0_CLK clkbuf_9_429_0_CLK/X _86122_/CLK sky130_fd_sc_hd__clkbuf_1
X_65425_ _65403_/A _65425_/B _65425_/X sky130_fd_sc_hd__and2_4
X_50651_ _50496_/A _50651_/X sky130_fd_sc_hd__buf_2
X_62637_ _62635_/Y _62593_/X _62636_/Y _84394_/D sky130_fd_sc_hd__a21oi_4
X_81471_ _81482_/CLK _81471_/D _81471_/Q sky130_fd_sc_hd__dfxtp_4
X_69193_ _69179_/A _87279_/Q _69193_/X sky130_fd_sc_hd__and2_4
X_83210_ _83231_/CLK _72629_/Y _79160_/B sky130_fd_sc_hd__dfxtp_4
X_80422_ _80422_/A _80422_/B _80423_/B sky130_fd_sc_hd__xor2_4
X_68144_ _67495_/X _68144_/X sky130_fd_sc_hd__buf_2
X_53370_ _85646_/Q _53351_/X _53369_/Y _53370_/Y sky130_fd_sc_hd__o21ai_4
X_65356_ _65353_/X _65355_/X _65277_/X _65359_/A sky130_fd_sc_hd__a21o_4
X_84190_ _83520_/CLK _65606_/X _84190_/Q sky130_fd_sc_hd__dfxtp_4
X_50582_ _50607_/A _48922_/B _50582_/Y sky130_fd_sc_hd__nand2_4
X_62568_ _61629_/B _62504_/X _62534_/X _62475_/X _62569_/D sky130_fd_sc_hd__nand4_4
X_52321_ _52318_/Y _52314_/X _52320_/X _52321_/Y sky130_fd_sc_hd__a21oi_4
X_64307_ _64295_/A _64307_/B _64307_/C _64307_/X sky130_fd_sc_hd__and3_4
X_83141_ _83141_/CLK _73673_/Y _70123_/A sky130_fd_sc_hd__dfxtp_4
X_80353_ _80353_/A _80353_/B _80353_/Y sky130_fd_sc_hd__nand2_4
X_61519_ _61516_/X _61517_/X _61518_/Y _61519_/Y sky130_fd_sc_hd__a21oi_4
X_68075_ _68444_/A _88212_/Q _68075_/X sky130_fd_sc_hd__and2_4
X_65287_ _64807_/A _65287_/X sky130_fd_sc_hd__buf_2
X_62499_ _62497_/Y _62467_/X _62498_/Y _84406_/D sky130_fd_sc_hd__a21oi_4
X_55040_ _55038_/Y _55024_/X _55039_/X _85330_/D sky130_fd_sc_hd__a21oi_4
X_67026_ _67025_/X _67026_/X sky130_fd_sc_hd__buf_2
X_52252_ _52198_/A _52267_/B sky130_fd_sc_hd__buf_2
X_64238_ _59456_/Y _64226_/X _64237_/Y _64238_/Y sky130_fd_sc_hd__o21ai_4
X_83072_ _83584_/CLK _74411_/Y _83072_/Q sky130_fd_sc_hd__dfxtp_4
X_80284_ _80280_/B _80280_/C _80284_/Y sky130_fd_sc_hd__nand2_4
X_51203_ _51191_/X _51203_/B _51197_/C _52895_/D _51203_/X sky130_fd_sc_hd__and4_4
X_86900_ _86900_/CLK _45086_/Y _64343_/B sky130_fd_sc_hd__dfxtp_4
X_82023_ _81990_/CLK _77774_/B _81991_/D sky130_fd_sc_hd__dfxtp_4
X_52183_ _52181_/Y _52170_/X _52182_/X _85873_/D sky130_fd_sc_hd__a21oi_4
X_64169_ _58207_/A _64192_/C _64180_/C _64192_/D _64169_/Y sky130_fd_sc_hd__nand4_4
X_87880_ _87883_/CLK _42403_/Y _87880_/Q sky130_fd_sc_hd__dfxtp_4
X_51134_ _51130_/A _52829_/B _51134_/Y sky130_fd_sc_hd__nand2_4
X_86831_ _87990_/CLK _45977_/X _86831_/Q sky130_fd_sc_hd__dfxtp_4
X_56991_ _56985_/D _56991_/Y sky130_fd_sc_hd__inv_2
X_68977_ _69021_/A _68977_/B _68977_/X sky130_fd_sc_hd__and2_4
X_58730_ _58605_/A _58730_/X sky130_fd_sc_hd__buf_2
X_51065_ _51039_/A _51065_/X sky130_fd_sc_hd__buf_2
X_55942_ _55939_/X _55941_/X _55615_/A _55945_/A sky130_fd_sc_hd__a21o_4
X_67928_ _87898_/Q _67831_/X _67879_/X _67927_/X _67928_/X sky130_fd_sc_hd__a211o_4
X_86762_ _80672_/CLK _86762_/D _86762_/Q sky130_fd_sc_hd__dfxtp_4
X_83974_ _83974_/CLK _83974_/D _83974_/Q sky130_fd_sc_hd__dfxtp_4
X_50016_ _50025_/A _49994_/X _50025_/C _53230_/D _50016_/X sky130_fd_sc_hd__and4_4
X_85713_ _84766_/CLK _53016_/Y _85713_/Q sky130_fd_sc_hd__dfxtp_4
X_58661_ _58631_/X _58659_/Y _58660_/Y _58650_/X _58636_/X _58661_/X
+ sky130_fd_sc_hd__o32a_4
X_82925_ _82925_/CLK _78211_/X _82925_/Q sky130_fd_sc_hd__dfxtp_4
X_55873_ _55873_/A _56073_/A sky130_fd_sc_hd__buf_2
X_67859_ _67854_/X _67857_/X _67858_/X _67859_/X sky130_fd_sc_hd__a21o_4
X_86693_ _86695_/CLK _86693_/D _58921_/A sky130_fd_sc_hd__dfxtp_4
X_57612_ _84969_/Q _57603_/X _57611_/Y _57612_/Y sky130_fd_sc_hd__o21ai_4
X_54824_ _85371_/Q _54812_/X _54823_/Y _54824_/Y sky130_fd_sc_hd__o21ai_4
X_85644_ _85738_/CLK _53385_/Y _85644_/Q sky130_fd_sc_hd__dfxtp_4
X_70870_ _51807_/B _70855_/X _70869_/Y _70870_/Y sky130_fd_sc_hd__o21ai_4
X_58592_ _58100_/X _85951_/Q _58568_/X _58592_/X sky130_fd_sc_hd__o21a_4
X_82856_ _82855_/CLK _78125_/B _40897_/A sky130_fd_sc_hd__dfxtp_4
X_57543_ _46399_/A _57543_/X sky130_fd_sc_hd__buf_2
X_81807_ _81807_/CLK _81807_/D _81807_/Q sky130_fd_sc_hd__dfxtp_4
X_69529_ _69520_/X _69050_/Y _69516_/X _69528_/Y _69529_/X sky130_fd_sc_hd__a211o_4
X_88363_ _88363_/CLK _88363_/D _88363_/Q sky130_fd_sc_hd__dfxtp_4
X_54755_ _54775_/A _54755_/B _54775_/C _47465_/A _54755_/X sky130_fd_sc_hd__and4_4
X_85575_ _86500_/CLK _53753_/Y _85575_/Q sky130_fd_sc_hd__dfxtp_4
X_51967_ _73707_/B _51960_/X _51966_/Y _51967_/Y sky130_fd_sc_hd__o21ai_4
X_82787_ _83238_/CLK _82787_/D _78318_/B sky130_fd_sc_hd__dfxtp_4
X_87314_ _83153_/CLK _43679_/X _87314_/Q sky130_fd_sc_hd__dfxtp_4
X_41720_ _41717_/X _41374_/A _41719_/X _41720_/Y sky130_fd_sc_hd__o21ai_4
X_53706_ _85584_/Q _53610_/X _53705_/Y _53706_/Y sky130_fd_sc_hd__o21ai_4
X_84526_ _84400_/CLK _61056_/X _61055_/C sky130_fd_sc_hd__dfxtp_4
X_72540_ _61295_/A _72540_/B _72510_/C _72540_/Y sky130_fd_sc_hd__nor3_4
X_50918_ _50918_/A _50941_/A sky130_fd_sc_hd__buf_2
X_81738_ _81783_/CLK _75982_/B _41406_/A sky130_fd_sc_hd__dfxtp_4
X_57474_ _74831_/A _56971_/B _57473_/Y _57474_/Y sky130_fd_sc_hd__o21ai_4
X_88294_ _87253_/CLK _41011_/Y _88294_/Q sky130_fd_sc_hd__dfxtp_4
X_54686_ _54683_/Y _54666_/X _54685_/X _54686_/Y sky130_fd_sc_hd__a21oi_4
X_51898_ _51887_/A _51898_/B _51893_/C _52724_/D _51898_/X sky130_fd_sc_hd__and4_4
X_59213_ _86672_/Q _59189_/B _59213_/Y sky130_fd_sc_hd__nor2_4
X_56425_ _56103_/X _56409_/X _56424_/Y _85199_/D sky130_fd_sc_hd__o21ai_4
X_41651_ _41651_/A _41651_/X sky130_fd_sc_hd__buf_2
X_87245_ _87766_/CLK _87245_/D _68530_/B sky130_fd_sc_hd__dfxtp_4
X_53637_ _53634_/Y _53619_/X _53636_/X _53637_/Y sky130_fd_sc_hd__a21oi_4
X_72471_ _72461_/A _72471_/B _72471_/Y sky130_fd_sc_hd__nor2_4
X_84457_ _84454_/CLK _84457_/D _78080_/B sky130_fd_sc_hd__dfxtp_4
X_50849_ _50768_/A _50849_/X sky130_fd_sc_hd__buf_2
X_81669_ _81288_/CLK _79949_/X _81637_/D sky130_fd_sc_hd__dfxtp_4
X_74210_ _86979_/Q _57092_/X _74209_/X _74210_/Y sky130_fd_sc_hd__o21ai_4
X_40602_ _40420_/A _47943_/A sky130_fd_sc_hd__buf_2
X_59144_ _57757_/A _72358_/A sky130_fd_sc_hd__buf_2
X_71422_ _70407_/C _71432_/B _71422_/C _71365_/X _71422_/X sky130_fd_sc_hd__and4_4
X_83408_ _83482_/CLK _71697_/Y _58283_/A sky130_fd_sc_hd__dfxtp_4
X_44370_ _44370_/A _87143_/D sky130_fd_sc_hd__inv_2
X_56356_ _56358_/A _56358_/B _55756_/B _56356_/Y sky130_fd_sc_hd__nand3_4
X_75190_ _75190_/A _75190_/B _75190_/C _75190_/Y sky130_fd_sc_hd__nand3_4
X_87176_ _87178_/CLK _44258_/Y _87176_/Q sky130_fd_sc_hd__dfxtp_4
X_41582_ _41457_/A _41582_/X sky130_fd_sc_hd__buf_2
X_53568_ _85611_/Q _53556_/X _53567_/Y _53568_/Y sky130_fd_sc_hd__o21ai_4
X_84388_ _84392_/CLK _62723_/Y _75918_/B sky130_fd_sc_hd__dfxtp_4
X_43321_ _43320_/Y _87483_/D sky130_fd_sc_hd__inv_2
X_55307_ _55306_/X _45672_/Y _55307_/Y sky130_fd_sc_hd__nor2_4
X_86127_ _86127_/CLK _50817_/Y _86127_/Q sky130_fd_sc_hd__dfxtp_4
X_74141_ _86982_/Q _73370_/B _74141_/Y sky130_fd_sc_hd__nor2_4
X_40533_ _40477_/X _40488_/X _40532_/X _88375_/Q _40492_/X _40534_/A
+ sky130_fd_sc_hd__o32ai_4
X_52519_ _65103_/B _52516_/X _52518_/Y _52519_/Y sky130_fd_sc_hd__o21ai_4
X_59075_ _59061_/X _86075_/Q _59074_/X _59075_/Y sky130_fd_sc_hd__o21ai_4
X_71353_ _71429_/A _71363_/D sky130_fd_sc_hd__buf_2
X_83339_ _83362_/CLK _83339_/D _83339_/Q sky130_fd_sc_hd__dfxtp_4
X_56287_ _56368_/A _56270_/B _56287_/C _56287_/Y sky130_fd_sc_hd__nand3_4
X_53499_ _53458_/A _50275_/B _53499_/Y sky130_fd_sc_hd__nand2_4
X_46040_ _46039_/Y _86799_/D sky130_fd_sc_hd__inv_2
X_58026_ _58070_/A _58026_/B _58026_/Y sky130_fd_sc_hd__nor2_4
X_70304_ _70296_/X _70297_/X _70304_/C _70301_/D _70304_/X sky130_fd_sc_hd__and4_4
X_43252_ _43251_/Y _87518_/D sky130_fd_sc_hd__inv_2
X_55238_ _55655_/A _83316_/Q _55655_/B _55243_/B sky130_fd_sc_hd__nand3_4
X_74072_ _41957_/Y _72888_/X _73551_/X _74071_/Y _74072_/X sky130_fd_sc_hd__a211o_4
X_86058_ _85645_/CLK _86058_/D _86058_/Q sky130_fd_sc_hd__dfxtp_4
X_40464_ _46526_/A _40784_/A sky130_fd_sc_hd__buf_2
X_71284_ _53213_/B _71264_/X _71283_/Y _83547_/D sky130_fd_sc_hd__o21ai_4
X_42203_ _42203_/A _42203_/Y sky130_fd_sc_hd__inv_2
X_73023_ _83168_/Q _72943_/X _73022_/Y _73023_/X sky130_fd_sc_hd__a21o_4
X_77900_ _82245_/Q _81957_/Q _77900_/Y sky130_fd_sc_hd__xnor2_4
X_85009_ _85037_/CLK _57412_/X _57409_/A sky130_fd_sc_hd__dfxtp_4
X_70235_ _70224_/X _83828_/Q _70234_/X _70235_/X sky130_fd_sc_hd__a21o_4
X_43183_ _43182_/Y _43217_/A sky130_fd_sc_hd__buf_2
X_55169_ _55159_/A _85004_/Q _55169_/X sky130_fd_sc_hd__and2_4
X_78880_ _78875_/Y _78854_/B _78879_/Y _78880_/Y sky130_fd_sc_hd__o21ai_4
X_40395_ _40394_/X _40395_/X sky130_fd_sc_hd__buf_2
X_42134_ _42120_/X _42116_/X _41125_/X _88017_/Q _42117_/X _42134_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77831_ _82157_/Q _77831_/B _77831_/X sky130_fd_sc_hd__xor2_4
X_70166_ _70158_/Y _70157_/X _70165_/Y _83849_/D sky130_fd_sc_hd__o21ai_4
X_47991_ _48044_/A _47991_/B _47991_/Y sky130_fd_sc_hd__nand2_4
X_59977_ _59977_/A _59977_/B _59977_/Y sky130_fd_sc_hd__nand2_4
X_49730_ _49716_/X _52944_/B _49730_/Y sky130_fd_sc_hd__nand2_4
X_46942_ _82399_/Q _46942_/Y sky130_fd_sc_hd__inv_2
X_58928_ _58928_/A _58928_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_50_0_CLK clkbuf_7_50_0_CLK/A clkbuf_7_50_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_42065_ _40935_/X _41907_/X _88051_/Q _41912_/X _88051_/D sky130_fd_sc_hd__a2bb2o_4
X_77762_ _82262_/Q _81974_/Q _81926_/D sky130_fd_sc_hd__xor2_4
X_74974_ _80763_/Q _74965_/B _74974_/Y sky130_fd_sc_hd__nand2_4
X_70097_ _82530_/D _70085_/X _70096_/X _70097_/X sky130_fd_sc_hd__a21bo_4
Xclkbuf_8_190_0_CLK clkbuf_7_95_0_CLK/X clkbuf_8_190_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_79501_ _84816_/Q _84136_/Q _79503_/A sky130_fd_sc_hd__xor2_4
X_41016_ _41016_/A _41016_/X sky130_fd_sc_hd__buf_2
X_76713_ _76713_/A _76713_/B _81545_/D sky130_fd_sc_hd__xor2_4
X_49661_ _49580_/A _49661_/X sky130_fd_sc_hd__buf_2
X_73925_ _44126_/X _85906_/Q _73925_/X sky130_fd_sc_hd__and2_4
X_46873_ _86694_/Q _46859_/X _46872_/Y _46873_/Y sky130_fd_sc_hd__o21ai_4
X_58859_ _58756_/X _85930_/Q _58793_/X _58859_/X sky130_fd_sc_hd__o21a_4
X_77693_ _77693_/A _77680_/X _77693_/C _77693_/D _77694_/A sky130_fd_sc_hd__and4_4
X_48612_ _48612_/A _48612_/X sky130_fd_sc_hd__buf_2
X_79432_ _79429_/X _79431_/Y _79432_/X sky130_fd_sc_hd__xor2_4
X_45824_ _57071_/B _45824_/B _45824_/Y sky130_fd_sc_hd__nor2_4
X_76644_ _76639_/Y _81377_/Q _76640_/Y _76644_/Y sky130_fd_sc_hd__nand3_4
X_49592_ _49571_/X _49592_/B _49577_/C _52805_/D _49592_/X sky130_fd_sc_hd__and4_4
X_61870_ _61948_/A _61870_/X sky130_fd_sc_hd__buf_2
X_73856_ _73854_/X _85621_/Q _73782_/X _73855_/X _73856_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_7_65_0_CLK clkbuf_6_32_0_CLK/X clkbuf_7_65_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_60821_ _64738_/A _64561_/A sky130_fd_sc_hd__buf_2
X_72807_ _72929_/A _65451_/B _72807_/X sky130_fd_sc_hd__and2_4
X_48543_ _48043_/X _49048_/B _48542_/Y _48544_/A sky130_fd_sc_hd__o21ai_4
X_79363_ _79363_/A _79363_/B _79369_/B sky130_fd_sc_hd__xor2_4
X_45755_ _57448_/A _45705_/X _45691_/X _45755_/X sky130_fd_sc_hd__o21a_4
X_76575_ _76574_/Y _76575_/Y sky130_fd_sc_hd__inv_2
X_42967_ _42944_/X _42945_/X _40426_/X _66808_/B _42954_/X _42968_/A
+ sky130_fd_sc_hd__o32ai_4
X_73787_ _73742_/A _66041_/B _73787_/X sky130_fd_sc_hd__and2_4
X_70999_ _50827_/B _70983_/X _70998_/Y _70999_/Y sky130_fd_sc_hd__o21ai_4
X_78314_ _78314_/A _82754_/D _82466_/D sky130_fd_sc_hd__xor2_4
X_44706_ _44686_/X _44687_/X _40672_/Y _44705_/Y _44689_/X _86992_/D
+ sky130_fd_sc_hd__o32ai_4
X_63540_ _63540_/A _63541_/D sky130_fd_sc_hd__buf_2
X_75526_ _75525_/X _75528_/A sky130_fd_sc_hd__inv_2
X_41918_ _41992_/A _42477_/A sky130_fd_sc_hd__buf_2
X_48474_ _48471_/X _82359_/Q _48473_/Y _74416_/A sky130_fd_sc_hd__o21ai_4
X_60752_ _60761_/A _60752_/B _84575_/Q _60752_/Y sky130_fd_sc_hd__nor3_4
X_72738_ _72729_/X _72733_/X _72737_/X _72738_/X sky130_fd_sc_hd__a21o_4
X_79294_ _79280_/Y _79277_/X _79294_/X sky130_fd_sc_hd__and2_4
X_45686_ _45668_/X _61551_/A _45685_/X _45686_/Y sky130_fd_sc_hd__o21ai_4
X_42898_ _42898_/A _87662_/D sky130_fd_sc_hd__inv_2
X_47425_ _81804_/Q _47426_/A sky130_fd_sc_hd__inv_2
X_78245_ _78253_/B _82496_/Q _78244_/Y _78245_/Y sky130_fd_sc_hd__a21oi_4
X_44637_ _41032_/A _44618_/X _87022_/Q _44619_/X _87022_/D sky130_fd_sc_hd__a2bb2o_4
X_63471_ _63471_/A _63496_/D sky130_fd_sc_hd__buf_2
X_75457_ _75457_/A _75457_/B _75457_/C _75458_/A sky130_fd_sc_hd__or3_4
X_41849_ _40507_/X _41847_/X _67136_/B _41848_/X _41849_/X sky130_fd_sc_hd__a2bb2o_4
X_60683_ _63540_/A _63699_/D sky130_fd_sc_hd__buf_2
X_72669_ _70210_/C _72658_/X _72668_/Y _83196_/D sky130_fd_sc_hd__a21bo_4
X_65210_ _65172_/X _86122_/Q _65127_/X _65209_/X _65210_/X sky130_fd_sc_hd__a211o_4
X_62422_ _62336_/A _62479_/A sky130_fd_sc_hd__buf_2
X_74408_ _74408_/A _53663_/B _74408_/Y sky130_fd_sc_hd__nand2_4
X_47356_ _47355_/Y _53003_/D sky130_fd_sc_hd__buf_2
X_66190_ _65721_/X _66135_/B _65724_/X _66190_/Y sky130_fd_sc_hd__nand3_4
X_78176_ _78166_/Y _78175_/X _78176_/Y sky130_fd_sc_hd__nand2_4
X_44568_ _44549_/A _44568_/X sky130_fd_sc_hd__buf_2
X_75388_ _75351_/A _75354_/A _75362_/X _75404_/A sky130_fd_sc_hd__a21o_4
X_46307_ _48499_/A _46308_/A sky130_fd_sc_hd__buf_2
X_65141_ _84213_/Q _65142_/C sky130_fd_sc_hd__inv_2
X_77127_ _77127_/A _77127_/B _77127_/Y sky130_fd_sc_hd__nor2_4
X_43519_ _43518_/X _43503_/X _41791_/X _87380_/Q _43506_/X _43519_/Y
+ sky130_fd_sc_hd__o32ai_4
X_62353_ _62342_/A _62341_/X _84416_/Q _62353_/Y sky130_fd_sc_hd__nor3_4
X_74339_ _70326_/A _74327_/X _74338_/Y _74339_/X sky130_fd_sc_hd__a21bo_4
X_47287_ _47147_/A _47287_/X sky130_fd_sc_hd__buf_2
X_44499_ _44496_/X _44497_/X _41244_/X _87079_/Q _44498_/X _44500_/A
+ sky130_fd_sc_hd__o32ai_4
X_49026_ _49007_/A _49025_/X _49026_/Y sky130_fd_sc_hd__nand2_4
X_61304_ _72563_/C _72583_/C sky130_fd_sc_hd__buf_2
X_46238_ _73939_/A _86754_/D sky130_fd_sc_hd__buf_2
X_65072_ _65047_/A _65047_/B _65072_/C _65072_/Y sky130_fd_sc_hd__nor3_4
X_77058_ _77052_/Y _77057_/X _77068_/A sky130_fd_sc_hd__nand2_4
X_62284_ _62282_/Y _62253_/X _62283_/Y _62284_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_8_143_0_CLK clkbuf_7_71_0_CLK/X clkbuf_9_286_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_68900_ _68897_/X _68899_/X _68806_/X _68900_/X sky130_fd_sc_hd__a21o_4
X_64023_ _64021_/X _63994_/X _64022_/Y _64023_/Y sky130_fd_sc_hd__a21oi_4
X_76009_ _76009_/A _76009_/B _76009_/Y sky130_fd_sc_hd__nand2_4
X_61235_ _61264_/B _61149_/X _61215_/Y _61264_/A _61234_/Y _61235_/Y
+ sky130_fd_sc_hd__a41oi_4
X_46169_ _46166_/A _46128_/D _46169_/C _46169_/Y sky130_fd_sc_hd__nand3_4
X_69880_ _69461_/Y _69732_/X _69870_/X _69879_/Y _69880_/X sky130_fd_sc_hd__a211o_4
X_68831_ _68827_/X _68830_/X _68806_/X _68831_/X sky130_fd_sc_hd__a21o_4
X_61166_ _61160_/Y _61162_/X _61254_/B _61163_/Y _61165_/Y _84516_/D
+ sky130_fd_sc_hd__a41oi_4
Xclkbuf_7_18_0_CLK clkbuf_6_9_0_CLK/X clkbuf_8_37_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_60117_ _62193_/A _62244_/D sky130_fd_sc_hd__buf_2
X_49928_ _49928_/A _53141_/B _49928_/Y sky130_fd_sc_hd__nand2_4
X_68762_ _68993_/A _68762_/X sky130_fd_sc_hd__buf_2
X_65974_ _44174_/A _68347_/A sky130_fd_sc_hd__buf_2
X_61097_ _61096_/X _61097_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_158_0_CLK clkbuf_7_79_0_CLK/X clkbuf_8_158_0_CLK/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_153_0_CLK clkbuf_9_76_0_CLK/X _81275_/CLK sky130_fd_sc_hd__clkbuf_1
X_67713_ _67354_/X _67713_/X sky130_fd_sc_hd__buf_2
X_64925_ _64797_/X _86741_/Q _64772_/X _64924_/X _64926_/B sky130_fd_sc_hd__a211o_4
X_60048_ _59727_/X _60059_/A _60044_/Y _60045_/Y _60047_/Y _84671_/D
+ sky130_fd_sc_hd__a41oi_4
X_49859_ _49864_/A _53072_/B _49859_/Y sky130_fd_sc_hd__nand2_4
X_80971_ _80931_/CLK _75655_/X _80959_/D sky130_fd_sc_hd__dfxtp_4
X_68693_ _68587_/X _68693_/B _68693_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_783_0_CLK clkbuf_9_391_0_CLK/X _82491_/CLK sky130_fd_sc_hd__clkbuf_1
X_82710_ _82803_/CLK _82710_/D _82710_/Q sky130_fd_sc_hd__dfxtp_4
X_67644_ _67615_/X _67644_/B _67644_/X sky130_fd_sc_hd__and2_4
X_52870_ _85739_/Q _52848_/X _52869_/Y _52870_/Y sky130_fd_sc_hd__o21ai_4
X_64856_ _64778_/A _85816_/Q _64856_/X sky130_fd_sc_hd__and2_4
X_83690_ _83690_/CLK _83690_/D _47212_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_274_0_CLK clkbuf_9_274_0_CLK/A clkbuf_9_274_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_51821_ _85940_/Q _51817_/X _51820_/Y _51821_/Y sky130_fd_sc_hd__o21ai_4
X_63807_ _60906_/X _63858_/C sky130_fd_sc_hd__buf_2
X_82641_ _82896_/CLK _83993_/Q _78940_/A sky130_fd_sc_hd__dfxtp_4
X_67575_ _67575_/A _67575_/B _67575_/X sky130_fd_sc_hd__and2_4
X_64787_ _60151_/X _64775_/Y _64786_/Y _64787_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_168_0_CLK clkbuf_9_84_0_CLK/X _81682_/CLK sky130_fd_sc_hd__clkbuf_1
X_61999_ _61997_/X _61999_/B _61971_/C _61971_/D _62000_/D sky130_fd_sc_hd__nand4_4
X_69314_ _83933_/Q _69299_/X _69313_/X _69314_/X sky130_fd_sc_hd__a21bo_4
X_54540_ _54540_/A _54540_/X sky130_fd_sc_hd__buf_2
X_66526_ _60371_/A _66526_/X sky130_fd_sc_hd__buf_2
X_85360_ _86289_/CLK _85360_/D _85360_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_798_0_CLK clkbuf_9_399_0_CLK/X _81216_/CLK sky130_fd_sc_hd__clkbuf_1
X_51752_ _51758_/A _46625_/X _51752_/Y sky130_fd_sc_hd__nand2_4
X_63738_ _84729_/Q _63738_/B _63738_/C _63738_/D _63738_/Y sky130_fd_sc_hd__nand4_4
X_82572_ _82604_/CLK _82572_/D _78145_/A sky130_fd_sc_hd__dfxtp_4
X_84311_ _84308_/CLK _63593_/Y _84311_/Q sky130_fd_sc_hd__dfxtp_4
X_50703_ _86150_/Q _50680_/X _50702_/Y _50703_/Y sky130_fd_sc_hd__o21ai_4
X_81523_ _81514_/CLK _81567_/Q _81523_/Q sky130_fd_sc_hd__dfxtp_4
X_69245_ _69245_/A _69245_/X sky130_fd_sc_hd__buf_2
X_54471_ _54453_/X _54471_/B _54471_/C _46971_/Y _54471_/X sky130_fd_sc_hd__and4_4
X_66457_ _82735_/D _66457_/Y sky130_fd_sc_hd__inv_2
X_85291_ _80670_/CLK _85291_/D _85291_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_289_0_CLK clkbuf_8_144_0_CLK/X clkbuf_9_289_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_51683_ _52593_/A _51695_/A sky130_fd_sc_hd__buf_2
X_63669_ _63665_/Y _63666_/X _63668_/X _58352_/A _63363_/X _63669_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56210_ _56194_/X _56210_/X sky130_fd_sc_hd__buf_2
X_87030_ _88301_/CLK _87030_/D _87030_/Q sky130_fd_sc_hd__dfxtp_4
X_53422_ _53405_/X _47195_/A _53422_/Y sky130_fd_sc_hd__nand2_4
X_65408_ _65408_/A _86434_/Q _65408_/X sky130_fd_sc_hd__and2_4
X_84242_ _84241_/CLK _64482_/Y _79637_/B sky130_fd_sc_hd__dfxtp_4
X_50634_ _50624_/A _53854_/B _50634_/Y sky130_fd_sc_hd__nand2_4
X_57190_ _57189_/Y _57190_/Y sky130_fd_sc_hd__inv_2
X_81454_ _81492_/CLK _76764_/B _81454_/Q sky130_fd_sc_hd__dfxtp_4
X_69176_ _69021_/A _69176_/B _69176_/X sky130_fd_sc_hd__and2_4
X_66388_ _79455_/B _66389_/C sky130_fd_sc_hd__inv_2
Xclkbuf_10_721_0_CLK clkbuf_9_360_0_CLK/X _88283_/CLK sky130_fd_sc_hd__clkbuf_1
X_56141_ _56112_/X _56139_/X _56140_/Y _56141_/Y sky130_fd_sc_hd__o21ai_4
X_80405_ _80406_/B _80406_/A _80405_/X sky130_fd_sc_hd__or2_4
X_68127_ _82072_/D _68120_/X _68126_/X _68127_/X sky130_fd_sc_hd__a21bo_4
X_53353_ _53353_/A _53353_/B _53353_/Y sky130_fd_sc_hd__nand2_4
X_65339_ _65336_/X _65338_/X _65287_/X _65339_/X sky130_fd_sc_hd__a21o_4
X_84173_ _82746_/CLK _84173_/D _65855_/C sky130_fd_sc_hd__dfxtp_4
X_50565_ _50607_/A _48889_/B _50565_/Y sky130_fd_sc_hd__nand2_4
Xpsn_inst_psn_buff_6 _71216_/A _71236_/A2 sky130_fd_sc_hd__buf_2
X_81385_ _83932_/CLK _81385_/D _76857_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_212_0_CLK clkbuf_8_106_0_CLK/X clkbuf_9_212_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_52304_ _64826_/B _52297_/X _52303_/Y _52304_/Y sky130_fd_sc_hd__o21ai_4
X_83124_ _83145_/CLK _74070_/Y _83124_/Q sky130_fd_sc_hd__dfxtp_4
X_80336_ _80336_/A _80329_/Y _80330_/Y _80336_/Y sky130_fd_sc_hd__nand3_4
X_56072_ _56058_/X _56070_/X _56071_/Y _56072_/Y sky130_fd_sc_hd__o21ai_4
X_68058_ _68377_/A _68059_/A sky130_fd_sc_hd__buf_2
X_53284_ _53293_/A _53274_/B _53293_/C _52771_/D _53284_/X sky130_fd_sc_hd__and4_4
X_50496_ _50496_/A _50526_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_106_0_CLK clkbuf_9_53_0_CLK/X _87174_/CLK sky130_fd_sc_hd__clkbuf_1
X_55023_ _85333_/Q _55020_/X _55022_/Y _55023_/Y sky130_fd_sc_hd__o21ai_4
X_59900_ _59899_/X _59901_/A sky130_fd_sc_hd__buf_2
X_67009_ _87425_/Q _66915_/X _66984_/X _67008_/X _67009_/X sky130_fd_sc_hd__a211o_4
X_52235_ _52220_/A _48851_/B _52235_/Y sky130_fd_sc_hd__nand2_4
X_83055_ _85566_/CLK _83055_/D _83055_/Q sky130_fd_sc_hd__dfxtp_4
X_87932_ _82886_/CLK _87932_/D _87932_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_736_0_CLK clkbuf_9_368_0_CLK/X _87373_/CLK sky130_fd_sc_hd__clkbuf_1
X_80267_ _80266_/B _80267_/Y sky130_fd_sc_hd__inv_2
X_70020_ _69702_/X _69704_/X _69994_/X _70020_/X sky130_fd_sc_hd__a21o_4
X_82006_ _82008_/CLK _82038_/Q _77149_/A sky130_fd_sc_hd__dfxtp_4
X_59831_ _44315_/A _59831_/X sky130_fd_sc_hd__buf_2
X_52166_ _52166_/A _52194_/B _52182_/C _52166_/X sky130_fd_sc_hd__and3_4
X_87863_ _87073_/CLK _87863_/D _87863_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_227_0_CLK clkbuf_8_113_0_CLK/X clkbuf_9_227_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_80198_ _80198_/A _80198_/B _80221_/B sky130_fd_sc_hd__and2_4
X_51117_ _51112_/A _52807_/B _51117_/Y sky130_fd_sc_hd__nand2_4
X_86814_ _86814_/CLK _46016_/Y _86814_/Q sky130_fd_sc_hd__dfxtp_4
X_59762_ _59761_/X _59762_/Y sky130_fd_sc_hd__inv_2
X_52097_ _51956_/X _52097_/X sky130_fd_sc_hd__buf_2
X_56974_ _45626_/Y _56952_/X _56973_/X _85106_/D sky130_fd_sc_hd__o21ai_4
X_87794_ _88097_/CLK _87794_/D _69147_/B sky130_fd_sc_hd__dfxtp_4
X_58713_ _58625_/X _85461_/Q _58712_/X _58713_/Y sky130_fd_sc_hd__o21ai_4
X_51048_ _51021_/A _51058_/A sky130_fd_sc_hd__buf_2
X_55925_ _83034_/Q _55607_/A _44101_/A _55924_/X _55926_/B sky130_fd_sc_hd__a211o_4
X_86745_ _85529_/CLK _86745_/D _86745_/Q sky130_fd_sc_hd__dfxtp_4
X_71971_ _71968_/Y _71969_/X _71970_/Y _71971_/Y sky130_fd_sc_hd__a21boi_4
X_59693_ _59692_/Y _62185_/B sky130_fd_sc_hd__buf_2
X_83957_ _83957_/CLK _68881_/X _83957_/Q sky130_fd_sc_hd__dfxtp_4
X_73710_ _73709_/X _73711_/A sky130_fd_sc_hd__buf_2
X_58644_ _58125_/X _85787_/Q _58126_/X _58644_/X sky130_fd_sc_hd__o21a_4
X_70922_ _51031_/B _70909_/X _70921_/Y _70922_/Y sky130_fd_sc_hd__o21ai_4
X_82908_ _82906_/CLK _78270_/B _82908_/Q sky130_fd_sc_hd__dfxtp_4
X_55856_ _85267_/Q _55489_/A _55469_/X _55855_/X _55856_/X sky130_fd_sc_hd__a211o_4
X_43870_ _43869_/X _43870_/X sky130_fd_sc_hd__buf_2
X_74690_ _74689_/X _82984_/D sky130_fd_sc_hd__inv_2
X_86676_ _86359_/CLK _86676_/D _86676_/Q sky130_fd_sc_hd__dfxtp_4
X_83888_ _82339_/CLK _69905_/X _83888_/Q sky130_fd_sc_hd__dfxtp_4
X_42821_ _42820_/X _42821_/X sky130_fd_sc_hd__buf_2
X_54807_ _54807_/A _54825_/A sky130_fd_sc_hd__buf_2
X_73641_ _73641_/A _86558_/Q _73641_/X sky130_fd_sc_hd__and2_4
X_85627_ _86237_/CLK _85627_/D _85627_/Q sky130_fd_sc_hd__dfxtp_4
X_70853_ _46685_/X _70830_/Y _70852_/Y _70853_/Y sky130_fd_sc_hd__o21ai_4
X_58575_ _84817_/Q _58095_/X _58567_/X _58574_/X _84817_/D sky130_fd_sc_hd__a2bb2oi_4
X_82839_ _82740_/CLK _82839_/D _82839_/Q sky130_fd_sc_hd__dfxtp_4
X_55787_ _55784_/X _55786_/X _44110_/X _55787_/X sky130_fd_sc_hd__a21o_4
X_52999_ _52999_/A _52999_/B _52999_/Y sky130_fd_sc_hd__nand2_4
X_45540_ _45536_/X _45539_/X _45523_/X _45540_/X sky130_fd_sc_hd__a21o_4
X_57526_ _57524_/Y _57506_/X _57525_/X _84986_/D sky130_fd_sc_hd__a21oi_4
X_76360_ _76340_/X _76358_/Y _76359_/Y _76360_/Y sky130_fd_sc_hd__a21oi_4
X_42752_ _42752_/A _42752_/Y sky130_fd_sc_hd__inv_2
X_88346_ _87851_/CLK _88346_/D _88346_/Q sky130_fd_sc_hd__dfxtp_4
X_54738_ _54656_/X _54755_/B sky130_fd_sc_hd__buf_2
X_73572_ _73559_/Y _73572_/B _73572_/Y sky130_fd_sc_hd__xnor2_4
X_85558_ _85558_/CLK _53840_/Y _85558_/Q sky130_fd_sc_hd__dfxtp_4
X_70784_ _70871_/A _70791_/B _70791_/C _70791_/D _70784_/Y sky130_fd_sc_hd__nand4_4
X_75311_ _80690_/Q _80990_/Q _75311_/Y sky130_fd_sc_hd__nor2_4
X_41703_ _41604_/A _41703_/B _41703_/X sky130_fd_sc_hd__or2_4
X_72523_ _61260_/X _61319_/X _72503_/A _72602_/A sky130_fd_sc_hd__a21boi_4
X_84509_ _84623_/CLK _61201_/X _61200_/C sky130_fd_sc_hd__dfxtp_4
X_45471_ _45389_/X _45471_/X sky130_fd_sc_hd__buf_2
X_57457_ _57456_/Y _85001_/D sky130_fd_sc_hd__inv_2
X_76291_ _76288_/Y _76309_/B _76291_/X sky130_fd_sc_hd__xor2_4
X_88277_ _82301_/CLK _88277_/D _69547_/B sky130_fd_sc_hd__dfxtp_4
X_42683_ _41064_/X _42679_/X _69452_/B _42681_/X _42683_/X sky130_fd_sc_hd__a2bb2o_4
X_54669_ _54649_/X _47313_/Y _54669_/Y sky130_fd_sc_hd__nand2_4
X_85489_ _85489_/CLK _85489_/D _85489_/Q sky130_fd_sc_hd__dfxtp_4
X_47210_ _47210_/A _47181_/B _47210_/C _51225_/D _47210_/X sky130_fd_sc_hd__and4_4
X_78030_ _78030_/A _78031_/B sky130_fd_sc_hd__inv_2
X_44422_ _44404_/X _44405_/X _41565_/X _87115_/Q _44406_/X _44422_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56408_ _56070_/X _56394_/X _56407_/Y _85205_/D sky130_fd_sc_hd__o21ai_4
X_87228_ _87487_/CLK _87228_/D _68944_/B sky130_fd_sc_hd__dfxtp_4
X_75242_ _75242_/A _75216_/Y _75243_/A sky130_fd_sc_hd__nor2_4
X_41634_ _40620_/X _41634_/B _41634_/X sky130_fd_sc_hd__or2_4
X_48190_ _48190_/A _51947_/B _48190_/Y sky130_fd_sc_hd__nand2_4
X_72454_ _83253_/Q _72445_/X _72448_/X _72453_/X _83253_/D sky130_fd_sc_hd__a2bb2oi_4
X_57388_ _57384_/X _56578_/X _85022_/Q _57385_/X _57388_/X sky130_fd_sc_hd__a2bb2o_4
X_47141_ _82378_/Q _54571_/D sky130_fd_sc_hd__inv_2
X_59127_ _59123_/Y _59126_/Y _59053_/X _59127_/X sky130_fd_sc_hd__a21o_4
X_71405_ _71397_/X _83511_/Q _71404_/Y _83511_/D sky130_fd_sc_hd__a21o_4
X_44353_ _44352_/X _44353_/X sky130_fd_sc_hd__buf_2
X_56339_ _56345_/A _56345_/B _56339_/C _56339_/Y sky130_fd_sc_hd__nand3_4
X_75173_ _75169_/Y _75171_/Y _75172_/Y _75178_/A sky130_fd_sc_hd__o21ai_4
X_87159_ _86935_/CLK _87159_/D _87159_/Q sky130_fd_sc_hd__dfxtp_4
X_41565_ _41564_/X _41565_/X sky130_fd_sc_hd__buf_2
X_72385_ _72299_/X _72382_/Y _72384_/Y _72337_/X _72303_/X _72385_/X
+ sky130_fd_sc_hd__o32a_4
X_43304_ _43166_/A _43305_/A sky130_fd_sc_hd__buf_2
X_74124_ _68959_/B _57376_/X _72798_/X _74123_/Y _74124_/X sky130_fd_sc_hd__a211o_4
X_40516_ _40477_/X _40488_/X _40515_/X _88379_/Q _40492_/X _40516_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47072_ _86673_/Q _47050_/X _47071_/Y _47072_/Y sky130_fd_sc_hd__o21ai_4
X_71336_ _50383_/B _71320_/A _71335_/Y _71336_/Y sky130_fd_sc_hd__o21ai_4
X_59058_ _59027_/X _59056_/Y _59057_/Y _59046_/X _59031_/X _59058_/X
+ sky130_fd_sc_hd__o32a_4
X_44284_ _44072_/Y _57650_/A _44284_/C _44284_/Y sky130_fd_sc_hd__nor3_4
X_79981_ _79965_/Y _79964_/A _79963_/Y _79981_/Y sky130_fd_sc_hd__a21boi_4
X_41496_ _41513_/A _82330_/Q _41496_/X sky130_fd_sc_hd__or2_4
X_46023_ _45975_/X _46023_/X sky130_fd_sc_hd__buf_2
X_58009_ _57996_/Y _57981_/X _58004_/X _58008_/X _84933_/D sky130_fd_sc_hd__a22oi_4
X_43235_ _43226_/X _43229_/X _41016_/X _87525_/Q _43232_/X _43236_/A
+ sky130_fd_sc_hd__o32ai_4
X_74055_ _74052_/X _74054_/X _73944_/X _74055_/X sky130_fd_sc_hd__a21o_4
X_78932_ _78918_/Y _78931_/X _78937_/A sky130_fd_sc_hd__nand2_4
X_40447_ _44736_/A _40447_/X sky130_fd_sc_hd__buf_2
X_71267_ _71266_/X _71268_/A sky130_fd_sc_hd__buf_2
X_61020_ _59508_/X _61020_/X sky130_fd_sc_hd__buf_2
X_73006_ _56274_/X _73006_/X sky130_fd_sc_hd__buf_2
X_70218_ _70233_/A _70229_/D sky130_fd_sc_hd__buf_2
X_43166_ _43166_/A _43167_/A sky130_fd_sc_hd__buf_2
X_78863_ _82841_/Q _82553_/Q _78877_/A sky130_fd_sc_hd__xor2_4
X_40378_ _40629_/A _47825_/A sky130_fd_sc_hd__buf_2
X_71198_ _48551_/X _71190_/X _71197_/Y _71198_/Y sky130_fd_sc_hd__o21ai_4
X_42117_ _42096_/A _42117_/X sky130_fd_sc_hd__buf_2
X_77814_ _82268_/Q _77814_/B _77814_/Y sky130_fd_sc_hd__xnor2_4
X_70149_ _70149_/A _70146_/Y _70147_/Y _70148_/Y _70149_/X sky130_fd_sc_hd__and4_4
X_47974_ _47971_/X _82932_/Q _47973_/X _47975_/B sky130_fd_sc_hd__o21ai_4
X_43097_ _43085_/X _43086_/X _40734_/X _43096_/Y _43090_/X _87577_/D
+ sky130_fd_sc_hd__o32ai_4
X_78794_ _78794_/A _78795_/B sky130_fd_sc_hd__inv_2
X_49713_ _49708_/A _49697_/B _49724_/C _52927_/D _49713_/X sky130_fd_sc_hd__and4_4
X_46925_ _46924_/Y _52750_/D sky130_fd_sc_hd__buf_2
X_42048_ _42035_/X _42010_/X _40899_/X _42047_/Y _42037_/X _88058_/D
+ sky130_fd_sc_hd__o32ai_4
X_77745_ _77743_/A _77741_/Y _77739_/Y _77745_/Y sky130_fd_sc_hd__a21oi_4
X_62971_ _62971_/A _64536_/C _60302_/X _62979_/D _62971_/X sky130_fd_sc_hd__and4_4
X_74957_ _80762_/Q _74957_/B _74971_/A sky130_fd_sc_hd__xor2_4
X_64710_ _64710_/A _64710_/B _64710_/X sky130_fd_sc_hd__and2_4
X_61922_ _84877_/Q _61922_/X sky130_fd_sc_hd__buf_2
X_49644_ _49638_/A _52859_/B _49644_/Y sky130_fd_sc_hd__nand2_4
X_73908_ _73954_/A _66119_/B _73908_/X sky130_fd_sc_hd__and2_4
X_46856_ _46856_/A _52716_/D sky130_fd_sc_hd__buf_2
X_65690_ _65638_/X _85584_/Q _65669_/X _65689_/X _65690_/X sky130_fd_sc_hd__a211o_4
X_77676_ _77676_/A _77673_/Y _77675_/Y _77676_/X sky130_fd_sc_hd__or3_4
X_74888_ _74888_/A _74887_/Y _74889_/A sky130_fd_sc_hd__and2_4
X_79415_ _79415_/A _79414_/X _79416_/B sky130_fd_sc_hd__xnor2_4
X_45807_ _45797_/X _45804_/Y _45806_/Y _45807_/Y sky130_fd_sc_hd__a21oi_4
X_64641_ _64564_/X _86143_/Q _64566_/X _64640_/X _64641_/X sky130_fd_sc_hd__a211o_4
X_76627_ _76624_/Y _76640_/A _76628_/A sky130_fd_sc_hd__nand2_4
X_49575_ _86362_/Q _49551_/X _49574_/Y _49575_/Y sky130_fd_sc_hd__o21ai_4
X_61853_ _61871_/A _61839_/B _61839_/C _63100_/B _61853_/X sky130_fd_sc_hd__and4_4
X_73839_ _73367_/A _73839_/X sky130_fd_sc_hd__buf_2
X_46787_ _54364_/B _50981_/B sky130_fd_sc_hd__buf_2
X_43999_ _59516_/A _59598_/A sky130_fd_sc_hd__buf_2
X_48526_ _74437_/B _48788_/B sky130_fd_sc_hd__buf_2
X_60804_ _63699_/D _60804_/B _60804_/C _60804_/Y sky130_fd_sc_hd__nor3_4
X_67360_ _67359_/X _67360_/X sky130_fd_sc_hd__buf_2
X_79346_ _79346_/A _79346_/B _79346_/X sky130_fd_sc_hd__or2_4
X_45738_ _85035_/Q _45738_/Y sky130_fd_sc_hd__inv_2
X_64572_ _58785_/A _64572_/B _64572_/X sky130_fd_sc_hd__and2_4
X_76558_ _76554_/X _76555_/Y _76560_/B _76559_/A sky130_fd_sc_hd__a21oi_4
X_61784_ _61752_/A _61723_/X _78077_/B _61784_/Y sky130_fd_sc_hd__nor3_4
X_66311_ _66236_/X _85605_/Q _66251_/X _66310_/X _66311_/X sky130_fd_sc_hd__a211o_4
X_63523_ _63523_/A _61939_/X _63523_/X sky130_fd_sc_hd__and2_4
X_75509_ _75509_/A _75481_/X _75509_/C _75458_/X _75509_/Y sky130_fd_sc_hd__nand4_4
X_48457_ _73016_/B _48419_/X _48456_/Y _48457_/Y sky130_fd_sc_hd__o21ai_4
X_60735_ _60720_/A _63400_/C sky130_fd_sc_hd__buf_2
X_67291_ _88373_/Q _67193_/X _67194_/X _67290_/X _67291_/X sky130_fd_sc_hd__a211o_4
X_79277_ _58856_/Y _66484_/Y _79276_/Y _79277_/X sky130_fd_sc_hd__o21a_4
X_45669_ _63206_/B _61542_/A sky130_fd_sc_hd__buf_2
X_76489_ _76489_/A _81541_/Q _76489_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_4_15_0_CLK clkbuf_3_7_1_CLK/X clkbuf_4_15_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_69030_ _69233_/A _69134_/A sky130_fd_sc_hd__buf_2
X_47408_ _47418_/A _47408_/B _47377_/X _53031_/D _47408_/X sky130_fd_sc_hd__and4_4
X_66242_ _66226_/A _66242_/B _66242_/X sky130_fd_sc_hd__and2_4
X_78228_ _78228_/A _78228_/B _78228_/Y sky130_fd_sc_hd__nand2_4
X_63454_ _63434_/X _63448_/X _63449_/X _63452_/X _63453_/Y _63454_/Y
+ sky130_fd_sc_hd__o41ai_4
X_48388_ _48388_/A _48364_/X _48354_/X _48388_/X sky130_fd_sc_hd__and3_4
X_60666_ _60665_/X _60667_/A sky130_fd_sc_hd__buf_2
X_62405_ _61490_/X _62420_/B _62420_/C _62404_/X _62405_/Y sky130_fd_sc_hd__nand4_4
X_47339_ _81813_/Q _54685_/D sky130_fd_sc_hd__inv_2
X_66173_ _66173_/A _66385_/B _66173_/C _66173_/Y sky130_fd_sc_hd__nand3_4
X_78159_ _78156_/Y _78159_/B _78160_/B sky130_fd_sc_hd__xor2_4
X_63385_ _58412_/A _63370_/X _61358_/A _63372_/X _63385_/X sky130_fd_sc_hd__a2bb2o_4
X_60597_ _79131_/A _60577_/X _60586_/D _60596_/Y _60597_/Y sky130_fd_sc_hd__a2bb2oi_4
X_65124_ _64924_/A _65124_/B _65124_/X sky130_fd_sc_hd__and2_4
X_50350_ _86218_/Q _50316_/X _50349_/Y _50350_/Y sky130_fd_sc_hd__o21ai_4
X_62336_ _62336_/A _62337_/A sky130_fd_sc_hd__buf_2
X_81170_ _82335_/CLK _74964_/B _81170_/Q sky130_fd_sc_hd__dfxtp_4
X_49009_ _49009_/A _49009_/B _49009_/Y sky130_fd_sc_hd__nor2_4
X_80121_ _80121_/A _80121_/B _80121_/Y sky130_fd_sc_hd__nand2_4
X_65055_ _64704_/X _86736_/Q _64707_/X _65054_/X _65055_/X sky130_fd_sc_hd__a211o_4
X_69932_ _69897_/A _69932_/B _69932_/Y sky130_fd_sc_hd__nor2_4
Xpsn_inst_psn_buff_13 _55686_/C _56892_/C sky130_fd_sc_hd__buf_2
X_50281_ _50278_/Y _50274_/X _50280_/Y _86232_/D sky130_fd_sc_hd__a21boi_4
X_62267_ _62267_/A _62267_/B _76998_/B _62267_/Y sky130_fd_sc_hd__nor3_4
Xpsn_inst_psn_buff_24 _53441_/A _53450_/A sky130_fd_sc_hd__buf_2
X_52020_ _66153_/B _51994_/X _52019_/Y _52020_/Y sky130_fd_sc_hd__o21ai_4
X_64006_ _64001_/X _63969_/X _64002_/Y _64003_/Y _64005_/X _64006_/X
+ sky130_fd_sc_hd__a41o_4
X_61218_ _61103_/X _61096_/X _72590_/A _61218_/Y sky130_fd_sc_hd__o21ai_4
X_80052_ _80030_/A _80052_/B _80052_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_1008_0_CLK clkbuf_9_504_0_CLK/X _83572_/CLK sky130_fd_sc_hd__clkbuf_1
X_69863_ _73323_/A _68377_/X _66574_/X _69862_/Y _69863_/X sky130_fd_sc_hd__a211o_4
X_62198_ _62237_/A _62198_/B _59985_/A _59943_/A _62198_/Y sky130_fd_sc_hd__nand4_4
X_68814_ _88001_/Q _68715_/X _68540_/X _68813_/X _68814_/X sky130_fd_sc_hd__a211o_4
X_61149_ _61148_/X _61149_/X sky130_fd_sc_hd__buf_2
X_84860_ _84358_/CLK _58395_/X _84860_/Q sky130_fd_sc_hd__dfxtp_4
X_69794_ _73198_/A _69751_/X _69779_/X _69793_/Y _69794_/X sky130_fd_sc_hd__a211o_4
X_83811_ _83813_/CLK _70286_/X _74756_/B sky130_fd_sc_hd__dfxtp_4
X_68745_ _68617_/A _68745_/X sky130_fd_sc_hd__buf_2
X_53971_ _53956_/X _53971_/B _53971_/Y sky130_fd_sc_hd__nand2_4
X_65957_ _64593_/A _85917_/Q _65957_/X sky130_fd_sc_hd__and2_4
X_84791_ _86697_/CLK _58908_/Y _84791_/Q sky130_fd_sc_hd__dfxtp_4
X_55710_ _83011_/Q _55710_/B _55710_/Y sky130_fd_sc_hd__nand2_4
X_86530_ _86530_/CLK _86530_/D _86530_/Q sky130_fd_sc_hd__dfxtp_4
X_64908_ _64905_/X _64907_/X _64729_/X _64908_/X sky130_fd_sc_hd__a21o_4
X_52922_ _52922_/A _52916_/B _52900_/C _47218_/D _52922_/X sky130_fd_sc_hd__and4_4
X_83742_ _86322_/CLK _70607_/Y _47323_/A sky130_fd_sc_hd__dfxtp_4
X_56690_ _46233_/Y _56691_/A sky130_fd_sc_hd__buf_2
X_80954_ _81197_/CLK _75424_/B _80954_/Q sky130_fd_sc_hd__dfxtp_4
X_68676_ _68750_/A _88359_/Q _68676_/X sky130_fd_sc_hd__and2_4
X_65888_ _65888_/A _65888_/B _65888_/C _65888_/Y sky130_fd_sc_hd__nor3_4
X_55641_ _55641_/A _55640_/Y _55641_/Y sky130_fd_sc_hd__nor2_4
X_67627_ _87911_/Q _67533_/X _67625_/X _67626_/X _67627_/X sky130_fd_sc_hd__a211o_4
X_86461_ _83623_/CLK _86461_/D _86461_/Q sky130_fd_sc_hd__dfxtp_4
X_52853_ _52853_/A _52853_/B _52853_/C _52853_/D _52853_/X sky130_fd_sc_hd__and4_4
X_64839_ _64825_/Y _64838_/Y _64839_/Y sky130_fd_sc_hd__nand2_4
X_83673_ _83673_/CLK _70889_/Y _46769_/A sky130_fd_sc_hd__dfxtp_4
X_80885_ _80854_/CLK _75748_/B _80885_/Q sky130_fd_sc_hd__dfxtp_4
X_88200_ _88133_/CLK _41517_/Y _88200_/Q sky130_fd_sc_hd__dfxtp_4
X_85412_ _85635_/CLK _85412_/D _85412_/Q sky130_fd_sc_hd__dfxtp_4
X_51804_ _51804_/A _51805_/A sky130_fd_sc_hd__buf_2
X_58360_ _58360_/A _58364_/B _58360_/Y sky130_fd_sc_hd__nand2_4
X_82624_ _82624_/CLK _79094_/X _82624_/Q sky130_fd_sc_hd__dfxtp_4
X_55572_ _44063_/X _55572_/X sky130_fd_sc_hd__buf_2
X_67558_ _67082_/A _67582_/A sky130_fd_sc_hd__buf_2
X_86392_ _86393_/CLK _49414_/Y _86392_/Q sky130_fd_sc_hd__dfxtp_4
X_52784_ _52757_/A _52784_/X sky130_fd_sc_hd__buf_2
X_57311_ _56730_/X _56766_/X _56785_/D _57318_/D _56767_/X _57311_/X
+ sky130_fd_sc_hd__a41o_4
X_88131_ _86796_/CLK _41832_/X _88131_/Q sky130_fd_sc_hd__dfxtp_4
X_54523_ _54519_/Y _54502_/X _54522_/X _54523_/Y sky130_fd_sc_hd__a21oi_4
X_66509_ _64867_/B _66501_/B _66509_/C _66509_/X sky130_fd_sc_hd__and3_4
X_85343_ _85375_/CLK _54975_/Y _85343_/Q sky130_fd_sc_hd__dfxtp_4
X_51735_ _52588_/A _51721_/X _51715_/C _53257_/D _51735_/X sky130_fd_sc_hd__and4_4
X_58291_ _84886_/Q _63672_/B sky130_fd_sc_hd__buf_2
X_82555_ _82596_/CLK _82555_/D _82555_/Q sky130_fd_sc_hd__dfxtp_4
X_67489_ _67486_/X _67488_/X _67442_/X _67489_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_10_660_0_CLK clkbuf_9_330_0_CLK/X _87116_/CLK sky130_fd_sc_hd__clkbuf_1
X_57242_ _44288_/X _56584_/X _45460_/A _57238_/X _85053_/D sky130_fd_sc_hd__a2bb2o_4
X_81506_ _83918_/CLK _76155_/B _81506_/Q sky130_fd_sc_hd__dfxtp_4
X_69228_ _69216_/X _69226_/Y _69095_/X _69227_/Y _69228_/X sky130_fd_sc_hd__a211o_4
X_88062_ _88062_/CLK _88062_/D _42036_/A sky130_fd_sc_hd__dfxtp_4
X_54454_ _54401_/A _54471_/C sky130_fd_sc_hd__buf_2
X_85274_ _85277_/CLK _56212_/Y _56211_/C sky130_fd_sc_hd__dfxtp_4
X_51666_ _85968_/Q _51647_/X _51665_/Y _51666_/Y sky130_fd_sc_hd__o21ai_4
X_82486_ _82485_/CLK _82486_/D _82862_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_151_0_CLK clkbuf_8_75_0_CLK/X clkbuf_9_151_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_87013_ _88288_/CLK _44657_/Y _87013_/Q sky130_fd_sc_hd__dfxtp_4
X_53405_ _53352_/A _53405_/X sky130_fd_sc_hd__buf_2
X_84225_ _84223_/CLK _84225_/D _84225_/Q sky130_fd_sc_hd__dfxtp_4
X_50617_ _50597_/A _48992_/X _50617_/Y sky130_fd_sc_hd__nand2_4
X_81437_ _82648_/CLK _81469_/Q _76116_/B sky130_fd_sc_hd__dfxtp_4
X_57173_ _85068_/Q _56997_/X _57173_/Y sky130_fd_sc_hd__nor2_4
X_69159_ _69146_/X _69109_/X _69157_/Y _69158_/Y _69159_/X sky130_fd_sc_hd__a211o_4
X_54385_ _54385_/A _54395_/B sky130_fd_sc_hd__buf_2
X_51597_ _85981_/Q _51594_/X _51596_/Y _51597_/Y sky130_fd_sc_hd__o21ai_4
X_56124_ _56131_/A _56140_/B _56124_/C _56124_/Y sky130_fd_sc_hd__nand3_4
X_41350_ _41350_/A _41325_/X _41350_/X sky130_fd_sc_hd__or2_4
X_53336_ _53332_/A _53336_/B _53336_/Y sky130_fd_sc_hd__nand2_4
X_72170_ _59368_/X _85981_/Q _72169_/X _72170_/Y sky130_fd_sc_hd__o21ai_4
X_84156_ _82177_/CLK _84156_/D _84156_/Q sky130_fd_sc_hd__dfxtp_4
X_50548_ _50546_/Y _50525_/X _50547_/X _86180_/D sky130_fd_sc_hd__a21oi_4
X_81368_ _81333_/CLK _81368_/D _76486_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_675_0_CLK clkbuf_9_337_0_CLK/X _87652_/CLK sky130_fd_sc_hd__clkbuf_1
X_71121_ _71112_/X _71076_/B _71119_/C _71121_/Y sky130_fd_sc_hd__nand3_4
X_83107_ _82998_/CLK _83107_/D _70285_/C sky130_fd_sc_hd__dfxtp_4
X_56055_ _56055_/A _56055_/X sky130_fd_sc_hd__buf_2
X_80319_ _80318_/Y _80319_/B _80320_/B sky130_fd_sc_hd__nand2_4
X_53267_ _53264_/Y _51904_/X _53266_/X _53267_/Y sky130_fd_sc_hd__a21oi_4
X_41281_ _41255_/X _40760_/A _41280_/X _41281_/Y sky130_fd_sc_hd__o21ai_4
X_84087_ _84087_/CLK _84087_/D _80911_/D sky130_fd_sc_hd__dfxtp_4
X_50479_ _52182_/A _50492_/B _50497_/C _50479_/X sky130_fd_sc_hd__and3_4
X_81299_ _81279_/CLK _76987_/X _81267_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_166_0_CLK clkbuf_8_83_0_CLK/X clkbuf_9_166_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_55006_ _55003_/Y _54998_/X _55005_/X _85337_/D sky130_fd_sc_hd__a21oi_4
X_43020_ _43020_/A _43024_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_93_0_CLK clkbuf_9_93_0_CLK/A clkbuf_9_93_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_52218_ _52218_/A _52198_/X _52218_/C _52218_/X sky130_fd_sc_hd__and3_4
X_71052_ _71055_/A _70942_/B _71055_/C _71052_/Y sky130_fd_sc_hd__nand3_4
X_87915_ _87915_/CLK _87915_/D _87915_/Q sky130_fd_sc_hd__dfxtp_4
X_83038_ _83001_/CLK _74548_/Y _74547_/C sky130_fd_sc_hd__dfxtp_4
X_53198_ _53172_/A _53198_/X sky130_fd_sc_hd__buf_2
X_70003_ _69943_/X _68525_/Y _69984_/X _70002_/Y _70003_/X sky130_fd_sc_hd__a211o_4
X_59814_ _60341_/A _59814_/X sky130_fd_sc_hd__buf_2
X_52149_ _73040_/B _52125_/X _52148_/Y _52149_/Y sky130_fd_sc_hd__o21ai_4
X_75860_ _75860_/A _75860_/B _75860_/X sky130_fd_sc_hd__xor2_4
X_87846_ _87850_/CLK _87846_/D _68692_/A sky130_fd_sc_hd__dfxtp_4
X_74811_ _83841_/Q _74731_/X _74804_/X _74805_/X _74810_/Y _74811_/X
+ sky130_fd_sc_hd__a2111o_4
X_59745_ _59651_/B _59745_/X sky130_fd_sc_hd__buf_2
X_44971_ _44904_/A _44972_/A sky130_fd_sc_hd__inv_2
X_56957_ _56602_/X _85113_/Q _56953_/X _56957_/Y sky130_fd_sc_hd__nor3_4
X_75791_ _75778_/A _75789_/Y _75790_/X _75791_/Y sky130_fd_sc_hd__o21ai_4
X_87777_ _87525_/CLK _42672_/Y _69381_/B sky130_fd_sc_hd__dfxtp_4
X_84989_ _84991_/CLK _84989_/D _84989_/Q sky130_fd_sc_hd__dfxtp_4
X_46710_ _83679_/Q _52632_/B sky130_fd_sc_hd__inv_2
X_77530_ _77518_/A _82114_/Q _77530_/Y sky130_fd_sc_hd__nand2_4
X_43922_ _43916_/X _43902_/X _41403_/X _67856_/B _43917_/X _43922_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55908_ _55908_/A _55908_/B _55908_/X sky130_fd_sc_hd__and2_4
X_86728_ _86121_/CLK _46541_/Y _86728_/Q sky130_fd_sc_hd__dfxtp_4
X_74742_ _70588_/A _74742_/B _71039_/D _74752_/A sky130_fd_sc_hd__nand3_4
X_47690_ _81232_/Q _47691_/A sky130_fd_sc_hd__inv_2
X_59676_ _59696_/A _66514_/B _80614_/A _59676_/Y sky130_fd_sc_hd__nor3_4
X_71954_ _56908_/A _71939_/X _71953_/Y _83315_/D sky130_fd_sc_hd__o21ai_4
X_56888_ _56572_/X _56886_/Y _56887_/Y _85126_/D sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_613_0_CLK clkbuf_9_306_0_CLK/X _80991_/CLK sky130_fd_sc_hd__clkbuf_1
X_46641_ _83686_/Q _52590_/B sky130_fd_sc_hd__inv_2
X_70905_ _70905_/A _70903_/B _70899_/C _70905_/D _70905_/Y sky130_fd_sc_hd__nand4_4
X_58627_ _58625_/X _85468_/Q _58626_/X _58627_/Y sky130_fd_sc_hd__o21ai_4
X_77461_ _77424_/Y _77426_/X _77449_/X _77461_/X sky130_fd_sc_hd__a21bo_4
X_43853_ _43852_/Y _87233_/D sky130_fd_sc_hd__inv_2
X_55839_ _56420_/C _44063_/X _55523_/X _55838_/X _55839_/X sky130_fd_sc_hd__a211o_4
X_74673_ _74673_/A _45713_/A _74673_/Y sky130_fd_sc_hd__nand2_4
X_86659_ _86665_/CLK _47211_/Y _59373_/A sky130_fd_sc_hd__dfxtp_4
X_71885_ _71863_/A _71783_/A _71783_/C _71883_/D _71885_/Y sky130_fd_sc_hd__nor4_4
Xclkbuf_9_104_0_CLK clkbuf_8_52_0_CLK/X clkbuf_9_104_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_79200_ _84789_/Q _66509_/C _79201_/A sky130_fd_sc_hd__nor2_4
X_76412_ _76408_/Y _76409_/Y _76411_/Y _76412_/X sky130_fd_sc_hd__or3_4
X_42804_ _41397_/X _42802_/X _87710_/Q _42803_/X _42804_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_9_31_0_CLK clkbuf_9_31_0_CLK/A clkbuf_9_31_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_49360_ _49415_/A _49360_/X sky130_fd_sc_hd__buf_2
X_73624_ _72978_/X _73624_/X sky130_fd_sc_hd__buf_2
X_70836_ _70863_/A _70846_/B _71066_/C _70841_/D _70836_/Y sky130_fd_sc_hd__nand4_4
X_46572_ _83780_/Q _52563_/B sky130_fd_sc_hd__inv_2
X_58558_ _58538_/X _83355_/Q _58557_/Y _84819_/D sky130_fd_sc_hd__o21a_4
X_77392_ _77392_/A _77394_/A sky130_fd_sc_hd__inv_2
X_43784_ _43774_/X _43781_/X _41016_/X _69332_/B _43776_/X _43784_/Y
+ sky130_fd_sc_hd__o32ai_4
X_40996_ _40944_/X _40946_/X _40994_/X _88296_/Q _40995_/X _40996_/Y
+ sky130_fd_sc_hd__o32ai_4
X_48311_ _66256_/B _48293_/X _48310_/Y _48311_/Y sky130_fd_sc_hd__o21ai_4
X_79131_ _79131_/A _79131_/B _79131_/X sky130_fd_sc_hd__xor2_4
X_45523_ _45678_/A _45523_/X sky130_fd_sc_hd__buf_2
X_57509_ _57499_/A _47880_/Y _57509_/Y sky130_fd_sc_hd__nand2_4
X_76343_ _76343_/A _81615_/D _76343_/X sky130_fd_sc_hd__xor2_4
X_88329_ _87288_/CLK _40816_/Y _88329_/Q sky130_fd_sc_hd__dfxtp_4
X_42735_ _42721_/X _42723_/X _41214_/X _68848_/B _42732_/X _42736_/A
+ sky130_fd_sc_hd__o32ai_4
X_49291_ _49232_/A _51320_/B _49291_/Y sky130_fd_sc_hd__nand2_4
X_73555_ _43587_/Y _73030_/X _73486_/X _73554_/Y _73555_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_628_0_CLK clkbuf_9_314_0_CLK/X _82131_/CLK sky130_fd_sc_hd__clkbuf_1
X_70767_ _52837_/B _70761_/X _70766_/Y _70767_/Y sky130_fd_sc_hd__o21ai_4
X_58489_ _84836_/Q _58490_/A sky130_fd_sc_hd__inv_2
X_48242_ _48186_/A _49223_/A sky130_fd_sc_hd__buf_2
X_60520_ _60359_/X _60517_/Y _60481_/A _60518_/X _60519_/Y _60520_/Y
+ sky130_fd_sc_hd__a41oi_4
X_72506_ _72516_/C _72535_/A _72506_/C _72535_/B _72506_/Y sky130_fd_sc_hd__nand4_4
X_79062_ _82654_/Q _79064_/A sky130_fd_sc_hd__inv_2
X_45454_ _45447_/X _45450_/X _45453_/Y _45454_/Y sky130_fd_sc_hd__a21oi_4
X_76274_ _76274_/A _81610_/D _76274_/X sky130_fd_sc_hd__xor2_4
X_42666_ _42592_/A _42666_/X sky130_fd_sc_hd__buf_2
X_73486_ _72857_/X _73486_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_119_0_CLK clkbuf_8_59_0_CLK/X clkbuf_9_119_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_70698_ _70698_/A _70698_/B _70699_/A sky130_fd_sc_hd__nor2_4
Xclkbuf_9_46_0_CLK clkbuf_9_47_0_CLK/A clkbuf_9_46_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_78013_ _77999_/B _78013_/Y sky130_fd_sc_hd__inv_2
X_44405_ _44382_/A _44405_/X sky130_fd_sc_hd__buf_2
X_75225_ _75226_/A _80985_/Q _75225_/Y sky130_fd_sc_hd__nor2_4
X_41617_ _41611_/X _41613_/X _41616_/X _67279_/B _41608_/X _41617_/Y
+ sky130_fd_sc_hd__o32ai_4
X_72437_ _86598_/Q _72428_/B _72437_/Y sky130_fd_sc_hd__nor2_4
X_48173_ _50048_/A _50224_/B _48173_/Y sky130_fd_sc_hd__nand2_4
X_60451_ _60408_/C _60408_/A _60439_/X _60440_/X _60588_/A _60572_/C
+ sky130_fd_sc_hd__a41o_4
X_45385_ _45377_/X _45382_/Y _45384_/Y _45385_/Y sky130_fd_sc_hd__a21oi_4
X_42597_ _42580_/A _42597_/X sky130_fd_sc_hd__buf_2
X_47124_ _53386_/B _52869_/B sky130_fd_sc_hd__buf_2
X_44336_ _44330_/X _44331_/X _41667_/X _87160_/Q _44332_/X _44336_/Y
+ sky130_fd_sc_hd__o32ai_4
X_63170_ _63053_/A _63170_/X sky130_fd_sc_hd__buf_2
X_75156_ _75151_/Y _75156_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_3_4_0_CLK clkbuf_2_2_2_CLK/X clkbuf_3_4_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_41548_ _41411_/X _41548_/X sky130_fd_sc_hd__buf_2
X_60382_ _60447_/A _60383_/A sky130_fd_sc_hd__buf_2
X_72368_ _72368_/A _72401_/B _72368_/Y sky130_fd_sc_hd__nor2_4
X_62121_ _61820_/A _62121_/X sky130_fd_sc_hd__buf_2
X_74107_ _72909_/A _74107_/X sky130_fd_sc_hd__buf_2
X_47055_ _86675_/Q _47050_/X _47054_/Y _47055_/Y sky130_fd_sc_hd__o21ai_4
X_71319_ _70428_/A _71319_/B _71320_/A sky130_fd_sc_hd__nor2_4
X_44267_ _44267_/A _44268_/A sky130_fd_sc_hd__inv_2
X_79964_ _79964_/A _79963_/Y _79964_/Y sky130_fd_sc_hd__nand2_4
X_75087_ _75086_/Y _75087_/Y sky130_fd_sc_hd__inv_2
X_41479_ _41478_/Y _41479_/X sky130_fd_sc_hd__buf_2
X_72299_ _59325_/A _72299_/X sky130_fd_sc_hd__buf_2
X_46006_ _46006_/A _46006_/Y sky130_fd_sc_hd__inv_2
X_43218_ _43218_/A _43218_/X sky130_fd_sc_hd__buf_2
X_62052_ _62050_/X _62090_/B _78060_/B _62052_/Y sky130_fd_sc_hd__nor3_4
X_78915_ _78903_/Y _82509_/D sky130_fd_sc_hd__inv_2
X_74038_ _74038_/A _85901_/Q _74038_/X sky130_fd_sc_hd__and2_4
X_44198_ _56953_/A _57043_/B sky130_fd_sc_hd__buf_2
X_79895_ _79895_/A _79895_/B _81090_/D sky130_fd_sc_hd__xnor2_4
X_61003_ _61003_/A _60865_/C _60865_/B _61003_/Y sky130_fd_sc_hd__nand3_4
X_43149_ _43017_/A _43149_/X sky130_fd_sc_hd__buf_2
X_66860_ _66625_/A _66912_/A sky130_fd_sc_hd__buf_2
X_78846_ _82839_/Q _82551_/Q _78857_/A sky130_fd_sc_hd__xor2_4
X_65811_ _65660_/A _65811_/X sky130_fd_sc_hd__buf_2
X_47957_ _47946_/A _47957_/B _47957_/X sky130_fd_sc_hd__and2_4
X_66791_ _66791_/A _66790_/X _66791_/Y sky130_fd_sc_hd__nand2_4
X_78777_ _78775_/Y _78777_/B _78778_/B sky130_fd_sc_hd__xor2_4
X_75989_ _75981_/A _75986_/A _75990_/B sky130_fd_sc_hd__and2_4
X_68530_ _68452_/A _68530_/B _68530_/X sky130_fd_sc_hd__and2_4
X_46908_ _46767_/A _46908_/X sky130_fd_sc_hd__buf_2
X_65742_ _65742_/A _65742_/B _65742_/Y sky130_fd_sc_hd__nand2_4
X_77728_ _77728_/A _77728_/B _77728_/X sky130_fd_sc_hd__xor2_4
X_62954_ _62950_/Y _62942_/X _62953_/Y _62954_/Y sky130_fd_sc_hd__a21oi_4
X_47888_ _47883_/Y _47846_/X _47887_/X _47888_/Y sky130_fd_sc_hd__a21oi_4
X_49627_ _49607_/X _52843_/B _49627_/Y sky130_fd_sc_hd__nand2_4
X_61905_ _61871_/A _61949_/B _61949_/C _63137_/B _61905_/X sky130_fd_sc_hd__and4_4
X_68461_ _68461_/A _68586_/A sky130_fd_sc_hd__buf_2
X_46839_ _46835_/Y _46798_/X _46838_/X _86698_/D sky130_fd_sc_hd__a21oi_4
X_65673_ _65673_/A _65825_/A sky130_fd_sc_hd__buf_2
X_77659_ _77660_/A _77656_/Y _77658_/Y _77693_/A sky130_fd_sc_hd__a21o_4
X_62885_ _63611_/A _62875_/X _62884_/Y _62885_/X sky130_fd_sc_hd__o21a_4
X_67412_ _86972_/Q _67311_/X _67313_/X _67411_/X _67413_/B sky130_fd_sc_hd__a211o_4
X_64624_ _64676_/A _85856_/Q _64624_/X sky130_fd_sc_hd__and2_4
X_49558_ _49558_/A _52773_/B _49558_/Y sky130_fd_sc_hd__nand2_4
X_61836_ _61834_/Y _61801_/X _61835_/Y _61836_/Y sky130_fd_sc_hd__a21oi_4
X_80670_ _80670_/CLK _80670_/D _80670_/Q sky130_fd_sc_hd__dfxtp_4
X_68392_ _68392_/A _69607_/A sky130_fd_sc_hd__buf_2
X_48509_ _48471_/X _47973_/A _48508_/Y _74431_/A sky130_fd_sc_hd__o21ai_4
X_67343_ _87923_/Q _67293_/X _67271_/X _67342_/X _67343_/X sky130_fd_sc_hd__a211o_4
X_79329_ _84800_/Q _84120_/Q _79331_/A sky130_fd_sc_hd__xor2_4
X_64555_ _64210_/A _64229_/X _64553_/Y _64554_/Y _64555_/Y sky130_fd_sc_hd__nand4_4
X_49489_ _49500_/A _49500_/B _49467_/C _52704_/D _49489_/X sky130_fd_sc_hd__and4_4
X_61767_ _61754_/X _61758_/X _61766_/Y _58154_/A _61719_/X _61767_/Y
+ sky130_fd_sc_hd__o32ai_4
X_51520_ _50946_/A _51629_/A sky130_fd_sc_hd__buf_2
X_63506_ _63495_/X _63496_/X _63499_/X _63503_/X _63505_/Y _63506_/Y
+ sky130_fd_sc_hd__o41ai_4
X_82340_ _82299_/CLK _77065_/X _48136_/A sky130_fd_sc_hd__dfxtp_4
X_60718_ _60707_/X _60709_/X _60820_/A _60714_/Y _60717_/Y _84581_/D
+ sky130_fd_sc_hd__a41oi_4
X_67274_ _66915_/A _67274_/X sky130_fd_sc_hd__buf_2
X_64486_ _61238_/C _64457_/C _64484_/Y _64485_/Y _64486_/Y sky130_fd_sc_hd__nand4_4
X_61698_ _61692_/Y _61694_/Y _61320_/Y _61695_/Y _61697_/Y _61698_/X
+ sky130_fd_sc_hd__a41o_4
X_69013_ _69009_/X _69012_/X _68922_/X _69013_/X sky130_fd_sc_hd__a21o_4
X_66225_ _65595_/X _66225_/X sky130_fd_sc_hd__buf_2
X_51451_ _51504_/A _51473_/B sky130_fd_sc_hd__buf_2
X_63437_ _63372_/A _63437_/X sky130_fd_sc_hd__buf_2
X_82271_ _82272_/CLK _82271_/D _82271_/Q sky130_fd_sc_hd__dfxtp_4
X_60649_ _60724_/B _60712_/B sky130_fd_sc_hd__buf_2
X_84010_ _84074_/CLK _68215_/X _82050_/D sky130_fd_sc_hd__dfxtp_4
X_50402_ _50399_/Y _50395_/X _50401_/X _86208_/D sky130_fd_sc_hd__a21oi_4
X_81222_ _85317_/CLK _81222_/D _81222_/Q sky130_fd_sc_hd__dfxtp_4
X_54170_ _85491_/Q _54167_/X _54169_/Y _54170_/Y sky130_fd_sc_hd__o21ai_4
X_66156_ _65300_/X _85616_/Q _44261_/X _66155_/X _66156_/X sky130_fd_sc_hd__a211o_4
X_51382_ _51364_/A _50870_/B _51382_/Y sky130_fd_sc_hd__nand2_4
X_63368_ _63368_/A _63368_/X sky130_fd_sc_hd__buf_2
X_53121_ _53147_/A _53121_/X sky130_fd_sc_hd__buf_2
X_65107_ _65104_/X _65106_/X _64959_/X _65107_/X sky130_fd_sc_hd__a21o_4
X_50333_ _50464_/A _50333_/X sky130_fd_sc_hd__buf_2
X_62319_ _62319_/A _63448_/B _62319_/C _62322_/C sky130_fd_sc_hd__nand3_4
X_81153_ _82284_/CLK _81153_/D _40558_/A sky130_fd_sc_hd__dfxtp_4
X_66087_ _66011_/X _66087_/B _66087_/X sky130_fd_sc_hd__and2_4
X_63299_ _58287_/Y _63250_/X _59430_/Y _60493_/A _63299_/X sky130_fd_sc_hd__o22a_4
X_80104_ _80117_/B _80103_/Y _80107_/A sky130_fd_sc_hd__xor2_4
X_53052_ _53048_/A _53063_/B _53058_/C _53052_/D _53052_/X sky130_fd_sc_hd__and4_4
X_65038_ _65035_/X _85553_/Q _65036_/X _65037_/X _65038_/X sky130_fd_sc_hd__a211o_4
X_69915_ _81959_/D _69894_/X _69914_/X _83887_/D sky130_fd_sc_hd__a21bo_4
X_50264_ _50251_/X _50264_/B _50264_/Y sky130_fd_sc_hd__nand2_4
X_85961_ _85961_/CLK _51706_/Y _85961_/Q sky130_fd_sc_hd__dfxtp_4
X_81084_ _81084_/CLK _75657_/A _81084_/Q sky130_fd_sc_hd__dfxtp_4
X_52003_ _51982_/X _50300_/B _52003_/Y sky130_fd_sc_hd__nand2_4
X_87700_ _87126_/CLK _42824_/X _68067_/B sky130_fd_sc_hd__dfxtp_4
X_80035_ _80013_/Y _80031_/X _80034_/Y _80035_/Y sky130_fd_sc_hd__a21oi_4
X_84912_ _84714_/CLK _84912_/D _58187_/A sky130_fd_sc_hd__dfxtp_4
X_57860_ _57824_/X _85496_/Q _57849_/X _57860_/X sky130_fd_sc_hd__o21a_4
X_69846_ _69832_/X _69844_/Y _69815_/X _69845_/Y _69846_/X sky130_fd_sc_hd__a211o_4
X_50195_ _50187_/X _50708_/B _50195_/Y sky130_fd_sc_hd__nand2_4
X_85892_ _86203_/CLK _85892_/D _74232_/B sky130_fd_sc_hd__dfxtp_4
X_56811_ _56713_/A _56810_/X _56811_/Y sky130_fd_sc_hd__nand2_4
X_87631_ _87888_/CLK _87631_/D _66676_/B sky130_fd_sc_hd__dfxtp_4
X_84843_ _84877_/CLK _84843_/D _84843_/Q sky130_fd_sc_hd__dfxtp_4
X_57791_ _57790_/X _57791_/X sky130_fd_sc_hd__buf_2
X_69777_ _68587_/X _69776_/Y _69777_/Y sky130_fd_sc_hd__nor2_4
X_66989_ _66942_/A _88194_/Q _66989_/X sky130_fd_sc_hd__and2_4
X_59530_ _59529_/X _61183_/A sky130_fd_sc_hd__buf_2
X_56742_ _56727_/X _56736_/X _56741_/Y _56742_/Y sky130_fd_sc_hd__o21ai_4
X_68728_ _69735_/A _68727_/Y _68728_/Y sky130_fd_sc_hd__nor2_4
X_87562_ _83158_/CLK _87562_/D _43137_/A sky130_fd_sc_hd__dfxtp_4
X_53954_ _53952_/Y _53948_/X _53953_/Y _85535_/D sky130_fd_sc_hd__a21boi_4
X_84774_ _86688_/CLK _84774_/D _84774_/Q sky130_fd_sc_hd__dfxtp_4
X_81986_ _82104_/CLK _81986_/D _81986_/Q sky130_fd_sc_hd__dfxtp_4
X_86513_ _85859_/CLK _48547_/Y _86513_/Q sky130_fd_sc_hd__dfxtp_4
X_52905_ _52910_/A _47184_/X _52905_/Y sky130_fd_sc_hd__nand2_4
X_59461_ _59442_/X _83462_/Q _59460_/Y _84726_/D sky130_fd_sc_hd__o21a_4
X_83725_ _85379_/CLK _83725_/D _47489_/A sky130_fd_sc_hd__dfxtp_4
X_56673_ _83328_/Q _57270_/A sky130_fd_sc_hd__buf_2
X_68659_ _87092_/Q _68580_/X _68630_/X _68658_/X _68659_/X sky130_fd_sc_hd__a211o_4
X_80937_ _80962_/CLK _80937_/D _80937_/Q sky130_fd_sc_hd__dfxtp_4
X_87493_ _88012_/CLK _43294_/X _87493_/Q sky130_fd_sc_hd__dfxtp_4
X_53885_ _53882_/Y _53829_/X _53884_/X _53885_/Y sky130_fd_sc_hd__a21oi_4
X_58412_ _58412_/A _58415_/B _58412_/Y sky130_fd_sc_hd__nand2_4
X_55624_ _55616_/X _55624_/B _55624_/X sky130_fd_sc_hd__and2_4
X_86444_ _86155_/CLK _86444_/D _65164_/B sky130_fd_sc_hd__dfxtp_4
X_40850_ _40835_/X _40836_/X _40849_/X _88323_/Q _40832_/X _40850_/Y
+ sky130_fd_sc_hd__o32ai_4
X_52836_ _52834_/Y _52809_/X _52835_/X _52836_/Y sky130_fd_sc_hd__a21oi_4
X_71670_ _71308_/A _71680_/A sky130_fd_sc_hd__buf_2
X_59392_ _59392_/A _58988_/B _59392_/Y sky130_fd_sc_hd__nand2_4
X_83656_ _85536_/CLK _70943_/Y _83656_/Q sky130_fd_sc_hd__dfxtp_4
X_80868_ _81125_/CLK _75597_/B _80868_/Q sky130_fd_sc_hd__dfxtp_4
X_70621_ _52999_/B _70583_/X _70620_/Y _83739_/D sky130_fd_sc_hd__o21ai_4
X_58343_ _84873_/Q _58344_/A sky130_fd_sc_hd__buf_2
X_82607_ _82575_/CLK _78927_/B _82607_/Q sky130_fd_sc_hd__dfxtp_4
X_55555_ _55524_/A _55555_/B _55555_/Y sky130_fd_sc_hd__nor2_4
X_86375_ _83663_/CLK _86375_/D _58896_/B sky130_fd_sc_hd__dfxtp_4
X_52767_ _52767_/A _52773_/A sky130_fd_sc_hd__buf_2
X_40781_ _40780_/Y _40781_/X sky130_fd_sc_hd__buf_2
X_83587_ _85593_/CLK _83587_/D _83587_/Q sky130_fd_sc_hd__dfxtp_4
X_80799_ _80817_/CLK _75855_/Y _75533_/B sky130_fd_sc_hd__dfxtp_4
X_88114_ _87834_/CLK _88114_/D _88114_/Q sky130_fd_sc_hd__dfxtp_4
X_54506_ _85429_/Q _54485_/X _54505_/Y _54506_/Y sky130_fd_sc_hd__o21ai_4
X_42520_ _42517_/X _42501_/X _40716_/X _42518_/Y _42519_/X _87836_/D
+ sky130_fd_sc_hd__o32ai_4
X_73340_ _83155_/Q _73318_/X _73339_/Y _83155_/D sky130_fd_sc_hd__a21o_4
X_85326_ _83550_/CLK _85326_/D _85326_/Q sky130_fd_sc_hd__dfxtp_4
X_51718_ _85958_/Q _51701_/X _51717_/Y _51718_/Y sky130_fd_sc_hd__o21ai_4
X_70552_ DATA_TO_HASH[4] _70552_/Y sky130_fd_sc_hd__inv_2
X_58274_ _58274_/A _58280_/B _58274_/Y sky130_fd_sc_hd__nand2_4
X_82538_ _82538_/CLK _82538_/D _79020_/B sky130_fd_sc_hd__dfxtp_4
X_55486_ _55482_/X _55485_/X _44112_/X _55491_/A sky130_fd_sc_hd__a21o_4
X_52698_ _52674_/X _52694_/B _52694_/C _52698_/D _52698_/X sky130_fd_sc_hd__and4_4
X_57225_ _56852_/A _57193_/D _57225_/Y sky130_fd_sc_hd__nor2_4
X_42451_ _42579_/A _42488_/A sky130_fd_sc_hd__buf_2
X_88045_ _88084_/CLK _42075_/X _88045_/Q sky130_fd_sc_hd__dfxtp_4
X_54437_ _54446_/A _52744_/B _54437_/Y sky130_fd_sc_hd__nand2_4
X_73271_ _73269_/X _73270_/Y _73221_/X _73271_/Y sky130_fd_sc_hd__a21oi_4
X_85257_ _85257_/CLK _56257_/Y _85257_/Q sky130_fd_sc_hd__dfxtp_4
X_51649_ _51671_/A _53174_/B _51649_/Y sky130_fd_sc_hd__nand2_4
X_70483_ _71706_/A _70483_/B _71435_/C _70483_/X sky130_fd_sc_hd__and3_4
X_82469_ _82924_/CLK _82469_/D _78273_/B sky130_fd_sc_hd__dfxtp_4
X_75010_ _75008_/X _75021_/B _75010_/Y sky130_fd_sc_hd__nand2_4
X_41402_ _41373_/X _82891_/Q _41401_/X _41402_/X sky130_fd_sc_hd__o21a_4
X_72222_ _72172_/X _72220_/Y _72221_/Y _72189_/X _72176_/X _72222_/X
+ sky130_fd_sc_hd__o32a_4
X_84208_ _85315_/CLK _84208_/D _65268_/C sky130_fd_sc_hd__dfxtp_4
X_45170_ _45167_/X _45169_/Y _45125_/X _45170_/Y sky130_fd_sc_hd__a21oi_4
X_57156_ _57129_/Y _57156_/X sky130_fd_sc_hd__buf_2
X_54368_ _54365_/Y _54366_/X _54367_/X _54368_/Y sky130_fd_sc_hd__a21oi_4
X_42382_ _42382_/A _87892_/D sky130_fd_sc_hd__inv_2
X_85188_ _85186_/CLK _56453_/Y _56452_/C sky130_fd_sc_hd__dfxtp_4
X_56107_ _55802_/X _55811_/X _56108_/B sky130_fd_sc_hd__and2_4
X_44121_ _44120_/Y _44196_/A sky130_fd_sc_hd__buf_2
X_41333_ _41235_/X _41333_/X sky130_fd_sc_hd__buf_2
X_53319_ _85655_/Q _53295_/X _53318_/Y _53319_/Y sky130_fd_sc_hd__o21ai_4
X_72153_ _59292_/X _85342_/Q _59365_/X _72153_/X sky130_fd_sc_hd__o21a_4
X_84139_ _82746_/CLK _84139_/D _84139_/Q sky130_fd_sc_hd__dfxtp_4
X_57087_ _57086_/X _57087_/X sky130_fd_sc_hd__buf_2
X_54299_ _54297_/Y _54285_/X _54298_/X _54299_/Y sky130_fd_sc_hd__a21oi_4
X_71104_ _71101_/X _71080_/B _71099_/C _71104_/Y sky130_fd_sc_hd__nand3_4
X_44052_ _44052_/A _44052_/X sky130_fd_sc_hd__buf_2
X_56038_ _56029_/X _56035_/X _56037_/Y _85307_/D sky130_fd_sc_hd__o21ai_4
X_41264_ _41264_/A _41264_/X sky130_fd_sc_hd__buf_2
X_72084_ _72075_/A _53910_/A _72084_/Y sky130_fd_sc_hd__nand2_4
X_76961_ _76828_/Y _76961_/Y sky130_fd_sc_hd__inv_2
X_43003_ _40524_/X _42994_/X _87609_/Q _42995_/X _87609_/D sky130_fd_sc_hd__a2bb2o_4
X_78700_ _78700_/A _78700_/Y sky130_fd_sc_hd__inv_2
X_71035_ _70786_/A _71181_/A sky130_fd_sc_hd__buf_2
X_75912_ _61192_/C _75912_/B _75912_/X sky130_fd_sc_hd__xor2_4
X_48860_ _48857_/Y _48840_/X _48859_/X _48860_/Y sky130_fd_sc_hd__a21oi_4
X_79680_ _79680_/A _84246_/Q _79681_/B sky130_fd_sc_hd__xor2_4
X_41195_ _41112_/X _41113_/X _41193_/X _68763_/B _41194_/X _41196_/A
+ sky130_fd_sc_hd__o32ai_4
X_76892_ _76884_/X _81500_/Q _76893_/A sky130_fd_sc_hd__and2_4
X_47811_ _86595_/Q _47806_/X _47810_/Y _47811_/Y sky130_fd_sc_hd__o21ai_4
X_78631_ _78630_/Y _78632_/C sky130_fd_sc_hd__inv_2
X_75843_ _75842_/Y _75843_/Y sky130_fd_sc_hd__inv_2
X_87829_ _87826_/CLK _87829_/D _87829_/Q sky130_fd_sc_hd__dfxtp_4
X_48791_ _48533_/A _48770_/X _48814_/C _48791_/X sky130_fd_sc_hd__and3_4
X_57989_ _58631_/A _57989_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_552_0_CLK clkbuf_9_276_0_CLK/X _88175_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_43_0_CLK clkbuf_6_43_0_CLK/A clkbuf_7_87_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_47742_ _47741_/Y _53219_/B sky130_fd_sc_hd__buf_2
X_59728_ _59689_/B _59689_/A _59666_/A _59728_/Y sky130_fd_sc_hd__a21oi_4
X_78562_ _78533_/X _78536_/X _78561_/Y _78562_/X sky130_fd_sc_hd__o21a_4
X_44954_ _44905_/X _61364_/B _44907_/X _44954_/Y sky130_fd_sc_hd__o21ai_4
X_75774_ _75761_/Y _75762_/Y _75773_/X _75774_/Y sky130_fd_sc_hd__a21oi_4
X_72986_ _73181_/A _85881_/Q _72986_/X sky130_fd_sc_hd__and2_4
X_77513_ _77502_/A _77501_/Y _77495_/Y _77514_/B sky130_fd_sc_hd__o21ai_4
X_43905_ _41352_/X _43886_/X _67616_/B _43887_/X _87207_/D sky130_fd_sc_hd__a2bb2o_4
X_74725_ _74723_/X _83794_/Q _74745_/D _74730_/B sky130_fd_sc_hd__nand3_4
X_47673_ _49379_/A _47692_/A sky130_fd_sc_hd__buf_2
X_71937_ _56816_/Y _71917_/X _71936_/Y _71937_/Y sky130_fd_sc_hd__o21ai_4
X_59659_ _59582_/B _59660_/D sky130_fd_sc_hd__buf_2
X_78493_ _78491_/X _78492_/Y _78494_/A sky130_fd_sc_hd__and2_4
X_44885_ _85185_/Q _44882_/X _44884_/X _44885_/X sky130_fd_sc_hd__o21a_4
X_49412_ _49493_/A _49420_/C sky130_fd_sc_hd__buf_2
X_46624_ _46624_/A _46624_/Y sky130_fd_sc_hd__inv_2
X_77444_ _77444_/A _77444_/B _77444_/Y sky130_fd_sc_hd__nor2_4
X_43836_ _41161_/X _43832_/X _68604_/B _43833_/X _43836_/X sky130_fd_sc_hd__a2bb2o_4
X_62670_ _62659_/Y _62660_/X _62661_/Y _62664_/Y _62669_/X _62670_/X
+ sky130_fd_sc_hd__a41o_4
X_74656_ _74685_/C _74656_/X sky130_fd_sc_hd__buf_2
X_71868_ _71847_/Y _83346_/Q _71867_/Y _83346_/D sky130_fd_sc_hd__a21o_4
Xclkbuf_10_567_0_CLK clkbuf_9_283_0_CLK/X _86807_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_58_0_CLK clkbuf_6_59_0_CLK/A clkbuf_6_58_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_49343_ _49341_/Y _49326_/X _49342_/Y _49343_/Y sky130_fd_sc_hd__a21boi_4
X_61621_ _84873_/Q _61323_/B _61621_/X sky130_fd_sc_hd__or2_4
X_73607_ _73607_/A _65932_/B _73607_/X sky130_fd_sc_hd__and2_4
X_70819_ _70819_/A _70952_/B sky130_fd_sc_hd__buf_2
X_46555_ _54073_/B _50862_/B sky130_fd_sc_hd__buf_2
X_77375_ _81932_/Q _82188_/D _77375_/X sky130_fd_sc_hd__xor2_4
X_43767_ _43005_/X _43760_/X _40977_/X _87275_/Q _43756_/X _43767_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74587_ _74549_/A _46228_/A _45156_/A _74587_/Y sky130_fd_sc_hd__nand3_4
X_40979_ _40978_/Y _40979_/Y sky130_fd_sc_hd__inv_2
X_71799_ _58209_/Y _71783_/Y _71798_/Y _83371_/D sky130_fd_sc_hd__o21ai_4
X_79114_ _79114_/A _79113_/Y _79114_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_1_1_2_CLK clkbuf_1_1_1_CLK/X clkbuf_2_3_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_45506_ _45502_/X _45505_/X _45446_/X _45506_/X sky130_fd_sc_hd__a21o_4
X_64340_ _79775_/B _64314_/X _64339_/X _64340_/X sky130_fd_sc_hd__a21o_4
X_76326_ _81358_/Q _76326_/B _76326_/X sky130_fd_sc_hd__xor2_4
X_42718_ _42681_/A _42718_/X sky130_fd_sc_hd__buf_2
X_49274_ _49270_/Y _49271_/X _49273_/Y _49274_/Y sky130_fd_sc_hd__a21boi_4
X_61552_ _58442_/A _61563_/B _61563_/C _61514_/D _61553_/A sky130_fd_sc_hd__nand4_4
X_73538_ _72829_/A _85570_/Q _73472_/X _73537_/X _73538_/X sky130_fd_sc_hd__a211o_4
X_46486_ _46485_/X _46487_/B sky130_fd_sc_hd__buf_2
X_43698_ _47834_/A _43698_/X sky130_fd_sc_hd__buf_2
X_48225_ _66041_/B _48203_/X _48224_/Y _48225_/Y sky130_fd_sc_hd__o21ai_4
X_60503_ _60502_/Y _60503_/X sky130_fd_sc_hd__buf_2
X_79045_ _79057_/A _79044_/Y _79045_/X sky130_fd_sc_hd__and2_4
X_45437_ _45428_/X _45432_/X _45436_/Y _45437_/Y sky130_fd_sc_hd__a21oi_4
X_64271_ _79837_/B _64255_/X _64270_/X _64271_/X sky130_fd_sc_hd__a21o_4
X_76257_ _76242_/Y _76236_/X _76237_/Y _76257_/Y sky130_fd_sc_hd__a21boi_4
X_42649_ _42647_/X _42648_/X _40977_/X _87787_/Q _42637_/X _42649_/Y
+ sky130_fd_sc_hd__o32ai_4
X_61483_ _61483_/A _61468_/B _61467_/X _61451_/D _61483_/Y sky130_fd_sc_hd__nand4_4
X_73469_ _87043_/Q _56550_/X _73468_/X _73481_/C sky130_fd_sc_hd__o21ai_4
X_66010_ _66007_/X _66009_/X _65937_/X _66010_/X sky130_fd_sc_hd__a21o_4
X_63222_ _79321_/A _63189_/X _63221_/Y _63222_/X sky130_fd_sc_hd__a21o_4
X_75208_ _75205_/Y _75207_/Y _75217_/B sky130_fd_sc_hd__nand2_4
X_60434_ _60516_/B _60435_/C sky130_fd_sc_hd__buf_2
X_48156_ _48734_/A _48156_/X sky130_fd_sc_hd__buf_2
X_45368_ _56670_/A _45369_/A sky130_fd_sc_hd__buf_2
X_76188_ _76189_/A _76187_/Y _76189_/B _76188_/X sky130_fd_sc_hd__a21o_4
X_47107_ _83701_/Q _53373_/B sky130_fd_sc_hd__inv_2
X_44319_ _43951_/B _44316_/X _44313_/A _44218_/X _44320_/A sky130_fd_sc_hd__o22a_4
X_63153_ _58554_/A _63131_/X _63117_/X _58331_/A _63118_/X _63153_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75139_ _75138_/Y _75142_/A sky130_fd_sc_hd__inv_2
X_48087_ _48075_/X _46528_/A _48086_/X _48088_/B sky130_fd_sc_hd__o21ai_4
X_60365_ _60477_/A _60519_/B _79581_/A _60365_/Y sky130_fd_sc_hd__nor3_4
X_45299_ _85255_/Q _45297_/X _45298_/X _45299_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_505_0_CLK clkbuf_9_252_0_CLK/X _83681_/CLK sky130_fd_sc_hd__clkbuf_1
X_62104_ _62037_/X _62021_/B _63655_/B _62020_/X _62104_/X sky130_fd_sc_hd__and4_4
X_47038_ _54509_/D _52818_/D sky130_fd_sc_hd__buf_2
X_63084_ _58429_/Y _63073_/X _63059_/X _59474_/A _63060_/X _63084_/Y
+ sky130_fd_sc_hd__o32ai_4
X_67961_ _67961_/A _67960_/X _67961_/Y sky130_fd_sc_hd__nand2_4
X_79947_ _79944_/Y _79946_/Y _79947_/Y sky130_fd_sc_hd__nand2_4
X_60296_ _60267_/A _60296_/X sky130_fd_sc_hd__buf_2
X_69700_ _69908_/A _69700_/B _69700_/Y sky130_fd_sc_hd__nor2_4
X_66912_ _66912_/A _87621_/Q _66912_/X sky130_fd_sc_hd__and2_4
X_62035_ _62031_/Y _62033_/X _62034_/Y _62035_/Y sky130_fd_sc_hd__a21oi_4
X_67892_ _87452_/Q _67868_/X _67821_/X _67891_/X _67892_/X sky130_fd_sc_hd__a211o_4
X_79878_ _79875_/Y _79858_/Y _79877_/X _79878_/Y sky130_fd_sc_hd__o21ai_4
X_69631_ _81981_/D _69564_/X _69630_/X _83909_/D sky130_fd_sc_hd__a21bo_4
X_66843_ _66606_/A _66843_/X sky130_fd_sc_hd__buf_2
X_78829_ _78829_/A _78828_/Y _78829_/Y sky130_fd_sc_hd__nand2_4
X_48989_ _48908_/A _53834_/B _48989_/X sky130_fd_sc_hd__and2_4
X_69562_ _69505_/X _46199_/X _69560_/Y _69561_/Y _69562_/X sky130_fd_sc_hd__a211o_4
X_81840_ _81857_/CLK _81840_/D _77423_/A sky130_fd_sc_hd__dfxtp_4
X_66774_ _66819_/A _86830_/Q _66774_/X sky130_fd_sc_hd__and2_4
X_63986_ _60909_/X _64050_/C sky130_fd_sc_hd__buf_2
X_68513_ _68507_/X _68511_/X _68512_/X _68513_/Y sky130_fd_sc_hd__a21oi_4
X_65725_ _65721_/X _65725_/B _65724_/X _65725_/Y sky130_fd_sc_hd__nand3_4
X_50951_ _86101_/Q _50936_/X _50950_/Y _50951_/Y sky130_fd_sc_hd__o21ai_4
X_62937_ _60291_/C _62982_/C sky130_fd_sc_hd__buf_2
X_81771_ _83987_/CLK _81771_/D _81771_/Q sky130_fd_sc_hd__dfxtp_4
X_69493_ _88025_/Q _69315_/X _69393_/X _69492_/X _69493_/X sky130_fd_sc_hd__a211o_4
X_83510_ _83507_/CLK _71407_/X _83510_/Q sky130_fd_sc_hd__dfxtp_4
X_80722_ _81084_/CLK _75908_/X _80690_/D sky130_fd_sc_hd__dfxtp_4
X_68444_ _68444_/A _88368_/Q _68444_/X sky130_fd_sc_hd__and2_4
X_53670_ _85591_/Q _53660_/X _53669_/Y _53670_/Y sky130_fd_sc_hd__o21ai_4
X_65656_ _65654_/X _86194_/Q _65576_/X _65655_/X _65656_/X sky130_fd_sc_hd__a211o_4
X_84490_ _84649_/CLK _61275_/Y _84490_/Q sky130_fd_sc_hd__dfxtp_4
X_50882_ _50819_/X _50882_/X sky130_fd_sc_hd__buf_2
X_62868_ _60273_/A _62935_/B sky130_fd_sc_hd__buf_2
X_52621_ _52648_/A _52643_/A sky130_fd_sc_hd__buf_2
X_64607_ _60109_/A _64608_/A sky130_fd_sc_hd__buf_2
X_83441_ _83338_/CLK _83441_/D _83441_/Q sky130_fd_sc_hd__dfxtp_4
X_61819_ _62851_/A _61820_/A sky130_fd_sc_hd__buf_2
X_80653_ _86772_/CLK _80653_/D _80653_/Q sky130_fd_sc_hd__dfxtp_4
X_68375_ _83977_/Q _68338_/X _68374_/X _83977_/D sky130_fd_sc_hd__a21bo_4
X_65587_ _65587_/A _65587_/B _65587_/Y sky130_fd_sc_hd__nand2_4
X_62799_ _62773_/X _62762_/B _61922_/X _62799_/Y sky130_fd_sc_hd__nand3_4
X_55340_ _55336_/X _83752_/Q _55365_/B _55445_/D sky130_fd_sc_hd__nand3_4
X_67326_ _67323_/X _67325_/X _67255_/X _67326_/Y sky130_fd_sc_hd__a21oi_4
X_86160_ _83306_/CLK _50653_/Y _86160_/Q sky130_fd_sc_hd__dfxtp_4
X_52552_ _65270_/B _52549_/X _52551_/Y _52552_/Y sky130_fd_sc_hd__o21ai_4
X_64538_ _58987_/Y _64226_/X _64537_/Y _64538_/Y sky130_fd_sc_hd__o21ai_4
X_83372_ _83372_/CLK _71797_/Y _83372_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_307 sky130_fd_sc_hd__decap_3
X_80584_ _80581_/X _80584_/B _82269_/D sky130_fd_sc_hd__xor2_4
XPHY_318 sky130_fd_sc_hd__decap_3
XPHY_329 sky130_fd_sc_hd__decap_3
X_85111_ _85089_/CLK _85111_/D _45549_/A sky130_fd_sc_hd__dfxtp_4
X_51503_ _51557_/A _51503_/X sky130_fd_sc_hd__buf_2
X_82323_ _82103_/CLK _77123_/B _82323_/Q sky130_fd_sc_hd__dfxtp_4
X_55271_ _55268_/X _55270_/X _44109_/X _55285_/A sky130_fd_sc_hd__a21o_4
X_67257_ _67141_/X _67247_/Y _67152_/X _67256_/Y _67257_/X sky130_fd_sc_hd__a211o_4
X_86091_ _86091_/CLK _86091_/D _86091_/Q sky130_fd_sc_hd__dfxtp_4
X_52483_ _52481_/Y _52462_/X _52482_/Y _52483_/Y sky130_fd_sc_hd__a21boi_4
X_64469_ _58274_/A _64423_/X _64468_/Y _64469_/Y sky130_fd_sc_hd__o21ai_4
X_57010_ _57010_/A _57010_/Y sky130_fd_sc_hd__inv_2
X_54222_ _54250_/A _54230_/A sky130_fd_sc_hd__buf_2
X_66208_ _65752_/X _66195_/B _65754_/X _66217_/A sky130_fd_sc_hd__nand3_4
X_85042_ _85042_/CLK _85042_/D _85042_/Q sky130_fd_sc_hd__dfxtp_4
X_51434_ _51432_/Y _51420_/X _51433_/X _86011_/D sky130_fd_sc_hd__a21oi_4
X_82254_ _85332_/CLK _80429_/X _82254_/Q sky130_fd_sc_hd__dfxtp_4
X_67188_ _67095_/A _67188_/B _67188_/X sky130_fd_sc_hd__and2_4
X_81205_ _84981_/CLK _75037_/X _49009_/A sky130_fd_sc_hd__dfxtp_4
X_54153_ _54149_/A _47324_/A _54153_/Y sky130_fd_sc_hd__nand2_4
X_66139_ _66164_/A _66164_/B _66138_/Y _66139_/Y sky130_fd_sc_hd__nor3_4
X_51365_ _65260_/B _51362_/X _51364_/Y _51365_/Y sky130_fd_sc_hd__o21ai_4
X_82185_ _84951_/CLK _82185_/D _82185_/Q sky130_fd_sc_hd__dfxtp_4
X_53104_ _53102_/Y _53082_/X _53103_/X _53104_/Y sky130_fd_sc_hd__a21oi_4
X_50316_ _50219_/X _50316_/X sky130_fd_sc_hd__buf_2
X_81136_ _80818_/CLK _81136_/D _81136_/Q sky130_fd_sc_hd__dfxtp_4
X_58961_ _58877_/A _58961_/X sky130_fd_sc_hd__buf_2
X_54084_ _54082_/Y _53472_/X _54083_/Y _85508_/D sky130_fd_sc_hd__a21boi_4
X_51296_ _51296_/A _49265_/B _51296_/Y sky130_fd_sc_hd__nand2_4
X_86993_ _86998_/CLK _86993_/D _86993_/Q sky130_fd_sc_hd__dfxtp_4
X_53035_ _53062_/A _53058_/C sky130_fd_sc_hd__buf_2
X_57912_ _84940_/Q _57912_/Y sky130_fd_sc_hd__inv_2
X_50247_ _53190_/A _50247_/X sky130_fd_sc_hd__buf_2
X_85944_ _82774_/CLK _85944_/D _85944_/Q sky130_fd_sc_hd__dfxtp_4
X_81067_ _83944_/CLK _81099_/Q _75201_/B sky130_fd_sc_hd__dfxtp_4
X_58892_ _58813_/X _85768_/Q _58838_/X _58892_/X sky130_fd_sc_hd__o21a_4
X_80018_ _84659_/Q _64100_/C _80018_/X sky130_fd_sc_hd__xor2_4
X_57843_ _57806_/X _86329_/Q _57843_/Y sky130_fd_sc_hd__nor2_4
X_69829_ _69403_/Y _69732_/X _69815_/X _69828_/Y _69829_/X sky130_fd_sc_hd__a211o_4
X_50178_ _65249_/B _50162_/X _50177_/Y _50178_/Y sky130_fd_sc_hd__o21ai_4
X_85875_ _86191_/CLK _52172_/Y _85875_/Q sky130_fd_sc_hd__dfxtp_4
X_87614_ _88128_/CLK _87614_/D _87614_/Q sky130_fd_sc_hd__dfxtp_4
X_72840_ _73535_/A _72840_/B _72840_/X sky130_fd_sc_hd__and2_4
X_84826_ _84829_/CLK _84826_/D _84826_/Q sky130_fd_sc_hd__dfxtp_4
X_57774_ _57773_/X _85725_/Q _44177_/X _57774_/X sky130_fd_sc_hd__o21a_4
X_54986_ _85340_/Q _54967_/X _54985_/Y _54986_/Y sky130_fd_sc_hd__o21ai_4
X_59513_ _43970_/A _59876_/B sky130_fd_sc_hd__buf_2
X_56725_ _57153_/A _56725_/B _56725_/Y sky130_fd_sc_hd__nand2_4
X_41951_ _42024_/A _41951_/X sky130_fd_sc_hd__buf_2
X_87545_ _87824_/CLK _43193_/Y _87545_/Q sky130_fd_sc_hd__dfxtp_4
X_53937_ _85538_/Q _53869_/X _53936_/Y _53937_/Y sky130_fd_sc_hd__o21ai_4
X_72771_ _72771_/A _72924_/B sky130_fd_sc_hd__buf_2
X_84757_ _84757_/CLK _59252_/Y _84757_/Q sky130_fd_sc_hd__dfxtp_4
X_81969_ _82558_/CLK _81969_/D _81969_/Q sky130_fd_sc_hd__dfxtp_4
X_74510_ _74508_/Y _74492_/X _74509_/X _74510_/Y sky130_fd_sc_hd__a21oi_4
X_40902_ _40877_/X _82855_/Q _40901_/X _40903_/A sky130_fd_sc_hd__o21ai_4
X_71722_ _58224_/Y _71718_/X _71721_/Y _83399_/D sky130_fd_sc_hd__o21ai_4
X_59444_ _59398_/A _59444_/X sky130_fd_sc_hd__buf_2
X_83708_ _83707_/CLK _83708_/D _83708_/Q sky130_fd_sc_hd__dfxtp_4
X_56656_ _83331_/Q _83330_/Q _56912_/A sky130_fd_sc_hd__nand2_4
X_44670_ _44669_/Y _87007_/D sky130_fd_sc_hd__inv_2
X_75490_ _75488_/Y _75491_/C _75491_/B _75493_/A sky130_fd_sc_hd__a21oi_4
X_87476_ _87749_/CLK _87476_/D _87476_/Q sky130_fd_sc_hd__dfxtp_4
X_53868_ _53866_/Y _53829_/X _53867_/X _53868_/Y sky130_fd_sc_hd__a21oi_4
X_41882_ _42000_/A _41882_/X sky130_fd_sc_hd__buf_2
X_84688_ _84329_/CLK _59854_/Y _84688_/Q sky130_fd_sc_hd__dfxtp_4
X_55607_ _55607_/A _45422_/Y _55607_/Y sky130_fd_sc_hd__nor2_4
X_43621_ _40640_/X _43609_/X _43620_/Y _43611_/X _43622_/A sky130_fd_sc_hd__a2bb2o_4
X_74441_ _72001_/A _74441_/X sky130_fd_sc_hd__buf_2
X_86427_ _86139_/CLK _86427_/D _64784_/B sky130_fd_sc_hd__dfxtp_4
X_40833_ _40758_/X _40759_/X _40831_/X _69740_/B _40832_/X _40833_/Y
+ sky130_fd_sc_hd__o32ai_4
X_52819_ _52814_/Y _52809_/X _52818_/X _52819_/Y sky130_fd_sc_hd__a21oi_4
X_83639_ _86127_/CLK _83639_/D _83639_/Q sky130_fd_sc_hd__dfxtp_4
X_59375_ _59364_/Y _59230_/X _59371_/X _59374_/X _84747_/D sky130_fd_sc_hd__a22oi_4
X_71653_ _58504_/Y _71649_/X _71652_/Y _71653_/Y sky130_fd_sc_hd__o21ai_4
X_56587_ _56764_/B _56587_/X sky130_fd_sc_hd__buf_2
X_53799_ _53838_/A _53799_/X sky130_fd_sc_hd__buf_2
X_46340_ _46288_/A _53978_/B _46340_/Y sky130_fd_sc_hd__nand2_4
X_70604_ _52979_/B _70584_/X _70603_/Y _83743_/D sky130_fd_sc_hd__o21ai_4
X_58326_ _58326_/A _58326_/B _58326_/Y sky130_fd_sc_hd__nand2_4
X_77160_ _77173_/A _77159_/Y _77161_/B sky130_fd_sc_hd__xor2_4
X_43552_ _43542_/X _43546_/X _40459_/X _87364_/Q _43549_/X _43553_/A
+ sky130_fd_sc_hd__o32ai_4
X_55538_ _45535_/A _55510_/X _44048_/X _55537_/Y _55538_/X sky130_fd_sc_hd__a211o_4
X_74372_ _74369_/Y _74370_/X _74371_/X _74372_/Y sky130_fd_sc_hd__a21oi_4
X_86358_ _86359_/CLK _86358_/D _86358_/Q sky130_fd_sc_hd__dfxtp_4
X_40764_ _40764_/A _88340_/D sky130_fd_sc_hd__inv_2
X_71584_ _71581_/X _83449_/Q _71583_/Y _83449_/D sky130_fd_sc_hd__a21o_4
X_76111_ _76107_/Y _76099_/B _76110_/X _76112_/B sky130_fd_sc_hd__o21ai_4
X_42503_ _42486_/X _42501_/X _40678_/X _42502_/Y _42489_/X _87843_/D
+ sky130_fd_sc_hd__o32ai_4
X_73323_ _73323_/A _73577_/B _73323_/Y sky130_fd_sc_hd__nor2_4
X_85309_ _85213_/CLK _85309_/D _56027_/C sky130_fd_sc_hd__dfxtp_4
X_46271_ _53951_/B _50738_/B sky130_fd_sc_hd__buf_2
X_70535_ _70534_/Y _71626_/A sky130_fd_sc_hd__buf_2
X_58257_ _58253_/X _83448_/Q _58256_/Y _58257_/X sky130_fd_sc_hd__o21a_4
X_77091_ _81998_/Q _81910_/Q _77091_/Y sky130_fd_sc_hd__nand2_4
X_43483_ _41697_/X _43465_/X _87399_/Q _43467_/X _87399_/D sky130_fd_sc_hd__a2bb2o_4
X_55469_ _44047_/X _55469_/X sky130_fd_sc_hd__buf_2
X_86289_ _86289_/CLK _86289_/D _86289_/Q sky130_fd_sc_hd__dfxtp_4
X_40695_ _40670_/X _40864_/A _40694_/X _40695_/Y sky130_fd_sc_hd__o21ai_4
X_48010_ _47867_/X _46436_/A _48009_/Y _48011_/A sky130_fd_sc_hd__o21ai_4
X_45222_ _45297_/A _45222_/X sky130_fd_sc_hd__buf_2
X_76042_ _81714_/D _76042_/B _76042_/Y sky130_fd_sc_hd__nand2_4
X_57208_ _57196_/Y _57055_/A _57208_/Y sky130_fd_sc_hd__nand2_4
X_88028_ _87767_/CLK _88028_/D _88028_/Q sky130_fd_sc_hd__dfxtp_4
X_42434_ _42373_/X _42434_/X sky130_fd_sc_hd__buf_2
X_73254_ _73248_/X _73253_/X _73200_/X _73270_/B sky130_fd_sc_hd__a21o_4
X_70466_ _70458_/X _70466_/Y sky130_fd_sc_hd__inv_2
X_58188_ _58187_/X _58184_/B _58188_/Y sky130_fd_sc_hd__nor2_4
X_72205_ _86618_/Q _72193_/B _72205_/Y sky130_fd_sc_hd__nor2_4
X_45153_ _45153_/A _45153_/X sky130_fd_sc_hd__buf_2
X_57139_ _56696_/A _57153_/B _57138_/Y _85073_/D sky130_fd_sc_hd__a21oi_4
X_42365_ _42365_/A _87899_/D sky130_fd_sc_hd__inv_2
X_73185_ _73182_/X _73184_/X _73067_/A _73188_/A sky130_fd_sc_hd__a21o_4
X_70397_ _70942_/A _74529_/A _70407_/C _70397_/Y sky130_fd_sc_hd__nand3_4
X_44104_ _44104_/A _44104_/Y sky130_fd_sc_hd__inv_2
X_79801_ _79793_/A _79793_/B _79800_/X _79801_/Y sky130_fd_sc_hd__o21ai_4
X_41316_ _41316_/A _41316_/X sky130_fd_sc_hd__buf_2
X_60150_ _60150_/A _65198_/A sky130_fd_sc_hd__buf_2
X_72136_ _83280_/Q _72115_/X _72130_/X _72135_/X _83280_/D sky130_fd_sc_hd__a2bb2oi_4
X_49961_ _48171_/X _49981_/A sky130_fd_sc_hd__buf_2
X_45084_ _64343_/B _61460_/B sky130_fd_sc_hd__buf_2
X_42296_ _41570_/X _42290_/X _87934_/Q _42291_/X _87934_/D sky130_fd_sc_hd__a2bb2o_4
X_77993_ _77993_/A _77993_/B _77994_/B sky130_fd_sc_hd__xor2_4
X_48912_ _48901_/A _48912_/B _48912_/Y sky130_fd_sc_hd__nand2_4
X_44035_ _65614_/A _59297_/A sky130_fd_sc_hd__buf_4
X_79732_ _84219_/Q _83267_/Q _79732_/X sky130_fd_sc_hd__xor2_4
X_41247_ _41246_/Y _41247_/Y sky130_fd_sc_hd__inv_2
X_60081_ _60081_/A _60081_/B _80082_/A _60081_/Y sky130_fd_sc_hd__nor3_4
X_72067_ _57563_/X _72068_/A sky130_fd_sc_hd__buf_2
X_76944_ _76941_/Y _76944_/B _81568_/D sky130_fd_sc_hd__nor2_4
X_49892_ _72128_/B _49880_/X _49891_/Y _49892_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_491_0_CLK clkbuf_9_245_0_CLK/X _85957_/CLK sky130_fd_sc_hd__clkbuf_1
X_71018_ _71168_/A _70620_/B _70925_/X _71018_/D _71018_/Y sky130_fd_sc_hd__nand4_4
X_48843_ _48851_/A _48843_/B _48843_/Y sky130_fd_sc_hd__nand2_4
X_79663_ _79647_/X _79664_/A _79663_/X sky130_fd_sc_hd__or2_4
X_41178_ _41143_/X _40659_/A _41177_/X _41178_/Y sky130_fd_sc_hd__o21ai_4
X_76875_ _76873_/Y _76874_/Y _76910_/C sky130_fd_sc_hd__xor2_4
X_78614_ _78617_/B _78614_/Y sky130_fd_sc_hd__inv_2
X_75826_ _75824_/A _81021_/Q _75824_/B _75827_/B sky130_fd_sc_hd__nand3_4
X_63840_ _61398_/B _63790_/X _63840_/C _63776_/X _63840_/Y sky130_fd_sc_hd__nand4_4
X_48774_ _65612_/B _48754_/X _48773_/Y _48774_/Y sky130_fd_sc_hd__o21ai_4
X_79594_ _79594_/A _79594_/B _79588_/Y _79594_/Y sky130_fd_sc_hd__nand3_4
X_45986_ _45985_/Y _86827_/D sky130_fd_sc_hd__inv_2
X_47725_ _47725_/A _54903_/B sky130_fd_sc_hd__inv_2
X_78545_ _82514_/Q _82770_/D _82482_/D sky130_fd_sc_hd__xor2_4
X_44937_ _74545_/C _44933_/X _44936_/X _44937_/Y sky130_fd_sc_hd__o21ai_4
X_63771_ _63749_/A _63772_/B sky130_fd_sc_hd__buf_2
X_75757_ _80917_/Q _75754_/Y _75756_/X _75757_/Y sky130_fd_sc_hd__o21ai_4
X_60983_ _64032_/A _63738_/B sky130_fd_sc_hd__buf_2
X_72969_ _72967_/X _72969_/B _72969_/C _72969_/Y sky130_fd_sc_hd__nand3_4
X_65510_ _65342_/X _83076_/Q _65391_/X _65509_/X _65510_/X sky130_fd_sc_hd__a211o_4
X_62722_ _62673_/A _62673_/B _75918_/B _62722_/Y sky130_fd_sc_hd__nor3_4
X_74708_ _74711_/A _74708_/Y sky130_fd_sc_hd__inv_2
X_47656_ _47650_/Y _47651_/X _47655_/X _86612_/D sky130_fd_sc_hd__a21oi_4
X_66490_ _66501_/A _66501_/B _66490_/C _66490_/X sky130_fd_sc_hd__and3_4
X_78476_ _78476_/A _78476_/Y sky130_fd_sc_hd__inv_2
X_44868_ _80670_/Q _45387_/A sky130_fd_sc_hd__inv_2
X_75688_ _75688_/A _80831_/Q _75688_/Y sky130_fd_sc_hd__xnor2_4
X_46607_ _52577_/B _51744_/B sky130_fd_sc_hd__buf_2
X_65441_ _65387_/A _65441_/B _65441_/X sky130_fd_sc_hd__and2_4
X_77427_ _77423_/Y _77426_/C _77422_/Y _77427_/Y sky130_fd_sc_hd__o21ai_4
X_43819_ _41108_/X _43817_/X _69555_/B _43818_/X _87252_/D sky130_fd_sc_hd__a2bb2o_4
X_62653_ _62653_/A _62653_/B _75923_/B _62653_/Y sky130_fd_sc_hd__nor3_4
X_74639_ _74638_/X _56589_/A _45479_/A _74633_/X _83004_/D sky130_fd_sc_hd__a2bb2o_4
X_47587_ _47595_/A _47595_/B _47595_/C _53133_/D _47587_/X sky130_fd_sc_hd__and4_4
X_44799_ _41432_/Y _44788_/X _86948_/Q _44789_/X _86948_/D sky130_fd_sc_hd__a2bb2o_4
X_49326_ _48193_/X _49326_/X sky130_fd_sc_hd__buf_2
X_61604_ _61476_/A _61634_/B sky130_fd_sc_hd__buf_2
X_68160_ _68160_/A _68160_/X sky130_fd_sc_hd__buf_2
X_46538_ _46525_/X _49140_/A _46537_/X _46539_/A sky130_fd_sc_hd__o21ai_4
X_65372_ _84204_/Q _65373_/C sky130_fd_sc_hd__inv_2
X_77358_ _77354_/X _77360_/C _77359_/A _77371_/A sky130_fd_sc_hd__a21boi_4
X_62584_ _62582_/Y _62540_/X _62583_/Y _62584_/Y sky130_fd_sc_hd__a21oi_4
X_67111_ _67087_/A _88125_/Q _67111_/X sky130_fd_sc_hd__and2_4
X_64323_ _64323_/A _64323_/X sky130_fd_sc_hd__buf_2
X_76309_ _76288_/Y _76309_/B _76309_/X sky130_fd_sc_hd__or2_4
X_61535_ _61476_/A _61546_/B sky130_fd_sc_hd__buf_2
X_49257_ _49261_/A _50777_/B _49257_/Y sky130_fd_sc_hd__nand2_4
X_68091_ _68088_/X _66559_/Y _68089_/X _68090_/Y _68091_/X sky130_fd_sc_hd__a211o_4
X_46469_ _48034_/B _46469_/B _46469_/Y sky130_fd_sc_hd__nand2_4
X_77289_ _77272_/Y _77270_/X _77288_/Y _77290_/B sky130_fd_sc_hd__a21oi_4
X_48208_ _48184_/A _48207_/X _48208_/Y sky130_fd_sc_hd__nand2_4
X_67042_ _87116_/Q _66988_/X _67040_/X _67041_/X _67042_/X sky130_fd_sc_hd__a211o_4
X_79028_ _82746_/Q _79028_/B _79028_/X sky130_fd_sc_hd__xor2_4
X_64254_ _79846_/B _63258_/X _64253_/X _64254_/X sky130_fd_sc_hd__a21o_4
X_49188_ _48934_/A _49405_/A sky130_fd_sc_hd__buf_2
X_61466_ _72528_/A _61468_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_444_0_CLK clkbuf_9_222_0_CLK/X _81224_/CLK sky130_fd_sc_hd__clkbuf_1
X_63205_ _63203_/X _64412_/C _63204_/X _63239_/D _63205_/X sky130_fd_sc_hd__and4_4
X_48139_ _48133_/Y _48109_/X _48138_/X _86564_/D sky130_fd_sc_hd__a21oi_4
X_60417_ _60417_/A _60515_/B sky130_fd_sc_hd__buf_2
X_64185_ _64181_/X _63741_/X _64182_/Y _64183_/Y _64184_/X _64185_/X
+ sky130_fd_sc_hd__a41o_4
X_61397_ _72515_/D _61398_/C sky130_fd_sc_hd__buf_2
X_51150_ _51160_/A _51160_/B _51141_/X _52841_/D _51150_/X sky130_fd_sc_hd__and4_4
X_63136_ _63342_/C _63147_/C sky130_fd_sc_hd__buf_2
X_60348_ _65680_/A _64939_/A sky130_fd_sc_hd__buf_2
X_68993_ _68993_/A _68993_/X sky130_fd_sc_hd__buf_2
X_50101_ _48979_/A _50082_/B _50059_/C _50101_/X sky130_fd_sc_hd__and3_4
X_51081_ _86077_/Q _51073_/X _51080_/Y _51081_/Y sky130_fd_sc_hd__o21ai_4
X_67944_ _86950_/Q _67942_/X _67872_/X _67943_/X _67944_/X sky130_fd_sc_hd__a211o_4
X_63067_ _63020_/A _63067_/X sky130_fd_sc_hd__buf_2
X_60279_ _60249_/X _60276_/Y _60299_/A _60277_/X _60278_/Y _60279_/Y
+ sky130_fd_sc_hd__a41oi_4
X_83990_ _84003_/CLK _83990_/D _82638_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_459_0_CLK clkbuf_9_229_0_CLK/X _86611_/CLK sky130_fd_sc_hd__clkbuf_1
X_50032_ _50028_/Y _50029_/X _50031_/X _86278_/D sky130_fd_sc_hd__a21oi_4
X_62018_ _62016_/Y _61959_/X _62017_/Y _62018_/Y sky130_fd_sc_hd__a21oi_4
X_82941_ _82369_/CLK _78096_/Y _82941_/Q sky130_fd_sc_hd__dfxtp_4
X_67875_ _68129_/A _67875_/X sky130_fd_sc_hd__buf_2
X_69614_ _69610_/X _69613_/X _69389_/X _69614_/Y sky130_fd_sc_hd__a21oi_4
X_54840_ _54758_/A _54850_/A sky130_fd_sc_hd__buf_2
X_66826_ _66499_/B _66815_/Y _66793_/X _66825_/Y _66826_/X sky130_fd_sc_hd__a211o_4
X_85660_ _85436_/CLK _53294_/Y _85660_/Q sky130_fd_sc_hd__dfxtp_4
X_82872_ _82675_/CLK _82496_/Q _82872_/Q sky130_fd_sc_hd__dfxtp_4
X_84611_ _84469_/CLK _60492_/Y _79151_/A sky130_fd_sc_hd__dfxtp_4
X_81823_ _81660_/CLK _81631_/Q _81823_/Q sky130_fd_sc_hd__dfxtp_4
X_69545_ _87509_/Q _69468_/X _59036_/A _69544_/X _69545_/X sky130_fd_sc_hd__a211o_4
X_54771_ _54769_/Y _54747_/X _54770_/X _54771_/Y sky130_fd_sc_hd__a21oi_4
X_66757_ _60371_/A _66757_/X sky130_fd_sc_hd__buf_2
X_85591_ _83068_/CLK _85591_/D _85591_/Q sky130_fd_sc_hd__dfxtp_4
X_51983_ _51982_/X _53504_/B _51983_/Y sky130_fd_sc_hd__nand2_4
X_63969_ _63741_/A _63969_/X sky130_fd_sc_hd__buf_2
X_56510_ _56510_/A _56520_/B _56510_/C _56510_/Y sky130_fd_sc_hd__nand3_4
X_87330_ _87333_/CLK _87330_/D _87330_/Q sky130_fd_sc_hd__dfxtp_4
X_53722_ _53846_/A _53722_/X sky130_fd_sc_hd__buf_2
X_65708_ _65825_/A _86511_/Q _65708_/X sky130_fd_sc_hd__and2_4
X_84542_ _84549_/CLK _84542_/D _76990_/A sky130_fd_sc_hd__dfxtp_4
X_50934_ _50941_/A _50941_/B _50948_/C _46707_/X _50934_/X sky130_fd_sc_hd__and4_4
X_57490_ _84993_/Q _47806_/X _57489_/Y _57490_/Y sky130_fd_sc_hd__o21ai_4
X_81754_ _81783_/CLK _76100_/B _81754_/Q sky130_fd_sc_hd__dfxtp_4
X_69476_ _69423_/X _69340_/X _69474_/Y _69475_/Y _69476_/X sky130_fd_sc_hd__a211o_4
X_66688_ _69245_/A _66688_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_503_0_CLK clkbuf_9_502_0_CLK/A clkbuf_9_503_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_56441_ _56139_/X _56439_/X _56440_/Y _56441_/Y sky130_fd_sc_hd__o21ai_4
X_80705_ _80681_/CLK _80737_/Q _75558_/A sky130_fd_sc_hd__dfxtp_4
X_68427_ _68405_/A _68427_/B _68427_/X sky130_fd_sc_hd__and2_4
X_87261_ _88034_/CLK _43800_/X _69443_/B sky130_fd_sc_hd__dfxtp_4
X_53653_ _53747_/A _53653_/X sky130_fd_sc_hd__buf_2
X_65639_ _65877_/A _65704_/A sky130_fd_sc_hd__buf_2
X_84473_ _82452_/CLK _61537_/Y _79141_/B sky130_fd_sc_hd__dfxtp_4
X_50865_ _50863_/Y _50849_/X _50864_/Y _86118_/D sky130_fd_sc_hd__a21boi_4
X_81685_ _81684_/CLK _81685_/D _81685_/Q sky130_fd_sc_hd__dfxtp_4
X_86212_ _86490_/CLK _50382_/Y _86212_/Q sky130_fd_sc_hd__dfxtp_4
X_52604_ _85788_/Q _52601_/X _52603_/Y _52604_/Y sky130_fd_sc_hd__o21ai_4
X_59160_ _58641_/A _59160_/X sky130_fd_sc_hd__buf_2
X_83424_ _83756_/CLK _71653_/Y _83424_/Q sky130_fd_sc_hd__dfxtp_4
X_56372_ _56439_/A _56372_/X sky130_fd_sc_hd__buf_2
X_80636_ _80636_/A _80635_/Y _80636_/Y sky130_fd_sc_hd__xnor2_4
X_68358_ _68823_/A _68358_/X sky130_fd_sc_hd__buf_2
X_87192_ _87189_/CLK _87192_/D _67975_/B sky130_fd_sc_hd__dfxtp_4
X_53584_ _53582_/Y _53537_/X _53583_/X _85608_/D sky130_fd_sc_hd__a21oi_4
X_50796_ _86131_/Q _50775_/X _50795_/Y _50796_/Y sky130_fd_sc_hd__o21ai_4
XPHY_104 sky130_fd_sc_hd__decap_3
X_58111_ _57983_/X _85380_/Q _58110_/X _58111_/Y sky130_fd_sc_hd__o21ai_4
XPHY_115 sky130_fd_sc_hd__decap_3
X_55323_ _55323_/A _85134_/Q _55323_/X sky130_fd_sc_hd__and2_4
X_67309_ _87348_/Q _67239_/X _67240_/X _67308_/X _67309_/X sky130_fd_sc_hd__a211o_4
X_86143_ _85536_/CLK _86143_/D _86143_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_126 sky130_fd_sc_hd__decap_3
X_52535_ _52501_/X _54054_/B _52535_/Y sky130_fd_sc_hd__nand2_4
X_59091_ _58864_/X _59089_/Y _59090_/Y _58943_/X _58868_/X _59091_/X
+ sky130_fd_sc_hd__o32a_4
X_83355_ _83761_/CLK _83355_/D _83355_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_137 sky130_fd_sc_hd__decap_3
X_80567_ _84772_/Q _84164_/Q _80567_/X sky130_fd_sc_hd__xor2_4
X_68289_ _68272_/X _67769_/Y _68287_/X _68288_/Y _68289_/X sky130_fd_sc_hd__a211o_4
XPHY_148 sky130_fd_sc_hd__decap_3
XPHY_159 sky130_fd_sc_hd__decap_3
X_58042_ _58017_/X _85386_/Q _58041_/X _58042_/Y sky130_fd_sc_hd__o21ai_4
X_70320_ _70337_/A _70320_/X sky130_fd_sc_hd__buf_2
X_82306_ _80835_/CLK _77002_/X _40546_/A sky130_fd_sc_hd__dfxtp_4
X_55254_ _55254_/A _83320_/Q _55253_/X _55290_/A sky130_fd_sc_hd__nand3_4
X_86074_ _85754_/CLK _86074_/D _86074_/Q sky130_fd_sc_hd__dfxtp_4
X_40480_ _40479_/X _40480_/X sky130_fd_sc_hd__buf_2
X_52466_ _52466_/A _53985_/B _52466_/Y sky130_fd_sc_hd__nand2_4
X_83286_ _85542_/CLK _83286_/D _83286_/Q sky130_fd_sc_hd__dfxtp_4
X_80498_ _80496_/X _80498_/B _80498_/Y sky130_fd_sc_hd__xnor2_4
Xclkbuf_8_71_0_CLK clkbuf_8_71_0_CLK/A clkbuf_8_71_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_54205_ _54215_/A _47420_/Y _54205_/Y sky130_fd_sc_hd__nand2_4
X_85025_ _85089_/CLK _85025_/D _45393_/A sky130_fd_sc_hd__dfxtp_4
X_51417_ _51414_/Y _51229_/X _51416_/X _86014_/D sky130_fd_sc_hd__a21oi_4
X_70251_ _70260_/A _70260_/B _70251_/C _70260_/D _70251_/X sky130_fd_sc_hd__and4_4
X_82237_ _82515_/CLK _82269_/Q _82237_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_3_0_CLK clkbuf_7_3_0_CLK/A clkbuf_8_7_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_55185_ _85037_/Q _55145_/A _55168_/X _55184_/X _55185_/X sky130_fd_sc_hd__a211o_4
X_52397_ _52324_/A _52397_/X sky130_fd_sc_hd__buf_2
X_42150_ _42162_/A _42150_/X sky130_fd_sc_hd__buf_2
X_54136_ _54217_/A _54160_/B sky130_fd_sc_hd__buf_2
X_51348_ _52528_/A _51352_/B _51352_/C _51348_/X sky130_fd_sc_hd__and3_4
X_70182_ _70180_/Y _70157_/X _70181_/Y _70182_/Y sky130_fd_sc_hd__o21ai_4
X_82168_ _84166_/CLK _84160_/Q _82168_/Q sky130_fd_sc_hd__dfxtp_4
X_59993_ _59951_/D _60129_/B _59974_/Y _59981_/Y _59992_/Y _84677_/D
+ sky130_fd_sc_hd__a41oi_4
X_41101_ _40932_/A _41102_/B sky130_fd_sc_hd__buf_2
X_81119_ _80697_/CLK _79868_/X _75688_/A sky130_fd_sc_hd__dfxtp_4
X_42081_ _42081_/A _43161_/A sky130_fd_sc_hd__buf_2
X_58944_ _58864_/X _58941_/Y _58942_/Y _58943_/X _58868_/X _58944_/X
+ sky130_fd_sc_hd__o32a_4
X_54067_ _54067_/A _54067_/X sky130_fd_sc_hd__buf_2
X_51279_ _51277_/Y _51263_/X _51278_/X _51279_/Y sky130_fd_sc_hd__a21oi_4
X_74990_ _74990_/A _74987_/C _74990_/X sky130_fd_sc_hd__and2_4
X_86976_ _87333_/CLK _86976_/D _86976_/Q sky130_fd_sc_hd__dfxtp_4
X_82099_ _82349_/CLK _77471_/B _82099_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_86_0_CLK clkbuf_8_87_0_CLK/A clkbuf_8_86_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_53018_ _85712_/Q _53010_/X _53017_/Y _53018_/Y sky130_fd_sc_hd__o21ai_4
X_41032_ _41032_/A _41032_/X sky130_fd_sc_hd__buf_2
X_73941_ _41941_/Y _56182_/X _73819_/X _73940_/Y _73941_/X sky130_fd_sc_hd__a211o_4
X_85927_ _85447_/CLK _85927_/D _85927_/Q sky130_fd_sc_hd__dfxtp_4
X_58875_ _58828_/X _58872_/Y _58873_/Y _58874_/X _58832_/X _58875_/X
+ sky130_fd_sc_hd__o32a_4
X_45840_ _85028_/Q _45824_/B _45840_/Y sky130_fd_sc_hd__nor2_4
X_57826_ _57811_/X _85403_/Q _57825_/X _57826_/Y sky130_fd_sc_hd__o21ai_4
X_76660_ _76662_/A _76658_/Y _76662_/C _76661_/A sky130_fd_sc_hd__a21oi_4
X_73872_ _73438_/B _73872_/X sky130_fd_sc_hd__buf_2
X_85858_ _83562_/CLK _52258_/Y _65890_/B sky130_fd_sc_hd__dfxtp_4
X_75611_ _80998_/Q _75611_/B _80966_/D sky130_fd_sc_hd__xor2_4
X_72823_ _72821_/X _72822_/Y _72766_/X _72823_/Y sky130_fd_sc_hd__a21oi_4
X_84809_ _85957_/CLK _84809_/D _84809_/Q sky130_fd_sc_hd__dfxtp_4
X_57757_ _57757_/A _58857_/A sky130_fd_sc_hd__buf_2
X_45771_ _85001_/Q _45705_/X _45691_/X _45771_/X sky130_fd_sc_hd__o21a_4
X_76591_ _76583_/Y _76616_/B _76591_/X sky130_fd_sc_hd__xor2_4
X_54969_ _54985_/A _47543_/Y _54969_/Y sky130_fd_sc_hd__nand2_4
X_42983_ _40469_/X _42962_/X _66948_/B _42963_/X _87619_/D sky130_fd_sc_hd__a2bb2o_4
X_85789_ _84807_/CLK _52600_/Y _85789_/Q sky130_fd_sc_hd__dfxtp_4
X_47510_ _47556_/A _47549_/B sky130_fd_sc_hd__buf_2
X_78330_ _78330_/A _78330_/B _78332_/A sky130_fd_sc_hd__nand2_4
X_56708_ _56708_/A _56707_/X _56708_/C _57284_/A sky130_fd_sc_hd__nand3_4
X_44722_ _44721_/Y _44722_/Y sky130_fd_sc_hd__inv_2
X_75542_ _80704_/Q _75554_/B _75543_/B sky130_fd_sc_hd__xor2_4
X_87528_ _87782_/CLK _87528_/D _87528_/Q sky130_fd_sc_hd__dfxtp_4
X_41934_ _41934_/A _41934_/Y sky130_fd_sc_hd__inv_2
X_48490_ _48483_/Y _48459_/X _48489_/X _86518_/D sky130_fd_sc_hd__a21oi_4
X_72754_ _72749_/X _72753_/X _72735_/X _72754_/X sky130_fd_sc_hd__a21o_4
X_57688_ _59629_/A _57689_/A sky130_fd_sc_hd__buf_2
X_47441_ _47434_/Y _47414_/X _47440_/X _86635_/D sky130_fd_sc_hd__a21oi_4
X_71705_ _58298_/Y _71695_/X _71704_/Y _83404_/D sky130_fd_sc_hd__o21ai_4
X_59427_ _59427_/A _59427_/Y sky130_fd_sc_hd__inv_2
X_78261_ _82683_/Q _78261_/B _78261_/X sky130_fd_sc_hd__xor2_4
X_44653_ _41069_/Y _44648_/X _87015_/Q _44650_/X _44653_/X sky130_fd_sc_hd__a2bb2o_4
X_56639_ _56638_/X _56639_/X sky130_fd_sc_hd__buf_2
X_75473_ _75473_/A _75477_/A sky130_fd_sc_hd__inv_2
X_87459_ _87149_/CLK _43362_/X _87459_/Q sky130_fd_sc_hd__dfxtp_4
X_41865_ _41902_/A _41877_/A sky130_fd_sc_hd__inv_2
X_72685_ _73078_/A _72686_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_24_0_CLK clkbuf_8_25_0_CLK/A clkbuf_9_49_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_77212_ _77207_/B _77210_/X _77211_/Y _77212_/Y sky130_fd_sc_hd__a21boi_4
X_43604_ _55102_/A _43604_/X sky130_fd_sc_hd__buf_2
X_74424_ _83069_/Q _74412_/X _74423_/Y _74424_/Y sky130_fd_sc_hd__o21ai_4
X_40816_ _40816_/A _40816_/Y sky130_fd_sc_hd__inv_2
X_59358_ _59208_/X _86052_/Q _59357_/X _59358_/Y sky130_fd_sc_hd__o21ai_4
X_47372_ _47372_/A _47372_/Y sky130_fd_sc_hd__inv_2
X_71636_ _59484_/Y _71628_/X _71635_/Y _71636_/Y sky130_fd_sc_hd__o21ai_4
X_78192_ _78192_/A _78191_/X _78192_/Y sky130_fd_sc_hd__nand2_4
X_44584_ _44554_/X _44555_/X _40903_/X _44583_/Y _44557_/X _87045_/D
+ sky130_fd_sc_hd__o32ai_4
XPHY_6 sky130_fd_sc_hd__decap_3
X_41796_ _40628_/X _82337_/Q _41795_/X _41796_/Y sky130_fd_sc_hd__o21ai_4
X_49111_ _40380_/X _81771_/Q _49110_/Y _49112_/A sky130_fd_sc_hd__o21ai_4
X_46323_ _46316_/Y _46300_/X _46322_/X _46323_/Y sky130_fd_sc_hd__a21oi_4
X_58309_ _58271_/X _83402_/Q _58308_/Y _84882_/D sky130_fd_sc_hd__o21a_4
X_77143_ _77141_/B _77143_/B _81916_/Q _77143_/Y sky130_fd_sc_hd__nand3_4
X_43535_ _40404_/X _43532_/X _87372_/Q _43533_/X _43535_/X sky130_fd_sc_hd__a2bb2o_4
X_74355_ _45954_/X _58334_/A _56158_/A _74355_/Y sky130_fd_sc_hd__nand3_4
X_40747_ _40817_/A _82852_/Q _40747_/X sky130_fd_sc_hd__or2_4
X_59289_ _59285_/Y _59288_/Y _59278_/X _59289_/X sky130_fd_sc_hd__a21o_4
X_71567_ _71585_/A _71583_/B sky130_fd_sc_hd__buf_2
X_49042_ _49022_/A _53858_/B _49042_/X sky130_fd_sc_hd__and2_4
X_61320_ _61317_/X _72575_/A _61260_/X _61319_/X _61277_/B _61320_/Y
+ sky130_fd_sc_hd__a41oi_4
X_73306_ _73306_/A _73426_/A sky130_fd_sc_hd__buf_2
X_46254_ _83656_/Q _53946_/B sky130_fd_sc_hd__inv_2
XPHY_660 sky130_fd_sc_hd__decap_3
X_70518_ _70511_/A _70949_/B _70508_/X _70518_/Y sky130_fd_sc_hd__nand3_4
X_77074_ _82092_/Q _77074_/B _82341_/D sky130_fd_sc_hd__xor2_4
X_43466_ _43182_/Y _43466_/X sky130_fd_sc_hd__buf_2
X_74286_ _72714_/A _72714_/B _74286_/C _74286_/Y sky130_fd_sc_hd__nand3_4
XPHY_671 sky130_fd_sc_hd__decap_3
Xclkbuf_8_39_0_CLK clkbuf_8_39_0_CLK/A clkbuf_9_79_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_40678_ _40678_/A _40678_/X sky130_fd_sc_hd__buf_2
X_71498_ _71308_/A _71815_/B _71496_/C _71498_/X sky130_fd_sc_hd__and3_4
XPHY_682 sky130_fd_sc_hd__decap_3
XPHY_693 sky130_fd_sc_hd__decap_3
X_45205_ _45192_/X _45201_/Y _45204_/Y _45205_/Y sky130_fd_sc_hd__a21oi_4
X_76025_ _76025_/A _81744_/D _76025_/X sky130_fd_sc_hd__xor2_4
X_42417_ _42417_/A _42417_/X sky130_fd_sc_hd__buf_2
X_61251_ _61131_/Y _61151_/Y _64454_/B _61249_/Y _61250_/Y _84498_/D
+ sky130_fd_sc_hd__a41oi_4
X_73237_ _73234_/X _73236_/X _73067_/X _73237_/X sky130_fd_sc_hd__a21o_4
X_70449_ _50302_/B _70421_/Y _70448_/Y _83771_/D sky130_fd_sc_hd__o21ai_4
X_46185_ _46183_/X _46150_/B _46184_/Y _46185_/X sky130_fd_sc_hd__and3_4
X_43397_ _43397_/A _43397_/X sky130_fd_sc_hd__buf_2
X_60202_ _60202_/A _60324_/C sky130_fd_sc_hd__buf_2
X_45136_ _85202_/Q _45102_/X _45135_/X _45136_/Y sky130_fd_sc_hd__o21ai_4
X_42348_ _42330_/X _42346_/X _41705_/X _87909_/Q _42347_/X _42348_/Y
+ sky130_fd_sc_hd__o32ai_4
X_61182_ _64250_/A _61182_/X sky130_fd_sc_hd__buf_2
X_73168_ _73168_/A _73167_/X _73169_/B sky130_fd_sc_hd__nand2_4
X_60133_ _60091_/C _59922_/C _60091_/A _60133_/Y sky130_fd_sc_hd__o21ai_4
X_72119_ _59325_/X _72116_/Y _72118_/Y _59342_/X _59329_/X _72119_/X
+ sky130_fd_sc_hd__o32a_4
X_49944_ _49941_/Y _49924_/X _49943_/X _86295_/D sky130_fd_sc_hd__a21oi_4
X_45067_ _45067_/A _45067_/B _45067_/Y sky130_fd_sc_hd__nand2_4
X_65990_ _65484_/A _65990_/X sky130_fd_sc_hd__buf_2
X_42279_ _42204_/X _42279_/X sky130_fd_sc_hd__buf_2
X_73099_ _53678_/B _73098_/Y _73099_/X sky130_fd_sc_hd__xor2_4
X_77976_ _78043_/A _77975_/A _77977_/A sky130_fd_sc_hd__nand2_4
X_44018_ _44146_/A _44019_/A sky130_fd_sc_hd__inv_2
X_79715_ _79711_/X _79714_/Y _79715_/X sky130_fd_sc_hd__xor2_4
X_64941_ _84221_/Q _64942_/C sky130_fd_sc_hd__inv_2
X_76927_ _76924_/A _81599_/Q _76927_/Y sky130_fd_sc_hd__nand2_4
X_60064_ _60064_/A _60081_/B _60064_/C _60064_/Y sky130_fd_sc_hd__nor3_4
X_49875_ _58130_/B _49853_/X _49874_/Y _49875_/Y sky130_fd_sc_hd__o21ai_4
X_48826_ _86475_/Q _48809_/X _48825_/Y _48826_/Y sky130_fd_sc_hd__o21ai_4
X_67660_ _87154_/Q _67585_/X _67633_/X _67659_/X _67660_/X sky130_fd_sc_hd__a211o_4
X_79646_ _79636_/X _79646_/B _79646_/Y sky130_fd_sc_hd__nand2_4
X_64872_ _64778_/A _85815_/Q _64872_/X sky130_fd_sc_hd__and2_4
X_76858_ _76858_/A _76857_/Y _76862_/A sky130_fd_sc_hd__xor2_4
X_66611_ _66607_/X _66610_/X _66411_/A _66611_/Y sky130_fd_sc_hd__a21oi_4
X_63823_ _63819_/Y _63823_/B _63821_/Y _63822_/Y _63823_/X sky130_fd_sc_hd__and4_4
X_75809_ _75810_/A _75810_/C _75810_/B _75811_/A sky130_fd_sc_hd__a21o_4
X_48757_ _48777_/A _50440_/B _48757_/Y sky130_fd_sc_hd__nand2_4
X_67591_ _67354_/X _67591_/X sky130_fd_sc_hd__buf_2
X_79577_ _79577_/A _79564_/Y _79578_/B sky130_fd_sc_hd__nand2_4
X_45969_ _40386_/Y _45963_/X _66644_/B _45964_/X _86835_/D sky130_fd_sc_hd__a2bb2o_4
X_76789_ _76786_/X _76788_/Y _76790_/B sky130_fd_sc_hd__xnor2_4
X_69330_ _69234_/A _87781_/Q _69330_/X sky130_fd_sc_hd__and2_4
X_47708_ _47661_/A _47749_/C sky130_fd_sc_hd__buf_2
X_66542_ _67816_/A _68614_/A sky130_fd_sc_hd__buf_2
X_78528_ _78528_/A _78528_/B _78528_/X sky130_fd_sc_hd__and2_4
X_63754_ _63724_/A _63757_/C sky130_fd_sc_hd__buf_2
X_48688_ _48652_/X _48136_/A _48687_/Y _74505_/A sky130_fd_sc_hd__o21ai_4
X_60966_ _60966_/A _60967_/A sky130_fd_sc_hd__inv_2
X_62705_ _62701_/Y _62660_/X _62702_/Y _62703_/Y _62704_/X _62705_/X
+ sky130_fd_sc_hd__a41o_4
X_69261_ _69442_/A _69261_/X sky130_fd_sc_hd__buf_2
X_47639_ _83629_/Q _47639_/Y sky130_fd_sc_hd__inv_2
X_66473_ _66501_/A _66419_/X _84116_/Q _66473_/X sky130_fd_sc_hd__and3_4
X_78459_ _78458_/A _82669_/D _78460_/A sky130_fd_sc_hd__nand2_4
X_63685_ _63697_/A _58201_/A _63537_/C _63685_/X sky130_fd_sc_hd__and3_4
X_60897_ _60891_/Y _60543_/B _60896_/Y _60897_/Y sky130_fd_sc_hd__nand3_4
X_68212_ _84011_/Q _68200_/X _68211_/X _68212_/X sky130_fd_sc_hd__a21bo_4
X_65424_ _65350_/X _86209_/Q _65400_/X _65423_/X _65424_/X sky130_fd_sc_hd__a211o_4
X_50650_ _86160_/Q _50563_/X _50649_/Y _50650_/Y sky130_fd_sc_hd__o21ai_4
X_62636_ _62653_/A _62653_/B _62636_/C _62636_/Y sky130_fd_sc_hd__nor3_4
X_81470_ _81482_/CLK _81470_/D _81470_/Q sky130_fd_sc_hd__dfxtp_4
X_69192_ _88047_/Q _68975_/X _68976_/X _69191_/X _69192_/X sky130_fd_sc_hd__a211o_4
X_49309_ _49307_/Y _49281_/X _49308_/X _86413_/D sky130_fd_sc_hd__a21oi_4
X_80421_ _59229_/A _84150_/Q _80423_/A sky130_fd_sc_hd__xor2_4
X_68143_ _84028_/Q _68140_/X _68142_/X _84028_/D sky130_fd_sc_hd__a21bo_4
X_65355_ _65272_/X _85540_/Q _65326_/X _65354_/X _65355_/X sky130_fd_sc_hd__a211o_4
X_50581_ _50576_/Y _50577_/X _50580_/Y _50581_/Y sky130_fd_sc_hd__a21boi_4
X_62567_ _62533_/A _63655_/B _62532_/X _62569_/C sky130_fd_sc_hd__nand3_4
Xclkbuf_10_383_0_CLK clkbuf_9_191_0_CLK/X _85761_/CLK sky130_fd_sc_hd__clkbuf_1
X_52320_ _52320_/A _48998_/A _52320_/X sky130_fd_sc_hd__and2_4
X_64306_ _64306_/A _64307_/B sky130_fd_sc_hd__buf_2
X_83140_ _83141_/CLK _83140_/D _83140_/Q sky130_fd_sc_hd__dfxtp_4
X_61518_ _61518_/A _61518_/B _79142_/B _61518_/Y sky130_fd_sc_hd__nor3_4
X_80352_ _80352_/A _80341_/Y _80353_/B sky130_fd_sc_hd__nand2_4
X_68074_ _68644_/A _68444_/A sky130_fd_sc_hd__buf_2
X_65286_ _65211_/X _85543_/Q _65212_/X _65285_/X _65286_/X sky130_fd_sc_hd__a211o_4
X_62498_ _62483_/X _62541_/B _62498_/C _62498_/Y sky130_fd_sc_hd__nor3_4
X_67025_ _57776_/A _67025_/X sky130_fd_sc_hd__buf_2
X_52251_ _85859_/Q _52239_/X _52250_/Y _52251_/Y sky130_fd_sc_hd__o21ai_4
X_83071_ _85884_/CLK _83071_/D _83071_/Q sky130_fd_sc_hd__dfxtp_4
X_64237_ _64250_/A _84855_/Q _64250_/C _64237_/Y sky130_fd_sc_hd__nand3_4
X_61449_ _61429_/A _61448_/X _61429_/C _61449_/Y sky130_fd_sc_hd__nand3_4
X_80283_ _80281_/Y _80282_/Y _80283_/Y sky130_fd_sc_hd__nor2_4
X_51202_ _51149_/A _51203_/B sky130_fd_sc_hd__buf_2
X_82022_ _81990_/CLK _77768_/B _82022_/Q sky130_fd_sc_hd__dfxtp_4
X_52182_ _52182_/A _52194_/B _52182_/C _52182_/X sky130_fd_sc_hd__and3_4
X_64168_ _61673_/B _64179_/B _64179_/C _64179_/D _64168_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_10_398_0_CLK clkbuf_9_199_0_CLK/X _82822_/CLK sky130_fd_sc_hd__clkbuf_1
X_51133_ _51131_/Y _51119_/X _51132_/X _86068_/D sky130_fd_sc_hd__a21oi_4
X_63119_ _58543_/Y _63073_/X _63117_/X _58320_/A _63118_/X _63119_/Y
+ sky130_fd_sc_hd__o32ai_4
X_86830_ _87990_/CLK _45978_/X _86830_/Q sky130_fd_sc_hd__dfxtp_4
X_56990_ _56943_/X _56988_/Y _56989_/Y _85104_/D sky130_fd_sc_hd__o21ai_4
X_68976_ _66180_/A _68976_/X sky130_fd_sc_hd__buf_2
X_64099_ _64094_/X _64048_/X _64095_/Y _64096_/Y _64098_/X _64099_/X
+ sky130_fd_sc_hd__a41o_4
X_51064_ _86080_/Q _51047_/X _51063_/Y _51064_/Y sky130_fd_sc_hd__o21ai_4
X_55941_ _56390_/C _55641_/A _55610_/X _55940_/X _55941_/X sky130_fd_sc_hd__a211o_4
X_67927_ _67972_/A _67927_/B _67927_/X sky130_fd_sc_hd__and2_4
X_86761_ _84287_/CLK _46205_/Y _57701_/A sky130_fd_sc_hd__dfxtp_4
X_83973_ _83973_/CLK _83973_/D _83973_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_321_0_CLK clkbuf_9_160_0_CLK/X _85727_/CLK sky130_fd_sc_hd__clkbuf_1
X_50015_ _86281_/Q _50012_/X _50014_/Y _50015_/Y sky130_fd_sc_hd__o21ai_4
X_85712_ _85712_/CLK _53020_/Y _85712_/Q sky130_fd_sc_hd__dfxtp_4
X_58660_ _58660_/A _58649_/B _58660_/Y sky130_fd_sc_hd__nor2_4
X_82924_ _82924_/CLK _78202_/X _82924_/Q sky130_fd_sc_hd__dfxtp_4
X_55872_ _55872_/A _55871_/X _55873_/A sky130_fd_sc_hd__and2_4
X_67858_ _68442_/A _67858_/X sky130_fd_sc_hd__buf_2
X_86692_ _86372_/CLK _46897_/Y _58942_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_951_0_CLK clkbuf_9_475_0_CLK/X _86535_/CLK sky130_fd_sc_hd__clkbuf_1
X_57611_ _57630_/A _48081_/Y _57611_/Y sky130_fd_sc_hd__nand2_4
X_54823_ _54823_/A _47582_/A _54823_/Y sky130_fd_sc_hd__nand2_4
X_66809_ _87881_/Q _66759_/X _66807_/X _66808_/X _66809_/X sky130_fd_sc_hd__a211o_4
X_85643_ _85643_/CLK _85643_/D _85643_/Q sky130_fd_sc_hd__dfxtp_4
X_58591_ _58703_/A _58591_/X sky130_fd_sc_hd__buf_2
X_82855_ _82855_/CLK _78108_/B _82855_/Q sky130_fd_sc_hd__dfxtp_4
X_67789_ _67312_/X _67789_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_442_0_CLK clkbuf_9_443_0_CLK/A clkbuf_9_442_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_57542_ _84982_/Q _57527_/X _57541_/Y _57542_/Y sky130_fd_sc_hd__o21ai_4
X_81806_ _81296_/CLK _81614_/Q _81806_/Q sky130_fd_sc_hd__dfxtp_4
X_69528_ _69525_/X _69527_/X _69389_/X _69528_/Y sky130_fd_sc_hd__a21oi_4
X_88362_ _87859_/CLK _40643_/Y _68595_/B sky130_fd_sc_hd__dfxtp_4
X_54754_ _54672_/X _54775_/C sky130_fd_sc_hd__buf_2
X_85574_ _83564_/CLK _53760_/Y _85574_/Q sky130_fd_sc_hd__dfxtp_4
X_51966_ _51961_/X _50264_/B _51966_/Y sky130_fd_sc_hd__nand2_4
X_82786_ _82786_/CLK _82818_/Q _82786_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_336_0_CLK clkbuf_9_168_0_CLK/X _86054_/CLK sky130_fd_sc_hd__clkbuf_1
X_87313_ _86534_/CLK _43680_/X _72800_/A sky130_fd_sc_hd__dfxtp_4
X_53705_ _53611_/X _48550_/Y _53705_/Y sky130_fd_sc_hd__nand2_4
X_84525_ _84292_/CLK _61058_/X _61057_/C sky130_fd_sc_hd__dfxtp_4
X_50917_ _86107_/Q _50910_/X _50916_/Y _50917_/Y sky130_fd_sc_hd__o21ai_4
X_57473_ _58273_/A _57473_/B _57473_/Y sky130_fd_sc_hd__nand2_4
X_81737_ _86807_/CLK _81737_/D _41414_/A sky130_fd_sc_hd__dfxtp_4
X_69459_ _69322_/A _88284_/Q _69459_/X sky130_fd_sc_hd__and2_4
X_88293_ _87253_/CLK _41018_/Y _88293_/Q sky130_fd_sc_hd__dfxtp_4
X_54685_ _54674_/A _54707_/B _54674_/C _54685_/D _54685_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_966_0_CLK clkbuf_9_483_0_CLK/X _83304_/CLK sky130_fd_sc_hd__clkbuf_1
X_51897_ _51843_/A _51898_/B sky130_fd_sc_hd__buf_2
X_59212_ _59154_/A _86352_/Q _59212_/Y sky130_fd_sc_hd__nor2_4
X_56424_ _56431_/A _56433_/B _56424_/C _56424_/Y sky130_fd_sc_hd__nand3_4
X_87244_ _88012_/CLK _43834_/X _68546_/B sky130_fd_sc_hd__dfxtp_4
X_41650_ _41588_/X _41304_/A _41649_/X _41651_/A sky130_fd_sc_hd__o21ai_4
X_53636_ _53636_/A _53658_/B _53667_/C _53636_/X sky130_fd_sc_hd__and3_4
X_72470_ _72467_/Y _72469_/Y _57718_/A _72470_/X sky130_fd_sc_hd__a21o_4
X_84456_ _84564_/CLK _61753_/Y _78079_/B sky130_fd_sc_hd__dfxtp_4
X_50848_ _86121_/Q _50804_/X _50847_/Y _50848_/Y sky130_fd_sc_hd__o21ai_4
X_81668_ _81668_/CLK _79932_/Y _81668_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_457_0_CLK clkbuf_8_228_0_CLK/X clkbuf_9_457_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_40601_ _49140_/B _40601_/X sky130_fd_sc_hd__buf_2
X_59143_ _59143_/A _59143_/Y sky130_fd_sc_hd__inv_2
X_71421_ _71418_/B _71432_/B sky130_fd_sc_hd__buf_2
X_83407_ _83380_/CLK _83407_/D _83407_/Q sky130_fd_sc_hd__dfxtp_4
X_56355_ _56144_/X _56350_/X _56354_/Y _56355_/Y sky130_fd_sc_hd__o21ai_4
X_80619_ _80607_/A _80607_/B _80618_/X _80619_/X sky130_fd_sc_hd__a21o_4
X_41581_ _41486_/A _41581_/X sky130_fd_sc_hd__buf_2
X_87175_ _87178_/CLK _44278_/Y _43986_/A sky130_fd_sc_hd__dfxtp_4
X_53567_ _53622_/A _53567_/B _53567_/Y sky130_fd_sc_hd__nand2_4
X_84387_ _84503_/CLK _84387_/D _84387_/Q sky130_fd_sc_hd__dfxtp_4
X_50779_ _50764_/A _53993_/B _50779_/Y sky130_fd_sc_hd__nand2_4
X_81599_ _81473_/CLK _65466_/C _81599_/Q sky130_fd_sc_hd__dfxtp_4
X_43320_ _43316_/X _43319_/X _41245_/X _87483_/Q _43308_/X _43320_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55306_ _55177_/A _55306_/X sky130_fd_sc_hd__buf_2
X_74140_ _74140_/A _74202_/A sky130_fd_sc_hd__buf_2
X_86126_ _86030_/CLK _86126_/D _86126_/Q sky130_fd_sc_hd__dfxtp_4
X_52518_ _52518_/A _46464_/Y _52518_/Y sky130_fd_sc_hd__nand2_4
X_40532_ _40531_/X _40532_/X sky130_fd_sc_hd__buf_2
X_71352_ _70959_/C _71429_/A sky130_fd_sc_hd__buf_2
X_59074_ _59073_/X _85755_/Q _59037_/X _59074_/X sky130_fd_sc_hd__o21a_4
X_83338_ _83338_/CLK _83338_/D _83338_/Q sky130_fd_sc_hd__dfxtp_4
X_56286_ _56347_/A _56368_/A sky130_fd_sc_hd__buf_2
X_53498_ _53696_/A _53498_/X sky130_fd_sc_hd__buf_2
X_70303_ _70337_/A _70303_/X sky130_fd_sc_hd__buf_2
X_58025_ _57896_/A _58025_/X sky130_fd_sc_hd__buf_2
X_43251_ _43241_/X _43244_/X _41054_/X _87518_/Q _43250_/X _43251_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55237_ _55655_/A _55655_/B _83316_/Q _55237_/Y sky130_fd_sc_hd__a21oi_4
X_74071_ _74071_/A _73152_/X _74071_/Y sky130_fd_sc_hd__nor2_4
X_86057_ _85738_/CLK _51193_/Y _86057_/Q sky130_fd_sc_hd__dfxtp_4
X_40463_ _40931_/A _40463_/X sky130_fd_sc_hd__buf_2
X_52449_ _64743_/B _52422_/X _52448_/Y _52449_/Y sky130_fd_sc_hd__o21ai_4
X_71283_ _71183_/A _71268_/A _71279_/C _71276_/D _71283_/Y sky130_fd_sc_hd__nand4_4
X_83269_ _85332_/CLK _83269_/D _83269_/Q sky130_fd_sc_hd__dfxtp_4
X_42202_ _42173_/X _42200_/X _41316_/X _87981_/Q _42201_/X _42203_/A
+ sky130_fd_sc_hd__o32ai_4
X_73022_ _73020_/X _73021_/Y _72970_/X _73022_/Y sky130_fd_sc_hd__a21oi_4
X_85008_ _85040_/CLK _85008_/D _57414_/A sky130_fd_sc_hd__dfxtp_4
X_70234_ _70239_/A _70239_/B _83188_/Q _70239_/D _70234_/X sky130_fd_sc_hd__and4_4
X_43182_ _46450_/A _51340_/A _43182_/B1 _43182_/Y sky130_fd_sc_hd__a21oi_4
X_55168_ _55168_/A _55168_/X sky130_fd_sc_hd__buf_2
X_40394_ _41061_/A _82332_/Q _40393_/X _40394_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_10_904_0_CLK clkbuf_9_452_0_CLK/X _87859_/CLK sky130_fd_sc_hd__clkbuf_1
X_54119_ _54123_/A _54123_/B _54118_/X _52948_/D _54119_/X sky130_fd_sc_hd__and4_4
X_42133_ _41121_/X _42125_/X _88018_/Q _42126_/X _88018_/D sky130_fd_sc_hd__a2bb2o_4
X_77830_ _77835_/B _77830_/B _77831_/B sky130_fd_sc_hd__xnor2_4
X_70165_ _70165_/A _70160_/X _70162_/X _70164_/X _70165_/Y sky130_fd_sc_hd__nand4_4
X_47990_ _46317_/A _48044_/A sky130_fd_sc_hd__buf_2
X_55099_ _47838_/X _55118_/A sky130_fd_sc_hd__buf_2
X_59976_ _59976_/A _59977_/A sky130_fd_sc_hd__buf_2
Xclkbuf_5_21_0_CLK clkbuf_4_10_1_CLK/X clkbuf_6_43_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_46941_ _46941_/A _46944_/B sky130_fd_sc_hd__buf_2
X_42064_ _42060_/X _42049_/X _40929_/X _42063_/Y _41872_/X _42064_/Y
+ sky130_fd_sc_hd__o32ai_4
X_58927_ _58925_/X _85445_/Q _58926_/X _58927_/Y sky130_fd_sc_hd__o21ai_4
X_77761_ _82149_/Q _77761_/B _77761_/X sky130_fd_sc_hd__xor2_4
X_74973_ _80763_/Q _74965_/B _74973_/Y sky130_fd_sc_hd__nor2_4
X_70096_ _69974_/Y _59834_/A _70081_/X _70095_/Y _70096_/X sky130_fd_sc_hd__a211o_4
X_86959_ _86965_/CLK _86959_/D _86959_/Q sky130_fd_sc_hd__dfxtp_4
X_79500_ _79494_/A _79494_/B _79499_/Y _79500_/Y sky130_fd_sc_hd__a21boi_4
X_41015_ _40991_/X _81715_/Q _41014_/X _41016_/A sky130_fd_sc_hd__o21a_4
X_76712_ _76712_/A _76711_/Y _76713_/B sky130_fd_sc_hd__xor2_4
X_49660_ _49632_/A _49660_/X sky130_fd_sc_hd__buf_2
X_73924_ _73916_/Y _73917_/Y _73923_/X _73924_/Y sky130_fd_sc_hd__o21ai_4
X_58858_ _58858_/A _58858_/X sky130_fd_sc_hd__buf_2
X_46872_ _46860_/X _51031_/B _46872_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_919_0_CLK clkbuf_9_459_0_CLK/X _86576_/CLK sky130_fd_sc_hd__clkbuf_1
X_77692_ _77689_/Y _77692_/B _77692_/Y sky130_fd_sc_hd__nor2_4
X_48611_ _48605_/Y _48585_/X _48610_/X _48611_/Y sky130_fd_sc_hd__a21oi_4
X_79431_ _79417_/Y _79422_/Y _79430_/X _79431_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_8_0_CLK clkbuf_9_4_0_CLK/X _85180_/CLK sky130_fd_sc_hd__clkbuf_1
X_45823_ _57217_/B _45823_/Y sky130_fd_sc_hd__inv_2
X_57809_ _57872_/A _57809_/X sky130_fd_sc_hd__buf_2
X_76643_ _76643_/A _76642_/Y _76645_/A sky130_fd_sc_hd__nand2_4
X_49591_ _86359_/Q _49579_/X _49590_/Y _49591_/Y sky130_fd_sc_hd__o21ai_4
X_73855_ _73829_/X _66084_/B _73855_/X sky130_fd_sc_hd__and2_4
X_58789_ _58787_/X _86096_/Q _58788_/X _58789_/Y sky130_fd_sc_hd__o21ai_4
X_48542_ _48642_/A _48542_/B _48542_/Y sky130_fd_sc_hd__nand2_4
X_60820_ _60820_/A _60820_/B _60820_/Y sky130_fd_sc_hd__nand2_4
X_72806_ _72806_/A _72806_/X sky130_fd_sc_hd__buf_2
X_79362_ _84803_/Q _66435_/A _79362_/X sky130_fd_sc_hd__xor2_4
X_45754_ _45752_/Y _45734_/X _45720_/X _45753_/Y _45754_/X sky130_fd_sc_hd__a211o_4
X_76574_ _81278_/Q _81546_/Q _76574_/Y sky130_fd_sc_hd__nand2_4
X_42966_ _40418_/X _42962_/X _66795_/B _42963_/X _87626_/D sky130_fd_sc_hd__a2bb2o_4
X_73786_ _72829_/A _73786_/X sky130_fd_sc_hd__buf_2
X_70998_ _70990_/A _71082_/B _70990_/C _70998_/Y sky130_fd_sc_hd__nand3_4
X_78313_ _82786_/Q _78312_/X _82754_/D sky130_fd_sc_hd__xor2_4
X_44705_ _44705_/A _44705_/Y sky130_fd_sc_hd__inv_2
X_75525_ _75523_/X _75524_/Y _75525_/X sky130_fd_sc_hd__and2_4
X_41917_ _41917_/A _41917_/Y sky130_fd_sc_hd__inv_2
X_60751_ _60558_/X _60761_/A sky130_fd_sc_hd__buf_2
X_48473_ _48473_/A _48485_/B _48473_/Y sky130_fd_sc_hd__nand2_4
X_72737_ _72737_/A _72737_/X sky130_fd_sc_hd__buf_2
X_79293_ _79277_/X _79280_/Y _79293_/X sky130_fd_sc_hd__or2_4
X_45685_ _45452_/A _45685_/X sky130_fd_sc_hd__buf_2
X_42897_ _42895_/X _42896_/X _41656_/X _87662_/Q _42881_/X _42898_/A
+ sky130_fd_sc_hd__o32ai_4
X_47424_ _47565_/A _47466_/C sky130_fd_sc_hd__buf_2
X_78244_ _78234_/Y _78237_/X _78252_/A _78244_/Y sky130_fd_sc_hd__a21boi_4
X_44636_ _41027_/Y _44618_/X _87023_/Q _44619_/X _87023_/D sky130_fd_sc_hd__a2bb2o_4
X_63470_ _63466_/Y _63455_/X _63469_/Y _63470_/Y sky130_fd_sc_hd__a21oi_4
X_75456_ _75456_/A _75457_/C sky130_fd_sc_hd__inv_2
X_41848_ _40755_/A _41848_/X sky130_fd_sc_hd__buf_2
X_60682_ _60682_/A _60804_/C sky130_fd_sc_hd__buf_2
X_72668_ _72668_/A _72668_/B _55467_/X _72668_/Y sky130_fd_sc_hd__nand3_4
X_62421_ _62406_/A _62421_/B _62421_/C _62421_/D _62421_/Y sky130_fd_sc_hd__nand4_4
X_74407_ _74404_/Y _74405_/X _74406_/X _83073_/D sky130_fd_sc_hd__a21oi_4
X_47355_ _47355_/A _47355_/Y sky130_fd_sc_hd__inv_2
X_71619_ _71603_/Y _83436_/Q _71618_/Y _83436_/D sky130_fd_sc_hd__a21o_4
X_78175_ _78167_/A _78172_/A _78175_/X sky130_fd_sc_hd__and2_4
X_44567_ _44567_/A _44567_/X sky130_fd_sc_hd__buf_2
X_75387_ _75362_/X _75359_/X _75404_/B sky130_fd_sc_hd__nand2_4
X_41779_ _41778_/X _41750_/X _88151_/Q _41751_/X _88151_/D sky130_fd_sc_hd__a2bb2o_4
X_72599_ _72522_/Y _72551_/X _72539_/Y _72597_/Y _72598_/Y _72599_/Y
+ sky130_fd_sc_hd__a41oi_4
X_46306_ _46610_/A _48499_/A sky130_fd_sc_hd__buf_2
X_65140_ _64915_/X _65126_/Y _65139_/Y _65140_/Y sky130_fd_sc_hd__o21ai_4
X_77126_ _77126_/A _77125_/X _77130_/A sky130_fd_sc_hd__nand2_4
X_43518_ _43518_/A _43518_/X sky130_fd_sc_hd__buf_2
X_74338_ _74338_/A _74338_/B _55801_/D _74338_/Y sky130_fd_sc_hd__nand3_4
X_62352_ _62345_/X _62347_/X _62351_/Y _84744_/Q _62300_/X _62352_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47286_ _47382_/A _47286_/X sky130_fd_sc_hd__buf_2
X_44498_ _44549_/A _44498_/X sky130_fd_sc_hd__buf_2
X_49025_ _53852_/B _49025_/X sky130_fd_sc_hd__buf_2
X_61303_ _61302_/Y _72563_/C sky130_fd_sc_hd__buf_2
X_46237_ _46237_/A _73939_/A sky130_fd_sc_hd__buf_2
X_65071_ _84216_/Q _65072_/C sky130_fd_sc_hd__inv_2
XPHY_490 sky130_fd_sc_hd__decap_3
X_77057_ _77041_/C _77053_/Y _77056_/Y _77057_/X sky130_fd_sc_hd__o21a_4
X_43449_ _43518_/A _43449_/X sky130_fd_sc_hd__buf_2
X_62283_ _62267_/A _62267_/B _84421_/Q _62283_/Y sky130_fd_sc_hd__nor3_4
X_74269_ _88340_/Q _72899_/X _73898_/X _74269_/X sky130_fd_sc_hd__o21a_4
X_64022_ _64074_/A _64074_/B _64022_/C _64022_/Y sky130_fd_sc_hd__nor3_4
X_76008_ _76008_/A _76005_/C _76009_/B sky130_fd_sc_hd__and2_4
X_61234_ _61234_/A _61250_/B _84502_/Q _61234_/Y sky130_fd_sc_hd__nor3_4
X_46168_ _46166_/A _46170_/C _46107_/A _46168_/Y sky130_fd_sc_hd__a21oi_4
X_45119_ _45114_/Y _45118_/Y _45063_/X _45119_/X sky130_fd_sc_hd__a21o_4
X_68830_ _73989_/A _68757_/X _68731_/X _68829_/Y _68830_/X sky130_fd_sc_hd__a211o_4
X_61165_ _61165_/A _61165_/B _61165_/C _61165_/Y sky130_fd_sc_hd__nor3_4
X_46099_ _80653_/Q _46099_/X sky130_fd_sc_hd__buf_2
X_60116_ _62534_/A _62193_/A sky130_fd_sc_hd__buf_2
X_49927_ _49923_/Y _49924_/X _49926_/X _86298_/D sky130_fd_sc_hd__a21oi_4
X_68761_ _68756_/X _68760_/X _68684_/X _68761_/X sky130_fd_sc_hd__a21o_4
X_65973_ _65685_/X _86236_/Q _65701_/X _65972_/X _65973_/X sky130_fd_sc_hd__a211o_4
X_61096_ _61083_/B _61096_/X sky130_fd_sc_hd__buf_2
X_77959_ _77954_/B _77954_/A _77960_/C sky130_fd_sc_hd__nand2_4
X_67712_ _81490_/D _67688_/X _67711_/X _67712_/X sky130_fd_sc_hd__a21bo_4
X_64924_ _64924_/A _86421_/Q _64924_/X sky130_fd_sc_hd__and2_4
X_60047_ _60064_/A _60081_/B _60047_/C _60047_/Y sky130_fd_sc_hd__nor3_4
X_49858_ _49856_/Y _49844_/X _49857_/X _86311_/D sky130_fd_sc_hd__a21oi_4
X_80970_ _80931_/CLK _75648_/X _80958_/D sky130_fd_sc_hd__dfxtp_4
X_68692_ _68692_/A _68693_/B sky130_fd_sc_hd__inv_2
X_48809_ _48836_/A _48809_/X sky130_fd_sc_hd__buf_2
X_67643_ _87974_/Q _67591_/X _67641_/X _67642_/X _67643_/X sky130_fd_sc_hd__a211o_4
X_79629_ _79629_/A _79629_/B _79629_/X sky130_fd_sc_hd__xor2_4
X_64855_ _64855_/A _64854_/X _64855_/Y sky130_fd_sc_hd__nand2_4
X_49789_ _49807_/A _49802_/B _49789_/C _53003_/D _49789_/X sky130_fd_sc_hd__and4_4
X_51820_ _51820_/A _46740_/X _51820_/Y sky130_fd_sc_hd__nand2_4
X_63806_ _60915_/X _63858_/B sky130_fd_sc_hd__buf_2
X_82640_ _82642_/CLK _82640_/D _78928_/A sky130_fd_sc_hd__dfxtp_4
X_67574_ _67571_/X _67573_/X _67502_/X _67577_/A sky130_fd_sc_hd__a21o_4
X_64786_ _64782_/X _64867_/B _64785_/X _64786_/Y sky130_fd_sc_hd__nand3_4
X_61998_ _61712_/X _61999_/B sky130_fd_sc_hd__buf_2
X_69313_ _69300_/X _69109_/X _69311_/Y _69312_/Y _69313_/X sky130_fd_sc_hd__a211o_4
X_66525_ _66522_/Y _59756_/X _66524_/X _84106_/D sky130_fd_sc_hd__a21o_4
X_51751_ _51745_/Y _51391_/X _51750_/X _51751_/Y sky130_fd_sc_hd__a21oi_4
X_63737_ _60882_/X _63738_/C sky130_fd_sc_hd__buf_2
X_82571_ _82570_/CLK _82571_/D _82571_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_2_2_1_CLK clkbuf_2_2_1_CLK/A clkbuf_2_2_2_CLK/A sky130_fd_sc_hd__clkbuf_1
X_60949_ _60864_/X _64182_/D sky130_fd_sc_hd__buf_2
X_84310_ _84314_/CLK _84310_/D _80422_/B sky130_fd_sc_hd__dfxtp_4
X_50702_ _50682_/A _50188_/B _50702_/Y sky130_fd_sc_hd__nand2_4
X_81522_ _81756_/CLK _81522_/D _81522_/Q sky130_fd_sc_hd__dfxtp_4
X_69244_ _83938_/Q _69230_/X _69243_/X _69244_/X sky130_fd_sc_hd__a21bo_4
X_54470_ _85436_/Q _54457_/X _54469_/Y _54470_/Y sky130_fd_sc_hd__o21ai_4
X_66456_ _84120_/Q _65296_/X _66455_/Y _84120_/D sky130_fd_sc_hd__a21o_4
X_85290_ _80670_/CLK _85290_/D _85290_/Q sky130_fd_sc_hd__dfxtp_4
X_51682_ _85965_/Q _51675_/X _51681_/Y _51682_/Y sky130_fd_sc_hd__o21ai_4
X_63668_ _62126_/D _60780_/X _63357_/X _60766_/X _63667_/Y _63668_/X
+ sky130_fd_sc_hd__a2111o_4
X_53421_ _53417_/Y _53408_/X _53420_/X _85637_/D sky130_fd_sc_hd__a21oi_4
X_65407_ _65407_/A _65407_/X sky130_fd_sc_hd__buf_2
X_84241_ _84241_/CLK _84241_/D _79629_/B sky130_fd_sc_hd__dfxtp_4
X_50633_ _86163_/Q _50626_/X _50632_/Y _50633_/Y sky130_fd_sc_hd__o21ai_4
X_62619_ _61685_/A _62597_/B _59913_/A _62597_/D _62619_/Y sky130_fd_sc_hd__nand4_4
X_69175_ _83943_/Q _69161_/X _69174_/X _69175_/X sky130_fd_sc_hd__a21bo_4
X_81453_ _81433_/CLK _76753_/B _81453_/Q sky130_fd_sc_hd__dfxtp_4
X_66387_ _66046_/A _66389_/A sky130_fd_sc_hd__buf_2
X_63599_ _61558_/B _63548_/X _63597_/X _63598_/Y _63599_/X sky130_fd_sc_hd__a211o_4
X_80404_ _80393_/X _80404_/B _80404_/X sky130_fd_sc_hd__and2_4
X_68126_ _68121_/X _66791_/Y _68110_/X _68125_/Y _68126_/X sky130_fd_sc_hd__a211o_4
X_56140_ _56140_/A _56140_/B _85289_/Q _56140_/Y sky130_fd_sc_hd__nand3_4
X_53352_ _53352_/A _53353_/A sky130_fd_sc_hd__buf_2
X_65338_ _65211_/X _85509_/Q _65212_/X _65337_/X _65338_/X sky130_fd_sc_hd__a211o_4
X_84172_ _81233_/CLK _84172_/D _84172_/Q sky130_fd_sc_hd__dfxtp_4
X_50564_ _50534_/A _50607_/A sky130_fd_sc_hd__buf_2
X_81384_ _83918_/CLK _81384_/D _76847_/B sky130_fd_sc_hd__dfxtp_4
Xpsn_inst_psn_buff_7 _71216_/A _71233_/A2 sky130_fd_sc_hd__buf_2
X_52303_ _52299_/A _48963_/X _52303_/Y sky130_fd_sc_hd__nand2_4
X_83123_ _86213_/CLK _83123_/D _70128_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_250_0_CLK clkbuf_8_251_0_CLK/A clkbuf_9_501_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_56071_ _56052_/A _56086_/B _55879_/B _56071_/Y sky130_fd_sc_hd__nand3_4
X_80335_ _80333_/Y _80336_/A sky130_fd_sc_hd__inv_2
X_68057_ _68057_/A _68377_/A sky130_fd_sc_hd__buf_2
X_53283_ _53311_/A _53293_/A sky130_fd_sc_hd__buf_2
X_65269_ _65267_/Y _65195_/X _65268_/X _84208_/D sky130_fd_sc_hd__a21o_4
X_50495_ _86189_/Q _50464_/X _50494_/Y _50495_/Y sky130_fd_sc_hd__o21ai_4
X_55022_ _55037_/A _47639_/Y _55022_/Y sky130_fd_sc_hd__nand2_4
X_67008_ _66961_/X _86788_/Q _67008_/X sky130_fd_sc_hd__and2_4
X_52234_ _52231_/Y _52232_/X _52233_/X _85863_/D sky130_fd_sc_hd__a21oi_4
X_83054_ _85566_/CLK _83054_/D _83054_/Q sky130_fd_sc_hd__dfxtp_4
X_87931_ _82886_/CLK _87931_/D _87931_/Q sky130_fd_sc_hd__dfxtp_4
X_80266_ _80265_/Y _80266_/B _80266_/Y sky130_fd_sc_hd__nand2_4
X_82005_ _82005_/CLK _82005_/D _77134_/A sky130_fd_sc_hd__dfxtp_4
X_59830_ _60175_/A _60353_/B _60312_/C _60312_/D _59830_/Y sky130_fd_sc_hd__nand4_4
X_52165_ _52198_/A _52194_/B sky130_fd_sc_hd__buf_2
X_87862_ _87348_/CLK _87862_/D _87862_/Q sky130_fd_sc_hd__dfxtp_4
X_80197_ _80209_/A _80209_/B _80197_/Y sky130_fd_sc_hd__xnor2_4
X_51116_ _51113_/Y _51093_/X _51115_/X _51116_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_260_0_CLK clkbuf_9_130_0_CLK/X _83457_/CLK sky130_fd_sc_hd__clkbuf_1
X_86813_ _81154_/CLK _46017_/X _67179_/B sky130_fd_sc_hd__dfxtp_4
X_59761_ _59761_/A _59761_/B _59761_/X sky130_fd_sc_hd__and2_4
X_56973_ _57043_/B _56971_/Y _56664_/Y _56972_/Y _56973_/X sky130_fd_sc_hd__a2bb2o_4
X_52096_ _65423_/B _52089_/X _52095_/Y _52096_/Y sky130_fd_sc_hd__o21ai_4
X_68959_ _68746_/A _68959_/B _68959_/Y sky130_fd_sc_hd__nor2_4
X_87793_ _87553_/CLK _42639_/Y _87793_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_890_0_CLK clkbuf_9_445_0_CLK/X _85542_/CLK sky130_fd_sc_hd__clkbuf_1
X_58712_ _58641_/X _85941_/Q _58664_/X _58712_/X sky130_fd_sc_hd__o21a_4
X_51047_ _51101_/A _51047_/X sky130_fd_sc_hd__buf_2
X_55924_ _55949_/A _56041_/C _55924_/X sky130_fd_sc_hd__and2_4
X_86744_ _85529_/CLK _86744_/D _86744_/Q sky130_fd_sc_hd__dfxtp_4
X_71970_ _71970_/A _71970_/B _71970_/Y sky130_fd_sc_hd__nand2_4
X_83956_ _83957_/CLK _83956_/D _83956_/Q sky130_fd_sc_hd__dfxtp_4
X_59692_ _59648_/A _59692_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_42_0_CLK clkbuf_9_21_0_CLK/X _83846_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_9_381_0_CLK clkbuf_8_190_0_CLK/X clkbuf_9_381_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_58643_ _58625_/X _85467_/Q _58642_/X _58643_/Y sky130_fd_sc_hd__o21ai_4
X_70921_ _70869_/A _70914_/B _70914_/C _70919_/D _70921_/Y sky130_fd_sc_hd__nand4_4
X_82907_ _87922_/CLK _78261_/B _41661_/A sky130_fd_sc_hd__dfxtp_4
X_55855_ _44079_/X _55855_/B _55855_/X sky130_fd_sc_hd__and2_4
X_86675_ _86353_/CLK _86675_/D _86675_/Q sky130_fd_sc_hd__dfxtp_4
X_83887_ _82339_/CLK _83887_/D _81959_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_275_0_CLK clkbuf_9_137_0_CLK/X _83761_/CLK sky130_fd_sc_hd__clkbuf_1
X_42820_ _51949_/A _42820_/X sky130_fd_sc_hd__buf_2
X_54806_ _85374_/Q _54784_/X _54805_/Y _54806_/Y sky130_fd_sc_hd__o21ai_4
X_73640_ _73637_/X _73639_/X _73612_/X _73643_/A sky130_fd_sc_hd__a21o_4
X_85626_ _85630_/CLK _53494_/Y _85626_/Q sky130_fd_sc_hd__dfxtp_4
X_70852_ _70905_/A _70890_/B _70852_/C _70860_/D _70852_/Y sky130_fd_sc_hd__nand4_4
X_58574_ _58570_/Y _58573_/Y _58105_/X _58574_/X sky130_fd_sc_hd__a21o_4
X_82838_ _84177_/CLK _82838_/D _82838_/Q sky130_fd_sc_hd__dfxtp_4
X_55786_ _85195_/Q _55747_/X _55300_/X _55785_/X _55786_/X sky130_fd_sc_hd__a211o_4
X_52998_ _52996_/Y _52975_/X _52997_/X _52998_/Y sky130_fd_sc_hd__a21oi_4
X_57525_ _47917_/A _49317_/X _46603_/X _57525_/X sky130_fd_sc_hd__and3_4
X_88345_ _88345_/CLK _40735_/X _69004_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_57_0_CLK clkbuf_9_28_0_CLK/X _85103_/CLK sky130_fd_sc_hd__clkbuf_1
X_42751_ _42739_/X _42740_/X _41245_/X _87739_/Q _42750_/X _42752_/A
+ sky130_fd_sc_hd__o32ai_4
X_54737_ _85387_/Q _54729_/X _54736_/Y _54737_/Y sky130_fd_sc_hd__o21ai_4
X_85557_ _85557_/CLK _53845_/Y _85557_/Q sky130_fd_sc_hd__dfxtp_4
X_73571_ _47830_/Y _73570_/Y _73572_/B sky130_fd_sc_hd__xor2_4
X_51949_ _51949_/A _52618_/A sky130_fd_sc_hd__buf_2
X_70783_ _70848_/A _70791_/B sky130_fd_sc_hd__buf_2
X_82769_ _82769_/CLK _82769_/D _82769_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_396_0_CLK clkbuf_8_198_0_CLK/X clkbuf_9_396_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_75310_ _80786_/Q _81042_/D _80754_/D sky130_fd_sc_hd__xor2_4
X_41702_ _41701_/X _41682_/X _67659_/B _41684_/X _88166_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_203_0_CLK clkbuf_8_203_0_CLK/A clkbuf_9_407_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_72522_ _61368_/D _72516_/A _72607_/C _72563_/C _72522_/Y sky130_fd_sc_hd__nand4_4
X_84508_ _84508_/CLK _84508_/D _61203_/C sky130_fd_sc_hd__dfxtp_4
X_45470_ _45470_/A _45470_/Y sky130_fd_sc_hd__inv_2
X_57456_ _57440_/X _57454_/X _57455_/Y _57456_/Y sky130_fd_sc_hd__o21ai_4
X_76290_ _81644_/Q _76290_/B _76309_/B sky130_fd_sc_hd__xnor2_4
X_42682_ _41059_/X _42679_/X _87773_/Q _42681_/X _87773_/D sky130_fd_sc_hd__a2bb2o_4
X_88276_ _88283_/CLK _41111_/X _69558_/B sky130_fd_sc_hd__dfxtp_4
X_54668_ _54665_/Y _54666_/X _54667_/X _54668_/Y sky130_fd_sc_hd__a21oi_4
X_85488_ _83736_/CLK _54187_/Y _85488_/Q sky130_fd_sc_hd__dfxtp_4
X_44421_ _41560_/X _44412_/X _87116_/Q _44413_/X _87116_/D sky130_fd_sc_hd__a2bb2o_4
X_56407_ _56397_/X _56399_/B _56407_/C _56407_/Y sky130_fd_sc_hd__nand3_4
X_75241_ _75237_/X _75240_/X _75241_/Y sky130_fd_sc_hd__xnor2_4
X_87227_ _87487_/CLK _43867_/Y _87227_/Q sky130_fd_sc_hd__dfxtp_4
X_53619_ _53747_/A _53619_/X sky130_fd_sc_hd__buf_2
X_41633_ _41632_/Y _88179_/D sky130_fd_sc_hd__inv_2
X_72453_ _72450_/Y _72452_/Y _57779_/X _72453_/X sky130_fd_sc_hd__a21o_4
X_84439_ _84441_/CLK _62018_/Y _78062_/B sky130_fd_sc_hd__dfxtp_4
X_57387_ _57384_/X _56575_/X _85023_/Q _57385_/X _57387_/X sky130_fd_sc_hd__a2bb2o_4
X_54599_ _54597_/Y _54584_/X _54598_/X _85413_/D sky130_fd_sc_hd__a21oi_4
X_47140_ _47140_/A _47143_/C sky130_fd_sc_hd__buf_2
X_71404_ _70676_/A _71404_/B _71411_/C _71404_/Y sky130_fd_sc_hd__nor3_4
X_59126_ _59061_/X _86071_/Q _59125_/X _59126_/Y sky130_fd_sc_hd__o21ai_4
X_44352_ _44624_/A _44352_/X sky130_fd_sc_hd__buf_2
X_56338_ _56351_/A _56345_/B sky130_fd_sc_hd__buf_2
X_75172_ _75175_/B _75172_/Y sky130_fd_sc_hd__inv_2
X_87158_ _87471_/CLK _87158_/D _87158_/Q sky130_fd_sc_hd__dfxtp_4
X_41564_ _41533_/X _40489_/A _41563_/X _41564_/X sky130_fd_sc_hd__o21a_4
X_72384_ _72384_/A _72428_/B _72384_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_8_218_0_CLK clkbuf_8_219_0_CLK/A clkbuf_8_218_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_43303_ _41203_/X _43300_/X _87490_/Q _43302_/X _87490_/D sky130_fd_sc_hd__a2bb2o_4
X_74123_ _74123_/A _73195_/A _74123_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_213_0_CLK clkbuf_9_106_0_CLK/X _84645_/CLK sky130_fd_sc_hd__clkbuf_1
X_86109_ _84807_/CLK _86109_/D _86109_/Q sky130_fd_sc_hd__dfxtp_4
X_40515_ _40514_/X _40515_/X sky130_fd_sc_hd__buf_2
X_47071_ _47063_/A _52837_/B _47071_/Y sky130_fd_sc_hd__nand2_4
X_59057_ _59057_/A _59008_/B _59057_/Y sky130_fd_sc_hd__nor2_4
X_71335_ _71335_/A _71335_/B _71313_/X _71335_/Y sky130_fd_sc_hd__nand3_4
X_56269_ _56245_/A _56270_/B sky130_fd_sc_hd__buf_2
X_44283_ _44282_/X _57650_/A sky130_fd_sc_hd__buf_2
X_79980_ _79980_/A _79980_/B _79982_/A sky130_fd_sc_hd__nand2_4
X_87089_ _88267_/CLK _44476_/X _87089_/Q sky130_fd_sc_hd__dfxtp_4
X_41495_ _41494_/Y _88205_/D sky130_fd_sc_hd__inv_2
Xclkbuf_10_843_0_CLK clkbuf_9_421_0_CLK/X _84166_/CLK sky130_fd_sc_hd__clkbuf_1
X_58008_ _57989_/X _58005_/Y _58006_/Y _58007_/X _57993_/X _58008_/X
+ sky130_fd_sc_hd__o32a_4
X_46022_ _45962_/X _46022_/X sky130_fd_sc_hd__buf_2
X_43234_ _43234_/A _43234_/Y sky130_fd_sc_hd__inv_2
X_74054_ _68888_/B _73872_/X _73920_/X _74053_/Y _74054_/X sky130_fd_sc_hd__a211o_4
X_78931_ _78919_/A _78931_/B _78931_/X sky130_fd_sc_hd__and2_4
X_40446_ _40445_/X _40446_/X sky130_fd_sc_hd__buf_2
X_71266_ _71266_/A _70733_/Y _71266_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_334_0_CLK clkbuf_9_335_0_CLK/A clkbuf_9_334_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_73005_ _73001_/X _73004_/X _72951_/X _73021_/B sky130_fd_sc_hd__a21o_4
X_70217_ _70232_/A _70229_/B sky130_fd_sc_hd__buf_2
X_43165_ _43014_/Y _43166_/A sky130_fd_sc_hd__buf_2
X_78862_ _78862_/A _78862_/B _78862_/X sky130_fd_sc_hd__xor2_4
X_40377_ _40376_/Y _40377_/Y sky130_fd_sc_hd__inv_2
X_71197_ _71197_/A _71076_/B _71197_/C _71197_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_228_0_CLK clkbuf_9_114_0_CLK/X _81859_/CLK sky130_fd_sc_hd__clkbuf_1
X_42116_ _42077_/A _42116_/X sky130_fd_sc_hd__buf_2
X_77813_ _77813_/A _77828_/A sky130_fd_sc_hd__inv_2
X_70148_ _83527_/Q _83175_/Q _83526_/Q _83174_/Q _70148_/Y sky130_fd_sc_hd__a22oi_4
X_47973_ _47973_/A _47973_/B _47973_/X sky130_fd_sc_hd__or2_4
X_59959_ _62475_/A _62621_/D sky130_fd_sc_hd__buf_2
X_43096_ _87577_/Q _43096_/Y sky130_fd_sc_hd__inv_2
X_78793_ _78793_/A _78793_/B _78794_/A sky130_fd_sc_hd__xor2_4
Xclkbuf_10_858_0_CLK clkbuf_9_429_0_CLK/X _86121_/CLK sky130_fd_sc_hd__clkbuf_1
X_49712_ _49657_/A _49724_/C sky130_fd_sc_hd__buf_2
X_46924_ _82401_/Q _46924_/Y sky130_fd_sc_hd__inv_2
X_42047_ _88058_/Q _42047_/Y sky130_fd_sc_hd__inv_2
X_77744_ _82147_/Q _77744_/B _82115_/D sky130_fd_sc_hd__xor2_4
X_62970_ _62968_/X _62942_/X _62969_/Y _62970_/Y sky130_fd_sc_hd__a21oi_4
X_74956_ _80945_/Q _74956_/B _81194_/D sky130_fd_sc_hd__xor2_4
X_70079_ _70079_/A _70078_/X _59787_/X _70079_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_9_349_0_CLK clkbuf_8_174_0_CLK/X clkbuf_9_349_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_49643_ _49639_/Y _49623_/X _49642_/X _49643_/Y sky130_fd_sc_hd__a21oi_4
X_61921_ _61479_/B _61953_/B _61860_/C _61860_/D _61921_/Y sky130_fd_sc_hd__nand4_4
X_73907_ _72829_/A _73907_/X sky130_fd_sc_hd__buf_2
X_46855_ _82952_/Q _46856_/A sky130_fd_sc_hd__inv_2
X_77675_ _77675_/A _77675_/Y sky130_fd_sc_hd__inv_2
X_74887_ _74887_/A _74887_/B _74887_/C _74887_/Y sky130_fd_sc_hd__nand3_4
X_79414_ _79414_/A _79414_/B _79414_/X sky130_fd_sc_hd__xor2_4
X_45806_ _45748_/X _61640_/A _45765_/X _45806_/Y sky130_fd_sc_hd__o21ai_4
X_64640_ _64611_/A _85823_/Q _64640_/X sky130_fd_sc_hd__and2_4
X_76626_ _76625_/Y _76623_/A _76640_/A sky130_fd_sc_hd__nand2_4
X_49574_ _49558_/A _52787_/B _49574_/Y sky130_fd_sc_hd__nand2_4
X_61852_ _61711_/X _61871_/A sky130_fd_sc_hd__buf_2
X_73838_ _73836_/X _73838_/B _73838_/C _73838_/Y sky130_fd_sc_hd__nand3_4
X_46786_ _46786_/A _54364_/B sky130_fd_sc_hd__inv_2
X_43998_ _43998_/A _59516_/A sky130_fd_sc_hd__buf_2
X_48525_ _83578_/Q _74437_/B sky130_fd_sc_hd__inv_2
X_60803_ _84563_/Q _60673_/X _60754_/X _60750_/X _60803_/Y sky130_fd_sc_hd__a2bb2oi_4
X_79345_ _79341_/Y _79344_/Y _79355_/B sky130_fd_sc_hd__xor2_4
X_45737_ _45733_/Y _45734_/X _45720_/X _45736_/Y _45737_/X sky130_fd_sc_hd__a211o_4
X_64571_ _64642_/A _64571_/X sky130_fd_sc_hd__buf_2
X_76557_ _76557_/A _76560_/B sky130_fd_sc_hd__inv_2
X_42949_ _42949_/A _42949_/Y sky130_fd_sc_hd__inv_2
X_61783_ _61770_/X _61773_/X _61782_/Y _84918_/Q _61719_/X _61783_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73769_ _70107_/C _73697_/X _73768_/X _73769_/Y sky130_fd_sc_hd__o21ai_4
X_66310_ _66237_/X _66310_/B _66310_/X sky130_fd_sc_hd__and2_4
X_63522_ _63398_/A _63523_/A sky130_fd_sc_hd__buf_2
X_75508_ _75508_/A _75508_/B _75510_/A sky130_fd_sc_hd__or2_4
X_48456_ _48469_/A _50440_/B _48456_/Y sky130_fd_sc_hd__nand2_4
X_60734_ _84578_/Q _60673_/X _60733_/Y _60723_/X _60734_/Y sky130_fd_sc_hd__a2bb2oi_4
X_67290_ _67266_/A _67290_/B _67290_/X sky130_fd_sc_hd__and2_4
X_79276_ _79266_/X _79276_/B _79276_/Y sky130_fd_sc_hd__nand2_4
X_45668_ _45668_/A _45668_/X sky130_fd_sc_hd__buf_2
X_76488_ _76489_/A _81541_/Q _76491_/B sky130_fd_sc_hd__nor2_4
X_47407_ _47407_/A _53031_/D sky130_fd_sc_hd__buf_2
X_66241_ _66235_/X _66239_/X _66240_/X _66244_/A sky130_fd_sc_hd__a21o_4
X_78227_ _82583_/Q _82495_/Q _78230_/A sky130_fd_sc_hd__xor2_4
X_44619_ _44603_/A _44619_/X sky130_fd_sc_hd__buf_2
X_75439_ _75466_/B _75438_/Y _75440_/B sky130_fd_sc_hd__xor2_4
X_63453_ _64292_/A _63465_/B _63465_/C _63465_/D _63453_/Y sky130_fd_sc_hd__nand4_4
X_48387_ _74375_/A _48388_/A sky130_fd_sc_hd__buf_2
X_60665_ _59539_/A _59705_/X _60665_/C _62640_/C _60665_/X sky130_fd_sc_hd__or4_4
X_45599_ _45599_/A _45599_/Y sky130_fd_sc_hd__inv_2
X_62404_ _62475_/A _62404_/X sky130_fd_sc_hd__buf_2
X_47338_ _47198_/X _47380_/A sky130_fd_sc_hd__buf_2
X_66172_ _66117_/X _84975_/Q _64707_/X _66171_/X _66173_/C sky130_fd_sc_hd__a211o_4
X_78158_ _78151_/Y _78152_/A _78157_/Y _78159_/B sky130_fd_sc_hd__a21boi_4
X_63384_ _63410_/A _63384_/B _63384_/C _63384_/D _63384_/X sky130_fd_sc_hd__and4_4
X_60596_ _60596_/A _60596_/B _60596_/Y sky130_fd_sc_hd__nor2_4
X_65123_ _65116_/X _65121_/X _65122_/X _65126_/A sky130_fd_sc_hd__a21o_4
X_77109_ _77109_/A _77109_/B _77110_/B sky130_fd_sc_hd__xor2_4
X_62335_ _62362_/A _62335_/B _62335_/C _62335_/D _62335_/Y sky130_fd_sc_hd__nand4_4
X_47269_ _47241_/X _52950_/B _47269_/Y sky130_fd_sc_hd__nand2_4
X_78089_ _78089_/A _78090_/B sky130_fd_sc_hd__inv_2
X_49008_ _86453_/Q _49003_/X _49007_/Y _49008_/Y sky130_fd_sc_hd__o21ai_4
X_80120_ _80114_/Y _80119_/Y _81684_/D sky130_fd_sc_hd__xor2_4
X_65054_ _65319_/A _65054_/B _65054_/X sky130_fd_sc_hd__and2_4
X_69931_ _73462_/A _69833_/X _69617_/X _69930_/Y _69931_/X sky130_fd_sc_hd__a211o_4
X_50280_ _50279_/X _53504_/B _50280_/Y sky130_fd_sc_hd__nand2_4
X_62266_ _62179_/X _62267_/B sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_14 _55686_/C _56647_/A4 sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_25 _41869_/Y _50212_/A sky130_fd_sc_hd__buf_8
X_64005_ _64053_/A _58434_/A _64071_/C _64005_/X sky130_fd_sc_hd__and3_4
X_61217_ _61169_/X _61214_/Y _61216_/Y _84506_/Q _59509_/X _61217_/X
+ sky130_fd_sc_hd__o32a_4
X_80051_ _80047_/X _80050_/Y _80073_/B sky130_fd_sc_hd__xor2_4
X_69862_ _69908_/A _69862_/B _69862_/Y sky130_fd_sc_hd__nor2_4
X_62197_ _62195_/Y _59951_/C _84729_/Q _62196_/X _62197_/X sky130_fd_sc_hd__a2bb2o_4
X_68813_ _68542_/X _87745_/Q _68813_/X sky130_fd_sc_hd__and2_4
X_61148_ _64210_/A _61147_/Y _61148_/X sky130_fd_sc_hd__and2_4
X_69793_ _69766_/A _69793_/B _69793_/Y sky130_fd_sc_hd__nor2_4
X_83810_ _83813_/CLK _83810_/D _74722_/A sky130_fd_sc_hd__dfxtp_4
X_68744_ _43068_/A _68414_/X _68741_/X _68743_/X _68744_/X sky130_fd_sc_hd__a211o_4
X_53970_ _53967_/Y _53892_/X _53969_/X _53970_/Y sky130_fd_sc_hd__a21oi_4
X_65956_ _65954_/Y _65915_/X _65955_/X _84166_/D sky130_fd_sc_hd__a21o_4
X_61079_ _61079_/A _61079_/Y sky130_fd_sc_hd__inv_2
X_84790_ _86695_/CLK _84790_/D _84790_/Q sky130_fd_sc_hd__dfxtp_4
X_52921_ _52893_/X _52922_/A sky130_fd_sc_hd__buf_2
X_64907_ _64828_/X _85558_/Q _64829_/X _64906_/X _64907_/X sky130_fd_sc_hd__a211o_4
X_83741_ _86322_/CLK _83741_/D _47334_/A sky130_fd_sc_hd__dfxtp_4
X_80953_ _81211_/CLK _80965_/Q _80953_/Q sky130_fd_sc_hd__dfxtp_4
X_68675_ _69651_/A _68750_/A sky130_fd_sc_hd__buf_2
X_65887_ _84171_/Q _65888_/C sky130_fd_sc_hd__inv_2
X_55640_ _55640_/A _55640_/Y sky130_fd_sc_hd__inv_2
X_67626_ _67675_/A _87655_/Q _67626_/X sky130_fd_sc_hd__and2_4
X_86460_ _85562_/CLK _48941_/Y _64759_/B sky130_fd_sc_hd__dfxtp_4
X_52852_ _52852_/A _52853_/B sky130_fd_sc_hd__buf_2
X_64838_ _64832_/X _64888_/B _64837_/X _64838_/Y sky130_fd_sc_hd__nand3_4
X_83672_ _83673_/CLK _70891_/Y _46778_/A sky130_fd_sc_hd__dfxtp_4
X_80884_ _80854_/CLK _75741_/B _80852_/D sky130_fd_sc_hd__dfxtp_4
X_85411_ _85635_/CLK _54608_/Y _85411_/Q sky130_fd_sc_hd__dfxtp_4
X_51803_ _53282_/A _51804_/A sky130_fd_sc_hd__buf_2
X_82623_ _82715_/CLK _82623_/D _82623_/Q sky130_fd_sc_hd__dfxtp_4
X_55571_ _55507_/X _55571_/X sky130_fd_sc_hd__buf_2
X_67557_ _87914_/Q _67533_/X _67508_/X _67556_/X _67557_/X sky130_fd_sc_hd__a211o_4
X_86391_ _83681_/CLK _86391_/D _58687_/B sky130_fd_sc_hd__dfxtp_4
X_52783_ _52783_/A _52783_/X sky130_fd_sc_hd__buf_2
X_64769_ _64769_/A _86267_/Q _64769_/X sky130_fd_sc_hd__and2_4
X_57310_ _57310_/A _85037_/D sky130_fd_sc_hd__inv_2
X_88130_ _88386_/CLK _88130_/D _66978_/B sky130_fd_sc_hd__dfxtp_4
X_54522_ _54509_/A _54526_/B _54509_/C _54522_/D _54522_/X sky130_fd_sc_hd__and4_4
X_66508_ _60371_/X _66315_/Y _66507_/Y _66508_/Y sky130_fd_sc_hd__o21ai_4
X_85342_ _85342_/CLK _54980_/Y _85342_/Q sky130_fd_sc_hd__dfxtp_4
X_51734_ _52593_/A _52588_/A sky130_fd_sc_hd__buf_2
X_58290_ _83406_/Q _58290_/Y sky130_fd_sc_hd__inv_2
X_82554_ _82558_/CLK _83874_/Q _82554_/Q sky130_fd_sc_hd__dfxtp_4
X_67488_ _87469_/Q _67394_/X _67462_/X _67487_/X _67488_/X sky130_fd_sc_hd__a211o_4
X_81505_ _81322_/CLK _81505_/D _81505_/Q sky130_fd_sc_hd__dfxtp_4
X_57241_ _44288_/X _56578_/X _45444_/A _57238_/X _85054_/D sky130_fd_sc_hd__a2bb2o_4
X_69227_ _68532_/X _68536_/X _69212_/X _69227_/Y sky130_fd_sc_hd__a21oi_4
X_88061_ _87813_/CLK _42040_/Y _73320_/A sky130_fd_sc_hd__dfxtp_4
X_54453_ _54399_/A _54453_/X sky130_fd_sc_hd__buf_2
X_66439_ _66435_/Y _64532_/X _66438_/X _84123_/D sky130_fd_sc_hd__o21ai_4
X_85273_ _85177_/CLK _56215_/Y _85273_/Q sky130_fd_sc_hd__dfxtp_4
X_51665_ _51671_/A _53187_/B _51665_/Y sky130_fd_sc_hd__nand2_4
X_82485_ _82485_/CLK _78594_/X _78154_/B sky130_fd_sc_hd__dfxtp_4
X_87012_ _87333_/CLK _87012_/D _87012_/Q sky130_fd_sc_hd__dfxtp_4
X_53404_ _53351_/A _53404_/X sky130_fd_sc_hd__buf_2
X_84224_ _81227_/CLK _64871_/X _84224_/Q sky130_fd_sc_hd__dfxtp_4
X_50616_ _50613_/Y _50577_/X _50615_/Y _50616_/Y sky130_fd_sc_hd__a21boi_4
X_57172_ _57169_/X _57170_/Y _74342_/A _57172_/Y sky130_fd_sc_hd__a21oi_4
X_81436_ _82648_/CLK _81468_/Q _76126_/C sky130_fd_sc_hd__dfxtp_4
X_69158_ _68407_/X _68410_/X _69061_/X _69158_/Y sky130_fd_sc_hd__a21oi_4
X_54384_ _54245_/A _54385_/A sky130_fd_sc_hd__buf_2
X_51596_ _51617_/A _53122_/B _51596_/Y sky130_fd_sc_hd__nand2_4
X_56123_ _56123_/A _56140_/B sky130_fd_sc_hd__buf_2
X_68109_ _84037_/Q _68101_/X _68108_/X _68109_/X sky130_fd_sc_hd__a21bo_4
X_53335_ _53333_/Y _53328_/X _53334_/X _53335_/Y sky130_fd_sc_hd__a21oi_4
X_84155_ _84166_/CLK _84155_/D _80481_/B sky130_fd_sc_hd__dfxtp_4
X_50547_ _48691_/A _50552_/B _50552_/C _50547_/X sky130_fd_sc_hd__and3_4
X_81367_ _81352_/CLK _81367_/D _81367_/Q sky130_fd_sc_hd__dfxtp_4
X_69089_ _69661_/A _69089_/B _69089_/Y sky130_fd_sc_hd__nor2_4
X_71120_ _49125_/X _71117_/X _71119_/Y _71120_/Y sky130_fd_sc_hd__o21ai_4
X_83106_ _83095_/CLK _83106_/D _83106_/Q sky130_fd_sc_hd__dfxtp_4
X_80318_ _80318_/A _80317_/B _80318_/Y sky130_fd_sc_hd__nand2_4
X_56054_ _56044_/X _56054_/B _56055_/A sky130_fd_sc_hd__xnor2_4
X_41280_ _81698_/Q _41280_/B _41280_/X sky130_fd_sc_hd__or2_4
X_53266_ _51914_/A _53274_/B _53266_/C _52750_/D _53266_/X sky130_fd_sc_hd__and4_4
X_84086_ _83918_/CLK _67045_/X _80910_/D sky130_fd_sc_hd__dfxtp_4
X_50478_ _86193_/Q _50464_/X _50477_/Y _50478_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_7_64_0_CLK clkbuf_6_32_0_CLK/X clkbuf_7_64_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_81298_ _81362_/CLK _76986_/X _81298_/Q sky130_fd_sc_hd__dfxtp_4
X_55005_ _55013_/A _55026_/B _55013_/C _55005_/D _55005_/X sky130_fd_sc_hd__and4_4
X_52217_ _85866_/Q _52214_/X _52216_/Y _52217_/Y sky130_fd_sc_hd__o21ai_4
X_71051_ _48878_/B _71047_/X _71050_/Y _71051_/Y sky130_fd_sc_hd__o21ai_4
X_83037_ _85213_/CLK _74556_/Y _44966_/A sky130_fd_sc_hd__dfxtp_4
X_87914_ _87653_/CLK _87914_/D _87914_/Q sky130_fd_sc_hd__dfxtp_4
X_80249_ _80247_/Y _80243_/X _80251_/A sky130_fd_sc_hd__nand2_4
X_53197_ _53194_/Y _53189_/X _53196_/X _85679_/D sky130_fd_sc_hd__a21oi_4
X_70002_ _69650_/X _69653_/X _70001_/X _70002_/Y sky130_fd_sc_hd__a21oi_4
X_59813_ _57689_/A _60341_/A sky130_fd_sc_hd__buf_2
X_52148_ _52127_/X _48763_/B _52148_/Y sky130_fd_sc_hd__nand2_4
X_87845_ _88097_/CLK _87845_/D _68727_/A sky130_fd_sc_hd__dfxtp_4
X_74810_ _74810_/A _74810_/B _74810_/C _74810_/D _74810_/Y sky130_fd_sc_hd__nand4_4
X_59744_ _59743_/Y _59754_/A _59816_/A _59744_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_7_79_0_CLK clkbuf_7_78_0_CLK/A clkbuf_7_79_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_44970_ _44966_/Y _45033_/B _44970_/Y sky130_fd_sc_hd__nand2_4
X_52079_ _52083_/A _52079_/B _52079_/Y sky130_fd_sc_hd__nand2_4
X_56956_ _56949_/X _56607_/X _45501_/A _56947_/X _85114_/D sky130_fd_sc_hd__a2bb2o_4
X_75790_ _75778_/Y _75779_/Y _80920_/Q _75781_/Y _75790_/X sky130_fd_sc_hd__a2bb2o_4
X_87776_ _87776_/CLK _87776_/D _87776_/Q sky130_fd_sc_hd__dfxtp_4
X_84988_ _84991_/CLK _84988_/D _84988_/Q sky130_fd_sc_hd__dfxtp_4
X_43921_ _41397_/X _43907_/X _67845_/B _43908_/X _87198_/D sky130_fd_sc_hd__a2bb2o_4
X_55907_ _55904_/X _55906_/X _44118_/B _55907_/X sky130_fd_sc_hd__a21o_4
X_74741_ _71753_/D _71268_/A _74735_/X _74736_/X _74740_/Y _74741_/X
+ sky130_fd_sc_hd__a2111o_4
X_86727_ _86119_/CLK _86727_/D _86727_/Q sky130_fd_sc_hd__dfxtp_4
X_71953_ _74531_/A _70766_/C _71349_/D _71894_/Y _71953_/Y sky130_fd_sc_hd__nand4_4
X_59675_ _66262_/A _66514_/B sky130_fd_sc_hd__buf_2
X_83939_ _81352_/CLK _69229_/X _83939_/Q sky130_fd_sc_hd__dfxtp_4
X_56887_ _56753_/A _56887_/B _56887_/Y sky130_fd_sc_hd__nand2_4
X_70904_ _51003_/B _70885_/A _70903_/Y _70904_/Y sky130_fd_sc_hd__o21ai_4
X_46640_ _46636_/Y _46598_/X _46639_/X _86719_/D sky130_fd_sc_hd__a21oi_4
X_58626_ _57997_/X _85948_/Q _58109_/X _58626_/X sky130_fd_sc_hd__o21a_4
X_77460_ _77459_/X _77460_/Y sky130_fd_sc_hd__inv_2
X_43852_ _43846_/X _43824_/X _41209_/X _68815_/B _43847_/X _43852_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55838_ _55836_/A _56510_/C _55838_/X sky130_fd_sc_hd__and2_4
X_74672_ _74672_/A _74672_/Y sky130_fd_sc_hd__inv_2
X_86658_ _86340_/CLK _47219_/Y _59377_/A sky130_fd_sc_hd__dfxtp_4
X_71884_ _71871_/X _59437_/B _71883_/Y _83341_/D sky130_fd_sc_hd__a21o_4
X_76411_ _76410_/Y _76411_/Y sky130_fd_sc_hd__inv_2
X_42803_ _42822_/A _42803_/X sky130_fd_sc_hd__buf_2
X_73623_ _70125_/A _86754_/D _73622_/X _83143_/D sky130_fd_sc_hd__o21ai_4
X_85609_ _86535_/CLK _85609_/D _85609_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_142_0_CLK clkbuf_7_71_0_CLK/X clkbuf_9_285_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_46571_ _46566_/Y _46523_/X _46570_/Y _86725_/D sky130_fd_sc_hd__a21boi_4
X_70835_ _70848_/A _70846_/B sky130_fd_sc_hd__buf_2
X_58557_ _58557_/A _58557_/B _58557_/Y sky130_fd_sc_hd__nand2_4
X_77391_ _77382_/A _77382_/B _77381_/A _77417_/A sky130_fd_sc_hd__o21a_4
X_55769_ _55159_/A _85289_/Q _55769_/X sky130_fd_sc_hd__and2_4
X_43783_ _43782_/Y _43783_/Y sky130_fd_sc_hd__inv_2
X_86589_ _86237_/CLK _47888_/Y _86589_/Q sky130_fd_sc_hd__dfxtp_4
X_40995_ _40995_/A _40995_/X sky130_fd_sc_hd__buf_2
X_48310_ _48319_/A _48310_/B _48310_/Y sky130_fd_sc_hd__nand2_4
X_79130_ _79130_/A _79130_/B _82438_/D sky130_fd_sc_hd__xor2_4
X_57508_ _57504_/Y _57506_/X _57507_/X _57508_/Y sky130_fd_sc_hd__a21oi_4
X_45522_ _45519_/Y _45489_/X _45520_/X _45521_/Y _45522_/X sky130_fd_sc_hd__a211o_4
X_76342_ _76356_/A _76342_/B _81615_/D sky130_fd_sc_hd__xor2_4
X_88328_ _87063_/CLK _40823_/X _88328_/Q sky130_fd_sc_hd__dfxtp_4
X_42734_ _42734_/A _87745_/D sky130_fd_sc_hd__inv_2
X_49290_ _49288_/Y _49271_/X _49289_/Y _49290_/Y sky130_fd_sc_hd__a21boi_4
X_73554_ _73554_/A _73577_/B _73554_/Y sky130_fd_sc_hd__nor2_4
X_70766_ _70860_/A _70779_/B _70766_/C _70769_/D _70766_/Y sky130_fd_sc_hd__nand4_4
X_58488_ _58467_/X _58485_/Y _58487_/Y _84837_/D sky130_fd_sc_hd__a21oi_4
X_48241_ _48169_/X _48241_/X sky130_fd_sc_hd__buf_2
X_72505_ _61302_/A _72503_/A _72535_/B sky130_fd_sc_hd__nand2_4
X_79061_ _79059_/X _79060_/Y _82717_/D sky130_fd_sc_hd__nand2_4
X_45453_ _45434_/X _61367_/A _45452_/X _45453_/Y sky130_fd_sc_hd__o21ai_4
X_57439_ _57439_/A _85004_/D sky130_fd_sc_hd__inv_2
X_76273_ _76273_/A _76272_/Y _81610_/D sky130_fd_sc_hd__xnor2_4
X_88259_ _87103_/CLK _88259_/D _68775_/B sky130_fd_sc_hd__dfxtp_4
X_42665_ _42590_/A _42665_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_17_0_CLK clkbuf_6_8_0_CLK/X clkbuf_8_35_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_73485_ _42057_/Y _72888_/X _72890_/X _73484_/Y _73485_/X sky130_fd_sc_hd__a211o_4
X_70697_ _70935_/A _70698_/B sky130_fd_sc_hd__inv_2
X_78012_ _78012_/A _78012_/Y sky130_fd_sc_hd__inv_2
X_44404_ _44381_/A _44404_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_157_0_CLK clkbuf_7_78_0_CLK/X clkbuf_9_315_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_75224_ _75224_/A _75224_/Y sky130_fd_sc_hd__inv_2
X_41616_ _41615_/X _41616_/X sky130_fd_sc_hd__buf_2
X_48172_ _48171_/X _50048_/A sky130_fd_sc_hd__buf_2
X_60450_ _60404_/Y _60588_/A sky130_fd_sc_hd__buf_2
X_72436_ _72414_/X _72436_/B _72436_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_152_0_CLK clkbuf_9_76_0_CLK/X _81631_/CLK sky130_fd_sc_hd__clkbuf_1
X_45384_ _45350_/X _61692_/B _45370_/X _45384_/Y sky130_fd_sc_hd__o21ai_4
X_42596_ _42596_/A _42596_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_782_0_CLK clkbuf_9_391_0_CLK/X _82702_/CLK sky130_fd_sc_hd__clkbuf_1
X_59109_ _59104_/Y _59108_/Y _58939_/X _59109_/X sky130_fd_sc_hd__a21o_4
X_47123_ _83699_/Q _53386_/B sky130_fd_sc_hd__inv_2
X_44335_ _41663_/X _44326_/X _87161_/Q _44327_/X _44335_/X sky130_fd_sc_hd__a2bb2o_4
X_75155_ _75151_/Y _75153_/Y _75154_/Y _75155_/Y sky130_fd_sc_hd__o21ai_4
X_41547_ _41547_/A _88195_/D sky130_fd_sc_hd__inv_2
X_60381_ _60381_/A _60447_/A sky130_fd_sc_hd__buf_2
X_72367_ _57790_/X _72401_/B sky130_fd_sc_hd__buf_2
X_62120_ _62120_/A _62144_/A sky130_fd_sc_hd__buf_2
X_74106_ _72908_/A _74106_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_273_0_CLK clkbuf_8_136_0_CLK/X clkbuf_9_273_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_47054_ _47063_/A _52829_/B _47054_/Y sky130_fd_sc_hd__nand2_4
X_71318_ _70454_/Y _71319_/B sky130_fd_sc_hd__buf_2
X_44266_ _44006_/X _44164_/X _44266_/C _44266_/Y sky130_fd_sc_hd__nand3_4
X_79963_ _79963_/A _79958_/A _79957_/Y _79963_/Y sky130_fd_sc_hd__nand3_4
X_75086_ _75086_/A _75079_/B _75086_/Y sky130_fd_sc_hd__nor2_4
X_41478_ _41449_/X _82333_/Q _41477_/X _41478_/Y sky130_fd_sc_hd__o21ai_4
X_72298_ _72286_/Y _72237_/X _72293_/X _72297_/X _83267_/D sky130_fd_sc_hd__a22oi_4
X_46005_ _45994_/X _46001_/X _40490_/X _86818_/Q _45995_/X _46006_/A
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_10_167_0_CLK clkbuf_9_83_0_CLK/X _81668_/CLK sky130_fd_sc_hd__clkbuf_1
X_43217_ _43217_/A _43218_/A sky130_fd_sc_hd__buf_2
X_62051_ _61820_/A _62090_/B sky130_fd_sc_hd__buf_2
X_74037_ _86987_/Q _73916_/B _74036_/X _74048_/C sky130_fd_sc_hd__o21ai_4
X_78914_ _78899_/Y _78913_/X _78914_/Y sky130_fd_sc_hd__nand2_4
X_40429_ _49140_/B _40429_/X sky130_fd_sc_hd__buf_2
X_71249_ _50232_/B _71239_/X _71248_/Y _71249_/Y sky130_fd_sc_hd__o21ai_4
X_44197_ _44196_/X _56953_/A sky130_fd_sc_hd__buf_2
X_79894_ _79531_/X _79532_/Y _79895_/B sky130_fd_sc_hd__nand2_4
Xclkbuf_10_797_0_CLK clkbuf_9_398_0_CLK/X _84115_/CLK sky130_fd_sc_hd__clkbuf_1
X_61002_ _60952_/X _60993_/Y _60995_/Y _60999_/X _61001_/X _84543_/D
+ sky130_fd_sc_hd__o41a_4
X_43148_ _43147_/Y _87558_/D sky130_fd_sc_hd__inv_2
X_78845_ _82726_/Q _78845_/B _78845_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_9_288_0_CLK clkbuf_8_144_0_CLK/X clkbuf_9_288_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_65810_ _65805_/X _65808_/X _65809_/X _65810_/X sky130_fd_sc_hd__a21o_4
X_47956_ _47904_/X _46380_/A _47955_/X _47957_/B sky130_fd_sc_hd__o21ai_4
X_43079_ _43053_/X _43054_/X _40696_/X _43078_/Y _43058_/X _43079_/Y
+ sky130_fd_sc_hd__o32ai_4
X_66790_ _87126_/Q _66715_/X _66717_/X _66789_/X _66790_/X sky130_fd_sc_hd__a211o_4
X_78776_ _78788_/A _82700_/Q _78777_/B sky130_fd_sc_hd__xor2_4
X_75988_ _81708_/D _81420_/Q _76005_/A sky130_fd_sc_hd__xor2_4
Xclkbuf_10_720_0_CLK clkbuf_9_360_0_CLK/X _88272_/CLK sky130_fd_sc_hd__clkbuf_1
X_46907_ _46901_/Y _46891_/X _46906_/X _86691_/D sky130_fd_sc_hd__a21oi_4
X_65741_ _65737_/X _65741_/B _65740_/X _65742_/B sky130_fd_sc_hd__nand3_4
X_77727_ _77725_/Y _78044_/A _77728_/B sky130_fd_sc_hd__xor2_4
X_74939_ _74942_/B _74939_/B _74940_/B sky130_fd_sc_hd__xnor2_4
X_62953_ _62988_/A _62988_/B _84367_/Q _62953_/Y sky130_fd_sc_hd__nor3_4
X_47887_ _47887_/A _47886_/X _47887_/X sky130_fd_sc_hd__and2_4
X_49626_ _49622_/Y _49623_/X _49625_/X _86353_/D sky130_fd_sc_hd__a21oi_4
X_61904_ _59605_/Y _61949_/C sky130_fd_sc_hd__buf_2
Xclkbuf_9_211_0_CLK clkbuf_9_210_0_CLK/A clkbuf_9_211_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_68460_ _83974_/Q _68338_/X _68459_/X _83974_/D sky130_fd_sc_hd__a21bo_4
X_46838_ _46830_/A _46830_/B _46830_/C _52704_/D _46838_/X sky130_fd_sc_hd__and4_4
X_65672_ _65668_/X _65671_/X _65642_/X _65676_/A sky130_fd_sc_hd__a21o_4
X_77658_ _77657_/X _77658_/Y sky130_fd_sc_hd__inv_2
X_62884_ _58487_/A _62841_/X _60197_/C _60202_/A _62884_/Y sky130_fd_sc_hd__nand4_4
X_67411_ _67364_/X _67411_/B _67411_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_105_0_CLK clkbuf_9_52_0_CLK/X _87169_/CLK sky130_fd_sc_hd__clkbuf_1
X_64623_ _64623_/A _64622_/X _64623_/Y sky130_fd_sc_hd__nand2_4
X_76609_ _76605_/X _76604_/Y _76609_/Y sky130_fd_sc_hd__nand2_4
X_49557_ _49555_/Y _49541_/X _49556_/X _86366_/D sky130_fd_sc_hd__a21oi_4
X_61835_ _61865_/A _61865_/B _78074_/B _61835_/Y sky130_fd_sc_hd__nor3_4
X_68391_ _68382_/X _68388_/X _68390_/X _68391_/X sky130_fd_sc_hd__a21o_4
X_46769_ _46769_/A _52663_/B sky130_fd_sc_hd__inv_2
X_77589_ _77584_/X _77587_/Y _77585_/Y _77590_/B sky130_fd_sc_hd__nand3_4
Xclkbuf_10_735_0_CLK clkbuf_9_367_0_CLK/X _88097_/CLK sky130_fd_sc_hd__clkbuf_1
X_48508_ _48508_/A _48485_/B _48508_/Y sky130_fd_sc_hd__nand2_4
X_79328_ _58792_/Y _66457_/Y _79327_/Y _79346_/A sky130_fd_sc_hd__o21a_4
X_67342_ _67342_/A _87667_/Q _67342_/X sky130_fd_sc_hd__and2_4
X_64554_ _61232_/X _61692_/B _61207_/X _64554_/Y sky130_fd_sc_hd__nand3_4
X_49488_ _49407_/A _49500_/A sky130_fd_sc_hd__buf_2
X_61766_ _61782_/A _61766_/B _61761_/Y _61766_/D _61766_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_9_226_0_CLK clkbuf_8_113_0_CLK/X clkbuf_9_226_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_63505_ _59403_/A _63491_/B _63514_/C _63491_/D _63505_/Y sky130_fd_sc_hd__nand4_4
X_48439_ _48043_/X _48958_/B _48438_/Y _48440_/A sky130_fd_sc_hd__o21ai_4
X_60717_ _60700_/A _60752_/B _60717_/C _60717_/Y sky130_fd_sc_hd__nor3_4
X_67273_ _87926_/Q _67176_/X _67271_/X _67272_/X _67273_/X sky130_fd_sc_hd__a211o_4
X_79259_ _79259_/A _83217_/Q _79260_/B sky130_fd_sc_hd__xor2_4
X_64485_ _61232_/X _61617_/B _61207_/X _64485_/Y sky130_fd_sc_hd__nand3_4
X_61697_ _61697_/A _61697_/Y sky130_fd_sc_hd__inv_2
X_69012_ _87481_/Q _68989_/X _69010_/X _69011_/X _69012_/X sky130_fd_sc_hd__a211o_4
X_66224_ _66221_/X _66223_/X _66057_/X _66224_/X sky130_fd_sc_hd__a21o_4
X_51450_ _52688_/A _51504_/A sky130_fd_sc_hd__buf_2
X_63436_ _63436_/A _63436_/X sky130_fd_sc_hd__buf_2
X_82270_ _82272_/CLK _82270_/D _82270_/Q sky130_fd_sc_hd__dfxtp_4
X_60648_ _60662_/A _60724_/B sky130_fd_sc_hd__buf_2
X_50401_ _52103_/A _50430_/B _50338_/X _50401_/X sky130_fd_sc_hd__and3_4
X_81221_ _84197_/CLK _81029_/Q _81221_/Q sky130_fd_sc_hd__dfxtp_4
X_66155_ _64694_/A _66155_/B _66155_/X sky130_fd_sc_hd__and2_4
X_51381_ _51379_/Y _51366_/X _51380_/X _51381_/Y sky130_fd_sc_hd__a21oi_4
X_63367_ _63357_/X _63368_/A sky130_fd_sc_hd__buf_2
X_60579_ _79136_/A _60577_/X _60578_/Y _60586_/D _84596_/D sky130_fd_sc_hd__a2bb2oi_4
X_53120_ _53172_/A _53120_/X sky130_fd_sc_hd__buf_2
X_65106_ _65035_/X _85518_/Q _65036_/X _65105_/X _65106_/X sky130_fd_sc_hd__a211o_4
X_50332_ _50329_/Y _50313_/X _50331_/X _50332_/Y sky130_fd_sc_hd__a21oi_4
X_62318_ _62203_/Y _62319_/A sky130_fd_sc_hd__buf_2
X_81152_ _81211_/CLK _80744_/Q _40571_/A sky130_fd_sc_hd__dfxtp_4
X_66086_ _66083_/X _66085_/X _65304_/X _66426_/A sky130_fd_sc_hd__a21o_4
X_63298_ _58976_/A _62999_/X _61636_/B _60608_/X _63298_/Y sky130_fd_sc_hd__a2bb2oi_4
X_80103_ _80101_/X _80108_/B _80103_/Y sky130_fd_sc_hd__xnor2_4
X_65037_ _65002_/A _65037_/B _65037_/X sky130_fd_sc_hd__and2_4
X_53051_ _85706_/Q _53038_/X _53050_/Y _53051_/Y sky130_fd_sc_hd__o21ai_4
X_69914_ _69499_/Y _69732_/X _69870_/X _69913_/Y _69914_/X sky130_fd_sc_hd__a211o_4
X_50263_ _50261_/Y _50227_/X _50262_/Y _50263_/Y sky130_fd_sc_hd__a21boi_4
X_62249_ _62249_/A _63384_/B _59987_/X _62251_/C sky130_fd_sc_hd__nand3_4
X_85960_ _85961_/CLK _85960_/D _85960_/Q sky130_fd_sc_hd__dfxtp_4
X_81083_ _81117_/CLK _75650_/A _81083_/Q sky130_fd_sc_hd__dfxtp_4
X_52002_ _66094_/B _51994_/X _52001_/Y _52002_/Y sky130_fd_sc_hd__o21ai_4
X_84911_ _84555_/CLK _58195_/Y _62124_/B sky130_fd_sc_hd__dfxtp_4
X_80034_ _80021_/X _80032_/X _80033_/X _80034_/Y sky130_fd_sc_hd__a21oi_4
X_69845_ _69413_/X _69416_/X _69816_/X _69845_/Y sky130_fd_sc_hd__a21oi_4
X_50194_ _50189_/Y _50191_/X _50193_/X _86246_/D sky130_fd_sc_hd__a21oi_4
X_85891_ _86490_/CLK _85891_/D _66334_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_opt_21_CLK _85555_/CLK _83300_/CLK sky130_fd_sc_hd__clkbuf_16
X_56810_ _56816_/A _56810_/X sky130_fd_sc_hd__buf_2
X_87630_ _87625_/CLK _87630_/D _66698_/B sky130_fd_sc_hd__dfxtp_4
X_84842_ _84299_/CLK _58466_/Y _84842_/Q sky130_fd_sc_hd__dfxtp_4
X_57790_ _64621_/A _57790_/X sky130_fd_sc_hd__buf_2
X_69776_ _87811_/Q _69776_/Y sky130_fd_sc_hd__inv_2
X_66988_ _66868_/A _66988_/X sky130_fd_sc_hd__buf_2
X_56741_ _56726_/X _56738_/X _56739_/X _56740_/X _45957_/A _56741_/Y
+ sky130_fd_sc_hd__a41oi_4
X_68727_ _68727_/A _68727_/Y sky130_fd_sc_hd__inv_2
X_87561_ _88326_/CLK _43140_/Y _73036_/A sky130_fd_sc_hd__dfxtp_4
X_53953_ _53949_/A _53953_/B _53953_/Y sky130_fd_sc_hd__nand2_4
X_65939_ _65896_/A _65939_/B _65939_/X sky130_fd_sc_hd__and2_4
X_84773_ _86686_/CLK _84773_/D _84773_/Q sky130_fd_sc_hd__dfxtp_4
X_81985_ _81985_/CLK _81985_/D _81985_/Q sky130_fd_sc_hd__dfxtp_4
X_86512_ _86498_/CLK _86512_/D _86512_/Q sky130_fd_sc_hd__dfxtp_4
X_52904_ _52903_/X _52910_/A sky130_fd_sc_hd__buf_2
X_59460_ _59460_/A _59444_/X _59460_/Y sky130_fd_sc_hd__nand2_4
X_83724_ _85375_/CLK _70687_/X _47497_/A sky130_fd_sc_hd__dfxtp_4
X_56672_ _83329_/Q _56672_/Y sky130_fd_sc_hd__inv_2
X_68658_ _68735_/A _68658_/B _68658_/X sky130_fd_sc_hd__and2_4
X_80936_ _80962_/CLK _75151_/B _80936_/Q sky130_fd_sc_hd__dfxtp_4
X_87492_ _87758_/CLK _43298_/Y _87492_/Q sky130_fd_sc_hd__dfxtp_4
X_53884_ _52365_/A _53875_/B _53888_/C _53884_/X sky130_fd_sc_hd__and3_4
X_58411_ _84855_/Q _58412_/A sky130_fd_sc_hd__inv_2
X_55623_ _83007_/Q _55689_/A _44102_/A _55622_/X _55624_/B sky130_fd_sc_hd__a211o_4
X_67609_ _87156_/Q _67585_/X _67516_/X _67608_/X _67609_/X sky130_fd_sc_hd__a211o_4
X_86443_ _85538_/CLK _86443_/D _86443_/Q sky130_fd_sc_hd__dfxtp_4
X_52835_ _52818_/A _52831_/B _52818_/C _52835_/D _52835_/X sky130_fd_sc_hd__and4_4
X_83655_ _85536_/CLK _70946_/Y _46270_/A sky130_fd_sc_hd__dfxtp_4
X_59391_ _59390_/Y _59392_/A sky130_fd_sc_hd__buf_2
X_80867_ _80818_/CLK _75587_/B _80835_/D sky130_fd_sc_hd__dfxtp_4
X_68589_ _68587_/X _68588_/Y _68589_/Y sky130_fd_sc_hd__nor2_4
X_70620_ _70724_/A _70620_/B _70620_/C _70620_/D _70620_/Y sky130_fd_sc_hd__nand4_4
X_58342_ _58342_/A _58342_/Y sky130_fd_sc_hd__inv_2
X_82606_ _82575_/CLK _78920_/B _82606_/Q sky130_fd_sc_hd__dfxtp_4
X_55554_ _45501_/A _55511_/X _55506_/X _55553_/Y _55554_/X sky130_fd_sc_hd__a211o_4
X_86374_ _83663_/CLK _86374_/D _86374_/Q sky130_fd_sc_hd__dfxtp_4
X_40780_ _40773_/X _82302_/Q _40779_/X _40780_/Y sky130_fd_sc_hd__o21ai_4
X_52766_ _52630_/A _52767_/A sky130_fd_sc_hd__buf_2
X_83586_ _85593_/CLK _83586_/D _83586_/Q sky130_fd_sc_hd__dfxtp_4
X_80798_ _80991_/CLK _80798_/D _75514_/A sky130_fd_sc_hd__dfxtp_4
X_88113_ _88108_/CLK _41884_/Y _73595_/A sky130_fd_sc_hd__dfxtp_4
X_54505_ _54486_/X _53332_/B _54505_/Y sky130_fd_sc_hd__nand2_4
X_85325_ _85354_/CLK _85325_/D _85325_/Q sky130_fd_sc_hd__dfxtp_4
X_51717_ _51717_/A _53240_/B _51717_/Y sky130_fd_sc_hd__nand2_4
X_70551_ _70533_/X _83751_/Q _70550_/Y _83751_/D sky130_fd_sc_hd__a21o_4
X_58273_ _58273_/A _58280_/B sky130_fd_sc_hd__buf_2
X_82537_ _82536_/CLK _82537_/D _82537_/Q sky130_fd_sc_hd__dfxtp_4
X_55485_ _85042_/Q _55468_/X _55458_/X _55484_/Y _55485_/X sky130_fd_sc_hd__a211o_4
X_52697_ _85771_/Q _52684_/X _52696_/Y _52697_/Y sky130_fd_sc_hd__o21ai_4
X_57224_ _57123_/Y _57220_/Y _57221_/X _57223_/X _85060_/D sky130_fd_sc_hd__a211o_4
X_88044_ _88044_/CLK _88044_/D _88044_/Q sky130_fd_sc_hd__dfxtp_4
X_42450_ _42449_/Y _42579_/A sky130_fd_sc_hd__inv_2
X_54436_ _54434_/Y _54422_/X _54435_/X _85443_/D sky130_fd_sc_hd__a21oi_4
X_73270_ _73268_/X _73270_/B _73270_/C _73270_/Y sky130_fd_sc_hd__nand3_4
X_85256_ _85190_/CLK _85256_/D _85256_/Q sky130_fd_sc_hd__dfxtp_4
X_51648_ _50222_/X _51671_/A sky130_fd_sc_hd__buf_2
X_70482_ DATA_TO_HASH[2] _71435_/C sky130_fd_sc_hd__buf_2
X_82468_ _82942_/CLK _78341_/X _78262_/B sky130_fd_sc_hd__dfxtp_4
X_41401_ _41743_/B _41379_/X _41401_/X sky130_fd_sc_hd__or2_4
X_72221_ _86617_/Q _72162_/B _72221_/Y sky130_fd_sc_hd__nor2_4
X_84207_ _84220_/CLK _84207_/D _65294_/C sky130_fd_sc_hd__dfxtp_4
X_57155_ _57141_/X _56739_/X _56800_/X _57155_/D _57158_/A sky130_fd_sc_hd__and4_4
X_81419_ _84049_/CLK _81451_/Q _75991_/B sky130_fd_sc_hd__dfxtp_4
X_42381_ _42378_/X _42369_/X _41791_/X _87892_/Q _42370_/X _42382_/A
+ sky130_fd_sc_hd__o32ai_4
X_54367_ _54362_/A _54362_/B _54362_/C _46790_/Y _54367_/X sky130_fd_sc_hd__and4_4
X_85187_ _85186_/CLK _56455_/Y _56454_/C sky130_fd_sc_hd__dfxtp_4
X_51579_ _51552_/A _51603_/C sky130_fd_sc_hd__buf_2
X_82399_ _82965_/CLK _82207_/Q _82399_/Q sky130_fd_sc_hd__dfxtp_4
X_44120_ _44091_/Y _44102_/X _44119_/Y _44120_/Y sky130_fd_sc_hd__a21oi_4
X_56106_ _56082_/X _56103_/X _56105_/Y _56106_/Y sky130_fd_sc_hd__o21ai_4
X_41332_ _41331_/X _41332_/X sky130_fd_sc_hd__buf_2
X_53318_ _53298_/A _47016_/A _53318_/Y sky130_fd_sc_hd__nand2_4
X_72152_ _72358_/A _72152_/X sky130_fd_sc_hd__buf_2
X_84138_ _82177_/CLK _84138_/D _84138_/Q sky130_fd_sc_hd__dfxtp_4
X_57086_ _57126_/A _57086_/X sky130_fd_sc_hd__buf_2
X_54298_ _54312_/A _54298_/B _54312_/C _54298_/D _54298_/X sky130_fd_sc_hd__and4_4
X_71103_ _50144_/B _71095_/X _71102_/Y _83607_/D sky130_fd_sc_hd__o21ai_4
X_44051_ _44051_/A _44052_/A sky130_fd_sc_hd__buf_2
X_56037_ _56023_/A _56052_/B _55934_/B _56037_/Y sky130_fd_sc_hd__nand3_4
X_41263_ _41261_/X _81702_/Q _41262_/X _41264_/A sky130_fd_sc_hd__o21ai_4
X_53249_ _53243_/X _53244_/B _53266_/C _53249_/D _53249_/X sky130_fd_sc_hd__and4_4
X_72083_ _72083_/A _72083_/X sky130_fd_sc_hd__buf_2
X_76960_ _76804_/Y _81363_/D sky130_fd_sc_hd__inv_2
X_84069_ _81428_/CLK _67448_/X _84069_/Q sky130_fd_sc_hd__dfxtp_4
X_43002_ _40520_/X _42994_/X _87610_/Q _42995_/X _87610_/D sky130_fd_sc_hd__a2bb2o_4
X_71034_ _53161_/B _71013_/X _71033_/Y _71034_/Y sky130_fd_sc_hd__o21ai_4
X_75911_ _61200_/C _62806_/C _80725_/D sky130_fd_sc_hd__xor2_4
X_41194_ _40995_/A _41194_/X sky130_fd_sc_hd__buf_2
X_76891_ _81596_/Q _81468_/D _76891_/X sky130_fd_sc_hd__xor2_4
X_47810_ _47819_/A _53255_/B _47810_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_opt_12_CLK _84914_/CLK _84884_/CLK sky130_fd_sc_hd__clkbuf_16
X_78630_ _78630_/A _82692_/Q _78630_/Y sky130_fd_sc_hd__nand2_4
X_75842_ _75830_/A _75830_/B _75842_/Y sky130_fd_sc_hd__nor2_4
X_87828_ _87288_/CLK _87828_/D _69110_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_14_0_CLK clkbuf_3_7_1_CLK/X clkbuf_4_14_1_CLK/A sky130_fd_sc_hd__clkbuf_1
X_48790_ _48790_/A _48814_/C sky130_fd_sc_hd__buf_2
X_57988_ _57985_/Y _57987_/Y _57889_/X _57988_/X sky130_fd_sc_hd__a21o_4
X_47741_ _83546_/Q _47741_/Y sky130_fd_sc_hd__inv_2
X_59727_ _66377_/A _59727_/X sky130_fd_sc_hd__buf_2
X_78561_ _78561_/A _78561_/B _78561_/Y sky130_fd_sc_hd__nand2_4
X_44953_ _64246_/B _61364_/B sky130_fd_sc_hd__buf_2
X_56939_ _72732_/B _56939_/X sky130_fd_sc_hd__buf_2
X_75773_ _75751_/A _75750_/Y _75761_/Y _75762_/Y _75773_/X sky130_fd_sc_hd__o22a_4
X_87759_ _87260_/CLK _42707_/X _68480_/B sky130_fd_sc_hd__dfxtp_4
X_72985_ _72905_/A _72985_/X sky130_fd_sc_hd__buf_2
X_77512_ _77512_/A _77512_/B _77514_/A sky130_fd_sc_hd__xor2_4
X_43904_ _43903_/Y _87208_/D sky130_fd_sc_hd__inv_2
X_74724_ _70735_/X _74745_/D sky130_fd_sc_hd__buf_2
X_47672_ _49406_/A _49379_/A sky130_fd_sc_hd__buf_2
X_71936_ _74533_/A _74518_/B _71940_/C _71945_/D _71936_/Y sky130_fd_sc_hd__nand4_4
X_59658_ _59582_/A _59660_/C sky130_fd_sc_hd__buf_2
X_78492_ _78488_/Y _78490_/Y _78487_/Y _78492_/Y sky130_fd_sc_hd__o21ai_4
X_44884_ _45389_/A _44884_/X sky130_fd_sc_hd__buf_2
X_49411_ _86392_/Q _49388_/X _49410_/Y _49411_/Y sky130_fd_sc_hd__o21ai_4
X_58609_ _58140_/X _86110_/Q _58608_/X _58609_/Y sky130_fd_sc_hd__o21ai_4
X_46623_ _46623_/A _46651_/A sky130_fd_sc_hd__buf_2
X_77443_ _77443_/A _77447_/A sky130_fd_sc_hd__inv_2
X_43835_ _41157_/X _43832_/X _87243_/Q _43833_/X _43835_/X sky130_fd_sc_hd__a2bb2o_4
X_74655_ _45951_/Y _56642_/Y _82995_/Q _74630_/X _82995_/D sky130_fd_sc_hd__a2bb2o_4
X_71867_ _71867_/A _71867_/B _70884_/B _71711_/A _71867_/Y sky130_fd_sc_hd__nor4_4
X_59589_ _59588_/Y _61948_/A sky130_fd_sc_hd__buf_2
X_49342_ _49327_/X _54075_/B _49342_/Y sky130_fd_sc_hd__nand2_4
X_61620_ _63280_/B _61611_/B _61611_/C _61572_/D _61620_/Y sky130_fd_sc_hd__nand4_4
X_73606_ _73306_/A _73607_/A sky130_fd_sc_hd__buf_2
X_46554_ _83782_/Q _54073_/B sky130_fd_sc_hd__inv_2
X_70818_ _70804_/A _71219_/A sky130_fd_sc_hd__buf_2
X_77374_ _77396_/B _77374_/B _82188_/D sky130_fd_sc_hd__xor2_4
X_43766_ _43766_/A _43766_/Y sky130_fd_sc_hd__inv_2
X_74586_ _45141_/A _74582_/X _74585_/X _83026_/D sky130_fd_sc_hd__o21ai_4
X_40978_ _40944_/X _40946_/X _40977_/X _88299_/Q _40916_/X _40978_/Y
+ sky130_fd_sc_hd__o32ai_4
X_71798_ _70804_/A _71313_/X _71716_/B _71798_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_1007_0_CLK clkbuf_9_503_0_CLK/X _86196_/CLK sky130_fd_sc_hd__clkbuf_1
X_79113_ _79110_/A _82753_/Q _79110_/B _79113_/Y sky130_fd_sc_hd__nand3_4
X_45505_ _55555_/B _45489_/X _45443_/X _45504_/Y _45505_/X sky130_fd_sc_hd__a211o_4
X_76325_ _76325_/A _76324_/Y _76326_/B sky130_fd_sc_hd__xnor2_4
X_42717_ _42651_/X _42717_/X sky130_fd_sc_hd__buf_2
X_61551_ _61551_/A _61542_/B _61542_/C _61512_/X _61551_/Y sky130_fd_sc_hd__nand4_4
X_49273_ _49273_/A _46407_/X _49273_/Y sky130_fd_sc_hd__nand2_4
X_73537_ _73516_/A _86466_/Q _73537_/X sky130_fd_sc_hd__and2_4
X_46485_ _48499_/A _46485_/X sky130_fd_sc_hd__buf_2
X_70749_ _70753_/A _70719_/A _70749_/Y sky130_fd_sc_hd__nand2_4
X_43697_ _40820_/X _43695_/X _73056_/A _43696_/X _43697_/X sky130_fd_sc_hd__a2bb2o_4
X_60502_ _60502_/A _60500_/Y _60501_/Y _60502_/Y sky130_fd_sc_hd__nor3_4
X_48224_ _48204_/X _47932_/B _48224_/Y sky130_fd_sc_hd__nand2_4
X_79044_ _79044_/A _79044_/B _79044_/C _79044_/Y sky130_fd_sc_hd__nand3_4
X_45436_ _45434_/X _61358_/A _45370_/X _45436_/Y sky130_fd_sc_hd__o21ai_4
X_64270_ _64257_/Y _64268_/X _64269_/X _64270_/X sky130_fd_sc_hd__o21a_4
X_76256_ _76253_/Y _76255_/Y _76268_/D sky130_fd_sc_hd__nor2_4
X_42648_ _42592_/A _42648_/X sky130_fd_sc_hd__buf_2
X_61482_ _61482_/A _61481_/X _61482_/C _61482_/Y sky130_fd_sc_hd__nand3_4
X_73468_ _69935_/B _73279_/X _73202_/X _73468_/X sky130_fd_sc_hd__o21a_4
X_63221_ _63218_/Y _63220_/X _63172_/X _63221_/Y sky130_fd_sc_hd__a21oi_4
X_75207_ _75207_/A _75207_/B _75201_/Y _75207_/Y sky130_fd_sc_hd__nand3_4
X_48155_ _86562_/Q _48150_/X _48154_/Y _48155_/Y sky130_fd_sc_hd__o21ai_4
X_60433_ _60433_/A _60417_/A _60438_/A _60443_/A _60516_/B sky130_fd_sc_hd__nand4_4
X_72419_ _57759_/X _72419_/X sky130_fd_sc_hd__buf_2
X_45367_ _64545_/B _61682_/B sky130_fd_sc_hd__buf_2
X_76187_ _76187_/A _81553_/Q _76187_/Y sky130_fd_sc_hd__nand2_4
X_42579_ _42579_/A _42580_/A sky130_fd_sc_hd__buf_2
X_73399_ _88314_/Q _73059_/X _73007_/X _73399_/Y sky130_fd_sc_hd__o21ai_4
X_47106_ _47101_/Y _47081_/X _47105_/X _86670_/D sky130_fd_sc_hd__a21oi_4
X_44318_ _44318_/A _44317_/X _87169_/D sky130_fd_sc_hd__nor2_4
X_63152_ _79385_/A _63130_/X _63151_/Y _84349_/D sky130_fd_sc_hd__a21o_4
X_75138_ _75138_/A _75138_/B _75138_/Y sky130_fd_sc_hd__nor2_4
X_60364_ _60525_/A _60519_/B sky130_fd_sc_hd__buf_2
X_48086_ _48086_/A _48086_/B _48086_/X sky130_fd_sc_hd__or2_4
X_45298_ _55756_/B _45281_/X _45237_/X _45298_/X sky130_fd_sc_hd__o21a_4
X_62103_ _62100_/Y _62101_/X _62102_/Y _62103_/Y sky130_fd_sc_hd__a21oi_4
X_47037_ _82389_/Q _54509_/D sky130_fd_sc_hd__inv_2
X_44249_ _44174_/A _68385_/A sky130_fd_sc_hd__buf_2
X_63083_ _79447_/A _63072_/X _63082_/Y _84355_/D sky130_fd_sc_hd__a21o_4
X_67960_ _86949_/Q _67906_/X _67908_/X _67959_/X _67960_/X sky130_fd_sc_hd__a211o_4
X_75069_ _75067_/Y _75069_/B _75069_/Y sky130_fd_sc_hd__nand2_4
X_79946_ _79946_/A _79934_/A _79946_/Y sky130_fd_sc_hd__nand2_4
X_60295_ _60249_/X _60325_/B _60290_/Y _60337_/A _60294_/Y _60295_/Y
+ sky130_fd_sc_hd__a41oi_4
X_66911_ _66794_/A _66911_/X sky130_fd_sc_hd__buf_2
X_62034_ _62002_/A _62002_/B _78061_/B _62034_/Y sky130_fd_sc_hd__nor3_4
X_67891_ _67891_/A _67891_/B _67891_/X sky130_fd_sc_hd__and2_4
X_79877_ _79861_/X _79865_/B _79876_/X _79877_/X sky130_fd_sc_hd__a21o_4
X_69630_ _69198_/Y _69603_/X _69604_/X _69629_/Y _69630_/X sky130_fd_sc_hd__a211o_4
X_66842_ _87368_/Q _66797_/X _66747_/X _66841_/X _66842_/X sky130_fd_sc_hd__a211o_4
X_78828_ _78828_/A _78828_/B _78828_/C _78828_/Y sky130_fd_sc_hd__nand3_4
X_48988_ _48988_/A _53834_/B sky130_fd_sc_hd__buf_2
X_69561_ _69127_/X _69130_/X _69500_/X _69561_/Y sky130_fd_sc_hd__a21oi_4
X_47939_ _83775_/Q _57537_/B sky130_fd_sc_hd__inv_2
Xclkbuf_9_150_0_CLK clkbuf_8_75_0_CLK/X clkbuf_9_150_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_66773_ _87883_/Q _66697_/X _66675_/X _66772_/X _66773_/X sky130_fd_sc_hd__a211o_4
X_78759_ _78770_/B _78770_/D _78759_/X sky130_fd_sc_hd__and2_4
X_63985_ _63979_/Y _63980_/Y _63981_/Y _63985_/D _63985_/X sky130_fd_sc_hd__and4_4
X_68512_ _68208_/X _68512_/X sky130_fd_sc_hd__buf_2
X_65724_ _65660_/X _83062_/Q _65568_/X _65723_/X _65724_/X sky130_fd_sc_hd__a211o_4
X_50950_ _50938_/X _51812_/B _50950_/Y sky130_fd_sc_hd__nand2_4
X_62936_ _62646_/B _62936_/X sky130_fd_sc_hd__buf_2
X_81770_ _82896_/CLK _76032_/X _81770_/Q sky130_fd_sc_hd__dfxtp_4
X_69492_ _69580_/A _87769_/Q _69492_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_674_0_CLK clkbuf_9_337_0_CLK/X _87150_/CLK sky130_fd_sc_hd__clkbuf_1
X_49609_ _59167_/B _49606_/X _49608_/Y _49609_/Y sky130_fd_sc_hd__o21ai_4
X_80721_ _80721_/CLK _75907_/X _80721_/Q sky130_fd_sc_hd__dfxtp_4
X_68443_ _68438_/X _68441_/X _68442_/X _68446_/A sky130_fd_sc_hd__a21o_4
X_65655_ _65731_/A _85874_/Q _65655_/X sky130_fd_sc_hd__and2_4
X_50881_ _50879_/Y _50839_/X _50880_/X _86114_/D sky130_fd_sc_hd__a21oi_4
X_62867_ _63586_/A _60337_/D _62866_/Y _62867_/X sky130_fd_sc_hd__o21a_4
X_52620_ _52620_/A _52648_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_165_0_CLK clkbuf_8_82_0_CLK/X clkbuf_9_165_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_64606_ _64561_/X _64582_/Y _64605_/Y _64606_/Y sky130_fd_sc_hd__o21ai_4
X_83440_ _83491_/CLK _83440_/D _83440_/Q sky130_fd_sc_hd__dfxtp_4
X_61818_ _59770_/A _62851_/A sky130_fd_sc_hd__buf_2
X_80652_ _80657_/CLK _80652_/D _46094_/A sky130_fd_sc_hd__dfxtp_4
X_68374_ _68357_/Y _68358_/X _68326_/X _68373_/Y _68374_/X sky130_fd_sc_hd__a211o_4
X_65586_ _65582_/X _65663_/B _65585_/X _65587_/B sky130_fd_sc_hd__nand3_4
Xclkbuf_9_92_0_CLK clkbuf_9_93_0_CLK/A clkbuf_9_92_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_62798_ _57670_/A _62749_/X _62768_/X _62759_/X _62797_/X _62798_/Y
+ sky130_fd_sc_hd__a41oi_4
X_67325_ _87104_/Q _67230_/X _67278_/X _67324_/X _67325_/X sky130_fd_sc_hd__a211o_4
X_52551_ _52567_/A _54069_/B _52551_/Y sky130_fd_sc_hd__nand2_4
X_64537_ _64455_/X _84732_/Q _61102_/X _64537_/Y sky130_fd_sc_hd__nand3_4
X_83371_ _83372_/CLK _83371_/D _83371_/Q sky130_fd_sc_hd__dfxtp_4
X_61749_ _61744_/X _61749_/B _61765_/C _61748_/X _61749_/Y sky130_fd_sc_hd__nand4_4
X_80583_ _80570_/Y _80574_/Y _80582_/X _80584_/B sky130_fd_sc_hd__o21ai_4
XPHY_308 sky130_fd_sc_hd__decap_3
Xclkbuf_10_689_0_CLK clkbuf_9_344_0_CLK/X _87436_/CLK sky130_fd_sc_hd__clkbuf_1
X_85110_ _85114_/CLK _85110_/D _45572_/A sky130_fd_sc_hd__dfxtp_4
XPHY_319 sky130_fd_sc_hd__decap_3
X_51502_ _85998_/Q _51485_/X _51501_/Y _51502_/Y sky130_fd_sc_hd__o21ai_4
X_82322_ _82327_/CLK _77118_/B _82322_/Q sky130_fd_sc_hd__dfxtp_4
X_55270_ _45808_/A _55272_/A _44044_/X _55269_/X _55270_/X sky130_fd_sc_hd__a211o_4
X_67256_ _67252_/X _67254_/X _67255_/X _67256_/Y sky130_fd_sc_hd__a21oi_4
X_86090_ _85770_/CLK _86090_/D _86090_/Q sky130_fd_sc_hd__dfxtp_4
X_52482_ _52468_/A _52482_/B _52482_/Y sky130_fd_sc_hd__nand2_4
X_64468_ _64515_/A _84859_/Q _64515_/C _64468_/Y sky130_fd_sc_hd__nand3_4
X_54221_ _47832_/X _54250_/A sky130_fd_sc_hd__buf_2
X_66207_ _66204_/Y _66205_/X _66206_/X _84149_/D sky130_fd_sc_hd__a21o_4
X_85041_ _85041_/CLK _85041_/D _45647_/A sky130_fd_sc_hd__dfxtp_4
X_51433_ _51410_/X _51421_/X _51438_/C _52963_/D _51433_/X sky130_fd_sc_hd__and4_4
X_63419_ _63368_/X _63410_/X _63411_/X _63415_/X _63418_/Y _63419_/Y
+ sky130_fd_sc_hd__o41ai_4
X_82253_ _82253_/CLK _80418_/X _82253_/Q sky130_fd_sc_hd__dfxtp_4
X_67187_ _84080_/Q _67092_/X _67186_/X _84080_/D sky130_fd_sc_hd__a21bo_4
X_64399_ _58434_/A _64418_/B _64399_/Y sky130_fd_sc_hd__nor2_4
X_81204_ _81211_/CLK _75028_/X _49019_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_612_0_CLK clkbuf_9_306_0_CLK/X _80818_/CLK sky130_fd_sc_hd__clkbuf_1
X_54152_ _54150_/Y _54144_/X _54151_/X _85495_/D sky130_fd_sc_hd__a21oi_4
X_66138_ _66138_/A _66138_/Y sky130_fd_sc_hd__inv_2
X_51364_ _51364_/A _50852_/B _51364_/Y sky130_fd_sc_hd__nand2_4
X_82184_ _85407_/CLK _82184_/D _82184_/Q sky130_fd_sc_hd__dfxtp_4
X_53103_ _53107_/A _53113_/B _53107_/C _53103_/D _53103_/X sky130_fd_sc_hd__and4_4
X_50315_ _50311_/Y _50313_/X _50314_/X _86225_/D sky130_fd_sc_hd__a21oi_4
X_81135_ _83957_/CLK _81135_/D _40689_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_103_0_CLK clkbuf_8_51_0_CLK/X clkbuf_9_103_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_58960_ _58918_/X _58957_/Y _58958_/Y _58959_/X _58923_/X _58960_/X
+ sky130_fd_sc_hd__o32a_4
X_54083_ _53801_/B _52565_/B _54083_/Y sky130_fd_sc_hd__nand2_4
X_66069_ _64593_/A _73827_/B _66069_/X sky130_fd_sc_hd__and2_4
X_51295_ _51293_/Y _51289_/X _51294_/X _51295_/Y sky130_fd_sc_hd__a21oi_4
X_86992_ _82536_/CLK _86992_/D _44705_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_30_0_CLK clkbuf_9_31_0_CLK/A clkbuf_9_30_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_53034_ _85709_/Q _53010_/X _53033_/Y _53034_/Y sky130_fd_sc_hd__o21ai_4
X_57911_ _84941_/Q _57896_/X _57900_/X _57910_/X _84941_/D sky130_fd_sc_hd__a2bb2oi_4
X_50246_ _50537_/A _53190_/A sky130_fd_sc_hd__buf_2
X_85943_ _82768_/CLK _51806_/Y _85943_/Q sky130_fd_sc_hd__dfxtp_4
X_81066_ _81065_/CLK _81098_/Q _75186_/B sky130_fd_sc_hd__dfxtp_4
X_58891_ _59061_/A _58891_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_627_0_CLK clkbuf_9_313_0_CLK/X _81996_/CLK sky130_fd_sc_hd__clkbuf_1
X_80017_ _84931_/Q _84179_/Q _80019_/A sky130_fd_sc_hd__xor2_4
X_57842_ _84946_/Q _57819_/X _57834_/X _57841_/X _84946_/D sky130_fd_sc_hd__a2bb2oi_4
X_69828_ _69825_/X _69827_/X _69742_/X _69828_/Y sky130_fd_sc_hd__a21oi_4
X_50177_ _50169_/A _49135_/X _50177_/Y sky130_fd_sc_hd__nand2_4
X_85874_ _86193_/CLK _85874_/D _85874_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_118_0_CLK clkbuf_8_59_0_CLK/X clkbuf_9_118_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_87613_ _82888_/CLK _87613_/D _67104_/B sky130_fd_sc_hd__dfxtp_4
X_84825_ _84960_/CLK _58537_/X _58535_/A sky130_fd_sc_hd__dfxtp_4
X_57773_ _57947_/A _57773_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_45_0_CLK clkbuf_8_22_0_CLK/X clkbuf_9_45_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_69759_ _69334_/X _69336_/X _69728_/X _69759_/Y sky130_fd_sc_hd__a21oi_4
X_54985_ _54985_/A _47572_/Y _54985_/Y sky130_fd_sc_hd__nand2_4
X_59512_ _59512_/A _59512_/X sky130_fd_sc_hd__buf_2
X_56724_ _56724_/A _56723_/Y _57153_/A sky130_fd_sc_hd__nand2_4
X_87544_ _87544_/CLK _87544_/D _73440_/A sky130_fd_sc_hd__dfxtp_4
X_41950_ _41950_/A _41950_/Y sky130_fd_sc_hd__inv_2
X_53936_ _53871_/X _53936_/B _53936_/Y sky130_fd_sc_hd__nand2_4
X_72770_ _41983_/Y _72723_/X _72725_/X _72769_/Y _72770_/X sky130_fd_sc_hd__a211o_4
X_84756_ _84757_/CLK _84756_/D _84756_/Q sky130_fd_sc_hd__dfxtp_4
X_81968_ _82558_/CLK _81968_/D _81968_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_3_3_0_CLK clkbuf_3_3_0_CLK/A clkbuf_3_3_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_40901_ _46469_/B _40901_/B _40901_/X sky130_fd_sc_hd__or2_4
X_83707_ _83707_/CLK _83707_/D _83707_/Q sky130_fd_sc_hd__dfxtp_4
X_71721_ _70526_/A _71223_/B _70954_/C _71721_/Y sky130_fd_sc_hd__nand3_4
X_59443_ _59443_/A _59445_/A sky130_fd_sc_hd__inv_2
X_56655_ _56655_/A _56655_/Y sky130_fd_sc_hd__inv_2
X_80919_ _84105_/CLK _80919_/D _80919_/Q sky130_fd_sc_hd__dfxtp_4
X_87475_ _87675_/CLK _87475_/D _87475_/Q sky130_fd_sc_hd__dfxtp_4
X_41881_ _41881_/A _42000_/A sky130_fd_sc_hd__buf_2
X_53867_ _50142_/A _53806_/B _53806_/C _53867_/X sky130_fd_sc_hd__and3_4
X_84687_ _84329_/CLK _84687_/D _80347_/A sky130_fd_sc_hd__dfxtp_4
X_81899_ _81975_/CLK _81899_/D _77013_/B sky130_fd_sc_hd__dfxtp_4
X_43620_ _87338_/Q _43620_/Y sky130_fd_sc_hd__inv_2
X_55606_ _44106_/C _55607_/A sky130_fd_sc_hd__buf_2
X_74440_ _74438_/Y _72107_/X _74439_/Y _83066_/D sky130_fd_sc_hd__a21boi_4
X_86426_ _85818_/CLK _49244_/Y _64798_/B sky130_fd_sc_hd__dfxtp_4
X_40832_ _40832_/A _40832_/X sky130_fd_sc_hd__buf_2
X_52818_ _52818_/A _52818_/B _52818_/C _52818_/D _52818_/X sky130_fd_sc_hd__and4_4
X_59374_ _59237_/X _59372_/Y _59373_/Y _59301_/X _59241_/X _59374_/X
+ sky130_fd_sc_hd__o32a_4
X_71652_ _71650_/A _71246_/B _71644_/C _71652_/Y sky130_fd_sc_hd__nand3_4
X_83638_ _86424_/CLK _70996_/Y _83638_/Q sky130_fd_sc_hd__dfxtp_4
X_56586_ _56567_/Y _56764_/B sky130_fd_sc_hd__buf_2
X_53798_ _53798_/A _53838_/A sky130_fd_sc_hd__buf_2
X_70603_ _70714_/A _70613_/B _74533_/D _70594_/X _70603_/Y sky130_fd_sc_hd__nand4_4
X_58325_ _84877_/Q _58326_/A sky130_fd_sc_hd__inv_2
X_43551_ _43550_/Y _43551_/Y sky130_fd_sc_hd__inv_2
X_55537_ _55462_/X _45533_/Y _55537_/Y sky130_fd_sc_hd__nor2_4
X_86357_ _83046_/CLK _49604_/Y _86357_/Q sky130_fd_sc_hd__dfxtp_4
X_74371_ _74371_/A _72113_/B _74366_/C _74371_/X sky130_fd_sc_hd__and3_4
X_40763_ _40758_/X _40759_/X _40762_/X _88340_/Q _40744_/X _40764_/A
+ sky130_fd_sc_hd__o32ai_4
X_52749_ _85761_/Q _52737_/X _52748_/Y _52749_/Y sky130_fd_sc_hd__o21ai_4
X_83569_ _86500_/CLK _71218_/Y _83569_/Q sky130_fd_sc_hd__dfxtp_4
X_71583_ _71626_/A _71583_/B _71582_/X _71583_/Y sky130_fd_sc_hd__nor3_4
X_76110_ _76093_/A _76108_/Y _76109_/Y _76110_/X sky130_fd_sc_hd__a21o_4
X_42502_ _73940_/A _42502_/Y sky130_fd_sc_hd__inv_2
X_85308_ _85213_/CLK _56033_/Y _55943_/B sky130_fd_sc_hd__dfxtp_4
X_73322_ _44305_/X _73577_/B sky130_fd_sc_hd__buf_2
X_46270_ _46270_/A _53951_/B sky130_fd_sc_hd__inv_2
X_70534_ DATA_TO_HASH[7] _70534_/Y sky130_fd_sc_hd__inv_2
X_58256_ _58254_/Y _58268_/B _58256_/Y sky130_fd_sc_hd__nand2_4
X_77090_ _77098_/A _82287_/D _77096_/B sky130_fd_sc_hd__xor2_4
X_43482_ _41693_/X _43465_/X _87400_/Q _43467_/X _43482_/X sky130_fd_sc_hd__a2bb2o_4
X_55468_ _55454_/X _55468_/X sky130_fd_sc_hd__buf_2
X_86288_ _86289_/CLK _86288_/D _86288_/Q sky130_fd_sc_hd__dfxtp_4
X_40694_ _40694_/A _40710_/B _40694_/X sky130_fd_sc_hd__or2_4
X_45221_ _45213_/X _45217_/Y _45220_/Y _45221_/Y sky130_fd_sc_hd__a21oi_4
X_57207_ _56873_/X _57153_/B _57206_/Y _57207_/X sky130_fd_sc_hd__a21o_4
X_76041_ _81339_/Q _76041_/B _76047_/B sky130_fd_sc_hd__xor2_4
X_42433_ _40520_/X _42414_/X _87866_/Q _42415_/X _87866_/D sky130_fd_sc_hd__a2bb2o_4
X_88027_ _87273_/CLK _42115_/X _88027_/Q sky130_fd_sc_hd__dfxtp_4
X_54419_ _54425_/A _52726_/B _54419_/Y sky130_fd_sc_hd__nand2_4
X_73253_ _69823_/B _73250_/X _73251_/X _73252_/Y _73253_/X sky130_fd_sc_hd__a211o_4
X_85239_ _85269_/CLK _56316_/Y _85239_/Q sky130_fd_sc_hd__dfxtp_4
X_70465_ _58342_/Y _70458_/X _70464_/Y _70465_/Y sky130_fd_sc_hd__o21ai_4
X_58187_ _58187_/A _58187_/X sky130_fd_sc_hd__buf_2
X_55399_ _55409_/A _55397_/Y _55398_/Y _55399_/X sky130_fd_sc_hd__a21o_4
X_72204_ _72277_/A _86298_/Q _72204_/Y sky130_fd_sc_hd__nor2_4
X_45152_ _45149_/Y _45151_/Y _45137_/X _45152_/X sky130_fd_sc_hd__a21o_4
X_57138_ _57136_/Y _57137_/X _57087_/X _57138_/Y sky130_fd_sc_hd__a21oi_4
X_42364_ _42350_/X _42346_/X _41757_/X _87899_/Q _42347_/X _42365_/A
+ sky130_fd_sc_hd__o32ai_4
X_73184_ _72988_/X _85585_/Q _73092_/A _73183_/X _73184_/X sky130_fd_sc_hd__a211o_4
X_70396_ _70370_/A _70407_/C sky130_fd_sc_hd__buf_2
X_44103_ _86841_/Q _45938_/A sky130_fd_sc_hd__inv_2
X_79800_ _79782_/X _79785_/Y _79800_/X sky130_fd_sc_hd__or2_4
X_41315_ _41242_/X _41661_/A _41314_/X _41316_/A sky130_fd_sc_hd__o21a_4
X_72135_ _72132_/Y _72134_/Y _59351_/X _72135_/X sky130_fd_sc_hd__a21o_4
X_49960_ _49906_/A _49960_/X sky130_fd_sc_hd__buf_2
X_45083_ _45080_/X _45082_/Y _45049_/X _45083_/Y sky130_fd_sc_hd__a21oi_4
X_57069_ _56850_/X _56976_/X _57069_/Y sky130_fd_sc_hd__nor2_4
X_42295_ _42294_/Y _42295_/Y sky130_fd_sc_hd__inv_2
X_77992_ _77950_/B _77989_/X _77991_/X _77993_/B sky130_fd_sc_hd__a21boi_4
X_48911_ _71972_/B _48912_/B sky130_fd_sc_hd__buf_2
X_44034_ _64850_/A _65614_/A sky130_fd_sc_hd__buf_2
X_79731_ _79721_/X _79722_/X _79730_/Y _79731_/Y sky130_fd_sc_hd__a21boi_4
X_41246_ _41239_/X _41241_/X _41245_/X _68970_/B _41236_/X _41246_/Y
+ sky130_fd_sc_hd__o32ai_4
X_72066_ _72001_/A _72066_/X sky130_fd_sc_hd__buf_2
X_76943_ _76942_/Y _76944_/B sky130_fd_sc_hd__inv_2
X_60080_ _60162_/A _72625_/B sky130_fd_sc_hd__buf_2
X_49891_ _49901_/A _53105_/B _49891_/Y sky130_fd_sc_hd__nand2_4
X_71017_ _71039_/D _71018_/D sky130_fd_sc_hd__buf_2
X_48842_ _48839_/Y _48840_/X _48841_/X _86473_/D sky130_fd_sc_hd__a21oi_4
X_79662_ _79651_/X _79639_/X _79662_/X sky130_fd_sc_hd__and2_4
X_41177_ _41007_/B _41145_/B _41177_/X sky130_fd_sc_hd__or2_4
X_76874_ _76874_/A _76874_/B _76874_/Y sky130_fd_sc_hd__xnor2_4
X_78613_ _78613_/A _78616_/B sky130_fd_sc_hd__inv_2
X_75825_ _75824_/A _75824_/B _81021_/Q _75825_/X sky130_fd_sc_hd__a21o_4
X_48773_ _48777_/A _52158_/B _48773_/Y sky130_fd_sc_hd__nand2_4
X_79593_ _79591_/Y _79594_/A sky130_fd_sc_hd__inv_2
X_45985_ _45980_/X _44865_/X _40431_/X _86827_/Q _45982_/X _45985_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47724_ _47719_/Y _47698_/X _47723_/X _86605_/D sky130_fd_sc_hd__a21oi_4
X_78544_ _78561_/B _78561_/A _82770_/D sky130_fd_sc_hd__xor2_4
X_44936_ _85311_/Q _44935_/X _45757_/A _44936_/X sky130_fd_sc_hd__o21a_4
X_75756_ _75742_/Y _75743_/Y _75732_/A _80788_/D _75756_/X sky130_fd_sc_hd__a2bb2o_4
X_63770_ _63766_/X _63744_/X _63769_/Y _84296_/D sky130_fd_sc_hd__a21oi_4
X_60982_ _60982_/A _64032_/A sky130_fd_sc_hd__buf_2
X_72968_ _72969_/B _72969_/C _72967_/X _72968_/X sky130_fd_sc_hd__a21o_4
X_62721_ _62893_/A _62721_/X sky130_fd_sc_hd__buf_2
X_74707_ MACRO_RD_SELECT _74711_/A sky130_fd_sc_hd__buf_2
X_47655_ _47655_/A _47692_/B _47614_/X _53170_/D _47655_/X sky130_fd_sc_hd__and4_4
X_71919_ _56672_/Y _71917_/X _71918_/Y _83329_/D sky130_fd_sc_hd__o21ai_4
X_78475_ _78475_/A _78475_/B _78476_/A sky130_fd_sc_hd__nor2_4
X_44867_ _44867_/A _86912_/D sky130_fd_sc_hd__inv_2
X_75687_ _75687_/A _75689_/A sky130_fd_sc_hd__inv_2
X_72899_ _72899_/A _72899_/X sky130_fd_sc_hd__buf_2
X_46606_ _83689_/Q _52577_/B sky130_fd_sc_hd__inv_2
X_65440_ _65438_/X _86208_/Q _65182_/X _65439_/X _65440_/X sky130_fd_sc_hd__a211o_4
X_77426_ _77422_/Y _77423_/Y _77426_/C _77426_/X sky130_fd_sc_hd__or3_4
X_43818_ _43802_/A _43818_/X sky130_fd_sc_hd__buf_2
X_62652_ _62395_/X _62652_/X sky130_fd_sc_hd__buf_2
X_74638_ _45951_/Y _74638_/X sky130_fd_sc_hd__buf_2
X_47586_ _47586_/A _53133_/D sky130_fd_sc_hd__buf_2
X_44798_ _41428_/Y _44788_/X _86949_/Q _44789_/X _86949_/D sky130_fd_sc_hd__a2bb2o_4
X_61603_ _61413_/A _61634_/A sky130_fd_sc_hd__buf_2
X_49325_ _86409_/Q _49285_/X _49324_/Y _49325_/Y sky130_fd_sc_hd__o21ai_4
X_46537_ _82920_/Q _46527_/X _46537_/X sky130_fd_sc_hd__or2_4
X_65371_ _65045_/A _65397_/B sky130_fd_sc_hd__buf_2
X_77357_ _77339_/B _77339_/A _77356_/Y _77359_/A sky130_fd_sc_hd__a21boi_4
X_43749_ _40929_/X _43736_/X _69967_/B _43737_/X _87284_/D sky130_fd_sc_hd__a2bb2o_4
X_62583_ _62551_/X _62553_/X _84399_/Q _62583_/Y sky130_fd_sc_hd__nor3_4
X_74569_ _74552_/X _74569_/X sky130_fd_sc_hd__buf_2
X_67110_ _66868_/A _67110_/X sky130_fd_sc_hd__buf_2
X_64322_ _64263_/A _64336_/A sky130_fd_sc_hd__buf_2
X_76308_ _76299_/Y _76321_/A _76311_/A sky130_fd_sc_hd__xor2_4
X_49256_ _48535_/A _49261_/A sky130_fd_sc_hd__buf_2
X_61534_ _61413_/A _61546_/A sky130_fd_sc_hd__buf_2
X_68090_ _66580_/X _66584_/X _67897_/X _68090_/Y sky130_fd_sc_hd__a21oi_4
X_46468_ _82926_/Q _48034_/B sky130_fd_sc_hd__inv_2
X_77288_ _77274_/B _77288_/Y sky130_fd_sc_hd__inv_2
X_48207_ _47895_/B _48207_/X sky130_fd_sc_hd__buf_2
X_67041_ _66942_/A _67041_/B _67041_/X sky130_fd_sc_hd__and2_4
X_79027_ _79027_/A _79027_/B _79028_/B sky130_fd_sc_hd__xor2_4
X_45419_ _63017_/B _61338_/A sky130_fd_sc_hd__buf_2
X_64253_ _64242_/Y _64252_/X _72577_/B _64253_/X sky130_fd_sc_hd__o21a_4
X_76239_ _76238_/X _76239_/X sky130_fd_sc_hd__buf_2
X_49187_ _65392_/B _49153_/X _49186_/Y _49187_/Y sky130_fd_sc_hd__o21ai_4
X_61465_ _61308_/A _72528_/A sky130_fd_sc_hd__buf_2
X_46399_ _46399_/A _46399_/X sky130_fd_sc_hd__buf_2
X_63204_ _60606_/X _63204_/X sky130_fd_sc_hd__buf_2
X_48138_ _48138_/A _48342_/A _48138_/X sky130_fd_sc_hd__and2_4
X_60416_ _60447_/B _60417_/A sky130_fd_sc_hd__buf_2
X_64184_ _64184_/A _58370_/A _64184_/C _64184_/X sky130_fd_sc_hd__and3_4
X_61396_ _61393_/X _61394_/X _61395_/Y _84484_/D sky130_fd_sc_hd__a21oi_4
X_63135_ _63088_/A _84830_/Q _63087_/X _63135_/D _63135_/X sky130_fd_sc_hd__and4_4
X_48069_ _52050_/A _48069_/B _48723_/C _48069_/X sky130_fd_sc_hd__and3_4
X_60347_ _60069_/Y _60343_/Y _60337_/D _60344_/Y _60346_/Y _60347_/Y
+ sky130_fd_sc_hd__a41oi_4
X_68992_ _68988_/X _68991_/X _68922_/X _68992_/X sky130_fd_sc_hd__a21o_4
X_50100_ _86264_/Q _50088_/X _50099_/Y _50100_/Y sky130_fd_sc_hd__o21ai_4
X_51080_ _51097_/A _52773_/B _51080_/Y sky130_fd_sc_hd__nand2_4
X_67943_ _67992_/A _88218_/Q _67943_/X sky130_fd_sc_hd__and2_4
X_79929_ _79928_/Y _79929_/Y sky130_fd_sc_hd__inv_2
X_63066_ _63041_/A _63066_/B _63030_/C _63066_/D _63066_/X sky130_fd_sc_hd__and4_4
X_60278_ _60244_/A _60244_/B _79806_/A _60278_/Y sky130_fd_sc_hd__nor3_4
X_50031_ _50050_/A _50040_/B _50025_/C _53244_/D _50031_/X sky130_fd_sc_hd__and4_4
X_62017_ _62002_/A _62002_/B _78062_/B _62017_/Y sky130_fd_sc_hd__nor3_4
X_82940_ _81198_/CLK _78086_/X _82940_/Q sky130_fd_sc_hd__dfxtp_4
X_67874_ _87145_/Q _67825_/X _67872_/X _67873_/X _67874_/X sky130_fd_sc_hd__a211o_4
X_69613_ _87068_/Q _69485_/X _69611_/X _69612_/X _69613_/X sky130_fd_sc_hd__a211o_4
X_66825_ _66821_/X _66824_/X _66658_/X _66825_/Y sky130_fd_sc_hd__a21oi_4
X_82871_ _82498_/CLK _82495_/Q _82871_/Q sky130_fd_sc_hd__dfxtp_4
X_84610_ _83216_/CLK _60498_/Y _79150_/A sky130_fd_sc_hd__dfxtp_4
X_81822_ _81275_/CLK _81630_/Q _81822_/Q sky130_fd_sc_hd__dfxtp_4
X_69544_ _69626_/A _69544_/B _69544_/X sky130_fd_sc_hd__and2_4
X_54770_ _54775_/A _54788_/B _54775_/C _47494_/A _54770_/X sky130_fd_sc_hd__and4_4
X_66756_ _84098_/Q _66734_/X _66755_/X _84098_/D sky130_fd_sc_hd__a21bo_4
X_85590_ _85590_/CLK _53677_/Y _85590_/Q sky130_fd_sc_hd__dfxtp_4
X_51982_ _52407_/A _51982_/X sky130_fd_sc_hd__buf_2
X_63968_ _60967_/A _61502_/A _63962_/X _63965_/Y _63967_/Y _63968_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_53721_ _53719_/Y _53715_/X _53720_/X _53721_/Y sky130_fd_sc_hd__a21oi_4
X_65707_ _65407_/A _65707_/X sky130_fd_sc_hd__buf_2
X_84541_ _84534_/CLK _84541_/D _76989_/A sky130_fd_sc_hd__dfxtp_4
X_50933_ _86104_/Q _50910_/X _50932_/Y _50933_/Y sky130_fd_sc_hd__o21ai_4
X_62919_ _84842_/Q _62642_/B _62919_/Y sky130_fd_sc_hd__nor2_4
X_81753_ _81756_/CLK _76090_/B _41326_/A sky130_fd_sc_hd__dfxtp_4
X_69475_ _68969_/X _68971_/X _69418_/X _69475_/Y sky130_fd_sc_hd__a21oi_4
X_66687_ _84101_/Q _66614_/X _66686_/X _66687_/X sky130_fd_sc_hd__a21bo_4
X_63899_ _61451_/A _63853_/B _63947_/C _63866_/X _63899_/Y sky130_fd_sc_hd__nand4_4
X_56440_ _56446_/A _56446_/B _85193_/Q _56440_/Y sky130_fd_sc_hd__nand3_4
X_68426_ _88017_/Q _68402_/X _68359_/X _68425_/X _68426_/X sky130_fd_sc_hd__a211o_4
X_80704_ _81104_/CLK _80704_/D _80704_/Q sky130_fd_sc_hd__dfxtp_4
X_87260_ _87260_/CLK _87260_/D _87260_/Q sky130_fd_sc_hd__dfxtp_4
X_65638_ _65118_/A _65638_/X sky130_fd_sc_hd__buf_2
X_53652_ _85594_/Q _53626_/X _53651_/Y _53652_/Y sky130_fd_sc_hd__o21ai_4
X_84472_ _82452_/CLK _61547_/Y _61546_/C sky130_fd_sc_hd__dfxtp_4
X_50864_ _50845_/A _54075_/B _50864_/Y sky130_fd_sc_hd__nand2_4
X_81684_ _81684_/CLK _81684_/D _81684_/Q sky130_fd_sc_hd__dfxtp_4
X_86211_ _86203_/CLK _86211_/D _86211_/Q sky130_fd_sc_hd__dfxtp_4
X_52603_ _52624_/A _46662_/A _52603_/Y sky130_fd_sc_hd__nand2_4
X_83423_ _84945_/CLK _71657_/Y _58508_/A sky130_fd_sc_hd__dfxtp_4
X_56371_ _56370_/Y _56439_/A sky130_fd_sc_hd__buf_2
X_80635_ _80270_/X _80271_/Y _80635_/Y sky130_fd_sc_hd__nand2_4
X_68357_ _68352_/X _68356_/X _68357_/Y sky130_fd_sc_hd__nand2_4
X_87191_ _87189_/CLK _87191_/D _68000_/B sky130_fd_sc_hd__dfxtp_4
X_53583_ _50360_/A _53620_/B _53620_/C _53583_/X sky130_fd_sc_hd__and3_4
X_65569_ _65416_/X _73016_/B _65569_/X sky130_fd_sc_hd__and2_4
X_50795_ _50777_/A _46412_/B _50795_/Y sky130_fd_sc_hd__nand2_4
X_58110_ _57997_/X _85476_/Q _58109_/X _58110_/X sky130_fd_sc_hd__o21a_4
XPHY_105 sky130_fd_sc_hd__decap_3
X_55322_ _55318_/X _55321_/X _55309_/X _55322_/X sky130_fd_sc_hd__a21o_4
X_67308_ _67308_/A _86807_/Q _67308_/X sky130_fd_sc_hd__and2_4
X_86142_ _85535_/CLK _86142_/D _86142_/Q sky130_fd_sc_hd__dfxtp_4
X_52534_ _52531_/Y _52532_/X _52533_/X _85803_/D sky130_fd_sc_hd__a21oi_4
XPHY_116 sky130_fd_sc_hd__decap_3
X_59090_ _59090_/A _59090_/B _59090_/Y sky130_fd_sc_hd__nor2_4
X_83354_ _83761_/CLK _71844_/X _83354_/Q sky130_fd_sc_hd__dfxtp_4
X_80566_ _80560_/A _80560_/B _80565_/Y _80566_/Y sky130_fd_sc_hd__a21boi_4
X_68288_ _67775_/X _67778_/X _68260_/X _68288_/Y sky130_fd_sc_hd__a21oi_4
XPHY_127 sky130_fd_sc_hd__decap_3
XPHY_138 sky130_fd_sc_hd__decap_3
XPHY_149 sky130_fd_sc_hd__decap_3
X_58041_ _58030_/X _85482_/Q _57962_/X _58041_/X sky130_fd_sc_hd__o21a_4
X_82305_ _82557_/CLK _82305_/D _82305_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_551_0_CLK clkbuf_9_275_0_CLK/X _81783_/CLK sky130_fd_sc_hd__clkbuf_1
X_55253_ _82984_/Q _44059_/A _55140_/X _55252_/X _55253_/X sky130_fd_sc_hd__a211o_4
X_67239_ _67120_/X _67239_/X sky130_fd_sc_hd__buf_2
X_86073_ _85754_/CLK _51106_/Y _86073_/Q sky130_fd_sc_hd__dfxtp_4
X_52465_ _52461_/Y _52462_/X _52464_/Y _52465_/Y sky130_fd_sc_hd__a21boi_4
Xclkbuf_6_42_0_CLK clkbuf_6_43_0_CLK/A clkbuf_7_85_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_83285_ _86149_/CLK _83285_/D _83285_/Q sky130_fd_sc_hd__dfxtp_4
X_80497_ _80497_/A _63517_/C _80498_/B sky130_fd_sc_hd__xor2_4
X_54204_ _54202_/Y _54197_/X _54203_/X _85485_/D sky130_fd_sc_hd__a21oi_4
X_85024_ _83008_/CLK _85024_/D _85024_/Q sky130_fd_sc_hd__dfxtp_4
X_51416_ _51410_/X _51230_/X _51438_/C _52942_/D _51416_/X sky130_fd_sc_hd__and4_4
X_70250_ _70249_/X _70260_/D sky130_fd_sc_hd__buf_2
X_82236_ _82515_/CLK _82268_/Q _82236_/Q sky130_fd_sc_hd__dfxtp_4
X_55184_ _55711_/A _57430_/A _55184_/X sky130_fd_sc_hd__and2_4
X_52396_ _52394_/Y _52390_/X _52395_/X _52396_/Y sky130_fd_sc_hd__a21oi_4
X_54135_ _85497_/Q _54113_/X _54134_/Y _54135_/Y sky130_fd_sc_hd__o21ai_4
X_51347_ _51265_/A _51352_/B sky130_fd_sc_hd__buf_2
X_70181_ _70181_/A _70160_/X _70162_/X _70164_/X _70181_/Y sky130_fd_sc_hd__nand4_4
X_82167_ _82009_/CLK _84159_/Q _82167_/Q sky130_fd_sc_hd__dfxtp_4
X_59992_ _59873_/A _59873_/B _59992_/C _59992_/Y sky130_fd_sc_hd__nor3_4
X_41100_ _40931_/A _41100_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_566_0_CLK clkbuf_9_283_0_CLK/X _87348_/CLK sky130_fd_sc_hd__clkbuf_1
X_81118_ _81048_/CLK _79859_/X _81118_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_6_57_0_CLK clkbuf_6_57_0_CLK/A clkbuf_6_57_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_42080_ _42080_/A _88044_/D sky130_fd_sc_hd__inv_2
X_58943_ _58766_/A _58943_/X sky130_fd_sc_hd__buf_2
X_54066_ _54064_/Y _54060_/X _54065_/Y _85512_/D sky130_fd_sc_hd__a21boi_4
X_51278_ _51278_/A _51278_/B _51278_/X sky130_fd_sc_hd__and2_4
X_86975_ _87416_/CLK _86975_/D _86975_/Q sky130_fd_sc_hd__dfxtp_4
X_82098_ _82860_/CLK _77468_/B _77118_/A sky130_fd_sc_hd__dfxtp_4
X_41031_ _41024_/X _81712_/Q _41030_/X _41032_/A sky130_fd_sc_hd__o21ai_4
X_53017_ _53025_/A _53017_/B _53017_/Y sky130_fd_sc_hd__nand2_4
X_50229_ _50228_/X _50230_/A sky130_fd_sc_hd__buf_2
X_73940_ _73940_/A _74244_/B _73940_/Y sky130_fd_sc_hd__nor2_4
X_85926_ _85447_/CLK _51899_/Y _85926_/Q sky130_fd_sc_hd__dfxtp_4
X_81049_ _84269_/CLK _75421_/X _81049_/Q sky130_fd_sc_hd__dfxtp_4
X_58874_ _58603_/A _58874_/X sky130_fd_sc_hd__buf_2
Xclkbuf_1_0_2_CLK clkbuf_1_0_2_CLK/A clkbuf_2_1_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_57825_ _57824_/X _85499_/Q _57736_/X _57825_/X sky130_fd_sc_hd__o21a_4
X_85857_ _83311_/CLK _52264_/Y _85857_/Q sky130_fd_sc_hd__dfxtp_4
X_73871_ _68693_/B _73674_/X _73819_/X _73870_/Y _73871_/X sky130_fd_sc_hd__a211o_4
X_75610_ _75640_/A _75609_/Y _75611_/B sky130_fd_sc_hd__xor2_4
X_84808_ _84807_/CLK _84808_/D _84808_/Q sky130_fd_sc_hd__dfxtp_4
X_72822_ _72820_/X _72802_/X _72822_/C _72822_/Y sky130_fd_sc_hd__nand3_4
X_45770_ _45768_/Y _45734_/X _45720_/X _45769_/Y _45770_/X sky130_fd_sc_hd__a211o_4
X_57756_ _59801_/A _57757_/A sky130_fd_sc_hd__buf_2
X_76590_ _76516_/Y _76584_/X _76589_/Y _76616_/B sky130_fd_sc_hd__a21oi_4
X_42982_ _42981_/Y _87620_/D sky130_fd_sc_hd__inv_2
X_54968_ _54250_/A _54985_/A sky130_fd_sc_hd__buf_2
X_85788_ _85786_/CLK _85788_/D _85788_/Q sky130_fd_sc_hd__dfxtp_4
X_44721_ _44712_/X _44713_/X _40702_/X _86987_/Q _44714_/X _44721_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56707_ _46234_/Y _56707_/X sky130_fd_sc_hd__buf_2
X_75541_ _75541_/A _75543_/A sky130_fd_sc_hd__inv_2
X_87527_ _87782_/CLK _43231_/Y _87527_/Q sky130_fd_sc_hd__dfxtp_4
X_41933_ _41932_/X _41927_/X _40667_/X _73892_/A _41928_/X _41934_/A
+ sky130_fd_sc_hd__o32ai_4
X_53919_ _53902_/A _53919_/B _53919_/Y sky130_fd_sc_hd__nand2_4
X_72753_ _72750_/X _85601_/Q _44130_/X _72752_/X _72753_/X sky130_fd_sc_hd__a211o_4
X_84739_ _83451_/CLK _84739_/D _84739_/Q sky130_fd_sc_hd__dfxtp_4
X_57687_ _57687_/A _59629_/A sky130_fd_sc_hd__inv_2
X_54899_ _85357_/Q _54892_/X _54898_/Y _54899_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_504_0_CLK clkbuf_9_252_0_CLK/X _86393_/CLK sky130_fd_sc_hd__clkbuf_1
X_47440_ _47437_/X _47415_/X _47466_/C _53048_/D _47440_/X sky130_fd_sc_hd__and4_4
X_71704_ _71338_/A _71685_/X _71333_/C _71704_/Y sky130_fd_sc_hd__nand3_4
X_59426_ _74831_/A _59426_/X sky130_fd_sc_hd__buf_2
X_78260_ _78263_/A _78259_/Y _78261_/B sky130_fd_sc_hd__xor2_4
X_44652_ _41064_/A _44648_/X _87016_/Q _44650_/X _44652_/X sky130_fd_sc_hd__a2bb2o_4
X_56638_ _55467_/X _56638_/B _56638_/X sky130_fd_sc_hd__xor2_4
X_87458_ _87720_/CLK _87458_/D _87458_/Q sky130_fd_sc_hd__dfxtp_4
X_75472_ _75472_/A _81052_/D _75472_/X sky130_fd_sc_hd__xor2_4
X_41864_ _42626_/A _41902_/A sky130_fd_sc_hd__buf_2
X_72684_ _83190_/Q _72672_/X _72683_/Y _72684_/X sky130_fd_sc_hd__a21bo_4
X_77211_ _77200_/A _82302_/D _77211_/Y sky130_fd_sc_hd__nand2_4
X_43603_ _43602_/X _55102_/A sky130_fd_sc_hd__buf_2
X_74423_ _74413_/X _53678_/B _74423_/Y sky130_fd_sc_hd__nand2_4
X_86409_ _85800_/CLK _49329_/Y _86409_/Q sky130_fd_sc_hd__dfxtp_4
X_40815_ _40758_/X _40759_/X _40814_/X _88329_/Q _40744_/X _40816_/A
+ sky130_fd_sc_hd__o32ai_4
X_47371_ _47362_/Y _47364_/X _47370_/X _86642_/D sky130_fd_sc_hd__a21oi_4
X_59357_ _59219_/X _85732_/Q _59220_/X _59357_/X sky130_fd_sc_hd__o21a_4
X_71635_ _71637_/A _71223_/B _71637_/C _71635_/Y sky130_fd_sc_hd__nand3_4
X_78191_ _78191_/A _78191_/B _78191_/C _78191_/X sky130_fd_sc_hd__and3_4
X_44583_ _44583_/A _44583_/Y sky130_fd_sc_hd__inv_2
X_56569_ _56558_/X _72641_/C _56564_/B _56569_/X sky130_fd_sc_hd__and3_4
X_87389_ _87195_/CLK _87389_/D _87389_/Q sky130_fd_sc_hd__dfxtp_4
X_41795_ _40620_/X _81185_/Q _41795_/X sky130_fd_sc_hd__or2_4
XPHY_7 sky130_fd_sc_hd__decap_3
X_49110_ _49110_/A _46348_/A _49110_/Y sky130_fd_sc_hd__nand2_4
X_46322_ _50755_/A _46428_/B _46428_/C _46322_/X sky130_fd_sc_hd__and3_4
X_58308_ _63348_/A _58280_/B _58308_/Y sky130_fd_sc_hd__nand2_4
X_77142_ _77142_/A _77142_/B _77142_/Y sky130_fd_sc_hd__nand2_4
X_43534_ _40400_/X _43532_/X _87373_/Q _43533_/X _87373_/D sky130_fd_sc_hd__a2bb2o_4
X_74354_ _83086_/Q _73050_/A _74353_/Y _83086_/D sky130_fd_sc_hd__a21o_4
X_40746_ _40746_/A _88343_/D sky130_fd_sc_hd__inv_2
X_71566_ _71557_/X _83454_/Q _71565_/Y _71566_/X sky130_fd_sc_hd__a21o_4
X_59288_ _59286_/X _86058_/Q _59287_/X _59288_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_519_0_CLK clkbuf_9_259_0_CLK/X _81322_/CLK sky130_fd_sc_hd__clkbuf_1
X_49041_ _49041_/A _53858_/B sky130_fd_sc_hd__buf_2
X_73305_ _73257_/X _86188_/Q _73205_/X _73304_/X _73305_/X sky130_fd_sc_hd__a211o_4
X_46253_ _46280_/A _46272_/A sky130_fd_sc_hd__buf_2
X_70517_ _57663_/Y _70501_/X _70516_/Y _83758_/D sky130_fd_sc_hd__o21ai_4
XPHY_650 sky130_fd_sc_hd__decap_3
X_58239_ _58219_/X _58236_/Y _58238_/Y _58239_/Y sky130_fd_sc_hd__a21oi_4
X_77073_ _77073_/A _77084_/A _77074_/B sky130_fd_sc_hd__xor2_4
X_43465_ _43513_/A _43465_/X sky130_fd_sc_hd__buf_2
X_74285_ _70267_/C _72702_/X _74284_/Y _74285_/X sky130_fd_sc_hd__a21bo_4
XPHY_661 sky130_fd_sc_hd__decap_3
X_40677_ _40670_/X _82865_/Q _40676_/X _40678_/A sky130_fd_sc_hd__o21ai_4
X_71497_ _71487_/X _83478_/Q _71496_/X _71497_/X sky130_fd_sc_hd__a21o_4
XPHY_672 sky130_fd_sc_hd__decap_3
XPHY_683 sky130_fd_sc_hd__decap_3
X_45204_ _45202_/X _61558_/B _45144_/X _45204_/Y sky130_fd_sc_hd__o21ai_4
X_76024_ _76024_/A _76023_/Y _81744_/D sky130_fd_sc_hd__xor2_4
X_42416_ _40469_/X _42414_/X _87875_/Q _42415_/X _42416_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_694 sky130_fd_sc_hd__decap_3
X_61250_ _61262_/A _61250_/B _61250_/C _61250_/Y sky130_fd_sc_hd__nor3_4
X_73236_ _73210_/X _85583_/Q _73092_/X _73235_/X _73236_/X sky130_fd_sc_hd__a211o_4
X_46184_ _46195_/A _46128_/A _46133_/B _46184_/Y sky130_fd_sc_hd__nand3_4
X_70448_ _71650_/A _70954_/B _71194_/C _70448_/Y sky130_fd_sc_hd__nand3_4
X_43396_ _43396_/A _43396_/X sky130_fd_sc_hd__buf_2
X_60201_ _60227_/A _60202_/A sky130_fd_sc_hd__buf_2
X_45135_ _55848_/B _45134_/X _45116_/X _45135_/X sky130_fd_sc_hd__o21a_4
X_42347_ _41872_/A _42347_/X sky130_fd_sc_hd__buf_2
X_73167_ _73163_/X _83066_/Q _72880_/X _73166_/X _73167_/X sky130_fd_sc_hd__a211o_4
X_61181_ _64263_/A _64250_/A sky130_fd_sc_hd__buf_2
X_70379_ _70366_/X _74523_/A _70375_/C _70379_/Y sky130_fd_sc_hd__nand3_4
X_60132_ _60132_/A _60132_/X sky130_fd_sc_hd__buf_2
X_72118_ _86625_/Q _72193_/B _72118_/Y sky130_fd_sc_hd__nor2_4
X_49943_ _49925_/X _49943_/B _49953_/C _53155_/D _49943_/X sky130_fd_sc_hd__and4_4
X_45066_ _83031_/Q _45067_/A sky130_fd_sc_hd__inv_2
X_42278_ _42277_/Y _87944_/D sky130_fd_sc_hd__inv_2
X_73098_ _73098_/A _73097_/X _73098_/Y sky130_fd_sc_hd__nand2_4
X_77975_ _77975_/A _78043_/A _77975_/Y sky130_fd_sc_hd__nor2_4
X_44017_ _57848_/A _57736_/A sky130_fd_sc_hd__buf_2
X_79714_ _79712_/X _79719_/B _79714_/Y sky130_fd_sc_hd__xnor2_4
X_41229_ _41184_/X _40710_/A _41228_/X _41230_/A sky130_fd_sc_hd__o21ai_4
X_64940_ _64739_/A _65047_/A sky130_fd_sc_hd__buf_2
X_60063_ _60062_/X _60063_/Y sky130_fd_sc_hd__inv_2
X_72049_ _49069_/A _72043_/X _72048_/X _72049_/X sky130_fd_sc_hd__and3_4
X_76926_ _81471_/D _76926_/B _76928_/A sky130_fd_sc_hd__nand2_4
X_49874_ _49864_/A _53086_/B _49874_/Y sky130_fd_sc_hd__nand2_4
X_48825_ _48831_/A _50508_/B _48825_/Y sky130_fd_sc_hd__nand2_4
X_79645_ _79639_/X _79645_/B _79645_/X sky130_fd_sc_hd__xor2_4
X_64871_ _64868_/Y _64814_/X _64870_/Y _64871_/X sky130_fd_sc_hd__a21o_4
X_76857_ _81673_/Q _76857_/B _76857_/Y sky130_fd_sc_hd__xnor2_4
X_66610_ _88402_/Q _66608_/X _46212_/A _66609_/X _66610_/X sky130_fd_sc_hd__a211o_4
X_63822_ _58237_/X _63858_/B _63858_/C _63793_/D _63822_/Y sky130_fd_sc_hd__nand4_4
X_75808_ _75832_/B _75810_/B sky130_fd_sc_hd__inv_2
X_48756_ _48837_/A _48777_/A sky130_fd_sc_hd__buf_2
X_67590_ _84063_/Q _67568_/X _67589_/X _67590_/X sky130_fd_sc_hd__a21bo_4
X_79576_ _79576_/A _79576_/B _79577_/A sky130_fd_sc_hd__nand2_4
X_45968_ _45967_/Y _86836_/D sky130_fd_sc_hd__inv_2
X_76788_ _76781_/Y _76774_/X _76787_/Y _76788_/Y sky130_fd_sc_hd__a21oi_4
X_47707_ _86606_/Q _47666_/X _47706_/Y _47707_/Y sky130_fd_sc_hd__o21ai_4
X_66541_ _44019_/A _67816_/A sky130_fd_sc_hd__buf_2
X_78527_ _78526_/B _78526_/C _78522_/Y _78528_/B sky130_fd_sc_hd__o21ai_4
X_44919_ _45153_/A _44919_/X sky130_fd_sc_hd__buf_2
X_63753_ _63369_/B _64177_/B _63753_/C _64177_/D _63759_/B sky130_fd_sc_hd__nand4_4
X_75739_ _75723_/B _75736_/X _75738_/Y _75740_/B sky130_fd_sc_hd__a21oi_4
X_48687_ _48687_/A _48632_/B _48687_/Y sky130_fd_sc_hd__nand2_4
X_60965_ _60930_/A _60855_/X _60930_/C _60966_/A sky130_fd_sc_hd__nand3_4
X_45899_ _44039_/X _46159_/A sky130_fd_sc_hd__buf_2
X_62704_ _62669_/A _63054_/A _62704_/C _62669_/D _62704_/X sky130_fd_sc_hd__and4_4
X_69260_ _88042_/Q _69217_/X _69245_/X _69259_/X _69260_/X sky130_fd_sc_hd__a211o_4
X_47638_ _47634_/Y _47602_/X _47637_/X _86614_/D sky130_fd_sc_hd__a21oi_4
X_66472_ _60110_/X _65154_/Y _66471_/Y _66472_/Y sky130_fd_sc_hd__o21ai_4
X_78458_ _78458_/A _82669_/D _78458_/Y sky130_fd_sc_hd__nor2_4
X_63684_ _63696_/A _62151_/X _63684_/X sky130_fd_sc_hd__and2_4
X_60896_ _60895_/X _60896_/Y sky130_fd_sc_hd__inv_2
X_68211_ _68196_/X _67292_/Y _68207_/X _68210_/Y _68211_/X sky130_fd_sc_hd__a211o_4
X_65423_ _65401_/A _65423_/B _65423_/X sky130_fd_sc_hd__and2_4
X_77409_ _77409_/A _82095_/D _77412_/B sky130_fd_sc_hd__nor2_4
X_62635_ _62628_/X _62630_/X _62634_/Y _58374_/A _62212_/A _62635_/Y
+ sky130_fd_sc_hd__o32ai_4
X_69191_ _69191_/A _87791_/Q _69191_/X sky130_fd_sc_hd__and2_4
X_47569_ _47564_/Y _47555_/X _47568_/X _47569_/Y sky130_fd_sc_hd__a21oi_4
X_78389_ _78384_/Y _78390_/A sky130_fd_sc_hd__inv_2
X_49308_ _52524_/A _49283_/B _49234_/X _49308_/X sky130_fd_sc_hd__and3_4
X_80420_ _80412_/X _80413_/X _80419_/Y _80436_/A sky130_fd_sc_hd__a21boi_4
X_68142_ _68121_/X _66886_/Y _68128_/X _68141_/Y _68142_/X sky130_fd_sc_hd__a211o_4
X_65354_ _65403_/A _86244_/Q _65354_/X sky130_fd_sc_hd__and2_4
X_50580_ _50580_/A _71974_/B _50580_/Y sky130_fd_sc_hd__nand2_4
X_62566_ _61630_/A _62566_/B _62501_/X _62566_/D _62569_/B sky130_fd_sc_hd__nand4_4
X_64305_ _64275_/A _64305_/B _64274_/X _64305_/X sky130_fd_sc_hd__and3_4
X_49239_ _49220_/A _52454_/B _49239_/Y sky130_fd_sc_hd__nand2_4
X_61517_ _61394_/A _61517_/X sky130_fd_sc_hd__buf_2
X_80351_ _80350_/B _80350_/C _80352_/A sky130_fd_sc_hd__nand2_4
X_68073_ _68068_/X _68072_/X _67977_/X _68077_/A sky130_fd_sc_hd__a21o_4
X_65285_ _65285_/A _65285_/B _65285_/X sky130_fd_sc_hd__and2_4
X_62497_ _62488_/X _62493_/Y _62496_/X _84846_/Q _62440_/X _62497_/Y
+ sky130_fd_sc_hd__o32ai_4
X_67024_ _87360_/Q _66997_/X _66998_/X _67023_/X _67024_/X sky130_fd_sc_hd__a211o_4
X_52250_ _52250_/A _48695_/B _52250_/Y sky130_fd_sc_hd__nand2_4
X_64236_ _64248_/A _64225_/B _64236_/C _64236_/X sky130_fd_sc_hd__and3_4
X_83070_ _86516_/CLK _74422_/Y _83070_/Q sky130_fd_sc_hd__dfxtp_4
X_61448_ _58543_/A _61448_/X sky130_fd_sc_hd__buf_2
X_80282_ _80274_/Y _80282_/Y sky130_fd_sc_hd__inv_2
X_51201_ _51147_/A _51201_/X sky130_fd_sc_hd__buf_2
X_82021_ _81954_/CLK _77761_/B _81989_/D sky130_fd_sc_hd__dfxtp_4
X_52181_ _85873_/Q _52178_/X _52180_/Y _52181_/Y sky130_fd_sc_hd__o21ai_4
X_64167_ _63694_/B _64190_/B _64178_/C _64190_/D _64167_/Y sky130_fd_sc_hd__nand4_4
X_61379_ _61313_/A _61380_/A sky130_fd_sc_hd__buf_2
X_51132_ _51115_/A _51121_/B _51115_/C _52827_/D _51132_/X sky130_fd_sc_hd__and4_4
X_63118_ _63118_/A _63118_/X sky130_fd_sc_hd__buf_2
X_64098_ _64162_/A _58461_/A _64173_/C _64098_/X sky130_fd_sc_hd__and3_4
X_68975_ _69958_/A _68975_/X sky130_fd_sc_hd__buf_2
X_55940_ _55949_/A _85180_/Q _55940_/X sky130_fd_sc_hd__and2_4
X_51063_ _51058_/A _52752_/B _51063_/Y sky130_fd_sc_hd__nand2_4
X_67926_ _68637_/A _67972_/A sky130_fd_sc_hd__buf_2
X_63049_ _63038_/A _63049_/B _63085_/C _60541_/B _63049_/X sky130_fd_sc_hd__and4_4
X_86760_ _81990_/CLK _46216_/Y _44012_/A sky130_fd_sc_hd__dfxtp_4
X_83972_ _80931_/CLK _68515_/X _83972_/Q sky130_fd_sc_hd__dfxtp_4
X_50014_ _50027_/A _53227_/B _50014_/Y sky130_fd_sc_hd__nand2_4
X_85711_ _84766_/CLK _53024_/Y _85711_/Q sky130_fd_sc_hd__dfxtp_4
X_82923_ _82923_/CLK _78197_/X _82923_/Q sky130_fd_sc_hd__dfxtp_4
X_55871_ _45107_/A _55531_/X _55533_/X _55870_/X _55871_/X sky130_fd_sc_hd__a211o_4
X_67857_ _87453_/Q _67834_/X _67835_/X _67856_/X _67857_/X sky130_fd_sc_hd__a211o_4
X_86691_ _86372_/CLK _86691_/D _58953_/A sky130_fd_sc_hd__dfxtp_4
X_57610_ _57606_/Y _57581_/X _57609_/Y _57610_/Y sky130_fd_sc_hd__a21boi_4
X_54822_ _54819_/Y _54802_/X _54821_/X _85372_/D sky130_fd_sc_hd__a21oi_4
X_66808_ _66760_/A _66808_/B _66808_/X sky130_fd_sc_hd__and2_4
X_85642_ _85738_/CLK _53394_/Y _85642_/Q sky130_fd_sc_hd__dfxtp_4
X_58590_ _58585_/X _58587_/Y _58588_/Y _58098_/X _58589_/X _58590_/X
+ sky130_fd_sc_hd__o32a_4
X_82854_ _82855_/CLK _78102_/B _82854_/Q sky130_fd_sc_hd__dfxtp_4
X_67788_ _67550_/X _67788_/X sky130_fd_sc_hd__buf_2
X_57541_ _57528_/X _53514_/B _57541_/Y sky130_fd_sc_hd__nand2_4
X_81805_ _81620_/CLK _81613_/Q _81805_/Q sky130_fd_sc_hd__dfxtp_4
X_69527_ _87011_/Q _69485_/X _69361_/X _69526_/X _69527_/X sky130_fd_sc_hd__a211o_4
X_88361_ _82541_/CLK _88361_/D _88361_/Q sky130_fd_sc_hd__dfxtp_4
X_54753_ _54807_/A _54775_/A sky130_fd_sc_hd__buf_2
X_66739_ _87372_/Q _66642_/X _66643_/X _66738_/X _66739_/X sky130_fd_sc_hd__a211o_4
X_85573_ _83564_/CLK _85573_/D _85573_/Q sky130_fd_sc_hd__dfxtp_4
X_51965_ _51963_/Y _51934_/X _51964_/Y _85916_/D sky130_fd_sc_hd__a21boi_4
X_82785_ _82973_/CLK _82785_/D _82785_/Q sky130_fd_sc_hd__dfxtp_4
X_87312_ _86534_/CLK _43681_/X _72831_/A sky130_fd_sc_hd__dfxtp_4
X_53704_ _53700_/Y _53680_/X _53703_/X _85585_/D sky130_fd_sc_hd__a21oi_4
X_84524_ _81048_/CLK _84524_/D _84524_/Q sky130_fd_sc_hd__dfxtp_4
X_50916_ _50932_/A _51779_/B _50916_/Y sky130_fd_sc_hd__nand2_4
X_57472_ _57472_/A _84998_/D sky130_fd_sc_hd__inv_2
X_81736_ _82067_/CLK _81736_/D _41422_/A sky130_fd_sc_hd__dfxtp_4
X_69458_ _69183_/A _69458_/X sky130_fd_sc_hd__buf_2
X_88292_ _87790_/CLK _88292_/D _88292_/Q sky130_fd_sc_hd__dfxtp_4
X_54684_ _54656_/X _54707_/B sky130_fd_sc_hd__buf_2
X_51896_ _85926_/Q _51873_/X _51895_/Y _51896_/Y sky130_fd_sc_hd__o21ai_4
X_59211_ _59207_/Y _59210_/Y _59165_/X _59211_/X sky130_fd_sc_hd__a21o_4
X_56423_ _56436_/A _56433_/B sky130_fd_sc_hd__buf_2
X_68409_ _68409_/A _88274_/Q _68409_/X sky130_fd_sc_hd__and2_4
X_87243_ _87757_/CLK _43835_/X _87243_/Q sky130_fd_sc_hd__dfxtp_4
X_53635_ _53671_/A _53667_/C sky130_fd_sc_hd__buf_2
X_84455_ _84564_/CLK _61769_/Y _78078_/B sky130_fd_sc_hd__dfxtp_4
X_50847_ _50806_/A _51358_/B _50847_/Y sky130_fd_sc_hd__nand2_4
X_81667_ _81040_/CLK _80262_/X _81667_/Q sky130_fd_sc_hd__dfxtp_4
X_69389_ _68660_/X _69389_/X sky130_fd_sc_hd__buf_2
X_40600_ _40590_/X _40596_/X _88368_/Q _40599_/X _40600_/X sky130_fd_sc_hd__a2bb2o_4
X_71420_ _71419_/Y _71420_/X sky130_fd_sc_hd__buf_2
X_59142_ _84766_/Q _59129_/X _59134_/X _59141_/X _59142_/Y sky130_fd_sc_hd__a2bb2oi_4
X_83406_ _83482_/CLK _71701_/Y _83406_/Q sky130_fd_sc_hd__dfxtp_4
X_80618_ _80608_/A _80608_/B _80607_/A _80607_/B _80618_/X sky130_fd_sc_hd__o22a_4
X_56354_ _56358_/A _56358_/B _55748_/B _56354_/Y sky130_fd_sc_hd__nand3_4
X_87174_ _87174_/CLK _44281_/Y _87174_/Q sky130_fd_sc_hd__dfxtp_4
X_41580_ _41580_/A _41580_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_490_0_CLK clkbuf_9_245_0_CLK/X _85959_/CLK sky130_fd_sc_hd__clkbuf_1
X_53566_ _53564_/Y _53524_/X _53565_/Y _53566_/Y sky130_fd_sc_hd__a21boi_4
X_84386_ _84508_/CLK _84386_/D _84386_/Q sky130_fd_sc_hd__dfxtp_4
X_50778_ _86135_/Q _50775_/X _50777_/Y _50778_/Y sky130_fd_sc_hd__o21ai_4
X_81598_ _81482_/CLK _65481_/C _76915_/A sky130_fd_sc_hd__dfxtp_4
X_55305_ _55190_/X _55305_/X sky130_fd_sc_hd__buf_2
X_86125_ _86040_/CLK _86125_/D _86125_/Q sky130_fd_sc_hd__dfxtp_4
X_40531_ _40429_/X _82309_/Q _40530_/X _40531_/X sky130_fd_sc_hd__o21a_4
X_52517_ _52602_/A _52518_/A sky130_fd_sc_hd__buf_2
X_59073_ _58904_/A _59073_/X sky130_fd_sc_hd__buf_2
X_71351_ _70935_/A _71351_/X sky130_fd_sc_hd__buf_2
X_83337_ _83337_/CLK _83337_/D _83337_/Q sky130_fd_sc_hd__dfxtp_4
X_56285_ _56282_/Y _56347_/A sky130_fd_sc_hd__buf_2
X_80549_ _80547_/X _80549_/B _80549_/Y sky130_fd_sc_hd__xnor2_4
X_53497_ _53798_/A _53696_/A sky130_fd_sc_hd__buf_2
X_58024_ _84932_/Q _57896_/X _58016_/X _58023_/X _84932_/D sky130_fd_sc_hd__a2bb2oi_4
X_70302_ _70289_/X _74770_/A _70301_/X _83805_/D sky130_fd_sc_hd__a21o_4
X_55236_ _45847_/A _55244_/A _55158_/A _55235_/X _55655_/B sky130_fd_sc_hd__a211o_4
X_43250_ _43212_/A _43250_/X sky130_fd_sc_hd__buf_2
X_74070_ _70111_/Y _74003_/B _74069_/X _74070_/Y sky130_fd_sc_hd__o21ai_4
X_86056_ _85643_/CLK _86056_/D _86056_/Q sky130_fd_sc_hd__dfxtp_4
X_52448_ _52448_/A _46313_/Y _52448_/Y sky130_fd_sc_hd__nand2_4
X_40462_ _40380_/A _40931_/A sky130_fd_sc_hd__buf_2
X_71282_ _53209_/B _71264_/X _71281_/Y _83548_/D sky130_fd_sc_hd__o21ai_4
X_83268_ _83630_/CLK _83268_/D _83268_/Q sky130_fd_sc_hd__dfxtp_4
X_42201_ _42096_/A _42201_/X sky130_fd_sc_hd__buf_2
X_73021_ _73019_/X _73021_/B _73021_/C _73021_/Y sky130_fd_sc_hd__nand3_4
X_85007_ _85034_/CLK _85007_/D _57419_/A sky130_fd_sc_hd__dfxtp_4
X_70233_ _70233_/A _70239_/D sky130_fd_sc_hd__buf_2
X_82219_ _81928_/CLK _82251_/Q _77354_/A sky130_fd_sc_hd__dfxtp_4
X_43181_ _43013_/X _51340_/A sky130_fd_sc_hd__buf_2
X_55167_ _45719_/A _44059_/A _55165_/X _55166_/X _55167_/X sky130_fd_sc_hd__a211o_4
X_40393_ _40368_/X _81180_/Q _40393_/X sky130_fd_sc_hd__or2_4
X_52379_ _52373_/X _50169_/B _52379_/Y sky130_fd_sc_hd__nand2_4
X_83199_ _83835_/CLK _83199_/D _83199_/Q sky130_fd_sc_hd__dfxtp_4
X_42132_ _42132_/A _88019_/D sky130_fd_sc_hd__inv_2
X_54118_ _53357_/A _54118_/X sky130_fd_sc_hd__buf_2
X_70164_ _70348_/D _70164_/X sky130_fd_sc_hd__buf_2
X_55098_ _47841_/A _55098_/X sky130_fd_sc_hd__buf_2
X_59975_ _59910_/X _59976_/A sky130_fd_sc_hd__buf_2
X_58926_ _58877_/X _85925_/Q _58900_/X _58926_/X sky130_fd_sc_hd__o21a_4
X_46940_ _47081_/A _46940_/X sky130_fd_sc_hd__buf_2
X_42063_ _42063_/A _42063_/Y sky130_fd_sc_hd__inv_2
X_54049_ _54037_/A _46500_/Y _54049_/Y sky130_fd_sc_hd__nand2_4
X_77760_ _77757_/X _77759_/Y _77761_/B sky130_fd_sc_hd__xor2_4
X_86958_ _86965_/CLK _86958_/D _86958_/Q sky130_fd_sc_hd__dfxtp_4
X_74972_ _74963_/B _74972_/B _74972_/Y sky130_fd_sc_hd__nand2_4
X_70095_ _69117_/X _69119_/X _69156_/X _70095_/Y sky130_fd_sc_hd__a21oi_4
X_41014_ _41014_/A _41019_/B _41014_/X sky130_fd_sc_hd__or2_4
X_76711_ _76709_/X _76710_/Y _76711_/Y sky130_fd_sc_hd__nor2_4
X_85909_ _86549_/CLK _85909_/D _66082_/B sky130_fd_sc_hd__dfxtp_4
X_73923_ _73919_/X _73922_/X _73421_/X _73923_/X sky130_fd_sc_hd__a21o_4
X_46871_ _52722_/B _51031_/B sky130_fd_sc_hd__buf_2
X_58857_ _58857_/A _58857_/X sky130_fd_sc_hd__buf_2
X_77691_ _77690_/Y _77692_/B sky130_fd_sc_hd__inv_2
X_86889_ _86861_/CLK _45249_/Y _64466_/B sky130_fd_sc_hd__dfxtp_4
X_48610_ _50511_/A _48624_/B _48610_/C _48610_/X sky130_fd_sc_hd__and3_4
X_79430_ _79416_/A _79416_/B _79430_/X sky130_fd_sc_hd__or2_4
X_45822_ _45814_/X _45818_/Y _45821_/Y _86852_/D sky130_fd_sc_hd__a21oi_4
X_57808_ _86652_/Q _57833_/B _57808_/Y sky130_fd_sc_hd__nor2_4
X_76642_ _81377_/Q _76642_/Y sky130_fd_sc_hd__inv_2
X_49590_ _49580_/X _52803_/B _49590_/Y sky130_fd_sc_hd__nand2_4
X_73854_ _74012_/A _73854_/X sky130_fd_sc_hd__buf_2
X_58788_ _58682_/X _85776_/Q _58706_/X _58788_/X sky130_fd_sc_hd__o21a_4
X_48541_ _86513_/Q _48536_/X _48540_/Y _48541_/Y sky130_fd_sc_hd__o21ai_4
X_72805_ _44520_/Y _72775_/X _72804_/Y _72822_/C sky130_fd_sc_hd__a21o_4
Xclkbuf_10_443_0_CLK clkbuf_9_221_0_CLK/X _84194_/CLK sky130_fd_sc_hd__clkbuf_1
X_79361_ _58755_/Y _66445_/C _79360_/Y _79361_/X sky130_fd_sc_hd__o21a_4
X_45753_ _85066_/Q _45736_/B _45753_/Y sky130_fd_sc_hd__nor2_4
X_57739_ _57711_/X _57739_/X sky130_fd_sc_hd__buf_2
X_76573_ _81278_/Q _81546_/Q _76576_/B sky130_fd_sc_hd__nor2_4
X_42965_ _40408_/X _42962_/X _87627_/Q _42963_/X _87627_/D sky130_fd_sc_hd__a2bb2o_4
X_73785_ _73781_/X _73784_/X _73738_/X _73789_/A sky130_fd_sc_hd__a21o_4
X_70997_ _70997_/A _71082_/B sky130_fd_sc_hd__buf_2
X_78312_ _78312_/A _82658_/D _78312_/X sky130_fd_sc_hd__xor2_4
X_44704_ _44704_/A _86993_/D sky130_fd_sc_hd__inv_2
X_75524_ _75519_/X _75524_/B _75520_/Y _75524_/Y sky130_fd_sc_hd__nand3_4
X_41916_ _41894_/X _41879_/X _40641_/X _88106_/Q _41882_/X _41917_/A
+ sky130_fd_sc_hd__o32ai_4
X_48472_ _48472_/A _48473_/A sky130_fd_sc_hd__inv_2
X_60750_ _60727_/A _60132_/A _60749_/Y _60750_/X sky130_fd_sc_hd__and3_4
X_72736_ _72735_/X _72737_/A sky130_fd_sc_hd__buf_2
X_79292_ _79281_/X _79292_/B _79292_/X sky130_fd_sc_hd__and2_4
X_45684_ _63217_/B _61551_/A sky130_fd_sc_hd__buf_2
X_42896_ _42945_/A _42896_/X sky130_fd_sc_hd__buf_2
X_47423_ _86636_/Q _47382_/X _47422_/Y _47423_/Y sky130_fd_sc_hd__o21ai_4
X_59409_ _84740_/Q _63161_/A sky130_fd_sc_hd__inv_2
X_78243_ _78241_/X _78252_/C _78246_/A sky130_fd_sc_hd__nand2_4
X_44635_ _44634_/Y _87024_/D sky130_fd_sc_hd__inv_2
X_75455_ _80700_/Q _80956_/D _75456_/A sky130_fd_sc_hd__nand2_4
X_41847_ _48164_/A _41847_/X sky130_fd_sc_hd__buf_2
X_72667_ _83197_/Q _72658_/X _72666_/Y _83197_/D sky130_fd_sc_hd__a21bo_4
X_60681_ _60652_/X _60682_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_458_0_CLK clkbuf_9_229_0_CLK/X _83630_/CLK sky130_fd_sc_hd__clkbuf_1
X_74406_ _74406_/A _74395_/X _74421_/C _74406_/X sky130_fd_sc_hd__and3_4
X_62420_ _61500_/X _62420_/B _62420_/C _62404_/X _62421_/D sky130_fd_sc_hd__nand4_4
X_47354_ _86643_/Q _47332_/X _47353_/Y _47354_/Y sky130_fd_sc_hd__o21ai_4
X_71618_ _71863_/A _70667_/A _71614_/C _71622_/D _71618_/Y sky130_fd_sc_hd__nor4_4
X_78174_ _78193_/B _78174_/B _78191_/A sky130_fd_sc_hd__xor2_4
X_44566_ _42081_/A _44567_/A sky130_fd_sc_hd__buf_2
X_75386_ _75383_/X _75386_/B _75390_/A sky130_fd_sc_hd__nand2_4
X_41778_ _41777_/Y _41778_/X sky130_fd_sc_hd__buf_2
X_72598_ _72581_/A _72573_/B _79310_/B _72598_/Y sky130_fd_sc_hd__nor3_4
X_46305_ _53964_/A _51256_/A sky130_fd_sc_hd__buf_2
X_77125_ _77111_/X _77122_/A _77125_/X sky130_fd_sc_hd__and2_4
X_43517_ _43516_/Y _87381_/D sky130_fd_sc_hd__inv_2
X_62351_ _62634_/A _62351_/B _62351_/C _62351_/D _62351_/Y sky130_fd_sc_hd__nand4_4
X_74337_ _70323_/C _74327_/X _74336_/Y _74337_/X sky130_fd_sc_hd__a21bo_4
X_40729_ _40729_/A _40729_/X sky130_fd_sc_hd__buf_2
X_47285_ _47280_/Y _47271_/X _47284_/X _86651_/D sky130_fd_sc_hd__a21oi_4
X_71549_ _71530_/Y _83460_/Q _71548_/Y _71549_/X sky130_fd_sc_hd__a21o_4
X_44497_ _44548_/A _44497_/X sky130_fd_sc_hd__buf_2
X_49024_ _83611_/Q _53852_/B sky130_fd_sc_hd__inv_2
X_61302_ _61302_/A _61302_/Y sky130_fd_sc_hd__inv_2
X_46236_ _56777_/B _46237_/A sky130_fd_sc_hd__buf_2
X_65070_ _64939_/A _65070_/X sky130_fd_sc_hd__buf_2
XPHY_480 sky130_fd_sc_hd__decap_3
X_77056_ _77054_/A _82281_/D _77055_/Y _77056_/Y sky130_fd_sc_hd__a21oi_4
X_43448_ _41601_/X _43446_/X _87416_/Q _43447_/X _43448_/X sky130_fd_sc_hd__a2bb2o_4
X_62282_ _62271_/X _62275_/Y _62281_/X _58162_/A _62214_/X _62282_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74268_ _74265_/X _74267_/X _72741_/X _74268_/X sky130_fd_sc_hd__a21o_4
XPHY_491 sky130_fd_sc_hd__decap_3
X_76007_ _76005_/B _81708_/D _81420_/Q _76008_/A sky130_fd_sc_hd__nand3_4
X_64021_ _64017_/X _63969_/X _64018_/Y _64019_/Y _64020_/X _64021_/X
+ sky130_fd_sc_hd__a41o_4
X_61233_ _61232_/X _61107_/X _61176_/B _61264_/A sky130_fd_sc_hd__nand3_4
X_73219_ _73220_/B _73220_/C _73218_/X _73219_/X sky130_fd_sc_hd__a21o_4
X_46167_ _46167_/A _46167_/B _46159_/X _46167_/Y sky130_fd_sc_hd__nor3_4
X_43379_ _43367_/X _43375_/X _41408_/X _87452_/Q _43378_/X _43379_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74199_ _74199_/A _74198_/X _74200_/B sky130_fd_sc_hd__nand2_4
X_45118_ _56414_/C _45102_/X _45117_/X _45118_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_502_0_CLK clkbuf_9_502_0_CLK/A clkbuf_9_502_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_61164_ _72564_/A _61165_/B sky130_fd_sc_hd__buf_2
X_46098_ _46098_/A _40381_/X _46109_/A sky130_fd_sc_hd__nand2_4
X_60115_ _59971_/X _60049_/Y _60113_/Y _62203_/A _60114_/Y _84659_/D
+ sky130_fd_sc_hd__a41oi_4
X_49926_ _49925_/X _49915_/X _49904_/C _53139_/D _49926_/X sky130_fd_sc_hd__and4_4
X_45049_ _44972_/X _45049_/X sky130_fd_sc_hd__buf_2
X_68760_ _87492_/Q _68757_/X _68731_/X _68759_/X _68760_/X sky130_fd_sc_hd__a211o_4
X_65972_ _65702_/A _65972_/B _65972_/X sky130_fd_sc_hd__and2_4
X_61095_ _61153_/A _61095_/X sky130_fd_sc_hd__buf_2
X_77958_ _82171_/Q _77958_/B _77958_/X sky130_fd_sc_hd__xor2_4
X_67711_ _67496_/X _67698_/Y _67624_/X _67710_/Y _67711_/X sky130_fd_sc_hd__a211o_4
X_64923_ _64923_/A _64924_/A sky130_fd_sc_hd__buf_2
X_60046_ _59852_/A _60081_/B sky130_fd_sc_hd__buf_2
X_76909_ _76931_/A _76914_/A sky130_fd_sc_hd__inv_2
X_49857_ _49851_/A _49851_/B _49862_/C _53070_/D _49857_/X sky130_fd_sc_hd__and4_4
X_68691_ _69567_/A _68691_/X sky130_fd_sc_hd__buf_2
X_77889_ _82068_/Q _77891_/A sky130_fd_sc_hd__inv_2
X_48808_ _48808_/A _48836_/A sky130_fd_sc_hd__buf_2
X_67642_ _67569_/X _87718_/Q _67642_/X sky130_fd_sc_hd__and2_4
X_79628_ _84209_/Q _83257_/Q _79630_/A sky130_fd_sc_hd__xor2_4
X_64854_ _64797_/X _83304_/Q _64772_/X _64853_/X _64854_/X sky130_fd_sc_hd__a211o_4
X_49788_ _49678_/X _49807_/A sky130_fd_sc_hd__buf_2
X_63805_ _63049_/B _63790_/X _63757_/C _63776_/X _63805_/Y sky130_fd_sc_hd__nand4_4
X_48739_ _48801_/A _48416_/A _48739_/X sky130_fd_sc_hd__and2_4
Xclkbuf_8_70_0_CLK clkbuf_8_71_0_CLK/A clkbuf_8_70_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_67573_ _87401_/Q _67476_/X _67477_/X _67572_/X _67573_/X sky130_fd_sc_hd__a211o_4
X_79559_ _79548_/Y _79558_/Y _79559_/Y sky130_fd_sc_hd__nor2_4
X_64785_ _64657_/X _86747_/Q _64733_/X _64784_/X _64785_/X sky130_fd_sc_hd__a211o_4
X_61997_ _58254_/A _61997_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_2_0_CLK clkbuf_7_3_0_CLK/A clkbuf_8_5_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_69312_ _68685_/X _68687_/X _69295_/X _69312_/Y sky130_fd_sc_hd__a21oi_4
X_66524_ _64867_/B _66524_/B _66524_/C _66524_/X sky130_fd_sc_hd__and3_4
X_51750_ _51768_/A _51749_/X _51750_/C _52580_/D _51750_/X sky130_fd_sc_hd__and4_4
X_63736_ _64136_/B _63736_/X sky130_fd_sc_hd__buf_2
X_82570_ _82570_/CLK _82602_/Q _82570_/Q sky130_fd_sc_hd__dfxtp_4
X_60948_ _60933_/X _60938_/Y _61024_/B _60944_/Y _60947_/Y _84549_/D
+ sky130_fd_sc_hd__a41oi_4
X_50701_ _50698_/Y _50699_/X _50700_/Y _86151_/D sky130_fd_sc_hd__a21boi_4
X_81521_ _82642_/CLK _76366_/B _76032_/A sky130_fd_sc_hd__dfxtp_4
X_69243_ _68929_/X _68551_/Y _69231_/X _69242_/Y _69243_/X sky130_fd_sc_hd__a211o_4
X_66455_ _66453_/Y _66454_/Y _65842_/X _66455_/Y sky130_fd_sc_hd__a21oi_4
X_51681_ _51697_/A _53205_/B _51681_/Y sky130_fd_sc_hd__nand2_4
X_63667_ _58976_/A _60667_/A _60724_/A _62577_/Y _60663_/Y _63667_/Y
+ sky130_fd_sc_hd__o32ai_4
X_60879_ _60934_/A _60879_/B _60863_/X _60879_/D _60879_/Y sky130_fd_sc_hd__nand4_4
X_53420_ _53420_/A _53402_/B _53410_/C _51214_/D _53420_/X sky130_fd_sc_hd__and4_4
X_65406_ _44170_/A _65407_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_85_0_CLK clkbuf_8_85_0_CLK/A clkbuf_8_85_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_84240_ _82436_/CLK _84240_/D _84240_/Q sky130_fd_sc_hd__dfxtp_4
X_50632_ _50627_/X _49025_/X _50632_/Y sky130_fd_sc_hd__nand2_4
X_62618_ _62269_/X _58210_/X _62618_/C _62618_/D _62618_/X sky130_fd_sc_hd__and4_4
X_81452_ _81433_/CLK _76745_/B _81452_/Q sky130_fd_sc_hd__dfxtp_4
X_69174_ _69146_/X _69109_/X _69172_/Y _69173_/Y _69174_/X sky130_fd_sc_hd__a211o_4
X_66386_ _66282_/X _65983_/Y _66385_/Y _66386_/Y sky130_fd_sc_hd__o21ai_4
X_63598_ _63598_/A _63630_/B _63630_/C _63598_/Y sky130_fd_sc_hd__nor3_4
X_80403_ _80425_/A _80409_/A sky130_fd_sc_hd__inv_2
X_68125_ _66800_/X _66803_/X _68106_/X _68125_/Y sky130_fd_sc_hd__a21oi_4
X_53351_ _53351_/A _53351_/X sky130_fd_sc_hd__buf_2
X_65337_ _65285_/A _65337_/B _65337_/X sky130_fd_sc_hd__and2_4
X_84171_ _81233_/CLK _84171_/D _84171_/Q sky130_fd_sc_hd__dfxtp_4
X_50563_ _50506_/A _50563_/X sky130_fd_sc_hd__buf_2
X_62549_ _62549_/A _62561_/B _62548_/Y _62549_/Y sky130_fd_sc_hd__nand3_4
X_81383_ _83918_/CLK _81383_/D _76840_/B sky130_fd_sc_hd__dfxtp_4
Xpsn_inst_psn_buff_8 _71216_/A _71231_/A2 sky130_fd_sc_hd__buf_2
X_52302_ _52300_/Y _52289_/X _52301_/X _52302_/Y sky130_fd_sc_hd__a21oi_4
X_83122_ _86213_/CLK _83122_/D _83122_/Q sky130_fd_sc_hd__dfxtp_4
X_80334_ _80331_/Y _80333_/Y _80334_/Y sky130_fd_sc_hd__nand2_4
X_56070_ _56069_/Y _56070_/X sky130_fd_sc_hd__buf_2
X_68056_ _68052_/X _68055_/X _68033_/X _68056_/X sky130_fd_sc_hd__a21o_4
X_53282_ _53282_/A _53311_/A sky130_fd_sc_hd__buf_2
X_65268_ _65268_/A _65268_/B _65268_/C _65268_/X sky130_fd_sc_hd__and3_4
X_50494_ _50465_/X _48816_/B _50494_/Y sky130_fd_sc_hd__nand2_4
X_55021_ _54250_/A _55037_/A sky130_fd_sc_hd__buf_2
X_67007_ _87937_/Q _66935_/X _66911_/X _67006_/X _67007_/X sky130_fd_sc_hd__a211o_4
X_52233_ _48849_/A _52248_/B _52223_/C _52233_/X sky130_fd_sc_hd__and3_4
X_64219_ _63380_/A _64219_/B _64219_/Y sky130_fd_sc_hd__nor2_4
X_83053_ _83310_/CLK _74502_/Y _83053_/Q sky130_fd_sc_hd__dfxtp_4
X_87930_ _87110_/CLK _87930_/D _87930_/Q sky130_fd_sc_hd__dfxtp_4
X_80265_ _80268_/B _80265_/Y sky130_fd_sc_hd__inv_2
X_65199_ _64666_/A _65199_/X sky130_fd_sc_hd__buf_2
X_82004_ _82008_/CLK _82036_/Q _77143_/B sky130_fd_sc_hd__dfxtp_4
X_52164_ _85876_/Q _52152_/X _52163_/Y _52164_/Y sky130_fd_sc_hd__o21ai_4
X_87861_ _87348_/CLK _87861_/D _87861_/Q sky130_fd_sc_hd__dfxtp_4
X_80196_ _80196_/A _80195_/X _80209_/B sky130_fd_sc_hd__xnor2_4
X_51115_ _51115_/A _51115_/B _51115_/C _52805_/D _51115_/X sky130_fd_sc_hd__and4_4
X_86812_ _81182_/CLK _86812_/D _67201_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_23_0_CLK clkbuf_8_23_0_CLK/A clkbuf_9_47_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_59760_ _59699_/A _59761_/B sky130_fd_sc_hd__buf_2
X_52095_ _52100_/A _48358_/X _52095_/Y sky130_fd_sc_hd__nand2_4
X_56972_ _56972_/A _56650_/Y _56972_/Y sky130_fd_sc_hd__nand2_4
X_68958_ _68384_/A _68958_/X sky130_fd_sc_hd__buf_2
X_87792_ _88084_/CLK _42640_/X _69176_/B sky130_fd_sc_hd__dfxtp_4
X_58711_ _84805_/Q _58711_/Y sky130_fd_sc_hd__inv_2
X_51046_ _51044_/Y _51039_/X _51045_/X _51046_/Y sky130_fd_sc_hd__a21oi_4
X_55923_ _55920_/X _55922_/X _44118_/B _55926_/A sky130_fd_sc_hd__a21o_4
X_67909_ _67909_/A _67909_/B _67909_/X sky130_fd_sc_hd__and2_4
X_86743_ _85527_/CLK _46375_/Y _86743_/Q sky130_fd_sc_hd__dfxtp_4
X_59691_ _59816_/A _59691_/X sky130_fd_sc_hd__buf_2
X_83955_ _83957_/CLK _68928_/X _83955_/Q sky130_fd_sc_hd__dfxtp_4
X_68889_ _74053_/A _68493_/X _68494_/X _68888_/Y _68889_/X sky130_fd_sc_hd__a211o_4
X_70920_ _51026_/B _70909_/X _70919_/Y _83663_/D sky130_fd_sc_hd__o21ai_4
X_58642_ _58641_/X _85947_/Q _58109_/X _58642_/X sky130_fd_sc_hd__o21a_4
X_82906_ _82906_/CLK _78257_/B _41319_/B sky130_fd_sc_hd__dfxtp_4
X_55854_ _55853_/X _55854_/X sky130_fd_sc_hd__buf_2
X_86674_ _86353_/CLK _47068_/Y _59189_/A sky130_fd_sc_hd__dfxtp_4
X_83886_ _82339_/CLK _69928_/X _83886_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_38_0_CLK clkbuf_8_39_0_CLK/A clkbuf_8_38_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_54805_ _54790_/A _47552_/A _54805_/Y sky130_fd_sc_hd__nand2_4
X_85625_ _86235_/CLK _53500_/Y _85625_/Q sky130_fd_sc_hd__dfxtp_4
X_70851_ _70832_/A _70852_/C sky130_fd_sc_hd__buf_2
X_58573_ _58140_/X _86113_/Q _58572_/X _58573_/Y sky130_fd_sc_hd__o21ai_4
X_82837_ _84177_/CLK _82837_/D _82837_/Q sky130_fd_sc_hd__dfxtp_4
X_55785_ _55794_/A _56523_/C _55785_/X sky130_fd_sc_hd__and2_4
X_52997_ _52997_/A _52997_/B _52997_/C _52997_/D _52997_/X sky130_fd_sc_hd__and4_4
X_57524_ _84986_/Q _47806_/X _57523_/Y _57524_/Y sky130_fd_sc_hd__o21ai_4
X_88344_ _88345_/CLK _40740_/X _88344_/Q sky130_fd_sc_hd__dfxtp_4
X_54736_ _54731_/X _47431_/Y _54736_/Y sky130_fd_sc_hd__nand2_4
X_42750_ _42700_/A _42750_/X sky130_fd_sc_hd__buf_2
X_73570_ _73570_/A _73569_/X _73570_/Y sky130_fd_sc_hd__nand2_4
X_85556_ _85556_/CLK _85556_/D _85556_/Q sky130_fd_sc_hd__dfxtp_4
X_51948_ _73636_/B _51945_/X _51947_/Y _51948_/Y sky130_fd_sc_hd__o21ai_4
X_70782_ _70782_/A _70871_/A sky130_fd_sc_hd__buf_2
X_82768_ _82768_/CLK _82768_/D _82960_/D sky130_fd_sc_hd__dfxtp_4
X_41701_ _41700_/Y _41701_/X sky130_fd_sc_hd__buf_2
X_72521_ _79502_/B _61252_/X _72517_/Y _72520_/X _72521_/X sky130_fd_sc_hd__o22a_4
X_84507_ _84507_/CLK _84507_/D _75909_/A sky130_fd_sc_hd__dfxtp_4
X_81719_ _81532_/CLK _81719_/D _40984_/B sky130_fd_sc_hd__dfxtp_4
X_57455_ _57331_/A _57470_/B _57331_/C _57455_/Y sky130_fd_sc_hd__nand3_4
X_88275_ _88263_/CLK _88275_/D _88275_/Q sky130_fd_sc_hd__dfxtp_4
X_42681_ _42681_/A _42681_/X sky130_fd_sc_hd__buf_2
X_54667_ _54667_/A _54674_/B _54644_/X _47310_/A _54667_/X sky130_fd_sc_hd__and4_4
X_85487_ _83736_/CLK _54192_/Y _85487_/Q sky130_fd_sc_hd__dfxtp_4
X_51879_ _51876_/Y _51877_/X _51878_/X _85930_/D sky130_fd_sc_hd__a21oi_4
X_82699_ _84111_/CLK _82699_/D _82687_/D sky130_fd_sc_hd__dfxtp_4
X_44420_ _41556_/X _44412_/X _87117_/Q _44413_/X _44420_/X sky130_fd_sc_hd__a2bb2o_4
X_56406_ _56064_/X _56394_/X _56405_/Y _56406_/Y sky130_fd_sc_hd__o21ai_4
X_75240_ _75240_/A _75251_/A _75240_/X sky130_fd_sc_hd__xor2_4
X_41632_ _41611_/X _41613_/X _41631_/X _67349_/B _41608_/X _41632_/Y
+ sky130_fd_sc_hd__o32ai_4
X_87226_ _88002_/CLK _43871_/X _68980_/B sky130_fd_sc_hd__dfxtp_4
X_53618_ _53798_/A _53747_/A sky130_fd_sc_hd__buf_2
X_72452_ _57697_/X _85957_/Q _72451_/X _72452_/Y sky130_fd_sc_hd__o21ai_4
X_84438_ _84438_/CLK _62035_/Y _78061_/B sky130_fd_sc_hd__dfxtp_4
X_57386_ _57384_/X _56571_/X _85024_/Q _57385_/X _85024_/D sky130_fd_sc_hd__a2bb2o_4
X_54598_ _54589_/X _54585_/B _54591_/C _47189_/A _54598_/X sky130_fd_sc_hd__and4_4
X_59125_ _59073_/X _85751_/Q _59124_/X _59125_/X sky130_fd_sc_hd__o21a_4
X_71403_ _71342_/B _71411_/C sky130_fd_sc_hd__buf_2
X_56337_ _56350_/A _56337_/X sky130_fd_sc_hd__buf_2
X_44351_ _44382_/A _44351_/X sky130_fd_sc_hd__buf_2
X_75171_ _75175_/C _75171_/Y sky130_fd_sc_hd__inv_2
X_87157_ _87915_/CLK _44342_/Y _87157_/Q sky130_fd_sc_hd__dfxtp_4
X_41563_ _41563_/A _41563_/B _41563_/X sky130_fd_sc_hd__or2_4
X_72383_ _57696_/X _72428_/B sky130_fd_sc_hd__buf_2
X_53549_ _85615_/Q _53540_/X _53548_/Y _53549_/Y sky130_fd_sc_hd__o21ai_4
X_84369_ _84449_/CLK _84369_/D _84369_/Q sky130_fd_sc_hd__dfxtp_4
X_43302_ _43302_/A _43302_/X sky130_fd_sc_hd__buf_2
X_74122_ _68956_/B _44235_/X _72725_/A _74121_/Y _74122_/X sky130_fd_sc_hd__a211o_4
X_86108_ _85786_/CLK _50915_/Y _86108_/Q sky130_fd_sc_hd__dfxtp_4
X_40514_ _40512_/X _41584_/A _40513_/X _40514_/X sky130_fd_sc_hd__o21a_4
X_47070_ _53353_/B _52837_/B sky130_fd_sc_hd__buf_2
X_59056_ _59029_/A _86364_/Q _59056_/Y sky130_fd_sc_hd__nor2_4
X_71334_ _50378_/B _71320_/A _71333_/Y _71334_/Y sky130_fd_sc_hd__o21ai_4
X_44282_ _44038_/X _44282_/X sky130_fd_sc_hd__buf_2
X_56268_ _56164_/X _56188_/X _56267_/Y _56268_/Y sky130_fd_sc_hd__o21ai_4
X_41494_ _41489_/X _41490_/X _41493_/X _66718_/B _41474_/X _41494_/Y
+ sky130_fd_sc_hd__o32ai_4
X_87088_ _88263_/CLK _87088_/D _87088_/Q sky130_fd_sc_hd__dfxtp_4
X_46021_ _46021_/A _46021_/Y sky130_fd_sc_hd__inv_2
X_58007_ _58007_/A _58007_/X sky130_fd_sc_hd__buf_2
X_43233_ _43226_/X _43229_/X _41009_/X _87526_/Q _43232_/X _43234_/A
+ sky130_fd_sc_hd__o32ai_4
X_55219_ _55149_/A _55219_/B _55219_/X sky130_fd_sc_hd__and2_4
X_74053_ _74053_/A _72853_/X _74053_/Y sky130_fd_sc_hd__nor2_4
X_78930_ _78928_/Y _78930_/B _78938_/A sky130_fd_sc_hd__xor2_4
X_86039_ _85527_/CLK _86039_/D _64874_/B sky130_fd_sc_hd__dfxtp_4
X_40445_ _40429_/X _82324_/Q _40444_/X _40445_/X sky130_fd_sc_hd__o21a_4
X_71265_ _71264_/X _71265_/X sky130_fd_sc_hd__buf_2
X_56199_ _56188_/X _56016_/X _56198_/Y _85279_/D sky130_fd_sc_hd__o21ai_4
X_73004_ _43137_/Y _72830_/X _72799_/X _73003_/Y _73004_/X sky130_fd_sc_hd__a211o_4
X_70216_ _70231_/A _70229_/A sky130_fd_sc_hd__buf_2
X_43164_ _43164_/A _43164_/Y sky130_fd_sc_hd__inv_2
X_78861_ _78866_/A _78860_/Y _78862_/B sky130_fd_sc_hd__xor2_4
X_40376_ _57491_/A _40364_/X _40371_/X _88401_/Q _40375_/X _40376_/Y
+ sky130_fd_sc_hd__o32ai_4
X_71196_ _71196_/A _71197_/C sky130_fd_sc_hd__buf_2
X_42115_ _41070_/X _42103_/X _88027_/Q _42104_/X _42115_/X sky130_fd_sc_hd__a2bb2o_4
X_77812_ _82155_/Q _77812_/B _77812_/X sky130_fd_sc_hd__xor2_4
X_70147_ _83523_/Q _83171_/Q _83498_/Q _83146_/Q _70147_/Y sky130_fd_sc_hd__a22oi_4
X_47972_ _47972_/A _47973_/B sky130_fd_sc_hd__buf_2
X_43095_ _43085_/X _43086_/X _40729_/X _43094_/Y _43090_/X _43095_/Y
+ sky130_fd_sc_hd__o32ai_4
X_59958_ _62504_/A _62515_/A sky130_fd_sc_hd__buf_2
X_78792_ _82433_/Q _78792_/B _78793_/B sky130_fd_sc_hd__xnor2_4
X_49711_ _57692_/B _49687_/X _49710_/Y _49711_/Y sky130_fd_sc_hd__o21ai_4
X_46923_ _58997_/A _46908_/X _46922_/Y _46923_/Y sky130_fd_sc_hd__o21ai_4
X_42046_ _42046_/A _42046_/Y sky130_fd_sc_hd__inv_2
X_58909_ _58872_/A _86374_/Q _58909_/Y sky130_fd_sc_hd__nor2_4
X_77743_ _77743_/A _77742_/Y _77744_/B sky130_fd_sc_hd__xnor2_4
X_74955_ _74952_/Y _74954_/Y _74956_/B sky130_fd_sc_hd__xor2_4
X_70078_ _69910_/X _69912_/X _69994_/X _70078_/X sky130_fd_sc_hd__a21o_4
X_59889_ _59562_/B _59544_/A _59544_/B _59890_/C _60171_/B sky130_fd_sc_hd__nand4_4
X_49642_ _49625_/A _49642_/B _49629_/X _52857_/D _49642_/X sky130_fd_sc_hd__and4_4
X_73906_ _73902_/X _73905_/X _73857_/X _73910_/A sky130_fd_sc_hd__a21o_4
X_61920_ _61842_/A _61953_/B sky130_fd_sc_hd__buf_2
X_46854_ _46667_/A _46868_/C sky130_fd_sc_hd__buf_2
Xclkbuf_10_382_0_CLK clkbuf_9_191_0_CLK/X _85439_/CLK sky130_fd_sc_hd__clkbuf_1
X_77674_ _77674_/A _82123_/Q _77675_/A sky130_fd_sc_hd__nand2_4
X_74886_ _74887_/A _74887_/C _74887_/B _74888_/A sky130_fd_sc_hd__a21o_4
X_79413_ _84808_/Q _66415_/C _79415_/A sky130_fd_sc_hd__xor2_4
X_45805_ _62126_/D _61640_/A sky130_fd_sc_hd__buf_2
X_76625_ _76615_/Y _76616_/B _76624_/B _76625_/Y sky130_fd_sc_hd__o21ai_4
X_49573_ _49568_/Y _49570_/X _49572_/X _86363_/D sky130_fd_sc_hd__a21oi_4
X_61851_ _61823_/A _61823_/B _63459_/B _61788_/X _61851_/X sky130_fd_sc_hd__and4_4
X_73837_ _73838_/B _73838_/C _73836_/X _73837_/X sky130_fd_sc_hd__a21o_4
X_46785_ _46781_/Y _46751_/X _46784_/X _86704_/D sky130_fd_sc_hd__a21oi_4
X_43997_ _43994_/A _43998_/A sky130_fd_sc_hd__inv_2
X_48524_ _48516_/Y _48517_/X _48523_/X _86515_/D sky130_fd_sc_hd__a21oi_4
X_60802_ _78059_/A _60673_/X _60675_/Y _60801_/X _84564_/D sky130_fd_sc_hd__a2bb2oi_4
X_79344_ _79342_/X _79344_/B _79344_/Y sky130_fd_sc_hd__xnor2_4
X_45736_ _57179_/B _45736_/B _45736_/Y sky130_fd_sc_hd__nor2_4
X_64570_ _64564_/X _86145_/Q _64566_/X _64569_/X _64570_/X sky130_fd_sc_hd__a211o_4
X_76556_ _76531_/Y _76535_/B _76533_/Y _76557_/A sky130_fd_sc_hd__o21a_4
X_42948_ _42944_/X _42945_/X _41791_/X _68078_/B _42934_/X _42949_/A
+ sky130_fd_sc_hd__o32ai_4
X_61782_ _61782_/A _61776_/Y _61779_/Y _61781_/Y _61782_/Y sky130_fd_sc_hd__nand4_4
X_73768_ _73766_/X _73767_/Y _73720_/X _73768_/X sky130_fd_sc_hd__a21o_4
X_75507_ _75507_/A _75462_/X _75481_/X _75482_/Y _75508_/A sky130_fd_sc_hd__nand4_4
X_63521_ _58554_/A _63497_/X _61492_/A _63498_/X _63521_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_10_397_0_CLK clkbuf_9_198_0_CLK/X _82272_/CLK sky130_fd_sc_hd__clkbuf_1
X_48455_ _53663_/B _50440_/B sky130_fd_sc_hd__buf_2
X_60733_ _63410_/A _60714_/A _60732_/Y _60733_/Y sky130_fd_sc_hd__a21boi_4
X_72719_ _83178_/Q _72709_/X _72718_/X _72719_/X sky130_fd_sc_hd__a21o_4
X_79275_ _79292_/B _79275_/B _79275_/X sky130_fd_sc_hd__xor2_4
X_45667_ _45666_/Y _44975_/A _45667_/X sky130_fd_sc_hd__and2_4
X_76487_ _81657_/Q _76487_/Y sky130_fd_sc_hd__inv_2
X_42879_ _42874_/X _42875_/X _41606_/X _67248_/B _42858_/X _42879_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73699_ _73699_/A _73624_/X _73699_/Y sky130_fd_sc_hd__nor2_4
X_47406_ _81806_/Q _47407_/A sky130_fd_sc_hd__inv_2
X_66240_ _65880_/A _66240_/X sky130_fd_sc_hd__buf_2
X_78226_ _78226_/A _78226_/B _78226_/X sky130_fd_sc_hd__xor2_4
X_44618_ _44618_/A _44618_/X sky130_fd_sc_hd__buf_2
X_63452_ _61417_/B _63426_/X _63450_/X _63451_/X _63452_/X sky130_fd_sc_hd__a211o_4
X_75438_ _75436_/Y _75406_/Y _75437_/X _75438_/Y sky130_fd_sc_hd__o21ai_4
X_60664_ _60663_/Y _60671_/B sky130_fd_sc_hd__buf_2
X_48386_ _48372_/X _82367_/Q _48385_/Y _74375_/A sky130_fd_sc_hd__o21ai_4
X_45598_ _45595_/Y _45596_/X _45548_/X _45597_/Y _45598_/X sky130_fd_sc_hd__a211o_4
X_62403_ _62448_/A _63520_/B _62375_/C _62406_/C sky130_fd_sc_hd__nand3_4
X_47337_ _86645_/Q _47332_/X _47336_/Y _47337_/Y sky130_fd_sc_hd__o21ai_4
X_66171_ _64710_/A _66171_/B _66171_/X sky130_fd_sc_hd__and2_4
X_78157_ _78145_/A _82860_/D _78157_/Y sky130_fd_sc_hd__nand2_4
X_44549_ _44549_/A _44549_/X sky130_fd_sc_hd__buf_2
X_63383_ _63381_/Y _63284_/X _63382_/Y _84328_/D sky130_fd_sc_hd__a21oi_4
X_75369_ _75365_/Y _75345_/B _75368_/X _75369_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_320_0_CLK clkbuf_9_160_0_CLK/X _86655_/CLK sky130_fd_sc_hd__clkbuf_1
X_60595_ _60570_/B _60570_/C _60595_/C _60596_/B sky130_fd_sc_hd__nor3_4
X_65122_ _64851_/A _65122_/X sky130_fd_sc_hd__buf_2
X_77108_ _77113_/A _77112_/A _77107_/Y _77109_/B sky130_fd_sc_hd__a21boi_4
X_62334_ _61428_/X _59898_/A _62233_/C _62334_/D _62335_/D sky130_fd_sc_hd__nand4_4
Xclkbuf_10_950_0_CLK clkbuf_9_475_0_CLK/X _83153_/CLK sky130_fd_sc_hd__clkbuf_1
X_47268_ _54121_/B _52950_/B sky130_fd_sc_hd__buf_2
X_78088_ _78088_/A _78088_/B _78089_/A sky130_fd_sc_hd__nand2_4
X_49007_ _49007_/A _49006_/X _49007_/Y sky130_fd_sc_hd__nand2_4
X_46219_ _46217_/Y _46215_/B _46218_/Y _46220_/A sky130_fd_sc_hd__nand3_4
X_65053_ _65050_/X _65052_/X _64701_/X _65053_/X sky130_fd_sc_hd__a21o_4
X_69930_ _69791_/A _69929_/Y _69930_/Y sky130_fd_sc_hd__nor2_4
X_77039_ _77038_/X _77041_/B sky130_fd_sc_hd__inv_2
X_62265_ _62120_/A _62267_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_441_0_CLK clkbuf_9_441_0_CLK/A clkbuf_9_441_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_47199_ _47198_/X _47210_/A sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_15 _55686_/C _56175_/B sky130_fd_sc_hd__buf_2
X_64004_ _63733_/X _64071_/C sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_26 _50212_/A _41870_/B1 sky130_fd_sc_hd__buf_2
X_80050_ _80048_/X _80057_/B _80050_/Y sky130_fd_sc_hd__xnor2_4
X_61216_ _61215_/Y _61238_/C _61216_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_335_0_CLK clkbuf_9_167_0_CLK/X _84757_/CLK sky130_fd_sc_hd__clkbuf_1
X_69861_ _73320_/A _44299_/A _68933_/X _69860_/Y _69861_/X sky130_fd_sc_hd__a211o_4
X_62196_ _62196_/A _62196_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_965_0_CLK clkbuf_9_482_0_CLK/X _83594_/CLK sky130_fd_sc_hd__clkbuf_1
X_68812_ _80816_/D _68713_/X _68811_/X _68812_/X sky130_fd_sc_hd__a21bo_4
X_61147_ _61153_/A _64523_/D _64523_/B _61147_/Y sky130_fd_sc_hd__nand3_4
X_69792_ _73196_/A _69747_/X _68691_/X _69791_/Y _69792_/X sky130_fd_sc_hd__a211o_4
X_49909_ _72174_/B _49906_/X _49908_/Y _49909_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_456_0_CLK clkbuf_8_228_0_CLK/X clkbuf_9_456_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_68743_ _69067_/A _73921_/A _68743_/X sky130_fd_sc_hd__and2_4
X_65955_ _65916_/A _65970_/B _84166_/Q _65955_/X sky130_fd_sc_hd__and3_4
X_61078_ _59657_/A _61078_/B _60615_/A _61079_/A sky130_fd_sc_hd__nand3_4
X_52920_ _52892_/A _52920_/X sky130_fd_sc_hd__buf_2
X_64906_ _64883_/A _86262_/Q _64906_/X sky130_fd_sc_hd__and2_4
X_60029_ _62198_/B _60091_/A sky130_fd_sc_hd__buf_2
X_83740_ _86322_/CLK _83740_/D _47343_/A sky130_fd_sc_hd__dfxtp_4
X_80952_ _81211_/CLK _75393_/B _80952_/Q sky130_fd_sc_hd__dfxtp_4
X_68674_ _68670_/X _68673_/X _68390_/X _68674_/X sky130_fd_sc_hd__a21o_4
X_65886_ _65700_/X _65884_/Y _65885_/Y _65886_/Y sky130_fd_sc_hd__o21ai_4
X_67625_ _67270_/X _67625_/X sky130_fd_sc_hd__buf_2
X_52851_ _85743_/Q _52848_/X _52850_/Y _52851_/Y sky130_fd_sc_hd__o21ai_4
X_64837_ _64835_/X _83305_/Q _44171_/X _64836_/X _64837_/X sky130_fd_sc_hd__a211o_4
X_83671_ _83673_/CLK _70894_/Y _46786_/A sky130_fd_sc_hd__dfxtp_4
X_80883_ _81130_/CLK _75731_/B _80851_/D sky130_fd_sc_hd__dfxtp_4
X_85410_ _86655_/CLK _54613_/Y _85410_/Q sky130_fd_sc_hd__dfxtp_4
X_51802_ _53097_/A _53282_/A sky130_fd_sc_hd__buf_2
X_82622_ _82715_/CLK _79071_/B _82622_/Q sky130_fd_sc_hd__dfxtp_4
X_55570_ _55504_/Y _55536_/X _55552_/X _55570_/D _55570_/X sky130_fd_sc_hd__and4_4
X_67556_ _67460_/A _67556_/B _67556_/X sky130_fd_sc_hd__and2_4
X_86390_ _83676_/CLK _49426_/Y _58699_/B sky130_fd_sc_hd__dfxtp_4
X_52782_ _85755_/Q _52765_/X _52781_/Y _52782_/Y sky130_fd_sc_hd__o21ai_4
X_64768_ _64666_/X _86171_/Q _64766_/X _64767_/X _64768_/X sky130_fd_sc_hd__a211o_4
X_54521_ _54521_/A _54526_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_903_0_CLK clkbuf_9_451_0_CLK/X _88363_/CLK sky130_fd_sc_hd__clkbuf_1
X_66507_ _65339_/X _66521_/B _65344_/X _66507_/Y sky130_fd_sc_hd__nand3_4
X_85341_ _85375_/CLK _54984_/Y _85341_/Q sky130_fd_sc_hd__dfxtp_4
X_51733_ _85955_/Q _50220_/X _51732_/Y _51733_/Y sky130_fd_sc_hd__o21ai_4
X_63719_ _63717_/Y _63679_/X _63718_/Y _63719_/Y sky130_fd_sc_hd__a21oi_4
X_82553_ _82553_/CLK _82553_/D _82553_/Q sky130_fd_sc_hd__dfxtp_4
X_67487_ _67513_/A _87213_/Q _67487_/X sky130_fd_sc_hd__and2_4
X_64699_ _65836_/A _86045_/Q _64699_/X sky130_fd_sc_hd__and2_4
X_57240_ _44288_/X _56575_/X _45426_/A _57238_/X _85055_/D sky130_fd_sc_hd__a2bb2o_4
X_81504_ _81322_/CLK _81504_/D _76946_/B sky130_fd_sc_hd__dfxtp_4
X_69226_ _69222_/X _69226_/B _69226_/Y sky130_fd_sc_hd__nand2_4
X_88060_ _88060_/CLK _88060_/D _42041_/A sky130_fd_sc_hd__dfxtp_4
X_54452_ _85439_/Q _54431_/X _54451_/Y _54452_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_5_20_0_CLK clkbuf_4_10_1_CLK/X clkbuf_6_41_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_66438_ _66436_/Y _66437_/Y _63317_/X _66438_/X sky130_fd_sc_hd__a21o_4
X_85272_ _85241_/CLK _85272_/D _56216_/C sky130_fd_sc_hd__dfxtp_4
X_51664_ _51661_/Y _51639_/X _51663_/X _85969_/D sky130_fd_sc_hd__a21oi_4
X_82484_ _82580_/CLK _82484_/D _82860_/D sky130_fd_sc_hd__dfxtp_4
X_87011_ _87011_/CLK _87011_/D _87011_/Q sky130_fd_sc_hd__dfxtp_4
X_53403_ _53400_/Y _53382_/X _53402_/X _85640_/D sky130_fd_sc_hd__a21oi_4
X_84223_ _84223_/CLK _84223_/D _84223_/Q sky130_fd_sc_hd__dfxtp_4
X_50615_ _50624_/A _53834_/B _50615_/Y sky130_fd_sc_hd__nand2_4
X_81435_ _84064_/CLK _81467_/Q _76109_/B sky130_fd_sc_hd__dfxtp_4
X_57171_ _56995_/A _74342_/A sky130_fd_sc_hd__buf_2
X_69157_ _69152_/X _69155_/X _69156_/X _69157_/Y sky130_fd_sc_hd__a21oi_4
X_54383_ _85452_/Q _54376_/X _54382_/Y _54383_/Y sky130_fd_sc_hd__o21ai_4
X_66369_ _66318_/X _66415_/B _84136_/Q _66369_/X sky130_fd_sc_hd__and3_4
X_51595_ _51622_/A _51617_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_918_0_CLK clkbuf_9_459_0_CLK/X _83561_/CLK sky130_fd_sc_hd__clkbuf_1
X_56122_ _45369_/A _56123_/A sky130_fd_sc_hd__buf_2
X_68108_ _68088_/X _66671_/Y _68089_/X _68107_/Y _68108_/X sky130_fd_sc_hd__a211o_4
X_53334_ _53330_/A _53330_/B _53330_/C _52818_/D _53334_/X sky130_fd_sc_hd__and4_4
X_84154_ _82746_/CLK _84154_/D _66138_/A sky130_fd_sc_hd__dfxtp_4
X_50546_ _86180_/Q _50533_/X _50545_/Y _50546_/Y sky130_fd_sc_hd__o21ai_4
X_81366_ _83940_/CLK _76961_/Y _81366_/Q sky130_fd_sc_hd__dfxtp_4
X_69088_ _69088_/A _69088_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_7_0_CLK clkbuf_9_3_0_CLK/X _85279_/CLK sky130_fd_sc_hd__clkbuf_1
X_83105_ _83095_/CLK _74307_/X _83105_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_409_0_CLK clkbuf_9_409_0_CLK/A clkbuf_9_409_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_56053_ _56029_/X _56050_/X _56052_/Y _85305_/D sky130_fd_sc_hd__o21ai_4
X_80317_ _80306_/Y _80317_/B _80318_/A _80320_/A sky130_fd_sc_hd__nand3_4
X_68039_ _84044_/Q _67925_/X _68038_/X _84044_/D sky130_fd_sc_hd__a21bo_4
X_53265_ _51843_/A _53274_/B sky130_fd_sc_hd__buf_2
X_84085_ _84087_/CLK _67068_/X _84085_/Q sky130_fd_sc_hd__dfxtp_4
X_50477_ _50465_/X _48540_/B _50477_/Y sky130_fd_sc_hd__nand2_4
X_81297_ _81811_/CLK _76985_/X _81265_/D sky130_fd_sc_hd__dfxtp_4
X_55004_ _54927_/A _55026_/B sky130_fd_sc_hd__buf_2
X_52216_ _52220_/A _52216_/B _52216_/Y sky130_fd_sc_hd__nand2_4
X_71050_ _71055_/A _71073_/B _71055_/C _71050_/Y sky130_fd_sc_hd__nand3_4
X_87913_ _87188_/CLK _42340_/Y _87913_/Q sky130_fd_sc_hd__dfxtp_4
X_83036_ _85213_/CLK _74558_/Y _44989_/A sky130_fd_sc_hd__dfxtp_4
X_80248_ _80243_/X _80247_/Y _80248_/X sky130_fd_sc_hd__xor2_4
X_53196_ _53211_/A _53181_/B _53195_/X _53196_/D _53196_/X sky130_fd_sc_hd__and4_4
X_70001_ _70001_/A _70001_/X sky130_fd_sc_hd__buf_2
X_59812_ _59758_/X _59654_/X _59811_/Y _59812_/Y sky130_fd_sc_hd__nand3_4
X_52147_ _52144_/Y _52145_/X _52146_/X _85880_/D sky130_fd_sc_hd__a21oi_4
X_87844_ _87588_/CLK _87844_/D _42499_/A sky130_fd_sc_hd__dfxtp_4
X_80179_ _80151_/Y _80169_/B _80164_/Y _80167_/Y _80179_/X sky130_fd_sc_hd__o22a_4
X_59743_ _59608_/A _59743_/B _59743_/Y sky130_fd_sc_hd__nor2_4
X_52078_ _85893_/Q _52075_/X _52077_/Y _52078_/Y sky130_fd_sc_hd__o21ai_4
X_56955_ _56600_/X _56952_/X _56954_/Y _85115_/D sky130_fd_sc_hd__a21oi_4
X_87775_ _87789_/CLK _87775_/D _69409_/B sky130_fd_sc_hd__dfxtp_4
X_84987_ _84991_/CLK _57522_/Y _84987_/Q sky130_fd_sc_hd__dfxtp_4
X_43920_ _41393_/X _43907_/X _67810_/B _43908_/X _43920_/X sky130_fd_sc_hd__a2bb2o_4
X_51029_ _51029_/A _51029_/B _51029_/C _52720_/D _51029_/X sky130_fd_sc_hd__and4_4
X_55906_ _85209_/Q _44106_/C _55627_/X _55905_/X _55906_/X sky130_fd_sc_hd__a211o_4
X_74740_ _71012_/B _74740_/B _71507_/B _74739_/Y _74740_/Y sky130_fd_sc_hd__nand4_4
X_86726_ _86119_/CLK _86726_/D _86726_/Q sky130_fd_sc_hd__dfxtp_4
X_71952_ _71942_/Y _83316_/Q _71951_/Y _83316_/D sky130_fd_sc_hd__a21o_4
X_59674_ _60036_/A _66262_/A sky130_fd_sc_hd__buf_2
X_83938_ _83932_/CLK _69244_/X _83938_/Q sky130_fd_sc_hd__dfxtp_4
X_56886_ _56880_/X _56886_/B _56886_/Y sky130_fd_sc_hd__xnor2_4
Xclkbuf_6_9_0_CLK clkbuf_6_9_0_CLK/A clkbuf_6_9_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_58625_ _58858_/A _58625_/X sky130_fd_sc_hd__buf_2
X_70903_ _70903_/A _70903_/B _70899_/C _70899_/D _70903_/Y sky130_fd_sc_hd__nand4_4
X_55837_ _85264_/Q _55475_/X _44048_/X _55836_/X _55837_/X sky130_fd_sc_hd__a211o_4
X_43851_ _41203_/X _43842_/X _68793_/B _43843_/X _87234_/D sky130_fd_sc_hd__a2bb2o_4
X_74671_ _74673_/A _56752_/A _74670_/Y _74672_/A sky130_fd_sc_hd__o21ai_4
X_86657_ _85727_/CLK _86657_/D _57698_/A sky130_fd_sc_hd__dfxtp_4
X_71883_ _71883_/A _71883_/B _71873_/X _71883_/D _71883_/Y sky130_fd_sc_hd__nor4_4
X_83869_ _82553_/CLK _70028_/X _82549_/D sky130_fd_sc_hd__dfxtp_4
X_76410_ _76410_/A _81568_/Q _76410_/Y sky130_fd_sc_hd__nand2_4
X_42802_ _42745_/A _42802_/X sky130_fd_sc_hd__buf_2
X_73622_ _73620_/X _73621_/Y _73546_/X _73622_/X sky130_fd_sc_hd__a21o_4
X_85608_ _85601_/CLK _85608_/D _85608_/Q sky130_fd_sc_hd__dfxtp_4
X_46570_ _46531_/A _54079_/B _46570_/Y sky130_fd_sc_hd__nand2_4
X_70834_ _51744_/B _70831_/X _70833_/Y _83689_/D sky130_fd_sc_hd__o21ai_4
X_58556_ _84819_/Q _58557_/A sky130_fd_sc_hd__inv_2
X_77390_ _77390_/A _82189_/D _77390_/X sky130_fd_sc_hd__xor2_4
X_43782_ _43774_/X _43781_/X _41009_/X _69318_/B _43776_/X _43782_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55768_ _55765_/X _55767_/X _44108_/X _55768_/X sky130_fd_sc_hd__a21o_4
X_86588_ _86237_/CLK _47896_/Y _65977_/B sky130_fd_sc_hd__dfxtp_4
X_40994_ _40994_/A _40994_/X sky130_fd_sc_hd__buf_2
X_45521_ _57254_/B _45490_/B _45521_/Y sky130_fd_sc_hd__nor2_4
X_57507_ _47871_/A _49317_/X _46603_/X _57507_/X sky130_fd_sc_hd__and3_4
X_76341_ _76324_/Y _76339_/X _76340_/X _76342_/B sky130_fd_sc_hd__a21boi_4
X_42733_ _42721_/X _42723_/X _41209_/X _87745_/Q _42732_/X _42734_/A
+ sky130_fd_sc_hd__o32ai_4
X_88327_ _88327_/CLK _40828_/Y _69725_/B sky130_fd_sc_hd__dfxtp_4
X_54719_ _85390_/Q _54703_/X _54718_/Y _54719_/Y sky130_fd_sc_hd__o21ai_4
X_73553_ _68361_/Y _73319_/X _73551_/X _73552_/Y _73553_/X sky130_fd_sc_hd__a211o_4
X_85539_ _85826_/CLK _85539_/D _85539_/Q sky130_fd_sc_hd__dfxtp_4
X_70765_ _70772_/A _70766_/C sky130_fd_sc_hd__buf_2
X_58487_ _58487_/A _58502_/B _58487_/Y sky130_fd_sc_hd__nor2_4
X_55699_ _74541_/C _55690_/X _44102_/X _55698_/X _55700_/B sky130_fd_sc_hd__a211o_4
X_48240_ _48237_/Y _48226_/X _48239_/Y _86550_/D sky130_fd_sc_hd__a21boi_4
X_72504_ _72516_/B _72535_/A sky130_fd_sc_hd__inv_2
X_79060_ _79058_/A _82749_/Q _79058_/B _79060_/Y sky130_fd_sc_hd__nand3_4
X_57438_ _57408_/X _57436_/X _57437_/Y _57439_/A sky130_fd_sc_hd__o21ai_4
X_45452_ _45452_/A _45452_/X sky130_fd_sc_hd__buf_2
X_76272_ _76268_/Y _76211_/Y _76271_/X _76272_/Y sky130_fd_sc_hd__o21ai_4
X_88258_ _87103_/CLK _41204_/X _68796_/B sky130_fd_sc_hd__dfxtp_4
X_42664_ _42663_/Y _42664_/Y sky130_fd_sc_hd__inv_2
X_73484_ _73484_/A _72892_/B _73484_/Y sky130_fd_sc_hd__nor2_4
X_70696_ _70758_/A _70696_/B _70758_/B _70935_/A sky130_fd_sc_hd__nor3_4
X_78011_ _78011_/A _78011_/Y sky130_fd_sc_hd__inv_2
X_44403_ _41511_/X _44394_/X _87125_/Q _44395_/X _44403_/X sky130_fd_sc_hd__a2bb2o_4
X_87209_ _87210_/CLK _43901_/Y _87209_/Q sky130_fd_sc_hd__dfxtp_4
X_75223_ _75214_/B _81068_/Q _75222_/Y _75223_/Y sky130_fd_sc_hd__a21boi_4
X_41615_ _41533_/X _82308_/Q _41614_/X _41615_/X sky130_fd_sc_hd__o21a_4
X_48171_ _48186_/A _48171_/X sky130_fd_sc_hd__buf_2
X_72435_ _83255_/Q _72381_/X _72429_/X _72434_/X _83255_/D sky130_fd_sc_hd__a2bb2oi_4
X_45383_ _62629_/A _61692_/B sky130_fd_sc_hd__buf_2
X_57369_ _57244_/X _45870_/Y _57369_/Y sky130_fd_sc_hd__nand2_4
X_88189_ _87116_/CLK _41576_/Y _67100_/B sky130_fd_sc_hd__dfxtp_4
X_42595_ _42590_/X _42592_/X _40866_/X _87808_/Q _42580_/X _42596_/A
+ sky130_fd_sc_hd__o32ai_4
X_47122_ _47118_/Y _47081_/X _47121_/X _47122_/Y sky130_fd_sc_hd__a21oi_4
X_59108_ _59085_/X _86072_/Q _59107_/X _59108_/Y sky130_fd_sc_hd__o21ai_4
X_44334_ _44333_/Y _87162_/D sky130_fd_sc_hd__inv_2
X_75154_ _75157_/B _75154_/Y sky130_fd_sc_hd__inv_2
X_41546_ _41540_/X _41541_/X _41545_/X _66966_/B _41537_/X _41547_/A
+ sky130_fd_sc_hd__o32ai_4
X_60380_ _59775_/X _60380_/B _60392_/A _60392_/C _60381_/A sky130_fd_sc_hd__and4_4
X_72366_ _72366_/A _72366_/B _72366_/Y sky130_fd_sc_hd__nor2_4
X_74105_ _74080_/X _86218_/Q _74103_/X _74104_/X _74105_/X sky130_fd_sc_hd__a211o_4
X_47053_ _47053_/A _52829_/B sky130_fd_sc_hd__buf_2
X_71317_ _48073_/B _71289_/Y _71316_/Y _83538_/D sky130_fd_sc_hd__o21ai_4
X_59039_ _59001_/X _86078_/Q _59038_/X _59039_/Y sky130_fd_sc_hd__o21ai_4
X_44265_ _65880_/A _44261_/X _57837_/A _44265_/D _44265_/Y sky130_fd_sc_hd__nor4_4
X_79962_ _79960_/Y _79963_/A sky130_fd_sc_hd__inv_2
X_75085_ _75082_/X _75085_/B _75102_/B _75102_/A sky130_fd_sc_hd__nand3_4
X_41477_ _81181_/Q _41459_/B _41477_/X sky130_fd_sc_hd__or2_4
X_72297_ _72270_/X _72294_/Y _72295_/Y _72296_/X _72274_/X _72297_/X
+ sky130_fd_sc_hd__o32a_4
X_46004_ _40484_/Y _45974_/X _67023_/B _45976_/X _86819_/D sky130_fd_sc_hd__a2bb2o_4
X_43216_ _43180_/A _43216_/X sky130_fd_sc_hd__buf_2
X_62050_ _61722_/A _62050_/X sky130_fd_sc_hd__buf_2
X_74036_ _88351_/Q _72899_/X _73898_/X _74036_/X sky130_fd_sc_hd__o21a_4
X_78913_ _78900_/A _78908_/A _78913_/X sky130_fd_sc_hd__and2_4
X_40428_ _40428_/A _40428_/Y sky130_fd_sc_hd__inv_2
X_71248_ _71252_/A _71223_/B _71248_/C _71248_/Y sky130_fd_sc_hd__nand3_4
X_44196_ _44196_/A _44196_/B _72899_/A _44196_/D _44196_/X sky130_fd_sc_hd__and4_4
X_79893_ _79547_/A _79546_/Y _79893_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_2_1_1_CLK clkbuf_2_1_0_CLK/X clkbuf_2_1_1_CLK/X sky130_fd_sc_hd__clkbuf_1
X_61001_ _60969_/X _61000_/X _84543_/Q _61001_/X sky130_fd_sc_hd__or3_4
X_43147_ _43146_/X _43110_/X _40831_/X _73108_/A _43121_/X _43147_/Y
+ sky130_fd_sc_hd__o32ai_4
X_78844_ _78874_/A _78854_/B _78845_/B sky130_fd_sc_hd__xor2_4
X_40359_ _44587_/A _44528_/A sky130_fd_sc_hd__buf_2
X_71179_ _52158_/B _71165_/X _71178_/Y _71179_/Y sky130_fd_sc_hd__o21ai_4
X_47955_ _47955_/A _47963_/B _47955_/X sky130_fd_sc_hd__or2_4
X_43078_ _87584_/Q _43078_/Y sky130_fd_sc_hd__inv_2
X_78775_ _82816_/Q _78775_/Y sky130_fd_sc_hd__inv_2
X_75987_ _81515_/Q _81739_/D _75987_/X sky130_fd_sc_hd__xor2_4
X_46906_ _46868_/A _46896_/B _46926_/C _52742_/D _46906_/X sky130_fd_sc_hd__and4_4
X_42029_ _42028_/X _42024_/X _40861_/X _73225_/A _42025_/X _42029_/Y
+ sky130_fd_sc_hd__o32ai_4
X_65740_ _64599_/X _83061_/Q _65015_/X _65739_/X _65740_/X sky130_fd_sc_hd__a211o_4
X_77726_ _82258_/Q _77732_/B _78044_/A sky130_fd_sc_hd__xnor2_4
X_62952_ _63306_/A _62988_/B sky130_fd_sc_hd__buf_2
X_74938_ _74933_/Y _74942_/A _74937_/Y _74939_/B sky130_fd_sc_hd__a21boi_4
X_47886_ _47886_/A _47886_/X sky130_fd_sc_hd__buf_2
X_61903_ _59684_/X _61949_/B sky130_fd_sc_hd__buf_2
X_49625_ _49625_/A _49614_/X _49615_/C _52841_/D _49625_/X sky130_fd_sc_hd__and4_4
X_46837_ _54395_/D _52704_/D sky130_fd_sc_hd__buf_2
X_65671_ _65638_/X _85585_/Q _65669_/X _65670_/X _65671_/X sky130_fd_sc_hd__a211o_4
X_77657_ _77629_/Y _77633_/B _77632_/A _77657_/X sky130_fd_sc_hd__o21a_4
X_62883_ _62881_/X _62838_/X _62882_/Y _84374_/D sky130_fd_sc_hd__a21oi_4
X_74869_ _81126_/D _74869_/B _74897_/A sky130_fd_sc_hd__xor2_4
X_67410_ _67407_/X _67409_/X _67383_/X _67410_/X sky130_fd_sc_hd__a21o_4
X_64622_ _64577_/X _86752_/Q _64579_/X _64621_/X _64622_/X sky130_fd_sc_hd__a211o_4
X_76608_ _76608_/A _76603_/X _76611_/A sky130_fd_sc_hd__nand2_4
X_49556_ _49561_/A _49537_/B _49548_/X _52771_/D _49556_/X sky130_fd_sc_hd__and4_4
X_61834_ _61823_/X _61828_/X _61833_/Y _84915_/Q _61815_/X _61834_/Y
+ sky130_fd_sc_hd__o32ai_4
X_68390_ _69678_/A _68390_/X sky130_fd_sc_hd__buf_2
X_46768_ _46720_/A _46806_/A sky130_fd_sc_hd__buf_2
X_77588_ _77584_/X _77585_/Y _77587_/Y _77590_/A sky130_fd_sc_hd__a21o_4
X_48507_ _81780_/Q _48508_/A sky130_fd_sc_hd__inv_2
X_67341_ _67222_/A _67342_/A sky130_fd_sc_hd__buf_2
X_79327_ _79320_/X _79322_/B _79327_/Y sky130_fd_sc_hd__nand2_4
X_45719_ _45719_/A _45719_/Y sky130_fd_sc_hd__inv_2
X_64553_ _64474_/X _64525_/B _84882_/Q _64553_/Y sky130_fd_sc_hd__nand3_4
X_76539_ _76535_/X _76540_/C _76540_/B _76541_/A sky130_fd_sc_hd__a21o_4
X_61765_ _61762_/X _61765_/B _61765_/C _61748_/X _61766_/D sky130_fd_sc_hd__nand4_4
X_49487_ _49434_/A _49487_/X sky130_fd_sc_hd__buf_2
X_46699_ _46695_/Y _46654_/X _46698_/X _86713_/D sky130_fd_sc_hd__a21oi_4
X_63504_ _63443_/A _63514_/C sky130_fd_sc_hd__buf_2
X_60716_ _60715_/X _60752_/B sky130_fd_sc_hd__buf_2
X_48438_ _48642_/A _48438_/B _48438_/Y sky130_fd_sc_hd__nand2_4
X_79258_ _84793_/Q _66490_/C _79258_/X sky130_fd_sc_hd__xor2_4
X_67272_ _67248_/A _87670_/Q _67272_/X sky130_fd_sc_hd__and2_4
X_64484_ _64474_/X _61169_/X _62097_/X _64484_/Y sky130_fd_sc_hd__nand3_4
X_61696_ _84866_/Q _61321_/Y _61697_/A sky130_fd_sc_hd__or2_4
X_69011_ _69011_/A _69011_/B _69011_/X sky130_fd_sc_hd__and2_4
X_66223_ _66053_/X _85611_/Q _66096_/X _66222_/X _66223_/X sky130_fd_sc_hd__a211o_4
X_78209_ _78209_/A _78208_/X _78210_/B sky130_fd_sc_hd__nand2_4
X_63435_ _63448_/A _59501_/X _63410_/C _63410_/D _63435_/X sky130_fd_sc_hd__and4_4
X_48369_ _48392_/A _48368_/X _48369_/Y sky130_fd_sc_hd__nand2_4
X_60647_ _60820_/B _60646_/Y _59787_/X _60647_/Y sky130_fd_sc_hd__o21ai_4
X_79189_ _79189_/A _79189_/B _79189_/Y sky130_fd_sc_hd__nor2_4
X_50400_ _53511_/A _50430_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_41_0_CLK clkbuf_9_20_0_CLK/X _83095_/CLK sky130_fd_sc_hd__clkbuf_1
X_81220_ _85317_/CLK _81028_/Q _81220_/Q sky130_fd_sc_hd__dfxtp_4
X_66154_ _64589_/X _86224_/Q _45922_/X _66153_/X _66154_/X sky130_fd_sc_hd__a211o_4
X_51380_ _51367_/X _51380_/B _51380_/X sky130_fd_sc_hd__and2_4
X_63366_ _63364_/Y _63284_/X _63365_/Y _63366_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_380_0_CLK clkbuf_8_190_0_CLK/X clkbuf_9_380_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_60578_ _60515_/B _60476_/C _63280_/C _60578_/Y sky130_fd_sc_hd__nand3_4
X_65105_ _65002_/A _65105_/B _65105_/X sky130_fd_sc_hd__and2_4
X_50331_ _48287_/A _50331_/B _50247_/X _50331_/X sky130_fd_sc_hd__and3_4
X_81151_ _82327_/CLK _75062_/A _40579_/A sky130_fd_sc_hd__dfxtp_4
X_62317_ _61421_/A _62631_/B _62631_/C _62332_/D _62317_/Y sky130_fd_sc_hd__nand4_4
X_66085_ _65733_/X _85621_/Q _65734_/X _66084_/X _66085_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_274_0_CLK clkbuf_9_137_0_CLK/X _83414_/CLK sky130_fd_sc_hd__clkbuf_1
X_63297_ _79245_/A _63258_/X _63296_/Y _84336_/D sky130_fd_sc_hd__a21o_4
X_80102_ _60067_/C _80102_/B _80108_/B sky130_fd_sc_hd__xor2_4
X_53050_ _53040_/X _53050_/B _53050_/Y sky130_fd_sc_hd__nand2_4
X_65036_ _64679_/A _65036_/X sky130_fd_sc_hd__buf_2
X_69913_ _69910_/X _69912_/X _69742_/X _69913_/Y sky130_fd_sc_hd__a21oi_4
X_50262_ _50230_/A _48207_/X _50262_/Y sky130_fd_sc_hd__nand2_4
X_62248_ _61358_/A _62247_/X _62576_/C _62560_/D _62251_/B sky130_fd_sc_hd__nand4_4
X_81082_ _81082_/CLK _75637_/A _81082_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_56_0_CLK clkbuf_9_28_0_CLK/X _85075_/CLK sky130_fd_sc_hd__clkbuf_1
X_52001_ _52027_/A _47969_/B _52001_/Y sky130_fd_sc_hd__nand2_4
X_80033_ _80019_/Y _80016_/Y _80033_/X sky130_fd_sc_hd__and2_4
X_84910_ _84714_/CLK _58199_/Y _84910_/Q sky130_fd_sc_hd__dfxtp_4
X_69844_ _69840_/X _69843_/X _69844_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_395_0_CLK clkbuf_9_395_0_CLK/A clkbuf_9_395_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_50193_ _51242_/A _53919_/B _50193_/X sky130_fd_sc_hd__and2_4
X_85890_ _85888_/CLK _85890_/D _85890_/Q sky130_fd_sc_hd__dfxtp_4
X_62179_ _62851_/A _62179_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_202_0_CLK clkbuf_8_203_0_CLK/A clkbuf_8_202_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_289_0_CLK clkbuf_9_144_0_CLK/X _84727_/CLK sky130_fd_sc_hd__clkbuf_1
X_84841_ _84841_/CLK _84841_/D _84841_/Q sky130_fd_sc_hd__dfxtp_4
X_69775_ _83898_/Q _69763_/X _69774_/X _69775_/X sky130_fd_sc_hd__a21bo_4
X_66987_ _66983_/X _66986_/X _66964_/X _66987_/X sky130_fd_sc_hd__a21o_4
X_56740_ _56735_/X _56740_/X sky130_fd_sc_hd__buf_2
X_68726_ _44148_/A _69735_/A sky130_fd_sc_hd__buf_2
X_87560_ _87820_/CLK _87560_/D _43141_/A sky130_fd_sc_hd__dfxtp_4
X_53952_ _85535_/Q _53921_/X _53951_/Y _53952_/Y sky130_fd_sc_hd__o21ai_4
X_65938_ _65933_/X _65936_/X _65937_/X _65938_/X sky130_fd_sc_hd__a21o_4
X_84772_ _86686_/CLK _84772_/D _84772_/Q sky130_fd_sc_hd__dfxtp_4
X_81984_ _81975_/CLK _83912_/Q _81984_/Q sky130_fd_sc_hd__dfxtp_4
X_86511_ _86500_/CLK _86511_/D _86511_/Q sky130_fd_sc_hd__dfxtp_4
X_52903_ _52630_/A _52903_/X sky130_fd_sc_hd__buf_2
X_83723_ _85372_/CLK _83723_/D _47505_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_217_0_CLK clkbuf_8_217_0_CLK/A clkbuf_9_435_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_56671_ _56852_/A _56671_/X sky130_fd_sc_hd__buf_2
X_80935_ _81061_/CLK _75138_/B _74879_/A sky130_fd_sc_hd__dfxtp_4
X_68657_ _69014_/A _68735_/A sky130_fd_sc_hd__buf_2
X_87491_ _87749_/CLK _43299_/X _87491_/Q sky130_fd_sc_hd__dfxtp_4
X_53883_ _53763_/A _53888_/C sky130_fd_sc_hd__buf_2
X_65869_ _65789_/X _65359_/Y _65868_/Y _65869_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_212_0_CLK clkbuf_9_106_0_CLK/X _84649_/CLK sky130_fd_sc_hd__clkbuf_1
X_58410_ _58406_/X _83368_/Q _58409_/Y _84856_/D sky130_fd_sc_hd__o21a_4
X_55622_ _55691_/A _55622_/B _55622_/X sky130_fd_sc_hd__and2_4
X_67608_ _67539_/X _67608_/B _67608_/X sky130_fd_sc_hd__and2_4
X_86442_ _86154_/CLK _86442_/D _86442_/Q sky130_fd_sc_hd__dfxtp_4
X_52834_ _85746_/Q _52821_/X _52833_/Y _52834_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_842_0_CLK clkbuf_9_421_0_CLK/X _84161_/CLK sky130_fd_sc_hd__clkbuf_1
X_59390_ _84744_/Q _59390_/Y sky130_fd_sc_hd__inv_2
X_83654_ _85822_/CLK _70948_/Y _83654_/Q sky130_fd_sc_hd__dfxtp_4
X_80866_ _80818_/CLK _75571_/B _80834_/D sky130_fd_sc_hd__dfxtp_4
X_68588_ _68588_/A _68588_/Y sky130_fd_sc_hd__inv_2
X_58341_ _58341_/A _58341_/X sky130_fd_sc_hd__buf_2
X_82605_ _82604_/CLK _78909_/B _82605_/Q sky130_fd_sc_hd__dfxtp_4
X_55553_ _55524_/A _45500_/Y _55553_/Y sky130_fd_sc_hd__nor2_4
X_67539_ _67062_/X _67539_/X sky130_fd_sc_hd__buf_2
X_86373_ _83660_/CLK _86373_/D _58920_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_333_0_CLK clkbuf_8_166_0_CLK/X clkbuf_9_333_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_52765_ _52684_/A _52765_/X sky130_fd_sc_hd__buf_2
X_83585_ _83584_/CLK _71169_/Y _48444_/A sky130_fd_sc_hd__dfxtp_4
X_80797_ _81111_/CLK _75886_/Y _75491_/B sky130_fd_sc_hd__dfxtp_4
X_88112_ _87070_/CLK _41892_/Y _88112_/Q sky130_fd_sc_hd__dfxtp_4
X_54504_ _54501_/Y _54502_/X _54503_/X _54504_/Y sky130_fd_sc_hd__a21oi_4
X_85324_ _85354_/CLK _85324_/D _85324_/Q sky130_fd_sc_hd__dfxtp_4
X_51716_ _51713_/Y _51693_/X _51715_/X _51716_/Y sky130_fd_sc_hd__a21oi_4
X_70550_ _71698_/A _70549_/X _70538_/X _70550_/D _70550_/Y sky130_fd_sc_hd__nor4_4
X_58272_ _84891_/Q _58274_/A sky130_fd_sc_hd__inv_2
X_82536_ _82536_/CLK _82536_/D _82536_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_227_0_CLK clkbuf_9_113_0_CLK/X _80676_/CLK sky130_fd_sc_hd__clkbuf_1
X_55484_ _55453_/X _55483_/Y _55484_/Y sky130_fd_sc_hd__nor2_4
X_52696_ _52706_/A _52696_/B _52696_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_857_0_CLK clkbuf_9_428_0_CLK/X _85514_/CLK sky130_fd_sc_hd__clkbuf_1
X_57223_ _57222_/Y _45904_/X _46237_/A _57223_/D _57223_/X sky130_fd_sc_hd__and4_4
X_69209_ _69073_/A _69209_/B _69209_/X sky130_fd_sc_hd__and2_4
X_88043_ _88044_/CLK _42085_/Y _88043_/Q sky130_fd_sc_hd__dfxtp_4
X_54435_ _54435_/A _54417_/B _54429_/C _54435_/D _54435_/X sky130_fd_sc_hd__and4_4
X_85255_ _85221_/CLK _85255_/D _85255_/Q sky130_fd_sc_hd__dfxtp_4
X_51647_ _51621_/A _51647_/X sky130_fd_sc_hd__buf_2
X_70481_ _70466_/Y _83765_/Q _70480_/X _70481_/X sky130_fd_sc_hd__a21o_4
X_82467_ _82924_/CLK _82467_/D _82467_/Q sky130_fd_sc_hd__dfxtp_4
X_41400_ _41490_/A _41400_/X sky130_fd_sc_hd__buf_2
X_72220_ _72220_/A _72220_/B _72220_/Y sky130_fd_sc_hd__nor2_4
X_84206_ _85315_/CLK _84206_/D _84206_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_348_0_CLK clkbuf_8_174_0_CLK/X clkbuf_9_348_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_81418_ _81532_/CLK _81418_/D _75972_/B sky130_fd_sc_hd__dfxtp_4
X_57154_ _44256_/A _57152_/X _57153_/Y _85071_/D sky130_fd_sc_hd__o21ai_4
X_42380_ _42379_/Y _87893_/D sky130_fd_sc_hd__inv_2
X_54366_ _54366_/A _54366_/X sky130_fd_sc_hd__buf_2
X_85186_ _85186_/CLK _56459_/Y _56458_/C sky130_fd_sc_hd__dfxtp_4
X_51578_ _85984_/Q _51566_/X _51577_/Y _51578_/Y sky130_fd_sc_hd__o21ai_4
X_82398_ _82965_/CLK _82206_/Q _82398_/Q sky130_fd_sc_hd__dfxtp_4
X_56105_ _56131_/A _56115_/B _55826_/B _56105_/Y sky130_fd_sc_hd__nand3_4
X_41331_ _41242_/X _41679_/A _41330_/X _41331_/X sky130_fd_sc_hd__o21a_4
X_53317_ _53315_/Y _53301_/X _53316_/X _53317_/Y sky130_fd_sc_hd__a21oi_4
X_72151_ _83278_/Q _72151_/Y sky130_fd_sc_hd__inv_2
X_84137_ _82177_/CLK _84137_/D _66364_/C sky130_fd_sc_hd__dfxtp_4
X_50529_ _86183_/Q _50506_/X _50528_/Y _50529_/Y sky130_fd_sc_hd__o21ai_4
X_57085_ _56989_/A _57083_/X _57084_/Y _57085_/X sky130_fd_sc_hd__o21a_4
X_81349_ _84105_/CLK _81349_/D _81349_/Q sky130_fd_sc_hd__dfxtp_4
X_54297_ _85468_/Q _54294_/X _54296_/Y _54297_/Y sky130_fd_sc_hd__o21ai_4
X_71102_ _71101_/X _71055_/B _71099_/C _71102_/Y sky130_fd_sc_hd__nand3_4
X_44050_ _44049_/X _44051_/A sky130_fd_sc_hd__buf_2
X_56036_ _45765_/A _56052_/B sky130_fd_sc_hd__buf_2
X_53248_ _53302_/A _53266_/C sky130_fd_sc_hd__buf_2
X_41262_ _41159_/A _40737_/A _41262_/X sky130_fd_sc_hd__or2_4
X_72082_ _83288_/Q _72051_/X _72081_/Y _72082_/Y sky130_fd_sc_hd__o21ai_4
X_84068_ _82648_/CLK _84068_/D _81500_/D sky130_fd_sc_hd__dfxtp_4
X_43001_ _43001_/A _43001_/Y sky130_fd_sc_hd__inv_2
X_71033_ _71178_/A _71030_/B _71030_/C _71018_/D _71033_/Y sky130_fd_sc_hd__nand4_4
X_75910_ _61203_/C _62816_/C _75910_/X sky130_fd_sc_hd__xor2_4
X_83019_ _80670_/CLK _74604_/Y _45244_/A sky130_fd_sc_hd__dfxtp_4
X_41193_ _41192_/X _41193_/X sky130_fd_sc_hd__buf_2
X_53179_ _53187_/A _53179_/B _53179_/Y sky130_fd_sc_hd__nand2_4
X_76890_ _76889_/X _81468_/D sky130_fd_sc_hd__buf_2
X_75841_ _75841_/A _75841_/Y sky130_fd_sc_hd__inv_2
X_87827_ _87826_/CLK _87827_/D _72728_/A sky130_fd_sc_hd__dfxtp_4
X_57987_ _57926_/X _85998_/Q _57986_/X _57987_/Y sky130_fd_sc_hd__o21ai_4
X_47740_ _47736_/Y _47698_/X _47739_/X _47740_/Y sky130_fd_sc_hd__a21oi_4
X_59726_ _66064_/A _66377_/A sky130_fd_sc_hd__buf_2
X_78560_ _78560_/A _78560_/B _78563_/A sky130_fd_sc_hd__nand2_4
X_44952_ _44950_/Y _45590_/B _44952_/X sky130_fd_sc_hd__and2_4
X_56938_ _72771_/A _72732_/B sky130_fd_sc_hd__buf_2
X_75772_ _75759_/A _75766_/A _75772_/X sky130_fd_sc_hd__and2_4
X_87758_ _87758_/CLK _42709_/Y _87758_/Q sky130_fd_sc_hd__dfxtp_4
X_72984_ _72973_/Y _72975_/Y _72983_/X _72984_/Y sky130_fd_sc_hd__o21ai_4
X_77511_ _77511_/A _77510_/Y _77512_/B sky130_fd_sc_hd__and2_4
X_43903_ _43895_/X _43902_/X _41347_/X _67596_/B _43897_/X _43903_/Y
+ sky130_fd_sc_hd__o32ai_4
X_86709_ _86711_/CLK _86709_/D _58722_/A sky130_fd_sc_hd__dfxtp_4
X_74723_ _70576_/X _74723_/X sky130_fd_sc_hd__buf_2
X_47671_ _72302_/A _47666_/X _47670_/Y _47671_/Y sky130_fd_sc_hd__o21ai_4
X_71935_ _71170_/A _74518_/B sky130_fd_sc_hd__buf_2
X_59657_ _59657_/A _60353_/B sky130_fd_sc_hd__buf_2
X_78491_ _78487_/Y _78488_/Y _78490_/Y _78491_/X sky130_fd_sc_hd__or3_4
X_44883_ _80671_/Q _45389_/A sky130_fd_sc_hd__inv_2
X_56869_ _56868_/X _56869_/Y sky130_fd_sc_hd__inv_2
X_87689_ _87888_/CLK _87689_/D _66817_/B sky130_fd_sc_hd__dfxtp_4
X_49410_ _49410_/A _46701_/X _49410_/Y sky130_fd_sc_hd__nand2_4
X_46622_ _46719_/A _46622_/X sky130_fd_sc_hd__buf_2
X_58608_ _58571_/X _85790_/Q _58594_/X _58608_/X sky130_fd_sc_hd__o21a_4
X_77442_ _77422_/Y _77423_/Y _77424_/Y _77442_/X sky130_fd_sc_hd__o21a_4
X_43834_ _41151_/X _43832_/X _68546_/B _43833_/X _43834_/X sky130_fd_sc_hd__a2bb2o_4
X_74654_ _45951_/Y _56638_/X _45604_/A _74645_/X _74654_/X sky130_fd_sc_hd__a2bb2o_4
X_71866_ _71847_/Y _83347_/Q _71865_/Y _83347_/D sky130_fd_sc_hd__a21o_4
X_59588_ _59662_/B _59633_/A _59634_/B _59588_/Y sky130_fd_sc_hd__o21ai_4
X_49341_ _65310_/B _49334_/X _49340_/Y _49341_/Y sky130_fd_sc_hd__o21ai_4
X_73605_ _73355_/A _73605_/X sky130_fd_sc_hd__buf_2
X_70817_ _47184_/X _70802_/X _70816_/Y _83693_/D sky130_fd_sc_hd__o21ai_4
X_46553_ _46548_/Y _46523_/X _46552_/Y _86727_/D sky130_fd_sc_hd__a21boi_4
X_58539_ _84824_/Q _58541_/A sky130_fd_sc_hd__inv_2
X_77373_ _77351_/B _77371_/Y _77372_/Y _77374_/B sky130_fd_sc_hd__a21oi_4
X_43765_ _43005_/X _43760_/X _40972_/X _69236_/B _43756_/X _43766_/A
+ sky130_fd_sc_hd__o32ai_4
X_74585_ _74575_/X _74583_/X _56084_/Y _74584_/X _74585_/X sky130_fd_sc_hd__a211o_4
X_40977_ _40976_/X _40977_/X sky130_fd_sc_hd__buf_2
X_71797_ _58204_/Y _71783_/Y _71796_/Y _71797_/Y sky130_fd_sc_hd__o21ai_4
X_79112_ _82625_/D _79112_/B _79114_/A sky130_fd_sc_hd__nand2_4
X_45504_ _45504_/A _45490_/B _45504_/Y sky130_fd_sc_hd__nor2_4
X_76324_ _76319_/Y _76295_/Y _76323_/X _76324_/Y sky130_fd_sc_hd__o21ai_4
X_42716_ _41165_/X _42710_/X _68624_/B _42711_/X _87753_/D sky130_fd_sc_hd__a2bb2o_4
X_49272_ _48995_/A _49273_/A sky130_fd_sc_hd__buf_2
X_61550_ _61541_/A _61549_/X _61541_/C _61550_/Y sky130_fd_sc_hd__nand3_4
X_73536_ _72721_/X _86178_/Q _44194_/X _73535_/X _73536_/X sky130_fd_sc_hd__a211o_4
X_46484_ _54043_/A _52524_/A sky130_fd_sc_hd__buf_2
X_70748_ _53115_/B _70738_/X _70747_/Y _70748_/Y sky130_fd_sc_hd__o21ai_4
X_43696_ _43673_/A _43696_/X sky130_fd_sc_hd__buf_2
X_48223_ _48220_/Y _48175_/X _48222_/Y _86553_/D sky130_fd_sc_hd__a21boi_4
X_60501_ _60501_/A _60501_/Y sky130_fd_sc_hd__inv_2
X_79043_ _79044_/A _79044_/C _79044_/B _79057_/A sky130_fd_sc_hd__a21o_4
X_45435_ _63030_/B _61358_/A sky130_fd_sc_hd__buf_2
X_76255_ _76255_/A _76255_/Y sky130_fd_sc_hd__inv_2
X_42647_ _42590_/A _42647_/X sky130_fd_sc_hd__buf_2
X_61481_ _84821_/Q _61481_/X sky130_fd_sc_hd__buf_2
X_73467_ _73463_/X _73466_/X _73347_/X _73481_/B sky130_fd_sc_hd__a21o_4
X_70679_ _70679_/A _70676_/B _70676_/C _70679_/Y sky130_fd_sc_hd__nor3_4
X_63220_ _58440_/Y _63170_/X _63295_/C _63267_/D _63220_/X sky130_fd_sc_hd__or4_4
X_75206_ _75203_/Y _75207_/A sky130_fd_sc_hd__inv_2
X_72418_ _72413_/X _72415_/Y _72416_/Y _72337_/X _72417_/X _72418_/X
+ sky130_fd_sc_hd__o32a_4
X_48154_ _48725_/A _50389_/B _48154_/Y sky130_fd_sc_hd__nand2_4
X_60432_ _60482_/A _60443_/A sky130_fd_sc_hd__buf_2
X_45366_ _45363_/X _45365_/Y _45348_/X _45366_/Y sky130_fd_sc_hd__a21oi_4
X_76186_ _76186_/A _76189_/A sky130_fd_sc_hd__inv_2
X_42578_ _42578_/A _87814_/D sky130_fd_sc_hd__inv_2
X_73398_ _73395_/X _73397_/X _73347_/X _73412_/B sky130_fd_sc_hd__a21o_4
X_47105_ _47113_/A _47082_/X _47091_/X _52857_/D _47105_/X sky130_fd_sc_hd__and4_4
X_44317_ _44153_/X _44313_/A _44210_/X _43975_/B _44316_/X _44317_/X
+ sky130_fd_sc_hd__o32a_4
X_63151_ _63148_/Y _63150_/X _63114_/X _63151_/Y sky130_fd_sc_hd__a21oi_4
X_75137_ _80774_/Q _81030_/D _80742_/D sky130_fd_sc_hd__xor2_4
X_41529_ _41529_/A _41529_/X sky130_fd_sc_hd__buf_2
X_48085_ _47857_/X _48138_/A sky130_fd_sc_hd__buf_2
X_60363_ _62678_/A _60273_/X _60263_/C _60363_/Y sky130_fd_sc_hd__a21oi_4
X_72349_ _72299_/X _72347_/Y _72348_/Y _72337_/X _72303_/X _72349_/X
+ sky130_fd_sc_hd__o32a_4
X_45297_ _45297_/A _45297_/X sky130_fd_sc_hd__buf_2
X_62102_ _62050_/X _62090_/B _78056_/B _62102_/Y sky130_fd_sc_hd__nor3_4
X_47036_ _46941_/A _47039_/B sky130_fd_sc_hd__buf_2
X_44248_ _58602_/A _72296_/A sky130_fd_sc_hd__buf_2
X_75068_ _80744_/Q _75061_/B _75069_/B sky130_fd_sc_hd__nand2_4
X_79945_ _79945_/A _79945_/B _79946_/A sky130_fd_sc_hd__nand2_4
X_63082_ _63080_/Y _63081_/X _63056_/X _63082_/Y sky130_fd_sc_hd__a21oi_4
X_60294_ _60317_/A _60244_/B _79784_/A _60294_/Y sky130_fd_sc_hd__nor3_4
X_74019_ _72877_/A _74019_/X sky130_fd_sc_hd__buf_2
X_66910_ _66910_/A _66910_/X sky130_fd_sc_hd__buf_2
X_62033_ _62033_/A _62033_/X sky130_fd_sc_hd__buf_2
X_44179_ _45924_/A _64713_/A sky130_fd_sc_hd__buf_2
X_67890_ _87964_/Q _67888_/X _67865_/X _67889_/X _67890_/X sky130_fd_sc_hd__a211o_4
X_79876_ _79844_/X _79866_/B _79861_/X _79865_/B _79876_/X sky130_fd_sc_hd__o22a_4
X_66841_ _66840_/X _86827_/Q _66841_/X sky130_fd_sc_hd__and2_4
X_78827_ _78828_/A _78828_/C _78828_/B _78829_/A sky130_fd_sc_hd__a21o_4
X_48987_ _48946_/X _48473_/A _48986_/Y _48988_/A sky130_fd_sc_hd__a21o_4
X_69560_ _69557_/X _69559_/X _69433_/X _69560_/Y sky130_fd_sc_hd__a21oi_4
X_47938_ _47933_/Y _47903_/X _47937_/X _86584_/D sky130_fd_sc_hd__a21oi_4
X_78758_ _78758_/A _78756_/Y _78758_/C _78770_/D sky130_fd_sc_hd__nand3_4
X_66772_ _66795_/A _87627_/Q _66772_/X sky130_fd_sc_hd__and2_4
X_63984_ _57683_/X _64046_/B _64046_/C _64016_/D _63985_/D sky130_fd_sc_hd__nand4_4
X_68511_ _87098_/Q _68455_/X _68509_/X _68510_/X _68511_/X sky130_fd_sc_hd__a211o_4
X_65723_ _65769_/A _86510_/Q _65723_/X sky130_fd_sc_hd__and2_4
X_77709_ _77675_/A _77676_/X _77700_/X _77709_/X sky130_fd_sc_hd__a21o_4
X_62935_ _62965_/A _62935_/B _62113_/X _62935_/Y sky130_fd_sc_hd__nand3_4
X_69491_ _69190_/A _69580_/A sky130_fd_sc_hd__buf_2
X_47869_ _47869_/A _47915_/B _47869_/Y sky130_fd_sc_hd__nand2_4
X_78689_ _78689_/A _78689_/Y sky130_fd_sc_hd__inv_2
X_49608_ _49607_/X _51130_/B _49608_/Y sky130_fd_sc_hd__nand2_4
X_80720_ _80720_/CLK _75906_/X _80688_/D sky130_fd_sc_hd__dfxtp_4
X_68442_ _68442_/A _68442_/X sky130_fd_sc_hd__buf_2
X_65654_ _58876_/A _65654_/X sky130_fd_sc_hd__buf_2
X_50880_ _51396_/A _50825_/B _50830_/C _50880_/X sky130_fd_sc_hd__and3_4
X_62866_ _58478_/A _62841_/X _60309_/C _60254_/B _62866_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_7_63_0_CLK clkbuf_7_63_0_CLK/A clkbuf_7_63_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_64605_ _64595_/X _64633_/B _64604_/X _64605_/Y sky130_fd_sc_hd__nand3_4
X_49539_ _49546_/A _52752_/B _49539_/Y sky130_fd_sc_hd__nand2_4
X_80651_ _86757_/CLK _80651_/D _46111_/A sky130_fd_sc_hd__dfxtp_4
X_61817_ _61722_/A _61865_/A sky130_fd_sc_hd__buf_2
X_68373_ _68369_/X _68372_/X _68327_/X _68373_/Y sky130_fd_sc_hd__a21oi_4
X_65585_ _65524_/X _83071_/Q _65568_/X _65584_/X _65585_/X sky130_fd_sc_hd__a211o_4
X_62797_ _62819_/A _84829_/Q _62819_/C _62782_/X _62797_/X sky130_fd_sc_hd__and4_4
X_67324_ _67324_/A _67324_/B _67324_/X sky130_fd_sc_hd__and2_4
X_52550_ _52177_/A _52567_/A sky130_fd_sc_hd__buf_2
X_64536_ _64546_/A _64525_/B _64536_/C _64536_/X sky130_fd_sc_hd__and3_4
X_83370_ _83367_/CLK _83370_/D _83370_/Q sky130_fd_sc_hd__dfxtp_4
X_61748_ _61747_/X _61748_/X sky130_fd_sc_hd__buf_2
X_80582_ _80566_/Y _80570_/B _80582_/X sky130_fd_sc_hd__or2_4
XPHY_309 sky130_fd_sc_hd__decap_3
X_51501_ _51491_/A _53025_/B _51501_/Y sky130_fd_sc_hd__nand2_4
X_82321_ _82327_/CLK _77110_/B _82321_/Q sky130_fd_sc_hd__dfxtp_4
X_67255_ _67014_/X _67255_/X sky130_fd_sc_hd__buf_2
X_52481_ _85813_/Q _52470_/X _52480_/Y _52481_/Y sky130_fd_sc_hd__o21ai_4
X_64467_ _64474_/A _64421_/X _64467_/C _64467_/X sky130_fd_sc_hd__and3_4
X_61679_ _61673_/Y _61675_/Y _61594_/X _61676_/Y _61678_/Y _61679_/X
+ sky130_fd_sc_hd__a41o_4
Xclkbuf_7_78_0_CLK clkbuf_7_78_0_CLK/A clkbuf_7_78_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_54220_ _54249_/A _54220_/X sky130_fd_sc_hd__buf_2
X_66206_ _66123_/A _66151_/B _80419_/B _66206_/X sky130_fd_sc_hd__and3_4
X_85040_ _85040_/CLK _85040_/D _57283_/B sky130_fd_sc_hd__dfxtp_4
X_51432_ _86011_/Q _51429_/X _51431_/Y _51432_/Y sky130_fd_sc_hd__o21ai_4
X_63418_ _64257_/A _63465_/B _63418_/C _63465_/D _63418_/Y sky130_fd_sc_hd__nand4_4
X_82252_ _83278_/CLK _80409_/X _82252_/Q sky130_fd_sc_hd__dfxtp_4
X_67186_ _67166_/X _67175_/Y _67152_/X _67185_/Y _67186_/X sky130_fd_sc_hd__a211o_4
X_64398_ _79722_/B _64373_/X _64397_/X _64398_/X sky130_fd_sc_hd__a21o_4
X_81203_ _81197_/CLK _75024_/X _49029_/A sky130_fd_sc_hd__dfxtp_4
X_54151_ _54127_/X _54160_/B _54146_/X _52982_/D _54151_/X sky130_fd_sc_hd__and4_4
X_66137_ _66065_/A _66137_/X sky130_fd_sc_hd__buf_2
X_51363_ _51790_/A _51364_/A sky130_fd_sc_hd__buf_2
X_63349_ _59448_/A _60493_/A _64190_/A _60555_/A _63349_/X sky130_fd_sc_hd__a2bb2o_4
X_82183_ _84951_/CLK _82183_/D _82183_/Q sky130_fd_sc_hd__dfxtp_4
X_53102_ _85697_/Q _53093_/X _53101_/Y _53102_/Y sky130_fd_sc_hd__o21ai_4
X_50314_ _50314_/A _74509_/C _50247_/X _50314_/X sky130_fd_sc_hd__and3_4
X_81134_ _81134_/CLK _81134_/D _40694_/A sky130_fd_sc_hd__dfxtp_4
X_54082_ _85508_/Q _54067_/X _54081_/Y _54082_/Y sky130_fd_sc_hd__o21ai_4
X_66068_ _65516_/A _66068_/X sky130_fd_sc_hd__buf_2
X_51294_ _51298_/A _51294_/B _51294_/X sky130_fd_sc_hd__and2_4
X_86991_ _86982_/CLK _86991_/D _44709_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_141_0_CLK clkbuf_7_70_0_CLK/X clkbuf_9_283_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_53033_ _53025_/A _53033_/B _53033_/Y sky130_fd_sc_hd__nand2_4
X_57910_ _57905_/Y _57907_/Y _57909_/X _57910_/X sky130_fd_sc_hd__a21o_4
X_65019_ _65019_/A _65018_/Y _65019_/Y sky130_fd_sc_hd__nand2_4
X_50245_ _50256_/A _50537_/A sky130_fd_sc_hd__buf_2
X_85942_ _82768_/CLK _51811_/Y _85942_/Q sky130_fd_sc_hd__dfxtp_4
X_81065_ _81065_/CLK _81097_/Q _75175_/B sky130_fd_sc_hd__dfxtp_4
X_58890_ _58835_/X _85448_/Q _58889_/X _58890_/Y sky130_fd_sc_hd__o21ai_4
X_80016_ _80005_/X _80006_/X _80015_/Y _80016_/Y sky130_fd_sc_hd__a21boi_4
X_57841_ _57836_/Y _57840_/Y _57829_/X _57841_/X sky130_fd_sc_hd__a21o_4
X_69827_ _87052_/Q _66608_/X _58827_/A _69826_/X _69827_/X sky130_fd_sc_hd__a211o_4
X_50176_ _50174_/Y _50166_/X _50175_/X _50176_/Y sky130_fd_sc_hd__a21oi_4
X_85873_ _85859_/CLK _85873_/D _85873_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_16_0_CLK clkbuf_6_8_0_CLK/X clkbuf_7_16_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_87612_ _82899_/CLK _87612_/D _87612_/Q sky130_fd_sc_hd__dfxtp_4
X_84824_ _83438_/CLK _84824_/D _84824_/Q sky130_fd_sc_hd__dfxtp_4
X_57772_ _57965_/A _57947_/A sky130_fd_sc_hd__buf_2
X_69758_ _69758_/A _69758_/B _69758_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_156_0_CLK clkbuf_7_78_0_CLK/X clkbuf_9_313_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_54984_ _54982_/Y _54971_/X _54983_/X _54984_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_151_0_CLK clkbuf_9_75_0_CLK/X _81689_/CLK sky130_fd_sc_hd__clkbuf_1
X_59511_ _69814_/A _59512_/A sky130_fd_sc_hd__buf_2
X_56723_ _56609_/X _56723_/B _56723_/Y sky130_fd_sc_hd__nand2_4
X_68709_ _87090_/Q _68707_/X _68630_/X _68708_/X _68709_/X sky130_fd_sc_hd__a211o_4
X_87543_ _87544_/CLK _43198_/Y _73465_/A sky130_fd_sc_hd__dfxtp_4
X_53935_ _53933_/Y _53914_/X _53934_/Y _85539_/D sky130_fd_sc_hd__a21boi_4
X_84755_ _84757_/CLK _84755_/D _84755_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_781_0_CLK clkbuf_9_390_0_CLK/X _82711_/CLK sky130_fd_sc_hd__clkbuf_1
X_81967_ _82558_/CLK _81967_/D _81967_/Q sky130_fd_sc_hd__dfxtp_4
X_69689_ _69686_/X _69688_/X _69678_/X _69689_/X sky130_fd_sc_hd__a21o_4
X_40900_ _40899_/X _40821_/X _88314_/Q _40822_/X _40900_/X sky130_fd_sc_hd__a2bb2o_4
X_71720_ _58220_/Y _71718_/X _71719_/Y _83400_/D sky130_fd_sc_hd__o21ai_4
X_59442_ _58982_/A _59442_/X sky130_fd_sc_hd__buf_2
X_83706_ _83707_/CLK _83706_/D _83706_/Q sky130_fd_sc_hd__dfxtp_4
X_80918_ _81507_/CLK _80918_/D _80918_/Q sky130_fd_sc_hd__dfxtp_4
X_56654_ _57131_/A _56653_/Y _56655_/A sky130_fd_sc_hd__nor2_4
X_87474_ _88180_/CLK _87474_/D _87474_/Q sky130_fd_sc_hd__dfxtp_4
X_41880_ _41880_/A _41881_/A sky130_fd_sc_hd__buf_2
X_53866_ _85552_/Q _53784_/X _53865_/Y _53866_/Y sky130_fd_sc_hd__o21ai_4
X_84686_ _84713_/CLK _59861_/Y _80323_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_272_0_CLK clkbuf_8_136_0_CLK/X clkbuf_9_272_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_81898_ _82116_/CLK _81898_/D _82274_/D sky130_fd_sc_hd__dfxtp_4
X_55605_ _44116_/B _55605_/X sky130_fd_sc_hd__buf_2
X_86425_ _86424_/CLK _86425_/D _86425_/Q sky130_fd_sc_hd__dfxtp_4
X_40831_ _40831_/A _40831_/X sky130_fd_sc_hd__buf_2
X_52817_ _52845_/A _52818_/C sky130_fd_sc_hd__buf_2
X_59373_ _59373_/A _59226_/B _59373_/Y sky130_fd_sc_hd__nor2_4
X_71651_ _58500_/Y _71649_/X _71650_/Y _83425_/D sky130_fd_sc_hd__o21ai_4
X_83637_ _86424_/CLK _70999_/Y _46476_/A sky130_fd_sc_hd__dfxtp_4
X_56585_ _56568_/X _56584_/X _55590_/B _56572_/X _56585_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_10_166_0_CLK clkbuf_9_83_0_CLK/X _81250_/CLK sky130_fd_sc_hd__clkbuf_1
X_80849_ _80849_/CLK _80881_/Q _80849_/Q sky130_fd_sc_hd__dfxtp_4
X_53797_ _85566_/Q _53722_/X _53796_/Y _53797_/Y sky130_fd_sc_hd__o21ai_4
X_70602_ _70771_/A _70714_/A sky130_fd_sc_hd__buf_2
X_58324_ _58310_/X _83454_/Q _58323_/Y _84878_/D sky130_fd_sc_hd__o21a_4
X_43550_ _43542_/X _43546_/X _40452_/X _87365_/Q _43549_/X _43550_/Y
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_10_796_0_CLK clkbuf_9_398_0_CLK/X _82692_/CLK sky130_fd_sc_hd__clkbuf_1
X_55536_ _55536_/A _55526_/X _55536_/C _55536_/D _55536_/X sky130_fd_sc_hd__and4_4
X_74370_ _71978_/A _74370_/X sky130_fd_sc_hd__buf_2
X_86356_ _86359_/CLK _49611_/Y _59167_/B sky130_fd_sc_hd__dfxtp_4
X_40762_ _40762_/A _40762_/X sky130_fd_sc_hd__buf_2
X_52748_ _52744_/A _52748_/B _52748_/Y sky130_fd_sc_hd__nand2_4
X_71582_ _71189_/B _71582_/X sky130_fd_sc_hd__buf_2
X_83568_ _86500_/CLK _71220_/Y _48638_/A sky130_fd_sc_hd__dfxtp_4
X_42501_ _41993_/A _42501_/X sky130_fd_sc_hd__buf_2
X_73321_ _69860_/B _73319_/X _72890_/X _73320_/Y _73321_/X sky130_fd_sc_hd__a211o_4
X_85307_ _85213_/CLK _85307_/D _55934_/B sky130_fd_sc_hd__dfxtp_4
X_70533_ _70532_/Y _70533_/X sky130_fd_sc_hd__buf_2
X_58255_ _58273_/A _58268_/B sky130_fd_sc_hd__buf_2
X_82519_ _82518_/CLK _82519_/D _82519_/Q sky130_fd_sc_hd__dfxtp_4
X_43481_ _43480_/Y _87401_/D sky130_fd_sc_hd__inv_2
Xclkbuf_9_287_0_CLK clkbuf_9_286_0_CLK/A clkbuf_9_287_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_55467_ _55466_/X _55467_/X sky130_fd_sc_hd__buf_2
X_86287_ _86610_/CLK _49985_/Y _86287_/Q sky130_fd_sc_hd__dfxtp_4
X_40693_ _40692_/Y _88353_/D sky130_fd_sc_hd__inv_2
X_52679_ _52679_/A _52708_/A sky130_fd_sc_hd__buf_2
X_83499_ _81233_/CLK _71438_/X _83499_/Q sky130_fd_sc_hd__dfxtp_4
X_45220_ _45202_/X _61568_/B _45219_/X _45220_/Y sky130_fd_sc_hd__o21ai_4
X_57206_ _57204_/X _57205_/Y _57112_/X _57206_/Y sky130_fd_sc_hd__a21oi_4
X_76040_ _81522_/Q _76040_/B _81771_/D sky130_fd_sc_hd__xor2_4
X_88026_ _87776_/CLK _42119_/Y _88026_/Q sky130_fd_sc_hd__dfxtp_4
X_42432_ _42432_/A _42432_/Y sky130_fd_sc_hd__inv_2
X_54418_ _54416_/Y _54394_/X _54417_/X _85446_/D sky130_fd_sc_hd__a21oi_4
X_73252_ _73252_/A _73228_/B _73252_/Y sky130_fd_sc_hd__nor2_4
X_85238_ _85269_/CLK _85238_/D _56317_/C sky130_fd_sc_hd__dfxtp_4
X_70464_ _71323_/A _71500_/C _71672_/C _70464_/Y sky130_fd_sc_hd__nand3_4
X_58186_ _83376_/Q _58186_/Y sky130_fd_sc_hd__inv_2
X_55398_ _55298_/A _55398_/Y sky130_fd_sc_hd__inv_2
X_72203_ _83275_/Q _72115_/X _72195_/X _72202_/X _83275_/D sky130_fd_sc_hd__a2bb2oi_4
X_45151_ _85201_/Q _45102_/X _45150_/X _45151_/Y sky130_fd_sc_hd__o21ai_4
X_57137_ _57137_/A _45888_/A _57137_/X sky130_fd_sc_hd__or2_4
X_54349_ _54320_/A _54349_/X sky130_fd_sc_hd__buf_2
X_42363_ _41749_/X _42356_/X _87900_/Q _42357_/X _87900_/D sky130_fd_sc_hd__a2bb2o_4
X_73183_ _73183_/A _86481_/Q _73183_/X sky130_fd_sc_hd__and2_4
X_85169_ _85168_/CLK _85169_/D _55833_/B sky130_fd_sc_hd__dfxtp_4
X_70395_ _70786_/A _74529_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_210_0_CLK clkbuf_9_210_0_CLK/A clkbuf_9_210_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_44102_ _44102_/A _44102_/X sky130_fd_sc_hd__buf_2
X_41314_ _41314_/A _41275_/B _41314_/X sky130_fd_sc_hd__or2_4
X_72134_ _59381_/X _85984_/Q _72133_/X _72134_/Y sky130_fd_sc_hd__o21ai_4
X_45082_ _45082_/A _45067_/B _45082_/Y sky130_fd_sc_hd__nand2_4
X_57068_ _56649_/X _57067_/Y _56892_/B _57068_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_8_109_0_CLK clkbuf_7_54_0_CLK/X clkbuf_9_219_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_42294_ _42279_/X _42275_/X _41565_/X _87935_/Q _42276_/X _42294_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77991_ _77977_/Y _77975_/Y _77967_/C _77967_/B _77990_/Y _77991_/X
+ sky130_fd_sc_hd__o41a_4
Xclkbuf_10_104_0_CLK clkbuf_9_52_0_CLK/X _85071_/CLK sky130_fd_sc_hd__clkbuf_1
X_48910_ _83622_/Q _71972_/B sky130_fd_sc_hd__inv_2
X_44033_ _44012_/A _64850_/A sky130_fd_sc_hd__buf_2
X_56019_ _55966_/X _56019_/B _56019_/Y sky130_fd_sc_hd__xnor2_4
X_79730_ _84218_/Q _83266_/Q _79730_/Y sky130_fd_sc_hd__nand2_4
X_41245_ _41244_/X _41245_/X sky130_fd_sc_hd__buf_2
X_72065_ _72063_/Y _72059_/X _72064_/X _72065_/Y sky130_fd_sc_hd__a21oi_4
X_76942_ _76939_/X _76942_/B _76953_/A _76942_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_734_0_CLK clkbuf_9_367_0_CLK/X _87790_/CLK sky130_fd_sc_hd__clkbuf_1
X_49890_ _49887_/Y _49870_/X _49889_/X _49890_/Y sky130_fd_sc_hd__a21oi_4
X_71016_ _71016_/A _71039_/D sky130_fd_sc_hd__buf_2
X_48841_ _48841_/A _48849_/B _48849_/C _48841_/X sky130_fd_sc_hd__and3_4
X_79661_ _79660_/X _79667_/A sky130_fd_sc_hd__inv_2
X_41176_ _41176_/A _41176_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_9_225_0_CLK clkbuf_8_112_0_CLK/X clkbuf_9_225_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_76873_ _76873_/A _76873_/Y sky130_fd_sc_hd__inv_2
X_78612_ _78611_/A _82679_/D _78613_/A sky130_fd_sc_hd__nand2_4
X_75824_ _75824_/A _75824_/B _75824_/Y sky130_fd_sc_hd__nand2_4
X_48772_ _48769_/Y _48760_/X _48771_/X _86486_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_119_0_CLK clkbuf_9_59_0_CLK/X _84555_/CLK sky130_fd_sc_hd__clkbuf_1
X_79592_ _79592_/A _79591_/Y _79592_/Y sky130_fd_sc_hd__nand2_4
X_45984_ _45984_/A _45984_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_749_0_CLK clkbuf_9_374_0_CLK/X _87249_/CLK sky130_fd_sc_hd__clkbuf_1
X_47723_ _47758_/A _47739_/B _47749_/C _53207_/D _47723_/X sky130_fd_sc_hd__and4_4
X_59709_ _57754_/X _63055_/A sky130_fd_sc_hd__buf_2
X_78543_ _78539_/Y _78519_/B _78542_/X _78561_/A sky130_fd_sc_hd__o21ai_4
X_44935_ _45705_/A _44935_/X sky130_fd_sc_hd__buf_2
X_75755_ _75733_/Y _80788_/D sky130_fd_sc_hd__inv_2
X_60981_ _60926_/X _60930_/A _60982_/A sky130_fd_sc_hd__nor2_4
X_72967_ _53651_/B _72967_/B _72967_/X sky130_fd_sc_hd__xor2_4
X_62720_ _61348_/A _62893_/A sky130_fd_sc_hd__buf_2
X_74706_ _74630_/X _57083_/X _74705_/Y _74706_/X sky130_fd_sc_hd__o21a_4
X_47654_ _55031_/D _53170_/D sky130_fd_sc_hd__buf_2
X_71918_ _70368_/X _70979_/C _71902_/X _71928_/D _71918_/Y sky130_fd_sc_hd__nand4_4
X_78474_ _78474_/A _78473_/X _78482_/A sky130_fd_sc_hd__xnor2_4
X_44866_ _44857_/X _44865_/X _41790_/X _86912_/Q _44858_/X _44867_/A
+ sky130_fd_sc_hd__o32ai_4
X_75686_ _81006_/Q _75686_/B _75686_/X sky130_fd_sc_hd__xor2_4
X_72898_ _72893_/X _72897_/X _72862_/X _72898_/X sky130_fd_sc_hd__a21o_4
X_46605_ _46597_/Y _46598_/X _46604_/X _86722_/D sky130_fd_sc_hd__a21oi_4
X_77425_ _77424_/Y _77426_/C sky130_fd_sc_hd__inv_2
X_43817_ _43752_/A _43817_/X sky130_fd_sc_hd__buf_2
X_62651_ _62638_/Y _62642_/Y _62648_/X _58147_/A _62650_/X _62651_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74637_ _45952_/X _56583_/X _83005_/Q _74633_/X _83005_/D sky130_fd_sc_hd__a2bb2o_4
X_47585_ _47585_/A _47586_/A sky130_fd_sc_hd__inv_2
X_71849_ _71846_/A _71867_/B sky130_fd_sc_hd__buf_2
X_44797_ _44797_/A _44797_/Y sky130_fd_sc_hd__inv_2
X_49324_ _49287_/A _51358_/B _49324_/Y sky130_fd_sc_hd__nand2_4
X_61602_ _61590_/Y _61593_/Y _61594_/X _61597_/Y _61601_/Y _61602_/X
+ sky130_fd_sc_hd__a41o_4
X_46536_ _86728_/Q _46430_/X _46535_/Y _46536_/Y sky130_fd_sc_hd__o21ai_4
X_65370_ _65198_/X _65359_/Y _65369_/Y _65370_/Y sky130_fd_sc_hd__o21ai_4
X_77356_ _77338_/A _77338_/B _77356_/Y sky130_fd_sc_hd__nand2_4
X_62582_ _62576_/X _62578_/X _62581_/Y _58352_/A _62572_/X _62582_/Y
+ sky130_fd_sc_hd__o32ai_4
X_43748_ _40925_/X _43736_/X _73509_/A _43737_/X _43748_/X sky130_fd_sc_hd__a2bb2o_4
X_74568_ _74549_/Y _74568_/X sky130_fd_sc_hd__buf_2
X_64321_ _64295_/A _64307_/B _84832_/Q _64321_/X sky130_fd_sc_hd__and3_4
X_76307_ _76306_/X _76321_/A sky130_fd_sc_hd__buf_2
X_49255_ _48548_/A _49255_/X sky130_fd_sc_hd__buf_2
X_73519_ _73476_/A _86499_/Q _73519_/X sky130_fd_sc_hd__and2_4
X_61533_ _61521_/Y _61524_/Y _61525_/X _61528_/Y _61532_/Y _61533_/X
+ sky130_fd_sc_hd__a41o_4
X_46467_ _86734_/Q _46292_/X _46466_/Y _46467_/Y sky130_fd_sc_hd__o21ai_4
X_77287_ _77287_/A _77286_/Y _77318_/A sky130_fd_sc_hd__nor2_4
X_43679_ _40771_/X _43671_/X _87314_/Q _43673_/X _43679_/X sky130_fd_sc_hd__a2bb2o_4
X_74499_ _46272_/A _48672_/A _74499_/Y sky130_fd_sc_hd__nand2_4
X_48206_ _73689_/B _48203_/X _48205_/Y _48206_/Y sky130_fd_sc_hd__o21ai_4
X_67040_ _67039_/X _67040_/X sky130_fd_sc_hd__buf_2
X_79026_ _79022_/Y _79010_/B _79025_/Y _79027_/B sky130_fd_sc_hd__o21ai_4
X_45418_ _45416_/Y _45417_/Y _44901_/X _45418_/X sky130_fd_sc_hd__o21a_4
X_64252_ _64245_/X _64246_/X _64248_/X _64251_/Y _64229_/X _64252_/X
+ sky130_fd_sc_hd__o41a_4
X_76238_ _76236_/X _76237_/Y _76238_/X sky130_fd_sc_hd__and2_4
X_49186_ _49156_/X _50716_/B _49186_/Y sky130_fd_sc_hd__nand2_4
X_61464_ _61334_/A _61464_/X sky130_fd_sc_hd__buf_2
X_46398_ _44803_/A _46399_/A sky130_fd_sc_hd__buf_2
X_63203_ _60503_/X _63203_/X sky130_fd_sc_hd__buf_2
X_48137_ _48134_/X _82916_/Q _48136_/X _48342_/A sky130_fd_sc_hd__o21ai_4
X_60415_ _60606_/A _60447_/B sky130_fd_sc_hd__inv_2
X_45349_ _45344_/X _45347_/Y _45348_/X _45349_/Y sky130_fd_sc_hd__a21oi_4
X_76169_ _76169_/A _81603_/D sky130_fd_sc_hd__buf_2
X_64183_ _61683_/X _64172_/B _64172_/C _64172_/D _64183_/Y sky130_fd_sc_hd__nand4_4
X_61395_ _61384_/A _61384_/B _79152_/B _61395_/Y sky130_fd_sc_hd__nor3_4
X_63134_ _60458_/X _63135_/D sky130_fd_sc_hd__buf_2
X_48068_ _48790_/A _48723_/C sky130_fd_sc_hd__buf_2
X_60346_ _60477_/A _60319_/X _60346_/C _60346_/Y sky130_fd_sc_hd__nor3_4
X_68991_ _41963_/A _68989_/X _68555_/X _68990_/Y _68991_/X sky130_fd_sc_hd__a211o_4
X_47019_ _82391_/Q _54498_/D sky130_fd_sc_hd__inv_2
X_67942_ _67466_/X _67942_/X sky130_fd_sc_hd__buf_2
X_63065_ _60484_/A _63066_/D sky130_fd_sc_hd__buf_2
X_79928_ _79928_/A _79928_/B _79928_/Y sky130_fd_sc_hd__nor2_4
X_60277_ _60344_/C _60268_/C _60344_/B _60324_/C _60277_/X sky130_fd_sc_hd__a211o_4
X_50030_ _46308_/A _50050_/A sky130_fd_sc_hd__buf_2
X_62016_ _62004_/X _62006_/X _62015_/Y _84847_/Q _61973_/X _62016_/Y
+ sky130_fd_sc_hd__o32ai_4
X_79859_ _79859_/A _79858_/Y _79859_/X sky130_fd_sc_hd__xor2_4
X_67873_ _67873_/A _67873_/B _67873_/X sky130_fd_sc_hd__and2_4
X_69612_ _69612_/A _69612_/B _69612_/X sky130_fd_sc_hd__and2_4
X_66824_ _87125_/Q _66751_/X _66801_/X _66823_/X _66824_/X sky130_fd_sc_hd__a211o_4
X_82870_ _82498_/CLK _78228_/B _82870_/Q sky130_fd_sc_hd__dfxtp_4
X_81821_ _81275_/CLK _81821_/D _81821_/Q sky130_fd_sc_hd__dfxtp_4
X_69543_ _88021_/Q _69424_/X _69465_/X _69542_/X _69543_/X sky130_fd_sc_hd__a211o_4
X_66755_ _66499_/B _66743_/Y _66672_/X _66754_/Y _66755_/X sky130_fd_sc_hd__a211o_4
X_51981_ _51934_/A _51981_/X sky130_fd_sc_hd__buf_2
X_63967_ _63966_/Y _63967_/Y sky130_fd_sc_hd__inv_2
X_53720_ _52204_/A _53720_/B _53734_/C _53720_/X sky130_fd_sc_hd__and3_4
X_65706_ _65703_/X _65705_/X _65642_/X _65710_/A sky130_fd_sc_hd__a21o_4
X_84540_ _84292_/CLK _61015_/Y _84540_/Q sky130_fd_sc_hd__dfxtp_4
X_50932_ _50932_/A _46701_/X _50932_/Y sky130_fd_sc_hd__nand2_4
X_62918_ _58498_/A _60304_/A _64473_/A _62875_/X _62918_/X sky130_fd_sc_hd__o22a_4
X_81752_ _81756_/CLK _76083_/B _41330_/A sky130_fd_sc_hd__dfxtp_4
X_69474_ _69471_/X _69473_/X _69433_/X _69474_/Y sky130_fd_sc_hd__a21oi_4
X_66686_ _66526_/X _66671_/Y _66672_/X _66685_/Y _66686_/X sky130_fd_sc_hd__a211o_4
X_63898_ _63896_/X _63833_/X _63897_/Y _63898_/Y sky130_fd_sc_hd__a21oi_4
X_68425_ _68403_/A _68425_/B _68425_/X sky130_fd_sc_hd__and2_4
X_80703_ _81121_/CLK _80703_/D _80703_/Q sky130_fd_sc_hd__dfxtp_4
X_53651_ _53656_/A _53651_/B _53651_/Y sky130_fd_sc_hd__nand2_4
X_65637_ _65484_/X _86195_/Q _65534_/X _65636_/X _65637_/X sky130_fd_sc_hd__a211o_4
X_84471_ _82822_/CLK _61556_/Y _84471_/Q sky130_fd_sc_hd__dfxtp_4
X_50863_ _86118_/Q _50856_/X _50862_/Y _50863_/Y sky130_fd_sc_hd__o21ai_4
X_62849_ _62843_/X _62831_/X _62844_/Y _62846_/Y _62848_/X _62849_/X
+ sky130_fd_sc_hd__a41o_4
X_81683_ _81697_/CLK _81683_/D _76656_/B sky130_fd_sc_hd__dfxtp_4
X_86210_ _86210_/CLK _50392_/Y _86210_/Q sky130_fd_sc_hd__dfxtp_4
X_52602_ _52602_/A _52624_/A sky130_fd_sc_hd__buf_2
X_83422_ _84945_/CLK _71659_/Y _58513_/A sky130_fd_sc_hd__dfxtp_4
X_80634_ _80632_/Y _80633_/Y _80634_/Y sky130_fd_sc_hd__nand2_4
X_56370_ _56183_/X _56460_/B _56370_/C _56460_/D _56370_/Y sky130_fd_sc_hd__nand4_4
X_68356_ _87103_/Q _68353_/X _68354_/X _68355_/X _68356_/X sky130_fd_sc_hd__a211o_4
X_87190_ _87221_/CLK _43937_/Y _87190_/Q sky130_fd_sc_hd__dfxtp_4
X_53582_ _85608_/Q _53556_/X _53581_/Y _53582_/Y sky130_fd_sc_hd__o21ai_4
X_65568_ _65768_/A _65568_/X sky130_fd_sc_hd__buf_2
X_50794_ _50791_/Y _50792_/X _50793_/Y _86132_/D sky130_fd_sc_hd__a21boi_4
X_55321_ _85102_/Q _55305_/X _44045_/X _55320_/Y _55321_/X sky130_fd_sc_hd__a211o_4
X_86141_ _86045_/CLK _50752_/Y _86141_/Q sky130_fd_sc_hd__dfxtp_4
X_67307_ _87860_/Q _67236_/X _67284_/X _67306_/X _67307_/X sky130_fd_sc_hd__a211o_4
XPHY_106 sky130_fd_sc_hd__decap_3
X_52533_ _52533_/A _52509_/B _50918_/A _52533_/X sky130_fd_sc_hd__and3_4
X_64519_ _79581_/B _64429_/X _64518_/X _64519_/X sky130_fd_sc_hd__a21o_4
X_83353_ _83480_/CLK _83353_/D _83353_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_117 sky130_fd_sc_hd__decap_3
X_80565_ _84771_/Q _84163_/Q _80565_/Y sky130_fd_sc_hd__nand2_4
X_68287_ _68447_/A _68287_/X sky130_fd_sc_hd__buf_2
X_65499_ _65496_/Y _65448_/X _65498_/Y _84197_/D sky130_fd_sc_hd__a21o_4
XPHY_128 sky130_fd_sc_hd__decap_3
Xclkbuf_4_13_0_CLK clkbuf_3_6_1_CLK/X clkbuf_4_13_0_CLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_139 sky130_fd_sc_hd__decap_3
X_58040_ _58010_/X _58038_/Y _58039_/Y _58028_/X _58015_/X _58040_/X
+ sky130_fd_sc_hd__o32a_4
X_82304_ _82349_/CLK _77222_/B _82304_/Q sky130_fd_sc_hd__dfxtp_4
X_55252_ _55252_/A _85128_/Q _55252_/X sky130_fd_sc_hd__and2_4
X_67238_ _87863_/Q _67236_/X _67167_/X _67237_/X _67238_/X sky130_fd_sc_hd__a211o_4
X_86072_ _85751_/CLK _86072_/D _86072_/Q sky130_fd_sc_hd__dfxtp_4
X_52464_ _52468_/A _53983_/B _52464_/Y sky130_fd_sc_hd__nand2_4
X_83284_ _86149_/CLK _72104_/Y _83284_/Q sky130_fd_sc_hd__dfxtp_4
X_80496_ _59143_/A _84157_/Q _80496_/X sky130_fd_sc_hd__xor2_4
X_54203_ _54191_/A _54191_/B _54209_/C _53036_/D _54203_/X sky130_fd_sc_hd__and4_4
X_85023_ _83008_/CLK _57387_/X _85023_/Q sky130_fd_sc_hd__dfxtp_4
X_51415_ _51170_/A _51438_/C sky130_fd_sc_hd__buf_2
X_82235_ _82515_/CLK _82267_/Q _77599_/A sky130_fd_sc_hd__dfxtp_4
X_55183_ _55245_/A _55711_/A sky130_fd_sc_hd__buf_2
X_67169_ _87930_/Q _67117_/X _67167_/X _67168_/X _67169_/X sky130_fd_sc_hd__a211o_4
X_52395_ _52385_/A _52395_/B _52395_/X sky130_fd_sc_hd__and2_4
X_54134_ _54134_/A _47297_/Y _54134_/Y sky130_fd_sc_hd__nand2_4
X_51346_ _65147_/B _51332_/X _51345_/Y _51346_/Y sky130_fd_sc_hd__o21ai_4
X_70180_ _83846_/Q _70180_/Y sky130_fd_sc_hd__inv_2
X_82166_ _86553_/CLK _84158_/Q _82166_/Q sky130_fd_sc_hd__dfxtp_4
X_59991_ _59990_/X _60129_/B sky130_fd_sc_hd__inv_2
X_81117_ _81117_/CLK _79842_/X _75669_/A sky130_fd_sc_hd__dfxtp_4
X_58942_ _58942_/A _59090_/B _58942_/Y sky130_fd_sc_hd__nor2_4
X_54065_ _54031_/A _50854_/B _54065_/Y sky130_fd_sc_hd__nand2_4
X_51277_ _64820_/B _51259_/X _51276_/Y _51277_/Y sky130_fd_sc_hd__o21ai_4
X_86974_ _88180_/CLK _44752_/X _86974_/Q sky130_fd_sc_hd__dfxtp_4
X_82097_ _82604_/CLK _77444_/B _77110_/A sky130_fd_sc_hd__dfxtp_4
X_41030_ _40852_/B _41091_/B _41030_/X sky130_fd_sc_hd__or2_4
X_53016_ _53013_/Y _53001_/X _53015_/X _53016_/Y sky130_fd_sc_hd__a21oi_4
X_50228_ _50638_/A _50228_/X sky130_fd_sc_hd__buf_2
X_85925_ _85444_/CLK _51906_/Y _85925_/Q sky130_fd_sc_hd__dfxtp_4
X_81048_ _81048_/CLK _75407_/X _81048_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_1006_0_CLK clkbuf_9_503_0_CLK/X _85879_/CLK sky130_fd_sc_hd__clkbuf_1
X_58873_ _86697_/Q _58873_/B _58873_/Y sky130_fd_sc_hd__nor2_4
X_57824_ _44181_/X _57824_/X sky130_fd_sc_hd__buf_2
X_50159_ _86252_/Q _50137_/X _50158_/Y _50159_/Y sky130_fd_sc_hd__o21ai_4
X_73870_ _88102_/Q _73869_/X _73870_/Y sky130_fd_sc_hd__nor2_4
X_85856_ _83311_/CLK _52268_/Y _85856_/Q sky130_fd_sc_hd__dfxtp_4
X_72821_ _72802_/X _72822_/C _72820_/X _72821_/X sky130_fd_sc_hd__a21o_4
X_84807_ _84807_/CLK _58695_/Y _84807_/Q sky130_fd_sc_hd__dfxtp_4
X_57755_ _57754_/X _59801_/A sky130_fd_sc_hd__buf_2
X_42981_ _42970_/X _42971_/X _40459_/X _87620_/Q _42976_/X _42981_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54967_ _55072_/A _54967_/X sky130_fd_sc_hd__buf_2
X_85787_ _85786_/CLK _52611_/Y _85787_/Q sky130_fd_sc_hd__dfxtp_4
X_82999_ _83001_/CLK _82999_/D _45558_/A sky130_fd_sc_hd__dfxtp_4
X_44720_ _44707_/X _44708_/X _40695_/Y _44719_/Y _44710_/X _86988_/D
+ sky130_fd_sc_hd__o32ai_4
X_56706_ _56702_/X _56703_/X _56705_/Y _56706_/X sky130_fd_sc_hd__a21bo_4
X_75540_ _75519_/A _75516_/Y _75517_/Y _75540_/X sky130_fd_sc_hd__o21a_4
X_87526_ _87782_/CLK _43234_/Y _87526_/Q sky130_fd_sc_hd__dfxtp_4
X_41932_ _42013_/A _41932_/X sky130_fd_sc_hd__buf_2
X_53918_ _85542_/Q _53896_/X _53917_/Y _53918_/Y sky130_fd_sc_hd__o21ai_4
X_72752_ _73535_/A _65425_/B _72752_/X sky130_fd_sc_hd__and2_4
X_84738_ _83457_/CLK _84738_/D _84738_/Q sky130_fd_sc_hd__dfxtp_4
X_57686_ _57686_/A _57701_/A _57687_/A sky130_fd_sc_hd__nor2_4
X_54898_ _54893_/X _54898_/B _54898_/Y sky130_fd_sc_hd__nand2_4
X_71703_ _58294_/Y _71695_/X _71702_/Y _83405_/D sky130_fd_sc_hd__o21ai_4
X_59425_ _59417_/X _83345_/Q _59424_/Y _84737_/D sky130_fd_sc_hd__o21a_4
X_44651_ _41058_/Y _44648_/X _87017_/Q _44650_/X _87017_/D sky130_fd_sc_hd__a2bb2o_4
X_56637_ _56650_/B _55646_/X _56638_/B sky130_fd_sc_hd__nand2_4
X_75471_ _75465_/Y _75470_/Y _81052_/D sky130_fd_sc_hd__xor2_4
X_87457_ _87720_/CLK _43366_/Y _87457_/Q sky130_fd_sc_hd__dfxtp_4
X_53849_ _85556_/Q _53846_/X _53848_/Y _53849_/Y sky130_fd_sc_hd__o21ai_4
X_41863_ _41863_/A _41862_/Y _42626_/A sky130_fd_sc_hd__nor2_4
X_72683_ _72683_/A _72683_/B _55378_/X _72683_/Y sky130_fd_sc_hd__nand3_4
X_84669_ _84498_/CLK _60060_/X _84669_/Q sky130_fd_sc_hd__dfxtp_4
X_77210_ _77200_/A _82302_/D _77210_/X sky130_fd_sc_hd__or2_4
X_43602_ _43583_/Y _43602_/X sky130_fd_sc_hd__buf_2
X_74422_ _74419_/Y _74405_/X _74421_/X _74422_/Y sky130_fd_sc_hd__a21oi_4
X_86408_ _85800_/CLK _49333_/Y _86408_/Q sky130_fd_sc_hd__dfxtp_4
X_40814_ _40814_/A _40814_/X sky130_fd_sc_hd__buf_2
X_47370_ _47380_/A _47408_/B _47370_/C _53008_/D _47370_/X sky130_fd_sc_hd__and4_4
X_71634_ _71241_/A _71637_/A sky130_fd_sc_hd__buf_2
X_59356_ _59231_/X _85412_/Q _59355_/X _59356_/Y sky130_fd_sc_hd__o21ai_4
X_78190_ _78199_/A _78199_/B _78204_/A sky130_fd_sc_hd__xor2_4
X_44582_ _44554_/X _44555_/X _40898_/Y _44581_/Y _44557_/X _87046_/D
+ sky130_fd_sc_hd__o32ai_4
X_56568_ _56567_/Y _56568_/X sky130_fd_sc_hd__buf_2
X_41794_ _41793_/Y _41794_/Y sky130_fd_sc_hd__inv_2
X_87388_ _87195_/CLK _43502_/X _87388_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_8 sky130_fd_sc_hd__decap_3
X_46321_ _53969_/A _50755_/A sky130_fd_sc_hd__buf_2
X_58307_ _84882_/Q _63348_/A sky130_fd_sc_hd__inv_2
X_77141_ _77141_/A _77141_/B _77141_/C _77142_/B sky130_fd_sc_hd__and3_4
X_43533_ _43466_/X _43533_/X sky130_fd_sc_hd__buf_2
X_55519_ _55498_/X _55524_/A sky130_fd_sc_hd__buf_2
X_74353_ _56127_/B _73050_/A _74353_/Y sky130_fd_sc_hd__nor2_4
X_86339_ _86340_/CLK _49702_/Y _59372_/B sky130_fd_sc_hd__dfxtp_4
X_40745_ _40687_/X _40688_/X _40743_/X _88343_/Q _40744_/X _40746_/A
+ sky130_fd_sc_hd__o32ai_4
X_59287_ _59199_/X _85738_/Q _59263_/X _59287_/X sky130_fd_sc_hd__o21a_4
X_71565_ _71859_/A _71553_/B _71558_/X _71565_/Y sky130_fd_sc_hd__nor3_4
X_56499_ _56528_/A _56499_/X sky130_fd_sc_hd__buf_2
X_49040_ _49018_/X _48529_/Y _49039_/Y _49041_/A sky130_fd_sc_hd__a21o_4
X_73304_ _73206_/X _85868_/Q _73304_/X sky130_fd_sc_hd__and2_4
X_46252_ _57563_/A _46280_/A sky130_fd_sc_hd__buf_2
X_70516_ _70511_/A _70947_/B _70508_/X _70516_/Y sky130_fd_sc_hd__nand3_4
X_58238_ _58237_/X _58238_/B _58238_/Y sky130_fd_sc_hd__nor2_4
XPHY_640 sky130_fd_sc_hd__decap_3
X_77072_ _77068_/Y _77072_/B _77084_/A sky130_fd_sc_hd__nand2_4
X_43464_ _41647_/X _43446_/X _87408_/Q _43447_/X _87408_/D sky130_fd_sc_hd__a2bb2o_4
X_74284_ _72714_/A _72714_/B _74284_/C _74284_/Y sky130_fd_sc_hd__nand3_4
XPHY_651 sky130_fd_sc_hd__decap_3
X_40676_ _40676_/A _40710_/B _40676_/X sky130_fd_sc_hd__or2_4
X_71496_ _71488_/X _70476_/X _71496_/C _71496_/X sky130_fd_sc_hd__and3_4
XPHY_662 sky130_fd_sc_hd__decap_3
XPHY_673 sky130_fd_sc_hd__decap_3
X_45203_ _64434_/B _61558_/B sky130_fd_sc_hd__buf_2
X_76023_ _76023_/A _76023_/B _76023_/Y sky130_fd_sc_hd__nand2_4
X_88009_ _88006_/CLK _88009_/D _88009_/Q sky130_fd_sc_hd__dfxtp_4
X_42415_ _41911_/A _42415_/X sky130_fd_sc_hd__buf_2
XPHY_684 sky130_fd_sc_hd__decap_3
X_73235_ _73260_/A _86479_/Q _73235_/X sky130_fd_sc_hd__and2_4
X_46183_ _86764_/Q _46195_/A _46183_/X sky130_fd_sc_hd__or2_4
X_70447_ _71005_/A _70954_/B sky130_fd_sc_hd__buf_2
X_58169_ _58153_/X _83492_/Q _58168_/Y _58169_/X sky130_fd_sc_hd__o21a_4
XPHY_695 sky130_fd_sc_hd__decap_3
X_43395_ _41465_/X _43386_/X _87442_/Q _43388_/X _87442_/D sky130_fd_sc_hd__a2bb2o_4
X_60200_ _60199_/X _60227_/A sky130_fd_sc_hd__buf_2
X_45134_ _45284_/A _45134_/X sky130_fd_sc_hd__buf_2
X_42346_ _42397_/A _42346_/X sky130_fd_sc_hd__buf_2
X_61180_ _61180_/A _64263_/A sky130_fd_sc_hd__buf_2
X_73166_ _73386_/A _86514_/Q _73166_/X sky130_fd_sc_hd__and2_4
X_70378_ _71054_/A _74523_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_673_0_CLK clkbuf_9_336_0_CLK/X _88158_/CLK sky130_fd_sc_hd__clkbuf_1
X_60131_ _59875_/X _62194_/A _60129_/Y _59969_/X _60130_/X _84657_/D
+ sky130_fd_sc_hd__o41a_4
X_72117_ _57696_/X _72193_/B sky130_fd_sc_hd__buf_2
X_49942_ _49915_/A _49943_/B sky130_fd_sc_hd__buf_2
X_45065_ _55900_/B _45044_/X _45004_/X _45065_/X sky130_fd_sc_hd__o21a_4
X_42277_ _42252_/X _42275_/X _41515_/X _87944_/Q _42276_/X _42277_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77974_ _82253_/Q _81965_/Q _78043_/A sky130_fd_sc_hd__xnor2_4
X_73097_ _72963_/X _83069_/Q _73015_/X _73096_/X _73097_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_9_164_0_CLK clkbuf_8_82_0_CLK/X clkbuf_9_164_0_CLK/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_9_91_0_CLK clkbuf_8_45_0_CLK/X clkbuf_9_91_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_44016_ _68617_/A _57848_/A sky130_fd_sc_hd__buf_2
X_79713_ _79713_/A _79713_/B _79719_/B sky130_fd_sc_hd__xor2_4
X_41228_ _41228_/A _41197_/B _41228_/X sky130_fd_sc_hd__or2_4
X_60062_ _59977_/A _60091_/B _59938_/Y _60062_/X sky130_fd_sc_hd__o21a_4
X_72048_ _71964_/A _72048_/X sky130_fd_sc_hd__buf_2
X_76925_ _81599_/Q _76926_/B sky130_fd_sc_hd__inv_2
X_49873_ _49869_/Y _49870_/X _49872_/X _86308_/D sky130_fd_sc_hd__a21oi_4
X_48824_ _48821_/Y _48813_/X _48823_/X _48824_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_688_0_CLK clkbuf_9_344_0_CLK/X _88215_/CLK sky130_fd_sc_hd__clkbuf_1
X_79644_ _79642_/Y _79624_/B _79643_/X _79645_/B sky130_fd_sc_hd__o21ai_4
X_41159_ _41159_/A _40639_/A _41159_/X sky130_fd_sc_hd__or2_4
X_64870_ _64870_/A _64870_/B _64870_/C _64870_/Y sky130_fd_sc_hd__nor3_4
X_76856_ _81497_/Q _76858_/A sky130_fd_sc_hd__inv_2
X_63821_ _61386_/B _63790_/X _63757_/C _63776_/X _63821_/Y sky130_fd_sc_hd__nand4_4
X_75807_ _75807_/A _80796_/D _75832_/B sky130_fd_sc_hd__xor2_4
X_48755_ _48755_/A _48837_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_179_0_CLK clkbuf_8_89_0_CLK/X clkbuf_9_179_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_79575_ _79565_/Y _79576_/B _79576_/A _79575_/Y sky130_fd_sc_hd__nand3_4
X_45967_ _44857_/X _44865_/X _40370_/X _66618_/B _44858_/X _45967_/Y
+ sky130_fd_sc_hd__o32ai_4
X_76787_ _76772_/Y _76773_/Y _76787_/Y sky130_fd_sc_hd__nor2_4
X_73999_ _73930_/X _84975_/Q _45885_/X _73998_/X _73999_/X sky130_fd_sc_hd__a211o_4
X_47706_ _47696_/A _53200_/B _47706_/Y sky130_fd_sc_hd__nand2_4
X_66540_ _66540_/A _66540_/X sky130_fd_sc_hd__buf_2
X_78526_ _78522_/Y _78526_/B _78526_/C _78528_/A sky130_fd_sc_hd__or3_4
X_44918_ _80672_/Q _45153_/A sky130_fd_sc_hd__buf_2
X_63752_ _63751_/X _64177_/D sky130_fd_sc_hd__buf_2
X_75738_ _75727_/A _75726_/Y _75737_/X _75738_/Y sky130_fd_sc_hd__a21oi_4
X_48686_ _81764_/Q _48687_/A sky130_fd_sc_hd__inv_2
X_60964_ _60901_/B _60993_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_611_0_CLK clkbuf_9_305_0_CLK/X _80835_/CLK sky130_fd_sc_hd__clkbuf_1
X_45898_ _45897_/X _45898_/X sky130_fd_sc_hd__buf_2
X_62703_ _61376_/X _62694_/B _62694_/C _62664_/D _62703_/Y sky130_fd_sc_hd__nand4_4
X_47637_ _47655_/A _47645_/B _47614_/X _53159_/D _47637_/X sky130_fd_sc_hd__and4_4
X_66471_ _66216_/A _66397_/X _66216_/C _66471_/Y sky130_fd_sc_hd__nand3_4
X_78457_ _82797_/Q _78461_/A sky130_fd_sc_hd__inv_2
X_44849_ _45964_/A _44849_/X sky130_fd_sc_hd__buf_2
X_75669_ _75669_/A _75669_/B _75669_/Y sky130_fd_sc_hd__xnor2_4
X_63683_ _59436_/Y _63626_/X _61666_/A _63627_/X _63683_/X sky130_fd_sc_hd__a2bb2o_4
X_60895_ _60894_/X _60895_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_102_0_CLK clkbuf_8_51_0_CLK/X clkbuf_9_102_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_68210_ _67298_/X _67301_/X _68209_/X _68210_/Y sky130_fd_sc_hd__a21oi_4
X_65422_ _65420_/Y _65347_/X _65421_/X _84202_/D sky130_fd_sc_hd__a21o_4
X_77408_ _82223_/Q _77412_/A sky130_fd_sc_hd__inv_2
X_62634_ _62634_/A _62634_/B _62634_/C _62633_/Y _62634_/Y sky130_fd_sc_hd__nand4_4
X_69190_ _69190_/A _69191_/A sky130_fd_sc_hd__buf_2
X_47568_ _47530_/X _47595_/B _47595_/C _53125_/D _47568_/X sky130_fd_sc_hd__and4_4
X_78388_ _78384_/Y _78386_/Y _78387_/Y _78394_/A sky130_fd_sc_hd__o21ai_4
X_49307_ _65124_/B _49300_/X _49306_/Y _49307_/Y sky130_fd_sc_hd__o21ai_4
X_68141_ _66891_/X _66893_/X _68133_/X _68141_/Y sky130_fd_sc_hd__a21oi_4
X_46519_ _83785_/Q _54058_/B sky130_fd_sc_hd__inv_2
X_65353_ _65350_/X _86148_/Q _65224_/X _65352_/X _65353_/X sky130_fd_sc_hd__a211o_4
X_77339_ _77339_/A _77339_/B _77339_/X sky130_fd_sc_hd__or2_4
Xclkbuf_10_626_0_CLK clkbuf_9_313_0_CLK/X _80961_/CLK sky130_fd_sc_hd__clkbuf_1
X_62565_ _62487_/X _58187_/X _62565_/C _62608_/D _62565_/X sky130_fd_sc_hd__and4_4
X_47499_ _47517_/A _53080_/B _47499_/Y sky130_fd_sc_hd__nand2_4
X_64304_ _64304_/A _64303_/X _84961_/Q _64304_/D _64304_/X sky130_fd_sc_hd__and4_4
X_61516_ _61509_/Y _61511_/Y _61464_/X _61513_/Y _61515_/Y _61516_/X
+ sky130_fd_sc_hd__a41o_4
X_49238_ _64784_/B _49222_/X _49237_/Y _49238_/Y sky130_fd_sc_hd__o21ai_4
X_80350_ _80350_/A _80350_/B _80350_/C _80353_/A sky130_fd_sc_hd__nand3_4
X_68072_ _87444_/Q _68069_/X _68070_/X _68071_/X _68072_/X sky130_fd_sc_hd__a211o_4
X_65284_ _65158_/A _65285_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_117_0_CLK clkbuf_8_58_0_CLK/X clkbuf_9_117_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_62496_ _61558_/B _62462_/X _62436_/X _62478_/X _62495_/X _62496_/X
+ sky130_fd_sc_hd__a41o_4
Xclkbuf_9_44_0_CLK clkbuf_8_22_0_CLK/X clkbuf_9_44_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_67023_ _67023_/A _67023_/B _67023_/X sky130_fd_sc_hd__and2_4
X_79009_ _78993_/B _79006_/X _79008_/Y _79010_/B sky130_fd_sc_hd__a21oi_4
X_64235_ _64223_/A _64235_/B _64223_/C _64235_/X sky130_fd_sc_hd__and3_4
X_49169_ _86437_/Q _49153_/X _49168_/Y _49169_/Y sky130_fd_sc_hd__o21ai_4
X_61447_ _61437_/A _61447_/B _61398_/C _61447_/Y sky130_fd_sc_hd__nand3_4
X_80281_ _84747_/Q _84139_/Q _80281_/Y sky130_fd_sc_hd__nor2_4
X_51200_ _86055_/Q _51183_/X _51199_/Y _51200_/Y sky130_fd_sc_hd__o21ai_4
X_82020_ _82104_/CLK _77754_/B _81988_/D sky130_fd_sc_hd__dfxtp_4
X_52180_ _52210_/A _48540_/B _52180_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_3_2_0_CLK clkbuf_3_3_0_CLK/A clkbuf_3_2_1_CLK/A sky130_fd_sc_hd__clkbuf_1
X_64166_ _61676_/A _64177_/B _64189_/D _64177_/D _64166_/Y sky130_fd_sc_hd__nand4_4
X_61378_ _61378_/A _61367_/B _61367_/C _61367_/D _61378_/Y sky130_fd_sc_hd__nand4_4
X_51131_ _86068_/Q _51128_/X _51130_/Y _51131_/Y sky130_fd_sc_hd__o21ai_4
X_63117_ _60523_/A _63117_/X sky130_fd_sc_hd__buf_2
X_60329_ _57757_/A _65296_/A sky130_fd_sc_hd__buf_2
X_68974_ _80809_/D _68954_/X _68973_/X _83953_/D sky130_fd_sc_hd__a21bo_4
X_64097_ _63733_/X _64173_/C sky130_fd_sc_hd__buf_2
Xclkbuf_9_59_0_CLK clkbuf_9_59_0_CLK/A clkbuf_9_59_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_51062_ _51059_/Y _51039_/X _51061_/X _51062_/Y sky130_fd_sc_hd__a21oi_4
X_67925_ _68120_/A _67925_/X sky130_fd_sc_hd__buf_2
X_63048_ _60466_/X _63085_/C sky130_fd_sc_hd__buf_2
X_83971_ _80931_/CLK _83971_/D _80827_/D sky130_fd_sc_hd__dfxtp_4
X_50013_ _48171_/X _50027_/A sky130_fd_sc_hd__buf_2
X_85710_ _82390_/CLK _53032_/Y _85710_/Q sky130_fd_sc_hd__dfxtp_4
X_82922_ _82931_/CLK _78189_/X _82922_/Q sky130_fd_sc_hd__dfxtp_4
X_67856_ _67955_/A _67856_/B _67856_/X sky130_fd_sc_hd__and2_4
X_55870_ _44081_/X _55870_/B _55870_/X sky130_fd_sc_hd__and2_4
X_86690_ _86372_/CLK _86690_/D _86690_/Q sky130_fd_sc_hd__dfxtp_4
X_54821_ _54825_/A _54843_/B _54831_/C _53129_/D _54821_/X sky130_fd_sc_hd__and4_4
X_85641_ _85738_/CLK _85641_/D _85641_/Q sky130_fd_sc_hd__dfxtp_4
X_66807_ _69245_/A _66807_/X sky130_fd_sc_hd__buf_2
X_82853_ _82299_/CLK _78103_/B _82853_/Q sky130_fd_sc_hd__dfxtp_4
X_67787_ _67784_/X _67786_/X _67742_/X _67792_/A sky130_fd_sc_hd__a21o_4
X_64999_ _64817_/A _64999_/X sky130_fd_sc_hd__buf_2
X_57540_ _57538_/Y _57515_/X _57539_/Y _84983_/D sky130_fd_sc_hd__a21boi_4
X_81804_ _81362_/CLK _81612_/Q _81804_/Q sky130_fd_sc_hd__dfxtp_4
X_69526_ _69612_/A _69526_/B _69526_/X sky130_fd_sc_hd__and2_4
X_88360_ _88363_/CLK _40653_/X _68645_/B sky130_fd_sc_hd__dfxtp_4
X_54752_ _54344_/A _54807_/A sky130_fd_sc_hd__buf_2
X_66738_ _66664_/X _86831_/Q _66738_/X sky130_fd_sc_hd__and2_4
X_85572_ _83564_/CLK _85572_/D _85572_/Q sky130_fd_sc_hd__dfxtp_4
X_51964_ _51941_/A _48207_/X _51964_/Y sky130_fd_sc_hd__nand2_4
X_82784_ _82973_/CLK _78784_/Y _82784_/Q sky130_fd_sc_hd__dfxtp_4
X_87311_ _88327_/CLK _87311_/D _87311_/Q sky130_fd_sc_hd__dfxtp_4
X_53703_ _52182_/A _53720_/B _53734_/C _53703_/X sky130_fd_sc_hd__and3_4
X_84523_ _84287_/CLK _61062_/Y _76971_/A sky130_fd_sc_hd__dfxtp_4
X_50915_ _50913_/Y _50902_/X _50914_/X _50915_/Y sky130_fd_sc_hd__a21oi_4
X_81735_ _86807_/CLK _75955_/B _41427_/A sky130_fd_sc_hd__dfxtp_4
X_57471_ _57372_/X _57469_/X _57470_/Y _57472_/A sky130_fd_sc_hd__o21ai_4
X_69457_ _69457_/A _69457_/X sky130_fd_sc_hd__buf_2
X_88291_ _87022_/CLK _41029_/X _69362_/B sky130_fd_sc_hd__dfxtp_4
X_54683_ _85397_/Q _54676_/X _54682_/Y _54683_/Y sky130_fd_sc_hd__o21ai_4
X_66669_ _66669_/A _88207_/Q _66669_/X sky130_fd_sc_hd__and2_4
X_51895_ _51875_/A _51031_/B _51895_/Y sky130_fd_sc_hd__nand2_4
X_59210_ _59208_/X _86064_/Q _59209_/X _59210_/Y sky130_fd_sc_hd__o21ai_4
X_56422_ _56435_/A _56431_/A sky130_fd_sc_hd__buf_2
X_68408_ _67657_/X _68409_/A sky130_fd_sc_hd__buf_2
X_87242_ _88012_/CLK _43836_/X _68604_/B sky130_fd_sc_hd__dfxtp_4
X_53634_ _85598_/Q _53626_/X _53633_/Y _53634_/Y sky130_fd_sc_hd__o21ai_4
X_84454_ _84454_/CLK _61785_/Y _78077_/B sky130_fd_sc_hd__dfxtp_4
X_50846_ _50843_/Y _50792_/X _50845_/Y _86122_/D sky130_fd_sc_hd__a21boi_4
X_81666_ _81040_/CLK _80264_/Y _81666_/Q sky130_fd_sc_hd__dfxtp_4
X_69388_ _87021_/Q _69239_/X _69361_/X _69387_/X _69388_/X sky130_fd_sc_hd__a211o_4
X_59141_ _59137_/Y _59139_/Y _59140_/X _59141_/X sky130_fd_sc_hd__a21o_4
X_83405_ _83491_/CLK _83405_/D _83405_/Q sky130_fd_sc_hd__dfxtp_4
X_56353_ _56139_/X _56350_/X _56352_/Y _56353_/Y sky130_fd_sc_hd__o21ai_4
X_80617_ _80617_/A _80607_/X _80617_/Y sky130_fd_sc_hd__nand2_4
X_68339_ _68082_/X _68084_/X _68327_/X _68339_/Y sky130_fd_sc_hd__a21oi_4
X_87173_ _87169_/CLK _44289_/X _44072_/A sky130_fd_sc_hd__dfxtp_4
X_53565_ _53565_/A _48297_/X _53565_/Y sky130_fd_sc_hd__nand2_4
X_84385_ _84518_/CLK _62758_/Y _75915_/B sky130_fd_sc_hd__dfxtp_4
X_50777_ _50777_/A _50777_/B _50777_/Y sky130_fd_sc_hd__nand2_4
X_81597_ _81433_/CLK _84197_/Q _81597_/Q sky130_fd_sc_hd__dfxtp_4
X_55304_ _85039_/Q _44060_/X _55301_/X _55303_/X _55304_/X sky130_fd_sc_hd__a211o_4
X_86124_ _86040_/CLK _86124_/D _86124_/Q sky130_fd_sc_hd__dfxtp_4
X_40530_ _40368_/X _40530_/B _40530_/X sky130_fd_sc_hd__or2_4
X_52516_ _52515_/X _52516_/X sky130_fd_sc_hd__buf_2
X_71350_ _71344_/X _83529_/Q _71349_/X _83529_/D sky130_fd_sc_hd__a21o_4
X_59072_ _59033_/X _85435_/Q _59071_/X _59072_/Y sky130_fd_sc_hd__o21ai_4
X_83336_ _83333_/CLK _83336_/D _83336_/Q sky130_fd_sc_hd__dfxtp_4
X_80548_ _80548_/A _84322_/Q _80549_/B sky130_fd_sc_hd__xor2_4
X_56284_ _56350_/A _56284_/X sky130_fd_sc_hd__buf_2
X_53496_ _85625_/Q _53476_/X _53495_/Y _53496_/Y sky130_fd_sc_hd__o21ai_4
X_58023_ _58019_/Y _58022_/Y _57909_/X _58023_/X sky130_fd_sc_hd__a21o_4
X_70301_ _70296_/X _70297_/X _70301_/C _70301_/D _70301_/X sky130_fd_sc_hd__and4_4
X_55235_ _55235_/A _56898_/A _55235_/X sky130_fd_sc_hd__and2_4
X_86055_ _85735_/CLK _51204_/Y _86055_/Q sky130_fd_sc_hd__dfxtp_4
X_40461_ _40461_/A _40461_/Y sky130_fd_sc_hd__inv_2
X_52447_ _52445_/Y _52415_/X _52446_/X _85821_/D sky130_fd_sc_hd__a21oi_4
X_71281_ _71181_/A _71268_/A _71279_/C _71276_/D _71281_/Y sky130_fd_sc_hd__nand4_4
X_83267_ _85332_/CLK _83267_/D _83267_/Q sky130_fd_sc_hd__dfxtp_4
X_80479_ _80471_/B _80471_/A _80478_/X _80480_/B sky130_fd_sc_hd__a21boi_4
X_42200_ _42199_/X _42200_/X sky130_fd_sc_hd__buf_2
X_73020_ _73021_/B _73021_/C _73019_/X _73020_/X sky130_fd_sc_hd__a21o_4
X_85006_ _85034_/CLK _85006_/D _55317_/B sky130_fd_sc_hd__dfxtp_4
X_70232_ _70232_/A _70239_/B sky130_fd_sc_hd__buf_2
X_82218_ _81928_/CLK _82250_/Q _77339_/A sky130_fd_sc_hd__dfxtp_4
X_43180_ _43180_/A _43180_/X sky130_fd_sc_hd__buf_2
X_55166_ _55159_/A _85068_/Q _55166_/X sky130_fd_sc_hd__and2_4
X_40392_ _40391_/X _40342_/X _88399_/Q _40355_/X _40392_/X sky130_fd_sc_hd__a2bb2o_4
X_52378_ _52375_/Y _52364_/X _52377_/X _52378_/Y sky130_fd_sc_hd__a21oi_4
X_83198_ _85049_/CLK _83198_/D _70205_/C sky130_fd_sc_hd__dfxtp_4
X_42131_ _42120_/X _42116_/X _41116_/X _88019_/Q _42117_/X _42132_/A
+ sky130_fd_sc_hd__o32ai_4
X_54117_ _53436_/X _54117_/X sky130_fd_sc_hd__buf_2
X_51329_ _65105_/B _51309_/X _51328_/Y _51329_/Y sky130_fd_sc_hd__o21ai_4
X_70163_ _70134_/X _70348_/D sky130_fd_sc_hd__buf_2
X_82149_ _82746_/CLK _66319_/C _82149_/Q sky130_fd_sc_hd__dfxtp_4
X_55097_ _55094_/Y _55076_/X _55096_/X _55097_/Y sky130_fd_sc_hd__a21oi_4
X_59974_ _59995_/A _62621_/D _59950_/B _59977_/B _59974_/Y sky130_fd_sc_hd__nand4_4
X_42062_ _42060_/X _42049_/X _40925_/X _42061_/Y _41872_/X _42062_/Y
+ sky130_fd_sc_hd__o32ai_4
X_58925_ _59033_/A _58925_/X sky130_fd_sc_hd__buf_2
X_54048_ _54046_/Y _54015_/X _54047_/X _85516_/D sky130_fd_sc_hd__a21oi_4
X_74971_ _74971_/A _74971_/B _74972_/B sky130_fd_sc_hd__and2_4
X_70094_ _82531_/D _70085_/X _70093_/X _70094_/X sky130_fd_sc_hd__a21bo_4
X_86957_ _88224_/CLK _44783_/Y _86957_/Q sky130_fd_sc_hd__dfxtp_4
X_41013_ _41013_/A _41019_/B sky130_fd_sc_hd__buf_2
X_76710_ _76697_/Y _76704_/Y _76710_/Y sky130_fd_sc_hd__nor2_4
X_73922_ _43068_/Y _72888_/X _73920_/X _73921_/Y _73922_/X sky130_fd_sc_hd__a211o_4
X_85908_ _86549_/CLK _85908_/D _66094_/B sky130_fd_sc_hd__dfxtp_4
X_46870_ _83662_/Q _52722_/B sky130_fd_sc_hd__inv_2
X_58856_ _84794_/Q _58856_/Y sky130_fd_sc_hd__inv_2
X_77690_ _77687_/Y _77690_/B _77688_/Y _77690_/Y sky130_fd_sc_hd__nand3_4
X_86888_ _86861_/CLK _45262_/Y _62544_/A sky130_fd_sc_hd__dfxtp_4
X_45821_ _45819_/X _61655_/A _45765_/X _45821_/Y sky130_fd_sc_hd__o21ai_4
X_57807_ _57806_/X _86332_/Q _57807_/Y sky130_fd_sc_hd__nor2_4
X_76641_ _76639_/Y _76640_/Y _76643_/A sky130_fd_sc_hd__nand2_4
X_73853_ _73850_/X _86229_/Q _73804_/X _73852_/X _73853_/X sky130_fd_sc_hd__a211o_4
X_85839_ _86256_/CLK _85839_/D _85839_/Q sky130_fd_sc_hd__dfxtp_4
X_58787_ _59061_/A _58787_/X sky130_fd_sc_hd__buf_2
X_55999_ _55997_/X _74312_/C _55928_/B _55928_/C _55999_/X sky130_fd_sc_hd__and4_4
X_48540_ _48604_/A _48540_/B _48540_/Y sky130_fd_sc_hd__nand2_4
X_72804_ _69597_/B _72803_/X _72776_/X _72804_/Y sky130_fd_sc_hd__o21ai_4
X_79360_ _79351_/X _79360_/B _79360_/Y sky130_fd_sc_hd__nand2_4
X_45752_ _85098_/Q _45752_/Y sky130_fd_sc_hd__inv_2
X_57738_ _46224_/X _85407_/Q _57737_/X _57738_/Y sky130_fd_sc_hd__o21ai_4
X_76572_ _76572_/A _76572_/Y sky130_fd_sc_hd__inv_2
X_42964_ _40404_/X _42962_/X _87628_/Q _42963_/X _42964_/X sky130_fd_sc_hd__a2bb2o_4
X_73784_ _73735_/X _85624_/Q _73782_/X _73783_/X _73784_/X sky130_fd_sc_hd__a211o_4
X_70996_ _51328_/B _70983_/X _70995_/Y _70996_/Y sky130_fd_sc_hd__o21ai_4
X_78311_ _78308_/Y _78310_/Y _78311_/Y sky130_fd_sc_hd__nor2_4
X_44703_ _44679_/X _44680_/X _40667_/X _86993_/Q _44681_/X _44704_/A
+ sky130_fd_sc_hd__o32ai_4
X_75523_ _75519_/X _75520_/Y _75524_/B _75523_/X sky130_fd_sc_hd__a21o_4
X_87509_ _87790_/CLK _87509_/D _87509_/Q sky130_fd_sc_hd__dfxtp_4
X_41915_ _41887_/X _41888_/X _40633_/X _41914_/Y _41891_/X _88107_/D
+ sky130_fd_sc_hd__o32ai_4
X_72735_ _73262_/A _72735_/X sky130_fd_sc_hd__buf_2
X_48471_ _48471_/A _48471_/X sky130_fd_sc_hd__buf_2
X_79291_ _79291_/A _79297_/A sky130_fd_sc_hd__inv_2
X_45683_ _45680_/X _45682_/Y _45561_/X _45683_/Y sky130_fd_sc_hd__a21oi_4
X_57669_ _84957_/Q _57670_/A sky130_fd_sc_hd__buf_2
X_42895_ _42846_/X _42895_/X sky130_fd_sc_hd__buf_2
X_47422_ _47404_/A _53041_/B _47422_/Y sky130_fd_sc_hd__nand2_4
X_59408_ _59394_/X _83485_/Q _59407_/Y _84741_/D sky130_fd_sc_hd__o21a_4
X_78242_ _78241_/A _78241_/B _78252_/C sky130_fd_sc_hd__nand2_4
X_44634_ _44622_/X _44623_/X _41021_/A _87024_/Q _44625_/X _44634_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75454_ _80700_/Q _80956_/D _75457_/B sky130_fd_sc_hd__nor2_4
X_41846_ _41846_/A _88125_/D sky130_fd_sc_hd__inv_2
X_60680_ _63630_/B _60732_/C sky130_fd_sc_hd__buf_2
X_72666_ _72668_/A _72668_/B _55503_/D _72666_/Y sky130_fd_sc_hd__nand3_4
X_74405_ _74492_/A _74405_/X sky130_fd_sc_hd__buf_2
X_47353_ _47333_/X _52999_/B _47353_/Y sky130_fd_sc_hd__nand2_4
X_59339_ _59043_/A _59339_/X sky130_fd_sc_hd__buf_2
X_71617_ _71604_/X _83437_/Q _71616_/Y _83437_/D sky130_fd_sc_hd__a21o_4
X_78173_ _78173_/A _78173_/B _78173_/X sky130_fd_sc_hd__xor2_4
X_44565_ _44547_/A _44565_/X sky130_fd_sc_hd__buf_2
X_75385_ _75384_/X _75386_/B sky130_fd_sc_hd__inv_2
X_41777_ _40621_/X _41435_/A _41776_/X _41777_/Y sky130_fd_sc_hd__o21ai_4
X_72597_ _72528_/Y _72597_/B _72597_/C _72597_/Y sky130_fd_sc_hd__nand3_4
X_46304_ _46301_/X _82941_/Q _46303_/Y _53964_/A sky130_fd_sc_hd__o21ai_4
X_77124_ _77143_/B _81916_/Q _77141_/A sky130_fd_sc_hd__xor2_4
X_43516_ _43495_/X _43503_/X _41786_/X _87381_/Q _43506_/X _43516_/Y
+ sky130_fd_sc_hd__o32ai_4
X_62350_ _61438_/X _62309_/B _62309_/C _62225_/X _62351_/D sky130_fd_sc_hd__nand4_4
X_74336_ _74338_/A _74338_/B _55811_/X _74336_/Y sky130_fd_sc_hd__nand3_4
X_40728_ _40670_/X _40897_/A _40727_/X _40729_/A sky130_fd_sc_hd__o21ai_4
X_47284_ _47246_/X _47311_/B _47321_/C _52963_/D _47284_/X sky130_fd_sc_hd__and4_4
X_71548_ _71411_/A _71546_/B _71536_/A _71548_/Y sky130_fd_sc_hd__nor3_4
X_44496_ _44547_/A _44496_/X sky130_fd_sc_hd__buf_2
X_49023_ _49017_/Y _48985_/X _49022_/X _49023_/Y sky130_fd_sc_hd__a21oi_4
X_61301_ _84857_/Q _61301_/X sky130_fd_sc_hd__buf_2
X_46235_ _46234_/Y _56777_/B sky130_fd_sc_hd__buf_2
XPHY_470 sky130_fd_sc_hd__decap_3
X_77055_ _77047_/B _77055_/B _77055_/Y sky130_fd_sc_hd__nor2_4
X_43447_ _43397_/A _43447_/X sky130_fd_sc_hd__buf_2
X_62281_ _61375_/B _62278_/X _60027_/A _60011_/X _62280_/X _62281_/X
+ sky130_fd_sc_hd__a41o_4
X_74267_ _69114_/B _73124_/B _73920_/X _74266_/Y _74267_/X sky130_fd_sc_hd__a211o_4
XPHY_481 sky130_fd_sc_hd__decap_3
X_40659_ _40659_/A _40654_/B _40659_/X sky130_fd_sc_hd__or2_4
X_71479_ _71827_/A _71479_/B _71435_/C _71716_/D _71479_/X sky130_fd_sc_hd__and4_4
XPHY_492 sky130_fd_sc_hd__decap_3
X_64020_ _64053_/A _58438_/A _64071_/C _64020_/X sky130_fd_sc_hd__and3_4
X_76006_ _75994_/Y _76006_/B _76009_/A sky130_fd_sc_hd__nand2_4
X_61232_ _64223_/A _61232_/X sky130_fd_sc_hd__buf_2
X_73218_ _48550_/Y _73217_/Y _73218_/X sky130_fd_sc_hd__xor2_4
X_46166_ _46166_/A _45886_/X _46166_/C _46167_/A sky130_fd_sc_hd__and3_4
X_43378_ _43329_/X _43378_/X sky130_fd_sc_hd__buf_2
X_74198_ _74155_/X _84966_/Q _72992_/X _74197_/X _74198_/X sky130_fd_sc_hd__a211o_4
X_45117_ _55857_/B _45060_/X _45116_/X _45117_/X sky130_fd_sc_hd__o21a_4
X_42329_ _43161_/A _42417_/A sky130_fd_sc_hd__buf_2
X_61163_ _61095_/X _61109_/X _59691_/X _61163_/Y sky130_fd_sc_hd__a21oi_4
X_73149_ _73149_/A _72896_/B _73149_/Y sky130_fd_sc_hd__nor2_4
X_46097_ _46097_/A _46098_/A sky130_fd_sc_hd__buf_2
X_60114_ _60125_/A _60103_/B _84659_/Q _60114_/Y sky130_fd_sc_hd__nor3_4
X_49925_ _49925_/A _49925_/X sky130_fd_sc_hd__buf_2
X_45048_ _45046_/Y _45067_/B _45048_/Y sky130_fd_sc_hd__nand2_4
X_65971_ _65968_/Y _65915_/X _65970_/X _84165_/D sky130_fd_sc_hd__a21o_4
X_61094_ _61107_/A _61153_/A sky130_fd_sc_hd__buf_2
X_77957_ _77957_/A _77956_/Y _77958_/B sky130_fd_sc_hd__xnor2_4
X_67710_ _67705_/X _67708_/X _67709_/X _67710_/Y sky130_fd_sc_hd__a21oi_4
X_64922_ _64917_/X _64921_/X _64851_/X _64926_/A sky130_fd_sc_hd__a21o_4
X_76908_ _76906_/Y _76934_/A _76931_/A sky130_fd_sc_hd__xor2_4
X_60045_ _60058_/B _60079_/B _60027_/X _60045_/Y sky130_fd_sc_hd__nand3_4
X_49856_ _58070_/B _49853_/X _49855_/Y _49856_/Y sky130_fd_sc_hd__o21ai_4
X_68690_ _80821_/D _68586_/X _68689_/X _68690_/X sky130_fd_sc_hd__a21bo_4
X_77888_ _82163_/Q _77888_/B _82131_/D sky130_fd_sc_hd__xor2_4
X_48807_ _47832_/X _48808_/A sky130_fd_sc_hd__buf_2
X_67641_ _67997_/A _67641_/X sky130_fd_sc_hd__buf_2
X_79627_ _79626_/Y _79627_/Y sky130_fd_sc_hd__inv_2
X_64853_ _64773_/A _86456_/Q _64853_/X sky130_fd_sc_hd__and2_4
X_76839_ _76839_/A _76841_/A sky130_fd_sc_hd__inv_2
X_49787_ _49787_/A _49787_/X sky130_fd_sc_hd__buf_2
X_46999_ _46999_/A _52797_/D sky130_fd_sc_hd__buf_2
Xclkbuf_10_550_0_CLK clkbuf_9_275_0_CLK/X _81746_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_41_0_CLK clkbuf_6_41_0_CLK/A clkbuf_7_83_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_63804_ _63410_/B _63820_/B _63753_/C _63820_/D _63804_/Y sky130_fd_sc_hd__nand4_4
X_48738_ _72911_/B _48730_/X _48737_/Y _48738_/Y sky130_fd_sc_hd__o21ai_4
X_67572_ _67572_/A _86933_/Q _67572_/X sky130_fd_sc_hd__and2_4
X_79558_ _79558_/A _79558_/B _79558_/Y sky130_fd_sc_hd__nand2_4
X_64784_ _64810_/A _64784_/B _64784_/X sky130_fd_sc_hd__and2_4
X_61996_ _61538_/B _61995_/X _61953_/C _61937_/X _62000_/C sky130_fd_sc_hd__nand4_4
X_69311_ _69307_/X _69310_/X _69171_/X _69311_/Y sky130_fd_sc_hd__a21oi_4
X_66523_ _65464_/A _66524_/B sky130_fd_sc_hd__buf_2
X_78509_ _78505_/X _78510_/C _78508_/Y _78511_/A sky130_fd_sc_hd__a21o_4
X_63735_ _63735_/A _64136_/B sky130_fd_sc_hd__buf_2
X_48669_ _48612_/A _48669_/X sky130_fd_sc_hd__buf_2
X_60947_ _60946_/X _60838_/X _60947_/C _60947_/Y sky130_fd_sc_hd__nor3_4
X_79489_ _79489_/A _79488_/Y _82846_/D sky130_fd_sc_hd__xor2_4
X_50700_ _50695_/A _50183_/B _50700_/Y sky130_fd_sc_hd__nand2_4
X_81520_ _88175_/CLK _81564_/Q _76025_/A sky130_fd_sc_hd__dfxtp_4
X_69242_ _69238_/X _69241_/X _69142_/X _69242_/Y sky130_fd_sc_hd__a21oi_4
X_66454_ _65053_/X _66423_/B _65055_/X _66454_/Y sky130_fd_sc_hd__nand3_4
X_51680_ _51678_/Y _51667_/X _51679_/X _85966_/D sky130_fd_sc_hd__a21oi_4
X_63666_ _58194_/A _60798_/X _63384_/C _60703_/Y _62129_/X _63666_/X
+ sky130_fd_sc_hd__a32o_4
Xclkbuf_10_565_0_CLK clkbuf_9_282_0_CLK/X _82067_/CLK sky130_fd_sc_hd__clkbuf_1
X_60878_ _60853_/X _60879_/D sky130_fd_sc_hd__buf_2
Xclkbuf_6_56_0_CLK clkbuf_6_57_0_CLK/A clkbuf_6_56_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_65405_ _65402_/X _65404_/X _65277_/X _65410_/A sky130_fd_sc_hd__a21o_4
X_50631_ _50629_/Y _50619_/X _50630_/Y _50631_/Y sky130_fd_sc_hd__a21boi_4
X_62617_ _62615_/Y _62593_/X _62616_/Y _62617_/Y sky130_fd_sc_hd__a21oi_4
X_81451_ _84049_/CLK _76733_/B _81451_/Q sky130_fd_sc_hd__dfxtp_4
X_69173_ _68430_/X _68432_/X _69061_/X _69173_/Y sky130_fd_sc_hd__a21oi_4
X_66385_ _64747_/X _66385_/B _64750_/X _66385_/Y sky130_fd_sc_hd__nand3_4
X_63597_ _63657_/A _62027_/X _63597_/X sky130_fd_sc_hd__and2_4
X_80402_ _80416_/A _80416_/B _80425_/A sky130_fd_sc_hd__xor2_4
X_68124_ _82073_/D _68120_/X _68123_/X _84033_/D sky130_fd_sc_hd__a21bo_4
X_53350_ _48755_/A _53351_/A sky130_fd_sc_hd__buf_2
X_65336_ _65334_/X _86117_/Q _65256_/X _65335_/X _65336_/X sky130_fd_sc_hd__a211o_4
X_84170_ _82748_/CLK _84170_/D _65901_/C sky130_fd_sc_hd__dfxtp_4
X_50562_ _50559_/Y _50551_/X _50561_/X _86177_/D sky130_fd_sc_hd__a21oi_4
X_62548_ _61609_/X _62548_/B _62548_/C _62548_/D _62548_/Y sky130_fd_sc_hd__nand4_4
X_81382_ _84087_/CLK _81382_/D _76828_/B sky130_fd_sc_hd__dfxtp_4
X_52301_ _50599_/A _50599_/B _52280_/X _52301_/X sky130_fd_sc_hd__o21a_4
X_83121_ _86213_/CLK _83121_/D _70128_/C sky130_fd_sc_hd__dfxtp_4
Xpsn_inst_psn_buff_9 _44195_/Y _44196_/D sky130_fd_sc_hd__buf_8
X_80333_ _80315_/A _80313_/Y _80332_/Y _80333_/Y sky130_fd_sc_hd__a21oi_4
X_68055_ _87381_/Q _67987_/X _68053_/X _68054_/X _68055_/X sky130_fd_sc_hd__a211o_4
X_53281_ _85662_/Q _53268_/X _53280_/Y _53281_/Y sky130_fd_sc_hd__o21ai_4
X_65267_ _65198_/X _65255_/Y _65266_/Y _65267_/Y sky130_fd_sc_hd__o21ai_4
X_50493_ _50490_/Y _50491_/X _50492_/X _86190_/D sky130_fd_sc_hd__a21oi_4
X_62479_ _62479_/A _63585_/B _62479_/C _62463_/X _62479_/X sky130_fd_sc_hd__and4_4
X_55020_ _55072_/A _55020_/X sky130_fd_sc_hd__buf_2
X_67006_ _67057_/A _87681_/Q _67006_/X sky130_fd_sc_hd__and2_4
X_52232_ _52203_/A _52232_/X sky130_fd_sc_hd__buf_2
X_64218_ _64315_/A _64219_/B sky130_fd_sc_hd__buf_2
X_83052_ _85566_/CLK _74506_/Y _83052_/Q sky130_fd_sc_hd__dfxtp_4
X_80264_ _80264_/A _80264_/B _80264_/Y sky130_fd_sc_hd__xnor2_4
X_65198_ _65198_/A _65198_/X sky130_fd_sc_hd__buf_2
X_82003_ _82008_/CLK _82035_/Q _77127_/A sky130_fd_sc_hd__dfxtp_4
X_52163_ _52168_/A _52163_/B _52163_/Y sky130_fd_sc_hd__nand2_4
X_64149_ _62140_/X _64182_/B _64095_/C _64095_/D _64149_/Y sky130_fd_sc_hd__nand4_4
X_87860_ _87348_/CLK _42444_/X _87860_/Q sky130_fd_sc_hd__dfxtp_4
X_80195_ _80195_/A _84292_/Q _80195_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_10_503_0_CLK clkbuf_9_251_0_CLK/X _85459_/CLK sky130_fd_sc_hd__clkbuf_1
X_51114_ _51141_/A _51115_/C sky130_fd_sc_hd__buf_2
X_86811_ _81154_/CLK _46019_/X _67215_/B sky130_fd_sc_hd__dfxtp_4
X_52094_ _52092_/Y _52049_/X _52093_/X _85890_/D sky130_fd_sc_hd__a21oi_4
X_56971_ _58547_/A _56971_/B _56971_/C _56971_/Y sky130_fd_sc_hd__nor3_4
X_68957_ _74121_/A _68883_/X _68884_/X _68956_/Y _68957_/X sky130_fd_sc_hd__a211o_4
X_87791_ _87544_/CLK _87791_/D _87791_/Q sky130_fd_sc_hd__dfxtp_4
X_58710_ _84806_/Q _58599_/X _58702_/X _58709_/X _58710_/Y sky130_fd_sc_hd__a2bb2oi_4
X_51045_ _51029_/A _51045_/B _51045_/C _52735_/D _51045_/X sky130_fd_sc_hd__and4_4
X_55922_ _56395_/C _44070_/B _55627_/X _55921_/X _55922_/X sky130_fd_sc_hd__a211o_4
X_86742_ _85527_/CLK _46384_/Y _86742_/Q sky130_fd_sc_hd__dfxtp_4
X_67908_ _69797_/A _67908_/X sky130_fd_sc_hd__buf_2
X_59690_ _59801_/A _59816_/A sky130_fd_sc_hd__buf_2
X_83954_ _80821_/CLK _83954_/D _83954_/Q sky130_fd_sc_hd__dfxtp_4
X_68888_ _68746_/A _68888_/B _68888_/Y sky130_fd_sc_hd__nor2_4
X_58641_ _58641_/A _58641_/X sky130_fd_sc_hd__buf_2
X_82905_ _82906_/CLK _78247_/B _41674_/A sky130_fd_sc_hd__dfxtp_4
X_55853_ _55850_/X _55853_/B _55853_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_518_0_CLK clkbuf_9_259_0_CLK/X _81482_/CLK sky130_fd_sc_hd__clkbuf_1
X_67839_ _68644_/A _67909_/A sky130_fd_sc_hd__buf_2
X_86673_ _86353_/CLK _86673_/D _86673_/Q sky130_fd_sc_hd__dfxtp_4
X_83885_ _82301_/CLK _83885_/D _81957_/D sky130_fd_sc_hd__dfxtp_4
X_54804_ _54801_/Y _54802_/X _54803_/X _85375_/D sky130_fd_sc_hd__a21oi_4
X_85624_ _86235_/CLK _85624_/D _85624_/Q sky130_fd_sc_hd__dfxtp_4
X_70850_ _51779_/B _70830_/Y _70849_/Y _70850_/Y sky130_fd_sc_hd__o21ai_4
X_58572_ _58571_/X _85793_/Q _58089_/X _58572_/X sky130_fd_sc_hd__o21a_4
X_82836_ _84177_/CLK _82836_/D _82836_/Q sky130_fd_sc_hd__dfxtp_4
X_55784_ _56250_/C _55747_/X _55165_/X _55783_/X _55784_/X sky130_fd_sc_hd__a211o_4
X_52996_ _85716_/Q _52984_/X _52995_/Y _52996_/Y sky130_fd_sc_hd__o21ai_4
X_57523_ _47819_/A _57523_/B _57523_/Y sky130_fd_sc_hd__nand2_4
X_69509_ _69454_/A _69509_/B _69509_/X sky130_fd_sc_hd__and2_4
X_88343_ _87850_/CLK _88343_/D _88343_/Q sky130_fd_sc_hd__dfxtp_4
X_54735_ _54733_/Y _54720_/X _54734_/X _54735_/Y sky130_fd_sc_hd__a21oi_4
X_85555_ _85555_/CLK _53855_/Y _85555_/Q sky130_fd_sc_hd__dfxtp_4
X_51947_ _51947_/A _51947_/B _51947_/Y sky130_fd_sc_hd__nand2_4
X_70781_ _70387_/A _70782_/A sky130_fd_sc_hd__buf_2
X_82767_ _82769_/CLK _82767_/D _82767_/Q sky130_fd_sc_hd__dfxtp_4
X_41700_ _41577_/X _82900_/Q _41699_/X _41700_/Y sky130_fd_sc_hd__o21ai_4
X_72520_ _72597_/B _72597_/C _72583_/C _72510_/C _59789_/A _72520_/X
+ sky130_fd_sc_hd__a41o_4
X_84506_ _84501_/CLK _61217_/X _84506_/Q sky130_fd_sc_hd__dfxtp_4
X_57454_ _57441_/X _56758_/X _57453_/X _57454_/X sky130_fd_sc_hd__o21a_4
X_81718_ _81532_/CLK _81718_/D _81718_/Q sky130_fd_sc_hd__dfxtp_4
X_88274_ _88272_/CLK _41122_/X _88274_/Q sky130_fd_sc_hd__dfxtp_4
X_54666_ _54558_/A _54666_/X sky130_fd_sc_hd__buf_2
X_42680_ _42680_/A _42681_/A sky130_fd_sc_hd__buf_2
X_85486_ _86317_/CLK _54200_/Y _85486_/Q sky130_fd_sc_hd__dfxtp_4
X_51878_ _51870_/A _51870_/B _51870_/C _52704_/D _51878_/X sky130_fd_sc_hd__and4_4
X_82698_ _84111_/CLK _82698_/D _82686_/D sky130_fd_sc_hd__dfxtp_4
X_56405_ _56397_/X _56399_/B _85206_/Q _56405_/Y sky130_fd_sc_hd__nand3_4
X_87225_ _87225_/CLK _87225_/D _69011_/B sky130_fd_sc_hd__dfxtp_4
X_41631_ _41630_/X _41631_/X sky130_fd_sc_hd__buf_2
X_53617_ _85601_/Q _53556_/X _53616_/Y _53617_/Y sky130_fd_sc_hd__o21ai_4
X_72451_ _65308_/X _85669_/Q _72422_/X _72451_/X sky130_fd_sc_hd__o21a_4
X_84437_ _84438_/CLK _62053_/Y _78060_/B sky130_fd_sc_hd__dfxtp_4
X_50829_ _50538_/A _50830_/C sky130_fd_sc_hd__buf_2
X_81649_ _81811_/CLK _81681_/Q _76365_/A sky130_fd_sc_hd__dfxtp_4
X_57385_ _57380_/X _57385_/X sky130_fd_sc_hd__buf_2
X_54597_ _85413_/Q _54593_/X _54596_/Y _54597_/Y sky130_fd_sc_hd__o21ai_4
X_59124_ _59037_/A _59124_/X sky130_fd_sc_hd__buf_2
X_71402_ _71397_/X _83512_/Q _71401_/Y _83512_/D sky130_fd_sc_hd__a21o_4
X_44350_ _44381_/A _44350_/X sky130_fd_sc_hd__buf_2
X_56336_ _56103_/X _56321_/X _56335_/Y _56336_/Y sky130_fd_sc_hd__o21ai_4
X_75170_ _80681_/Q _80937_/D _75175_/C sky130_fd_sc_hd__nand2_4
X_87156_ _86934_/CLK _87156_/D _87156_/Q sky130_fd_sc_hd__dfxtp_4
X_41562_ _40586_/A _41563_/B sky130_fd_sc_hd__buf_2
X_53548_ _53548_/A _48022_/Y _53548_/Y sky130_fd_sc_hd__nand2_4
X_72382_ _72347_/A _86283_/Q _72382_/Y sky130_fd_sc_hd__nor2_4
X_84368_ _84449_/CLK _84368_/D _62943_/C sky130_fd_sc_hd__dfxtp_4
X_43301_ _43217_/A _43302_/A sky130_fd_sc_hd__buf_2
X_74121_ _74121_/A _73372_/B _74121_/Y sky130_fd_sc_hd__nor2_4
X_86107_ _85786_/CLK _50920_/Y _86107_/Q sky130_fd_sc_hd__dfxtp_4
X_40513_ _82313_/Q _40471_/X _40513_/X sky130_fd_sc_hd__or2_4
X_59055_ _84773_/Q _59043_/X _59047_/X _59054_/X _84773_/D sky130_fd_sc_hd__a2bb2oi_4
X_71333_ _71335_/A _71335_/B _71333_/C _71333_/Y sky130_fd_sc_hd__nand3_4
X_83319_ _83316_/CLK _83319_/D _55671_/A sky130_fd_sc_hd__dfxtp_4
X_44281_ _44279_/Y _44280_/Y _44277_/X _44281_/Y sky130_fd_sc_hd__a21oi_4
X_56267_ _56194_/X _56263_/B _56267_/C _56267_/Y sky130_fd_sc_hd__nand3_4
X_87087_ _87103_/CLK _44479_/X _87087_/Q sky130_fd_sc_hd__dfxtp_4
X_41493_ _41492_/X _41493_/X sky130_fd_sc_hd__buf_2
X_53479_ _85629_/Q _53476_/X _53478_/Y _53479_/Y sky130_fd_sc_hd__o21ai_4
X_84299_ _84299_/CLK _63711_/Y _80279_/B sky130_fd_sc_hd__dfxtp_4
X_46020_ _46013_/X _46001_/X _40531_/X _86810_/Q _46014_/X _46021_/A
+ sky130_fd_sc_hd__o32ai_4
X_58006_ _86637_/Q _57954_/X _58006_/Y sky130_fd_sc_hd__nor2_4
X_43232_ _43212_/A _43232_/X sky130_fd_sc_hd__buf_2
X_55218_ _72718_/C _83314_/Q _72718_/D _55218_/Y sky130_fd_sc_hd__nand3_4
X_86038_ _85527_/CLK _51295_/Y _86038_/Q sky130_fd_sc_hd__dfxtp_4
X_74052_ _68886_/B _73891_/X _73962_/X _74051_/Y _74052_/X sky130_fd_sc_hd__a211o_4
X_40444_ _40368_/X _41523_/A _40444_/X sky130_fd_sc_hd__or2_4
X_71264_ _71264_/A _71264_/X sky130_fd_sc_hd__buf_2
X_56198_ _56280_/A _56192_/B _56198_/C _56198_/Y sky130_fd_sc_hd__nand3_4
X_73003_ _87306_/Q _73003_/B _73003_/Y sky130_fd_sc_hd__nor2_4
X_70215_ _70209_/X _83834_/Q _70214_/X _83834_/D sky130_fd_sc_hd__a21o_4
X_43163_ _43162_/X _43149_/X _40866_/X _73252_/A _43154_/X _43164_/A
+ sky130_fd_sc_hd__o32ai_4
X_55149_ _55149_/A _55224_/A sky130_fd_sc_hd__buf_2
X_78860_ _78854_/Y _78855_/X _78859_/Y _78860_/Y sky130_fd_sc_hd__a21oi_4
X_40375_ _44736_/A _40375_/X sky130_fd_sc_hd__buf_2
X_71195_ _48540_/B _71190_/X _71194_/Y _83577_/D sky130_fd_sc_hd__o21ai_4
X_42114_ _41064_/X _42103_/X _88028_/Q _42104_/X _88028_/D sky130_fd_sc_hd__a2bb2o_4
X_77811_ _77808_/X _77811_/B _77812_/B sky130_fd_sc_hd__xnor2_4
X_70146_ _83522_/Q _83170_/Q _83503_/Q _83151_/Q _70146_/Y sky130_fd_sc_hd__a22oi_4
X_47971_ _47904_/A _47971_/X sky130_fd_sc_hd__buf_2
X_43094_ _87578_/Q _43094_/Y sky130_fd_sc_hd__inv_2
X_59957_ _59885_/Y _61205_/B sky130_fd_sc_hd__inv_2
X_78791_ _82817_/Q _78791_/B _78792_/B sky130_fd_sc_hd__xor2_4
X_87989_ _87993_/CLK _87989_/D _87989_/Q sky130_fd_sc_hd__dfxtp_4
X_49710_ _49699_/A _52924_/B _49710_/Y sky130_fd_sc_hd__nand2_4
X_46922_ _46948_/A _52748_/B _46922_/Y sky130_fd_sc_hd__nand2_4
X_42045_ _42028_/X _42043_/X _40894_/X _73372_/A _42044_/X _42046_/A
+ sky130_fd_sc_hd__o32ai_4
X_58908_ _84791_/Q _58871_/X _58899_/X _58907_/X _58908_/Y sky130_fd_sc_hd__a2bb2oi_4
X_77742_ _77742_/A _77741_/Y _77742_/Y sky130_fd_sc_hd__nand2_4
X_74954_ _81136_/D _74960_/C _74953_/Y _74954_/Y sky130_fd_sc_hd__a21oi_4
X_70077_ _69003_/X _69005_/X _69992_/X _70079_/A sky130_fd_sc_hd__a21o_4
X_59888_ _59585_/A _60593_/B sky130_fd_sc_hd__buf_2
X_49641_ _49641_/A _49642_/B sky130_fd_sc_hd__buf_2
X_73905_ _73854_/X _85619_/Q _73903_/X _73904_/X _73905_/X sky130_fd_sc_hd__a211o_4
X_58839_ _58813_/X _85772_/Q _58838_/X _58839_/X sky130_fd_sc_hd__o21a_4
X_46853_ _58887_/A _46813_/X _46852_/Y _46853_/Y sky130_fd_sc_hd__o21ai_4
X_77673_ _77674_/A _82123_/Q _77673_/Y sky130_fd_sc_hd__nor2_4
X_74885_ _74899_/A _74887_/B sky130_fd_sc_hd__inv_2
X_79412_ _79404_/X _79405_/X _79411_/Y _79416_/A sky130_fd_sc_hd__a21boi_4
X_45804_ _45799_/X _45802_/Y _45803_/X _45804_/Y sky130_fd_sc_hd__a21oi_4
X_76624_ _76616_/X _76624_/B _76624_/C _76624_/Y sky130_fd_sc_hd__nand3_4
X_49572_ _49571_/X _49561_/B _49548_/X _52785_/D _49572_/X sky130_fd_sc_hd__and4_4
X_61850_ _61848_/Y _61801_/X _61849_/Y _61850_/Y sky130_fd_sc_hd__a21oi_4
X_73836_ _53514_/B _73836_/B _73836_/X sky130_fd_sc_hd__xor2_4
X_46784_ _46784_/A _46784_/B _46784_/C _46783_/X _46784_/X sky130_fd_sc_hd__and4_4
X_43996_ _59571_/C _60665_/C _59563_/A _59584_/C sky130_fd_sc_hd__nand3_4
X_48523_ _50469_/A _48500_/X _48533_/C _48523_/X sky130_fd_sc_hd__and3_4
X_60801_ _60804_/B _60725_/B _60785_/Y _60801_/X sky130_fd_sc_hd__o21a_4
X_79343_ _79343_/A _79343_/B _79344_/B sky130_fd_sc_hd__xor2_4
X_45735_ _45705_/A _45736_/B sky130_fd_sc_hd__buf_2
X_76555_ _76554_/B _76554_/C _76550_/Y _76555_/Y sky130_fd_sc_hd__o21ai_4
X_42947_ _42946_/Y _87637_/D sky130_fd_sc_hd__inv_2
X_61781_ _61780_/X _61765_/B _61765_/C _61748_/X _61781_/Y sky130_fd_sc_hd__nand4_4
X_73767_ _73765_/X _73767_/B _73767_/C _73767_/Y sky130_fd_sc_hd__nand3_4
X_70979_ _70976_/A _71066_/B _70979_/C _70979_/Y sky130_fd_sc_hd__nand3_4
X_63520_ _63496_/A _63520_/B _63520_/C _63496_/D _63520_/X sky130_fd_sc_hd__and4_4
X_75506_ _75466_/A _75466_/B _75506_/C _75506_/D _75506_/X sky130_fd_sc_hd__and4_4
X_60732_ _60711_/X _60660_/X _60732_/C _60732_/Y sky130_fd_sc_hd__nand3_4
X_48454_ _83584_/Q _53663_/B sky130_fd_sc_hd__inv_2
X_72718_ _45893_/C _44907_/A _72718_/C _72718_/D _72718_/X sky130_fd_sc_hd__and4_4
X_79274_ _79272_/Y _79253_/Y _79273_/X _79275_/B sky130_fd_sc_hd__o21ai_4
X_45666_ _82992_/Q _45388_/X _45665_/X _45666_/Y sky130_fd_sc_hd__o21ai_4
X_76486_ _76486_/A _76485_/X _81336_/D sky130_fd_sc_hd__xor2_4
X_42878_ _41601_/X _42866_/X _67223_/B _42867_/X _87672_/D sky130_fd_sc_hd__a2bb2o_4
X_73698_ _73343_/X _73698_/X sky130_fd_sc_hd__buf_2
X_47405_ _86638_/Q _47382_/X _47404_/Y _47405_/Y sky130_fd_sc_hd__o21ai_4
X_78225_ _78225_/A _78234_/A _78226_/B sky130_fd_sc_hd__xor2_4
X_44617_ _46298_/A _44618_/A sky130_fd_sc_hd__buf_2
X_63451_ _63463_/A _84898_/Q _63463_/C _63451_/X sky130_fd_sc_hd__and3_4
X_75437_ _75401_/Y _75435_/D _75435_/B _75437_/X sky130_fd_sc_hd__a21bo_4
X_41829_ _41829_/A _41829_/Y sky130_fd_sc_hd__inv_2
X_48385_ _48384_/Y _48449_/B _48385_/Y sky130_fd_sc_hd__nand2_4
X_60663_ _60720_/A _60687_/A _60632_/A _60702_/C _60663_/Y sky130_fd_sc_hd__nand4_4
X_72649_ _70188_/C _72645_/X _72648_/Y _72649_/X sky130_fd_sc_hd__a21bo_4
X_45597_ _45597_/A _45597_/B _45597_/Y sky130_fd_sc_hd__nor2_4
X_62402_ _62203_/Y _62448_/A sky130_fd_sc_hd__buf_2
X_47336_ _47333_/X _52991_/B _47336_/Y sky130_fd_sc_hd__nand2_4
X_66170_ _66167_/X _66169_/X _65961_/X _66173_/A sky130_fd_sc_hd__a21o_4
X_78156_ _78154_/X _78162_/C _78156_/Y sky130_fd_sc_hd__nand2_4
X_44548_ _44548_/A _44548_/X sky130_fd_sc_hd__buf_2
X_63382_ _63305_/X _63392_/B _80614_/B _63382_/Y sky130_fd_sc_hd__nor3_4
X_75368_ _75347_/X _75366_/Y _75367_/Y _75368_/X sky130_fd_sc_hd__a21bo_4
X_60594_ _60594_/A _60596_/A sky130_fd_sc_hd__inv_2
X_65121_ _65118_/X _85517_/Q _64919_/X _65120_/X _65121_/X sky130_fd_sc_hd__a211o_4
X_77107_ _77114_/B _82288_/D _77107_/Y sky130_fd_sc_hd__nand2_4
X_62333_ _62319_/A _63459_/B _62319_/C _62335_/C sky130_fd_sc_hd__nand3_4
X_74319_ _74325_/A _74325_/B _56073_/A _74319_/Y sky130_fd_sc_hd__nand3_4
X_47267_ _83388_/Q _54121_/B sky130_fd_sc_hd__inv_2
X_78087_ _78088_/A _78088_/B _78087_/Y sky130_fd_sc_hd__nor2_4
X_44479_ _41198_/Y _44474_/X _87087_/Q _44475_/X _44479_/X sky130_fd_sc_hd__a2bb2o_4
X_75299_ _75299_/A _75299_/Y sky130_fd_sc_hd__inv_2
X_49006_ _53841_/B _49006_/X sky130_fd_sc_hd__buf_2
X_46218_ _44031_/X _46098_/A _46214_/C _46214_/D _46218_/Y sky130_fd_sc_hd__nand4_4
X_65052_ _64696_/X _85520_/Q _64697_/X _65051_/X _65052_/X sky130_fd_sc_hd__a211o_4
X_77038_ _81992_/Q _82280_/D _77038_/X sky130_fd_sc_hd__xor2_4
X_62264_ _62256_/X _62258_/X _62263_/Y _84918_/Q _62214_/X _62264_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47198_ _46725_/A _47198_/X sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_16 _44273_/Y _44274_/D sky130_fd_sc_hd__buf_8
X_64003_ _61522_/X _64052_/B _64003_/C _64052_/D _64003_/Y sky130_fd_sc_hd__nand4_4
X_61215_ _61112_/X _61096_/X _61103_/X _61205_/A _60528_/A _61215_/Y
+ sky130_fd_sc_hd__a41oi_4
Xpsn_inst_psn_buff_27 _50212_/A _41909_/B1 sky130_fd_sc_hd__buf_2
X_46149_ _46120_/A _46120_/B _49380_/C _46149_/Y sky130_fd_sc_hd__nand3_4
X_69860_ _68934_/X _69860_/B _69860_/Y sky130_fd_sc_hd__nor2_4
X_62195_ _62195_/A _62195_/Y sky130_fd_sc_hd__inv_2
X_68811_ _68798_/Y _68358_/X _68649_/X _68810_/Y _68811_/X sky130_fd_sc_hd__a211o_4
X_61146_ _61145_/X _64523_/D sky130_fd_sc_hd__buf_2
X_69791_ _69791_/A _69790_/Y _69791_/Y sky130_fd_sc_hd__nor2_4
X_78989_ _78967_/Y _82516_/D sky130_fd_sc_hd__inv_2
X_49908_ _49928_/A _53122_/B _49908_/Y sky130_fd_sc_hd__nand2_4
X_68742_ _68742_/A _69067_/A sky130_fd_sc_hd__buf_2
X_65954_ _65903_/X _65477_/Y _65953_/Y _65954_/Y sky130_fd_sc_hd__o21ai_4
X_61077_ _61144_/A _61083_/C sky130_fd_sc_hd__inv_2
X_64905_ _64752_/X _86166_/Q _64902_/X _64904_/X _64905_/X sky130_fd_sc_hd__a211o_4
X_60028_ _62194_/D _60091_/C _60027_/X _60028_/Y sky130_fd_sc_hd__nand3_4
X_49839_ _49830_/A _49851_/B _49830_/C _53052_/D _49839_/X sky130_fd_sc_hd__and4_4
X_80951_ _81996_/CLK _75376_/B _80951_/Q sky130_fd_sc_hd__dfxtp_4
X_68673_ _73845_/A _68493_/X _68494_/X _68672_/Y _68673_/X sky130_fd_sc_hd__a211o_4
X_65885_ _65390_/X _65828_/B _65393_/X _65885_/Y sky130_fd_sc_hd__nand3_4
X_67624_ _67863_/A _67624_/X sky130_fd_sc_hd__buf_2
X_52850_ _52850_/A _52850_/B _52850_/Y sky130_fd_sc_hd__nand2_4
X_64836_ _64836_/A _86457_/Q _64836_/X sky130_fd_sc_hd__and2_4
X_83670_ _83673_/CLK _70898_/Y _46794_/A sky130_fd_sc_hd__dfxtp_4
X_80882_ _81130_/CLK _75724_/B _80882_/Q sky130_fd_sc_hd__dfxtp_4
X_51801_ _85943_/Q _51789_/X _51800_/Y _51801_/Y sky130_fd_sc_hd__o21ai_4
X_82621_ _82589_/CLK _82621_/D _82621_/Q sky130_fd_sc_hd__dfxtp_4
X_67555_ _67555_/A _67555_/B _67555_/Y sky130_fd_sc_hd__nand2_4
X_52781_ _52773_/A _52781_/B _52781_/Y sky130_fd_sc_hd__nand2_4
X_64767_ _64767_/A _85851_/Q _64767_/X sky130_fd_sc_hd__and2_4
X_61979_ _61962_/X _61945_/X _63557_/B _61947_/D _61979_/X sky130_fd_sc_hd__and4_4
X_54520_ _54245_/A _54521_/A sky130_fd_sc_hd__buf_2
X_66506_ _66504_/Y _66483_/X _66505_/X _84110_/D sky130_fd_sc_hd__a21o_4
X_85340_ _85372_/CLK _54988_/Y _85340_/Q sky130_fd_sc_hd__dfxtp_4
X_51732_ _51737_/A _53255_/B _51732_/Y sky130_fd_sc_hd__nand2_4
X_63718_ _63701_/A _63701_/B _80268_/B _63718_/Y sky130_fd_sc_hd__nor3_4
X_82552_ _83133_/CLK _82552_/D _82552_/Q sky130_fd_sc_hd__dfxtp_4
X_67486_ _87981_/Q _67414_/X _67391_/X _67485_/X _67486_/X sky130_fd_sc_hd__a211o_4
X_64698_ _64616_/A _65836_/A sky130_fd_sc_hd__buf_2
X_81503_ _81461_/CLK _84071_/Q _81503_/Q sky130_fd_sc_hd__dfxtp_4
X_69225_ _87033_/Q _69182_/X _69183_/X _69224_/X _69226_/B sky130_fd_sc_hd__a211o_4
X_54451_ _54446_/A _54451_/B _54451_/Y sky130_fd_sc_hd__nand2_4
X_66437_ _64978_/X _66518_/B _64982_/X _66437_/Y sky130_fd_sc_hd__nand3_4
X_85271_ _85270_/CLK _85271_/D _56219_/C sky130_fd_sc_hd__dfxtp_4
X_51663_ _51657_/X _51651_/B _51684_/C _53185_/D _51663_/X sky130_fd_sc_hd__and4_4
X_63649_ _58184_/A _60798_/X _63384_/C _60703_/Y _62097_/X _63649_/X
+ sky130_fd_sc_hd__a32o_4
X_82483_ _82532_/CLK _78564_/X _82483_/Q sky130_fd_sc_hd__dfxtp_4
X_87010_ _88283_/CLK _44664_/X _87010_/Q sky130_fd_sc_hd__dfxtp_4
X_53402_ _53397_/A _53402_/B _53388_/C _52887_/D _53402_/X sky130_fd_sc_hd__and4_4
X_84222_ _85315_/CLK _84222_/D _84222_/Q sky130_fd_sc_hd__dfxtp_4
X_50614_ _50572_/A _50624_/A sky130_fd_sc_hd__buf_2
X_57170_ _57170_/A _57170_/B _56800_/X _57156_/X _57170_/Y sky130_fd_sc_hd__nand4_4
X_81434_ _82648_/CLK _81466_/Q _76092_/B sky130_fd_sc_hd__dfxtp_4
X_69156_ _69156_/A _69156_/X sky130_fd_sc_hd__buf_2
X_54382_ _54378_/A _52692_/B _54382_/Y sky130_fd_sc_hd__nand2_4
X_66368_ _66366_/X _64623_/Y _66367_/Y _66368_/Y sky130_fd_sc_hd__o21ai_4
X_51594_ _51621_/A _51594_/X sky130_fd_sc_hd__buf_2
X_68107_ _66681_/X _66684_/X _68106_/X _68107_/Y sky130_fd_sc_hd__a21oi_4
X_56121_ _56121_/A _56121_/X sky130_fd_sc_hd__buf_2
X_53333_ _85653_/Q _53324_/X _53332_/Y _53333_/Y sky130_fd_sc_hd__o21ai_4
X_65319_ _65319_/A _65319_/B _65319_/X sky130_fd_sc_hd__and2_4
X_84153_ _82746_/CLK _66152_/X _84153_/Q sky130_fd_sc_hd__dfxtp_4
X_50545_ _50541_/A _48684_/B _50545_/Y sky130_fd_sc_hd__nand2_4
X_81365_ _81461_/CLK _76832_/Y _81365_/Q sky130_fd_sc_hd__dfxtp_4
X_69087_ _87573_/Q _68636_/X _68517_/X _69086_/X _69087_/X sky130_fd_sc_hd__a211o_4
X_66299_ _66236_/X _85606_/Q _66251_/X _66298_/X _66299_/X sky130_fd_sc_hd__a211o_4
X_83104_ _83846_/CLK _74309_/X _70292_/C sky130_fd_sc_hd__dfxtp_4
X_56052_ _56052_/A _56052_/B _55913_/B _56052_/Y sky130_fd_sc_hd__nand3_4
X_80316_ _80313_/Y _80314_/Y _80315_/A _80318_/A sky130_fd_sc_hd__a21o_4
X_68038_ _67782_/X _68027_/Y _67983_/X _68037_/Y _68038_/X sky130_fd_sc_hd__a211o_4
X_53264_ _85665_/Q _51900_/X _53263_/Y _53264_/Y sky130_fd_sc_hd__o21ai_4
X_84084_ _83918_/CLK _84084_/D _84084_/Q sky130_fd_sc_hd__dfxtp_4
X_50476_ _50472_/Y _50474_/X _50475_/Y _50476_/Y sky130_fd_sc_hd__a21boi_4
X_81296_ _81296_/CLK _76984_/X _81264_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_442_0_CLK clkbuf_9_221_0_CLK/X _84197_/CLK sky130_fd_sc_hd__clkbuf_1
X_55003_ _85337_/Q _54994_/X _55002_/Y _55003_/Y sky130_fd_sc_hd__o21ai_4
X_52215_ _52215_/A _52220_/A sky130_fd_sc_hd__buf_2
X_83035_ _85213_/CLK _83035_/D _83035_/Q sky130_fd_sc_hd__dfxtp_4
X_87912_ _86932_/CLK _42341_/X _87912_/Q sky130_fd_sc_hd__dfxtp_4
X_80247_ _80244_/Y _80227_/Y _80246_/X _80247_/Y sky130_fd_sc_hd__o21ai_4
X_53195_ _53195_/A _53195_/X sky130_fd_sc_hd__buf_2
X_70000_ _82556_/D _69988_/X _69999_/X _83876_/D sky130_fd_sc_hd__a21bo_4
X_59811_ _59810_/Y _59811_/Y sky130_fd_sc_hd__inv_2
X_52146_ _50443_/A _52140_/X _52156_/C _52146_/X sky130_fd_sc_hd__and3_4
X_87843_ _88104_/CLK _87843_/D _73940_/A sky130_fd_sc_hd__dfxtp_4
X_80178_ _80178_/A _80178_/B _80178_/Y sky130_fd_sc_hd__nand2_4
X_69989_ _69610_/X _69613_/X _69939_/X _69989_/Y sky130_fd_sc_hd__a21oi_4
X_59742_ _59742_/A _59742_/Y sky130_fd_sc_hd__inv_2
X_52077_ _52121_/A _48335_/B _52077_/Y sky130_fd_sc_hd__nand2_4
X_56954_ _56602_/X _85115_/Q _56953_/X _56954_/Y sky130_fd_sc_hd__nor3_4
X_87774_ _87525_/CLK _42678_/Y _87774_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_457_0_CLK clkbuf_9_228_0_CLK/X _86297_/CLK sky130_fd_sc_hd__clkbuf_1
X_84986_ _86558_/CLK _84986_/D _84986_/Q sky130_fd_sc_hd__dfxtp_4
X_55905_ _55903_/A _56488_/C _55905_/X sky130_fd_sc_hd__and2_4
X_51028_ _50973_/A _51029_/A sky130_fd_sc_hd__buf_2
X_86725_ _86119_/CLK _86725_/D _86725_/Q sky130_fd_sc_hd__dfxtp_4
X_71951_ _71570_/X _70538_/X _71598_/C _71951_/Y sky130_fd_sc_hd__nor3_4
X_83937_ _84087_/CLK _69258_/X _83937_/Q sky130_fd_sc_hd__dfxtp_4
X_59673_ _59770_/A _60036_/A sky130_fd_sc_hd__buf_2
X_56885_ _56885_/A _56884_/Y _56886_/B sky130_fd_sc_hd__and2_4
X_70902_ _50998_/B _70885_/A _70901_/Y _70902_/Y sky130_fd_sc_hd__o21ai_4
X_58624_ _58857_/A _58624_/X sky130_fd_sc_hd__buf_2
X_43850_ _41199_/X _43842_/X _87235_/Q _43843_/X _43850_/X sky130_fd_sc_hd__a2bb2o_4
X_55836_ _55836_/A _55836_/B _55836_/X sky130_fd_sc_hd__and2_4
X_74670_ _74679_/A _45697_/A _74670_/Y sky130_fd_sc_hd__nand2_4
X_86656_ _85727_/CLK _47238_/Y _57722_/A sky130_fd_sc_hd__dfxtp_4
X_71882_ _71871_/X _83342_/Q _71881_/Y _71882_/X sky130_fd_sc_hd__a21o_4
X_83868_ _82541_/CLK _70032_/X _83868_/Q sky130_fd_sc_hd__dfxtp_4
X_42801_ _41393_/X _42787_/X _67808_/B _42788_/X _42801_/X sky130_fd_sc_hd__a2bb2o_4
X_73621_ _73619_/X _73601_/X _73604_/Y _73621_/Y sky130_fd_sc_hd__nand3_4
X_85607_ _86535_/CLK _85607_/D _85607_/Q sky130_fd_sc_hd__dfxtp_4
X_70833_ _70860_/A _70791_/B _71066_/C _70841_/D _70833_/Y sky130_fd_sc_hd__nand4_4
X_58555_ _58538_/X _83356_/Q _58554_/Y _58555_/X sky130_fd_sc_hd__o21a_4
X_82819_ _82786_/CLK _79523_/X _82787_/D sky130_fd_sc_hd__dfxtp_4
X_43781_ _43760_/A _43781_/X sky130_fd_sc_hd__buf_2
X_55767_ _85193_/Q _55152_/X _55168_/A _55766_/X _55767_/X sky130_fd_sc_hd__a211o_4
X_86587_ _86587_/CLK _86587_/D _73711_/B sky130_fd_sc_hd__dfxtp_4
X_40993_ _40991_/X _81718_/Q _40992_/X _40994_/A sky130_fd_sc_hd__o21a_4
X_52979_ _52979_/A _52979_/B _52979_/Y sky130_fd_sc_hd__nand2_4
X_83799_ _83842_/CLK _70319_/Y _70317_/A sky130_fd_sc_hd__dfxtp_4
X_45520_ _45395_/X _45520_/X sky130_fd_sc_hd__buf_2
X_57506_ _71978_/A _57506_/X sky130_fd_sc_hd__buf_2
X_76340_ _76302_/Y _76306_/A _76317_/B _76340_/X sky130_fd_sc_hd__a21o_4
X_88326_ _88326_/CLK _88326_/D _69740_/B sky130_fd_sc_hd__dfxtp_4
X_42732_ _42700_/A _42732_/X sky130_fd_sc_hd__buf_2
X_54718_ _54718_/A _47403_/A _54718_/Y sky130_fd_sc_hd__nand2_4
X_85538_ _85538_/CLK _85538_/D _85538_/Q sky130_fd_sc_hd__dfxtp_4
X_73552_ _73552_/A _73438_/B _73552_/Y sky130_fd_sc_hd__nor2_4
X_70764_ _70764_/A _70772_/A sky130_fd_sc_hd__buf_2
X_58486_ _84837_/Q _58487_/A sky130_fd_sc_hd__buf_2
X_55698_ _55698_/A _55990_/C _55698_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_501_0_CLK clkbuf_9_501_0_CLK/A clkbuf_9_501_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_72503_ _72503_/A _61302_/A _72516_/B sky130_fd_sc_hd__nor2_4
X_45451_ _63041_/B _61367_/A sky130_fd_sc_hd__buf_2
X_57437_ _56797_/A _57445_/B _56796_/Y _57437_/Y sky130_fd_sc_hd__nand3_4
X_76271_ _76241_/X _76269_/Y _76270_/X _76271_/X sky130_fd_sc_hd__o21a_4
X_88257_ _87083_/CLK _88257_/D _68820_/B sky130_fd_sc_hd__dfxtp_4
X_42663_ _42647_/X _42648_/X _41016_/X _87781_/Q _42658_/X _42663_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54649_ _54594_/X _54649_/X sky130_fd_sc_hd__buf_2
X_73483_ _83149_/Q _73437_/X _73482_/Y _73483_/X sky130_fd_sc_hd__a21o_4
X_85469_ _82206_/CLK _54293_/Y _85469_/Q sky130_fd_sc_hd__dfxtp_4
X_70695_ _70695_/A _70698_/A sky130_fd_sc_hd__buf_2
X_78010_ _78010_/A _77998_/A _78011_/A sky130_fd_sc_hd__and2_4
X_44402_ _41507_/X _44394_/X _87126_/Q _44395_/X _44402_/X sky130_fd_sc_hd__a2bb2o_4
X_75222_ _80684_/Q _80984_/Q _75222_/Y sky130_fd_sc_hd__nand2_4
X_87208_ _87720_/CLK _87208_/D _67596_/B sky130_fd_sc_hd__dfxtp_4
X_41614_ _40536_/B _41563_/B _41614_/X sky130_fd_sc_hd__or2_4
X_48170_ _48169_/X _48170_/X sky130_fd_sc_hd__buf_2
X_72434_ _72431_/Y _72433_/Y _57779_/X _72434_/X sky130_fd_sc_hd__a21o_4
X_45382_ _45379_/X _45381_/Y _45348_/X _45382_/Y sky130_fd_sc_hd__a21oi_4
X_57368_ _57368_/A _85027_/D sky130_fd_sc_hd__inv_2
X_88188_ _87110_/CLK _88188_/D _67128_/B sky130_fd_sc_hd__dfxtp_4
X_42594_ _42593_/Y _87809_/D sky130_fd_sc_hd__inv_2
X_47121_ _47113_/A _47082_/X _47091_/X _52867_/D _47121_/X sky130_fd_sc_hd__and4_4
X_59107_ _59105_/X _85752_/Q _59106_/X _59107_/X sky130_fd_sc_hd__o21a_4
X_44333_ _44330_/X _44331_/X _41656_/X _87162_/Q _44332_/X _44333_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56319_ _56309_/A _56312_/X _55874_/B _56319_/Y sky130_fd_sc_hd__nand3_4
X_87139_ _88215_/CLK _87139_/D _87139_/Q sky130_fd_sc_hd__dfxtp_4
X_75153_ _75153_/A _75153_/Y sky130_fd_sc_hd__inv_2
X_41545_ _41544_/X _41545_/X sky130_fd_sc_hd__buf_2
X_72365_ _72360_/Y _72364_/Y _72292_/X _72365_/X sky130_fd_sc_hd__a21o_4
X_57299_ _57427_/A _57340_/C _56750_/Y _57299_/Y sky130_fd_sc_hd__nand3_4
X_74104_ _73583_/A _74104_/B _74104_/X sky130_fd_sc_hd__and2_4
X_47052_ _47052_/A _47053_/A sky130_fd_sc_hd__inv_2
X_59038_ _59013_/X _85758_/Q _59037_/X _59038_/X sky130_fd_sc_hd__o21a_4
X_71316_ _71500_/A _71314_/B _71779_/B _71316_/Y sky130_fd_sc_hd__nand3_4
X_44264_ _44263_/X _57837_/A sky130_fd_sc_hd__buf_2
X_79961_ _79961_/A _79960_/Y _79964_/A sky130_fd_sc_hd__nand2_4
X_75084_ _75082_/X _75102_/B _75085_/B _75091_/A sky130_fd_sc_hd__a21o_4
X_41476_ _41476_/A _88208_/D sky130_fd_sc_hd__inv_2
X_72296_ _72296_/A _72296_/X sky130_fd_sc_hd__buf_2
X_46003_ _46002_/Y _86820_/D sky130_fd_sc_hd__inv_2
X_43215_ _40964_/X _43180_/X _87534_/Q _43185_/X _87534_/D sky130_fd_sc_hd__a2bb2o_4
X_74035_ _74032_/X _74034_/X _73944_/X _74048_/B sky130_fd_sc_hd__a21o_4
X_78912_ _78912_/A _78912_/B _78919_/A sky130_fd_sc_hd__xor2_4
X_40427_ _57491_/A _40364_/X _40426_/X _88393_/Q _40375_/X _40428_/A
+ sky130_fd_sc_hd__o32ai_4
X_71247_ _50224_/B _71239_/X _71246_/Y _71247_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_7_1_0_CLK clkbuf_6_0_0_CLK/X clkbuf_8_3_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_44195_ _72739_/A _44194_/X _44195_/Y sky130_fd_sc_hd__nor2_4
X_79892_ _79890_/Y _79891_/Y _79892_/Y sky130_fd_sc_hd__nand2_4
X_61000_ _60422_/A _61000_/X sky130_fd_sc_hd__buf_2
X_43146_ _43146_/A _43146_/X sky130_fd_sc_hd__buf_2
X_78843_ _78837_/B _78841_/Y _78842_/Y _78854_/B sky130_fd_sc_hd__a21oi_4
X_40358_ _40435_/A _44587_/A sky130_fd_sc_hd__buf_2
X_71178_ _71178_/A _71185_/B _71181_/C _71178_/D _71178_/Y sky130_fd_sc_hd__nand4_4
X_70129_ _70129_/A _70129_/B _70131_/B sky130_fd_sc_hd__nor2_4
X_47954_ _47846_/A _47954_/X sky130_fd_sc_hd__buf_2
X_43077_ _43076_/Y _87585_/D sky130_fd_sc_hd__inv_2
X_78774_ _78749_/Y _78753_/B _78752_/A _78778_/A sky130_fd_sc_hd__o21a_4
X_75986_ _75986_/A _75986_/B _81739_/D sky130_fd_sc_hd__xnor2_4
Xclkbuf_8_84_0_CLK clkbuf_8_85_0_CLK/A clkbuf_8_84_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_46905_ _54435_/D _52742_/D sky130_fd_sc_hd__buf_2
X_42028_ _42013_/A _42028_/X sky130_fd_sc_hd__buf_2
X_77725_ _82050_/Q _77725_/Y sky130_fd_sc_hd__inv_2
X_62951_ _62791_/X _62988_/A sky130_fd_sc_hd__buf_2
X_74937_ _81134_/D _74928_/B _74937_/Y sky130_fd_sc_hd__nand2_4
X_47885_ _40877_/X _82365_/Q _47884_/X _47886_/A sky130_fd_sc_hd__o21ai_4
X_49624_ _49571_/A _49625_/A sky130_fd_sc_hd__buf_2
X_61902_ _59668_/B _61902_/X sky130_fd_sc_hd__buf_2
X_46836_ _82954_/Q _54395_/D sky130_fd_sc_hd__inv_2
X_65670_ _65704_/A _86481_/Q _65670_/X sky130_fd_sc_hd__and2_4
X_77656_ _77652_/Y _77654_/Y _77655_/A _77656_/Y sky130_fd_sc_hd__o21ai_4
X_62882_ _62894_/A _62852_/X _84374_/Q _62882_/Y sky130_fd_sc_hd__nor3_4
X_74868_ _80933_/Q _74868_/B _74868_/X sky130_fd_sc_hd__xor2_4
X_64621_ _64621_/A _86432_/Q _64621_/X sky130_fd_sc_hd__and2_4
X_76607_ _76605_/X _76608_/A sky130_fd_sc_hd__inv_2
X_61833_ _61863_/A _61829_/Y _61830_/Y _61832_/Y _61833_/Y sky130_fd_sc_hd__nand4_4
X_49555_ _86366_/Q _49551_/X _49554_/Y _49555_/Y sky130_fd_sc_hd__o21ai_4
X_73819_ _73343_/X _73819_/X sky130_fd_sc_hd__buf_2
X_46767_ _46767_/A _46767_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_99_0_CLK clkbuf_8_99_0_CLK/A clkbuf_8_99_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_77587_ _77586_/X _77587_/Y sky130_fd_sc_hd__inv_2
X_43979_ _43979_/A _43978_/Y _43979_/Y sky130_fd_sc_hd__nor2_4
X_74799_ _74716_/A _70637_/A _74799_/C _74739_/B _74799_/X sky130_fd_sc_hd__and4_4
X_48506_ _86516_/Q _48478_/X _48505_/Y _48506_/Y sky130_fd_sc_hd__o21ai_4
X_67340_ _67340_/A _67339_/X _67340_/Y sky130_fd_sc_hd__nand2_4
X_79326_ _79334_/A _79325_/Y _82831_/D sky130_fd_sc_hd__xnor2_4
X_45718_ _45708_/X _45715_/Y _45717_/Y _45718_/Y sky130_fd_sc_hd__a21oi_4
X_64552_ _63713_/A _61226_/X _64552_/Y sky130_fd_sc_hd__nor2_4
X_76538_ _76537_/X _76540_/B sky130_fd_sc_hd__inv_2
X_49486_ _86378_/Q _49470_/X _49485_/Y _49486_/Y sky130_fd_sc_hd__o21ai_4
X_61764_ _61856_/A _61765_/B sky130_fd_sc_hd__buf_2
X_46698_ _46717_/A _46682_/B _46682_/C _52622_/D _46698_/X sky130_fd_sc_hd__and4_4
X_63503_ _61460_/B _63487_/X _63500_/X _63502_/X _63503_/X sky130_fd_sc_hd__a211o_4
X_48437_ _46317_/A _48642_/A sky130_fd_sc_hd__buf_2
X_60715_ _60036_/A _60715_/X sky130_fd_sc_hd__buf_2
X_67271_ _67270_/X _67271_/X sky130_fd_sc_hd__buf_2
X_79257_ _79256_/Y _79257_/Y sky130_fd_sc_hd__inv_2
X_45649_ _45647_/Y _45632_/X _45616_/X _45648_/Y _45649_/X sky130_fd_sc_hd__a211o_4
X_64483_ _61140_/X _64523_/B _58184_/A _61153_/C _64483_/X sky130_fd_sc_hd__and4_4
X_76469_ _81367_/Q _76469_/B _76469_/X sky130_fd_sc_hd__xor2_4
X_61695_ _61695_/A _61653_/X _61654_/X _61368_/D _61695_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_8_22_0_CLK clkbuf_8_23_0_CLK/A clkbuf_8_22_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_69010_ _69371_/A _69010_/X sky130_fd_sc_hd__buf_2
X_66222_ _66054_/X _74083_/B _66222_/X sky130_fd_sc_hd__and2_4
X_78208_ _78199_/Y _78206_/Y _78207_/Y _78208_/X sky130_fd_sc_hd__o21a_4
X_63434_ _63368_/A _63434_/X sky130_fd_sc_hd__buf_2
X_48368_ _48367_/Y _48368_/X sky130_fd_sc_hd__buf_2
X_60646_ _60662_/A _60687_/A _60646_/Y sky130_fd_sc_hd__nor2_4
X_79188_ _79188_/A _79188_/B _79189_/B sky130_fd_sc_hd__nand2_4
X_47319_ _81815_/Q _47320_/A sky130_fd_sc_hd__inv_2
X_66153_ _64593_/A _66153_/B _66153_/X sky130_fd_sc_hd__and2_4
X_78139_ _82666_/Q _78139_/B _78139_/X sky130_fd_sc_hd__xor2_4
X_63365_ _63305_/X _63392_/B _63365_/C _63365_/Y sky130_fd_sc_hd__nor3_4
X_48299_ _48296_/Y _48273_/X _48298_/Y _86540_/D sky130_fd_sc_hd__a21boi_4
X_60577_ _72250_/A _60577_/X sky130_fd_sc_hd__buf_2
X_65104_ _64999_/X _86126_/Q _64927_/X _65103_/X _65104_/X sky130_fd_sc_hd__a211o_4
X_50330_ _53511_/A _50331_/B sky130_fd_sc_hd__buf_2
X_62316_ _62471_/A _62332_/D sky130_fd_sc_hd__buf_2
X_81150_ _82284_/CLK _81150_/D _40588_/A sky130_fd_sc_hd__dfxtp_4
X_66084_ _44263_/X _66084_/B _66084_/X sky130_fd_sc_hd__and2_4
Xclkbuf_8_37_0_CLK clkbuf_8_37_0_CLK/A clkbuf_8_37_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_63296_ _63293_/Y _63295_/X _63231_/X _63296_/Y sky130_fd_sc_hd__a21oi_4
X_80101_ _84939_/Q _84187_/Q _80101_/X sky130_fd_sc_hd__xor2_4
X_69912_ _44583_/A _66608_/X _58827_/A _69911_/X _69912_/X sky130_fd_sc_hd__a211o_4
X_65035_ _65859_/A _65035_/X sky130_fd_sc_hd__buf_2
X_50261_ _86236_/Q _50250_/X _50260_/Y _50261_/Y sky130_fd_sc_hd__o21ai_4
X_62247_ _62623_/A _62247_/X sky130_fd_sc_hd__buf_2
X_81081_ _80696_/CLK _81113_/Q _75409_/A sky130_fd_sc_hd__dfxtp_4
X_52000_ _51998_/Y _51981_/X _51999_/Y _85909_/D sky130_fd_sc_hd__a21boi_4
X_80032_ _80016_/Y _80019_/Y _80032_/X sky130_fd_sc_hd__or2_4
X_69843_ _87051_/Q _69796_/X _69797_/X _69842_/X _69843_/X sky130_fd_sc_hd__a211o_4
X_50192_ _50105_/A _51242_/A sky130_fd_sc_hd__buf_2
X_62178_ _62120_/A _62181_/A sky130_fd_sc_hd__buf_2
X_61129_ _64303_/A _64523_/B sky130_fd_sc_hd__buf_2
X_84840_ _84840_/CLK _84840_/D _64412_/C sky130_fd_sc_hd__dfxtp_4
X_69774_ _69746_/X _69772_/Y _69733_/X _69773_/Y _69774_/X sky130_fd_sc_hd__a211o_4
X_66986_ _87426_/Q _66915_/X _66984_/X _66985_/X _66986_/X sky130_fd_sc_hd__a211o_4
X_68725_ _68720_/X _68724_/X _68725_/Y sky130_fd_sc_hd__nand2_4
X_53951_ _53951_/A _53951_/B _53951_/Y sky130_fd_sc_hd__nand2_4
X_65937_ _64729_/A _65937_/X sky130_fd_sc_hd__buf_2
X_84771_ _86686_/CLK _84771_/D _84771_/Q sky130_fd_sc_hd__dfxtp_4
X_81983_ _81933_/CLK _81983_/D _81983_/Q sky130_fd_sc_hd__dfxtp_4
X_86510_ _86499_/CLK _48580_/Y _86510_/Q sky130_fd_sc_hd__dfxtp_4
X_52902_ _52821_/A _52902_/X sky130_fd_sc_hd__buf_2
X_83722_ _85378_/CLK _70693_/X _47515_/A sky130_fd_sc_hd__dfxtp_4
X_56670_ _56670_/A _56852_/A sky130_fd_sc_hd__buf_2
X_68656_ _68653_/X _68655_/X _68558_/X _68656_/X sky130_fd_sc_hd__a21o_4
X_80934_ _81059_/CLK _75124_/B _74874_/A sky130_fd_sc_hd__dfxtp_4
X_87490_ _87235_/CLK _87490_/D _87490_/Q sky130_fd_sc_hd__dfxtp_4
X_53882_ _85549_/Q _53869_/X _53881_/Y _53882_/Y sky130_fd_sc_hd__o21ai_4
X_65868_ _65863_/X _65868_/B _65867_/X _65868_/Y sky130_fd_sc_hd__nand3_4
X_55621_ _55947_/A _55691_/A sky130_fd_sc_hd__buf_2
X_67607_ _67604_/X _67606_/X _67561_/X _67607_/X sky130_fd_sc_hd__a21o_4
X_86441_ _86154_/CLK _49133_/Y _86441_/Q sky130_fd_sc_hd__dfxtp_4
X_52833_ _52843_/A _52833_/B _52833_/Y sky130_fd_sc_hd__nand2_4
X_64819_ _64817_/X _86137_/Q _64776_/X _64818_/X _64819_/X sky130_fd_sc_hd__a211o_4
X_83653_ _85822_/CLK _83653_/D _46294_/A sky130_fd_sc_hd__dfxtp_4
X_80865_ _81990_/CLK _80897_/Q _80865_/Q sky130_fd_sc_hd__dfxtp_4
X_68587_ _64665_/A _68587_/X sky130_fd_sc_hd__buf_2
X_65799_ _65796_/X _65725_/B _65798_/X _65799_/Y sky130_fd_sc_hd__nand3_4
X_58340_ _58328_/X _83450_/Q _58339_/Y _84874_/D sky130_fd_sc_hd__o21a_4
X_82604_ _82604_/CLK _78901_/B _82572_/D sky130_fd_sc_hd__dfxtp_4
X_55552_ _55552_/A _55552_/X sky130_fd_sc_hd__buf_2
X_67538_ _67535_/X _67537_/X _67442_/X _67538_/X sky130_fd_sc_hd__a21o_4
X_86372_ _86372_/CLK _86372_/D _86372_/Q sky130_fd_sc_hd__dfxtp_4
X_52764_ _52761_/Y _52755_/X _52763_/X _52764_/Y sky130_fd_sc_hd__a21oi_4
X_83584_ _83584_/CLK _83584_/D _83584_/Q sky130_fd_sc_hd__dfxtp_4
X_80796_ _83957_/CLK _80796_/D _75472_/A sky130_fd_sc_hd__dfxtp_4
X_88111_ _88111_/CLK _41896_/Y _73650_/A sky130_fd_sc_hd__dfxtp_4
X_54503_ _54483_/A _54503_/B _54483_/C _54503_/D _54503_/X sky130_fd_sc_hd__and4_4
X_85323_ _85354_/CLK _85323_/D _85323_/Q sky130_fd_sc_hd__dfxtp_4
X_51715_ _51709_/X _51715_/B _51715_/C _53238_/D _51715_/X sky130_fd_sc_hd__and4_4
X_58271_ _58328_/A _58271_/X sky130_fd_sc_hd__buf_2
X_82535_ _82541_/CLK _82535_/D _82535_/Q sky130_fd_sc_hd__dfxtp_4
X_55483_ _55483_/A _55483_/Y sky130_fd_sc_hd__inv_2
X_67469_ _87162_/Q _67467_/X _67398_/X _67468_/X _67469_/X sky130_fd_sc_hd__a211o_4
X_52695_ _52693_/Y _52673_/X _52694_/X _52695_/Y sky130_fd_sc_hd__a21oi_4
X_57222_ _55657_/Y _57222_/Y sky130_fd_sc_hd__inv_2
X_69208_ _69204_/X _69207_/X _69116_/X _69208_/X sky130_fd_sc_hd__a21o_4
X_88042_ _87789_/CLK _42086_/X _88042_/Q sky130_fd_sc_hd__dfxtp_4
X_54434_ _85443_/Q _54431_/X _54433_/Y _54434_/Y sky130_fd_sc_hd__o21ai_4
X_85254_ _85190_/CLK _85254_/D _85254_/Q sky130_fd_sc_hd__dfxtp_4
X_51646_ _51644_/Y _51639_/X _51645_/X _85972_/D sky130_fd_sc_hd__a21oi_4
X_70480_ _71706_/A _70483_/B _71815_/B _70480_/X sky130_fd_sc_hd__and3_4
X_82466_ _82595_/CLK _82466_/D _78248_/B sky130_fd_sc_hd__dfxtp_4
X_84205_ _85315_/CLK _84205_/D _65348_/C sky130_fd_sc_hd__dfxtp_4
X_57153_ _57153_/A _57153_/B _57153_/Y sky130_fd_sc_hd__nand2_4
X_81417_ _81575_/CLK _81449_/Q _75976_/B sky130_fd_sc_hd__dfxtp_4
X_69139_ _69135_/X _69137_/X _69138_/X _69139_/X sky130_fd_sc_hd__a21o_4
X_54365_ _85455_/Q _54349_/X _54364_/Y _54365_/Y sky130_fd_sc_hd__o21ai_4
X_85185_ _85249_/CLK _85185_/D _85185_/Q sky130_fd_sc_hd__dfxtp_4
X_51577_ _51590_/A _53105_/B _51577_/Y sky130_fd_sc_hd__nand2_4
X_82397_ _82965_/CLK _82205_/Q _82397_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_381_0_CLK clkbuf_9_190_0_CLK/X _85757_/CLK sky130_fd_sc_hd__clkbuf_1
X_56104_ _56104_/A _56131_/A sky130_fd_sc_hd__buf_2
X_53316_ _53330_/A _53293_/B _53302_/X _52801_/D _53316_/X sky130_fd_sc_hd__and4_4
X_41330_ _41330_/A _41275_/B _41330_/X sky130_fd_sc_hd__or2_4
X_72150_ _83279_/Q _72115_/X _72142_/X _72149_/X _83279_/D sky130_fd_sc_hd__a2bb2oi_4
X_84136_ _82177_/CLK _84136_/D _84136_/Q sky130_fd_sc_hd__dfxtp_4
X_50528_ _50513_/A _48847_/B _50528_/Y sky130_fd_sc_hd__nand2_4
X_57084_ _57084_/A _57084_/B _57084_/Y sky130_fd_sc_hd__nand2_4
X_81348_ _84105_/CLK _76968_/Y _81348_/Q sky130_fd_sc_hd__dfxtp_4
X_54296_ _54314_/A _46662_/A _54296_/Y sky130_fd_sc_hd__nand2_4
X_71101_ _71071_/A _71101_/X sky130_fd_sc_hd__buf_2
X_56035_ _56035_/A _56035_/X sky130_fd_sc_hd__buf_2
X_41261_ _41061_/A _41261_/X sky130_fd_sc_hd__buf_2
X_53247_ _85669_/Q _53225_/X _53246_/Y _53247_/Y sky130_fd_sc_hd__o21ai_4
X_72081_ _72053_/A _49135_/A _72081_/Y sky130_fd_sc_hd__nand2_4
X_84067_ _82648_/CLK _84067_/D _81499_/D sky130_fd_sc_hd__dfxtp_4
X_50459_ _86196_/Q _50437_/X _50458_/Y _50459_/Y sky130_fd_sc_hd__o21ai_4
X_81279_ _81279_/CLK _81311_/Q _76595_/A sky130_fd_sc_hd__dfxtp_4
X_43000_ _42984_/X _42985_/X _40515_/X _67142_/B _42463_/A _43001_/A
+ sky130_fd_sc_hd__o32ai_4
X_71032_ _70997_/A _71178_/A sky130_fd_sc_hd__buf_2
X_83018_ _80670_/CLK _83018_/D _45257_/A sky130_fd_sc_hd__dfxtp_4
X_53178_ _53175_/Y _53163_/X _53177_/X _85683_/D sky130_fd_sc_hd__a21oi_4
X_41192_ _41042_/X _81714_/Q _41191_/X _41192_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_10_396_0_CLK clkbuf_9_198_0_CLK/X _84481_/CLK sky130_fd_sc_hd__clkbuf_1
X_52129_ _65519_/B _52125_/X _52128_/Y _52129_/Y sky130_fd_sc_hd__o21ai_4
X_75840_ _75838_/Y _75840_/B _75841_/A sky130_fd_sc_hd__xor2_4
X_87826_ _87826_/CLK _87826_/D _72769_/A sky130_fd_sc_hd__dfxtp_4
X_57986_ _57947_/X _85710_/Q _57948_/X _57986_/X sky130_fd_sc_hd__o21a_4
X_59725_ _80559_/A _59339_/X _59710_/Y _59724_/Y _84707_/D sky130_fd_sc_hd__a2bb2oi_4
X_44951_ _45819_/A _45590_/B sky130_fd_sc_hd__buf_2
X_56937_ _72978_/A _72771_/A sky130_fd_sc_hd__buf_2
X_75771_ _75771_/A _75771_/Y sky130_fd_sc_hd__inv_2
X_87757_ _87757_/CLK _87757_/D _68528_/B sky130_fd_sc_hd__dfxtp_4
X_72983_ _72977_/X _72981_/X _72982_/X _72983_/X sky130_fd_sc_hd__a21o_4
X_84969_ _86535_/CLK _57614_/Y _84969_/Q sky130_fd_sc_hd__dfxtp_4
X_77510_ _77509_/B _77508_/Y _77505_/Y _77510_/Y sky130_fd_sc_hd__o21ai_4
X_43902_ _43854_/A _43902_/X sky130_fd_sc_hd__buf_2
X_74722_ _74722_/A _74775_/A _71867_/B _70662_/X _74722_/Y sky130_fd_sc_hd__nand4_4
X_86708_ _86711_/CLK _86708_/D _58727_/A sky130_fd_sc_hd__dfxtp_4
X_47670_ _47696_/A _53179_/B _47670_/Y sky130_fd_sc_hd__nand2_4
X_71934_ _56808_/Y _71917_/X _71933_/Y _83323_/D sky130_fd_sc_hd__o21ai_4
X_59656_ _59775_/A _60414_/B sky130_fd_sc_hd__buf_2
X_78490_ _78489_/Y _78490_/Y sky130_fd_sc_hd__inv_2
X_44882_ _45281_/A _44882_/X sky130_fd_sc_hd__buf_2
X_56868_ _56868_/A _56868_/B _56868_/X sky130_fd_sc_hd__and2_4
X_87688_ _87126_/CLK _87688_/D _66828_/B sky130_fd_sc_hd__dfxtp_4
X_46621_ _46609_/Y _46598_/X _46620_/X _46621_/Y sky130_fd_sc_hd__a21oi_4
X_58607_ _58591_/X _85470_/Q _58606_/X _58607_/Y sky130_fd_sc_hd__o21ai_4
X_77441_ _77441_/A _82192_/D _77441_/X sky130_fd_sc_hd__xor2_4
X_43833_ _43802_/A _43833_/X sky130_fd_sc_hd__buf_2
X_55819_ _55816_/X _55818_/X _55819_/X sky130_fd_sc_hd__and2_4
X_86639_ _86640_/CLK _86639_/D _86639_/Q sky130_fd_sc_hd__dfxtp_4
X_74653_ _74638_/X _56633_/X _82997_/Q _74645_/X _74653_/X sky130_fd_sc_hd__a2bb2o_4
X_71865_ _71865_/A _71867_/B _70884_/B _71711_/A _71865_/Y sky130_fd_sc_hd__nor4_4
X_59587_ _59586_/X _59634_/B sky130_fd_sc_hd__buf_2
X_56799_ _44163_/B _56792_/X _56798_/Y _56799_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_440_0_CLK clkbuf_9_441_0_CLK/A clkbuf_9_440_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_49340_ _49352_/A _50862_/B _49340_/Y sky130_fd_sc_hd__nand2_4
X_73604_ _87005_/Q _56550_/X _73603_/X _73604_/Y sky130_fd_sc_hd__o21ai_4
X_46552_ _46531_/A _54071_/B _46552_/Y sky130_fd_sc_hd__nand2_4
X_70816_ _70810_/A _70949_/B _70810_/C _70816_/Y sky130_fd_sc_hd__nand3_4
X_58538_ _58423_/A _58538_/X sky130_fd_sc_hd__buf_2
X_77372_ _77361_/A _77345_/B _77371_/A _77372_/Y sky130_fd_sc_hd__a21oi_4
X_43764_ _40968_/X _43752_/X _87277_/Q _43753_/X _43764_/X sky130_fd_sc_hd__a2bb2o_4
X_74584_ _74600_/A _74584_/X sky130_fd_sc_hd__buf_2
X_40976_ _40512_/X _81721_/Q _40975_/X _40976_/X sky130_fd_sc_hd__o21a_4
X_71796_ _70804_/A _71333_/C _71716_/B _71796_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_334_0_CLK clkbuf_9_167_0_CLK/X _85718_/CLK sky130_fd_sc_hd__clkbuf_1
X_79111_ _82753_/Q _79112_/B sky130_fd_sc_hd__inv_2
X_45503_ _85018_/Q _55555_/B sky130_fd_sc_hd__inv_2
X_76323_ _76309_/X _76321_/Y _76322_/Y _76323_/X sky130_fd_sc_hd__a21o_4
X_88309_ _87068_/CLK _40926_/X _69961_/B sky130_fd_sc_hd__dfxtp_4
X_42715_ _41161_/X _42710_/X _87754_/Q _42711_/X _42715_/X sky130_fd_sc_hd__a2bb2o_4
X_49271_ _49247_/A _49271_/X sky130_fd_sc_hd__buf_2
X_73535_ _73535_/A _65890_/B _73535_/X sky130_fd_sc_hd__and2_4
X_70747_ _70753_/A _70717_/A _70747_/Y sky130_fd_sc_hd__nand2_4
X_46483_ _46423_/X _81197_/Q _46482_/Y _54043_/A sky130_fd_sc_hd__o21ai_4
X_58469_ _84841_/Q _63557_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_964_0_CLK clkbuf_9_482_0_CLK/X _85826_/CLK sky130_fd_sc_hd__clkbuf_1
X_43695_ _43685_/A _43695_/X sky130_fd_sc_hd__buf_2
X_48222_ _48184_/A _50275_/B _48222_/Y sky130_fd_sc_hd__nand2_4
X_60500_ _60440_/A _60500_/Y sky130_fd_sc_hd__inv_2
X_79042_ _79042_/A _79044_/B sky130_fd_sc_hd__inv_2
X_45434_ _45668_/A _45434_/X sky130_fd_sc_hd__buf_2
X_76254_ _76254_/A _76254_/B _76252_/Y _76255_/A sky130_fd_sc_hd__nand3_4
X_42646_ _42645_/Y _42646_/Y sky130_fd_sc_hd__inv_2
X_61480_ _61355_/A _61482_/A sky130_fd_sc_hd__buf_2
X_73466_ _69932_/B _73250_/X _73464_/X _73465_/Y _73466_/X sky130_fd_sc_hd__a211o_4
X_70678_ _70552_/Y _70679_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_455_0_CLK clkbuf_9_455_0_CLK/A clkbuf_9_455_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_75205_ _75205_/A _75205_/Y sky130_fd_sc_hd__inv_2
X_48153_ _48153_/A _50389_/B sky130_fd_sc_hd__buf_2
X_60431_ _60430_/Y _60438_/A sky130_fd_sc_hd__buf_2
X_72417_ _72417_/A _72417_/X sky130_fd_sc_hd__buf_2
X_45365_ _45365_/A _45381_/B _45365_/Y sky130_fd_sc_hd__nand2_4
X_76185_ _76187_/A _81553_/Q _76186_/A sky130_fd_sc_hd__nor2_4
X_42577_ _42573_/X _42574_/X _40831_/X _69734_/A _42540_/X _42578_/A
+ sky130_fd_sc_hd__o32ai_4
X_73397_ _43190_/Y _73298_/X _73251_/X _73396_/Y _73397_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_349_0_CLK clkbuf_9_174_0_CLK/X _85745_/CLK sky130_fd_sc_hd__clkbuf_1
X_47104_ _47103_/Y _52857_/D sky130_fd_sc_hd__buf_2
X_44316_ _58631_/A _44031_/X _57811_/A _58007_/A _44253_/X _44316_/X
+ sky130_fd_sc_hd__a41o_4
X_75136_ _75133_/Y _75135_/Y _81030_/D sky130_fd_sc_hd__xnor2_4
X_63150_ _63150_/A _63113_/B _63103_/C _63149_/X _63150_/X sky130_fd_sc_hd__or4_4
X_41528_ _41261_/X _81171_/Q _41527_/X _41529_/A sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_979_0_CLK clkbuf_9_489_0_CLK/X _85554_/CLK sky130_fd_sc_hd__clkbuf_1
X_48084_ _74129_/B _48049_/X _48083_/Y _48084_/Y sky130_fd_sc_hd__o21ai_4
X_60362_ _60362_/A _62678_/A sky130_fd_sc_hd__buf_2
X_72348_ _86606_/Q _72348_/B _72348_/Y sky130_fd_sc_hd__nor2_4
X_45296_ _45288_/X _45292_/Y _45295_/Y _45296_/Y sky130_fd_sc_hd__a21oi_4
X_62101_ _62033_/A _62101_/X sky130_fd_sc_hd__buf_2
X_47035_ _47081_/A _47035_/X sky130_fd_sc_hd__buf_2
X_44247_ _44247_/A _58602_/A sky130_fd_sc_hd__buf_2
X_63081_ _63081_/A _63081_/B _63081_/C _63033_/D _63081_/X sky130_fd_sc_hd__or4_4
X_75067_ _75067_/A _75067_/B _75067_/Y sky130_fd_sc_hd__nand2_4
X_79944_ _79944_/A _79945_/B _79945_/A _79944_/Y sky130_fd_sc_hd__nand3_4
X_41459_ _81185_/Q _41459_/B _41459_/X sky130_fd_sc_hd__or2_4
X_60293_ _60105_/X _60317_/A sky130_fd_sc_hd__buf_2
X_72279_ _72137_/X _72277_/Y _72278_/Y _72194_/X _72141_/X _72279_/X
+ sky130_fd_sc_hd__o32a_4
X_62032_ _61348_/A _62033_/A sky130_fd_sc_hd__buf_2
X_74018_ _74016_/X _85614_/Q _73903_/X _74017_/X _74018_/X sky130_fd_sc_hd__a211o_4
X_44178_ _44146_/A _45924_/A sky130_fd_sc_hd__buf_2
X_79875_ _79875_/A _79875_/B _79875_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_902_0_CLK clkbuf_9_451_0_CLK/X _82538_/CLK sky130_fd_sc_hd__clkbuf_1
X_43129_ _43129_/A _43129_/X sky130_fd_sc_hd__buf_2
X_66840_ _68721_/A _66840_/X sky130_fd_sc_hd__buf_2
X_78826_ _82628_/Q _78828_/B sky130_fd_sc_hd__inv_2
X_48986_ _48986_/A _49009_/B _48986_/Y sky130_fd_sc_hd__nor2_4
X_47937_ _47946_/A _47937_/B _47937_/X sky130_fd_sc_hd__and2_4
X_66771_ _66771_/A _66770_/X _66771_/Y sky130_fd_sc_hd__nand2_4
X_78757_ _78758_/A _78758_/C _78756_/Y _78770_/B sky130_fd_sc_hd__a21o_4
X_63983_ _60906_/X _64046_/C sky130_fd_sc_hd__buf_2
X_75969_ _75964_/A _75969_/B _75969_/Y sky130_fd_sc_hd__nand2_4
X_68510_ _68409_/A _88270_/Q _68510_/X sky130_fd_sc_hd__and2_4
X_65722_ _64683_/A _65725_/B sky130_fd_sc_hd__buf_2
X_77708_ _81952_/Q _77707_/A _77708_/Y sky130_fd_sc_hd__xnor2_4
X_62934_ _58187_/X _62808_/X _62827_/X _62818_/X _62933_/X _62934_/Y
+ sky130_fd_sc_hd__a41oi_4
Xclkbuf_10_917_0_CLK clkbuf_9_458_0_CLK/X _86549_/CLK sky130_fd_sc_hd__clkbuf_1
X_69490_ _81384_/D _69439_/X _69489_/X _83920_/D sky130_fd_sc_hd__a21bo_4
X_47868_ _82366_/Q _47869_/A sky130_fd_sc_hd__inv_2
X_78688_ _82523_/Q _82779_/D _82491_/D sky130_fd_sc_hd__xor2_4
X_49607_ _49580_/A _49607_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_6_0_CLK clkbuf_9_3_0_CLK/X _85177_/CLK sky130_fd_sc_hd__clkbuf_1
X_68441_ _88112_/Q _68069_/X _68439_/X _68440_/Y _68441_/X sky130_fd_sc_hd__a211o_4
X_46819_ _46915_/A _46830_/A sky130_fd_sc_hd__buf_2
X_65653_ _65014_/X _65653_/B _65017_/X _65664_/A sky130_fd_sc_hd__nand3_4
X_77639_ _77633_/X _77636_/Y _77634_/Y _77639_/Y sky130_fd_sc_hd__nand3_4
X_62865_ _62863_/X _62838_/X _62864_/Y _84376_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_408_0_CLK clkbuf_9_409_0_CLK/A clkbuf_9_408_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_47799_ _47799_/A _51728_/B _47799_/Y sky130_fd_sc_hd__nand2_4
X_64604_ _64599_/X _83313_/Q _64600_/X _64603_/X _64604_/X sky130_fd_sc_hd__a211o_4
X_49538_ _49536_/Y _49514_/X _49537_/X _49538_/Y sky130_fd_sc_hd__a21oi_4
X_61816_ _61805_/X _61807_/X _61814_/Y _58166_/A _61815_/X _61816_/Y
+ sky130_fd_sc_hd__o32ai_4
X_80650_ _74811_/X _74714_/Y DATA_FROM_HASH[7] sky130_fd_sc_hd__ebufn_2
X_68372_ _87007_/Q _68059_/X _68370_/X _68371_/X _68372_/X sky130_fd_sc_hd__a211o_4
X_65584_ _65769_/A _65584_/B _65584_/X sky130_fd_sc_hd__and2_4
X_62796_ _60179_/A _62819_/C sky130_fd_sc_hd__buf_2
X_67323_ _67318_/X _67321_/X _67322_/X _67323_/X sky130_fd_sc_hd__a21o_4
X_79309_ _84798_/Q _84118_/Q _79309_/X sky130_fd_sc_hd__xor2_4
X_64535_ _64545_/A _64535_/B _64545_/C _64535_/X sky130_fd_sc_hd__and3_4
X_49469_ _49002_/A _49496_/A sky130_fd_sc_hd__buf_2
X_61747_ _59721_/A _61747_/X sky130_fd_sc_hd__buf_2
X_80581_ _80596_/A _80596_/B _80581_/X sky130_fd_sc_hd__xor2_4
X_51500_ _51497_/Y _51477_/X _51499_/X _85999_/D sky130_fd_sc_hd__a21oi_4
X_82320_ _82327_/CLK _77103_/B _82320_/Q sky130_fd_sc_hd__dfxtp_4
X_67254_ _87107_/Q _67230_/X _67160_/X _67253_/X _67254_/X sky130_fd_sc_hd__a211o_4
X_52480_ _52476_/A _52480_/B _52480_/Y sky130_fd_sc_hd__nand2_4
X_64466_ _64494_/A _64466_/B _64207_/A _64466_/X sky130_fd_sc_hd__and3_4
X_61678_ _61678_/A _61678_/Y sky130_fd_sc_hd__inv_2
X_66205_ _66065_/A _66205_/X sky130_fd_sc_hd__buf_2
X_51431_ _51430_/X _52959_/B _51431_/Y sky130_fd_sc_hd__nand2_4
X_63417_ _63417_/A _63465_/D sky130_fd_sc_hd__buf_2
X_82251_ _82251_/CLK _82251_/D _82251_/Q sky130_fd_sc_hd__dfxtp_4
X_60629_ _60628_/Y _60629_/Y sky130_fd_sc_hd__inv_2
X_67185_ _67181_/X _67184_/X _67113_/X _67185_/Y sky130_fd_sc_hd__a21oi_4
X_64397_ _64389_/Y _64396_/X _64386_/X _64397_/X sky130_fd_sc_hd__o21a_4
X_81202_ _81198_/CLK _75014_/X _49039_/A sky130_fd_sc_hd__dfxtp_4
X_54150_ _85495_/Q _54140_/X _54149_/Y _54150_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_6_8_0_CLK clkbuf_6_9_0_CLK/A clkbuf_6_8_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_66136_ _66020_/X _66134_/Y _66135_/Y _66136_/Y sky130_fd_sc_hd__o21ai_4
X_51362_ _51259_/A _51362_/X sky130_fd_sc_hd__buf_2
X_63348_ _63348_/A _63250_/X _63348_/Y sky130_fd_sc_hd__nor2_4
X_82182_ _86655_/CLK _82182_/D _82374_/D sky130_fd_sc_hd__dfxtp_4
X_53101_ _53115_/A _53101_/B _53101_/Y sky130_fd_sc_hd__nand2_4
X_50313_ _50491_/A _50313_/X sky130_fd_sc_hd__buf_2
X_81133_ _81130_/CLK _80757_/Q _40700_/A sky130_fd_sc_hd__dfxtp_4
X_54081_ _54068_/X _52563_/B _54081_/Y sky130_fd_sc_hd__nand2_4
X_66067_ _66063_/Y _66065_/X _66066_/X _66067_/X sky130_fd_sc_hd__a21o_4
X_51293_ _86038_/Q _51285_/X _51292_/Y _51293_/Y sky130_fd_sc_hd__o21ai_4
X_63279_ _58279_/Y _63250_/X _59423_/Y _60493_/X _63279_/X sky130_fd_sc_hd__o22a_4
X_86990_ _86989_/CLK _86990_/D _86990_/Q sky130_fd_sc_hd__dfxtp_4
X_53032_ _53026_/Y _53028_/X _53031_/X _53032_/Y sky130_fd_sc_hd__a21oi_4
X_65018_ _65014_/X _64888_/B _65017_/X _65018_/Y sky130_fd_sc_hd__nand3_4
X_50244_ _53874_/A _74509_/C sky130_fd_sc_hd__buf_2
X_85941_ _82768_/CLK _51816_/Y _85941_/Q sky130_fd_sc_hd__dfxtp_4
X_81064_ _80681_/CLK _81096_/Q _75157_/B sky130_fd_sc_hd__dfxtp_4
X_80015_ _84930_/Q _84178_/Q _80015_/Y sky130_fd_sc_hd__nand2_4
X_57840_ _57838_/X _86010_/Q _57839_/X _57840_/Y sky130_fd_sc_hd__o21ai_4
X_69826_ _69865_/A _69826_/B _69826_/X sky130_fd_sc_hd__and2_4
X_50175_ _50131_/A _72079_/B _50175_/X sky130_fd_sc_hd__and2_4
X_85872_ _83562_/CLK _85872_/D _85872_/Q sky130_fd_sc_hd__dfxtp_4
X_87611_ _82888_/CLK _43001_/Y _67142_/B sky130_fd_sc_hd__dfxtp_4
X_84823_ _84823_/CLK _58545_/X _58543_/A sky130_fd_sc_hd__dfxtp_4
X_57771_ _58796_/A _72476_/B sky130_fd_sc_hd__buf_2
X_69757_ _87057_/Q _69664_/X _69665_/X _69756_/X _69758_/B sky130_fd_sc_hd__a211o_4
X_54983_ _54964_/A _54978_/X _54974_/C _47567_/A _54983_/X sky130_fd_sc_hd__and4_4
X_66969_ _66947_/X _66958_/Y _66910_/X _66968_/Y _66969_/X sky130_fd_sc_hd__a211o_4
X_59510_ _57754_/X _69814_/A sky130_fd_sc_hd__buf_2
X_56722_ _56684_/C _56721_/Y _56723_/B sky130_fd_sc_hd__xor2_4
X_68708_ _68735_/A _68708_/B _68708_/X sky130_fd_sc_hd__and2_4
X_87542_ _87542_/CLK _87542_/D _43199_/A sky130_fd_sc_hd__dfxtp_4
X_53934_ _53949_/A _50719_/B _53934_/Y sky130_fd_sc_hd__nand2_4
X_84754_ _84757_/CLK _84754_/D _84754_/Q sky130_fd_sc_hd__dfxtp_4
X_81966_ _82299_/CLK _81966_/D _81966_/Q sky130_fd_sc_hd__dfxtp_4
X_69688_ _88074_/Q _69607_/X _68617_/X _69687_/Y _69688_/X sky130_fd_sc_hd__a211o_4
X_59441_ _59417_/X _83340_/Q _59440_/Y _59441_/X sky130_fd_sc_hd__o21a_4
X_83705_ _85428_/CLK _70767_/Y _47069_/A sky130_fd_sc_hd__dfxtp_4
X_56653_ _56808_/A _83322_/Q _56653_/Y sky130_fd_sc_hd__nand2_4
X_80917_ _81507_/CLK _80917_/D _80917_/Q sky130_fd_sc_hd__dfxtp_4
X_68639_ _43057_/A _68636_/X _68517_/X _68638_/X _68639_/X sky130_fd_sc_hd__a211o_4
X_87473_ _87473_/CLK _87473_/D _87473_/Q sky130_fd_sc_hd__dfxtp_4
X_53865_ _53786_/A _49055_/A _53865_/Y sky130_fd_sc_hd__nand2_4
X_84685_ _84713_/CLK _59865_/Y _80308_/B sky130_fd_sc_hd__dfxtp_4
X_81897_ _82047_/CLK _77337_/X _82305_/D sky130_fd_sc_hd__dfxtp_4
X_55604_ _55603_/X _56564_/A sky130_fd_sc_hd__buf_2
X_86424_ _86424_/CLK _49254_/Y _86424_/Q sky130_fd_sc_hd__dfxtp_4
X_52816_ _53221_/A _52845_/A sky130_fd_sc_hd__buf_2
X_40830_ _40324_/X _82868_/Q _40829_/X _40831_/A sky130_fd_sc_hd__o21a_4
X_71650_ _71650_/A _71217_/B _71644_/C _71650_/Y sky130_fd_sc_hd__nand3_4
X_83636_ _86424_/CLK _83636_/D _83636_/Q sky130_fd_sc_hd__dfxtp_4
X_59372_ _59238_/X _59372_/B _59372_/Y sky130_fd_sc_hd__nor2_4
X_56584_ _56583_/X _56584_/X sky130_fd_sc_hd__buf_2
X_80848_ _80849_/CLK _80880_/Q _74960_/C sky130_fd_sc_hd__dfxtp_4
X_53796_ _53791_/A _71972_/B _53796_/Y sky130_fd_sc_hd__nand2_4
X_70601_ DATA_TO_HASH[5] _70771_/A sky130_fd_sc_hd__buf_2
X_58323_ _58322_/Y _58326_/B _58323_/Y sky130_fd_sc_hd__nand2_4
X_55535_ _45558_/A _55531_/X _55533_/X _55534_/X _55536_/D sky130_fd_sc_hd__a211o_4
X_86355_ _85428_/CLK _49616_/Y _86355_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_2_0_1_CLK clkbuf_2_0_1_CLK/A clkbuf_2_0_2_CLK/A sky130_fd_sc_hd__clkbuf_1
X_40761_ _40698_/X _40927_/A _40760_/X _40762_/A sky130_fd_sc_hd__o21a_4
X_52747_ _52745_/Y _52728_/X _52746_/X _52747_/Y sky130_fd_sc_hd__a21oi_4
X_71581_ _71581_/A _71581_/X sky130_fd_sc_hd__buf_2
X_83567_ _86500_/CLK _71224_/Y _83567_/Q sky130_fd_sc_hd__dfxtp_4
X_80779_ _80754_/CLK _75661_/Y _80779_/Q sky130_fd_sc_hd__dfxtp_4
X_42500_ _42486_/X _42472_/X _40673_/X _68746_/B _42489_/X _87844_/D
+ sky130_fd_sc_hd__o32ai_4
X_73320_ _73320_/A _73438_/B _73320_/Y sky130_fd_sc_hd__nor2_4
X_85306_ _85180_/CLK _56042_/Y _56041_/C sky130_fd_sc_hd__dfxtp_4
X_70532_ _70531_/Y _70532_/Y sky130_fd_sc_hd__inv_2
X_58254_ _58254_/A _58254_/Y sky130_fd_sc_hd__inv_2
X_82518_ _82518_/CLK _79117_/Y _82518_/Q sky130_fd_sc_hd__dfxtp_4
X_55466_ _55461_/X _55465_/X _55466_/X sky130_fd_sc_hd__and2_4
X_43480_ _43472_/X _43475_/X _41688_/X _87401_/Q _43479_/X _43480_/Y
+ sky130_fd_sc_hd__o32ai_4
X_86286_ _86610_/CLK _86286_/D _72347_/B sky130_fd_sc_hd__dfxtp_4
X_52678_ _85774_/Q _52656_/X _52677_/Y _52678_/Y sky130_fd_sc_hd__o21ai_4
X_40692_ _40687_/X _40688_/X _40691_/X _88353_/Q _40683_/X _40692_/Y
+ sky130_fd_sc_hd__o32ai_4
X_83498_ _83498_/CLK _71440_/X _83498_/Q sky130_fd_sc_hd__dfxtp_4
X_57205_ _57179_/A _85063_/Q _57205_/Y sky130_fd_sc_hd__nand2_4
X_88025_ _87776_/CLK _88025_/D _88025_/Q sky130_fd_sc_hd__dfxtp_4
X_54417_ _54399_/X _54417_/B _54402_/C _54417_/D _54417_/X sky130_fd_sc_hd__and4_4
X_42431_ _42417_/X _42430_/X _40515_/X _87867_/Q _41967_/A _42432_/A
+ sky130_fd_sc_hd__o32ai_4
X_73251_ _56934_/X _73251_/X sky130_fd_sc_hd__buf_2
X_85237_ _86900_/CLK _85237_/D _55874_/B sky130_fd_sc_hd__dfxtp_4
X_51629_ _51629_/A _51629_/X sky130_fd_sc_hd__buf_2
X_70463_ DATA_TO_HASH[7] _71672_/C sky130_fd_sc_hd__buf_2
X_58185_ _57677_/X _58181_/Y _58184_/Y _58185_/Y sky130_fd_sc_hd__a21oi_4
X_82449_ _82452_/CLK _79141_/X _82449_/Q sky130_fd_sc_hd__dfxtp_4
X_55397_ _55164_/X _55397_/Y sky130_fd_sc_hd__inv_2
X_72202_ _72198_/Y _72200_/Y _72201_/X _72202_/X sky130_fd_sc_hd__a21o_4
X_45150_ _55833_/B _45134_/X _45116_/X _45150_/X sky130_fd_sc_hd__o21a_4
X_57136_ _57132_/Y _57135_/Y _46178_/X _57136_/Y sky130_fd_sc_hd__o21ai_4
X_42362_ _41745_/X _42356_/X _87901_/Q _42357_/X _87901_/D sky130_fd_sc_hd__a2bb2o_4
X_54348_ _54342_/Y _54338_/X _54347_/X _54348_/Y sky130_fd_sc_hd__a21oi_4
X_73182_ _72988_/X _86193_/Q _72985_/X _73181_/X _73182_/X sky130_fd_sc_hd__a211o_4
X_85168_ _85168_/CLK _85168_/D _56510_/C sky130_fd_sc_hd__dfxtp_4
X_70394_ _70819_/A _70786_/A sky130_fd_sc_hd__buf_2
X_44101_ _44101_/A _44102_/A sky130_fd_sc_hd__buf_2
X_41313_ _41312_/X _41307_/X _67456_/B _41308_/X _88238_/D sky130_fd_sc_hd__a2bb2o_4
X_72133_ _72123_/X _85696_/Q _59334_/X _72133_/X sky130_fd_sc_hd__o21a_4
X_84119_ _84119_/CLK _84119_/D _82735_/D sky130_fd_sc_hd__dfxtp_4
X_45081_ _45081_/A _45082_/A sky130_fd_sc_hd__inv_2
X_57067_ _56893_/Y _57289_/B _56866_/A _56860_/X _57067_/Y sky130_fd_sc_hd__a22oi_4
X_42293_ _41560_/X _42290_/X _87936_/Q _42291_/X _87936_/D sky130_fd_sc_hd__a2bb2o_4
X_54279_ _54286_/A _54298_/B _54286_/C _46638_/A _54279_/X sky130_fd_sc_hd__and4_4
X_77990_ _77971_/X _77977_/A _77975_/Y _77990_/Y sky130_fd_sc_hd__a21oi_4
X_85099_ _85096_/CLK _57031_/Y _57027_/A sky130_fd_sc_hd__dfxtp_4
X_44032_ _58834_/A _57811_/A sky130_fd_sc_hd__buf_2
X_56018_ _55688_/X _56016_/X _56017_/Y _56018_/Y sky130_fd_sc_hd__o21ai_4
X_41244_ _41242_/X _40722_/A _41243_/X _41244_/X sky130_fd_sc_hd__o21a_4
X_76941_ _76939_/X _76953_/A _76942_/B _76941_/Y sky130_fd_sc_hd__a21oi_4
X_72064_ _49099_/A _72043_/X _72048_/X _72064_/X sky130_fd_sc_hd__and3_4
X_71015_ _71263_/D _71016_/A sky130_fd_sc_hd__buf_2
X_48840_ _48840_/A _48840_/X sky130_fd_sc_hd__buf_2
X_79660_ _79660_/A _79659_/Y _79660_/X sky130_fd_sc_hd__xor2_4
X_41175_ _41112_/X _41113_/X _41174_/X _68686_/B _41088_/X _41176_/A
+ sky130_fd_sc_hd__o32ai_4
X_76872_ _76872_/A _81466_/D _81562_/D sky130_fd_sc_hd__xor2_4
X_78611_ _78611_/A _82679_/D _78616_/A sky130_fd_sc_hd__nor2_4
X_75823_ _75811_/A _75815_/Y _75823_/C _75824_/B sky130_fd_sc_hd__nand3_4
X_87809_ _87553_/CLK _87809_/D _69804_/A sky130_fd_sc_hd__dfxtp_4
X_48771_ _52156_/A _48770_/X _48786_/C _48771_/X sky130_fd_sc_hd__and3_4
X_79591_ _79569_/Y _79573_/B _79590_/Y _79591_/Y sky130_fd_sc_hd__a21oi_4
X_45983_ _45980_/X _44865_/X _40425_/X _66810_/B _45982_/X _45984_/A
+ sky130_fd_sc_hd__o32ai_4
X_57969_ _57964_/Y _57968_/Y _57909_/X _57969_/X sky130_fd_sc_hd__a21o_4
X_47722_ _47722_/A _53207_/D sky130_fd_sc_hd__buf_2
X_59708_ _59544_/A _59741_/A sky130_fd_sc_hd__buf_2
X_78542_ _78540_/X _78510_/Y _78541_/Y _78542_/X sky130_fd_sc_hd__a21o_4
X_44934_ _80670_/Q _45705_/A sky130_fd_sc_hd__buf_2
X_75754_ _75743_/Y _75754_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_40_0_CLK clkbuf_9_20_0_CLK/X _82998_/CLK sky130_fd_sc_hd__clkbuf_1
X_60980_ _60908_/X _61012_/C _59691_/X _60980_/Y sky130_fd_sc_hd__a21oi_4
X_72966_ _72966_/A _72965_/X _72967_/B sky130_fd_sc_hd__nand2_4
X_74705_ _74673_/A _45876_/A _74705_/Y sky130_fd_sc_hd__nand2_4
X_47653_ _47653_/A _55031_/D sky130_fd_sc_hd__inv_2
X_71917_ _71916_/Y _71917_/X sky130_fd_sc_hd__buf_2
X_59639_ _59639_/A _60403_/A sky130_fd_sc_hd__buf_2
X_78473_ _78473_/A _78472_/X _78473_/X sky130_fd_sc_hd__xor2_4
X_44865_ _46001_/A _44865_/X sky130_fd_sc_hd__buf_2
X_75685_ _75685_/A _75684_/Y _75686_/B sky130_fd_sc_hd__xor2_4
X_72897_ _43126_/Y _72895_/X _72858_/X _72896_/Y _72897_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_273_0_CLK clkbuf_9_136_0_CLK/X _84951_/CLK sky130_fd_sc_hd__clkbuf_1
X_46604_ _51396_/A _46487_/B _46603_/X _46604_/X sky130_fd_sc_hd__and3_4
X_77424_ _77423_/A _82096_/D _77424_/Y sky130_fd_sc_hd__nand2_4
X_43816_ _41104_/X _43801_/X _69544_/B _43802_/X _87253_/D sky130_fd_sc_hd__a2bb2o_4
X_74636_ _45952_/X _56577_/Y _45448_/A _74633_/X _83006_/D sky130_fd_sc_hd__a2bb2o_4
X_62650_ _62949_/B _62650_/X sky130_fd_sc_hd__buf_2
X_47584_ _72193_/A _47570_/X _47583_/Y _47584_/Y sky130_fd_sc_hd__o21ai_4
X_71848_ _71847_/Y _71848_/X sky130_fd_sc_hd__buf_2
X_44796_ _44512_/A _41887_/A _41423_/X _86950_/Q _44516_/A _44797_/A
+ sky130_fd_sc_hd__o32ai_4
X_49323_ _49321_/Y _49271_/X _49322_/Y _86410_/D sky130_fd_sc_hd__a21boi_4
X_61601_ _61600_/Y _61601_/Y sky130_fd_sc_hd__inv_2
X_46535_ _46434_/A _50852_/B _46535_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_55_0_CLK clkbuf_9_27_0_CLK/X _85096_/CLK sky130_fd_sc_hd__clkbuf_1
X_77355_ _77354_/B _77354_/A _77360_/C sky130_fd_sc_hd__nand2_4
X_43747_ _40921_/X _43736_/X _73487_/A _43737_/X _43747_/X sky130_fd_sc_hd__a2bb2o_4
X_62581_ _62579_/Y _62561_/B _62580_/Y _62581_/Y sky130_fd_sc_hd__nand3_4
X_74567_ _45046_/Y _74551_/X _74566_/X _74567_/Y sky130_fd_sc_hd__o21ai_4
X_40959_ _40959_/A _40959_/X sky130_fd_sc_hd__buf_2
X_71779_ _71779_/A _71779_/B _70986_/A _71779_/X sky130_fd_sc_hd__and3_4
Xclkbuf_9_394_0_CLK clkbuf_9_395_0_CLK/A clkbuf_9_394_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_64320_ _64319_/X _64320_/B _64274_/X _64320_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_201_0_CLK clkbuf_8_201_0_CLK/A clkbuf_9_402_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_76306_ _76306_/A _76305_/Y _76306_/X sky130_fd_sc_hd__and2_4
X_49254_ _49252_/Y _49247_/X _49253_/Y _49254_/Y sky130_fd_sc_hd__a21boi_4
X_61532_ _61532_/A _61532_/Y sky130_fd_sc_hd__inv_2
X_73518_ _73515_/X _73517_/X _72949_/X _73521_/A sky130_fd_sc_hd__a21o_4
X_46466_ _46421_/A _51328_/B _46466_/Y sky130_fd_sc_hd__nand2_4
X_77286_ _77286_/A _77286_/Y sky130_fd_sc_hd__inv_2
X_43678_ _40767_/X _43671_/X _87315_/Q _43673_/X _43678_/X sky130_fd_sc_hd__a2bb2o_4
X_74498_ _74496_/Y _74492_/X _74497_/X _83054_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_288_0_CLK clkbuf_9_144_0_CLK/X _84903_/CLK sky130_fd_sc_hd__clkbuf_1
X_48205_ _48204_/X _50260_/B _48205_/Y sky130_fd_sc_hd__nand2_4
X_79025_ _79012_/A _79023_/Y _79024_/X _79025_/Y sky130_fd_sc_hd__o21ai_4
X_45417_ _85152_/Q _45876_/B _44919_/X _45417_/Y sky130_fd_sc_hd__o21ai_4
X_76237_ _76231_/Y _76233_/Y _76235_/Y _76237_/Y sky130_fd_sc_hd__nand3_4
X_64251_ _59460_/A _64249_/X _64250_/Y _64251_/Y sky130_fd_sc_hd__o21ai_4
X_42629_ _42743_/A _52754_/A sky130_fd_sc_hd__buf_2
X_49185_ _53932_/B _50716_/B sky130_fd_sc_hd__buf_2
X_61463_ _61429_/A _61461_/X _61482_/C _61463_/Y sky130_fd_sc_hd__nand3_4
X_73449_ _72908_/A _73449_/X sky130_fd_sc_hd__buf_2
X_46397_ _86740_/Q _46364_/X _46396_/Y _46397_/Y sky130_fd_sc_hd__o21ai_4
X_63202_ _63154_/X _64411_/B _63165_/X _63192_/D _63202_/X sky130_fd_sc_hd__and4_4
X_48136_ _48136_/A _48136_/B _48136_/X sky130_fd_sc_hd__or2_4
X_60414_ _60413_/X _60414_/B _60414_/Y sky130_fd_sc_hd__nand2_4
X_45348_ _45714_/A _45348_/X sky130_fd_sc_hd__buf_2
X_64182_ _62174_/X _64182_/B _64182_/C _64182_/D _64182_/Y sky130_fd_sc_hd__nand4_4
X_76168_ _76166_/X _76168_/B _76169_/A sky130_fd_sc_hd__and2_4
X_61394_ _61394_/A _61394_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_216_0_CLK clkbuf_8_217_0_CLK/A clkbuf_8_216_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_211_0_CLK clkbuf_9_105_0_CLK/X _84493_/CLK sky130_fd_sc_hd__clkbuf_1
X_63133_ _63097_/A _64343_/B _63108_/C _63121_/D _63133_/X sky130_fd_sc_hd__and4_4
X_75119_ _75116_/X _75120_/B _75120_/A _75119_/X sky130_fd_sc_hd__a21o_4
X_60345_ _60105_/X _60477_/A sky130_fd_sc_hd__buf_2
X_48067_ _48067_/A _52050_/A sky130_fd_sc_hd__buf_2
X_45279_ _45277_/X _61617_/B _45219_/X _45279_/Y sky130_fd_sc_hd__o21ai_4
X_68990_ _69648_/A _42525_/Y _68990_/Y sky130_fd_sc_hd__nor2_4
X_76099_ _76099_/A _76099_/B _76100_/B sky130_fd_sc_hd__xnor2_4
Xclkbuf_10_841_0_CLK clkbuf_9_420_0_CLK/X _82746_/CLK sky130_fd_sc_hd__clkbuf_1
X_47018_ _59118_/A _47004_/X _47017_/Y _47018_/Y sky130_fd_sc_hd__o21ai_4
X_67941_ _67937_/X _67940_/X _67917_/X _67941_/X sky130_fd_sc_hd__a21o_4
X_63064_ _63039_/A _64276_/C _63028_/X _63014_/D _63064_/X sky130_fd_sc_hd__and4_4
X_79927_ _79927_/A _79927_/B _79928_/B sky130_fd_sc_hd__nand2_4
X_60276_ _60331_/D _60273_/X _60275_/X _60344_/B _60276_/Y sky130_fd_sc_hd__a22oi_4
Xclkbuf_9_332_0_CLK clkbuf_8_166_0_CLK/X clkbuf_9_332_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_62015_ _61957_/A _62015_/B _62012_/Y _62015_/D _62015_/Y sky130_fd_sc_hd__nand4_4
X_67872_ _68370_/A _67872_/X sky130_fd_sc_hd__buf_2
X_79858_ _79812_/Y _79852_/X _79857_/Y _79858_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_226_0_CLK clkbuf_9_113_0_CLK/X _81111_/CLK sky130_fd_sc_hd__clkbuf_1
X_69611_ _69611_/A _69611_/X sky130_fd_sc_hd__buf_2
X_66823_ _66823_/A _88201_/Q _66823_/X sky130_fd_sc_hd__and2_4
X_78809_ _78809_/A _82546_/Q _78809_/Y sky130_fd_sc_hd__nand2_4
X_48969_ _48969_/A _71998_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_856_0_CLK clkbuf_9_428_0_CLK/X _85800_/CLK sky130_fd_sc_hd__clkbuf_1
X_79789_ _79790_/B _79776_/Y _79789_/X sky130_fd_sc_hd__or2_4
X_81820_ _81275_/CLK _81628_/Q _81820_/Q sky130_fd_sc_hd__dfxtp_4
X_69542_ _69956_/A _69542_/B _69542_/X sky130_fd_sc_hd__and2_4
X_66754_ _66750_/X _66753_/X _66658_/X _66754_/Y sky130_fd_sc_hd__a21oi_4
X_51980_ _73780_/B _51960_/X _51979_/Y _51980_/Y sky130_fd_sc_hd__o21ai_4
X_63966_ _58528_/A _64191_/B _60889_/X _64191_/D _63966_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_9_347_0_CLK clkbuf_9_347_0_CLK/A clkbuf_9_347_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_65705_ _65638_/X _85583_/Q _65669_/X _65704_/X _65705_/X sky130_fd_sc_hd__a211o_4
X_50931_ _50927_/Y _50928_/X _50930_/X _86105_/D sky130_fd_sc_hd__a21oi_4
X_62917_ _62081_/B _64473_/A sky130_fd_sc_hd__inv_2
X_81751_ _81756_/CLK _76074_/B _41686_/B sky130_fd_sc_hd__dfxtp_4
X_69473_ _87015_/Q _69414_/X _69430_/X _69472_/X _69473_/X sky130_fd_sc_hd__a211o_4
X_66685_ _66681_/X _66684_/X _66411_/A _66685_/Y sky130_fd_sc_hd__a21oi_4
X_63897_ _63848_/X _63849_/X _63897_/C _63897_/Y sky130_fd_sc_hd__nor3_4
X_80702_ _82211_/CLK _80702_/D _80702_/Q sky130_fd_sc_hd__dfxtp_4
X_68424_ _68420_/X _68423_/X _68400_/X _68424_/Y sky130_fd_sc_hd__a21oi_4
X_53650_ _53648_/Y _53619_/X _53649_/X _85595_/D sky130_fd_sc_hd__a21oi_4
X_65636_ _65667_/A _85875_/Q _65636_/X sky130_fd_sc_hd__and2_4
X_84470_ _82452_/CLK _61567_/Y _79138_/B sky130_fd_sc_hd__dfxtp_4
X_50862_ _50857_/X _50862_/B _50862_/Y sky130_fd_sc_hd__nand2_4
X_62848_ _62847_/X _63198_/A _62848_/C _62880_/D _62848_/X sky130_fd_sc_hd__and4_4
X_81682_ _81682_/CLK _80098_/X _81682_/Q sky130_fd_sc_hd__dfxtp_4
X_52601_ _52515_/X _52601_/X sky130_fd_sc_hd__buf_2
X_83421_ _83421_/CLK _83421_/D _83421_/Q sky130_fd_sc_hd__dfxtp_4
X_80633_ _80624_/A _80623_/X _80633_/C _80633_/Y sky130_fd_sc_hd__nand3_4
X_68355_ _65381_/A _88275_/Q _68355_/X sky130_fd_sc_hd__and2_4
X_53581_ _53622_/A _57617_/B _53581_/Y sky130_fd_sc_hd__nand2_4
X_65567_ _65562_/X _65565_/X _65566_/X _66044_/A sky130_fd_sc_hd__a21o_4
X_50793_ _50787_/X _46407_/X _50793_/Y sky130_fd_sc_hd__nand2_4
X_62779_ _62893_/A _62779_/X sky130_fd_sc_hd__buf_2
X_55320_ _44059_/X _55320_/B _55320_/Y sky130_fd_sc_hd__nor2_4
X_67306_ _67259_/A _87604_/Q _67306_/X sky130_fd_sc_hd__and2_4
X_86140_ _86139_/CLK _50756_/Y _86140_/Q sky130_fd_sc_hd__dfxtp_4
X_52532_ _52496_/A _52532_/X sky130_fd_sc_hd__buf_2
X_64518_ _64511_/Y _64517_/X _64442_/X _64518_/X sky130_fd_sc_hd__o21a_4
X_83352_ _83480_/CLK _83352_/D _83352_/Q sky130_fd_sc_hd__dfxtp_4
X_80564_ _80561_/X _80564_/B _82267_/D sky130_fd_sc_hd__xnor2_4
XPHY_107 sky130_fd_sc_hd__decap_3
X_68286_ _82640_/D _68279_/X _68285_/X _83992_/D sky130_fd_sc_hd__a21bo_4
X_65498_ _65397_/A _65397_/B _65498_/C _65498_/Y sky130_fd_sc_hd__nor3_4
XPHY_118 sky130_fd_sc_hd__decap_3
XPHY_129 sky130_fd_sc_hd__decap_3
X_82303_ _82349_/CLK _77217_/B _82303_/Q sky130_fd_sc_hd__dfxtp_4
X_55251_ _55224_/A _55252_/A sky130_fd_sc_hd__buf_2
X_67237_ _67259_/A _87607_/Q _67237_/X sky130_fd_sc_hd__and2_4
X_86071_ _85751_/CLK _51116_/Y _86071_/Q sky130_fd_sc_hd__dfxtp_4
X_52463_ _52431_/A _52468_/A sky130_fd_sc_hd__buf_2
X_64449_ _64515_/A _84861_/Q _64515_/C _64449_/Y sky130_fd_sc_hd__nand3_4
X_83283_ _85826_/CLK _83283_/D _83283_/Q sky130_fd_sc_hd__dfxtp_4
X_80495_ _59159_/Y _66109_/C _80494_/Y _80495_/X sky130_fd_sc_hd__o21a_4
X_54202_ _85485_/Q _54193_/X _54201_/Y _54202_/Y sky130_fd_sc_hd__o21ai_4
X_85022_ _83008_/CLK _57388_/X _85022_/Q sky130_fd_sc_hd__dfxtp_4
X_51414_ _86014_/Q _51402_/X _51413_/Y _51414_/Y sky130_fd_sc_hd__o21ai_4
X_82234_ _82234_/CLK _82266_/Q _77580_/A sky130_fd_sc_hd__dfxtp_4
X_55182_ _55129_/A _55245_/A sky130_fd_sc_hd__buf_2
X_67168_ _67095_/A _87674_/Q _67168_/X sky130_fd_sc_hd__and2_4
X_52394_ _65282_/B _52372_/X _52393_/Y _52394_/Y sky130_fd_sc_hd__o21ai_4
X_54133_ _54131_/Y _54117_/X _54132_/X _85498_/D sky130_fd_sc_hd__a21oi_4
X_66119_ _64710_/A _66119_/B _66119_/X sky130_fd_sc_hd__and2_4
X_51345_ _51350_/A _50832_/B _51345_/Y sky130_fd_sc_hd__nand2_4
X_82165_ _83556_/CLK _84157_/Q _82165_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_809_0_CLK clkbuf_9_404_0_CLK/X _82349_/CLK sky130_fd_sc_hd__clkbuf_1
X_59990_ _59976_/A _62515_/C _62515_/A _59990_/X sky130_fd_sc_hd__o21a_4
X_67099_ _67096_/X _67098_/X _67026_/X _67099_/X sky130_fd_sc_hd__a21o_4
X_81116_ _81084_/CLK _79833_/X _75657_/A sky130_fd_sc_hd__dfxtp_4
X_58941_ _58941_/A _86372_/Q _58941_/Y sky130_fd_sc_hd__nor2_4
X_54064_ _85512_/Q _54018_/X _54063_/Y _54064_/Y sky130_fd_sc_hd__o21ai_4
X_51276_ _51280_/A _49245_/B _51276_/Y sky130_fd_sc_hd__nand2_4
X_86973_ _82906_/CLK _86973_/D _86973_/Q sky130_fd_sc_hd__dfxtp_4
X_82096_ _82860_/CLK _82096_/D _82096_/Q sky130_fd_sc_hd__dfxtp_4
X_53015_ _53019_/A _53036_/B _53019_/C _53015_/D _53015_/X sky130_fd_sc_hd__and4_4
X_50227_ _50227_/A _50227_/X sky130_fd_sc_hd__buf_2
X_85924_ _85444_/CLK _51910_/Y _85924_/Q sky130_fd_sc_hd__dfxtp_4
X_81047_ _80697_/CLK _75390_/X _81047_/Q sky130_fd_sc_hd__dfxtp_4
X_58872_ _58872_/A _86377_/Q _58872_/Y sky130_fd_sc_hd__nor2_4
X_57823_ _57801_/X _57820_/Y _57821_/Y _57822_/X _57809_/X _57823_/X
+ sky130_fd_sc_hd__o32a_4
X_69809_ _73228_/A _69751_/X _69779_/X _69808_/Y _69809_/X sky130_fd_sc_hd__a211o_4
X_50158_ _50153_/A _52367_/B _50158_/Y sky130_fd_sc_hd__nand2_4
X_85855_ _85566_/CLK _85855_/D _85855_/Q sky130_fd_sc_hd__dfxtp_4
X_72820_ _74373_/B _72820_/B _72820_/X sky130_fd_sc_hd__xor2_4
X_84806_ _84807_/CLK _58710_/Y _84806_/Q sky130_fd_sc_hd__dfxtp_4
X_57754_ _57687_/A _57754_/X sky130_fd_sc_hd__buf_2
X_42980_ _42979_/Y _87621_/D sky130_fd_sc_hd__inv_2
X_50089_ _50064_/A _50103_/A sky130_fd_sc_hd__buf_2
X_54966_ _48755_/A _55072_/A sky130_fd_sc_hd__buf_2
X_85786_ _85786_/CLK _52615_/Y _85786_/Q sky130_fd_sc_hd__dfxtp_4
X_82998_ _82998_/CLK _82998_/D _45575_/A sky130_fd_sc_hd__dfxtp_4
X_56705_ _56704_/X _56705_/B _56705_/Y sky130_fd_sc_hd__nand2_4
X_87525_ _87525_/CLK _87525_/D _87525_/Q sky130_fd_sc_hd__dfxtp_4
X_53917_ _53898_/A _53917_/B _53917_/Y sky130_fd_sc_hd__nand2_4
X_41931_ _42059_/A _42013_/A sky130_fd_sc_hd__buf_2
X_72751_ _73352_/A _73535_/A sky130_fd_sc_hd__buf_2
X_84737_ _83402_/CLK _84737_/D _59423_/A sky130_fd_sc_hd__dfxtp_4
X_81949_ _82124_/CLK _78043_/Y _81949_/Q sky130_fd_sc_hd__dfxtp_4
X_57685_ _57677_/X _57682_/Y _57684_/Y _84954_/D sky130_fd_sc_hd__a21oi_4
X_54897_ _54895_/Y _54882_/X _54896_/X _85358_/D sky130_fd_sc_hd__a21oi_4
X_71702_ _71338_/A _71685_/X _71815_/B _71702_/Y sky130_fd_sc_hd__nand3_4
X_59424_ _59423_/Y _59424_/B _59424_/Y sky130_fd_sc_hd__nand2_4
X_44650_ _44650_/A _44650_/X sky130_fd_sc_hd__buf_2
X_56636_ _56567_/Y _56636_/X sky130_fd_sc_hd__buf_2
X_75470_ _75438_/Y _75466_/X _75508_/B _75470_/Y sky130_fd_sc_hd__a21boi_4
X_41862_ _43012_/B _41862_/Y sky130_fd_sc_hd__inv_2
X_87456_ _87210_/CLK _87456_/D _87456_/Q sky130_fd_sc_hd__dfxtp_4
X_53848_ _53848_/A _53848_/B _53848_/Y sky130_fd_sc_hd__nand2_4
X_72682_ _70225_/C _72672_/X _72681_/Y _72682_/X sky130_fd_sc_hd__a21bo_4
X_84668_ _84668_/CLK _84668_/D _60064_/C sky130_fd_sc_hd__dfxtp_4
X_43601_ _43600_/X _43601_/Y sky130_fd_sc_hd__inv_2
X_74421_ _48487_/A _74420_/X _74421_/C _74421_/X sky130_fd_sc_hd__and3_4
X_86407_ _86119_/CLK _86407_/D _65279_/B sky130_fd_sc_hd__dfxtp_4
X_40813_ _40783_/X _82295_/Q _40812_/X _40814_/A sky130_fd_sc_hd__o21a_4
X_59355_ _59292_/X _85636_/Q _59205_/X _59355_/X sky130_fd_sc_hd__o21a_4
X_71633_ _59480_/Y _71628_/X _71632_/Y _71633_/Y sky130_fd_sc_hd__o21ai_4
X_83619_ _85566_/CLK _71065_/Y _83619_/Q sky130_fd_sc_hd__dfxtp_4
X_56567_ _44134_/X _56567_/Y sky130_fd_sc_hd__inv_2
X_44581_ _87046_/Q _44581_/Y sky130_fd_sc_hd__inv_2
X_87387_ _87141_/CLK _43505_/Y _87387_/Q sky130_fd_sc_hd__dfxtp_4
X_53779_ _53777_/Y _53696_/X _53778_/Y _85570_/D sky130_fd_sc_hd__a21boi_4
X_41793_ _41753_/X _41754_/X _41791_/X _88148_/Q _41792_/X _41793_/Y
+ sky130_fd_sc_hd__o32ai_4
X_84599_ _84606_/CLK _84599_/D _79139_/A sky130_fd_sc_hd__dfxtp_4
X_46320_ _46301_/X _82940_/Q _46319_/Y _53969_/A sky130_fd_sc_hd__o21ai_4
X_58306_ _58282_/X _58303_/Y _58305_/Y _58306_/Y sky130_fd_sc_hd__a21oi_4
X_77140_ _77149_/A _81918_/Q _77154_/A sky130_fd_sc_hd__xor2_4
X_55518_ _55509_/X _55515_/X _55517_/X _55536_/A sky130_fd_sc_hd__a21o_4
X_43532_ _53443_/A _43532_/X sky130_fd_sc_hd__buf_2
X_74352_ _83087_/Q _74340_/X _74351_/Y _74352_/X sky130_fd_sc_hd__a21bo_4
XPHY_9 sky130_fd_sc_hd__decap_3
X_86338_ _86340_/CLK _86338_/D _59376_/B sky130_fd_sc_hd__dfxtp_4
X_40744_ _40832_/A _40744_/X sky130_fd_sc_hd__buf_2
X_59286_ _59286_/A _59286_/X sky130_fd_sc_hd__buf_2
X_71564_ _71557_/X _83455_/Q _71563_/Y _71564_/X sky130_fd_sc_hd__a21o_4
X_56498_ _56070_/X _56483_/X _56497_/Y _85173_/D sky130_fd_sc_hd__o21ai_4
X_73303_ _44573_/Y _73006_/X _73302_/Y _73303_/X sky130_fd_sc_hd__a21o_4
X_46251_ _47002_/A _57563_/A sky130_fd_sc_hd__buf_2
XPHY_630 sky130_fd_sc_hd__decap_3
X_70515_ _57659_/Y _70501_/X _70514_/Y _83759_/D sky130_fd_sc_hd__o21ai_4
X_58237_ _84900_/Q _58237_/X sky130_fd_sc_hd__buf_2
X_77071_ _77062_/Y _77069_/Y _77070_/Y _77072_/B sky130_fd_sc_hd__o21a_4
X_43463_ _41643_/X _43446_/X _87409_/Q _43447_/X _87409_/D sky130_fd_sc_hd__a2bb2o_4
X_55449_ _55445_/A _55354_/Y _55445_/C _55449_/Y sky130_fd_sc_hd__a21boi_4
X_74283_ _70134_/C _74003_/B _74282_/X _83114_/D sky130_fd_sc_hd__o21ai_4
X_86269_ _85562_/CLK _86269_/D _86269_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_641 sky130_fd_sc_hd__decap_3
X_40675_ _40736_/A _40710_/B sky130_fd_sc_hd__buf_2
X_71495_ _71487_/X _83479_/Q _71494_/X _83479_/D sky130_fd_sc_hd__a21o_4
XPHY_652 sky130_fd_sc_hd__decap_3
XPHY_663 sky130_fd_sc_hd__decap_3
X_45202_ _45350_/A _45202_/X sky130_fd_sc_hd__buf_2
X_76022_ _76013_/Y _76020_/Y _76021_/Y _76023_/B sky130_fd_sc_hd__o21a_4
X_42414_ _42373_/X _42414_/X sky130_fd_sc_hd__buf_2
X_88008_ _88006_/CLK _42153_/X _88008_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_674 sky130_fd_sc_hd__decap_3
X_73234_ _73062_/X _86191_/Q _73205_/X _73233_/X _73234_/X sky130_fd_sc_hd__a211o_4
X_70446_ _47969_/B _70421_/Y _70445_/Y _70446_/Y sky130_fd_sc_hd__o21ai_4
X_46182_ _44905_/X _46162_/D _57657_/B _46181_/Y _86765_/D sky130_fd_sc_hd__a211o_4
X_58168_ _64272_/A _58160_/B _58168_/Y sky130_fd_sc_hd__nand2_4
XPHY_685 sky130_fd_sc_hd__decap_3
X_43394_ _41461_/X _43386_/X _87443_/Q _43388_/X _87443_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_696 sky130_fd_sc_hd__decap_3
X_45133_ _56233_/C _45073_/X _45132_/X _45133_/Y sky130_fd_sc_hd__o21ai_4
X_57119_ _57109_/X _56634_/X _85077_/Q _57110_/X _85077_/D sky130_fd_sc_hd__a2bb2o_4
X_42345_ _41701_/X _42342_/X _87910_/Q _42343_/X _87910_/D sky130_fd_sc_hd__a2bb2o_4
X_73165_ _73165_/A _73386_/A sky130_fd_sc_hd__buf_2
X_58099_ _58079_/X _58096_/Y _58097_/Y _58098_/X _58083_/X _58099_/X
+ sky130_fd_sc_hd__o32a_4
X_70377_ DATA_TO_HASH[5] _71054_/A sky130_fd_sc_hd__buf_2
Xclkbuf_opt_1_CLK _83246_/CLK _84897_/CLK sky130_fd_sc_hd__clkbuf_16
X_60130_ _60513_/A _61587_/B _79998_/A _60130_/X sky130_fd_sc_hd__or3_4
X_72116_ _59326_/X _72116_/B _72116_/Y sky130_fd_sc_hd__nor2_4
X_49941_ _86295_/Q _49934_/X _49940_/Y _49941_/Y sky130_fd_sc_hd__o21ai_4
X_45064_ _45058_/Y _45062_/Y _45063_/X _45064_/X sky130_fd_sc_hd__a21o_4
X_42276_ _42276_/A _42276_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_62_0_CLK clkbuf_7_63_0_CLK/A clkbuf_7_62_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_73096_ _73239_/A _73096_/B _73096_/X sky130_fd_sc_hd__and2_4
X_77973_ _82077_/Q _77975_/A sky130_fd_sc_hd__inv_2
X_44015_ _45920_/A _68617_/A sky130_fd_sc_hd__buf_2
X_79712_ _84217_/Q _72313_/A _79712_/X sky130_fd_sc_hd__xor2_4
X_41227_ _41227_/A _41227_/Y sky130_fd_sc_hd__inv_2
X_60061_ _59968_/A _59968_/B _59802_/X _60061_/Y sky130_fd_sc_hd__a21oi_4
X_72047_ _83295_/Q _72001_/X _72046_/Y _72047_/Y sky130_fd_sc_hd__o21ai_4
X_76924_ _76924_/A _81471_/D sky130_fd_sc_hd__inv_2
X_49872_ _49893_/A _49884_/B _49862_/C _53084_/D _49872_/X sky130_fd_sc_hd__and4_4
X_48823_ _50069_/A _48823_/B _48823_/X sky130_fd_sc_hd__and2_4
X_79643_ _79619_/A _79642_/D _79642_/B _79643_/X sky130_fd_sc_hd__a21bo_4
X_41158_ _41157_/X _41152_/X _88267_/Q _41153_/X _88267_/D sky130_fd_sc_hd__a2bb2o_4
X_76855_ _76855_/A _81464_/D _81560_/D sky130_fd_sc_hd__xor2_4
X_63820_ _63424_/B _63820_/B _63753_/C _63820_/D _63823_/B sky130_fd_sc_hd__nand4_4
X_75806_ _81100_/Q _75806_/B _80796_/D sky130_fd_sc_hd__xor2_4
X_48754_ _48781_/A _48754_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_77_0_CLK clkbuf_7_77_0_CLK/A clkbuf_7_77_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_79574_ _79573_/B _79572_/Y _79569_/Y _79576_/A sky130_fd_sc_hd__a21o_4
X_45966_ _40330_/Y _45963_/X _66602_/B _45964_/X _45966_/X sky130_fd_sc_hd__a2bb2o_4
X_41089_ _41040_/X _41041_/X _41087_/X _69513_/B _41088_/X _41090_/A
+ sky130_fd_sc_hd__o32ai_4
X_76786_ _76784_/Y _76785_/Y _76786_/X sky130_fd_sc_hd__xor2_4
X_73998_ _72758_/X _66171_/B _73998_/X sky130_fd_sc_hd__and2_4
X_47705_ _54894_/B _53200_/B sky130_fd_sc_hd__buf_2
X_78525_ _78525_/A _78526_/C sky130_fd_sc_hd__inv_2
X_44917_ _44917_/A _44894_/B _44917_/Y sky130_fd_sc_hd__nor2_4
X_75737_ _75715_/A _75714_/Y _75727_/A _75726_/Y _75737_/X sky130_fd_sc_hd__o22a_4
X_63751_ _60928_/X _63751_/X sky130_fd_sc_hd__buf_2
X_48685_ _86500_/Q _48669_/X _48684_/Y _48685_/Y sky130_fd_sc_hd__o21ai_4
X_60963_ _60962_/Y _60963_/X sky130_fd_sc_hd__buf_2
X_72949_ _72877_/A _72949_/X sky130_fd_sc_hd__buf_2
X_45897_ _45896_/X _45897_/X sky130_fd_sc_hd__buf_2
X_62702_ _62678_/A _62727_/B _61796_/X _62702_/Y sky130_fd_sc_hd__nand3_4
X_47636_ _47636_/A _53159_/D sky130_fd_sc_hd__buf_2
X_66470_ _66467_/Y _66449_/X _66469_/X _84117_/D sky130_fd_sc_hd__a21o_4
X_78456_ _78447_/B _82796_/Q _78455_/Y _78465_/A sky130_fd_sc_hd__a21boi_4
X_44848_ _43927_/X _44848_/X sky130_fd_sc_hd__buf_2
X_63682_ _63655_/A _58296_/A _63672_/C _60682_/A _63682_/X sky130_fd_sc_hd__and4_4
X_75668_ _80909_/Q _75670_/A sky130_fd_sc_hd__inv_2
X_60894_ _60865_/C _64180_/C _60894_/X sky130_fd_sc_hd__and2_4
X_65421_ _65268_/A _65294_/B _65421_/C _65421_/X sky130_fd_sc_hd__and3_4
X_77407_ _77394_/A _77405_/Y _77406_/Y _77416_/A sky130_fd_sc_hd__o21a_4
Xclkbuf_8_140_0_CLK clkbuf_7_70_0_CLK/X clkbuf_9_281_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_62633_ _61694_/B _62309_/B _62309_/C _62225_/X _62633_/Y sky130_fd_sc_hd__nand4_4
X_74619_ _58253_/A _74613_/X _56159_/A _74614_/X _74619_/X sky130_fd_sc_hd__a211o_4
X_47567_ _47567_/A _53125_/D sky130_fd_sc_hd__buf_2
X_78387_ _82792_/Q _78387_/Y sky130_fd_sc_hd__inv_2
X_44779_ _41370_/Y _44774_/X _86959_/Q _44775_/X _86959_/D sky130_fd_sc_hd__a2bb2o_4
X_75599_ _81109_/Q _75599_/B _75891_/A sky130_fd_sc_hd__xnor2_4
X_49306_ _49302_/A _50827_/B _49306_/Y sky130_fd_sc_hd__nand2_4
X_68140_ _68120_/A _68140_/X sky130_fd_sc_hd__buf_2
X_46518_ _46513_/Y _46399_/X _46517_/Y _86730_/D sky130_fd_sc_hd__a21boi_4
X_65352_ _65401_/A _85828_/Q _65352_/X sky130_fd_sc_hd__and2_4
X_77338_ _77338_/A _77338_/B _77339_/B sky130_fd_sc_hd__xor2_4
X_62564_ _62562_/Y _62540_/X _62563_/Y _84401_/D sky130_fd_sc_hd__a21oi_4
X_47498_ _54772_/B _53080_/B sky130_fd_sc_hd__buf_2
X_64303_ _64303_/A _64303_/X sky130_fd_sc_hd__buf_2
X_49237_ _49241_/A _50757_/B _49237_/Y sky130_fd_sc_hd__nand2_4
X_61515_ _61514_/Y _61515_/Y sky130_fd_sc_hd__inv_2
X_68071_ _68044_/A _68071_/B _68071_/X sky130_fd_sc_hd__and2_4
X_46449_ _46449_/A _50812_/A sky130_fd_sc_hd__buf_2
X_65283_ _65172_/X _86151_/Q _65256_/X _65282_/X _65283_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_7_15_0_CLK clkbuf_6_7_0_CLK/X clkbuf_8_31_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_77269_ _77268_/X _77269_/Y sky130_fd_sc_hd__inv_2
X_62495_ _62570_/A _62027_/X _62479_/C _62463_/X _62495_/X sky130_fd_sc_hd__and4_4
Xclkbuf_8_155_0_CLK clkbuf_7_77_0_CLK/X clkbuf_9_311_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_67022_ _67144_/A _67023_/A sky130_fd_sc_hd__buf_2
X_79008_ _78997_/A _78997_/B _79007_/X _79008_/Y sky130_fd_sc_hd__a21oi_4
X_64234_ _64234_/A _64234_/B _58225_/A _64221_/X _64234_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_150_0_CLK clkbuf_9_75_0_CLK/X _81632_/CLK sky130_fd_sc_hd__clkbuf_1
X_61446_ _61444_/X _61394_/X _61445_/Y _61446_/Y sky130_fd_sc_hd__a21oi_4
X_49168_ _49156_/X _50708_/B _49168_/Y sky130_fd_sc_hd__nand2_4
X_80280_ _80275_/Y _80280_/B _80280_/C _80280_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_780_0_CLK clkbuf_9_390_0_CLK/X _82580_/CLK sky130_fd_sc_hd__clkbuf_1
X_48119_ _48075_/X _82918_/Q _48118_/X _48329_/A sky130_fd_sc_hd__o21ai_4
X_64165_ _64163_/X _64129_/X _64164_/Y _64165_/Y sky130_fd_sc_hd__a21oi_4
X_49099_ _49099_/A _52370_/A sky130_fd_sc_hd__buf_2
X_61377_ _61377_/A _61376_/X _61377_/C _61377_/Y sky130_fd_sc_hd__nand3_4
X_51130_ _51130_/A _51130_/B _51130_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_271_0_CLK clkbuf_9_271_0_CLK/A clkbuf_9_271_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_63116_ _79414_/A _63072_/X _63115_/Y _84352_/D sky130_fd_sc_hd__a21o_4
X_60328_ _60235_/A _60327_/X _60198_/A _79691_/A _59814_/X _60328_/X
+ sky130_fd_sc_hd__o32a_4
X_68973_ _68907_/X _68882_/X _68964_/Y _68972_/Y _68973_/X sky130_fd_sc_hd__a211o_4
X_64096_ _61593_/B _64161_/B _64150_/C _64161_/D _64096_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_10_165_0_CLK clkbuf_9_82_0_CLK/X _81288_/CLK sky130_fd_sc_hd__clkbuf_1
X_51061_ _51056_/A _51045_/B _51071_/C _52750_/D _51061_/X sky130_fd_sc_hd__and4_4
X_67924_ _68461_/A _68120_/A sky130_fd_sc_hd__buf_2
X_63047_ _58418_/A _63010_/X _60523_/X _59463_/Y _60412_/X _63047_/Y
+ sky130_fd_sc_hd__o32ai_4
X_60259_ _60259_/A _60259_/B _60259_/Y sky130_fd_sc_hd__nand2_4
X_83970_ _80931_/CLK _83970_/D _80826_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_795_0_CLK clkbuf_9_397_0_CLK/X _82671_/CLK sky130_fd_sc_hd__clkbuf_1
X_50012_ _48169_/X _50012_/X sky130_fd_sc_hd__buf_2
X_82921_ _82923_/CLK _78182_/X _46528_/A sky130_fd_sc_hd__dfxtp_4
X_67855_ _66554_/X _67955_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_286_0_CLK clkbuf_9_286_0_CLK/A clkbuf_9_286_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_54820_ _54900_/A _54843_/B sky130_fd_sc_hd__buf_2
X_66806_ _84096_/Q _66734_/X _66805_/X _66806_/X sky130_fd_sc_hd__a21bo_4
X_85640_ _85643_/CLK _85640_/D _85640_/Q sky130_fd_sc_hd__dfxtp_4
X_82852_ _82596_/CLK _78088_/B _82852_/Q sky130_fd_sc_hd__dfxtp_4
X_67786_ _87392_/Q _67717_/X _67718_/X _67785_/X _67786_/X sky130_fd_sc_hd__a211o_4
X_64998_ _64995_/Y _64939_/X _64997_/Y _84219_/D sky130_fd_sc_hd__a21o_4
X_81803_ _81632_/CLK _81803_/D _81803_/Q sky130_fd_sc_hd__dfxtp_4
X_69525_ _69522_/X _69524_/X _69385_/X _69525_/X sky130_fd_sc_hd__a21o_4
X_54751_ _85384_/Q _54729_/X _54750_/Y _54751_/Y sky130_fd_sc_hd__o21ai_4
X_66737_ _87884_/Q _66639_/X _66688_/X _66736_/X _66737_/X sky130_fd_sc_hd__a211o_4
X_85571_ _85571_/CLK _53775_/Y _85571_/Q sky130_fd_sc_hd__dfxtp_4
X_51963_ _65972_/B _51960_/X _51962_/Y _51963_/Y sky130_fd_sc_hd__o21ai_4
X_63949_ _63520_/B _63934_/X _63949_/C _64027_/D _63949_/Y sky130_fd_sc_hd__nand4_4
X_82783_ _82975_/CLK _78762_/X _82783_/Q sky130_fd_sc_hd__dfxtp_4
X_87310_ _83158_/CLK _87310_/D _87310_/Q sky130_fd_sc_hd__dfxtp_4
X_53702_ _53763_/A _53734_/C sky130_fd_sc_hd__buf_2
X_84522_ _84292_/CLK _61065_/X _84522_/Q sky130_fd_sc_hd__dfxtp_4
X_50914_ _50908_/A _50919_/B _50897_/X _51777_/D _50914_/X sky130_fd_sc_hd__and4_4
X_57470_ _56885_/A _57470_/B _56884_/Y _57470_/Y sky130_fd_sc_hd__nand3_4
X_81734_ _82067_/CLK _81734_/D _81734_/Q sky130_fd_sc_hd__dfxtp_4
X_69456_ _69453_/X _69455_/X _69399_/X _69461_/A sky130_fd_sc_hd__a21o_4
X_88290_ _87022_/CLK _88290_/D _69376_/B sky130_fd_sc_hd__dfxtp_4
X_54682_ _54682_/A _47334_/Y _54682_/Y sky130_fd_sc_hd__nand2_4
X_66668_ _66663_/X _66666_/X _66667_/X _66668_/X sky130_fd_sc_hd__a21o_4
X_51894_ _51890_/Y _51877_/X _51893_/X _85927_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_8_108_0_CLK clkbuf_7_54_0_CLK/X clkbuf_9_217_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_56421_ _56099_/X _56409_/X _56420_/Y _85200_/D sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_103_0_CLK clkbuf_9_51_0_CLK/X _84529_/CLK sky130_fd_sc_hd__clkbuf_1
X_68407_ _68404_/X _68406_/X _68033_/X _68407_/X sky130_fd_sc_hd__a21o_4
X_87241_ _88012_/CLK _87241_/D _68627_/B sky130_fd_sc_hd__dfxtp_4
X_53633_ _53656_/A _48391_/A _53633_/Y sky130_fd_sc_hd__nand2_4
X_65619_ _65608_/Y _65619_/B _65619_/Y sky130_fd_sc_hd__nand2_4
X_84453_ _84454_/CLK _61803_/Y _78076_/B sky130_fd_sc_hd__dfxtp_4
X_50845_ _50845_/A _49322_/B _50845_/Y sky130_fd_sc_hd__nand2_4
X_81665_ _81682_/CLK _81697_/Q _76635_/A sky130_fd_sc_hd__dfxtp_4
X_69387_ _69612_/A _88289_/Q _69387_/X sky130_fd_sc_hd__and2_4
X_66599_ _87890_/Q _66562_/X _66564_/X _66598_/X _66599_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_733_0_CLK clkbuf_9_366_0_CLK/X _87333_/CLK sky130_fd_sc_hd__clkbuf_1
X_59140_ _59053_/A _59140_/X sky130_fd_sc_hd__buf_2
X_83404_ _83372_/CLK _83404_/D _58298_/A sky130_fd_sc_hd__dfxtp_4
X_80616_ _80623_/A _80615_/Y _80622_/B sky130_fd_sc_hd__xor2_4
X_56352_ _56358_/A _56358_/B _55764_/B _56352_/Y sky130_fd_sc_hd__nand3_4
X_68338_ _68338_/A _68338_/X sky130_fd_sc_hd__buf_2
X_87172_ _87174_/CLK _44295_/Y _44293_/B sky130_fd_sc_hd__dfxtp_4
X_53564_ _85612_/Q _53540_/X _53563_/Y _53564_/Y sky130_fd_sc_hd__o21ai_4
X_84384_ _84518_/CLK _62767_/Y _62766_/C sky130_fd_sc_hd__dfxtp_4
X_50776_ _50505_/A _50777_/A sky130_fd_sc_hd__buf_2
X_81596_ _81433_/CLK _84196_/Q _81596_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_224_0_CLK clkbuf_8_112_0_CLK/X clkbuf_9_224_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_55303_ _55317_/A _57419_/A _55303_/X sky130_fd_sc_hd__and2_4
X_86123_ _86029_/CLK _86123_/D _86123_/Q sky130_fd_sc_hd__dfxtp_4
X_52515_ _52515_/A _52515_/X sky130_fd_sc_hd__buf_2
X_59071_ _59048_/X _85659_/Q _59070_/X _59071_/X sky130_fd_sc_hd__o21a_4
X_83335_ _83335_/CLK _71901_/Y _83335_/Q sky130_fd_sc_hd__dfxtp_4
X_56283_ _56282_/Y _56350_/A sky130_fd_sc_hd__buf_2
X_80547_ _84770_/Q _84162_/Q _80547_/X sky130_fd_sc_hd__xor2_4
X_68269_ _67656_/X _67660_/X _68260_/X _68269_/Y sky130_fd_sc_hd__a21oi_4
X_53495_ _53478_/A _73765_/A _53495_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_118_0_CLK clkbuf_9_59_0_CLK/X _84392_/CLK sky130_fd_sc_hd__clkbuf_1
X_58022_ _57939_/X _85996_/Q _58021_/X _58022_/Y sky130_fd_sc_hd__o21ai_4
X_70300_ _70289_/X _74783_/A _70299_/X _70300_/X sky130_fd_sc_hd__a21o_4
X_55234_ _55129_/A _55235_/A sky130_fd_sc_hd__buf_2
X_86054_ _86054_/CLK _51208_/Y _86054_/Q sky130_fd_sc_hd__dfxtp_4
X_40460_ _40437_/X _40443_/X _40459_/X _88388_/Q _40447_/X _40461_/A
+ sky130_fd_sc_hd__o32ai_4
X_52446_ _51256_/A _52446_/B _52369_/X _52446_/X sky130_fd_sc_hd__and3_4
X_83266_ _86289_/CLK _72312_/Y _83266_/Q sky130_fd_sc_hd__dfxtp_4
X_71280_ _53205_/B _71265_/X _71279_/Y _71280_/Y sky130_fd_sc_hd__o21ai_4
X_80478_ _80478_/A _80478_/B _80478_/X sky130_fd_sc_hd__or2_4
Xclkbuf_10_748_0_CLK clkbuf_9_374_0_CLK/X _88001_/CLK sky130_fd_sc_hd__clkbuf_1
X_85005_ _85005_/CLK _57434_/Y _57430_/A sky130_fd_sc_hd__dfxtp_4
X_70231_ _70231_/A _70239_/A sky130_fd_sc_hd__buf_2
X_82217_ _83905_/CLK _82249_/Q _82217_/Q sky130_fd_sc_hd__dfxtp_4
X_55165_ _55134_/X _55165_/X sky130_fd_sc_hd__buf_2
X_40391_ _40390_/Y _40391_/X sky130_fd_sc_hd__buf_2
X_52377_ _50677_/A _52446_/B _52369_/X _52377_/X sky130_fd_sc_hd__and3_4
X_83197_ _85013_/CLK _83197_/D _83197_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_239_0_CLK clkbuf_9_239_0_CLK/A clkbuf_9_239_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_42130_ _41108_/X _42125_/X _88020_/Q _42126_/X _88020_/D sky130_fd_sc_hd__a2bb2o_4
X_54116_ _85501_/Q _54113_/X _54115_/Y _54116_/Y sky130_fd_sc_hd__o21ai_4
X_51328_ _51310_/X _51328_/B _51328_/Y sky130_fd_sc_hd__nand2_4
X_70162_ _70348_/B _70162_/X sky130_fd_sc_hd__buf_2
X_82148_ _84231_/CLK _84140_/Q _82148_/Q sky130_fd_sc_hd__dfxtp_4
X_55096_ _55112_/A _55104_/B _55083_/C _47776_/A _55096_/X sky130_fd_sc_hd__and4_4
X_59973_ _59973_/A _59977_/B sky130_fd_sc_hd__buf_2
X_42061_ _88053_/Q _42061_/Y sky130_fd_sc_hd__inv_2
X_58924_ _58918_/X _58920_/Y _58921_/Y _58874_/X _58923_/X _58924_/X
+ sky130_fd_sc_hd__o32a_4
X_54047_ _54047_/A _54043_/B _51749_/X _54047_/X sky130_fd_sc_hd__and3_4
X_51259_ _51259_/A _51259_/X sky130_fd_sc_hd__buf_2
X_74970_ _81140_/D _74989_/C _74987_/A sky130_fd_sc_hd__xor2_4
X_70093_ _70011_/X _69094_/Y _70081_/X _70092_/Y _70093_/X sky130_fd_sc_hd__a211o_4
X_86956_ _88224_/CLK _86956_/D _86956_/Q sky130_fd_sc_hd__dfxtp_4
X_82079_ _81169_/CLK _82079_/D _82079_/Q sky130_fd_sc_hd__dfxtp_4
X_41012_ _40321_/A _41013_/A sky130_fd_sc_hd__buf_2
X_73921_ _73921_/A _56181_/X _73921_/Y sky130_fd_sc_hd__nor2_4
X_85907_ _86549_/CLK _85907_/D _73901_/B sky130_fd_sc_hd__dfxtp_4
X_58855_ _58843_/Y _58739_/X _58850_/X _58854_/X _84795_/D sky130_fd_sc_hd__a22oi_4
X_86887_ _86887_/CLK _45280_/Y _62557_/A sky130_fd_sc_hd__dfxtp_4
X_57806_ _58080_/A _57806_/X sky130_fd_sc_hd__buf_2
X_45820_ _63314_/B _61655_/A sky130_fd_sc_hd__buf_2
X_76640_ _76640_/A _76640_/B _76637_/X _76640_/Y sky130_fd_sc_hd__nand3_4
X_73852_ _73949_/A _66082_/B _73852_/X sky130_fd_sc_hd__and2_4
X_85838_ _85536_/CLK _85838_/D _65094_/B sky130_fd_sc_hd__dfxtp_4
X_58786_ _64836_/A _59061_/A sky130_fd_sc_hd__buf_2
X_55998_ _55891_/X _74312_/C sky130_fd_sc_hd__buf_2
X_72803_ _72732_/B _72803_/X sky130_fd_sc_hd__buf_2
X_45751_ _45742_/X _45747_/Y _45750_/Y _45751_/Y sky130_fd_sc_hd__a21oi_4
X_57737_ _57705_/X _85503_/Q _57736_/X _57737_/X sky130_fd_sc_hd__o21a_4
X_76571_ _76568_/Y _76571_/B _81341_/D sky130_fd_sc_hd__nor2_4
X_42963_ _42951_/A _42963_/X sky130_fd_sc_hd__buf_2
X_54949_ _85347_/Q _53449_/X _54948_/Y _54949_/Y sky130_fd_sc_hd__o21ai_4
X_73783_ _73711_/A _66037_/B _73783_/X sky130_fd_sc_hd__and2_4
X_85769_ _85770_/CLK _52710_/Y _85769_/Q sky130_fd_sc_hd__dfxtp_4
X_70995_ _70990_/A _71080_/B _70990_/C _70995_/Y sky130_fd_sc_hd__nand3_4
X_78310_ _78309_/Y _78310_/Y sky130_fd_sc_hd__inv_2
X_44702_ _44702_/A _44702_/Y sky130_fd_sc_hd__inv_2
X_75522_ _75522_/A _75524_/B sky130_fd_sc_hd__inv_2
X_87508_ _87253_/CLK _43268_/X _87508_/Q sky130_fd_sc_hd__dfxtp_4
X_41914_ _41914_/A _41914_/Y sky130_fd_sc_hd__inv_2
X_48470_ _65584_/B _48419_/X _48469_/Y _48470_/Y sky130_fd_sc_hd__o21ai_4
X_72734_ _44131_/A _73262_/A sky130_fd_sc_hd__buf_2
X_79290_ _79286_/X _79304_/B _79291_/A sky130_fd_sc_hd__xor2_4
X_57668_ _57668_/A _57668_/Y sky130_fd_sc_hd__inv_2
X_45682_ _74667_/B _45654_/B _45682_/Y sky130_fd_sc_hd__nand2_4
X_42894_ _41651_/X _42886_/X _87663_/Q _42887_/X _87663_/D sky130_fd_sc_hd__a2bb2o_4
X_47421_ _47420_/Y _53041_/B sky130_fd_sc_hd__buf_2
X_59407_ _59407_/A _59399_/B _59407_/Y sky130_fd_sc_hd__nand2_4
X_78241_ _78241_/A _78241_/B _78241_/X sky130_fd_sc_hd__or2_4
X_44633_ _44633_/A _44633_/Y sky130_fd_sc_hd__inv_2
X_56619_ _56619_/A _56619_/X sky130_fd_sc_hd__buf_2
X_75453_ _81084_/Q _75457_/A sky130_fd_sc_hd__inv_2
X_87439_ _87484_/CLK _43402_/X _87439_/Q sky130_fd_sc_hd__dfxtp_4
X_41845_ _41839_/X _41841_/X _40501_/X _88125_/Q _41835_/X _41846_/A
+ sky130_fd_sc_hd__o32ai_4
X_72665_ _70205_/C _72658_/X _72664_/Y _83198_/D sky130_fd_sc_hd__a21bo_4
X_57599_ _57564_/X _53567_/B _57599_/Y sky130_fd_sc_hd__nand2_4
X_74404_ _83073_/Q _74377_/X _74403_/Y _74404_/Y sky130_fd_sc_hd__o21ai_4
X_47352_ _47352_/A _52999_/B sky130_fd_sc_hd__buf_2
X_59338_ _84750_/Q _59268_/X _59330_/X _59337_/X _59338_/Y sky130_fd_sc_hd__a2bb2oi_4
X_71616_ _70558_/X _70667_/A _71614_/C _71606_/X _71616_/Y sky130_fd_sc_hd__nor4_4
X_78172_ _78172_/A _78171_/Y _78173_/B sky130_fd_sc_hd__xnor2_4
X_44564_ _44564_/A _44564_/Y sky130_fd_sc_hd__inv_2
X_75384_ _75383_/B _75383_/C _75383_/A _75384_/X sky130_fd_sc_hd__o21a_4
X_41776_ _82885_/Q _46240_/A _41776_/X sky130_fd_sc_hd__or2_4
X_72596_ _79321_/B _60349_/X _72595_/X _72596_/X sky130_fd_sc_hd__o21a_4
X_46303_ _40842_/X _48924_/A _46303_/Y sky130_fd_sc_hd__nand2_4
X_77123_ _82099_/Q _77123_/B _77123_/X sky130_fd_sc_hd__xor2_4
X_43515_ _41782_/X _43513_/X _87382_/Q _43514_/X _87382_/D sky130_fd_sc_hd__a2bb2o_4
X_74335_ _70321_/C _74327_/X _74334_/Y _74335_/X sky130_fd_sc_hd__a21bo_4
X_40727_ _40727_/A _40710_/B _40727_/X sky130_fd_sc_hd__or2_4
X_59269_ _59256_/A _86347_/Q _59269_/Y sky130_fd_sc_hd__nor2_4
X_47283_ _47283_/A _52963_/D sky130_fd_sc_hd__buf_2
X_71547_ _71531_/X _83461_/Q _71546_/Y _83461_/D sky130_fd_sc_hd__a21o_4
X_44495_ _44495_/A _87080_/D sky130_fd_sc_hd__inv_2
X_61300_ _61355_/A _61305_/A sky130_fd_sc_hd__buf_2
X_49022_ _49022_/A _72025_/B _49022_/X sky130_fd_sc_hd__and2_4
X_46234_ _46233_/Y _46234_/Y sky130_fd_sc_hd__inv_2
XPHY_460 sky130_fd_sc_hd__decap_3
X_77054_ _77054_/A _82281_/D _77055_/B sky130_fd_sc_hd__nor2_4
X_43446_ _43513_/A _43446_/X sky130_fd_sc_hd__buf_2
X_62280_ _62597_/B _61796_/X _62237_/X _62280_/D _62280_/X sky130_fd_sc_hd__and4_4
X_74266_ _74266_/A _72853_/X _74266_/Y sky130_fd_sc_hd__nor2_4
XPHY_471 sky130_fd_sc_hd__decap_3
X_40658_ _40657_/Y _40658_/Y sky130_fd_sc_hd__inv_2
X_71478_ _71429_/A _71716_/D sky130_fd_sc_hd__buf_2
XPHY_482 sky130_fd_sc_hd__decap_3
XPHY_493 sky130_fd_sc_hd__decap_3
X_76005_ _76005_/A _76005_/B _76005_/C _76006_/B sky130_fd_sc_hd__and3_4
X_61231_ _61196_/A _64223_/A sky130_fd_sc_hd__buf_2
X_73217_ _73217_/A _73216_/X _73217_/Y sky130_fd_sc_hd__nand2_4
X_46165_ _46166_/A _46170_/C _46169_/C _46167_/B sky130_fd_sc_hd__a21boi_4
X_70429_ _71145_/A _71196_/A sky130_fd_sc_hd__buf_2
X_43377_ _43376_/Y _43377_/Y sky130_fd_sc_hd__inv_2
X_74197_ _74237_/A _66301_/B _74197_/X sky130_fd_sc_hd__and2_4
X_40589_ _40585_/X _82878_/Q _40588_/X _40590_/A sky130_fd_sc_hd__o21ai_4
X_45116_ _45265_/A _45116_/X sky130_fd_sc_hd__buf_2
X_42328_ _41651_/X _42325_/X _87919_/Q _42326_/X _87919_/D sky130_fd_sc_hd__a2bb2o_4
X_61162_ _61107_/X _61254_/C _61131_/Y _61162_/X sky130_fd_sc_hd__o21a_4
X_73148_ _42020_/Y _72888_/X _72890_/X _73147_/Y _73148_/X sky130_fd_sc_hd__a211o_4
X_46096_ _46162_/A _46090_/Y _46091_/Y _46096_/D _46097_/A sky130_fd_sc_hd__and4_4
X_60113_ _60058_/B _59913_/X _60027_/X _60110_/X _64638_/B _60113_/Y
+ sky130_fd_sc_hd__a32oi_4
X_49924_ _49924_/A _49924_/X sky130_fd_sc_hd__buf_2
X_45047_ _44968_/X _45067_/B sky130_fd_sc_hd__buf_2
X_42259_ _42259_/A _42259_/X sky130_fd_sc_hd__buf_2
X_65970_ _65970_/A _65970_/B _65970_/C _65970_/X sky130_fd_sc_hd__and3_4
X_61093_ _64243_/A _61107_/A sky130_fd_sc_hd__inv_2
X_73079_ _73193_/A _73079_/X sky130_fd_sc_hd__buf_2
X_77956_ _77961_/B _77944_/B _77955_/X _77956_/Y sky130_fd_sc_hd__a21oi_4
X_64921_ _64846_/X _85525_/Q _64919_/X _64920_/X _64921_/X sky130_fd_sc_hd__a211o_4
X_60044_ _60044_/A _60044_/Y sky130_fd_sc_hd__inv_2
X_76907_ _76907_/A _76907_/B _76934_/A sky130_fd_sc_hd__xnor2_4
X_49855_ _49864_/A _53067_/B _49855_/Y sky130_fd_sc_hd__nand2_4
X_77887_ _77887_/A _77886_/Y _77888_/B sky130_fd_sc_hd__xnor2_4
X_48806_ _48804_/Y _48785_/X _48805_/X _86479_/D sky130_fd_sc_hd__a21oi_4
X_67640_ _84061_/Q _67568_/X _67639_/X _84061_/D sky130_fd_sc_hd__a21bo_4
X_79626_ _79614_/X _79615_/X _79625_/Y _79626_/Y sky130_fd_sc_hd__a21boi_4
X_64852_ _64845_/X _64849_/X _64851_/X _64855_/A sky130_fd_sc_hd__a21o_4
Xclkbuf_4_12_0_CLK clkbuf_3_6_1_CLK/X clkbuf_4_12_1_CLK/A sky130_fd_sc_hd__clkbuf_1
X_76838_ _81590_/Q _76838_/B _81558_/D sky130_fd_sc_hd__xor2_4
X_49786_ _86323_/Q _49768_/X _49785_/Y _49786_/Y sky130_fd_sc_hd__o21ai_4
X_46998_ _82393_/Q _46999_/A sky130_fd_sc_hd__inv_2
X_63803_ _61378_/A _63772_/B _63803_/C _63787_/D _63809_/A sky130_fd_sc_hd__nand4_4
X_48737_ _48737_/A _52121_/B _48737_/Y sky130_fd_sc_hd__nand2_4
X_67571_ _87913_/Q _67473_/X _67524_/X _67570_/X _67571_/X sky130_fd_sc_hd__a211o_4
X_79557_ _79557_/A _79549_/Y _79550_/Y _79558_/B sky130_fd_sc_hd__nand3_4
X_45949_ _45918_/Y _45950_/B sky130_fd_sc_hd__inv_2
X_64783_ _64608_/A _64867_/B sky130_fd_sc_hd__buf_2
X_76769_ _76762_/Y _76763_/A _76768_/Y _76769_/Y sky130_fd_sc_hd__a21oi_4
X_61995_ _59692_/Y _61995_/X sky130_fd_sc_hd__buf_2
X_69310_ _87027_/Q _69153_/X _69168_/X _69309_/X _69310_/X sky130_fd_sc_hd__a211o_4
X_66522_ _60371_/X _66355_/Y _66521_/Y _66522_/Y sky130_fd_sc_hd__o21ai_4
X_78508_ _78508_/A _78508_/Y sky130_fd_sc_hd__inv_2
X_63734_ _63734_/A _63733_/X _63735_/A sky130_fd_sc_hd__nand2_4
X_60946_ _72543_/A _60946_/X sky130_fd_sc_hd__buf_2
X_48668_ _48662_/Y _48651_/X _48667_/X _48668_/Y sky130_fd_sc_hd__a21oi_4
X_79488_ _79442_/Y _79482_/X _79487_/Y _79488_/Y sky130_fd_sc_hd__a21oi_4
X_69241_ _87032_/Q _69239_/X _69103_/X _69240_/X _69241_/X sky130_fd_sc_hd__a211o_4
X_47619_ _47619_/A _47619_/X sky130_fd_sc_hd__buf_2
X_66453_ _66453_/A _65833_/B _66160_/X _66453_/Y sky130_fd_sc_hd__nand3_4
X_78439_ _78438_/Y _78439_/B _78439_/C _78439_/Y sky130_fd_sc_hd__nand3_4
X_63665_ _59430_/Y _63648_/B _63665_/Y sky130_fd_sc_hd__nor2_4
X_48599_ _48823_/B _50503_/B sky130_fd_sc_hd__buf_2
X_60877_ _60857_/X _60879_/B sky130_fd_sc_hd__buf_2
X_65404_ _65272_/X _85538_/Q _65326_/X _65403_/X _65404_/X sky130_fd_sc_hd__a211o_4
X_50630_ _50624_/A _72025_/B _50630_/Y sky130_fd_sc_hd__nand2_4
X_62616_ _62653_/A _62653_/B _62616_/C _62616_/Y sky130_fd_sc_hd__nor3_4
X_81450_ _81344_/CLK _81450_/D _81418_/D sky130_fd_sc_hd__dfxtp_4
X_69172_ _69167_/X _69170_/X _69171_/X _69172_/Y sky130_fd_sc_hd__a21oi_4
X_66384_ _84133_/Q _65296_/X _66383_/Y _84133_/D sky130_fd_sc_hd__a21o_4
X_63596_ _58385_/Y _63558_/X _61561_/A _63559_/X _63596_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_10_1005_0_CLK clkbuf_9_502_0_CLK/X _83068_/CLK sky130_fd_sc_hd__clkbuf_1
X_80401_ _80401_/A _80400_/X _80416_/B sky130_fd_sc_hd__xnor2_4
X_68123_ _68121_/X _66771_/Y _68110_/X _68122_/Y _68123_/X sky130_fd_sc_hd__a211o_4
X_65335_ _65258_/A _65335_/B _65335_/X sky130_fd_sc_hd__and2_4
X_50561_ _48885_/A _50560_/X _50552_/C _50561_/X sky130_fd_sc_hd__and3_4
X_81381_ _84087_/CLK _81381_/D _76821_/B sky130_fd_sc_hd__dfxtp_4
X_62547_ _62237_/X _62548_/C sky130_fd_sc_hd__buf_2
X_52300_ _85850_/Q _52297_/X _52299_/Y _52300_/Y sky130_fd_sc_hd__o21ai_4
X_83120_ _86213_/CLK _83120_/D _83120_/Q sky130_fd_sc_hd__dfxtp_4
X_80332_ _80314_/Y _80332_/Y sky130_fd_sc_hd__inv_2
X_68054_ _68405_/A _68054_/B _68054_/X sky130_fd_sc_hd__and2_4
X_53280_ _53276_/A _54460_/B _53280_/Y sky130_fd_sc_hd__nand2_4
X_65266_ _65262_/X _65111_/B _65265_/X _65266_/Y sky130_fd_sc_hd__nand3_4
X_50492_ _52199_/A _50492_/B _50497_/C _50492_/X sky130_fd_sc_hd__and3_4
X_62478_ _62478_/A _62478_/X sky130_fd_sc_hd__buf_2
X_67005_ _67001_/X _67004_/X _67005_/Y sky130_fd_sc_hd__nand2_4
X_52231_ _85863_/Q _52214_/X _52230_/Y _52231_/Y sky130_fd_sc_hd__o21ai_4
X_64217_ _64440_/A _64315_/A sky130_fd_sc_hd__buf_2
X_83051_ _83310_/CLK _74510_/Y _83051_/Q sky130_fd_sc_hd__dfxtp_4
X_61429_ _61429_/A _61428_/X _61429_/C _61429_/Y sky130_fd_sc_hd__nand3_4
X_80263_ _79900_/X _80263_/B _80264_/B sky130_fd_sc_hd__nand2_4
X_65197_ _65193_/Y _65195_/X _65196_/X _84211_/D sky130_fd_sc_hd__a21o_4
X_82002_ _82005_/CLK _82034_/Q _77111_/A sky130_fd_sc_hd__dfxtp_4
X_52162_ _52159_/Y _52145_/X _52161_/X _85877_/D sky130_fd_sc_hd__a21oi_4
X_64148_ _60982_/A _64182_/B sky130_fd_sc_hd__buf_2
X_80194_ _84948_/Q _84196_/Q _80196_/A sky130_fd_sc_hd__xor2_4
X_51113_ _86071_/Q _51101_/X _51112_/Y _51113_/Y sky130_fd_sc_hd__o21ai_4
X_86810_ _86814_/CLK _46021_/Y _86810_/Q sky130_fd_sc_hd__dfxtp_4
X_52093_ _52093_/A _52098_/B _52033_/X _52093_/X sky130_fd_sc_hd__and3_4
X_56970_ _56877_/X _56922_/X _56893_/B _56971_/C sky130_fd_sc_hd__o21ai_4
X_64079_ _58268_/A _60866_/A _64078_/X _64079_/Y sky130_fd_sc_hd__o21ai_4
X_68956_ _68669_/A _68956_/B _68956_/Y sky130_fd_sc_hd__nor2_4
X_87790_ _87790_/CLK _87790_/D _69203_/B sky130_fd_sc_hd__dfxtp_4
X_51044_ _86084_/Q _51020_/X _51043_/Y _51044_/Y sky130_fd_sc_hd__o21ai_4
X_55921_ _55903_/A _85178_/Q _55921_/X sky130_fd_sc_hd__and2_4
X_67907_ _64706_/A _69797_/A sky130_fd_sc_hd__buf_2
X_86741_ _85527_/CLK _46393_/Y _86741_/Q sky130_fd_sc_hd__dfxtp_4
X_83953_ _83957_/CLK _83953_/D _80809_/D sky130_fd_sc_hd__dfxtp_4
X_68887_ _74051_/A _68883_/X _68884_/X _68886_/Y _68887_/X sky130_fd_sc_hd__a211o_4
X_58640_ _64656_/A _58641_/A sky130_fd_sc_hd__buf_2
X_82904_ _87922_/CLK _78240_/B _41679_/A sky130_fd_sc_hd__dfxtp_4
X_55852_ _83026_/Q _55507_/X _44097_/X _55851_/X _55853_/B sky130_fd_sc_hd__a211o_4
X_67838_ _67833_/X _67837_/X _67742_/X _67842_/A sky130_fd_sc_hd__a21o_4
X_86672_ _86353_/CLK _86672_/D _86672_/Q sky130_fd_sc_hd__dfxtp_4
X_83884_ _82301_/CLK _83884_/D _81956_/D sky130_fd_sc_hd__dfxtp_4
X_54803_ _54798_/A _54816_/B _54798_/C _53113_/D _54803_/X sky130_fd_sc_hd__and4_4
X_85623_ _86235_/CLK _53513_/Y _85623_/Q sky130_fd_sc_hd__dfxtp_4
X_58571_ _58813_/A _58571_/X sky130_fd_sc_hd__buf_2
X_82835_ _83167_/CLK _82835_/D _82835_/Q sky130_fd_sc_hd__dfxtp_4
X_55783_ _55711_/X _55783_/B _55783_/X sky130_fd_sc_hd__and2_4
X_67769_ _67766_/X _67768_/X _67769_/Y sky130_fd_sc_hd__nand2_4
X_52995_ _52999_/A _52995_/B _52995_/Y sky130_fd_sc_hd__nand2_4
X_57522_ _57519_/Y _57515_/X _57521_/Y _57522_/Y sky130_fd_sc_hd__a21boi_4
X_69508_ _88024_/Q _69506_/X _69393_/X _69507_/X _69508_/X sky130_fd_sc_hd__a211o_4
X_88342_ _88345_/CLK _40750_/X _88342_/Q sky130_fd_sc_hd__dfxtp_4
X_54734_ _54748_/A _54734_/B _54748_/C _47426_/A _54734_/X sky130_fd_sc_hd__and4_4
X_85554_ _85554_/CLK _85554_/D _85554_/Q sky130_fd_sc_hd__dfxtp_4
X_51946_ _51922_/X _51947_/A sky130_fd_sc_hd__buf_2
X_82766_ _82769_/CLK _82766_/D _82766_/Q sky130_fd_sc_hd__dfxtp_4
X_70780_ _52855_/B _70761_/X _70779_/Y _83702_/D sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_672_0_CLK clkbuf_9_336_0_CLK/X _87149_/CLK sky130_fd_sc_hd__clkbuf_1
X_84505_ _84501_/CLK _84505_/D _84505_/Q sky130_fd_sc_hd__dfxtp_4
X_57453_ _85001_/Q _57463_/B _57453_/X sky130_fd_sc_hd__or2_4
X_81717_ _81514_/CLK _81717_/D _41002_/B sky130_fd_sc_hd__dfxtp_4
X_69439_ _69696_/A _69439_/X sky130_fd_sc_hd__buf_2
X_88273_ _88288_/CLK _41127_/Y _88273_/Q sky130_fd_sc_hd__dfxtp_4
X_54665_ _85400_/Q _54648_/X _54664_/Y _54665_/Y sky130_fd_sc_hd__o21ai_4
X_85485_ _85485_/CLK _85485_/D _85485_/Q sky130_fd_sc_hd__dfxtp_4
X_51877_ _51823_/A _51877_/X sky130_fd_sc_hd__buf_2
X_82697_ _82933_/CLK _78869_/X _82685_/D sky130_fd_sc_hd__dfxtp_4
X_56404_ _56060_/X _56394_/X _56403_/Y _85207_/D sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_163_0_CLK clkbuf_8_81_0_CLK/X clkbuf_9_163_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_41630_ _41628_/X _41286_/A _41629_/X _41630_/X sky130_fd_sc_hd__o21a_4
X_87224_ _87225_/CLK _43873_/X _69033_/B sky130_fd_sc_hd__dfxtp_4
X_53616_ _53622_/A _48357_/Y _53616_/Y sky130_fd_sc_hd__nand2_4
X_72450_ _72419_/X _85349_/Q _72449_/X _72450_/Y sky130_fd_sc_hd__o21ai_4
X_84436_ _84438_/CLK _62069_/Y _78059_/B sky130_fd_sc_hd__dfxtp_4
X_50828_ _86125_/Q _50820_/X _50827_/Y _50828_/Y sky130_fd_sc_hd__o21ai_4
X_57384_ _57484_/A _57384_/X sky130_fd_sc_hd__buf_2
X_81648_ _81265_/CLK _81680_/Q _81648_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_90_0_CLK clkbuf_8_45_0_CLK/X clkbuf_9_90_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_54596_ _54600_/A _47184_/A _54596_/Y sky130_fd_sc_hd__nand2_4
X_59123_ _59121_/X _85431_/Q _59122_/X _59123_/Y sky130_fd_sc_hd__o21ai_4
X_71401_ _70673_/A _71404_/B _71399_/C _71401_/Y sky130_fd_sc_hd__nor3_4
X_56335_ _56345_/A _56335_/B _55821_/B _56335_/Y sky130_fd_sc_hd__nand3_4
X_87155_ _86932_/CLK _87155_/D _87155_/Q sky130_fd_sc_hd__dfxtp_4
X_41561_ _41560_/X _41530_/X _67041_/B _41531_/X _88192_/D sky130_fd_sc_hd__a2bb2o_4
X_53547_ _53543_/Y _53524_/X _53546_/Y _85616_/D sky130_fd_sc_hd__a21boi_4
X_72381_ _72381_/A _72381_/X sky130_fd_sc_hd__buf_2
X_84367_ _84562_/CLK _62954_/Y _84367_/Q sky130_fd_sc_hd__dfxtp_4
X_50759_ _50740_/A _52454_/B _50759_/Y sky130_fd_sc_hd__nand2_4
X_81579_ _81352_/CLK _84179_/Q _76733_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_687_0_CLK clkbuf_9_343_0_CLK/X _87446_/CLK sky130_fd_sc_hd__clkbuf_1
X_43300_ _43287_/A _43300_/X sky130_fd_sc_hd__buf_2
X_86106_ _85786_/CLK _86106_/D _86106_/Q sky130_fd_sc_hd__dfxtp_4
X_74120_ _88347_/Q _73026_/X _73028_/X _74120_/Y sky130_fd_sc_hd__o21ai_4
X_40512_ _40783_/A _40512_/X sky130_fd_sc_hd__buf_2
X_59054_ _59050_/Y _59052_/Y _59053_/X _59054_/X sky130_fd_sc_hd__a21o_4
X_71332_ _48335_/B _71320_/X _71331_/Y _83533_/D sky130_fd_sc_hd__o21ai_4
X_83318_ _83316_/CLK _83318_/D _83318_/Q sky130_fd_sc_hd__dfxtp_4
X_44280_ _44268_/A _87174_/Q _44242_/C _44280_/Y sky130_fd_sc_hd__nand3_4
X_56266_ _56159_/X _56255_/X _56265_/Y _85253_/D sky130_fd_sc_hd__o21ai_4
X_41492_ _41421_/X _82331_/Q _41491_/X _41492_/X sky130_fd_sc_hd__o21a_4
X_87086_ _87086_/CLK _44480_/X _87086_/Q sky130_fd_sc_hd__dfxtp_4
X_53478_ _53478_/A _47880_/Y _53478_/Y sky130_fd_sc_hd__nand2_4
X_84298_ _84299_/CLK _63719_/Y _80268_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_178_0_CLK clkbuf_8_89_0_CLK/X clkbuf_9_178_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_58005_ _57991_/A _86317_/Q _58005_/Y sky130_fd_sc_hd__nor2_4
X_43231_ _43231_/A _43231_/Y sky130_fd_sc_hd__inv_2
X_55217_ _45875_/A _55152_/X _55158_/A _55216_/X _72718_/D sky130_fd_sc_hd__a211o_4
X_74051_ _74051_/A _73869_/X _74051_/Y sky130_fd_sc_hd__nor2_4
X_86037_ _85527_/CLK _51299_/Y _64920_/B sky130_fd_sc_hd__dfxtp_4
X_52429_ _85824_/Q _52184_/X _52428_/Y _52429_/Y sky130_fd_sc_hd__o21ai_4
X_40443_ _40363_/X _40443_/X sky130_fd_sc_hd__buf_2
X_71263_ _70630_/B _74515_/C _71735_/C _71263_/D _71264_/A sky130_fd_sc_hd__and4_4
X_83249_ _83248_/CLK _83249_/D _61980_/A sky130_fd_sc_hd__dfxtp_4
X_56197_ _56005_/X _56195_/X _56196_/Y _56197_/Y sky130_fd_sc_hd__o21ai_4
X_73002_ _72771_/A _73003_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_610_0_CLK clkbuf_9_305_0_CLK/X _81160_/CLK sky130_fd_sc_hd__clkbuf_1
X_70214_ _70214_/A _70214_/B _83194_/Q _70204_/X _70214_/X sky130_fd_sc_hd__and4_4
X_43162_ _43162_/A _43162_/X sky130_fd_sc_hd__buf_2
X_55148_ _55147_/X _55423_/B sky130_fd_sc_hd__buf_2
X_40374_ _44532_/A _44736_/A sky130_fd_sc_hd__buf_2
X_71194_ _71197_/A _71217_/B _71194_/C _71194_/Y sky130_fd_sc_hd__nand3_4
X_42113_ _41059_/X _42103_/X _88029_/Q _42104_/X _42113_/X sky130_fd_sc_hd__a2bb2o_4
X_77810_ _77817_/A _77795_/X _77809_/Y _77811_/B sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_101_0_CLK clkbuf_8_50_0_CLK/X clkbuf_9_101_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_70145_ _83511_/Q _83159_/Q _83508_/Q _83156_/Q _70149_/A sky130_fd_sc_hd__a22oi_4
X_47970_ _66097_/B _47948_/X _47969_/Y _47970_/Y sky130_fd_sc_hd__o21ai_4
X_55079_ _55075_/Y _55076_/X _55078_/X _85323_/D sky130_fd_sc_hd__a21oi_4
X_59956_ _59875_/X _59922_/X _59931_/X _59951_/Y _59955_/X _59956_/X
+ sky130_fd_sc_hd__o41a_4
X_43093_ _43092_/Y _87579_/D sky130_fd_sc_hd__inv_2
X_78790_ _78777_/B _82816_/Q _78789_/Y _78791_/B sky130_fd_sc_hd__a21oi_4
X_87988_ _87749_/CLK _87988_/D _87988_/Q sky130_fd_sc_hd__dfxtp_4
X_58907_ _58902_/Y _58906_/Y _58883_/X _58907_/X sky130_fd_sc_hd__a21o_4
X_46921_ _54442_/B _52748_/B sky130_fd_sc_hd__buf_2
X_42044_ _42025_/A _42044_/X sky130_fd_sc_hd__buf_2
X_77741_ _78045_/A _78045_/B _77738_/Y _77741_/Y sky130_fd_sc_hd__nand3_4
X_74953_ _74947_/A _74946_/X _74958_/A _74953_/Y sky130_fd_sc_hd__a21boi_4
X_86939_ _86941_/CLK _86939_/D _67429_/B sky130_fd_sc_hd__dfxtp_4
X_70076_ _82536_/D _70067_/X _70075_/X _83856_/D sky130_fd_sc_hd__a21bo_4
X_59887_ _59885_/Y _61277_/C _59887_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_625_0_CLK clkbuf_9_312_0_CLK/X _81994_/CLK sky130_fd_sc_hd__clkbuf_1
X_49640_ _49504_/A _49641_/A sky130_fd_sc_hd__buf_2
X_73904_ _73829_/X _73904_/B _73904_/X sky130_fd_sc_hd__and2_4
X_46852_ _46817_/A _51022_/B _46852_/Y sky130_fd_sc_hd__nand2_4
X_58838_ _58928_/A _58838_/X sky130_fd_sc_hd__buf_2
X_77672_ _82239_/Q _77676_/A sky130_fd_sc_hd__inv_2
X_74884_ _81128_/D _80840_/Q _74899_/A sky130_fd_sc_hd__xor2_4
Xclkbuf_9_116_0_CLK clkbuf_8_58_0_CLK/X clkbuf_9_116_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_79411_ _84807_/Q _66420_/C _79411_/Y sky130_fd_sc_hd__nand2_4
X_45803_ _45714_/A _45803_/X sky130_fd_sc_hd__buf_2
X_76623_ _76623_/A _76624_/C sky130_fd_sc_hd__inv_2
X_49571_ _49571_/A _49571_/X sky130_fd_sc_hd__buf_2
X_73835_ _73835_/A _73835_/B _73836_/B sky130_fd_sc_hd__nand2_4
Xclkbuf_9_43_0_CLK clkbuf_9_43_0_CLK/A clkbuf_9_43_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_46783_ _54362_/D _46783_/X sky130_fd_sc_hd__buf_2
X_58769_ _84801_/Q _58769_/Y sky130_fd_sc_hd__inv_2
X_43995_ _43995_/A _59563_/A sky130_fd_sc_hd__buf_2
X_60800_ _84565_/Q _60719_/X _60796_/Y _60799_/X _84565_/D sky130_fd_sc_hd__o22a_4
X_48522_ _48522_/A _50469_/A sky130_fd_sc_hd__buf_2
X_79342_ _84801_/Q _84121_/Q _79342_/X sky130_fd_sc_hd__xor2_4
X_45734_ _45734_/A _45734_/X sky130_fd_sc_hd__buf_2
X_76554_ _76550_/Y _76554_/B _76554_/C _76554_/X sky130_fd_sc_hd__or3_4
X_42946_ _42944_/X _42945_/X _41786_/X _68051_/B _42934_/X _42946_/Y
+ sky130_fd_sc_hd__o32ai_4
X_61780_ _84726_/Q _61780_/X sky130_fd_sc_hd__buf_2
X_73766_ _73767_/B _73767_/C _73765_/X _73766_/X sky130_fd_sc_hd__a21o_4
X_70978_ _71170_/A _70979_/C sky130_fd_sc_hd__buf_2
Xclkbuf_3_1_0_CLK clkbuf_2_0_2_CLK/X clkbuf_3_1_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_75505_ _75504_/X _75505_/Y sky130_fd_sc_hd__inv_2
X_48453_ _48447_/Y _48383_/X _48452_/X _48453_/Y sky130_fd_sc_hd__a21oi_4
X_60731_ _60731_/A _63410_/A sky130_fd_sc_hd__buf_2
X_72717_ _70260_/C _72702_/X _72716_/Y _83179_/D sky130_fd_sc_hd__a21bo_4
X_79273_ _79247_/X _79271_/Y _79270_/X _79273_/X sky130_fd_sc_hd__a21bo_4
X_45665_ _56705_/B _45507_/X _45429_/X _45665_/X sky130_fd_sc_hd__o21a_4
X_76485_ _76485_/A _76484_/Y _76485_/X sky130_fd_sc_hd__xor2_4
X_42877_ _42877_/A _87673_/D sky130_fd_sc_hd__inv_2
X_73697_ _73939_/A _73697_/X sky130_fd_sc_hd__buf_2
X_47404_ _47404_/A _53025_/B _47404_/Y sky130_fd_sc_hd__nand2_4
X_78224_ _78221_/Y _78223_/X _78234_/A sky130_fd_sc_hd__nand2_4
X_44616_ _44616_/A _87031_/D sky130_fd_sc_hd__inv_2
Xclkbuf_9_58_0_CLK clkbuf_9_59_0_CLK/A clkbuf_9_58_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_63450_ _63427_/A _61844_/X _63450_/X sky130_fd_sc_hd__and2_4
X_75436_ _75436_/A _75436_/Y sky130_fd_sc_hd__inv_2
X_41828_ _41824_/X _41825_/X _40452_/X _66920_/B _41821_/X _41829_/A
+ sky130_fd_sc_hd__o32ai_4
X_48384_ _48384_/A _48384_/Y sky130_fd_sc_hd__inv_2
X_72648_ _72656_/A _72656_/B _72648_/C _72648_/Y sky130_fd_sc_hd__nand3_4
X_60662_ _60662_/A _60720_/A sky130_fd_sc_hd__inv_2
X_45596_ _45596_/A _45596_/X sky130_fd_sc_hd__buf_2
X_62401_ _61492_/A _62332_/B _62386_/C _62431_/D _62401_/Y sky130_fd_sc_hd__nand4_4
X_47335_ _47334_/Y _52991_/B sky130_fd_sc_hd__buf_2
X_78155_ _78154_/A _78154_/B _78162_/C sky130_fd_sc_hd__nand2_4
X_44547_ _44547_/A _44547_/X sky130_fd_sc_hd__buf_2
X_63381_ _63368_/X _63369_/X _63373_/X _63377_/X _63380_/Y _63381_/Y
+ sky130_fd_sc_hd__o41ai_4
X_75367_ _75347_/X _75366_/Y _75339_/Y _75367_/Y sky130_fd_sc_hd__o21ai_4
X_41759_ _41759_/A _41759_/Y sky130_fd_sc_hd__inv_2
X_60593_ _60593_/A _60593_/B _60594_/A sky130_fd_sc_hd__nor2_4
X_72579_ _72579_/A _72579_/B _72579_/Y sky130_fd_sc_hd__nand2_4
X_65120_ _65227_/A _65120_/B _65120_/X sky130_fd_sc_hd__and2_4
X_77106_ _77106_/A _77112_/C _77109_/A sky130_fd_sc_hd__nand2_4
X_62332_ _61430_/A _62332_/B _62631_/C _62332_/D _62335_/B sky130_fd_sc_hd__nand4_4
X_74318_ _70301_/C _74314_/X _74317_/Y _74318_/X sky130_fd_sc_hd__a21bo_4
X_47266_ _47262_/Y _47224_/X _47265_/X _47266_/Y sky130_fd_sc_hd__a21oi_4
X_78086_ _82659_/Q _78085_/Y _78086_/X sky130_fd_sc_hd__xor2_4
X_44478_ _44478_/A _87088_/D sky130_fd_sc_hd__inv_2
X_75298_ _75287_/Y _75288_/Y _75289_/Y _75298_/X sky130_fd_sc_hd__o21a_4
X_49005_ _49005_/A _53841_/B sky130_fd_sc_hd__inv_2
X_65051_ _65836_/A _65051_/B _65051_/X sky130_fd_sc_hd__and2_4
X_46217_ _46222_/A _46217_/B _46217_/C _46217_/Y sky130_fd_sc_hd__nand3_4
X_77037_ _77030_/Y _77035_/Y _77036_/Y _77041_/C sky130_fd_sc_hd__a21o_4
XPHY_290 sky130_fd_sc_hd__decap_3
X_43429_ _41552_/X _43412_/X _87426_/Q _43413_/X _43429_/X sky130_fd_sc_hd__a2bb2o_4
X_62263_ _62212_/A _62260_/Y _62261_/Y _62262_/Y _62263_/Y sky130_fd_sc_hd__nand4_4
X_74249_ _88341_/Q _73801_/X _73087_/X _74249_/Y sky130_fd_sc_hd__o21ai_4
X_47197_ _59361_/A _47192_/X _47196_/Y _47197_/Y sky130_fd_sc_hd__o21ai_4
X_64002_ _63561_/B _63955_/X _64050_/C _64033_/D _64002_/Y sky130_fd_sc_hd__nand4_4
X_61214_ _61188_/C _61214_/Y sky130_fd_sc_hd__inv_2
Xpsn_inst_psn_buff_17 _44274_/D _44307_/D sky130_fd_sc_hd__buf_2
X_46148_ _49520_/A _49380_/C sky130_fd_sc_hd__buf_2
Xpsn_inst_psn_buff_28 _50212_/A _50218_/A sky130_fd_sc_hd__buf_2
X_62194_ _62194_/A _84905_/Q _62618_/D _62194_/D _62194_/X sky130_fd_sc_hd__and4_4
X_68810_ _68807_/X _68809_/X _68737_/X _68810_/Y sky130_fd_sc_hd__a21oi_4
X_61145_ _64221_/A _61145_/X sky130_fd_sc_hd__buf_2
X_46079_ _46067_/X _43046_/A _41615_/X _86777_/Q _46068_/X _46080_/A
+ sky130_fd_sc_hd__o32ai_4
X_69790_ _69790_/A _69790_/Y sky130_fd_sc_hd__inv_2
X_78988_ _78978_/B _82517_/D sky130_fd_sc_hd__inv_2
X_49907_ _49854_/A _49928_/A sky130_fd_sc_hd__buf_2
X_68741_ _69779_/A _68741_/X sky130_fd_sc_hd__buf_2
X_65953_ _65949_/X _65868_/B _65952_/X _65953_/Y sky130_fd_sc_hd__nand3_4
X_61076_ _61075_/X _60631_/D _61144_/A sky130_fd_sc_hd__and2_4
X_77939_ _77933_/A _77933_/B _77939_/Y sky130_fd_sc_hd__nor2_4
X_64904_ _64904_/A _64904_/B _64904_/X sky130_fd_sc_hd__and2_4
X_60027_ _60027_/A _60027_/X sky130_fd_sc_hd__buf_2
X_49838_ _58038_/B _49825_/X _49837_/Y _49838_/Y sky130_fd_sc_hd__o21ai_4
X_80950_ _81996_/CLK _80950_/D _74993_/A sky130_fd_sc_hd__dfxtp_4
X_68672_ _68746_/A _68672_/B _68672_/Y sky130_fd_sc_hd__nor2_4
X_65884_ _65884_/A _65884_/B _65884_/Y sky130_fd_sc_hd__nand2_4
X_67623_ _67623_/A _67623_/B _67623_/Y sky130_fd_sc_hd__nand2_4
X_79609_ _79609_/A _79609_/B _79610_/A sky130_fd_sc_hd__nand2_4
X_64835_ _64598_/X _64835_/X sky130_fd_sc_hd__buf_2
X_49769_ _49688_/X _49769_/X sky130_fd_sc_hd__buf_2
X_80881_ _80849_/CLK _75712_/B _80881_/Q sky130_fd_sc_hd__dfxtp_4
X_51800_ _51796_/A _51800_/B _51800_/Y sky130_fd_sc_hd__nand2_4
X_82620_ _82589_/CLK _79047_/B _82620_/Q sky130_fd_sc_hd__dfxtp_4
X_67554_ _86966_/Q _67551_/X _67552_/X _67553_/X _67555_/B sky130_fd_sc_hd__a211o_4
X_52780_ _52778_/Y _52755_/X _52779_/X _52780_/Y sky130_fd_sc_hd__a21oi_4
X_64766_ _64766_/A _64766_/X sky130_fd_sc_hd__buf_2
X_61978_ _61974_/Y _61959_/X _61977_/Y _84442_/D sky130_fd_sc_hd__a21oi_4
X_66505_ _64867_/B _66501_/B _84110_/Q _66505_/X sky130_fd_sc_hd__and3_4
X_51731_ _51729_/Y _51719_/X _51730_/X _85956_/D sky130_fd_sc_hd__a21oi_4
X_63717_ _63712_/Y _63715_/X _63716_/X _84866_/Q _63363_/A _63717_/Y
+ sky130_fd_sc_hd__o32ai_4
X_82551_ _82553_/CLK _83871_/Q _82551_/Q sky130_fd_sc_hd__dfxtp_4
X_60929_ _60928_/X _60930_/C sky130_fd_sc_hd__buf_2
X_67485_ _67460_/A _87725_/Q _67485_/X sky130_fd_sc_hd__and2_4
X_64697_ _64642_/A _64697_/X sky130_fd_sc_hd__buf_2
X_81502_ _81461_/CLK _81502_/D _76906_/A sky130_fd_sc_hd__dfxtp_4
X_69224_ _69253_/A _69224_/B _69224_/X sky130_fd_sc_hd__and2_4
X_54450_ _54447_/Y _54448_/X _54449_/X _85440_/D sky130_fd_sc_hd__a21oi_4
X_66436_ _66116_/X _66517_/B _66120_/X _66436_/Y sky130_fd_sc_hd__nand3_4
X_85270_ _85270_/CLK _85270_/D _56221_/C sky130_fd_sc_hd__dfxtp_4
X_51662_ _51608_/A _51684_/C sky130_fd_sc_hd__buf_2
X_63648_ _59423_/Y _63648_/B _63648_/Y sky130_fd_sc_hd__nor2_4
X_82482_ _82610_/CLK _82482_/D _82858_/D sky130_fd_sc_hd__dfxtp_4
X_53401_ _53347_/A _53402_/B sky130_fd_sc_hd__buf_2
X_84221_ _81224_/CLK _84221_/D _84221_/Q sky130_fd_sc_hd__dfxtp_4
X_50613_ _86167_/Q _50594_/X _50612_/Y _50613_/Y sky130_fd_sc_hd__o21ai_4
X_81433_ _81433_/CLK _81465_/Q _76085_/B sky130_fd_sc_hd__dfxtp_4
X_69155_ _87038_/Q _69153_/X _68891_/X _69154_/X _69155_/X sky130_fd_sc_hd__a211o_4
X_54381_ _54379_/Y _54366_/X _54380_/X _85453_/D sky130_fd_sc_hd__a21oi_4
X_66367_ _65923_/X _66367_/B _65927_/C _66367_/Y sky130_fd_sc_hd__nand3_4
X_51593_ _51591_/Y _51585_/X _51592_/X _51593_/Y sky130_fd_sc_hd__a21oi_4
X_63579_ _63554_/A _63554_/B _80442_/B _63579_/Y sky130_fd_sc_hd__nor3_4
X_56120_ _55801_/D _56120_/B _56121_/A sky130_fd_sc_hd__xor2_4
X_68106_ _68106_/A _68106_/X sky130_fd_sc_hd__buf_2
X_53332_ _53332_/A _53332_/B _53332_/Y sky130_fd_sc_hd__nand2_4
X_65318_ _72296_/A _66423_/B sky130_fd_sc_hd__buf_2
X_84152_ _81224_/CLK _66165_/X _84152_/Q sky130_fd_sc_hd__dfxtp_4
X_50544_ _50542_/Y _50525_/X _50543_/X _86181_/D sky130_fd_sc_hd__a21oi_4
X_81364_ _81461_/CLK _81364_/D _76424_/A sky130_fd_sc_hd__dfxtp_4
X_69086_ _69086_/A _87317_/Q _69086_/X sky130_fd_sc_hd__and2_4
X_66298_ _66237_/X _66298_/B _66298_/X sky130_fd_sc_hd__and2_4
X_83103_ _83095_/CLK _74311_/X _83103_/Q sky130_fd_sc_hd__dfxtp_4
X_80315_ _80315_/A _80313_/Y _80314_/Y _80317_/B sky130_fd_sc_hd__nand3_4
X_56051_ _56104_/A _56052_/A sky130_fd_sc_hd__buf_2
X_68037_ _68034_/X _68036_/X _67897_/X _68037_/Y sky130_fd_sc_hd__a21oi_4
X_53263_ _51902_/A _54442_/B _53263_/Y sky130_fd_sc_hd__nand2_4
X_65249_ _65227_/A _65249_/B _65249_/X sky130_fd_sc_hd__and2_4
X_84083_ _84105_/CLK _67116_/X _80907_/D sky130_fd_sc_hd__dfxtp_4
X_50475_ _48533_/A _50475_/B _50257_/X _50475_/Y sky130_fd_sc_hd__nand3_4
X_81295_ _81615_/CLK _76983_/X _81295_/Q sky130_fd_sc_hd__dfxtp_4
X_55002_ _55011_/A _47598_/A _55002_/Y sky130_fd_sc_hd__nand2_4
X_52214_ _52214_/A _52214_/X sky130_fd_sc_hd__buf_2
X_83034_ _85180_/CLK _74563_/Y _83034_/Q sky130_fd_sc_hd__dfxtp_4
X_87911_ _86930_/CLK _87911_/D _87911_/Q sky130_fd_sc_hd__dfxtp_4
X_80246_ _80230_/Y _80233_/Y _80245_/X _80246_/X sky130_fd_sc_hd__a21o_4
X_53194_ _85679_/Q _53172_/X _53193_/Y _53194_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_opt_24_CLK _86499_/CLK _86470_/CLK sky130_fd_sc_hd__clkbuf_16
X_59810_ _59810_/A _59743_/B _59810_/Y sky130_fd_sc_hd__nor2_4
X_52145_ _52203_/A _52145_/X sky130_fd_sc_hd__buf_2
X_87842_ _88097_/CLK _87842_/D _68801_/A sky130_fd_sc_hd__dfxtp_4
X_80177_ _80173_/Y _80176_/Y _80198_/A sky130_fd_sc_hd__xor2_4
X_69988_ _69988_/A _69988_/X sky130_fd_sc_hd__buf_2
X_59741_ _59741_/A _62669_/D _59741_/C _59742_/A sky130_fd_sc_hd__and3_4
X_52076_ _52185_/A _52121_/A sky130_fd_sc_hd__buf_2
X_56953_ _56953_/A _56953_/X sky130_fd_sc_hd__buf_2
X_68939_ _44727_/A _68818_/X _68819_/X _68938_/X _68940_/B sky130_fd_sc_hd__a211o_4
X_87773_ _87767_/CLK _87773_/D _87773_/Q sky130_fd_sc_hd__dfxtp_4
X_84985_ _85915_/CLK _84985_/D _84985_/Q sky130_fd_sc_hd__dfxtp_4
X_51027_ _86087_/Q _51020_/X _51026_/Y _51027_/Y sky130_fd_sc_hd__o21ai_4
X_55904_ _85273_/Q _44106_/C _44051_/A _55903_/X _55904_/X sky130_fd_sc_hd__a211o_4
X_86724_ _86404_/CLK _46584_/Y _86724_/Q sky130_fd_sc_hd__dfxtp_4
X_71950_ _55663_/Y _71939_/X _71949_/Y _71950_/Y sky130_fd_sc_hd__o21ai_4
X_59672_ _57701_/A _59770_/A sky130_fd_sc_hd__buf_2
X_83936_ _81346_/CLK _83936_/D _81400_/D sky130_fd_sc_hd__dfxtp_4
X_56884_ _56691_/A _56884_/B _56884_/C _56884_/Y sky130_fd_sc_hd__nand3_4
X_70901_ _70873_/A _70903_/B _70899_/C _70899_/D _70901_/Y sky130_fd_sc_hd__nand4_4
X_58623_ _58623_/A _58623_/Y sky130_fd_sc_hd__inv_2
X_55835_ _55832_/X _55834_/X _44113_/X _56088_/A sky130_fd_sc_hd__a21o_4
X_86655_ _86655_/CLK _86655_/D _57734_/A sky130_fd_sc_hd__dfxtp_4
X_71881_ _70552_/Y _71883_/B _71873_/X _71883_/D _71881_/Y sky130_fd_sc_hd__nor4_4
X_83867_ _82541_/CLK _70036_/X _82547_/D sky130_fd_sc_hd__dfxtp_4
X_42800_ _42799_/Y _87712_/D sky130_fd_sc_hd__inv_2
X_85606_ _86534_/CLK _85606_/D _85606_/Q sky130_fd_sc_hd__dfxtp_4
X_73620_ _73601_/X _73604_/Y _73619_/X _73620_/X sky130_fd_sc_hd__a21o_4
X_70832_ _70832_/A _71066_/C sky130_fd_sc_hd__buf_2
X_58554_ _58554_/A _58557_/B _58554_/Y sky130_fd_sc_hd__nand2_4
X_82818_ _82828_/CLK _82818_/D _82818_/Q sky130_fd_sc_hd__dfxtp_4
X_43780_ _43779_/Y _43780_/Y sky130_fd_sc_hd__inv_2
X_55766_ _55741_/A _85161_/Q _55766_/X sky130_fd_sc_hd__and2_4
X_86586_ _86554_/CLK _47921_/Y _66008_/B sky130_fd_sc_hd__dfxtp_4
X_40992_ _82294_/Q _40970_/B _40992_/X sky130_fd_sc_hd__or2_4
X_52978_ _52974_/Y _52975_/X _52977_/X _85720_/D sky130_fd_sc_hd__a21oi_4
X_83798_ _83819_/CLK _83798_/D _74782_/B sky130_fd_sc_hd__dfxtp_4
X_57505_ _47363_/A _71978_/A sky130_fd_sc_hd__buf_2
X_42731_ _41203_/X _42717_/X _68790_/B _42718_/X _87746_/D sky130_fd_sc_hd__a2bb2o_4
X_88325_ _88060_/CLK _88325_/D _69756_/B sky130_fd_sc_hd__dfxtp_4
X_54717_ _54715_/Y _54694_/X _54716_/X _54717_/Y sky130_fd_sc_hd__a21oi_4
X_73551_ _72889_/X _73551_/X sky130_fd_sc_hd__buf_2
X_85537_ _86145_/CLK _85537_/D _85537_/Q sky130_fd_sc_hd__dfxtp_4
X_51929_ _51928_/X _51929_/X sky130_fd_sc_hd__buf_2
X_70763_ _70763_/A _70860_/A sky130_fd_sc_hd__buf_2
X_82749_ _82748_/CLK _84133_/Q _82749_/Q sky130_fd_sc_hd__dfxtp_4
X_58485_ _83413_/Q _58485_/Y sky130_fd_sc_hd__inv_2
X_55697_ _55693_/X _55696_/X _55615_/X _55700_/A sky130_fd_sc_hd__a21o_4
X_72502_ _72502_/A _72516_/C sky130_fd_sc_hd__buf_2
X_45450_ _45448_/Y _45449_/Y _44901_/X _45450_/X sky130_fd_sc_hd__o21a_4
X_57436_ _57275_/X _57170_/A _57435_/X _57436_/X sky130_fd_sc_hd__o21a_4
X_76270_ _76237_/Y _76253_/Y _76255_/A _76270_/X sky130_fd_sc_hd__o21a_4
X_88256_ _87757_/CLK _41216_/Y _88256_/Q sky130_fd_sc_hd__dfxtp_4
X_42662_ _42661_/Y _42662_/Y sky130_fd_sc_hd__inv_2
X_54648_ _54729_/A _54648_/X sky130_fd_sc_hd__buf_2
X_73482_ _73480_/X _73481_/Y _73367_/X _73482_/Y sky130_fd_sc_hd__a21oi_4
X_85468_ _82206_/CLK _54299_/Y _85468_/Q sky130_fd_sc_hd__dfxtp_4
X_70694_ _70694_/A _70412_/X _70933_/B _70627_/A _70695_/A sky130_fd_sc_hd__nand4_4
X_44401_ _41503_/X _44394_/X _87127_/Q _44395_/X _87127_/D sky130_fd_sc_hd__a2bb2o_4
X_75221_ _80780_/Q _81036_/D _80748_/D sky130_fd_sc_hd__xor2_4
X_41613_ _41825_/A _41613_/X sky130_fd_sc_hd__buf_2
X_87207_ _87149_/CLK _87207_/D _67616_/B sky130_fd_sc_hd__dfxtp_4
X_72433_ _72352_/X _85959_/Q _72432_/X _72433_/Y sky130_fd_sc_hd__o21ai_4
X_84419_ _84538_/CLK _84419_/D _76995_/B sky130_fd_sc_hd__dfxtp_4
X_45381_ _45381_/A _45381_/B _45381_/Y sky130_fd_sc_hd__nand2_4
X_57367_ _57244_/X _56917_/A _57366_/Y _57368_/A sky130_fd_sc_hd__o21ai_4
X_88187_ _87110_/CLK _88187_/D _67161_/B sky130_fd_sc_hd__dfxtp_4
X_54579_ _85416_/Q _54567_/X _54578_/Y _54579_/Y sky130_fd_sc_hd__o21ai_4
X_42593_ _42590_/X _42592_/X _40861_/X _69804_/A _42580_/X _42593_/Y
+ sky130_fd_sc_hd__o32ai_4
X_85399_ _85492_/CLK _85399_/D _85399_/Q sky130_fd_sc_hd__dfxtp_4
X_47120_ _54559_/D _52867_/D sky130_fd_sc_hd__buf_2
X_59106_ _58847_/A _59106_/X sky130_fd_sc_hd__buf_2
X_44332_ _44736_/A _44332_/X sky130_fd_sc_hd__buf_2
X_56318_ _56064_/X _56305_/X _56317_/Y _85238_/D sky130_fd_sc_hd__o21ai_4
X_75152_ _80680_/Q _75151_/B _75153_/A sky130_fd_sc_hd__nand2_4
X_87138_ _87382_/CLK _87138_/D _87138_/Q sky130_fd_sc_hd__dfxtp_4
X_41544_ _41344_/X _81169_/Q _41543_/X _41544_/X sky130_fd_sc_hd__o21a_4
X_72364_ _72327_/X _85965_/Q _72363_/X _72364_/Y sky130_fd_sc_hd__o21ai_4
X_57298_ _57049_/A _85038_/Q _57326_/C _57298_/Y sky130_fd_sc_hd__nor3_4
X_74103_ _72905_/A _74103_/X sky130_fd_sc_hd__buf_2
X_47051_ _46909_/X _47063_/A sky130_fd_sc_hd__buf_2
X_59037_ _59037_/A _59037_/X sky130_fd_sc_hd__buf_2
X_71315_ _52047_/B _71289_/Y _71314_/Y _71315_/Y sky130_fd_sc_hd__o21ai_4
X_44263_ _64725_/A _44263_/X sky130_fd_sc_hd__buf_2
Xclkbuf_6_40_0_CLK clkbuf_6_41_0_CLK/A clkbuf_7_81_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_56249_ _56121_/X _56242_/X _56248_/Y _56249_/Y sky130_fd_sc_hd__o21ai_4
X_75083_ _80675_/Q _75082_/B _75102_/B sky130_fd_sc_hd__nand2_4
X_79960_ _79942_/A _79940_/Y _79959_/Y _79960_/Y sky130_fd_sc_hd__a21oi_4
X_41475_ _41399_/X _41400_/X _41473_/X _66656_/B _41474_/X _41476_/A
+ sky130_fd_sc_hd__o32ai_4
X_87069_ _88337_/CLK _44521_/Y _87069_/Q sky130_fd_sc_hd__dfxtp_4
X_72295_ _72295_/A _72332_/B _72295_/Y sky130_fd_sc_hd__nor2_4
X_46002_ _45994_/X _46001_/X _40479_/X _86820_/Q _45995_/X _46002_/Y
+ sky130_fd_sc_hd__o32ai_4
X_43214_ _43214_/A _87535_/D sky130_fd_sc_hd__inv_2
X_74034_ _68861_/B _73872_/X _73894_/X _74033_/Y _74034_/X sky130_fd_sc_hd__a211o_4
X_78911_ _82814_/D _82558_/Q _78912_/B sky130_fd_sc_hd__xnor2_4
X_40426_ _40425_/X _40426_/X sky130_fd_sc_hd__buf_2
X_71246_ _71252_/A _71246_/B _71248_/C _71246_/Y sky130_fd_sc_hd__nand3_4
X_44194_ _73948_/A _44194_/X sky130_fd_sc_hd__buf_2
X_79891_ _79882_/A _79881_/X _79889_/A _79891_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_opt_15_CLK _84518_/CLK _84640_/CLK sky130_fd_sc_hd__clkbuf_16
X_43145_ _43145_/A _43145_/Y sky130_fd_sc_hd__inv_2
X_78842_ _78841_/B _78833_/Y _78842_/Y sky130_fd_sc_hd__nor2_4
X_40357_ _40344_/A _40435_/A sky130_fd_sc_hd__inv_2
X_71177_ _71145_/A _71185_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_564_0_CLK clkbuf_9_282_0_CLK/X _84074_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_55_0_CLK clkbuf_6_55_0_CLK/A clkbuf_6_55_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_70128_ _70128_/A _83122_/Q _70128_/C _83120_/Q _70131_/A sky130_fd_sc_hd__nor4_4
X_47953_ _73830_/B _47948_/X _47952_/Y _47953_/Y sky130_fd_sc_hd__o21ai_4
X_43076_ _43072_/X _43075_/X _40691_/X _73989_/A _43061_/X _43076_/Y
+ sky130_fd_sc_hd__o32ai_4
X_59939_ _59918_/Y _62463_/A sky130_fd_sc_hd__buf_2
X_78773_ _78737_/Y _78770_/D _78770_/B _78773_/X sky130_fd_sc_hd__a21bo_4
X_75985_ _75980_/Y _75981_/A _75984_/Y _75986_/B sky130_fd_sc_hd__a21boi_4
X_46904_ _82947_/Q _54435_/D sky130_fd_sc_hd__inv_2
X_42027_ _42027_/A _42027_/Y sky130_fd_sc_hd__inv_2
X_77724_ _77724_/A _77724_/B _81921_/D sky130_fd_sc_hd__nand2_4
X_62950_ _62945_/Y _62946_/X _62949_/Y _58352_/A _62650_/X _62950_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74936_ _81135_/D _74945_/B _74942_/B sky130_fd_sc_hd__xor2_4
X_70059_ _82541_/D _70048_/X _70058_/X _70059_/X sky130_fd_sc_hd__a21bo_4
X_47884_ _47943_/A _82941_/Q _47884_/X sky130_fd_sc_hd__or2_4
X_61901_ _61915_/A _61915_/B _63496_/B _61915_/D _61901_/X sky130_fd_sc_hd__and4_4
X_49623_ _49570_/A _49623_/X sky130_fd_sc_hd__buf_2
X_46835_ _58867_/A _46813_/X _46834_/Y _46835_/Y sky130_fd_sc_hd__o21ai_4
X_77655_ _77655_/A _77652_/Y _77654_/Y _77660_/A sky130_fd_sc_hd__or3_4
X_62881_ _62877_/X _62831_/X _62878_/Y _62879_/Y _62880_/X _62881_/X
+ sky130_fd_sc_hd__a41o_4
X_74867_ _74867_/A _74866_/Y _74868_/B sky130_fd_sc_hd__xor2_4
Xclkbuf_10_579_0_CLK clkbuf_9_289_0_CLK/X _80804_/CLK sky130_fd_sc_hd__clkbuf_1
X_64620_ _64612_/X _64618_/X _64619_/X _64623_/A sky130_fd_sc_hd__a21o_4
X_76606_ _76604_/Y _76605_/X _81631_/D sky130_fd_sc_hd__xor2_4
X_49554_ _49558_/A _52768_/B _49554_/Y sky130_fd_sc_hd__nand2_4
X_61832_ _61831_/X _61765_/B _61846_/C _61846_/D _61832_/Y sky130_fd_sc_hd__nand4_4
X_73818_ _73939_/A _73818_/X sky130_fd_sc_hd__buf_2
X_46766_ _72052_/A _46767_/A sky130_fd_sc_hd__buf_2
X_77586_ _77570_/A _77567_/Y _77568_/Y _77586_/X sky130_fd_sc_hd__o21a_4
X_43978_ _44160_/B _43978_/Y sky130_fd_sc_hd__inv_2
X_74798_ _74794_/Y _74798_/B _74796_/Y _74798_/D _74798_/X sky130_fd_sc_hd__and4_4
X_48505_ _48515_/A _52163_/B _48505_/Y sky130_fd_sc_hd__nand2_4
X_79325_ _79316_/Y _79334_/B _79324_/X _79325_/Y sky130_fd_sc_hd__a21boi_4
X_45717_ _45668_/X _61572_/A _45685_/X _45717_/Y sky130_fd_sc_hd__o21ai_4
X_64551_ _64542_/Y _64532_/X _64550_/Y _84235_/D sky130_fd_sc_hd__o21ai_4
X_76537_ _76520_/Y _76521_/Y _76522_/Y _76537_/X sky130_fd_sc_hd__o21a_4
X_42929_ _41741_/X _42920_/X _67832_/B _42922_/X _87646_/D sky130_fd_sc_hd__a2bb2o_4
X_49485_ _49481_/A _51008_/B _49485_/Y sky130_fd_sc_hd__nand2_4
X_61763_ _61711_/X _61856_/A sky130_fd_sc_hd__buf_2
X_73749_ _70107_/B _73697_/X _73748_/X _73749_/Y sky130_fd_sc_hd__o21ai_4
X_46697_ _54312_/D _52622_/D sky130_fd_sc_hd__buf_2
Xclkbuf_10_502_0_CLK clkbuf_9_251_0_CLK/X _86100_/CLK sky130_fd_sc_hd__clkbuf_1
X_63502_ _63512_/A _57664_/A _63476_/C _63502_/X sky130_fd_sc_hd__and3_4
X_48436_ _86522_/Q _48419_/X _48435_/Y _48436_/Y sky130_fd_sc_hd__o21ai_4
X_60714_ _60714_/A _63417_/A _60725_/A _60714_/Y sky130_fd_sc_hd__nand3_4
X_67270_ _66673_/X _67270_/X sky130_fd_sc_hd__buf_2
X_79256_ _79244_/X _79246_/B _79255_/Y _79256_/Y sky130_fd_sc_hd__a21boi_4
X_45648_ _57409_/A _45354_/X _45648_/Y sky130_fd_sc_hd__nor2_4
X_64482_ _64480_/Y _64186_/X _64481_/Y _64482_/Y sky130_fd_sc_hd__a21oi_4
X_76468_ _76464_/Y _76468_/B _76469_/B sky130_fd_sc_hd__xor2_4
X_61694_ _61292_/A _61694_/B _61675_/C _61694_/Y sky130_fd_sc_hd__nand3_4
X_66221_ _66125_/X _86219_/Q _66180_/X _66220_/X _66221_/X sky130_fd_sc_hd__a211o_4
X_78207_ _78198_/A _82491_/Q _78207_/Y sky130_fd_sc_hd__nand2_4
X_63433_ _63431_/Y _63391_/X _63432_/Y _63433_/Y sky130_fd_sc_hd__a21oi_4
X_75419_ _75435_/B _75435_/D _75419_/X sky130_fd_sc_hd__and2_4
X_48367_ _83592_/Q _48367_/Y sky130_fd_sc_hd__inv_2
X_60645_ _60644_/X _60687_/A sky130_fd_sc_hd__buf_2
X_79187_ _79186_/Y _79180_/Y _79181_/Y _79188_/B sky130_fd_sc_hd__nand3_4
X_45579_ _45511_/X _61468_/A _45530_/X _45579_/Y sky130_fd_sc_hd__o21ai_4
X_76399_ _76399_/A _76400_/C sky130_fd_sc_hd__inv_2
X_47318_ _47130_/A _47349_/B sky130_fd_sc_hd__buf_2
X_66152_ _66149_/Y _66137_/X _66151_/X _66152_/X sky130_fd_sc_hd__a21o_4
X_78138_ _78129_/X _78137_/Y _78139_/B sky130_fd_sc_hd__xor2_4
X_63364_ _63354_/Y _63360_/X _63361_/X _58147_/A _63363_/X _63364_/Y
+ sky130_fd_sc_hd__o32ai_4
X_60576_ _58094_/A _72250_/A sky130_fd_sc_hd__buf_2
X_48298_ _48275_/X _48297_/X _48298_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_517_0_CLK clkbuf_9_258_0_CLK/X _81473_/CLK sky130_fd_sc_hd__clkbuf_1
X_65103_ _64929_/A _65103_/B _65103_/X sky130_fd_sc_hd__and2_4
X_62315_ _62304_/A _58248_/A _62315_/C _62286_/X _62315_/X sky130_fd_sc_hd__and4_4
X_47249_ _47246_/X _47228_/B _47234_/X _52938_/D _47249_/X sky130_fd_sc_hd__and4_4
X_66083_ _64598_/X _86229_/Q _65761_/X _66082_/X _66083_/X sky130_fd_sc_hd__a211o_4
X_78069_ _60755_/C _78069_/B _78069_/X sky130_fd_sc_hd__xor2_4
X_63295_ _63295_/A _63316_/B _63295_/C _63344_/D _63295_/X sky130_fd_sc_hd__or4_4
X_80100_ _80092_/A _80091_/X _80099_/Y _80117_/B sky130_fd_sc_hd__a21boi_4
X_65034_ _65034_/A _65859_/A sky130_fd_sc_hd__buf_2
X_69911_ _69865_/A _88313_/Q _69911_/X sky130_fd_sc_hd__and2_4
X_50260_ _50251_/X _50260_/B _50260_/Y sky130_fd_sc_hd__nand2_4
X_62246_ _59931_/X _61762_/X _62245_/X _62246_/X sky130_fd_sc_hd__a21o_4
X_81080_ _80696_/CLK _81112_/Q _75392_/A sky130_fd_sc_hd__dfxtp_4
X_80031_ _80023_/A _80008_/X _80031_/X sky130_fd_sc_hd__and2_4
X_69842_ _69900_/A _69842_/B _69842_/X sky130_fd_sc_hd__and2_4
X_50191_ _51263_/A _50191_/X sky130_fd_sc_hd__buf_2
X_62177_ _62169_/X _62171_/X _62176_/Y _84867_/Q _61782_/A _62177_/Y
+ sky130_fd_sc_hd__o32ai_4
X_61128_ _61128_/A _64303_/A sky130_fd_sc_hd__buf_2
X_69773_ _69347_/X _69349_/X _69728_/X _69773_/Y sky130_fd_sc_hd__a21oi_4
X_66985_ _66961_/X _66985_/B _66985_/X sky130_fd_sc_hd__and2_4
X_68724_ _87089_/Q _68353_/X _68354_/X _68723_/X _68724_/X sky130_fd_sc_hd__a211o_4
X_53950_ _53947_/Y _53948_/X _53949_/Y _53950_/Y sky130_fd_sc_hd__a21boi_4
X_65936_ _65859_/X _85631_/Q _65860_/X _65935_/X _65936_/X sky130_fd_sc_hd__a211o_4
X_61059_ _60994_/A _60998_/X _59846_/X _60992_/X _61059_/X sky130_fd_sc_hd__a211o_4
X_84770_ _85375_/CLK _59092_/Y _84770_/Q sky130_fd_sc_hd__dfxtp_4
X_81982_ _83906_/CLK _83910_/Q _77833_/B sky130_fd_sc_hd__dfxtp_4
X_52901_ _52898_/Y _52892_/X _52900_/X _52901_/Y sky130_fd_sc_hd__a21oi_4
X_83721_ _83721_/CLK _70709_/Y _46920_/A sky130_fd_sc_hd__dfxtp_4
X_68655_ _87496_/Q _68626_/X _68601_/X _68654_/X _68655_/X sky130_fd_sc_hd__a211o_4
X_80933_ _81061_/CLK _75109_/B _80933_/Q sky130_fd_sc_hd__dfxtp_4
X_53881_ _53871_/X _49083_/A _53881_/Y sky130_fd_sc_hd__nand2_4
X_65867_ _65811_/X _83052_/Q _65865_/X _65866_/X _65867_/X sky130_fd_sc_hd__a211o_4
X_55620_ _55620_/A _55947_/A sky130_fd_sc_hd__buf_2
X_67606_ _87400_/Q _67512_/X _67581_/X _67605_/X _67606_/X sky130_fd_sc_hd__a211o_4
X_86440_ _83594_/CLK _86440_/D _65253_/B sky130_fd_sc_hd__dfxtp_4
X_52832_ _52830_/Y _52809_/X _52831_/X _52832_/Y sky130_fd_sc_hd__a21oi_4
X_64818_ _64778_/A _85817_/Q _64818_/X sky130_fd_sc_hd__and2_4
X_83652_ _86139_/CLK _83652_/D _46313_/A sky130_fd_sc_hd__dfxtp_4
X_68586_ _68586_/A _68586_/X sky130_fd_sc_hd__buf_2
X_80864_ _81994_/CLK _80896_/Q _75061_/B sky130_fd_sc_hd__dfxtp_4
X_65798_ _65660_/X _83057_/Q _65768_/X _65797_/X _65798_/X sky130_fd_sc_hd__a211o_4
X_82603_ _82570_/CLK _78889_/B _82571_/D sky130_fd_sc_hd__dfxtp_4
X_67537_ _87403_/Q _67512_/X _67462_/X _67536_/X _67537_/X sky130_fd_sc_hd__a211o_4
X_55551_ _56616_/A _55546_/X _56616_/B _55550_/X _55552_/A sky130_fd_sc_hd__and4_4
X_86371_ _83660_/CLK _49529_/Y _86371_/Q sky130_fd_sc_hd__dfxtp_4
X_52763_ _52775_/A _52746_/B _52775_/C _52763_/D _52763_/X sky130_fd_sc_hd__and4_4
X_64749_ _64810_/A _64749_/B _64749_/X sky130_fd_sc_hd__and2_4
X_83583_ _83068_/CLK _71174_/Y _83583_/Q sky130_fd_sc_hd__dfxtp_4
X_80795_ _80818_/CLK _80795_/D _80795_/Q sky130_fd_sc_hd__dfxtp_4
X_88110_ _88111_/CLK _88110_/D _73675_/A sky130_fd_sc_hd__dfxtp_4
X_54502_ _54475_/A _54502_/X sky130_fd_sc_hd__buf_2
X_85322_ _85351_/CLK _85322_/D _85322_/Q sky130_fd_sc_hd__dfxtp_4
X_51714_ _51608_/A _51715_/C sky130_fd_sc_hd__buf_2
X_58270_ _46155_/A _58328_/A sky130_fd_sc_hd__buf_2
X_82534_ _82536_/CLK _83854_/Q _82534_/Q sky130_fd_sc_hd__dfxtp_4
X_55482_ _85106_/Q _55468_/X _55469_/X _55481_/Y _55482_/X sky130_fd_sc_hd__a211o_4
X_67468_ _67517_/A _67468_/B _67468_/X sky130_fd_sc_hd__and2_4
X_52694_ _52674_/X _52694_/B _52694_/C _52694_/D _52694_/X sky130_fd_sc_hd__and4_4
X_57221_ _57221_/A _85060_/Q _57221_/X sky130_fd_sc_hd__and2_4
X_69207_ _87534_/Q _69205_/X _69113_/X _69206_/X _69207_/X sky130_fd_sc_hd__a211o_4
X_88041_ _87789_/CLK _42087_/X _88041_/Q sky130_fd_sc_hd__dfxtp_4
X_54433_ _54446_/A _52739_/B _54433_/Y sky130_fd_sc_hd__nand2_4
X_66419_ _66003_/A _66419_/X sky130_fd_sc_hd__buf_2
X_85253_ _85221_/CLK _85253_/D _85253_/Q sky130_fd_sc_hd__dfxtp_4
X_51645_ _51629_/X _51651_/B _51651_/C _53170_/D _51645_/X sky130_fd_sc_hd__and4_4
X_82465_ _82443_/CLK _82465_/D _82465_/Q sky130_fd_sc_hd__dfxtp_4
X_67399_ _67324_/A _67399_/B _67399_/X sky130_fd_sc_hd__and2_4
X_84204_ _84194_/CLK _84204_/D _84204_/Q sky130_fd_sc_hd__dfxtp_4
X_81416_ _81703_/CLK _81448_/Q _75968_/B sky130_fd_sc_hd__dfxtp_4
X_57152_ _45909_/A _45672_/Y _57151_/Y _57152_/X sky130_fd_sc_hd__o21a_4
X_69138_ _69035_/A _69138_/X sky130_fd_sc_hd__buf_2
X_54364_ _54355_/A _54364_/B _54364_/Y sky130_fd_sc_hd__nand2_4
X_85184_ _85184_/CLK _56470_/Y _56469_/C sky130_fd_sc_hd__dfxtp_4
X_51576_ _51573_/Y _51557_/X _51575_/X _51576_/Y sky130_fd_sc_hd__a21oi_4
X_82396_ _82965_/CLK _82204_/Q _82396_/Q sky130_fd_sc_hd__dfxtp_4
X_56103_ _56102_/X _56103_/X sky130_fd_sc_hd__buf_2
X_53315_ _85656_/Q _53295_/X _53314_/Y _53315_/Y sky130_fd_sc_hd__o21ai_4
X_84135_ _82177_/CLK _84135_/D _84135_/Q sky130_fd_sc_hd__dfxtp_4
X_50527_ _50522_/Y _50525_/X _50526_/X _50527_/Y sky130_fd_sc_hd__a21oi_4
X_57083_ _56927_/A _56927_/C _57083_/X sky130_fd_sc_hd__and2_4
X_81347_ _84079_/CLK _76966_/Y _81347_/Q sky130_fd_sc_hd__dfxtp_4
X_69069_ _69958_/A _42534_/Y _69069_/Y sky130_fd_sc_hd__nor2_4
X_54295_ _54295_/A _54314_/A sky130_fd_sc_hd__buf_2
X_71100_ _50649_/B _71095_/X _71099_/Y _83608_/D sky130_fd_sc_hd__o21ai_4
X_56034_ _55956_/B _55956_/A _56035_/A sky130_fd_sc_hd__xnor2_4
X_41260_ _41259_/X _41251_/X _88249_/Q _41253_/X _88249_/D sky130_fd_sc_hd__a2bb2o_4
X_72080_ _72078_/Y _72033_/X _72079_/Y _83289_/D sky130_fd_sc_hd__a21boi_4
X_53246_ _53246_/A _53246_/B _53246_/Y sky130_fd_sc_hd__nand2_4
X_84066_ _81749_/CLK _84066_/D _81498_/D sky130_fd_sc_hd__dfxtp_4
X_50458_ _50439_/X _52163_/B _50458_/Y sky130_fd_sc_hd__nand2_4
X_81278_ _81269_/CLK _81310_/Q _81278_/Q sky130_fd_sc_hd__dfxtp_4
X_71031_ _53157_/B _71013_/X _71030_/Y _71031_/Y sky130_fd_sc_hd__o21ai_4
X_83017_ _86887_/CLK _74609_/Y _83017_/Q sky130_fd_sc_hd__dfxtp_4
X_80229_ _84950_/Q _65481_/C _80229_/Y sky130_fd_sc_hd__nand2_4
X_41191_ _41007_/A _40671_/A _41191_/X sky130_fd_sc_hd__or2_4
X_53177_ _53181_/A _53181_/B _53169_/X _53177_/D _53177_/X sky130_fd_sc_hd__and4_4
X_50389_ _50481_/A _50389_/B _50389_/Y sky130_fd_sc_hd__nand2_4
X_52128_ _52127_/X _52128_/B _52128_/Y sky130_fd_sc_hd__nand2_4
X_87825_ _88081_/CLK _42549_/Y _42548_/A sky130_fd_sc_hd__dfxtp_4
X_57985_ _57983_/X _85390_/Q _57984_/X _57985_/Y sky130_fd_sc_hd__o21ai_4
X_59724_ _59724_/A _59724_/Y sky130_fd_sc_hd__inv_2
X_44950_ _74547_/C _44933_/X _44949_/X _44950_/Y sky130_fd_sc_hd__o21ai_4
X_56936_ _72720_/A _72978_/A sky130_fd_sc_hd__buf_2
X_52059_ _52057_/Y _52022_/X _52058_/Y _52059_/Y sky130_fd_sc_hd__a21boi_4
X_75770_ _75768_/Y _75769_/Y _75771_/A sky130_fd_sc_hd__xor2_4
X_87756_ _88012_/CLK _42713_/X _68543_/B sky130_fd_sc_hd__dfxtp_4
X_72982_ _56547_/X _72982_/X sky130_fd_sc_hd__buf_2
X_84968_ _86530_/CLK _57620_/Y _84968_/Q sky130_fd_sc_hd__dfxtp_4
X_43901_ _43901_/A _43901_/Y sky130_fd_sc_hd__inv_2
X_74721_ _71266_/X _74775_/A sky130_fd_sc_hd__buf_2
X_86707_ _86384_/CLK _86707_/D _58751_/A sky130_fd_sc_hd__dfxtp_4
X_71933_ _74531_/A _70979_/C _71940_/C _71945_/D _71933_/Y sky130_fd_sc_hd__nand4_4
X_59655_ _59654_/X _59655_/X sky130_fd_sc_hd__buf_2
X_83919_ _83918_/CLK _83919_/D _81383_/D sky130_fd_sc_hd__dfxtp_4
X_44881_ _80670_/Q _45281_/A sky130_fd_sc_hd__buf_2
X_56867_ _56856_/Y _56884_/B _56721_/D _56867_/X sky130_fd_sc_hd__a21bo_4
X_87687_ _88133_/CLK _42851_/Y _66852_/B sky130_fd_sc_hd__dfxtp_4
X_84899_ _84727_/CLK _84899_/D _64283_/C sky130_fd_sc_hd__dfxtp_4
X_46620_ _46620_/A _46647_/B _46659_/C _52580_/D _46620_/X sky130_fd_sc_hd__and4_4
X_58606_ _58605_/X _85950_/Q _58568_/X _58606_/X sky130_fd_sc_hd__o21a_4
X_77440_ _77433_/Y _77439_/Y _82192_/D sky130_fd_sc_hd__xor2_4
X_43832_ _43752_/A _43832_/X sky130_fd_sc_hd__buf_2
X_55818_ _45196_/A _55492_/X _55312_/X _55817_/X _55818_/X sky130_fd_sc_hd__a211o_4
X_74652_ _74638_/X _56630_/A _45575_/A _74645_/X _82998_/D sky130_fd_sc_hd__a2bb2o_4
X_86638_ _86637_/CLK _47409_/Y _86638_/Q sky130_fd_sc_hd__dfxtp_4
X_71864_ _71847_/Y _83348_/Q _71863_/Y _83348_/D sky130_fd_sc_hd__a21o_4
X_59586_ _59662_/C _59657_/A _59615_/A _59775_/A _59586_/X sky130_fd_sc_hd__and4_4
X_56798_ _56798_/A _56798_/B _56798_/Y sky130_fd_sc_hd__nand2_4
X_73603_ _88369_/Q _73279_/X _73602_/X _73603_/X sky130_fd_sc_hd__o21a_4
X_70815_ _47174_/X _70802_/X _70814_/Y _70815_/Y sky130_fd_sc_hd__o21ai_4
X_46551_ _51372_/B _54071_/B sky130_fd_sc_hd__buf_2
X_58537_ _58448_/X _83361_/Q _58536_/Y _58537_/X sky130_fd_sc_hd__o21a_4
X_77371_ _77371_/A _77361_/Y _77371_/C _77371_/Y sky130_fd_sc_hd__nor3_4
X_43763_ _40964_/X _43752_/X _69206_/B _43753_/X _87278_/D sky130_fd_sc_hd__a2bb2o_4
X_55749_ _85256_/Q _55747_/X _55165_/X _55748_/X _55749_/X sky130_fd_sc_hd__a211o_4
X_74583_ _74552_/X _74583_/X sky130_fd_sc_hd__buf_2
X_86569_ _86535_/CLK _48089_/Y _74129_/B sky130_fd_sc_hd__dfxtp_4
X_40975_ _82297_/Q _40970_/B _40975_/X sky130_fd_sc_hd__or2_4
X_71795_ _58200_/Y _71784_/X _71794_/Y _71795_/Y sky130_fd_sc_hd__o21ai_4
X_79110_ _79110_/A _79110_/B _82625_/D sky130_fd_sc_hd__nand2_4
X_45502_ _45500_/Y _45439_/X _45471_/X _45501_/Y _45502_/X sky130_fd_sc_hd__a211o_4
X_76322_ _76305_/Y _76306_/A _76299_/Y _76322_/Y sky130_fd_sc_hd__a21boi_4
X_42714_ _41157_/X _42710_/X _87755_/Q _42711_/X _87755_/D sky130_fd_sc_hd__a2bb2o_4
X_88308_ _88324_/CLK _88308_/D _69972_/B sky130_fd_sc_hd__dfxtp_4
X_49270_ _86420_/Q _49255_/X _49269_/Y _49270_/Y sky130_fd_sc_hd__o21ai_4
X_73534_ _44600_/Y _73420_/X _73533_/Y _73534_/X sky130_fd_sc_hd__a21o_4
X_46482_ _48044_/B _47915_/B _46482_/Y sky130_fd_sc_hd__nand2_4
X_70746_ _53109_/B _70738_/X _70745_/Y _83711_/D sky130_fd_sc_hd__o21ai_4
X_58468_ _83417_/Q _58468_/Y sky130_fd_sc_hd__inv_2
X_43694_ _43693_/X _87305_/D sky130_fd_sc_hd__inv_2
X_48221_ _48221_/A _50275_/B sky130_fd_sc_hd__buf_2
X_79041_ _79048_/B _82524_/D _79042_/A sky130_fd_sc_hd__xor2_4
X_57419_ _57419_/A _57413_/X _57419_/X sky130_fd_sc_hd__or2_4
X_45433_ _44904_/A _45668_/A sky130_fd_sc_hd__buf_2
X_76253_ _76254_/A _76254_/B _76252_/Y _76253_/Y sky130_fd_sc_hd__a21oi_4
X_88239_ _87472_/CLK _41309_/X _67444_/B sky130_fd_sc_hd__dfxtp_4
X_42645_ _42614_/X _42615_/X _40972_/X _87788_/Q _42637_/X _42645_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73465_ _73465_/A _73228_/B _73465_/Y sky130_fd_sc_hd__nor2_4
X_70677_ _70664_/X _47468_/A _70676_/Y _83727_/D sky130_fd_sc_hd__a21o_4
X_58399_ _58399_/A _58400_/A sky130_fd_sc_hd__inv_2
X_75204_ _75207_/B _75201_/Y _75203_/Y _75205_/A sky130_fd_sc_hd__a21boi_4
X_48152_ _48152_/A _48153_/A sky130_fd_sc_hd__inv_2
X_60430_ _60447_/A _60430_/Y sky130_fd_sc_hd__inv_2
X_72416_ _86600_/Q _72428_/B _72416_/Y sky130_fd_sc_hd__nor2_4
X_45364_ _83011_/Q _45365_/A sky130_fd_sc_hd__inv_2
X_76184_ _81348_/Q _76183_/Y _76184_/X sky130_fd_sc_hd__xor2_4
X_42576_ _42576_/A _42576_/Y sky130_fd_sc_hd__inv_2
X_73396_ _87290_/Q _73003_/B _73396_/Y sky130_fd_sc_hd__nor2_4
X_47103_ _82382_/Q _47103_/Y sky130_fd_sc_hd__inv_2
X_44315_ _44315_/A _58007_/A sky130_fd_sc_hd__buf_2
X_75135_ _75120_/A _75116_/X _75134_/Y _75135_/Y sky130_fd_sc_hd__a21oi_4
X_41527_ _41358_/X _82323_/Q _41527_/X sky130_fd_sc_hd__or2_4
X_60361_ _60360_/X _60362_/A sky130_fd_sc_hd__buf_2
X_72347_ _72347_/A _72347_/B _72347_/Y sky130_fd_sc_hd__nor2_4
X_48083_ _48092_/A _48310_/B _48083_/Y sky130_fd_sc_hd__nand2_4
X_45295_ _45277_/X _61627_/B _45294_/X _45295_/Y sky130_fd_sc_hd__o21ai_4
X_62100_ _62093_/X _62095_/X _62099_/Y _58344_/A _62048_/X _62100_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47034_ _86677_/Q _47004_/X _47033_/Y _47034_/Y sky130_fd_sc_hd__o21ai_4
X_44246_ _44246_/A _58631_/A sky130_fd_sc_hd__buf_2
X_79943_ _79940_/Y _79941_/Y _79942_/A _79945_/A sky130_fd_sc_hd__a21o_4
X_63080_ _63074_/Y _63075_/X _63077_/X _63079_/X _63067_/X _63080_/Y
+ sky130_fd_sc_hd__o41ai_4
X_75066_ _80960_/Q _75066_/B _75066_/X sky130_fd_sc_hd__xor2_4
X_41458_ _41454_/X _41455_/X _88212_/Q _41457_/X _88212_/D sky130_fd_sc_hd__a2bb2o_4
X_60292_ _60292_/A _60337_/A sky130_fd_sc_hd__buf_2
X_72278_ _86612_/Q _72348_/B _72278_/Y sky130_fd_sc_hd__nor2_4
X_62031_ _62021_/X _62023_/X _62030_/Y _84846_/Q _61973_/X _62031_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74017_ _73972_/X _66183_/B _74017_/X sky130_fd_sc_hd__and2_4
X_40409_ _47363_/A _40409_/X sky130_fd_sc_hd__buf_2
X_71229_ _48673_/B _71216_/X _71228_/Y _71229_/Y sky130_fd_sc_hd__o21ai_4
X_44177_ _58126_/A _44177_/X sky130_fd_sc_hd__buf_2
X_79874_ _79870_/Y _79873_/Y _79874_/X sky130_fd_sc_hd__xor2_4
X_41389_ _41337_/X _41338_/X _41387_/X _67801_/B _41388_/X _41389_/Y
+ sky130_fd_sc_hd__o32ai_4
X_43128_ _43046_/X _43125_/X _40792_/X _43126_/Y _43127_/X _87566_/D
+ sky130_fd_sc_hd__o32ai_4
X_78825_ _78825_/A _82836_/Q _78828_/C sky130_fd_sc_hd__nand2_4
X_48985_ _48985_/A _48985_/X sky130_fd_sc_hd__buf_2
X_47936_ _47904_/X _82936_/Q _47935_/X _47937_/B sky130_fd_sc_hd__o21ai_4
X_43059_ _43053_/X _43054_/X _40650_/X _43057_/Y _43058_/X _87592_/D
+ sky130_fd_sc_hd__o32ai_4
X_66770_ _87127_/Q _66715_/X _66717_/X _66769_/X _66770_/X sky130_fd_sc_hd__a211o_4
X_78756_ _78755_/X _78756_/Y sky130_fd_sc_hd__inv_2
X_63982_ _63724_/A _64046_/B sky130_fd_sc_hd__buf_2
X_75968_ _81704_/D _75968_/B _75969_/B sky130_fd_sc_hd__nand2_4
X_65721_ _65716_/X _65720_/X _65566_/X _65721_/X sky130_fd_sc_hd__a21o_4
X_77707_ _77707_/A _82208_/D sky130_fd_sc_hd__inv_2
X_62933_ _62971_/A _84888_/Q _62819_/C _62979_/D _62933_/X sky130_fd_sc_hd__and4_4
X_74919_ _74912_/X _74930_/A _74920_/B sky130_fd_sc_hd__xor2_4
X_47867_ _47867_/A _47867_/X sky130_fd_sc_hd__buf_2
X_78687_ _78701_/A _78686_/Y _82779_/D sky130_fd_sc_hd__xnor2_4
X_75899_ _75899_/A _84369_/Q _75899_/X sky130_fd_sc_hd__xor2_4
X_49606_ _49632_/A _49606_/X sky130_fd_sc_hd__buf_2
X_68440_ _66053_/A _68440_/B _68440_/Y sky130_fd_sc_hd__nor2_4
X_46818_ _86700_/Q _46813_/X _46817_/Y _46818_/Y sky130_fd_sc_hd__o21ai_4
X_65652_ _65648_/Y _65602_/X _65651_/Y _84187_/D sky130_fd_sc_hd__a21o_4
X_77638_ _77666_/B _77638_/Y sky130_fd_sc_hd__inv_2
X_62864_ _62894_/A _62852_/X _62864_/C _62864_/Y sky130_fd_sc_hd__nor3_4
X_47798_ _47798_/A _51728_/B sky130_fd_sc_hd__buf_2
X_64603_ _64684_/A _86465_/Q _64603_/X sky130_fd_sc_hd__and2_4
X_49537_ _49537_/A _49537_/B _49522_/C _52750_/D _49537_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_441_0_CLK clkbuf_9_220_0_CLK/X _84150_/CLK sky130_fd_sc_hd__clkbuf_1
X_61815_ _61719_/A _61815_/X sky130_fd_sc_hd__buf_2
X_68371_ _68371_/A _88371_/Q _68371_/X sky130_fd_sc_hd__and2_4
X_46749_ _46733_/A _50961_/B _46749_/Y sky130_fd_sc_hd__nand2_4
X_65583_ _65782_/A _65769_/A sky130_fd_sc_hd__buf_2
X_77569_ _77568_/Y _77570_/C sky130_fd_sc_hd__inv_2
X_62795_ _62790_/X _62779_/X _62794_/Y _84382_/D sky130_fd_sc_hd__a21oi_4
X_67322_ _67203_/X _67322_/X sky130_fd_sc_hd__buf_2
X_79308_ _79302_/A _79301_/X _79307_/Y _79324_/A sky130_fd_sc_hd__a21boi_4
X_64534_ _64234_/A _64234_/B _64534_/C _64221_/X _64534_/X sky130_fd_sc_hd__and4_4
X_49468_ _49465_/Y _49460_/X _49467_/X _86382_/D sky130_fd_sc_hd__a21oi_4
X_61746_ _61966_/A _61765_/C sky130_fd_sc_hd__buf_2
X_80580_ _80580_/A _80580_/B _80596_/B sky130_fd_sc_hd__xnor2_4
X_48419_ _48478_/A _48419_/X sky130_fd_sc_hd__buf_2
X_79239_ _79239_/A _79240_/B sky130_fd_sc_hd__inv_2
X_67253_ _67183_/A _88183_/Q _67253_/X sky130_fd_sc_hd__and2_4
X_64465_ _63630_/A _64419_/B _64465_/Y sky130_fd_sc_hd__nor2_4
X_49399_ _49410_/A _46685_/X _49399_/Y sky130_fd_sc_hd__nand2_4
X_61677_ _58364_/A _61598_/X _61677_/C _72563_/B _61678_/A sky130_fd_sc_hd__nand4_4
Xclkbuf_10_456_0_CLK clkbuf_9_228_0_CLK/X _83275_/CLK sky130_fd_sc_hd__clkbuf_1
X_66204_ _66204_/A _66203_/Y _66204_/Y sky130_fd_sc_hd__nand2_4
X_51430_ _51211_/A _51430_/X sky130_fd_sc_hd__buf_2
X_63416_ _63416_/A _63465_/B sky130_fd_sc_hd__buf_2
X_82250_ _82253_/CLK _80387_/X _82250_/Q sky130_fd_sc_hd__dfxtp_4
X_60628_ _60628_/A _59552_/C _60628_/C _60628_/Y sky130_fd_sc_hd__nand3_4
X_67184_ _88378_/Q _67110_/X _67160_/X _67183_/X _67184_/X sky130_fd_sc_hd__a211o_4
X_64396_ _64390_/X _64392_/X _64393_/X _64395_/Y _64384_/X _64396_/X
+ sky130_fd_sc_hd__o41a_4
X_81201_ _84981_/CLK _75007_/X _49049_/A sky130_fd_sc_hd__dfxtp_4
X_66135_ _65659_/X _66135_/B _65662_/X _66135_/Y sky130_fd_sc_hd__nand3_4
X_51361_ _51359_/Y _51339_/X _51360_/X _86025_/D sky130_fd_sc_hd__a21oi_4
X_63347_ _60562_/B _61692_/B _63347_/C _60570_/A _63347_/X sky130_fd_sc_hd__and4_4
X_82181_ _84951_/CLK _77276_/Y _82181_/Q sky130_fd_sc_hd__dfxtp_4
X_60559_ _60558_/X _60612_/A sky130_fd_sc_hd__buf_2
X_53100_ _53096_/Y _53082_/X _53099_/X _85698_/D sky130_fd_sc_hd__a21oi_4
X_50312_ _50473_/A _50491_/A sky130_fd_sc_hd__buf_2
X_81132_ _80804_/CLK _81132_/D _40705_/A sky130_fd_sc_hd__dfxtp_4
X_54080_ _54078_/Y _54060_/X _54079_/Y _54080_/Y sky130_fd_sc_hd__a21boi_4
X_66066_ _65970_/A _66004_/B _84159_/Q _66066_/X sky130_fd_sc_hd__and3_4
X_51292_ _51296_/A _50781_/B _51292_/Y sky130_fd_sc_hd__nand2_4
X_63278_ _58970_/A _62999_/X _61617_/B _60608_/X _63278_/Y sky130_fd_sc_hd__a2bb2oi_4
X_53031_ _53048_/A _53036_/B _53019_/C _53031_/D _53031_/X sky130_fd_sc_hd__and4_4
X_65017_ _64835_/X _83298_/Q _65015_/X _65016_/X _65017_/X sky130_fd_sc_hd__a211o_4
X_50243_ _50768_/A _50243_/X sky130_fd_sc_hd__buf_2
X_62229_ _62632_/A _63369_/B _62319_/C _62229_/Y sky130_fd_sc_hd__nand3_4
X_85940_ _86100_/CLK _51825_/Y _85940_/Q sky130_fd_sc_hd__dfxtp_4
X_81063_ _81061_/CLK _81095_/Q _81063_/Q sky130_fd_sc_hd__dfxtp_4
X_80014_ _80008_/X _80013_/Y _81674_/D sky130_fd_sc_hd__xor2_4
Xclkbuf_9_500_0_CLK clkbuf_9_501_0_CLK/A clkbuf_9_500_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_69825_ _69822_/X _69824_/X _66579_/X _69825_/X sky130_fd_sc_hd__a21o_4
X_50174_ _86249_/Q _50162_/X _50173_/Y _50174_/Y sky130_fd_sc_hd__o21ai_4
X_85871_ _86500_/CLK _85871_/D _85871_/Q sky130_fd_sc_hd__dfxtp_4
X_87610_ _82899_/CLK _87610_/D _87610_/Q sky130_fd_sc_hd__dfxtp_4
X_84822_ _84869_/CLK _58549_/Y _58546_/A sky130_fd_sc_hd__dfxtp_4
X_57770_ _57770_/A _58796_/A sky130_fd_sc_hd__buf_2
X_69756_ _69770_/A _69756_/B _69756_/X sky130_fd_sc_hd__and2_4
X_54982_ _85341_/Q _54967_/X _54981_/Y _54982_/Y sky130_fd_sc_hd__o21ai_4
X_66968_ _66965_/X _66967_/X _66658_/X _66968_/Y sky130_fd_sc_hd__a21oi_4
X_56721_ _56721_/A _56651_/Y _56655_/Y _56721_/D _56721_/Y sky130_fd_sc_hd__nor4_4
X_68707_ _68059_/A _68707_/X sky130_fd_sc_hd__buf_2
X_87541_ _88085_/CLK _87541_/D _43201_/A sky130_fd_sc_hd__dfxtp_4
X_53933_ _85539_/Q _53921_/X _53932_/Y _53933_/Y sky130_fd_sc_hd__o21ai_4
X_65919_ _65763_/A _73583_/B _65919_/X sky130_fd_sc_hd__and2_4
X_84753_ _84760_/CLK _59303_/Y _84753_/Q sky130_fd_sc_hd__dfxtp_4
X_81965_ _82299_/CLK _83893_/Q _81965_/Q sky130_fd_sc_hd__dfxtp_4
X_69687_ _69687_/A _42564_/Y _69687_/Y sky130_fd_sc_hd__nor2_4
X_66899_ _66898_/X _66899_/X sky130_fd_sc_hd__buf_2
X_83704_ _85428_/CLK _70770_/Y _47077_/A sky130_fd_sc_hd__dfxtp_4
X_59440_ _59439_/Y _59424_/B _59440_/Y sky130_fd_sc_hd__nand2_4
X_80916_ _81507_/CLK _80916_/D _75732_/A sky130_fd_sc_hd__dfxtp_4
X_56652_ _83325_/Q _83324_/Q _57131_/A sky130_fd_sc_hd__nand2_4
X_87472_ _87472_/CLK _87472_/D _87472_/Q sky130_fd_sc_hd__dfxtp_4
X_68638_ _69086_/A _73822_/A _68638_/X sky130_fd_sc_hd__and2_4
X_53864_ _53861_/Y _53862_/X _53863_/Y _53864_/Y sky130_fd_sc_hd__a21boi_4
X_84684_ _84329_/CLK _59869_/Y _80294_/B sky130_fd_sc_hd__dfxtp_4
X_81896_ _82139_/CLK _77322_/X _77222_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_409_0_CLK clkbuf_9_204_0_CLK/X _83514_/CLK sky130_fd_sc_hd__clkbuf_1
X_55603_ _55570_/X _72648_/C _72643_/C _72641_/C _55603_/X sky130_fd_sc_hd__and4_4
X_86423_ _86422_/CLK _49260_/Y _86423_/Q sky130_fd_sc_hd__dfxtp_4
X_52815_ _49793_/A _53221_/A sky130_fd_sc_hd__buf_2
X_59371_ _59367_/Y _59370_/Y _59297_/X _59371_/X sky130_fd_sc_hd__a21o_4
X_83635_ _86122_/CLK _71007_/Y _83635_/Q sky130_fd_sc_hd__dfxtp_4
X_56583_ _72643_/C _56583_/B _56583_/X sky130_fd_sc_hd__xor2_4
X_80847_ _81130_/CLK _80847_/D _74945_/B sky130_fd_sc_hd__dfxtp_4
X_68569_ _68566_/X _68568_/X _68442_/X _68574_/A sky130_fd_sc_hd__a21o_4
X_53795_ _53792_/Y _53696_/X _53794_/Y _85567_/D sky130_fd_sc_hd__a21boi_4
Xclkbuf_7_0_0_CLK clkbuf_6_0_0_CLK/X clkbuf_8_1_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_70600_ _52973_/B _70584_/X _70599_/Y _83744_/D sky130_fd_sc_hd__o21ai_4
X_58322_ _58322_/A _58322_/Y sky130_fd_sc_hd__inv_2
X_55534_ _55534_/A _56627_/B _55534_/X sky130_fd_sc_hd__and2_4
X_86354_ _86353_/CLK _86354_/D _86354_/Q sky130_fd_sc_hd__dfxtp_4
X_40760_ _40760_/A _40760_/B _40760_/X sky130_fd_sc_hd__or2_4
X_52746_ _52729_/X _52746_/B _52746_/C _52746_/D _52746_/X sky130_fd_sc_hd__and4_4
X_71580_ _71580_/A _71581_/A sky130_fd_sc_hd__inv_2
X_83566_ _83311_/CLK _71227_/Y _48659_/A sky130_fd_sc_hd__dfxtp_4
X_80778_ _80849_/CLK _75662_/Y _80778_/Q sky130_fd_sc_hd__dfxtp_4
X_85305_ _85241_/CLK _85305_/D _55913_/B sky130_fd_sc_hd__dfxtp_4
X_70531_ _71507_/A _70530_/Y _70361_/A _70531_/Y sky130_fd_sc_hd__nor3_4
X_82517_ _82532_/CLK _82517_/D _82517_/Q sky130_fd_sc_hd__dfxtp_4
X_58253_ _58253_/A _58253_/X sky130_fd_sc_hd__buf_2
X_55465_ _45604_/A _55462_/X _44096_/X _55464_/X _55465_/X sky130_fd_sc_hd__a211o_4
X_86285_ _86282_/CLK _86285_/D _72366_/B sky130_fd_sc_hd__dfxtp_4
X_40691_ _40691_/A _40691_/X sky130_fd_sc_hd__buf_2
X_52677_ _52657_/X _52677_/B _52677_/Y sky130_fd_sc_hd__nand2_4
X_83497_ _84939_/CLK _71443_/Y _83497_/Q sky130_fd_sc_hd__dfxtp_4
X_57204_ _56857_/X _57129_/A _56863_/X _57198_/B _57204_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_8_83_0_CLK clkbuf_8_83_0_CLK/A clkbuf_8_83_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_88024_ _87249_/CLK _88024_/D _88024_/Q sky130_fd_sc_hd__dfxtp_4
X_42430_ _42574_/A _42430_/X sky130_fd_sc_hd__buf_2
X_54416_ _85446_/Q _54404_/X _54415_/Y _54416_/Y sky130_fd_sc_hd__o21ai_4
X_73250_ _73250_/A _73250_/X sky130_fd_sc_hd__buf_2
X_85236_ _86900_/CLK _85236_/D _55865_/B sky130_fd_sc_hd__dfxtp_4
X_51628_ _85975_/Q _51621_/X _51627_/Y _51628_/Y sky130_fd_sc_hd__o21ai_4
X_70462_ _71483_/B _71500_/C sky130_fd_sc_hd__buf_2
X_58184_ _58184_/A _58184_/B _58184_/Y sky130_fd_sc_hd__nor2_4
X_82448_ _82828_/CLK _79140_/X _82448_/Q sky130_fd_sc_hd__dfxtp_4
X_55396_ _55373_/Y _55396_/B _55409_/A sky130_fd_sc_hd__nand2_4
X_72201_ _72201_/A _72201_/X sky130_fd_sc_hd__buf_2
X_57135_ _57134_/Y _56685_/X _57135_/Y sky130_fd_sc_hd__nor2_4
X_42361_ _41741_/X _42356_/X _87902_/Q _42357_/X _87902_/D sky130_fd_sc_hd__a2bb2o_4
X_54347_ _54362_/A _54353_/B _54362_/C _46753_/Y _54347_/X sky130_fd_sc_hd__and4_4
X_73181_ _73181_/A _85873_/Q _73181_/X sky130_fd_sc_hd__and2_4
X_85167_ _85167_/CLK _56514_/Y _55823_/B sky130_fd_sc_hd__dfxtp_4
X_51559_ _51553_/A _51580_/B _51553_/C _53084_/D _51559_/X sky130_fd_sc_hd__and4_4
X_82379_ _86054_/CLK _82187_/Q _82379_/Q sky130_fd_sc_hd__dfxtp_4
X_70393_ DATA_TO_HASH[2] _70819_/A sky130_fd_sc_hd__buf_2
X_44100_ _44099_/X _44101_/A sky130_fd_sc_hd__buf_2
X_41312_ _41311_/Y _41312_/X sky130_fd_sc_hd__buf_2
X_72132_ _59331_/X _85376_/Q _72131_/X _72132_/Y sky130_fd_sc_hd__o21ai_4
X_84118_ _84166_/CLK _84118_/D _84118_/Q sky130_fd_sc_hd__dfxtp_4
X_45080_ _55889_/B _45044_/X _45079_/X _45080_/X sky130_fd_sc_hd__o21a_4
X_57066_ _56912_/A _57289_/B sky130_fd_sc_hd__buf_2
X_42292_ _41556_/X _42290_/X _87937_/Q _42291_/X _42292_/X sky130_fd_sc_hd__a2bb2o_4
X_54278_ _85471_/Q _54266_/X _54277_/Y _54278_/Y sky130_fd_sc_hd__o21ai_4
X_85098_ _85031_/CLK _85098_/D _85098_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_98_0_CLK clkbuf_8_99_0_CLK/A clkbuf_8_98_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_44031_ _72255_/A _44031_/X sky130_fd_sc_hd__buf_2
X_56017_ _56177_/A _56017_/B _85311_/Q _56017_/Y sky130_fd_sc_hd__nand3_4
X_41243_ _41068_/B _41223_/B _41243_/X sky130_fd_sc_hd__or2_4
X_53229_ _53282_/A _53244_/B sky130_fd_sc_hd__buf_2
X_72063_ _83292_/Q _72001_/X _72062_/Y _72063_/Y sky130_fd_sc_hd__o21ai_4
X_76940_ _76938_/B _76939_/A _76953_/A sky130_fd_sc_hd__nand2_4
X_84049_ _84049_/CLK _84049_/D _81481_/D sky130_fd_sc_hd__dfxtp_4
X_71014_ _70763_/A _71168_/A sky130_fd_sc_hd__buf_2
X_41174_ _41173_/X _41174_/X sky130_fd_sc_hd__buf_2
X_76871_ _76910_/A _76870_/Y _81466_/D sky130_fd_sc_hd__xor2_4
X_78610_ _78596_/Y _78608_/Y _78609_/Y _78610_/X sky130_fd_sc_hd__o21a_4
X_75822_ _75811_/A _75815_/Y _75823_/C _75824_/A sky130_fd_sc_hd__a21o_4
Xclkbuf_8_21_0_CLK clkbuf_8_21_0_CLK/A clkbuf_9_43_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_87808_ _87814_/CLK _42596_/Y _87808_/Q sky130_fd_sc_hd__dfxtp_4
X_48770_ _52573_/B _48770_/X sky130_fd_sc_hd__buf_2
X_79590_ _79572_/Y _79590_/Y sky130_fd_sc_hd__inv_2
X_45982_ _45981_/X _45982_/X sky130_fd_sc_hd__buf_2
X_57968_ _57939_/X _86000_/Q _57967_/X _57968_/Y sky130_fd_sc_hd__o21ai_4
X_47721_ _81229_/Q _47722_/A sky130_fd_sc_hd__inv_2
X_59707_ _63001_/A _63344_/B sky130_fd_sc_hd__buf_2
X_78541_ _78528_/A _78528_/B _78521_/X _78541_/Y sky130_fd_sc_hd__a21boi_4
X_44933_ _45252_/A _44933_/X sky130_fd_sc_hd__buf_2
X_56919_ _56636_/X _59498_/A _57193_/D _56921_/B sky130_fd_sc_hd__nand3_4
X_75753_ _75752_/X _75753_/Y sky130_fd_sc_hd__inv_2
X_87739_ _87487_/CLK _42752_/Y _87739_/Q sky130_fd_sc_hd__dfxtp_4
X_72965_ _72963_/X _83074_/Q _72785_/X _72964_/X _72965_/X sky130_fd_sc_hd__a211o_4
X_57899_ _58098_/A _57899_/X sky130_fd_sc_hd__buf_2
X_74704_ _74704_/A _74704_/Y sky130_fd_sc_hd__inv_2
X_47652_ _47792_/A _47692_/B sky130_fd_sc_hd__buf_2
X_71916_ _70554_/A _71386_/B _71916_/Y sky130_fd_sc_hd__nor2_4
X_59638_ _59638_/A _59651_/A sky130_fd_sc_hd__inv_2
X_78472_ _78472_/A _82670_/D _78472_/X sky130_fd_sc_hd__xor2_4
X_44864_ _44863_/Y _86913_/D sky130_fd_sc_hd__inv_2
X_75684_ _75684_/A _75684_/B _75684_/Y sky130_fd_sc_hd__nand2_4
X_72896_ _87310_/Q _72896_/B _72896_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_8_36_0_CLK clkbuf_8_37_0_CLK/A clkbuf_9_72_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_46603_ _53874_/A _46603_/X sky130_fd_sc_hd__buf_2
X_77423_ _77423_/A _82096_/D _77423_/Y sky130_fd_sc_hd__nor2_4
X_43815_ _41098_/X _43801_/X _87254_/Q _43802_/X _43815_/X sky130_fd_sc_hd__a2bb2o_4
X_74635_ _45952_/X _56574_/Y _83007_/Q _74633_/X _83007_/D sky130_fd_sc_hd__a2bb2o_4
X_47583_ _47574_/A _53131_/B _47583_/Y sky130_fd_sc_hd__nand2_4
X_71847_ _71846_/Y _71847_/Y sky130_fd_sc_hd__inv_2
X_59569_ _59568_/X _59570_/A sky130_fd_sc_hd__buf_2
X_44795_ _41415_/Y _44788_/X _86951_/Q _44789_/X _86951_/D sky130_fd_sc_hd__a2bb2o_4
X_49322_ _49273_/A _49322_/B _49322_/Y sky130_fd_sc_hd__nand2_4
X_61600_ _58461_/A _61598_/X _61677_/C _61563_/D _61600_/Y sky130_fd_sc_hd__nand4_4
X_46534_ _52545_/B _50852_/B sky130_fd_sc_hd__buf_2
X_77354_ _77354_/A _77354_/B _77354_/X sky130_fd_sc_hd__or2_4
X_43746_ _43745_/X _87287_/D sky130_fd_sc_hd__inv_2
X_74566_ _74559_/X _74553_/X _56055_/A _74554_/X _74566_/X sky130_fd_sc_hd__a211o_4
X_62580_ _61637_/X _62560_/B _62560_/C _62560_/D _62580_/Y sky130_fd_sc_hd__nand4_4
X_40958_ _40512_/X _81725_/Q _40957_/X _40959_/A sky130_fd_sc_hd__o21a_4
X_71778_ _71761_/Y _83379_/Q _71777_/X _83379_/D sky130_fd_sc_hd__a21o_4
X_76305_ _76301_/Y _76303_/Y _76300_/Y _76305_/Y sky130_fd_sc_hd__o21ai_4
X_49253_ _49263_/A _52468_/B _49253_/Y sky130_fd_sc_hd__nand2_4
X_61531_ _58434_/A _61563_/B _61563_/C _61514_/D _61532_/A sky130_fd_sc_hd__nand4_4
X_73517_ _73355_/X _85571_/Q _73472_/X _73516_/X _73517_/X sky130_fd_sc_hd__a211o_4
X_46465_ _46464_/Y _51328_/B sky130_fd_sc_hd__buf_2
X_70729_ _70668_/D _71266_/A sky130_fd_sc_hd__buf_2
X_77285_ _77285_/A _77280_/X _77285_/C _77286_/A sky130_fd_sc_hd__nand3_4
X_43677_ _43677_/A _43677_/Y sky130_fd_sc_hd__inv_2
X_74497_ _48666_/A _74501_/B _74501_/C _74497_/X sky130_fd_sc_hd__and3_4
X_40889_ _40585_/X _82282_/Q _40888_/X _40889_/Y sky130_fd_sc_hd__o21ai_4
X_48204_ _48171_/X _48204_/X sky130_fd_sc_hd__buf_2
X_79024_ _79012_/Y _79014_/B _82648_/Q _82520_/D _79024_/X sky130_fd_sc_hd__a2bb2o_4
X_45416_ _45416_/A _44894_/B _45416_/Y sky130_fd_sc_hd__nor2_4
X_64250_ _64250_/A _84854_/Q _64250_/C _64250_/Y sky130_fd_sc_hd__nand3_4
X_76236_ _76231_/Y _76233_/Y _76235_/Y _76236_/X sky130_fd_sc_hd__a21o_4
X_42628_ _52274_/A _42743_/A sky130_fd_sc_hd__inv_2
X_61462_ _61400_/X _61482_/C sky130_fd_sc_hd__buf_2
X_73448_ _73378_/X _86182_/Q _73446_/X _73447_/X _73448_/X sky130_fd_sc_hd__a211o_4
X_49184_ _49184_/A _53932_/B sky130_fd_sc_hd__inv_2
X_46396_ _46387_/A _46396_/B _46396_/Y sky130_fd_sc_hd__nand2_4
X_63201_ _58380_/A _63190_/X _63175_/X _58254_/Y _63176_/X _63201_/Y
+ sky130_fd_sc_hd__o32ai_4
X_60413_ _60412_/X _60413_/X sky130_fd_sc_hd__buf_2
X_48135_ _48135_/A _48136_/B sky130_fd_sc_hd__buf_2
X_45347_ _45347_/A _45381_/B _45347_/Y sky130_fd_sc_hd__nand2_4
X_64181_ _64181_/A _64181_/B _64181_/C _64181_/D _64181_/X sky130_fd_sc_hd__and4_4
X_76167_ _76160_/X _76165_/X _76161_/Y _76168_/B sky130_fd_sc_hd__nand3_4
X_42559_ _42554_/X _42547_/X _40798_/X _42558_/Y _42556_/X _42559_/Y
+ sky130_fd_sc_hd__o32ai_4
X_61393_ _61386_/Y _61388_/Y _61334_/X _61390_/Y _61392_/Y _61393_/X
+ sky130_fd_sc_hd__a41o_4
X_73379_ _73495_/A _85865_/Q _73379_/X sky130_fd_sc_hd__and2_4
X_63132_ _58546_/Y _63131_/X _63117_/X _58322_/Y _63118_/X _63132_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75118_ _75107_/A _75106_/A _75105_/A _75120_/A sky130_fd_sc_hd__o21ai_4
X_48066_ _47867_/X _82923_/Q _48065_/Y _48067_/A sky130_fd_sc_hd__o21ai_4
X_60344_ _60344_/A _60344_/B _60344_/C _60344_/Y sky130_fd_sc_hd__nand3_4
X_45278_ _62557_/A _61617_/B sky130_fd_sc_hd__buf_2
X_76098_ _76081_/Y _76095_/X _76097_/Y _76099_/B sky130_fd_sc_hd__a21oi_4
X_47017_ _47008_/A _52803_/B _47017_/Y sky130_fd_sc_hd__nand2_4
X_44229_ _44228_/X _56995_/A sky130_fd_sc_hd__buf_2
X_67940_ _87450_/Q _67868_/X _67938_/X _67939_/X _67940_/X sky130_fd_sc_hd__a211o_4
X_63063_ _63038_/A _64275_/B _63085_/C _63085_/D _63063_/X sky130_fd_sc_hd__and4_4
X_75049_ _75049_/A _75048_/Y _75051_/A sky130_fd_sc_hd__or2_4
X_79926_ _79926_/A _79918_/Y _79919_/Y _79927_/B sky130_fd_sc_hd__nand3_4
X_60275_ _60189_/Y _60274_/X _60253_/A _60275_/X sky130_fd_sc_hd__and3_4
X_62014_ _63585_/B _61999_/B _61971_/C _61971_/D _62015_/D sky130_fd_sc_hd__nand4_4
X_67871_ _67867_/X _67870_/X _67799_/X _67871_/X sky130_fd_sc_hd__a21o_4
X_79857_ _79856_/X _79857_/Y sky130_fd_sc_hd__inv_2
X_69610_ _69606_/X _69609_/X _69385_/X _69610_/X sky130_fd_sc_hd__a21o_4
X_66822_ _68474_/A _66823_/A sky130_fd_sc_hd__buf_2
X_78808_ _82834_/Q _78809_/A sky130_fd_sc_hd__inv_2
X_48968_ _48946_/X _48449_/A _48967_/Y _48969_/A sky130_fd_sc_hd__a21o_4
X_79788_ _79777_/X _79766_/X _79788_/X sky130_fd_sc_hd__and2_4
X_69541_ _81380_/D _69504_/X _69540_/X _83916_/D sky130_fd_sc_hd__a21bo_4
X_47919_ _48790_/A _47919_/X sky130_fd_sc_hd__buf_2
X_78739_ _78739_/A _78747_/A sky130_fd_sc_hd__inv_2
X_66753_ _87128_/Q _66751_/X _66682_/X _66752_/X _66753_/X sky130_fd_sc_hd__a211o_4
X_63965_ _63964_/Y _63965_/Y sky130_fd_sc_hd__inv_2
X_48899_ _83623_/Q _48899_/Y sky130_fd_sc_hd__inv_2
X_65704_ _65704_/A _86479_/Q _65704_/X sky130_fd_sc_hd__and2_4
X_50930_ _50941_/A _50941_/B _50948_/C _52622_/D _50930_/X sky130_fd_sc_hd__and4_4
X_62916_ _62916_/A _62916_/Y sky130_fd_sc_hd__inv_2
X_81750_ _81514_/CLK _76069_/B _81750_/Q sky130_fd_sc_hd__dfxtp_4
X_69472_ _69309_/A _69472_/B _69472_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_380_0_CLK clkbuf_9_190_0_CLK/X _85436_/CLK sky130_fd_sc_hd__clkbuf_1
X_66684_ _88399_/Q _66633_/X _66682_/X _66683_/X _66684_/X sky130_fd_sc_hd__a211o_4
X_63896_ _63889_/X _63890_/X _63892_/Y _63894_/Y _63895_/X _63896_/X
+ sky130_fd_sc_hd__a41o_4
X_80701_ _84276_/CLK _80733_/Q _75475_/A sky130_fd_sc_hd__dfxtp_4
X_68423_ _87005_/Q _68394_/X _68421_/X _68422_/X _68423_/X sky130_fd_sc_hd__a211o_4
X_65635_ _65632_/Y _65602_/X _65634_/Y _84188_/D sky130_fd_sc_hd__a21o_4
X_50861_ _50859_/Y _50849_/X _50860_/Y _86119_/D sky130_fd_sc_hd__a21boi_4
X_62847_ _62847_/A _62847_/X sky130_fd_sc_hd__buf_2
X_81681_ _81684_/CLK _81681_/D _81681_/Q sky130_fd_sc_hd__dfxtp_4
X_52600_ _52597_/Y _52592_/X _52599_/X _52600_/Y sky130_fd_sc_hd__a21oi_4
X_83420_ _83421_/CLK _83420_/D _58522_/A sky130_fd_sc_hd__dfxtp_4
X_80632_ _80632_/A _80632_/B _80632_/Y sky130_fd_sc_hd__nand2_4
X_68354_ _64980_/A _68354_/X sky130_fd_sc_hd__buf_2
X_53580_ _53578_/Y _53574_/X _53579_/Y _85609_/D sky130_fd_sc_hd__a21boi_4
X_65566_ _64807_/A _65566_/X sky130_fd_sc_hd__buf_2
X_50792_ _50768_/A _50792_/X sky130_fd_sc_hd__buf_2
X_62778_ _62771_/Y _62772_/X _62774_/Y _62775_/Y _62777_/X _62778_/X
+ sky130_fd_sc_hd__a41o_4
X_67305_ _64608_/A _67305_/X sky130_fd_sc_hd__buf_2
X_52531_ _85803_/Q _52516_/X _52530_/Y _52531_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_395_0_CLK clkbuf_9_197_0_CLK/X _82452_/CLK sky130_fd_sc_hd__clkbuf_1
X_64517_ _64512_/X _64513_/X _64514_/X _64516_/Y _64440_/X _64517_/X
+ sky130_fd_sc_hd__o41a_4
X_83351_ _83480_/CLK _83351_/D _83351_/Q sky130_fd_sc_hd__dfxtp_4
X_61729_ _59766_/X _62183_/D sky130_fd_sc_hd__buf_2
X_80563_ _80550_/A _80549_/Y _80562_/Y _80564_/B sky130_fd_sc_hd__o21a_4
X_68285_ _68254_/X _67746_/Y _68268_/X _68284_/Y _68285_/X sky130_fd_sc_hd__a211o_4
X_65497_ _84197_/Q _65498_/C sky130_fd_sc_hd__inv_2
XPHY_108 sky130_fd_sc_hd__decap_3
XPHY_119 sky130_fd_sc_hd__decap_3
X_82302_ _82343_/CLK _82302_/D _82302_/Q sky130_fd_sc_hd__dfxtp_4
X_55250_ _55247_/X _55249_/X _55138_/X _55254_/A sky130_fd_sc_hd__a21o_4
X_67236_ _66758_/X _67236_/X sky130_fd_sc_hd__buf_2
X_86070_ _85751_/CLK _51122_/Y _86070_/Q sky130_fd_sc_hd__dfxtp_4
X_52462_ _52462_/A _52462_/X sky130_fd_sc_hd__buf_2
X_64448_ _64402_/X _64421_/X _84837_/Q _64448_/X sky130_fd_sc_hd__and3_4
X_83282_ _83282_/CLK _72114_/Y _83282_/Q sky130_fd_sc_hd__dfxtp_4
X_80494_ _80494_/A _80494_/B _80494_/Y sky130_fd_sc_hd__nand2_4
X_54201_ _54215_/A _47411_/A _54201_/Y sky130_fd_sc_hd__nand2_4
X_85021_ _83008_/CLK _57389_/X _85021_/Q sky130_fd_sc_hd__dfxtp_4
X_51413_ _51403_/X _52940_/B _51413_/Y sky130_fd_sc_hd__nand2_4
X_82233_ _82531_/CLK _82265_/Q _82233_/Q sky130_fd_sc_hd__dfxtp_4
X_55181_ _55179_/X _55181_/B _55298_/A sky130_fd_sc_hd__and2_4
X_67167_ _67046_/A _67167_/X sky130_fd_sc_hd__buf_2
X_52393_ _52373_/X _49144_/X _52393_/Y sky130_fd_sc_hd__nand2_4
X_64379_ _64344_/X _64379_/B _64379_/C _64379_/X sky130_fd_sc_hd__and3_4
X_54132_ _54127_/X _54123_/B _54118_/X _52967_/D _54132_/X sky130_fd_sc_hd__and4_4
X_66118_ _64980_/A _66118_/X sky130_fd_sc_hd__buf_2
X_51344_ _51336_/Y _51339_/X _51343_/X _86029_/D sky130_fd_sc_hd__a21oi_4
X_82164_ _84166_/CLK _84156_/Q _82164_/Q sky130_fd_sc_hd__dfxtp_4
X_67098_ _87421_/Q _66997_/X _66998_/X _67097_/X _67098_/X sky130_fd_sc_hd__a211o_4
X_81115_ _81117_/CLK _79822_/Y _75650_/A sky130_fd_sc_hd__dfxtp_4
X_58940_ _58936_/Y _58938_/Y _58939_/X _58940_/X sky130_fd_sc_hd__a21o_4
X_54063_ _54020_/A _52545_/B _54063_/Y sky130_fd_sc_hd__nand2_4
X_66049_ _66045_/Y _65987_/X _66048_/Y _84160_/D sky130_fd_sc_hd__a21o_4
X_51275_ _51273_/Y _51263_/X _51274_/X _51275_/Y sky130_fd_sc_hd__a21oi_4
X_86972_ _87473_/CLK _44756_/X _86972_/Q sky130_fd_sc_hd__dfxtp_4
X_82095_ _82015_/CLK _82095_/D _82095_/Q sky130_fd_sc_hd__dfxtp_4
X_53014_ _53069_/A _53036_/B sky130_fd_sc_hd__buf_2
X_50226_ _50473_/A _50227_/A sky130_fd_sc_hd__buf_2
X_85923_ _85444_/CLK _51915_/Y _85923_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_333_0_CLK clkbuf_9_166_0_CLK/X _86665_/CLK sky130_fd_sc_hd__clkbuf_1
X_81046_ _81082_/CLK _75370_/X _81046_/Q sky130_fd_sc_hd__dfxtp_4
X_58871_ _58599_/A _58871_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_963_0_CLK clkbuf_9_481_0_CLK/X _85630_/CLK sky130_fd_sc_hd__clkbuf_1
X_57822_ _58098_/A _57822_/X sky130_fd_sc_hd__buf_2
X_69808_ _69897_/A _69808_/B _69808_/Y sky130_fd_sc_hd__nor2_4
X_50157_ _50154_/Y _50141_/X _50156_/X _50157_/Y sky130_fd_sc_hd__a21oi_4
X_85854_ _85566_/CLK _52282_/Y _85854_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_454_0_CLK clkbuf_9_455_0_CLK/A clkbuf_9_454_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_84805_ _84150_/CLK _84805_/D _84805_/Q sky130_fd_sc_hd__dfxtp_4
X_57753_ _84949_/Q _57753_/Y sky130_fd_sc_hd__inv_2
X_69739_ _69736_/X _69738_/X _69678_/X _69739_/X sky130_fd_sc_hd__a21o_4
X_50088_ _48836_/A _50088_/X sky130_fd_sc_hd__buf_2
X_54965_ _54962_/Y _54253_/X _54964_/X _54965_/Y sky130_fd_sc_hd__a21oi_4
X_85785_ _82768_/CLK _85785_/D _85785_/Q sky130_fd_sc_hd__dfxtp_4
X_82997_ _85013_/CLK _74653_/X _82997_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_348_0_CLK clkbuf_9_174_0_CLK/X _85648_/CLK sky130_fd_sc_hd__clkbuf_1
X_56704_ _44290_/X _56704_/X sky130_fd_sc_hd__buf_2
X_87524_ _87782_/CLK _43238_/Y _87524_/Q sky130_fd_sc_hd__dfxtp_4
X_41930_ _41930_/A _41930_/Y sky130_fd_sc_hd__inv_2
X_53916_ _53913_/Y _53914_/X _53915_/Y _85543_/D sky130_fd_sc_hd__a21boi_4
X_72750_ _73257_/A _72750_/X sky130_fd_sc_hd__buf_2
X_84736_ _84829_/CLK _84736_/D _59427_/A sky130_fd_sc_hd__dfxtp_4
X_57684_ _57683_/X _57666_/B _57684_/Y sky130_fd_sc_hd__nor2_4
X_81948_ _81970_/CLK _81948_/D _77628_/A sky130_fd_sc_hd__dfxtp_4
X_54896_ _54910_/A _54883_/B _54910_/C _53203_/D _54896_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_978_0_CLK clkbuf_9_489_0_CLK/X _83613_/CLK sky130_fd_sc_hd__clkbuf_1
X_71701_ _58290_/Y _71695_/X _71700_/Y _71701_/Y sky130_fd_sc_hd__o21ai_4
X_59423_ _59423_/A _59423_/Y sky130_fd_sc_hd__inv_2
X_56635_ _56587_/X _56634_/X _55499_/B _56590_/X _85141_/D sky130_fd_sc_hd__a2bb2o_4
X_87455_ _87720_/CLK _87455_/D _87455_/Q sky130_fd_sc_hd__dfxtp_4
X_41861_ _40363_/X _57491_/B sky130_fd_sc_hd__buf_2
X_53847_ _53956_/A _53848_/A sky130_fd_sc_hd__buf_2
X_72681_ _72683_/A _72683_/B _55387_/X _72681_/Y sky130_fd_sc_hd__nand3_4
X_84667_ _84660_/CLK _84667_/D _60067_/C sky130_fd_sc_hd__dfxtp_4
X_81879_ _82221_/CLK _78070_/X _81879_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_469_0_CLK clkbuf_9_469_0_CLK/A clkbuf_9_469_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_43600_ _40581_/A _43586_/X _68418_/B _43593_/X _43600_/X sky130_fd_sc_hd__a2bb2o_4
X_74420_ _74453_/A _74420_/X sky130_fd_sc_hd__buf_2
X_86406_ _83783_/CLK _49343_/Y _65310_/B sky130_fd_sc_hd__dfxtp_4
X_40812_ _82871_/Q _40847_/B _40812_/X sky130_fd_sc_hd__or2_4
X_83618_ _85562_/CLK _71067_/Y _83618_/Q sky130_fd_sc_hd__dfxtp_4
X_71632_ _71258_/A _71246_/B _71637_/C _71632_/Y sky130_fd_sc_hd__nand3_4
X_59354_ _84748_/Q _59354_/Y sky130_fd_sc_hd__inv_2
X_44580_ _44579_/Y _87047_/D sky130_fd_sc_hd__inv_2
X_56566_ _55640_/Y _56553_/Y _56565_/Y _85153_/D sky130_fd_sc_hd__o21ai_4
X_41792_ _41607_/X _41792_/X sky130_fd_sc_hd__buf_2
X_87386_ _86920_/CLK _87386_/D _87386_/Q sky130_fd_sc_hd__dfxtp_4
X_53778_ _53778_/A _50556_/B _53778_/Y sky130_fd_sc_hd__nand2_4
X_84598_ _84606_/CLK _60569_/Y _79138_/A sky130_fd_sc_hd__dfxtp_4
X_58305_ _63703_/B _58344_/B _58305_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_901_0_CLK clkbuf_9_450_0_CLK/X _82541_/CLK sky130_fd_sc_hd__clkbuf_1
X_43531_ _43178_/X _53443_/A sky130_fd_sc_hd__buf_2
X_55517_ _55516_/X _55517_/X sky130_fd_sc_hd__buf_2
X_74351_ _74351_/A _74342_/X _56117_/C _74351_/Y sky130_fd_sc_hd__nand3_4
X_86337_ _86655_/CLK _49714_/Y _57692_/B sky130_fd_sc_hd__dfxtp_4
X_40743_ _40742_/X _40743_/X sky130_fd_sc_hd__buf_2
X_52729_ _52648_/A _52729_/X sky130_fd_sc_hd__buf_2
X_59285_ _59260_/X _85418_/Q _59284_/X _59285_/Y sky130_fd_sc_hd__o21ai_4
X_71563_ _71698_/A _71553_/B _71558_/X _71563_/Y sky130_fd_sc_hd__nor3_4
X_83549_ _83550_/CLK _71280_/Y _47716_/A sky130_fd_sc_hd__dfxtp_4
X_56497_ _56487_/X _56507_/B _55876_/B _56497_/Y sky130_fd_sc_hd__nand3_4
X_73302_ _88318_/Q _73059_/X _73007_/X _73302_/Y sky130_fd_sc_hd__o21ai_4
X_46250_ _46279_/A _46250_/X sky130_fd_sc_hd__buf_2
X_70514_ _70511_/A _70945_/B _70508_/X _70514_/Y sky130_fd_sc_hd__nand3_4
XPHY_620 sky130_fd_sc_hd__decap_3
X_58236_ _83396_/Q _58236_/Y sky130_fd_sc_hd__inv_2
X_77070_ _77069_/A _82283_/D _77070_/Y sky130_fd_sc_hd__nand2_4
X_43462_ _41636_/X _43446_/X _87410_/Q _43447_/X _43462_/X sky130_fd_sc_hd__a2bb2o_4
X_55448_ _55446_/A _55448_/Y sky130_fd_sc_hd__inv_2
X_86268_ _83306_/CLK _50083_/Y _64755_/B sky130_fd_sc_hd__dfxtp_4
X_74282_ _74280_/X _74281_/Y _72630_/X _74282_/X sky130_fd_sc_hd__a21o_4
XPHY_631 sky130_fd_sc_hd__decap_3
X_40674_ _40673_/X _40651_/X _68750_/B _40652_/X _88356_/D sky130_fd_sc_hd__a2bb2o_4
X_71494_ _71488_/X _71427_/C _71496_/C _71494_/X sky130_fd_sc_hd__and3_4
XPHY_642 sky130_fd_sc_hd__decap_3
XPHY_653 sky130_fd_sc_hd__decap_3
X_45201_ _45195_/X _45199_/Y _45200_/X _45201_/Y sky130_fd_sc_hd__a21oi_4
X_76021_ _81711_/D _76021_/B _76021_/Y sky130_fd_sc_hd__nand2_4
X_88007_ _87249_/CLK _88007_/D _88007_/Q sky130_fd_sc_hd__dfxtp_4
X_42413_ _42412_/Y _42413_/Y sky130_fd_sc_hd__inv_2
XPHY_664 sky130_fd_sc_hd__decap_3
X_73233_ _73206_/X _85871_/Q _73233_/X sky130_fd_sc_hd__and2_4
X_85219_ _85186_/CLK _85219_/D _55713_/B sky130_fd_sc_hd__dfxtp_4
X_46181_ _46098_/A _46181_/Y sky130_fd_sc_hd__inv_2
X_70445_ _71650_/A _74529_/A _71194_/C _70445_/Y sky130_fd_sc_hd__nand3_4
X_58167_ _63069_/A _64272_/A sky130_fd_sc_hd__buf_2
XPHY_675 sky130_fd_sc_hd__decap_3
X_43393_ _41454_/X _43386_/X _87444_/Q _43388_/X _87444_/D sky130_fd_sc_hd__a2bb2o_4
X_55379_ _55378_/X _55379_/Y sky130_fd_sc_hd__inv_2
X_86199_ _86196_/CLK _86199_/D _86199_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_686 sky130_fd_sc_hd__decap_3
XPHY_697 sky130_fd_sc_hd__decap_3
Xclkbuf_10_916_0_CLK clkbuf_9_458_0_CLK/X _84980_/CLK sky130_fd_sc_hd__clkbuf_1
X_45132_ _55846_/B _45131_/X _45087_/X _45132_/X sky130_fd_sc_hd__o21a_4
X_57118_ _57109_/X _56630_/X _85078_/Q _57110_/X _85078_/D sky130_fd_sc_hd__a2bb2o_4
X_42344_ _41697_/X _42342_/X _87911_/Q _42343_/X _87911_/D sky130_fd_sc_hd__a2bb2o_4
X_73164_ _72814_/A _73165_/A sky130_fd_sc_hd__buf_2
X_70376_ _50852_/B _70364_/X _70375_/Y _70376_/Y sky130_fd_sc_hd__o21ai_4
X_58098_ _58098_/A _58098_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_5_0_CLK clkbuf_9_2_0_CLK/X _85297_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_9_407_0_CLK clkbuf_9_407_0_CLK/A clkbuf_9_407_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_72115_ _72250_/A _72115_/X sky130_fd_sc_hd__buf_2
X_49940_ _49955_/A _53153_/B _49940_/Y sky130_fd_sc_hd__nand2_4
X_45063_ _45212_/A _45063_/X sky130_fd_sc_hd__buf_2
X_57049_ _57049_/A _85096_/Q _56953_/A _57049_/Y sky130_fd_sc_hd__nor3_4
X_42275_ _42199_/X _42275_/X sky130_fd_sc_hd__buf_2
X_73095_ _73091_/X _73094_/X _73067_/X _73098_/A sky130_fd_sc_hd__a21o_4
X_77972_ _77971_/X _77972_/Y sky130_fd_sc_hd__inv_2
X_44014_ _44174_/A _45920_/A sky130_fd_sc_hd__inv_2
X_79711_ _65072_/C _72323_/Y _79710_/Y _79711_/X sky130_fd_sc_hd__o21a_4
X_41226_ _41205_/X _41206_/X _41225_/X _88254_/Q _41194_/X _41227_/A
+ sky130_fd_sc_hd__o32ai_4
X_60060_ _84669_/Q _60053_/X _60059_/Y _60060_/X sky130_fd_sc_hd__o21a_4
X_72046_ _72040_/A _49064_/A _72046_/Y sky130_fd_sc_hd__nand2_4
X_76923_ _76919_/Y _76922_/Y _76924_/A sky130_fd_sc_hd__xor2_4
X_49871_ _49925_/A _49893_/A sky130_fd_sc_hd__buf_2
X_48822_ _50105_/A _50069_/A sky130_fd_sc_hd__buf_2
X_79642_ _79619_/A _79642_/B _79619_/B _79642_/D _79642_/Y sky130_fd_sc_hd__nand4_4
X_41157_ _41157_/A _41157_/X sky130_fd_sc_hd__buf_2
X_76854_ _76854_/A _76854_/B _81464_/D sky130_fd_sc_hd__xor2_4
X_75805_ _75802_/B _75796_/Y _75804_/Y _75810_/C sky130_fd_sc_hd__o21a_4
X_48753_ _48751_/Y _48734_/X _48752_/X _48753_/Y sky130_fd_sc_hd__a21oi_4
X_79573_ _79569_/Y _79573_/B _79572_/Y _79576_/B sky130_fd_sc_hd__nand3_4
X_45965_ _41797_/X _45963_/X _66577_/B _45964_/X _45965_/X sky130_fd_sc_hd__a2bb2o_4
X_41088_ _40995_/A _41088_/X sky130_fd_sc_hd__buf_2
X_76785_ _81697_/Q _76785_/B _76785_/Y sky130_fd_sc_hd__xnor2_4
X_73997_ _73994_/X _73996_/X _72735_/X _74000_/A sky130_fd_sc_hd__a21o_4
X_47704_ _47704_/A _54894_/B sky130_fd_sc_hd__inv_2
X_78524_ _78524_/A _82673_/D _78525_/A sky130_fd_sc_hd__nand2_4
X_44916_ _44913_/Y _44915_/Y _44889_/X _44916_/X sky130_fd_sc_hd__a21o_4
X_63750_ _60996_/B _63753_/C sky130_fd_sc_hd__buf_2
X_75736_ _75723_/A _75736_/B _75736_/X sky130_fd_sc_hd__and2_4
X_60962_ _60962_/A _60962_/Y sky130_fd_sc_hd__inv_2
X_48684_ _48695_/A _48684_/B _48684_/Y sky130_fd_sc_hd__nand2_4
X_72948_ _43133_/Y _72830_/X _72799_/X _72947_/Y _72948_/X sky130_fd_sc_hd__a211o_4
X_45896_ _73948_/A _45896_/X sky130_fd_sc_hd__buf_2
Xclkbuf_6_7_0_CLK clkbuf_6_7_0_CLK/A clkbuf_6_7_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_62701_ _58232_/X _62689_/X _60205_/X _62699_/X _62700_/X _62701_/Y
+ sky130_fd_sc_hd__a41oi_4
X_47635_ _81238_/Q _47636_/A sky130_fd_sc_hd__inv_2
X_78455_ _78455_/A _82668_/D _78455_/Y sky130_fd_sc_hd__nand2_4
X_44847_ _41741_/A _44838_/X _67836_/B _44839_/X _86922_/D sky130_fd_sc_hd__a2bb2o_4
X_63681_ _63678_/Y _63679_/X _63680_/Y _63681_/Y sky130_fd_sc_hd__a21oi_4
X_75667_ _81004_/Q _75667_/B _75667_/X sky130_fd_sc_hd__xor2_4
X_60893_ _60892_/Y _64180_/C sky130_fd_sc_hd__buf_2
X_72879_ _72784_/A _72880_/A sky130_fd_sc_hd__buf_2
X_65420_ _65399_/X _65410_/Y _65419_/Y _65420_/Y sky130_fd_sc_hd__o21ai_4
X_77406_ _77406_/A _82094_/D _77406_/Y sky130_fd_sc_hd__nand2_4
X_62632_ _62632_/A _84882_/Q _62632_/C _62634_/C sky130_fd_sc_hd__nand3_4
X_74618_ _45319_/A _74612_/X _74617_/X _83014_/D sky130_fd_sc_hd__o21ai_4
X_47566_ _81245_/Q _47567_/A sky130_fd_sc_hd__inv_2
X_78386_ _78385_/Y _78386_/Y sky130_fd_sc_hd__inv_2
X_44778_ _41366_/Y _44774_/X _86960_/Q _44775_/X _86960_/D sky130_fd_sc_hd__a2bb2o_4
X_75598_ _75598_/A _75607_/B sky130_fd_sc_hd__inv_2
X_49305_ _49303_/Y _49281_/X _49304_/X _49305_/Y sky130_fd_sc_hd__a21oi_4
X_46517_ _46408_/A _49322_/B _46517_/Y sky130_fd_sc_hd__nand2_4
X_65351_ _64667_/A _65401_/A sky130_fd_sc_hd__buf_2
X_77337_ _81929_/Q _82185_/D _77337_/X sky130_fd_sc_hd__xor2_4
X_43729_ _40885_/A _43716_/X _69862_/B _43718_/X _43729_/X sky130_fd_sc_hd__a2bb2o_4
X_62563_ _62551_/X _62553_/X _84401_/Q _62563_/Y sky130_fd_sc_hd__nor3_4
X_74549_ _74549_/A _45955_/X _74549_/Y sky130_fd_sc_hd__nand2_4
X_47497_ _47497_/A _54772_/B sky130_fd_sc_hd__inv_2
X_64302_ _64243_/A _64304_/A sky130_fd_sc_hd__buf_2
X_49236_ _49233_/Y _49189_/X _49235_/X _49236_/Y sky130_fd_sc_hd__a21oi_4
X_61514_ _59421_/A _61484_/B _61484_/C _61514_/D _61514_/Y sky130_fd_sc_hd__nand4_4
X_68070_ _69779_/A _68070_/X sky130_fd_sc_hd__buf_2
X_46448_ _46301_/X _82928_/Q _46447_/Y _46449_/A sky130_fd_sc_hd__o21ai_4
X_65282_ _65258_/A _65282_/B _65282_/X sky130_fd_sc_hd__and2_4
X_77268_ _77254_/Y _77250_/A _77253_/A _77268_/X sky130_fd_sc_hd__o21a_4
X_62494_ _62336_/A _62570_/A sky130_fd_sc_hd__buf_2
X_67021_ _66553_/X _67144_/A sky130_fd_sc_hd__buf_2
X_79007_ _78998_/A _78998_/B _78997_/A _78997_/B _79007_/X sky130_fd_sc_hd__o22a_4
X_64233_ _63389_/A _64219_/B _64233_/Y sky130_fd_sc_hd__nor2_4
X_76219_ _76219_/A _76201_/Y _76219_/Y sky130_fd_sc_hd__nand2_4
X_49167_ _49166_/Y _50708_/B sky130_fd_sc_hd__buf_2
X_61445_ _61434_/A _61434_/B _79148_/B _61445_/Y sky130_fd_sc_hd__nor3_4
X_46379_ _86742_/Q _46364_/X _46378_/Y _46379_/Y sky130_fd_sc_hd__o21ai_4
X_77199_ _82109_/Q _77199_/B _77199_/X sky130_fd_sc_hd__xor2_4
X_48118_ _82342_/Q _48086_/B _48118_/X sky130_fd_sc_hd__or2_4
X_64164_ _64187_/A _64187_/B _79937_/B _64164_/Y sky130_fd_sc_hd__nor3_4
X_49098_ _48881_/X _81772_/Q _49097_/Y _49099_/A sky130_fd_sc_hd__o21ai_4
X_61376_ _84853_/Q _61376_/X sky130_fd_sc_hd__buf_2
X_63115_ _63111_/Y _63113_/X _63114_/X _63115_/Y sky130_fd_sc_hd__a21oi_4
X_48049_ _47840_/A _48049_/X sky130_fd_sc_hd__buf_2
X_60327_ _60255_/B _60228_/A _60781_/A _60327_/X sky130_fd_sc_hd__a21o_4
X_68972_ _68969_/X _68971_/X _68878_/X _68972_/Y sky130_fd_sc_hd__a21oi_4
X_64095_ _63629_/B _64095_/B _64095_/C _64095_/D _64095_/Y sky130_fd_sc_hd__nand4_4
X_51060_ _51141_/A _51071_/C sky130_fd_sc_hd__buf_2
X_67923_ _81481_/D _67806_/X _67922_/X _84049_/D sky130_fd_sc_hd__a21bo_4
X_63046_ _79476_/A _63008_/X _63045_/Y _63046_/X sky130_fd_sc_hd__a21o_4
X_79909_ _79909_/A _79913_/A _79913_/B _79915_/A sky130_fd_sc_hd__nand3_4
X_60258_ _60257_/X _60259_/A sky130_fd_sc_hd__buf_2
X_50011_ _50008_/Y _50003_/X _50010_/X _86282_/D sky130_fd_sc_hd__a21oi_4
X_82920_ _82931_/CLK _78173_/X _82920_/Q sky130_fd_sc_hd__dfxtp_4
X_67854_ _87965_/Q _67831_/X _67761_/X _67853_/X _67854_/X sky130_fd_sc_hd__a211o_4
X_60189_ _60189_/A _60189_/Y sky130_fd_sc_hd__inv_2
X_66805_ _66757_/X _66791_/Y _66793_/X _66804_/Y _66805_/X sky130_fd_sc_hd__a211o_4
X_82851_ _82563_/CLK _78091_/B _40923_/A sky130_fd_sc_hd__dfxtp_4
X_67785_ _67739_/X _86924_/Q _67785_/X sky130_fd_sc_hd__and2_4
X_64997_ _65047_/A _64870_/B _64997_/C _64997_/Y sky130_fd_sc_hd__nor3_4
X_81802_ _83184_/CLK _81802_/D _81802_/Q sky130_fd_sc_hd__dfxtp_4
X_69524_ _87511_/Q _69356_/X _69371_/X _69523_/X _69524_/X sky130_fd_sc_hd__a211o_4
X_54750_ _54731_/X _47459_/A _54750_/Y sky130_fd_sc_hd__nand2_4
X_66736_ _66760_/A _87628_/Q _66736_/X sky130_fd_sc_hd__and2_4
X_85570_ _83572_/CLK _85570_/D _85570_/Q sky130_fd_sc_hd__dfxtp_4
X_51962_ _51961_/X _50260_/B _51962_/Y sky130_fd_sc_hd__nand2_4
X_63948_ _60930_/C _64027_/D sky130_fd_sc_hd__buf_2
X_82782_ _82975_/CLK _82782_/D _82782_/Q sky130_fd_sc_hd__dfxtp_4
X_53701_ _51842_/A _53763_/A sky130_fd_sc_hd__buf_2
X_84521_ _84623_/CLK _61091_/Y _61089_/C sky130_fd_sc_hd__dfxtp_4
X_50913_ _86108_/Q _50910_/X _50912_/Y _50913_/Y sky130_fd_sc_hd__o21ai_4
X_81733_ _84020_/CLK _75944_/B _41435_/A sky130_fd_sc_hd__dfxtp_4
X_69455_ _87516_/Q _69442_/X _69396_/X _69454_/X _69455_/X sky130_fd_sc_hd__a211o_4
X_54681_ _54679_/Y _54666_/X _54680_/X _54681_/Y sky130_fd_sc_hd__a21oi_4
X_66667_ _66547_/A _66667_/X sky130_fd_sc_hd__buf_2
X_51893_ _51887_/A _51870_/B _51893_/C _52720_/D _51893_/X sky130_fd_sc_hd__and4_4
X_63879_ _63874_/X _63810_/X _63876_/Y _63877_/Y _63878_/X _63879_/X
+ sky130_fd_sc_hd__a41o_4
X_56420_ _56418_/A _56418_/B _56420_/C _56420_/Y sky130_fd_sc_hd__nand3_4
X_68406_ _87506_/Q _68365_/X _68053_/X _68405_/X _68406_/X sky130_fd_sc_hd__a211o_4
X_87240_ _88012_/CLK _43838_/X _87240_/Q sky130_fd_sc_hd__dfxtp_4
X_53632_ _53629_/Y _53619_/X _53631_/X _53632_/Y sky130_fd_sc_hd__a21oi_4
X_65618_ _65615_/X _65663_/B _65617_/X _65619_/B sky130_fd_sc_hd__nand3_4
X_84452_ _84452_/CLK _61822_/Y _78075_/B sky130_fd_sc_hd__dfxtp_4
X_50844_ _50638_/A _50845_/A sky130_fd_sc_hd__buf_2
X_81664_ _81587_/CLK _76773_/A _81664_/Q sky130_fd_sc_hd__dfxtp_4
X_69386_ _69382_/X _69384_/X _69385_/X _69386_/X sky130_fd_sc_hd__a21o_4
X_66598_ _69454_/A _66598_/B _66598_/X sky130_fd_sc_hd__and2_4
X_83403_ _83372_/CLK _83403_/D _58303_/A sky130_fd_sc_hd__dfxtp_4
X_80615_ _80613_/X _80614_/X _80615_/Y sky130_fd_sc_hd__xnor2_4
X_68337_ _83979_/Q _68318_/X _68336_/X _83979_/D sky130_fd_sc_hd__a21bo_4
X_56351_ _56351_/A _56358_/B sky130_fd_sc_hd__buf_2
X_87171_ _87169_/CLK _44311_/Y _43987_/A sky130_fd_sc_hd__dfxtp_4
X_65549_ _65184_/A _85881_/Q _65549_/X sky130_fd_sc_hd__and2_4
X_53563_ _53548_/A _48051_/Y _53563_/Y sky130_fd_sc_hd__nand2_4
X_84383_ _84520_/CLK _84383_/D _84383_/Q sky130_fd_sc_hd__dfxtp_4
X_50775_ _50742_/A _50775_/X sky130_fd_sc_hd__buf_2
X_81595_ _84064_/CLK _65531_/C _81595_/Q sky130_fd_sc_hd__dfxtp_4
X_55302_ _55192_/A _55317_/A sky130_fd_sc_hd__buf_2
X_86122_ _86122_/CLK _86122_/D _86122_/Q sky130_fd_sc_hd__dfxtp_4
X_52514_ _52512_/Y _52486_/X _52513_/Y _52514_/Y sky130_fd_sc_hd__a21boi_4
X_59070_ _58810_/A _59070_/X sky130_fd_sc_hd__buf_2
X_83334_ _83335_/CLK _83334_/D _83334_/Q sky130_fd_sc_hd__dfxtp_4
X_56282_ _73024_/B _56460_/B _56278_/A _56460_/D _56282_/Y sky130_fd_sc_hd__nand4_4
X_80546_ _80538_/X _80540_/B _80545_/Y _80550_/A sky130_fd_sc_hd__a21boi_4
X_68268_ _68447_/A _68268_/X sky130_fd_sc_hd__buf_2
X_53494_ _53491_/Y _53472_/X _53493_/X _53494_/Y sky130_fd_sc_hd__a21oi_4
X_58021_ _57966_/X _85708_/Q _58020_/X _58021_/X sky130_fd_sc_hd__o21a_4
X_55233_ _55230_/X _55232_/X _55138_/A _55655_/A sky130_fd_sc_hd__a21o_4
X_67219_ _88376_/Q _67193_/X _67194_/X _67218_/X _67219_/X sky130_fd_sc_hd__a211o_4
X_86053_ _86054_/CLK _86053_/D _86053_/Q sky130_fd_sc_hd__dfxtp_4
X_52445_ _64694_/B _52422_/X _52444_/Y _52445_/Y sky130_fd_sc_hd__o21ai_4
X_83265_ _81233_/CLK _83265_/D _72313_/A sky130_fd_sc_hd__dfxtp_4
X_80477_ _80489_/A _80489_/B _80480_/A sky130_fd_sc_hd__xor2_4
X_68199_ _84014_/Q _68180_/X _68198_/X _68199_/X sky130_fd_sc_hd__a21bo_4
X_85004_ _85034_/CLK _85004_/D _85004_/Q sky130_fd_sc_hd__dfxtp_4
X_70230_ _70224_/X _83829_/Q _70229_/X _83829_/D sky130_fd_sc_hd__a21o_4
X_82216_ _82084_/CLK _82248_/Q _77308_/A sky130_fd_sc_hd__dfxtp_4
X_55164_ _83747_/Q _55423_/B _55163_/Y _55164_/X sky130_fd_sc_hd__o21a_4
X_40390_ _40381_/X _81181_/Q _40389_/X _40390_/Y sky130_fd_sc_hd__o21ai_4
X_52376_ _52309_/A _52446_/B sky130_fd_sc_hd__buf_2
X_83196_ _83191_/CLK _83196_/D _70210_/C sky130_fd_sc_hd__dfxtp_4
X_54115_ _54134_/A _47260_/A _54115_/Y sky130_fd_sc_hd__nand2_4
X_51327_ _51325_/Y _51313_/X _51326_/X _51327_/Y sky130_fd_sc_hd__a21oi_4
X_70161_ _70154_/X _70348_/B sky130_fd_sc_hd__buf_2
X_82147_ _82147_/CLK _84139_/Q _82147_/Q sky130_fd_sc_hd__dfxtp_4
X_55095_ _46614_/X _55112_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_272_0_CLK clkbuf_9_136_0_CLK/X _83415_/CLK sky130_fd_sc_hd__clkbuf_1
X_59972_ _62534_/A _59995_/A sky130_fd_sc_hd__buf_2
X_58923_ _58923_/A _58923_/X sky130_fd_sc_hd__buf_2
X_54046_ _85516_/Q _54035_/X _54045_/Y _54046_/Y sky130_fd_sc_hd__o21ai_4
X_42060_ _43129_/A _42060_/X sky130_fd_sc_hd__buf_2
X_51258_ _48808_/A _51259_/A sky130_fd_sc_hd__buf_2
X_70092_ _69960_/X _69962_/X _68400_/X _70092_/Y sky130_fd_sc_hd__a21oi_4
X_86955_ _88232_/CLK _86955_/D _86955_/Q sky130_fd_sc_hd__dfxtp_4
X_82078_ _81169_/CLK _82078_/D _82078_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_54_0_CLK clkbuf_9_27_0_CLK/X _85100_/CLK sky130_fd_sc_hd__clkbuf_1
X_41011_ _41010_/Y _41011_/Y sky130_fd_sc_hd__inv_2
X_50209_ _50209_/A _51256_/B _50147_/C _50209_/X sky130_fd_sc_hd__and3_4
X_73920_ _72979_/X _73920_/X sky130_fd_sc_hd__buf_2
X_85906_ _86554_/CLK _52012_/Y _85906_/Q sky130_fd_sc_hd__dfxtp_4
X_81029_ _84197_/CLK _75122_/Y _81029_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_393_0_CLK clkbuf_9_393_0_CLK/A clkbuf_9_393_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_58854_ _58748_/X _58851_/Y _58853_/Y _58766_/X _58752_/X _58854_/X
+ sky130_fd_sc_hd__o32a_4
X_51189_ _51184_/X _52881_/B _51189_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_200_0_CLK clkbuf_8_201_0_CLK/A clkbuf_8_200_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_86886_ _80664_/CLK _45296_/Y _64494_/B sky130_fd_sc_hd__dfxtp_4
X_57805_ _58697_/A _58080_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_287_0_CLK clkbuf_9_143_0_CLK/X _85492_/CLK sky130_fd_sc_hd__clkbuf_1
X_73851_ _73709_/X _73949_/A sky130_fd_sc_hd__buf_2
X_85837_ _85837_/CLK _52366_/Y _65130_/B sky130_fd_sc_hd__dfxtp_4
X_58785_ _58785_/A _64836_/A sky130_fd_sc_hd__buf_2
X_55997_ _55996_/X _55997_/X sky130_fd_sc_hd__buf_2
X_72802_ _72797_/X _72801_/X _72737_/X _72802_/X sky130_fd_sc_hd__a21o_4
X_57736_ _57736_/A _57736_/X sky130_fd_sc_hd__buf_2
X_45750_ _45748_/X _61597_/A _45685_/X _45750_/Y sky130_fd_sc_hd__o21ai_4
X_76570_ _76569_/Y _76571_/B sky130_fd_sc_hd__inv_2
X_42962_ _42962_/A _42962_/X sky130_fd_sc_hd__buf_2
X_54948_ _53460_/A _47809_/A _54948_/Y sky130_fd_sc_hd__nand2_4
X_85768_ _85770_/CLK _52717_/Y _85768_/Q sky130_fd_sc_hd__dfxtp_4
X_73782_ _73284_/A _73782_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_69_0_CLK clkbuf_9_34_0_CLK/X _80657_/CLK sky130_fd_sc_hd__clkbuf_1
X_70994_ _70994_/A _71080_/B sky130_fd_sc_hd__buf_2
X_44701_ _44679_/X _44680_/X _40661_/X _86994_/Q _44681_/X _44702_/A
+ sky130_fd_sc_hd__o32ai_4
X_87507_ _87520_/CLK _43271_/Y _87507_/Q sky130_fd_sc_hd__dfxtp_4
X_75521_ _75498_/A _75495_/Y _75497_/A _75522_/A sky130_fd_sc_hd__o21a_4
X_41913_ _40626_/X _41907_/X _88108_/Q _41912_/X _41913_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_8_215_0_CLK clkbuf_8_215_0_CLK/A clkbuf_9_430_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_72733_ _43113_/Y _72731_/X _56935_/X _72732_/Y _72733_/X sky130_fd_sc_hd__a211o_4
X_84719_ _84903_/CLK _59487_/Y _64236_/C sky130_fd_sc_hd__dfxtp_4
X_45681_ _45681_/A _74667_/B sky130_fd_sc_hd__inv_2
X_57667_ _57650_/X _57663_/Y _57666_/Y _57667_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_210_0_CLK clkbuf_9_105_0_CLK/X _84503_/CLK sky130_fd_sc_hd__clkbuf_1
X_42893_ _41647_/X _42886_/X _67415_/B _42887_/X _87664_/D sky130_fd_sc_hd__a2bb2o_4
X_54879_ _54877_/Y _54856_/X _54878_/X _85361_/D sky130_fd_sc_hd__a21oi_4
X_85699_ _86688_/CLK _53091_/Y _85699_/Q sky130_fd_sc_hd__dfxtp_4
X_47420_ _83732_/Q _47420_/Y sky130_fd_sc_hd__inv_2
X_59406_ _63150_/A _59407_/A sky130_fd_sc_hd__buf_2
X_78240_ _78240_/A _78240_/B _78240_/X sky130_fd_sc_hd__xor2_4
X_44632_ _44622_/X _44623_/X _41016_/A _87025_/Q _44625_/X _44633_/A
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_10_840_0_CLK clkbuf_9_420_0_CLK/X _82177_/CLK sky130_fd_sc_hd__clkbuf_1
X_56618_ _72656_/C _56618_/B _56619_/A sky130_fd_sc_hd__xor2_4
X_75452_ _80795_/Q _75451_/Y _80763_/D sky130_fd_sc_hd__xor2_4
X_41844_ _40497_/X _41813_/X _88126_/Q _41814_/X _88126_/D sky130_fd_sc_hd__a2bb2o_4
X_87438_ _87484_/CLK _43403_/X _87438_/Q sky130_fd_sc_hd__dfxtp_4
X_72664_ _72668_/A _72668_/B _72664_/C _72664_/Y sky130_fd_sc_hd__nand3_4
X_57598_ _57596_/Y _57581_/X _57597_/Y _84972_/D sky130_fd_sc_hd__a21boi_4
X_74403_ _74408_/A _74403_/B _74403_/Y sky130_fd_sc_hd__nand2_4
X_47351_ _83739_/Q _47352_/A sky130_fd_sc_hd__inv_2
X_71615_ _71604_/X _83438_/Q _71614_/Y _83438_/D sky130_fd_sc_hd__a21o_4
X_59337_ _59333_/Y _59336_/Y _59278_/X _59337_/X sky130_fd_sc_hd__a21o_4
X_78171_ _78166_/Y _78167_/A _78170_/Y _78171_/Y sky130_fd_sc_hd__a21boi_4
X_44563_ _44547_/X _44548_/X _40861_/X _87053_/Q _44549_/X _44564_/A
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_9_331_0_CLK clkbuf_9_331_0_CLK/A clkbuf_9_331_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_56549_ _56548_/X _56549_/X sky130_fd_sc_hd__buf_2
X_87369_ _87373_/CLK _87369_/D _87369_/Q sky130_fd_sc_hd__dfxtp_4
X_75383_ _75383_/A _75383_/B _75383_/C _75383_/X sky130_fd_sc_hd__or3_4
X_41775_ _41775_/A _88152_/D sky130_fd_sc_hd__inv_2
X_72595_ _72607_/B _72549_/B _59846_/X _72597_/C _72595_/X sky130_fd_sc_hd__a211o_4
X_46302_ _46302_/A _48924_/A sky130_fd_sc_hd__inv_2
X_77122_ _77122_/A _77121_/Y _77123_/B sky130_fd_sc_hd__xnor2_4
X_43514_ _43466_/X _43514_/X sky130_fd_sc_hd__buf_2
X_74334_ _74338_/A _74338_/B _56108_/A _74334_/Y sky130_fd_sc_hd__nand3_4
X_40726_ _40726_/A _40726_/Y sky130_fd_sc_hd__inv_2
X_47282_ _81819_/Q _47283_/A sky130_fd_sc_hd__inv_2
Xclkbuf_10_225_0_CLK clkbuf_9_112_0_CLK/X _80708_/CLK sky130_fd_sc_hd__clkbuf_1
X_59268_ _59043_/A _59268_/X sky130_fd_sc_hd__buf_2
X_71546_ _70682_/A _71546_/B _71546_/C _71546_/Y sky130_fd_sc_hd__nor3_4
X_44494_ _44481_/X _44482_/X _41233_/X _87080_/Q _44484_/X _44495_/A
+ sky130_fd_sc_hd__o32ai_4
X_49021_ _49021_/A _72025_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_855_0_CLK clkbuf_9_427_0_CLK/X _82965_/CLK sky130_fd_sc_hd__clkbuf_1
X_46233_ _44120_/Y HASH_EN _46233_/Y sky130_fd_sc_hd__nand2_4
X_58219_ _58341_/A _58219_/X sky130_fd_sc_hd__buf_2
XPHY_450 sky130_fd_sc_hd__decap_3
X_77053_ _77038_/X _77045_/X _77053_/Y sky130_fd_sc_hd__nand2_4
X_43445_ _43178_/X _43513_/A sky130_fd_sc_hd__buf_2
X_74265_ _69110_/Y _73891_/X _45897_/X _74264_/Y _74265_/X sky130_fd_sc_hd__a211o_4
XPHY_461 sky130_fd_sc_hd__decap_3
X_40657_ _40635_/X _40638_/X _40656_/X _88359_/Q _40612_/X _40657_/Y
+ sky130_fd_sc_hd__o32ai_4
X_71477_ _71464_/X _83485_/Q _71476_/X _83485_/D sky130_fd_sc_hd__a21o_4
X_59199_ _58904_/A _59199_/X sky130_fd_sc_hd__buf_2
XPHY_472 sky130_fd_sc_hd__decap_3
XPHY_483 sky130_fd_sc_hd__decap_3
X_76004_ _81710_/D _76013_/B _76010_/A sky130_fd_sc_hd__xor2_4
X_73216_ _73214_/X _83064_/Q _73015_/X _73215_/X _73216_/X sky130_fd_sc_hd__a211o_4
XPHY_494 sky130_fd_sc_hd__decap_3
X_61230_ _61109_/X _61271_/A _61230_/C _61264_/B sky130_fd_sc_hd__nand3_4
Xclkbuf_9_346_0_CLK clkbuf_9_347_0_CLK/A clkbuf_9_346_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_46164_ _46164_/A _46188_/A _46169_/C sky130_fd_sc_hd__nor2_4
X_70428_ _70428_/A _71145_/A sky130_fd_sc_hd__inv_2
X_43376_ _43367_/X _43375_/X _41403_/X _87453_/Q _43353_/X _43376_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74196_ _74193_/X _74195_/X _56547_/X _74199_/A sky130_fd_sc_hd__a21o_4
X_40588_ _40588_/A _40588_/B _40588_/X sky130_fd_sc_hd__or2_4
X_45115_ _45389_/A _45265_/A sky130_fd_sc_hd__buf_2
X_42327_ _41647_/X _42325_/X _87920_/Q _42326_/X _87920_/D sky130_fd_sc_hd__a2bb2o_4
X_61161_ _61179_/A _61153_/C _64456_/C _61254_/C sky130_fd_sc_hd__nand3_4
X_73147_ _42583_/A _72892_/B _73147_/Y sky130_fd_sc_hd__nor2_4
X_46095_ _46092_/X _46121_/A _46094_/X _46096_/D sky130_fd_sc_hd__nor3_4
X_70359_ HASH_ADDR[1] _70907_/B sky130_fd_sc_hd__buf_2
X_60112_ _60111_/X _64638_/B sky130_fd_sc_hd__buf_2
X_49923_ _86298_/Q _49906_/X _49922_/Y _49923_/Y sky130_fd_sc_hd__o21ai_4
X_45046_ _45046_/A _45046_/Y sky130_fd_sc_hd__inv_2
X_42258_ _42258_/A _42258_/X sky130_fd_sc_hd__buf_2
X_73078_ _73078_/A _73193_/A sky130_fd_sc_hd__buf_2
X_77955_ _77950_/B _77950_/A _77955_/X sky130_fd_sc_hd__and2_4
X_61092_ _64361_/A _64243_/A sky130_fd_sc_hd__buf_2
X_41209_ _41209_/A _41209_/X sky130_fd_sc_hd__buf_2
X_64920_ _64948_/A _64920_/B _64920_/X sky130_fd_sc_hd__and2_4
X_60043_ _59922_/C _60091_/A _59985_/X _60044_/A sky130_fd_sc_hd__and3_4
X_72029_ _72025_/A _53854_/B _72029_/Y sky130_fd_sc_hd__nand2_4
X_76906_ _76906_/A _76906_/Y sky130_fd_sc_hd__inv_2
X_49854_ _49854_/A _49864_/A sky130_fd_sc_hd__buf_2
X_42189_ _42189_/A _87989_/D sky130_fd_sc_hd__inv_2
X_77886_ _77880_/B _77880_/A _77885_/Y _77886_/Y sky130_fd_sc_hd__a21oi_4
X_48805_ _52194_/A _48829_/B _48814_/C _48805_/X sky130_fd_sc_hd__and3_4
X_79625_ _65268_/C _83256_/Q _79625_/Y sky130_fd_sc_hd__nand2_4
X_64851_ _64851_/A _64851_/X sky130_fd_sc_hd__buf_2
X_76837_ _76837_/A _76837_/B _76838_/B sky130_fd_sc_hd__xor2_4
X_49785_ _49769_/X _52999_/B _49785_/Y sky130_fd_sc_hd__nand2_4
X_46997_ _46903_/A _47029_/C sky130_fd_sc_hd__buf_2
X_63802_ _60920_/A _63803_/C sky130_fd_sc_hd__buf_2
X_48736_ _48733_/Y _48734_/X _48735_/X _86493_/D sky130_fd_sc_hd__a21oi_4
X_67570_ _67569_/X _87657_/Q _67570_/X sky130_fd_sc_hd__and2_4
X_79556_ _79555_/B _79555_/C _79557_/A sky130_fd_sc_hd__nand2_4
X_45948_ _45918_/Y _45947_/Y _86840_/Q _45948_/Y sky130_fd_sc_hd__a21boi_4
X_64782_ _64779_/X _64781_/X _64629_/X _64782_/X sky130_fd_sc_hd__a21o_4
X_76768_ _76768_/A _76755_/Y _76768_/Y sky130_fd_sc_hd__nor2_4
X_61994_ _61541_/B _61933_/X _61967_/C _61952_/D _62000_/B sky130_fd_sc_hd__nand4_4
X_66521_ _65415_/X _66521_/B _65418_/X _66521_/Y sky130_fd_sc_hd__nand3_4
X_78507_ _78487_/Y _78488_/Y _78489_/Y _78508_/A sky130_fd_sc_hd__o21a_4
X_63733_ _61278_/A _63733_/X sky130_fd_sc_hd__buf_2
X_75719_ _75695_/Y _75719_/Y sky130_fd_sc_hd__inv_2
X_48667_ _48667_/A _48657_/B _48657_/C _48667_/X sky130_fd_sc_hd__and3_4
X_60945_ _65515_/A _72543_/A sky130_fd_sc_hd__buf_2
X_79487_ _79487_/A _79487_/Y sky130_fd_sc_hd__inv_2
X_45879_ _45819_/X _61695_/A _45836_/X _45879_/Y sky130_fd_sc_hd__o21ai_4
X_76699_ _76691_/A _81351_/D _76699_/X sky130_fd_sc_hd__or2_4
Xclkbuf_10_808_0_CLK clkbuf_9_404_0_CLK/X _82343_/CLK sky130_fd_sc_hd__clkbuf_1
X_69240_ _69128_/X _88300_/Q _69240_/X sky130_fd_sc_hd__and2_4
X_47618_ _47612_/Y _47602_/X _47617_/X _86616_/D sky130_fd_sc_hd__a21oi_4
X_66452_ _66448_/Y _66449_/X _66451_/Y _84121_/D sky130_fd_sc_hd__a21o_4
X_78438_ _78436_/Y _78438_/Y sky130_fd_sc_hd__inv_2
X_63664_ _63662_/Y _63635_/X _63663_/Y _63664_/Y sky130_fd_sc_hd__a21oi_4
X_48598_ _46423_/X _48056_/A _48597_/X _48823_/B sky130_fd_sc_hd__o21ai_4
X_60876_ _60909_/A _60934_/A sky130_fd_sc_hd__inv_2
X_65403_ _65403_/A _86242_/Q _65403_/X sky130_fd_sc_hd__and2_4
X_62615_ _62608_/X _62610_/X _62614_/Y _84868_/Q _62572_/X _62615_/Y
+ sky130_fd_sc_hd__o32ai_4
X_69171_ _69156_/A _69171_/X sky130_fd_sc_hd__buf_2
X_47549_ _47530_/X _47549_/B _47519_/X _53113_/D _47549_/X sky130_fd_sc_hd__and4_4
X_66383_ _66381_/Y _66382_/Y _65842_/X _66383_/Y sky130_fd_sc_hd__a21oi_4
X_78369_ _78369_/A _78369_/B _82758_/D sky130_fd_sc_hd__xnor2_4
X_63595_ _63546_/A _58483_/A _63581_/X _63595_/D _63595_/X sky130_fd_sc_hd__and4_4
X_80400_ _80400_/A _80400_/B _80400_/X sky130_fd_sc_hd__xor2_4
X_68122_ _66776_/X _66778_/X _68106_/X _68122_/Y sky130_fd_sc_hd__a21oi_4
X_65334_ _64752_/A _65334_/X sky130_fd_sc_hd__buf_2
X_50560_ _50496_/A _50560_/X sky130_fd_sc_hd__buf_2
X_62546_ _60056_/A _84834_/Q _59936_/X _62081_/B _62549_/A sky130_fd_sc_hd__a22oi_4
X_81380_ _83918_/CLK _81380_/D _76811_/B sky130_fd_sc_hd__dfxtp_4
X_49219_ _64647_/B _48548_/X _49218_/Y _49219_/Y sky130_fd_sc_hd__o21ai_4
X_80331_ _80329_/Y _80330_/Y _80331_/Y sky130_fd_sc_hd__nand2_4
X_68053_ _68450_/A _68053_/X sky130_fd_sc_hd__buf_2
X_65265_ _65178_/X _86728_/Q _65239_/X _65264_/X _65265_/X sky130_fd_sc_hd__a211o_4
X_50491_ _50491_/A _50491_/X sky130_fd_sc_hd__buf_2
X_62477_ _62493_/A _62472_/Y _62477_/C _62476_/Y _62477_/Y sky130_fd_sc_hd__nand4_4
X_67004_ _88385_/Q _66954_/X _66955_/X _67003_/X _67004_/X sky130_fd_sc_hd__a211o_4
X_52230_ _52220_/A _48847_/B _52230_/Y sky130_fd_sc_hd__nand2_4
X_64216_ _64214_/Y _64186_/X _64215_/Y _64216_/Y sky130_fd_sc_hd__a21oi_4
X_83050_ _86498_/CLK _83050_/D _83050_/Q sky130_fd_sc_hd__dfxtp_4
X_61428_ _58535_/A _61428_/X sky130_fd_sc_hd__buf_2
X_80262_ _79902_/Y _80262_/B _80262_/X sky130_fd_sc_hd__xor2_4
X_65196_ _65196_/A _65268_/B _84211_/Q _65196_/X sky130_fd_sc_hd__and3_4
X_82001_ _82288_/CLK _82001_/D _77105_/A sky130_fd_sc_hd__dfxtp_4
X_52161_ _52161_/A _52140_/X _52182_/C _52161_/X sky130_fd_sc_hd__and3_4
X_64147_ _64142_/Y _64144_/Y _64145_/Y _64146_/Y _64147_/X sky130_fd_sc_hd__and4_4
X_61359_ _63389_/A _61368_/B _61368_/C _61368_/D _61359_/Y sky130_fd_sc_hd__nand4_4
X_80193_ _80187_/A _80186_/X _80192_/Y _80209_/A sky130_fd_sc_hd__a21boi_4
X_51112_ _51112_/A _52803_/B _51112_/Y sky130_fd_sc_hd__nand2_4
X_52092_ _85890_/Q _52089_/X _52091_/Y _52092_/Y sky130_fd_sc_hd__o21ai_4
X_64078_ _58393_/Y _61003_/Y _58490_/A _60962_/A _64078_/X sky130_fd_sc_hd__o22a_4
X_68955_ _68955_/A _68956_/B sky130_fd_sc_hd__inv_2
X_51043_ _51022_/A _51043_/B _51043_/Y sky130_fd_sc_hd__nand2_4
X_55920_ _56211_/C _44087_/B _44052_/A _55919_/X _55920_/X sky130_fd_sc_hd__a211o_4
X_67906_ _67550_/X _67906_/X sky130_fd_sc_hd__buf_2
X_63029_ _63039_/A _64236_/C _63028_/X _63014_/D _63029_/X sky130_fd_sc_hd__and4_4
X_86740_ _85527_/CLK _46409_/Y _86740_/Q sky130_fd_sc_hd__dfxtp_4
X_83952_ _80776_/CLK _83952_/D _80808_/D sky130_fd_sc_hd__dfxtp_4
X_68886_ _68669_/A _68886_/B _68886_/Y sky130_fd_sc_hd__nor2_4
X_82903_ _81783_/CLK _78231_/B _82903_/Q sky130_fd_sc_hd__dfxtp_4
X_55851_ _55477_/A _55851_/B _55851_/X sky130_fd_sc_hd__and2_4
X_67837_ _87390_/Q _67834_/X _67835_/X _67836_/X _67837_/X sky130_fd_sc_hd__a211o_4
X_86671_ _86353_/CLK _86671_/D _59226_/A sky130_fd_sc_hd__dfxtp_4
X_83883_ _82301_/CLK _83883_/D _83883_/Q sky130_fd_sc_hd__dfxtp_4
X_54802_ _54693_/X _54802_/X sky130_fd_sc_hd__buf_2
X_85622_ _86235_/CLK _53517_/Y _85622_/Q sky130_fd_sc_hd__dfxtp_4
X_58570_ _58085_/X _85473_/Q _58569_/X _58570_/Y sky130_fd_sc_hd__o21ai_4
X_82834_ _84119_/CLK _82834_/D _82834_/Q sky130_fd_sc_hd__dfxtp_4
X_55782_ _55781_/X _55801_/B sky130_fd_sc_hd__buf_2
X_67768_ _86957_/Q _67670_/X _67671_/X _67767_/X _67768_/X sky130_fd_sc_hd__a211o_4
X_52994_ _52992_/Y _52975_/X _52993_/X _52994_/Y sky130_fd_sc_hd__a21oi_4
X_57521_ _57531_/A _53488_/B _57521_/Y sky130_fd_sc_hd__nand2_4
X_69507_ _69580_/A _87768_/Q _69507_/X sky130_fd_sc_hd__and2_4
X_88341_ _88337_/CLK _88341_/D _88341_/Q sky130_fd_sc_hd__dfxtp_4
X_54733_ _85388_/Q _54729_/X _54732_/Y _54733_/Y sky130_fd_sc_hd__o21ai_4
X_66719_ _87129_/Q _66715_/X _66717_/X _66718_/X _66719_/X sky130_fd_sc_hd__a211o_4
X_85553_ _85553_/CLK _53864_/Y _85553_/Q sky130_fd_sc_hd__dfxtp_4
X_51945_ _52152_/A _51945_/X sky130_fd_sc_hd__buf_2
X_82765_ _82769_/CLK _82765_/D _82957_/D sky130_fd_sc_hd__dfxtp_4
X_67699_ _67222_/A _67793_/A sky130_fd_sc_hd__buf_2
X_84504_ _84493_/CLK _84504_/D _61223_/C sky130_fd_sc_hd__dfxtp_4
X_81716_ _81514_/CLK _81716_/D _41007_/B sky130_fd_sc_hd__dfxtp_4
X_57452_ _57452_/A _57452_/Y sky130_fd_sc_hd__inv_2
X_69438_ _70009_/A _69696_/A sky130_fd_sc_hd__buf_2
X_88272_ _88272_/CLK _41131_/X _88272_/Q sky130_fd_sc_hd__dfxtp_4
X_54664_ _54649_/X _47306_/A _54664_/Y sky130_fd_sc_hd__nand2_4
X_85484_ _85484_/CLK _85484_/D _85484_/Q sky130_fd_sc_hd__dfxtp_4
X_51876_ _85930_/Q _51873_/X _51875_/Y _51876_/Y sky130_fd_sc_hd__o21ai_4
X_82696_ _82933_/CLK _78862_/X _82684_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_61_0_CLK clkbuf_7_61_0_CLK/A clkbuf_7_61_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_56403_ _56397_/X _56399_/B _85207_/Q _56403_/Y sky130_fd_sc_hd__nand3_4
X_87223_ _88002_/CLK _43874_/X _69045_/B sky130_fd_sc_hd__dfxtp_4
X_53615_ _53613_/Y _53603_/X _53614_/Y _85602_/D sky130_fd_sc_hd__a21boi_4
X_84435_ _84438_/CLK _62080_/Y _78058_/B sky130_fd_sc_hd__dfxtp_4
X_50827_ _50822_/A _50827_/B _50827_/Y sky130_fd_sc_hd__nand2_4
X_57383_ _57465_/A _57484_/A sky130_fd_sc_hd__buf_2
X_81647_ _81361_/CLK _76917_/A _76330_/A sky130_fd_sc_hd__dfxtp_4
X_69369_ _69234_/A _87778_/Q _69369_/X sky130_fd_sc_hd__and2_4
X_54595_ _54594_/X _54600_/A sky130_fd_sc_hd__buf_2
X_59122_ _59048_/X _85655_/Q _59070_/X _59122_/X sky130_fd_sc_hd__o21a_4
X_71400_ _71397_/X _83513_/Q _71399_/Y _71400_/X sky130_fd_sc_hd__a21o_4
X_56334_ _56347_/A _56345_/A sky130_fd_sc_hd__buf_2
X_87154_ _87149_/CLK _87154_/D _87154_/Q sky130_fd_sc_hd__dfxtp_4
X_53546_ _53565_/A _50322_/B _53546_/Y sky130_fd_sc_hd__nand2_4
X_41560_ _41559_/Y _41560_/X sky130_fd_sc_hd__buf_2
X_72380_ _72371_/Y _72358_/X _72376_/X _72379_/X _83260_/D sky130_fd_sc_hd__a22oi_4
X_84366_ _84449_/CLK _84366_/D _84366_/Q sky130_fd_sc_hd__dfxtp_4
X_50758_ _86139_/Q _50742_/X _50757_/Y _50758_/Y sky130_fd_sc_hd__o21ai_4
X_81578_ _81344_/CLK _84178_/Q _76726_/A sky130_fd_sc_hd__dfxtp_4
X_86105_ _86104_/CLK _86105_/D _86105_/Q sky130_fd_sc_hd__dfxtp_4
X_40511_ _40507_/X _40508_/X _88380_/Q _40510_/X _88380_/D sky130_fd_sc_hd__a2bb2o_4
X_71331_ _71335_/A _71335_/B _71680_/C _71331_/Y sky130_fd_sc_hd__nand3_4
X_59053_ _59053_/A _59053_/X sky130_fd_sc_hd__buf_2
X_83317_ _85003_/CLK _71950_/Y _83317_/Q sky130_fd_sc_hd__dfxtp_4
X_80529_ _80551_/A _80529_/Y sky130_fd_sc_hd__inv_2
X_56265_ _56194_/X _56263_/B _85253_/Q _56265_/Y sky130_fd_sc_hd__nand3_4
X_41491_ _81179_/Q _41471_/B _41491_/X sky130_fd_sc_hd__or2_4
X_87085_ _88263_/CLK _44486_/Y _87085_/Q sky130_fd_sc_hd__dfxtp_4
X_53477_ _54919_/A _53478_/A sky130_fd_sc_hd__buf_2
X_84297_ _84293_/CLK _84297_/D _63745_/C sky130_fd_sc_hd__dfxtp_4
X_50689_ _50687_/Y _50644_/X _50688_/Y _86153_/D sky130_fd_sc_hd__a21boi_4
Xclkbuf_7_76_0_CLK clkbuf_7_77_0_CLK/A clkbuf_7_76_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_58004_ _57999_/Y _58001_/Y _58003_/X _58004_/X sky130_fd_sc_hd__a21o_4
X_43230_ _43226_/X _43229_/X _41004_/X _87527_/Q _43212_/X _43231_/A
+ sky130_fd_sc_hd__o32ai_4
X_55216_ _55741_/A _85122_/Q _55216_/X sky130_fd_sc_hd__and2_4
X_74050_ _70112_/C _73939_/X _74049_/X _74050_/Y sky130_fd_sc_hd__o21ai_4
X_86036_ _86040_/CLK _51303_/Y _86036_/Q sky130_fd_sc_hd__dfxtp_4
X_40442_ _40441_/Y _40442_/Y sky130_fd_sc_hd__inv_2
X_52428_ _52185_/X _53946_/B _52428_/Y sky130_fd_sc_hd__nand2_4
X_71262_ _50268_/B _71239_/A _71261_/Y _71262_/Y sky130_fd_sc_hd__o21ai_4
X_83248_ _83248_/CLK _83248_/D _83248_/Q sky130_fd_sc_hd__dfxtp_4
X_56196_ _56280_/A _56192_/B _56196_/C _56196_/Y sky130_fd_sc_hd__nand3_4
X_73001_ _42004_/Y _72921_/X _72944_/X _73000_/Y _73001_/X sky130_fd_sc_hd__a211o_4
X_70213_ _70209_/X _83835_/Q _70212_/X _83835_/D sky130_fd_sc_hd__a21o_4
X_55147_ _55139_/X _55146_/X _55147_/X sky130_fd_sc_hd__and2_4
X_43161_ _43161_/A _43162_/A sky130_fd_sc_hd__buf_2
X_40373_ _44624_/A _44532_/A sky130_fd_sc_hd__buf_2
X_71193_ _70984_/A _71217_/B sky130_fd_sc_hd__buf_2
X_52359_ _52319_/A _52385_/A sky130_fd_sc_hd__buf_2
X_83179_ _83820_/CLK _83179_/D _70260_/C sky130_fd_sc_hd__dfxtp_4
X_42112_ _42112_/A _42112_/Y sky130_fd_sc_hd__inv_2
X_70144_ _70144_/A _70144_/B _70144_/C _70144_/D _70144_/X sky130_fd_sc_hd__and4_4
X_43092_ _43072_/X _43075_/X _40724_/X _74123_/A _43080_/X _43092_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55078_ _55083_/A _55056_/X _55083_/C _55078_/D _55078_/X sky130_fd_sc_hd__and4_4
X_59955_ _60513_/A _61587_/B _84681_/Q _59955_/X sky130_fd_sc_hd__or3_4
X_87987_ _82317_/CLK _87987_/D _87987_/Q sky130_fd_sc_hd__dfxtp_4
X_46920_ _46920_/A _54442_/B sky130_fd_sc_hd__inv_2
X_42043_ _42024_/A _42043_/X sky130_fd_sc_hd__buf_2
X_58906_ _58891_/X _86087_/Q _58905_/X _58906_/Y sky130_fd_sc_hd__o21ai_4
X_54029_ _85519_/Q _54018_/X _54028_/Y _54029_/Y sky130_fd_sc_hd__o21ai_4
X_77740_ _77739_/Y _77742_/A sky130_fd_sc_hd__inv_2
X_74952_ _74958_/B _74961_/B _74952_/Y sky130_fd_sc_hd__nand2_4
X_70075_ _69603_/X _69902_/Y _70056_/X _70074_/Y _70075_/X sky130_fd_sc_hd__a211o_4
X_86938_ _83987_/CLK _44816_/Y _86938_/Q sky130_fd_sc_hd__dfxtp_4
X_59886_ _59615_/A _61277_/C sky130_fd_sc_hd__inv_2
X_73903_ _72909_/A _73903_/X sky130_fd_sc_hd__buf_2
X_46851_ _52713_/B _51022_/B sky130_fd_sc_hd__buf_2
X_58837_ _58835_/X _85452_/Q _58836_/X _58837_/Y sky130_fd_sc_hd__o21ai_4
X_77671_ _77671_/A _82206_/D _77671_/X sky130_fd_sc_hd__xor2_4
X_74883_ _74876_/Y _74881_/Y _74882_/Y _74887_/C sky130_fd_sc_hd__a21o_4
X_86869_ _86869_/CLK _86869_/D _63124_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_14_0_CLK clkbuf_6_7_0_CLK/X clkbuf_8_29_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_79410_ _79418_/A _79410_/B _82839_/D sky130_fd_sc_hd__xnor2_4
X_45802_ _74691_/B _45832_/B _45802_/Y sky130_fd_sc_hd__nand2_4
X_76622_ _76618_/X _76621_/X _76623_/A sky130_fd_sc_hd__xor2_4
X_49570_ _49570_/A _49570_/X sky130_fd_sc_hd__buf_2
X_73834_ _73786_/X _84982_/Q _73740_/X _73833_/X _73835_/B sky130_fd_sc_hd__a211o_4
X_46782_ _82960_/Q _54362_/D sky130_fd_sc_hd__inv_2
X_58768_ _58755_/Y _58739_/X _58762_/X _58767_/X _84802_/D sky130_fd_sc_hd__a22oi_4
Xclkbuf_8_154_0_CLK clkbuf_7_77_0_CLK/X clkbuf_8_154_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_43994_ _43994_/A _43995_/A sky130_fd_sc_hd__buf_2
X_48521_ _48471_/X _47982_/A _48520_/Y _48522_/A sky130_fd_sc_hd__o21ai_4
X_79341_ _79331_/A _79331_/B _79340_/Y _79341_/Y sky130_fd_sc_hd__a21boi_4
X_45733_ _57027_/A _45733_/Y sky130_fd_sc_hd__inv_2
X_57719_ _57707_/Y _57714_/Y _57718_/X _57719_/X sky130_fd_sc_hd__a21o_4
X_76553_ _76552_/Y _76554_/C sky130_fd_sc_hd__inv_2
X_42945_ _42945_/A _42945_/X sky130_fd_sc_hd__buf_2
X_73765_ _73765_/A _73765_/B _73765_/X sky130_fd_sc_hd__xor2_4
X_70977_ _46412_/B _70961_/A _70976_/Y _70977_/Y sky130_fd_sc_hd__o21ai_4
X_58699_ _58699_/A _58699_/B _58699_/Y sky130_fd_sc_hd__nor2_4
X_75504_ _75536_/A _75503_/Y _75504_/X sky130_fd_sc_hd__and2_4
X_48452_ _48752_/A _48489_/B _48476_/C _48452_/X sky130_fd_sc_hd__and3_4
X_72716_ _72714_/A _72714_/B _56907_/X _72716_/Y sky130_fd_sc_hd__nand3_4
X_60730_ _60632_/X _60624_/X _60731_/A sky130_fd_sc_hd__nor2_4
X_79272_ _79247_/X _79270_/X _79248_/Y _79271_/Y _79272_/Y sky130_fd_sc_hd__nand4_4
X_45664_ _45661_/X _45663_/Y _45602_/X _45664_/X sky130_fd_sc_hd__a21o_4
X_76484_ _76448_/B _76482_/X _76483_/Y _76484_/Y sky130_fd_sc_hd__a21oi_4
X_42876_ _42874_/X _42875_/X _41596_/X _67188_/B _42858_/X _42877_/A
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_9_270_0_CLK clkbuf_9_271_0_CLK/A clkbuf_9_270_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_73696_ _70125_/D _86754_/D _73695_/X _83140_/D sky130_fd_sc_hd__o21ai_4
Xclkbuf_7_29_0_CLK clkbuf_7_28_0_CLK/A clkbuf_8_59_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_47403_ _47403_/A _53025_/B sky130_fd_sc_hd__buf_2
X_78223_ _78222_/Y _78220_/C _78223_/X sky130_fd_sc_hd__and2_4
X_44615_ _44588_/X _44589_/X _40976_/X _87031_/Q _44590_/X _44616_/A
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_8_169_0_CLK clkbuf_7_84_0_CLK/X clkbuf_9_339_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_75435_ _75400_/X _75435_/B _75401_/Y _75435_/D _75436_/A sky130_fd_sc_hd__and4_4
X_41827_ _41826_/Y _88134_/D sky130_fd_sc_hd__inv_2
X_48383_ _48193_/X _48383_/X sky130_fd_sc_hd__buf_2
X_60661_ _60694_/B _60654_/X _60697_/B _60660_/X _60671_/A sky130_fd_sc_hd__nand4_4
X_72647_ _44231_/A _72656_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_164_0_CLK clkbuf_9_82_0_CLK/X _81671_/CLK sky130_fd_sc_hd__clkbuf_1
X_45595_ _45595_/A _45595_/Y sky130_fd_sc_hd__inv_2
X_62400_ _62471_/A _62431_/D sky130_fd_sc_hd__buf_2
X_47334_ _47334_/A _47334_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_794_0_CLK clkbuf_9_397_0_CLK/X _82589_/CLK sky130_fd_sc_hd__clkbuf_1
X_78154_ _78154_/A _78154_/B _78154_/X sky130_fd_sc_hd__or2_4
X_44546_ _44545_/Y _44546_/Y sky130_fd_sc_hd__inv_2
X_75366_ _75354_/X _75366_/Y sky130_fd_sc_hd__inv_2
X_63380_ _63380_/A _63389_/B _63418_/C _63389_/D _63380_/Y sky130_fd_sc_hd__nand4_4
X_41758_ _41753_/X _41754_/X _41757_/X _88155_/Q _41736_/X _41759_/A
+ sky130_fd_sc_hd__o32ai_4
X_72578_ _79385_/B _61252_/X _72570_/Y _72577_/Y _72578_/X sky130_fd_sc_hd__o22a_4
X_60592_ _60591_/X _84592_/D sky130_fd_sc_hd__inv_2
X_77105_ _77105_/A _81913_/Q _77112_/C sky130_fd_sc_hd__nand2_4
X_74317_ _74325_/A _74325_/B _74317_/C _74317_/Y sky130_fd_sc_hd__nand3_4
X_62331_ _62236_/A _62332_/B sky130_fd_sc_hd__buf_2
X_40709_ _40709_/A _40709_/Y sky130_fd_sc_hd__inv_2
X_47265_ _47246_/X _47228_/B _47234_/X _52948_/D _47265_/X sky130_fd_sc_hd__and4_4
Xclkbuf_9_285_0_CLK clkbuf_9_285_0_CLK/A clkbuf_9_285_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_71529_ _71528_/X _71137_/B _71530_/A sky130_fd_sc_hd__nor2_4
X_78085_ _78085_/A _78084_/X _78085_/Y sky130_fd_sc_hd__xnor2_4
X_44477_ _44447_/X _44448_/X _41192_/X _87088_/Q _44449_/X _44478_/A
+ sky130_fd_sc_hd__o32ai_4
X_75297_ _75297_/A _81041_/D _75297_/X sky130_fd_sc_hd__xor2_4
X_41689_ _41672_/X _41673_/X _41688_/X _67575_/B _41668_/X _41690_/A
+ sky130_fd_sc_hd__o32ai_4
X_49004_ _48898_/A _49007_/A sky130_fd_sc_hd__buf_2
X_46216_ _46216_/A _46216_/Y sky130_fd_sc_hd__inv_2
X_65050_ _64691_/X _86128_/Q _64972_/X _65049_/X _65050_/X sky130_fd_sc_hd__a211o_4
XPHY_280 sky130_fd_sc_hd__decap_3
X_77036_ _77036_/A _77036_/B _77036_/Y sky130_fd_sc_hd__nor2_4
X_43428_ _43428_/A _43428_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_179_0_CLK clkbuf_9_89_0_CLK/X _81284_/CLK sky130_fd_sc_hd__clkbuf_1
X_62262_ _61365_/X _62560_/B _62560_/C _62211_/D _62262_/Y sky130_fd_sc_hd__nand4_4
X_74248_ _74245_/X _74247_/X _72741_/X _74248_/X sky130_fd_sc_hd__a21o_4
XPHY_291 sky130_fd_sc_hd__decap_3
X_47196_ _47196_/A _47195_/X _47196_/Y sky130_fd_sc_hd__nand2_4
X_64001_ _63997_/Y _63998_/Y _63999_/Y _64001_/D _64001_/X sky130_fd_sc_hd__and4_4
X_61213_ _75909_/A _60719_/X _61208_/Y _61212_/Y _84507_/D sky130_fd_sc_hd__o22a_4
X_46147_ _49793_/A _49520_/A sky130_fd_sc_hd__buf_2
X_43359_ _41356_/X _43356_/X _87462_/Q _43357_/X _87462_/D sky130_fd_sc_hd__a2bb2o_4
Xpsn_inst_psn_buff_18 _44274_/D _56456_/A sky130_fd_sc_hd__buf_2
X_62193_ _62193_/A _62618_/D sky130_fd_sc_hd__buf_2
X_74179_ _74176_/X _74179_/B _74180_/B sky130_fd_sc_hd__nand2_4
Xpsn_inst_psn_buff_29 _50212_/A _50221_/A sky130_fd_sc_hd__buf_8
X_61144_ _61144_/A _64221_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_107_0_CLK clkbuf_7_53_0_CLK/X clkbuf_9_214_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_46078_ _46077_/Y _46078_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_102_0_CLK clkbuf_9_51_0_CLK/X _84534_/CLK sky130_fd_sc_hd__clkbuf_1
X_78987_ _78986_/X _78987_/Y sky130_fd_sc_hd__inv_2
X_49906_ _49906_/A _49906_/X sky130_fd_sc_hd__buf_2
X_45029_ _85209_/Q _45027_/X _45028_/X _45029_/Y sky130_fd_sc_hd__o21ai_4
X_68740_ _83963_/Q _68713_/X _68739_/X _83963_/D sky130_fd_sc_hd__a21bo_4
Xclkbuf_10_732_0_CLK clkbuf_9_366_0_CLK/X _87032_/CLK sky130_fd_sc_hd__clkbuf_1
X_65952_ _65924_/X _84990_/Q _65950_/X _65951_/X _65952_/X sky130_fd_sc_hd__a211o_4
X_61075_ _59639_/A _61075_/B _61075_/C _59552_/B _61075_/X sky130_fd_sc_hd__and4_4
X_77938_ _77927_/B _81944_/D sky130_fd_sc_hd__inv_2
X_64903_ _64903_/A _64904_/A sky130_fd_sc_hd__buf_2
X_60026_ _60025_/X _60027_/A sky130_fd_sc_hd__buf_2
X_49837_ _49827_/X _53050_/B _49837_/Y sky130_fd_sc_hd__nand2_4
X_68671_ _68386_/A _68746_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_223_0_CLK clkbuf_9_222_0_CLK/A clkbuf_9_223_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_65883_ _65824_/X _83051_/Q _65707_/X _65882_/X _65884_/B sky130_fd_sc_hd__a211o_4
X_77869_ _77869_/A _77868_/Y _82033_/D sky130_fd_sc_hd__xnor2_4
X_67622_ _86963_/Q _67551_/X _67552_/X _67621_/X _67623_/B sky130_fd_sc_hd__a211o_4
X_79608_ _79608_/A _79609_/A _79609_/B _79611_/A sky130_fd_sc_hd__nand3_4
X_64834_ _64834_/A _64888_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_117_0_CLK clkbuf_9_58_0_CLK/X _84906_/CLK sky130_fd_sc_hd__clkbuf_1
X_49768_ _49825_/A _49768_/X sky130_fd_sc_hd__buf_2
X_80880_ _80849_/CLK _75705_/B _80880_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_747_0_CLK clkbuf_9_373_0_CLK/X _87487_/CLK sky130_fd_sc_hd__clkbuf_1
X_48719_ _52103_/A _48099_/X _48723_/C _48719_/X sky130_fd_sc_hd__and3_4
X_67553_ _67575_/A _67553_/B _67553_/X sky130_fd_sc_hd__and2_4
X_79539_ _79538_/Y _64542_/A _79540_/C sky130_fd_sc_hd__nand2_4
X_64765_ _64762_/Y _64662_/X _64764_/Y _84228_/D sky130_fd_sc_hd__a21o_4
X_49699_ _49699_/A _51222_/B _49699_/Y sky130_fd_sc_hd__nand2_4
X_61977_ _62002_/A _62002_/B _78065_/B _61977_/Y sky130_fd_sc_hd__nor3_4
X_66504_ _66475_/X _66303_/Y _66503_/Y _66504_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_238_0_CLK clkbuf_9_239_0_CLK/A clkbuf_9_238_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_51730_ _51709_/X _51721_/X _51715_/C _53253_/D _51730_/X sky130_fd_sc_hd__and4_4
X_63716_ _61695_/A _63384_/D _60667_/Y _60758_/X _84882_/Q _63716_/X
+ sky130_fd_sc_hd__a32o_4
X_82550_ _82369_/CLK _82550_/D _78839_/B sky130_fd_sc_hd__dfxtp_4
X_60928_ _60928_/A _60928_/X sky130_fd_sc_hd__buf_2
X_67484_ _67484_/A _67483_/X _67484_/Y sky130_fd_sc_hd__nand2_4
X_64696_ _64696_/A _64696_/X sky130_fd_sc_hd__buf_2
X_81501_ _81428_/CLK _84069_/Q _76894_/A sky130_fd_sc_hd__dfxtp_4
X_69223_ _69223_/A _69253_/A sky130_fd_sc_hd__buf_2
X_66435_ _66435_/A _66435_/Y sky130_fd_sc_hd__inv_2
X_51661_ _85969_/Q _51647_/X _51660_/Y _51661_/Y sky130_fd_sc_hd__o21ai_4
X_63647_ _63642_/Y _63635_/X _63646_/Y _63647_/Y sky130_fd_sc_hd__a21oi_4
X_82481_ _82563_/CLK _82481_/D _78124_/B sky130_fd_sc_hd__dfxtp_4
X_60859_ _60915_/A _60865_/C sky130_fd_sc_hd__buf_2
X_53400_ _85640_/Q _53378_/X _53399_/Y _53400_/Y sky130_fd_sc_hd__o21ai_4
X_84220_ _84220_/CLK _64970_/X _84220_/Q sky130_fd_sc_hd__dfxtp_4
X_50612_ _50597_/A _48982_/X _50612_/Y sky130_fd_sc_hd__nand2_4
X_81432_ _81431_/CLK _81464_/Q _76075_/B sky130_fd_sc_hd__dfxtp_4
X_69154_ _69073_/A _88306_/Q _69154_/X sky130_fd_sc_hd__and2_4
X_54380_ _54395_/A _54362_/B _54395_/C _46809_/Y _54380_/X sky130_fd_sc_hd__and4_4
X_66366_ _66366_/A _66366_/X sky130_fd_sc_hd__buf_2
X_51592_ _51580_/A _51603_/B _51603_/C _53118_/D _51592_/X sky130_fd_sc_hd__and4_4
X_63578_ _63578_/A _63578_/X sky130_fd_sc_hd__buf_2
X_68105_ _67013_/X _68106_/A sky130_fd_sc_hd__buf_2
X_53331_ _53327_/Y _53328_/X _53330_/X _85654_/D sky130_fd_sc_hd__a21oi_4
X_65317_ _65314_/X _65316_/X _64701_/X _65317_/X sky130_fd_sc_hd__a21o_4
X_84151_ _81224_/CLK _84151_/D _84151_/Q sky130_fd_sc_hd__dfxtp_4
X_50543_ _48680_/A _50552_/B _50552_/C _50543_/X sky130_fd_sc_hd__and3_4
X_62529_ _62487_/X _83243_/Q _62628_/C _62219_/X _62529_/X sky130_fd_sc_hd__and4_4
X_81363_ _81811_/CLK _81363_/D _81363_/Q sky130_fd_sc_hd__dfxtp_4
X_69085_ _80804_/D _69066_/X _69084_/X _83948_/D sky130_fd_sc_hd__a21bo_4
X_66297_ _66266_/X _86214_/Q _66295_/X _66296_/X _66297_/X sky130_fd_sc_hd__a211o_4
X_83102_ _83095_/CLK _83102_/D _83102_/Q sky130_fd_sc_hd__dfxtp_4
X_56050_ _56049_/Y _56050_/X sky130_fd_sc_hd__buf_2
X_80314_ _84749_/Q _66319_/C _80314_/Y sky130_fd_sc_hd__nand2_4
X_68036_ _86946_/Q _67942_/X _67991_/X _68035_/X _68036_/X sky130_fd_sc_hd__a211o_4
X_53262_ _53260_/Y _53242_/X _53261_/X _53262_/Y sky130_fd_sc_hd__a21oi_4
X_65248_ _65199_/X _86152_/Q _65224_/X _65247_/X _65248_/X sky130_fd_sc_hd__a211o_4
X_84082_ _83933_/CLK _67140_/X _80906_/D sky130_fd_sc_hd__dfxtp_4
X_50474_ _50577_/A _50474_/X sky130_fd_sc_hd__buf_2
X_81294_ _81808_/CLK _76982_/X _81262_/D sky130_fd_sc_hd__dfxtp_4
X_55001_ _54997_/Y _54998_/X _55000_/X _55001_/Y sky130_fd_sc_hd__a21oi_4
X_52213_ _52211_/Y _52203_/X _52212_/X _52213_/Y sky130_fd_sc_hd__a21oi_4
X_87910_ _86930_/CLK _87910_/D _87910_/Q sky130_fd_sc_hd__dfxtp_4
X_83033_ _85241_/CLK _83033_/D _83033_/Q sky130_fd_sc_hd__dfxtp_4
X_80245_ _80213_/X _80216_/Y _80230_/Y _80233_/Y _80245_/X sky130_fd_sc_hd__o22a_4
X_53193_ _53187_/A _53193_/B _53193_/Y sky130_fd_sc_hd__nand2_4
X_65179_ _65164_/A _86411_/Q _65179_/X sky130_fd_sc_hd__and2_4
X_52144_ _85880_/Q _52125_/X _52143_/Y _52144_/Y sky130_fd_sc_hd__o21ai_4
X_87841_ _88097_/CLK _42508_/Y _87841_/Q sky130_fd_sc_hd__dfxtp_4
X_80176_ _80176_/A _80175_/X _80176_/Y sky130_fd_sc_hd__xnor2_4
X_69987_ _82559_/D _69955_/X _69986_/X _69987_/X sky130_fd_sc_hd__a21bo_4
X_59740_ _62717_/A _62669_/D sky130_fd_sc_hd__buf_2
X_52075_ _52438_/A _52075_/X sky130_fd_sc_hd__buf_2
X_56952_ _56952_/A _56952_/X sky130_fd_sc_hd__buf_2
X_68938_ _68938_/A _88348_/Q _68938_/X sky130_fd_sc_hd__and2_4
X_87772_ _87767_/CLK _42683_/X _69452_/B sky130_fd_sc_hd__dfxtp_4
X_84984_ _85915_/CLK _84984_/D _84984_/Q sky130_fd_sc_hd__dfxtp_4
X_51026_ _51022_/A _51026_/B _51026_/Y sky130_fd_sc_hd__nand2_4
X_55903_ _55903_/A _85241_/Q _55903_/X sky130_fd_sc_hd__and2_4
X_86723_ _86404_/CLK _46593_/Y _86723_/Q sky130_fd_sc_hd__dfxtp_4
X_59671_ _66046_/A _59696_/A sky130_fd_sc_hd__buf_2
X_83935_ _84087_/CLK _69284_/X _83935_/Q sky130_fd_sc_hd__dfxtp_4
X_56883_ _56866_/A _56859_/X _83334_/Q _56884_/C sky130_fd_sc_hd__a21o_4
X_68869_ _87999_/Q _68778_/X _68800_/X _68868_/X _68869_/X sky130_fd_sc_hd__a211o_4
X_70900_ _46805_/X _70885_/X _70899_/Y _70900_/Y sky130_fd_sc_hd__o21ai_4
X_58622_ _84813_/Q _58599_/X _58615_/X _58621_/X _84813_/D sky130_fd_sc_hd__a2bb2oi_4
X_55834_ _85201_/Q _55475_/X _55523_/X _55833_/X _55834_/X sky130_fd_sc_hd__a211o_4
X_86654_ _86655_/CLK _86654_/D _86654_/Q sky130_fd_sc_hd__dfxtp_4
X_71880_ _71871_/X _83343_/Q _71879_/Y _71880_/X sky130_fd_sc_hd__a21o_4
X_83866_ _82541_/CLK _83866_/D _83866_/Q sky130_fd_sc_hd__dfxtp_4
X_85605_ _85895_/CLK _85605_/D _85605_/Q sky130_fd_sc_hd__dfxtp_4
X_70831_ _70830_/Y _70831_/X sky130_fd_sc_hd__buf_2
X_58553_ _84820_/Q _58554_/A sky130_fd_sc_hd__inv_2
X_82817_ _82740_/CLK _82849_/Q _82817_/Q sky130_fd_sc_hd__dfxtp_4
X_55765_ _85257_/Q _55152_/X _44043_/X _55764_/X _55765_/X sky130_fd_sc_hd__a211o_4
X_86585_ _86587_/CLK _86585_/D _66024_/B sky130_fd_sc_hd__dfxtp_4
X_40991_ _40783_/A _40991_/X sky130_fd_sc_hd__buf_2
X_52977_ _52997_/A _52982_/B _52977_/C _52977_/D _52977_/X sky130_fd_sc_hd__and4_4
X_83797_ _81808_/CLK _83797_/D _74768_/B sky130_fd_sc_hd__dfxtp_4
X_57504_ _84990_/Q _47806_/X _57503_/Y _57504_/Y sky130_fd_sc_hd__o21ai_4
X_88324_ _88324_/CLK _88324_/D _88324_/Q sky130_fd_sc_hd__dfxtp_4
X_42730_ _41199_/X _42717_/X _68768_/B _42718_/X _42730_/X sky130_fd_sc_hd__a2bb2o_4
X_54716_ _54699_/X _54734_/B _54721_/C _47399_/A _54716_/X sky130_fd_sc_hd__and4_4
X_73550_ _74140_/A _74117_/A sky130_fd_sc_hd__buf_2
X_85536_ _85536_/CLK _53950_/Y _85536_/Q sky130_fd_sc_hd__dfxtp_4
X_51928_ _52126_/A _51928_/X sky130_fd_sc_hd__buf_2
X_70762_ DATA_TO_HASH[7] _70763_/A sky130_fd_sc_hd__buf_2
X_58484_ _58467_/X _58480_/Y _58483_/Y _84838_/D sky130_fd_sc_hd__a21oi_4
X_82748_ _82748_/CLK _79455_/B _82748_/Q sky130_fd_sc_hd__dfxtp_4
X_55696_ _85217_/Q _55690_/A _55611_/X _55695_/X _55696_/X sky130_fd_sc_hd__a211o_4
X_72501_ _46150_/B _83378_/Q _72500_/Y _83242_/D sky130_fd_sc_hd__o21a_4
X_57435_ _85004_/Q _57413_/X _57435_/X sky130_fd_sc_hd__or2_4
X_88255_ _87083_/CLK _41222_/Y _88255_/Q sky130_fd_sc_hd__dfxtp_4
X_54647_ _54034_/A _54729_/A sky130_fd_sc_hd__buf_2
X_42661_ _42647_/X _42648_/X _41009_/X _87782_/Q _42658_/X _42661_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73481_ _73479_/X _73481_/B _73481_/C _73481_/Y sky130_fd_sc_hd__nand3_4
X_85467_ _82206_/CLK _54304_/Y _85467_/Q sky130_fd_sc_hd__dfxtp_4
X_51859_ _51804_/A _51870_/A sky130_fd_sc_hd__buf_2
X_70693_ _70664_/A _47515_/A _70692_/Y _70693_/X sky130_fd_sc_hd__a21o_4
X_82679_ _81216_/CLK _82679_/D _78231_/A sky130_fd_sc_hd__dfxtp_4
X_44400_ _44400_/A _44400_/Y sky130_fd_sc_hd__inv_2
X_75220_ _75216_/Y _75219_/Y _81036_/D sky130_fd_sc_hd__xor2_4
X_87206_ _87149_/CLK _43906_/X _67644_/B sky130_fd_sc_hd__dfxtp_4
X_41612_ _40637_/A _41825_/A sky130_fd_sc_hd__buf_2
X_72432_ _72389_/X _85671_/Q _72422_/X _72432_/X sky130_fd_sc_hd__o21a_4
X_84418_ _84418_/CLK _84418_/D _62328_/C sky130_fd_sc_hd__dfxtp_4
X_45380_ _45380_/A _45381_/A sky130_fd_sc_hd__inv_2
X_57366_ _57244_/X _45856_/Y _57366_/Y sky130_fd_sc_hd__nand2_4
X_88186_ _87110_/CLK _41593_/X _88186_/Q sky130_fd_sc_hd__dfxtp_4
X_42592_ _42592_/A _42592_/X sky130_fd_sc_hd__buf_2
X_54578_ _54578_/A _54578_/B _54578_/Y sky130_fd_sc_hd__nand2_4
X_85398_ _85492_/CLK _54681_/Y _85398_/Q sky130_fd_sc_hd__dfxtp_4
X_59105_ _58846_/A _59105_/X sky130_fd_sc_hd__buf_2
X_44331_ _44382_/A _44331_/X sky130_fd_sc_hd__buf_2
X_56317_ _56309_/A _56312_/X _56317_/C _56317_/Y sky130_fd_sc_hd__nand3_4
X_75151_ _80680_/Q _75151_/B _75151_/Y sky130_fd_sc_hd__nor2_4
X_87137_ _87137_/CLK _44385_/Y _87137_/Q sky130_fd_sc_hd__dfxtp_4
X_41543_ _41604_/A _82321_/Q _41543_/X sky130_fd_sc_hd__or2_4
X_53529_ _53503_/X _48257_/B _53529_/Y sky130_fd_sc_hd__nand2_4
X_72363_ _72361_/X _85677_/Q _72362_/X _72363_/X sky130_fd_sc_hd__o21a_4
X_84349_ _84350_/CLK _84349_/D _79385_/A sky130_fd_sc_hd__dfxtp_4
X_57297_ _57296_/Y _57290_/X _45888_/A _57297_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_4_11_0_CLK clkbuf_3_5_1_CLK/X clkbuf_4_11_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_74102_ _74102_/A _74102_/B _74102_/Y sky130_fd_sc_hd__nand2_4
X_47050_ _47004_/A _47050_/X sky130_fd_sc_hd__buf_2
X_59036_ _59036_/A _59037_/A sky130_fd_sc_hd__buf_2
X_71314_ _71500_/A _71314_/B _71313_/X _71314_/Y sky130_fd_sc_hd__nand3_4
X_44262_ _64717_/A _64725_/A sky130_fd_sc_hd__buf_2
X_56248_ _56250_/A _56253_/B _85260_/Q _56248_/Y sky130_fd_sc_hd__nand3_4
X_75082_ _80675_/Q _75082_/B _75082_/X sky130_fd_sc_hd__or2_4
X_87068_ _87068_/CLK _87068_/D _87068_/Q sky130_fd_sc_hd__dfxtp_4
X_41474_ _41235_/X _41474_/X sky130_fd_sc_hd__buf_2
X_72294_ _72366_/A _72294_/B _72294_/Y sky130_fd_sc_hd__nor2_4
X_46001_ _46001_/A _46001_/X sky130_fd_sc_hd__buf_2
X_43213_ _43196_/X _43207_/X _40959_/X _87535_/Q _43212_/X _43214_/A
+ sky130_fd_sc_hd__o32ai_4
X_78910_ _82638_/Q _78912_/A sky130_fd_sc_hd__inv_2
X_86019_ _85953_/CLK _51393_/Y _86019_/Q sky130_fd_sc_hd__dfxtp_4
X_74033_ _74033_/A _73873_/B _74033_/Y sky130_fd_sc_hd__nor2_4
X_40425_ _40421_/X _81175_/Q _40424_/X _40425_/X sky130_fd_sc_hd__o21a_4
X_71245_ _70809_/A _71246_/B sky130_fd_sc_hd__buf_2
X_44193_ _72745_/A _73948_/A sky130_fd_sc_hd__buf_2
X_56179_ _44187_/A _73378_/A sky130_fd_sc_hd__buf_2
X_79890_ _79890_/A _79890_/B _79890_/Y sky130_fd_sc_hd__nand2_4
X_43144_ _43100_/X _43110_/X _40826_/X _73083_/A _43121_/X _43145_/A
+ sky130_fd_sc_hd__o32ai_4
X_78841_ _78833_/Y _78841_/B _78841_/Y sky130_fd_sc_hd__nand2_4
X_40356_ _40331_/X _40342_/X _88402_/Q _40355_/X _88402_/D sky130_fd_sc_hd__a2bb2o_4
X_71176_ _48482_/B _71165_/X _71175_/Y _71176_/Y sky130_fd_sc_hd__o21ai_4
X_70127_ _70118_/Y _70119_/Y _70127_/C _70127_/D _70127_/X sky130_fd_sc_hd__and4_4
X_47952_ _47988_/A _48236_/B _47952_/Y sky130_fd_sc_hd__nand2_4
X_43075_ _43017_/A _43075_/X sky130_fd_sc_hd__buf_2
X_59938_ _59887_/Y _59892_/Y _60165_/A _59881_/X _59884_/X _59938_/Y
+ sky130_fd_sc_hd__a32oi_4
X_78772_ _78772_/A _78746_/Y _78780_/A sky130_fd_sc_hd__or2_4
X_75984_ _81706_/D _75972_/B _75984_/Y sky130_fd_sc_hd__nand2_4
X_46903_ _46903_/A _46926_/C sky130_fd_sc_hd__buf_2
X_42026_ _42013_/X _42024_/X _40854_/X _73196_/A _42025_/X _42027_/A
+ sky130_fd_sc_hd__o32ai_4
X_77723_ _77723_/A _77721_/A _77723_/C _77724_/B sky130_fd_sc_hd__nand3_4
Xclkbuf_10_1004_0_CLK clkbuf_9_502_0_CLK/X _85590_/CLK sky130_fd_sc_hd__clkbuf_1
X_74935_ _74935_/A _74935_/B _81191_/D sky130_fd_sc_hd__xor2_4
X_70058_ _70040_/X _69844_/Y _70056_/X _70057_/Y _70058_/X sky130_fd_sc_hd__a211o_4
X_47883_ _86589_/Q _47840_/X _47882_/Y _47883_/Y sky130_fd_sc_hd__o21ai_4
X_59869_ _59850_/Y _59789_/Y _59724_/Y _59866_/Y _59868_/X _59869_/Y
+ sky130_fd_sc_hd__a32oi_4
X_49622_ _86353_/Q _49606_/X _49621_/Y _49622_/Y sky130_fd_sc_hd__o21ai_4
X_61900_ _61896_/Y _61881_/X _61899_/Y _61900_/Y sky130_fd_sc_hd__a21oi_4
X_46834_ _46817_/A _51008_/B _46834_/Y sky130_fd_sc_hd__nand2_4
X_77654_ _77653_/Y _77654_/Y sky130_fd_sc_hd__inv_2
X_62880_ _62847_/X _63230_/A _62911_/C _62880_/D _62880_/X sky130_fd_sc_hd__and4_4
X_74866_ _74860_/Y _74865_/Y _74856_/Y _74866_/Y sky130_fd_sc_hd__a21oi_4
X_76605_ _76583_/Y _76616_/B _76614_/C _76605_/X sky130_fd_sc_hd__o21a_4
X_49553_ _49580_/A _49558_/A sky130_fd_sc_hd__buf_2
X_61831_ _84723_/Q _61831_/X sky130_fd_sc_hd__buf_2
X_73817_ _70102_/A _73697_/X _73816_/X _83135_/D sky130_fd_sc_hd__o21ai_4
X_46765_ _46760_/Y _46751_/X _46764_/X _86706_/D sky130_fd_sc_hd__a21oi_4
X_77585_ _77584_/B _77584_/C _77584_/A _77585_/Y sky130_fd_sc_hd__o21ai_4
X_43977_ _43973_/X _43976_/X _80669_/Q _59899_/B sky130_fd_sc_hd__a21o_4
X_74797_ _74797_/A _74804_/A _74797_/C _71738_/X _74798_/D sky130_fd_sc_hd__nand4_4
X_48504_ _74428_/B _52163_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_1019_0_CLK clkbuf_9_509_0_CLK/X _85859_/CLK sky130_fd_sc_hd__clkbuf_1
X_79324_ _79324_/A _79324_/B _79324_/X sky130_fd_sc_hd__or2_4
X_45716_ _63241_/B _61572_/A sky130_fd_sc_hd__buf_2
X_64550_ _64543_/Y _64549_/X _60074_/X _64550_/Y sky130_fd_sc_hd__o21ai_4
X_76536_ _76535_/B _76534_/Y _76531_/Y _76540_/C sky130_fd_sc_hd__o21ai_4
X_42928_ _42927_/Y _87647_/D sky130_fd_sc_hd__inv_2
X_49484_ _49482_/Y _49460_/X _49483_/X _86379_/D sky130_fd_sc_hd__a21oi_4
X_61762_ _59456_/A _61762_/X sky130_fd_sc_hd__buf_2
X_73748_ _73746_/X _73747_/Y _73720_/X _73748_/X sky130_fd_sc_hd__a21o_4
X_46696_ _46696_/A _54312_/D sky130_fd_sc_hd__inv_2
X_63501_ _63375_/A _63512_/A sky130_fd_sc_hd__buf_2
X_60713_ _60713_/A _63417_/A sky130_fd_sc_hd__buf_2
X_48435_ _48469_/A _48435_/B _48435_/Y sky130_fd_sc_hd__nand2_4
X_79255_ _84792_/Q _66495_/C _79255_/Y sky130_fd_sc_hd__nand2_4
X_45647_ _45647_/A _45647_/Y sky130_fd_sc_hd__inv_2
X_76467_ _76448_/B _76482_/C _76482_/A _76468_/B sky130_fd_sc_hd__a21boi_4
X_64481_ _64490_/A _64490_/B _79637_/B _64481_/Y sky130_fd_sc_hd__nor3_4
X_42859_ _42847_/X _42849_/X _41545_/X _66959_/B _42858_/X _42860_/A
+ sky130_fd_sc_hd__o32ai_4
X_61693_ _84730_/Q _61694_/B sky130_fd_sc_hd__buf_2
X_73679_ _72951_/A _73679_/X sky130_fd_sc_hd__buf_2
X_66220_ _66181_/A _85899_/Q _66220_/X sky130_fd_sc_hd__and2_4
X_78206_ _78198_/A _82491_/Q _78206_/Y sky130_fd_sc_hd__nor2_4
X_63432_ _63456_/A _63456_/B _80568_/B _63432_/Y sky130_fd_sc_hd__nor3_4
X_75418_ _75413_/X _75416_/Y _75414_/Y _75435_/D sky130_fd_sc_hd__nand3_4
X_48366_ _48360_/Y _48302_/X _48365_/X _86529_/D sky130_fd_sc_hd__a21oi_4
X_60644_ _60642_/C _60616_/Y _60644_/C _60644_/X sky130_fd_sc_hd__and3_4
X_79186_ _79185_/B _79185_/C _79186_/Y sky130_fd_sc_hd__nand2_4
X_45578_ _63137_/B _61468_/A sky130_fd_sc_hd__buf_2
X_76398_ _76398_/A _81651_/Q _76399_/A sky130_fd_sc_hd__nand2_4
X_47317_ _47128_/A _47317_/X sky130_fd_sc_hd__buf_2
X_66151_ _66123_/A _66151_/B _84153_/Q _66151_/X sky130_fd_sc_hd__and3_4
X_78137_ _78131_/Y _78136_/X _78137_/Y sky130_fd_sc_hd__nand2_4
X_44529_ _44529_/A _44529_/X sky130_fd_sc_hd__buf_2
X_63363_ _63363_/A _63363_/X sky130_fd_sc_hd__buf_2
X_75349_ _80693_/Q _80949_/D _75349_/Y sky130_fd_sc_hd__nor2_4
X_60575_ _60570_/X _60571_/Y _60546_/A _60572_/X _60574_/X _60575_/X
+ sky130_fd_sc_hd__o41a_4
X_48297_ _48058_/B _48297_/X sky130_fd_sc_hd__buf_2
X_65102_ _65102_/A _65102_/B _65102_/Y sky130_fd_sc_hd__nand2_4
X_62314_ _62218_/A _62315_/C sky130_fd_sc_hd__buf_2
X_47248_ _54630_/D _52938_/D sky130_fd_sc_hd__buf_2
X_66082_ _65763_/A _66082_/B _66082_/X sky130_fd_sc_hd__and2_4
X_78068_ _84573_/Q _78068_/B _78068_/X sky130_fd_sc_hd__xor2_4
X_63294_ _63247_/A _63344_/D sky130_fd_sc_hd__buf_2
X_65033_ _64999_/X _86161_/Q _64927_/X _65032_/X _65033_/X sky130_fd_sc_hd__a211o_4
X_69910_ _69907_/X _69909_/X _66579_/X _69910_/X sky130_fd_sc_hd__a21o_4
X_77019_ _77019_/A _77019_/Y sky130_fd_sc_hd__inv_2
X_62245_ _62478_/A _59995_/A _64235_/B _60025_/X _62245_/X sky130_fd_sc_hd__and4_4
X_47179_ _82374_/Q _47180_/A sky130_fd_sc_hd__inv_2
X_80030_ _80030_/A _80030_/Y sky130_fd_sc_hd__inv_2
X_69841_ _69755_/A _69900_/A sky130_fd_sc_hd__buf_2
X_50190_ _48759_/A _51263_/A sky130_fd_sc_hd__buf_2
X_62176_ _61715_/A _62172_/Y _62173_/Y _62175_/Y _62176_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_10_671_0_CLK clkbuf_9_335_0_CLK/X _88394_/CLK sky130_fd_sc_hd__clkbuf_1
X_61127_ _61122_/B _61122_/C _61122_/A _61128_/A sky130_fd_sc_hd__a21oi_4
X_69772_ _69772_/A _69772_/B _69772_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_162_0_CLK clkbuf_8_81_0_CLK/X clkbuf_9_162_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_66984_ _66628_/X _66984_/X sky130_fd_sc_hd__buf_2
X_68723_ _68938_/A _68723_/B _68723_/X sky130_fd_sc_hd__and2_4
X_65935_ _65934_/X _65935_/B _65935_/X sky130_fd_sc_hd__and2_4
X_61058_ _60950_/Y _60963_/X _60935_/X _61025_/X _61057_/X _61058_/X
+ sky130_fd_sc_hd__o41a_4
X_81981_ _83906_/CLK _81981_/D _81981_/Q sky130_fd_sc_hd__dfxtp_4
X_52900_ _52895_/A _52879_/B _52900_/C _52900_/D _52900_/X sky130_fd_sc_hd__and4_4
X_60009_ _59938_/Y _60079_/B _60009_/Y sky130_fd_sc_hd__nand2_4
X_83720_ _85439_/CLK _70711_/Y _46928_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_686_0_CLK clkbuf_9_343_0_CLK/X _87708_/CLK sky130_fd_sc_hd__clkbuf_1
X_68654_ _68604_/A _87240_/Q _68654_/X sky130_fd_sc_hd__and2_4
X_80932_ _81933_/CLK _80932_/D _80932_/Q sky130_fd_sc_hd__dfxtp_4
X_53880_ _53878_/Y _53862_/X _53879_/Y _85550_/D sky130_fd_sc_hd__a21boi_4
X_65866_ _65812_/A _86500_/Q _65866_/X sky130_fd_sc_hd__and2_4
X_67605_ _67582_/A _67605_/B _67605_/X sky130_fd_sc_hd__and2_4
X_52831_ _52818_/A _52831_/B _52818_/C _52831_/D _52831_/X sky130_fd_sc_hd__and4_4
X_64817_ _64817_/A _64817_/X sky130_fd_sc_hd__buf_2
X_83651_ _85822_/CLK _70955_/Y _83651_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_177_0_CLK clkbuf_8_88_0_CLK/X clkbuf_9_177_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_80863_ _83967_/CLK _80895_/Q _75062_/B sky130_fd_sc_hd__dfxtp_4
X_68585_ _80825_/D _68462_/X _68584_/X _68585_/X sky130_fd_sc_hd__a21bo_4
X_65797_ _65812_/A _86505_/Q _65797_/X sky130_fd_sc_hd__and2_4
X_82602_ _82570_/CLK _78882_/B _82602_/Q sky130_fd_sc_hd__dfxtp_4
X_55550_ _45526_/A _55505_/X _55532_/X _55549_/X _55550_/X sky130_fd_sc_hd__a211o_4
X_67536_ _67513_/A _67536_/B _67536_/X sky130_fd_sc_hd__and2_4
X_86370_ _83660_/CLK _86370_/D _58957_/B sky130_fd_sc_hd__dfxtp_4
X_52762_ _52708_/A _52775_/C sky130_fd_sc_hd__buf_2
X_64748_ _64602_/A _64810_/A sky130_fd_sc_hd__buf_2
X_83582_ _86516_/CLK _71176_/Y _83582_/Q sky130_fd_sc_hd__dfxtp_4
X_80794_ _80821_/CLK _75786_/X _80794_/Q sky130_fd_sc_hd__dfxtp_4
X_54501_ _85430_/Q _54485_/X _54500_/Y _54501_/Y sky130_fd_sc_hd__o21ai_4
X_85321_ _85351_/CLK _85321_/D _85321_/Q sky130_fd_sc_hd__dfxtp_4
X_51713_ _85959_/Q _51701_/X _51712_/Y _51713_/Y sky130_fd_sc_hd__o21ai_4
X_82533_ _82532_/CLK _83853_/Q _82533_/Q sky130_fd_sc_hd__dfxtp_4
X_55481_ _55470_/A _55481_/B _55481_/Y sky130_fd_sc_hd__nor2_4
X_67467_ _67466_/X _67467_/X sky130_fd_sc_hd__buf_2
X_52693_ _85772_/Q _52684_/X _52692_/Y _52693_/Y sky130_fd_sc_hd__o21ai_4
X_64679_ _64679_/A _64679_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_100_0_CLK clkbuf_8_50_0_CLK/X clkbuf_9_100_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_57220_ _56645_/Y _56878_/Y _57221_/A _57220_/Y sky130_fd_sc_hd__a21oi_4
X_69206_ _69755_/A _69206_/B _69206_/X sky130_fd_sc_hd__and2_4
X_88040_ _88044_/CLK _88040_/D _88040_/Q sky130_fd_sc_hd__dfxtp_4
X_54432_ _54322_/A _54446_/A sky130_fd_sc_hd__buf_2
X_66418_ _66411_/X _66061_/Y _66417_/Y _66418_/Y sky130_fd_sc_hd__o21ai_4
X_85252_ _85156_/CLK _56268_/Y _56267_/C sky130_fd_sc_hd__dfxtp_4
X_51644_ _85972_/Q _51621_/X _51643_/Y _51644_/Y sky130_fd_sc_hd__o21ai_4
X_82464_ _82820_/CLK _79156_/X _82464_/Q sky130_fd_sc_hd__dfxtp_4
X_67398_ _67039_/X _67398_/X sky130_fd_sc_hd__buf_2
X_84203_ _84194_/CLK _84203_/D _84203_/Q sky130_fd_sc_hd__dfxtp_4
X_57151_ _56727_/X _57133_/X _57150_/Y _57151_/Y sky130_fd_sc_hd__o21ai_4
X_81415_ _81575_/CLK _81447_/Q _75957_/B sky130_fd_sc_hd__dfxtp_4
X_69137_ _87539_/Q _69098_/X _69124_/X _69136_/X _69137_/X sky130_fd_sc_hd__a211o_4
X_54363_ _54361_/Y _54338_/X _54362_/X _85456_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_624_0_CLK clkbuf_9_312_0_CLK/X _83967_/CLK sky130_fd_sc_hd__clkbuf_1
X_66349_ _65976_/A _66349_/X sky130_fd_sc_hd__buf_2
X_85183_ _85184_/CLK _56473_/Y _85183_/Q sky130_fd_sc_hd__dfxtp_4
X_51575_ _51580_/A _51580_/B _51553_/C _53103_/D _51575_/X sky130_fd_sc_hd__and4_4
X_82395_ _82965_/CLK _82395_/D _82395_/Q sky130_fd_sc_hd__dfxtp_4
X_56102_ _55994_/X _56102_/B _56102_/X sky130_fd_sc_hd__xor2_4
X_53314_ _53298_/A _47006_/Y _53314_/Y sky130_fd_sc_hd__nand2_4
X_84134_ _84166_/CLK _84134_/D _84134_/Q sky130_fd_sc_hd__dfxtp_4
X_50526_ _48845_/A _50526_/B _50526_/C _50526_/X sky130_fd_sc_hd__and3_4
X_57082_ _85091_/Q _57084_/A _57080_/X _57081_/Y _85091_/D sky130_fd_sc_hd__a211o_4
X_81346_ _81346_/CLK _76965_/Y _81346_/Q sky130_fd_sc_hd__dfxtp_4
X_69068_ _43103_/A _68883_/X _68741_/X _69067_/X _69068_/X sky130_fd_sc_hd__a211o_4
X_54294_ _54320_/A _54294_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_115_0_CLK clkbuf_8_57_0_CLK/X clkbuf_9_115_0_CLK/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_9_42_0_CLK clkbuf_9_43_0_CLK/A clkbuf_9_42_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_56033_ _56029_/X _56031_/X _56032_/Y _56033_/Y sky130_fd_sc_hd__o21ai_4
X_68019_ _87894_/Q _67950_/X _67997_/X _68018_/X _68019_/X sky130_fd_sc_hd__a211o_4
X_53245_ _53241_/Y _53242_/X _53244_/X _53245_/Y sky130_fd_sc_hd__a21oi_4
X_84065_ _81749_/CLK _84065_/D _84065_/Q sky130_fd_sc_hd__dfxtp_4
X_50457_ _50454_/Y _50455_/X _50456_/X _50457_/Y sky130_fd_sc_hd__a21oi_4
X_81277_ _81627_/CLK _81277_/D _76552_/A sky130_fd_sc_hd__dfxtp_4
X_71030_ _71175_/A _71030_/B _71030_/C _71018_/D _71030_/Y sky130_fd_sc_hd__nand4_4
X_83016_ _83016_/CLK _83016_/D _45290_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_639_0_CLK clkbuf_9_319_0_CLK/X _82103_/CLK sky130_fd_sc_hd__clkbuf_1
X_80228_ _80228_/A _80227_/Y _80228_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_3_0_0_CLK clkbuf_2_0_2_CLK/X clkbuf_3_0_1_CLK/A sky130_fd_sc_hd__clkbuf_1
X_41190_ _41189_/X _41181_/X _68723_/B _41182_/X _88261_/D sky130_fd_sc_hd__a2bb2o_4
X_53176_ _53097_/X _53181_/B sky130_fd_sc_hd__buf_2
X_50388_ _50500_/A _50481_/A sky130_fd_sc_hd__buf_2
X_52127_ _52215_/A _52127_/X sky130_fd_sc_hd__buf_2
X_87824_ _87824_/CLK _42551_/Y _42550_/A sky130_fd_sc_hd__dfxtp_4
X_80159_ _80145_/Y _80142_/X _80159_/X sky130_fd_sc_hd__and2_4
X_57984_ _57884_/X _85486_/Q _57923_/X _57984_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_9_57_0_CLK clkbuf_9_57_0_CLK/A clkbuf_9_57_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_59723_ _59721_/X _59722_/X _59724_/A sky130_fd_sc_hd__and2_4
X_52058_ _52058_/A _50356_/B _52058_/Y sky130_fd_sc_hd__nand2_4
X_56935_ _56934_/X _56935_/X sky130_fd_sc_hd__buf_2
X_87755_ _87757_/CLK _87755_/D _87755_/Q sky130_fd_sc_hd__dfxtp_4
X_72981_ _43135_/Y _72978_/X _72979_/X _72980_/Y _72981_/X sky130_fd_sc_hd__a211o_4
X_84967_ _86535_/CLK _57624_/Y _84967_/Q sky130_fd_sc_hd__dfxtp_4
X_51009_ _86090_/Q _50992_/X _51008_/Y _51009_/Y sky130_fd_sc_hd__o21ai_4
X_43900_ _43895_/X _43876_/X _41341_/X _87209_/Q _43897_/X _43901_/A
+ sky130_fd_sc_hd__o32ai_4
X_74720_ _70620_/D _74720_/B _74720_/C _74804_/D _74720_/X sky130_fd_sc_hd__and4_4
X_86706_ _86384_/CLK _86706_/D _86706_/Q sky130_fd_sc_hd__dfxtp_4
X_71932_ _71894_/Y _71945_/D sky130_fd_sc_hd__buf_2
X_83918_ _83918_/CLK _83918_/D _81382_/D sky130_fd_sc_hd__dfxtp_4
X_59654_ _66064_/A _59654_/X sky130_fd_sc_hd__buf_2
X_44880_ _45827_/B _44880_/X sky130_fd_sc_hd__buf_2
X_56866_ _56866_/A _83334_/Q _56859_/X _56884_/B sky130_fd_sc_hd__nand3_4
X_87686_ _87686_/CLK _87686_/D _66876_/B sky130_fd_sc_hd__dfxtp_4
X_84898_ _84732_/CLK _84898_/D _84898_/Q sky130_fd_sc_hd__dfxtp_4
X_58605_ _58605_/A _58605_/X sky130_fd_sc_hd__buf_2
X_43831_ _41147_/X _43817_/X _68530_/B _43818_/X _87245_/D sky130_fd_sc_hd__a2bb2o_4
X_55817_ _55817_/A _55817_/B _55817_/X sky130_fd_sc_hd__and2_4
X_74651_ _56626_/A _74641_/X _74650_/Y _82999_/D sky130_fd_sc_hd__a21boi_4
X_86637_ _86637_/CLK _86637_/D _86637_/Q sky130_fd_sc_hd__dfxtp_4
X_71863_ _71863_/A _71867_/B _70884_/B _71711_/A _71863_/Y sky130_fd_sc_hd__nor4_4
X_59585_ _59585_/A _59775_/A sky130_fd_sc_hd__inv_2
X_83849_ _83842_/CLK _83849_/D _83849_/Q sky130_fd_sc_hd__dfxtp_4
X_56797_ _56797_/A _56796_/Y _56798_/A sky130_fd_sc_hd__nand2_4
X_73602_ _72861_/X _73602_/X sky130_fd_sc_hd__buf_2
X_70814_ _70810_/A _70947_/B _70810_/C _70814_/Y sky130_fd_sc_hd__nand3_4
X_46550_ _46525_/X _49148_/A _46549_/X _51372_/B sky130_fd_sc_hd__o21ai_4
X_58536_ _58535_/Y _58498_/B _58536_/Y sky130_fd_sc_hd__nand2_4
X_77370_ _77369_/X _77396_/B sky130_fd_sc_hd__inv_2
X_55748_ _55794_/A _55748_/B _55748_/X sky130_fd_sc_hd__and2_4
X_43762_ _43762_/A _43762_/Y sky130_fd_sc_hd__inv_2
X_74582_ _74549_/Y _74582_/X sky130_fd_sc_hd__buf_2
X_86568_ _85599_/CLK _48101_/Y _86568_/Q sky130_fd_sc_hd__dfxtp_4
X_40974_ _40973_/Y _40974_/Y sky130_fd_sc_hd__inv_2
X_71794_ _70804_/A _71680_/C _71785_/X _71794_/Y sky130_fd_sc_hd__nand3_4
X_45501_ _45501_/A _45456_/X _45501_/Y sky130_fd_sc_hd__nor2_4
X_76321_ _76321_/A _76320_/Y _76321_/Y sky130_fd_sc_hd__nand2_4
X_88307_ _87851_/CLK _40936_/X _88307_/Q sky130_fd_sc_hd__dfxtp_4
X_42713_ _41151_/X _42710_/X _68543_/B _42711_/X _42713_/X sky130_fd_sc_hd__a2bb2o_4
X_85519_ _86127_/CLK _54032_/Y _85519_/Q sky130_fd_sc_hd__dfxtp_4
X_73533_ _69972_/B _73026_/X _73421_/X _73533_/Y sky130_fd_sc_hd__o21ai_4
X_46481_ _48461_/A _47915_/B sky130_fd_sc_hd__buf_2
X_70745_ _70753_/A _70714_/A _70745_/Y sky130_fd_sc_hd__nand2_4
X_58467_ _58341_/A _58467_/X sky130_fd_sc_hd__buf_2
X_43693_ _40814_/A _43659_/X _69700_/B _43661_/X _43693_/X sky130_fd_sc_hd__a2bb2o_4
X_55679_ _55669_/A _55289_/X _55678_/X _55680_/B sky130_fd_sc_hd__a21boi_4
X_86499_ _86499_/CLK _48703_/Y _86499_/Q sky130_fd_sc_hd__dfxtp_4
X_48220_ _66028_/B _48203_/X _48219_/Y _48220_/Y sky130_fd_sc_hd__o21ai_4
X_79040_ _82828_/Q _82540_/Q _82524_/D sky130_fd_sc_hd__xor2_4
X_45432_ _45431_/Y _45590_/B _45432_/X sky130_fd_sc_hd__and2_4
X_57418_ _57417_/Y _85008_/D sky130_fd_sc_hd__inv_2
X_76252_ _76230_/Y _76232_/A _76233_/C _76252_/Y sky130_fd_sc_hd__o21ai_4
X_88238_ _87472_/CLK _88238_/D _67456_/B sky130_fd_sc_hd__dfxtp_4
X_42644_ _40968_/X _42631_/X _69218_/B _42634_/X _87789_/D sky130_fd_sc_hd__a2bb2o_4
X_73464_ _56934_/X _73464_/X sky130_fd_sc_hd__buf_2
X_70676_ _70676_/A _70676_/B _70676_/C _70676_/Y sky130_fd_sc_hd__nor3_4
X_58398_ _58388_/X _83347_/Q _58397_/Y _58398_/X sky130_fd_sc_hd__o21a_4
X_75203_ _75186_/A _75186_/B _75202_/Y _75203_/Y sky130_fd_sc_hd__a21boi_4
X_72415_ _72414_/X _72415_/B _72415_/Y sky130_fd_sc_hd__nor2_4
X_48151_ _48731_/A _48725_/A sky130_fd_sc_hd__buf_2
X_45363_ _85283_/Q _45343_/X _45303_/X _45363_/X sky130_fd_sc_hd__o21a_4
X_57349_ _56824_/X _57349_/B _57349_/Y sky130_fd_sc_hd__nand2_4
X_76183_ _76168_/B _76182_/Y _76183_/Y sky130_fd_sc_hd__xnor2_4
X_88169_ _87188_/CLK _41690_/Y _67575_/B sky130_fd_sc_hd__dfxtp_4
X_42575_ _42573_/X _42574_/X _40826_/X _87815_/Q _42540_/X _42576_/A
+ sky130_fd_sc_hd__o32ai_4
X_73395_ _42047_/Y _72974_/X _73393_/X _73394_/Y _73395_/X sky130_fd_sc_hd__a211o_4
X_47102_ _46961_/X _47113_/A sky130_fd_sc_hd__buf_2
X_44314_ _44312_/Y _44313_/Y _44318_/A _44314_/Y sky130_fd_sc_hd__a21oi_4
X_75134_ _75120_/B _75134_/Y sky130_fd_sc_hd__inv_2
X_41526_ _41525_/X _41486_/X _88198_/Q _41487_/X _88198_/D sky130_fd_sc_hd__a2bb2o_4
X_48082_ _48081_/Y _48310_/B sky130_fd_sc_hd__buf_2
X_60360_ _60168_/A _60177_/X _60360_/X sky130_fd_sc_hd__and2_4
X_72346_ _83263_/Q _72250_/X _72338_/X _72345_/X _83263_/D sky130_fd_sc_hd__a2bb2oi_4
X_45294_ _45219_/A _45294_/X sky130_fd_sc_hd__buf_2
X_47033_ _47008_/A _52813_/B _47033_/Y sky130_fd_sc_hd__nand2_4
X_59019_ _59019_/A _59008_/B _59019_/Y sky130_fd_sc_hd__nor2_4
X_44245_ _44245_/A _44246_/A sky130_fd_sc_hd__buf_2
X_75065_ _75067_/B _75067_/A _75066_/B sky130_fd_sc_hd__xor2_4
X_79942_ _79942_/A _79940_/Y _79941_/Y _79945_/B sky130_fd_sc_hd__nand3_4
X_41457_ _41457_/A _41457_/X sky130_fd_sc_hd__buf_2
X_60291_ _60233_/Y _60251_/A _60291_/C _60292_/A sky130_fd_sc_hd__nand3_4
X_72277_ _72277_/A _72277_/B _72277_/Y sky130_fd_sc_hd__nor2_4
X_62030_ _62142_/A _62025_/Y _62026_/Y _62030_/D _62030_/Y sky130_fd_sc_hd__nand4_4
X_74016_ _73378_/A _74016_/X sky130_fd_sc_hd__buf_2
X_40408_ _40407_/Y _40408_/X sky130_fd_sc_hd__buf_2
X_71228_ _71232_/A _71228_/B _71232_/C _71228_/Y sky130_fd_sc_hd__nand3_4
X_44176_ _64679_/A _58126_/A sky130_fd_sc_hd__buf_2
X_79873_ _79871_/X _79873_/B _79873_/Y sky130_fd_sc_hd__xnor2_4
X_41388_ _41235_/X _41388_/X sky130_fd_sc_hd__buf_2
X_43127_ _43127_/A _43127_/X sky130_fd_sc_hd__buf_2
X_78824_ _82836_/Q _78825_/A _78828_/A sky130_fd_sc_hd__or2_4
X_40339_ _46259_/A _44362_/A sky130_fd_sc_hd__inv_2
X_71159_ _71225_/A _71173_/B sky130_fd_sc_hd__buf_2
X_48984_ _86455_/Q _48952_/X _48983_/Y _48984_/Y sky130_fd_sc_hd__o21ai_4
X_47935_ _82360_/Q _47963_/B _47935_/X sky130_fd_sc_hd__or2_4
X_43058_ _43058_/A _43058_/X sky130_fd_sc_hd__buf_2
X_78755_ _78732_/A _78732_/B _78731_/A _78755_/X sky130_fd_sc_hd__o21a_4
X_75967_ _75976_/A _75976_/B _75970_/A sky130_fd_sc_hd__xor2_4
X_63981_ _64392_/B _64029_/B _63951_/C _64015_/D _63981_/Y sky130_fd_sc_hd__nand4_4
X_42009_ _42009_/A _42009_/Y sky130_fd_sc_hd__inv_2
X_65720_ _65717_/X _85582_/Q _65718_/X _65719_/X _65720_/X sky130_fd_sc_hd__a211o_4
X_77706_ _77703_/Y _77710_/A _77707_/A sky130_fd_sc_hd__nand2_4
X_74918_ _74914_/Y _74917_/X _74930_/A sky130_fd_sc_hd__nand2_4
X_62932_ _60199_/X _62979_/D sky130_fd_sc_hd__buf_2
X_47866_ _73638_/B _47840_/X _47865_/Y _47866_/Y sky130_fd_sc_hd__o21ai_4
X_78686_ _78675_/B _78667_/X _78669_/B _78686_/Y sky130_fd_sc_hd__a21boi_4
X_75898_ _75898_/A _62943_/C _75898_/X sky130_fd_sc_hd__xor2_4
X_49605_ _49002_/A _49632_/A sky130_fd_sc_hd__buf_2
X_46817_ _46817_/A _50998_/B _46817_/Y sky130_fd_sc_hd__nand2_4
X_65651_ _65634_/A _65802_/B _65651_/C _65651_/Y sky130_fd_sc_hd__nor3_4
X_77637_ _77633_/X _77634_/Y _77636_/Y _77666_/B sky130_fd_sc_hd__a21oi_4
X_62863_ _62856_/X _62831_/X _62857_/Y _62860_/Y _62862_/X _62863_/X
+ sky130_fd_sc_hd__a41o_4
X_74849_ _80930_/Q _74849_/B _74849_/X sky130_fd_sc_hd__xor2_4
X_47797_ _47797_/A _47798_/A sky130_fd_sc_hd__inv_2
X_64602_ _64602_/A _64684_/A sky130_fd_sc_hd__buf_2
X_61814_ _61863_/A _61809_/Y _61810_/Y _61813_/Y _61814_/Y sky130_fd_sc_hd__nand4_4
X_49536_ _86369_/Q _49524_/X _49535_/Y _49536_/Y sky130_fd_sc_hd__o21ai_4
X_68370_ _68370_/A _68370_/X sky130_fd_sc_hd__buf_2
X_46748_ _52651_/B _50961_/B sky130_fd_sc_hd__buf_2
X_65582_ _65579_/X _65581_/X _65389_/X _65582_/X sky130_fd_sc_hd__a21o_4
X_77568_ _77568_/A _82105_/D _77568_/Y sky130_fd_sc_hd__nand2_4
X_62794_ _62792_/X _62839_/B _75912_/B _62794_/Y sky130_fd_sc_hd__nor3_4
X_79307_ _84797_/Q _66469_/C _79307_/Y sky130_fd_sc_hd__nand2_4
X_67321_ _87412_/Q _67274_/X _67226_/X _67320_/X _67321_/X sky130_fd_sc_hd__a211o_4
X_64533_ _58364_/A _64521_/X _64533_/Y sky130_fd_sc_hd__nor2_4
X_76519_ _76501_/Y _76502_/Y _76503_/Y _76519_/X sky130_fd_sc_hd__o21a_4
X_49467_ _49467_/A _49456_/B _49467_/C _52681_/D _49467_/X sky130_fd_sc_hd__and4_4
X_61745_ _61712_/X _61749_/B sky130_fd_sc_hd__buf_2
X_46679_ _74509_/B _46717_/A sky130_fd_sc_hd__buf_2
X_77499_ _77446_/A _77447_/X _77458_/B _77499_/X sky130_fd_sc_hd__a21o_4
X_48418_ _48413_/Y _48403_/X _48417_/Y _86524_/D sky130_fd_sc_hd__a21boi_4
X_67252_ _67249_/X _67251_/X _67204_/X _67252_/X sky130_fd_sc_hd__a21o_4
X_79238_ _79238_/A _79239_/A _79238_/Y sky130_fd_sc_hd__nand2_4
X_64464_ _58461_/A _64511_/B _64464_/Y sky130_fd_sc_hd__nor2_4
X_61676_ _61676_/A _61653_/X _61654_/X _61639_/X _61676_/Y sky130_fd_sc_hd__nand4_4
X_49398_ _49395_/Y _49378_/X _49397_/X _86395_/D sky130_fd_sc_hd__a21oi_4
X_66203_ _66200_/X _64633_/B _66203_/C _66203_/Y sky130_fd_sc_hd__nand3_4
X_63415_ _61375_/B _60834_/X _63412_/X _63414_/X _63415_/X sky130_fd_sc_hd__a211o_4
X_48349_ _48346_/Y _48322_/X _48348_/Y _86531_/D sky130_fd_sc_hd__a21boi_4
X_60627_ _60627_/A _60628_/C sky130_fd_sc_hd__inv_2
X_67183_ _67183_/A _67183_/B _67183_/X sky130_fd_sc_hd__and2_4
X_79169_ _79169_/A _79169_/B _79171_/B sky130_fd_sc_hd__nand2_4
X_64395_ _58338_/Y _64367_/X _64394_/Y _64395_/Y sky130_fd_sc_hd__o21ai_4
X_81200_ _82284_/CLK _74998_/X _46446_/A sky130_fd_sc_hd__dfxtp_4
X_66134_ _66134_/A _66133_/X _66134_/Y sky130_fd_sc_hd__nand2_4
X_51360_ _51306_/X _51360_/B _51360_/X sky130_fd_sc_hd__and2_4
X_63346_ _63338_/Y _63310_/X _63345_/X _63346_/Y sky130_fd_sc_hd__o21ai_4
X_82180_ _84951_/CLK _82180_/D _82180_/Q sky130_fd_sc_hd__dfxtp_4
X_60558_ _65515_/A _60558_/X sky130_fd_sc_hd__buf_2
X_50311_ _86225_/Q _50238_/X _50310_/Y _50311_/Y sky130_fd_sc_hd__o21ai_4
X_81131_ _80792_/CLK _81131_/D _40710_/A sky130_fd_sc_hd__dfxtp_4
X_66065_ _66065_/A _66065_/X sky130_fd_sc_hd__buf_2
X_51291_ _51288_/Y _51289_/X _51290_/X _86039_/D sky130_fd_sc_hd__a21oi_4
X_63277_ _63275_/X _62987_/X _63276_/Y _84338_/D sky130_fd_sc_hd__a21oi_4
X_60489_ _60588_/A _60489_/X sky130_fd_sc_hd__buf_2
X_65016_ _64836_/A _86450_/Q _65016_/X sky130_fd_sc_hd__and2_4
X_53030_ _53112_/A _53048_/A sky130_fd_sc_hd__buf_2
X_50242_ _50473_/A _50768_/A sky130_fd_sc_hd__buf_2
X_62228_ _62532_/A _62319_/C sky130_fd_sc_hd__buf_2
X_81062_ _81061_/CLK _81094_/Q _81062_/Q sky130_fd_sc_hd__dfxtp_4
X_80013_ _80011_/Y _79992_/Y _80012_/X _80013_/Y sky130_fd_sc_hd__o21ai_4
X_69824_ _73252_/A _68377_/X _66574_/X _69823_/Y _69824_/X sky130_fd_sc_hd__a211o_4
X_50173_ _50169_/A _49125_/X _50173_/Y sky130_fd_sc_hd__nand2_4
X_62159_ _58207_/A _62105_/X _62065_/D _62055_/A _62158_/X _62159_/X
+ sky130_fd_sc_hd__a41o_4
X_85870_ _86500_/CLK _85870_/D _85870_/Q sky130_fd_sc_hd__dfxtp_4
X_84821_ _84823_/CLK _84821_/D _84821_/Q sky130_fd_sc_hd__dfxtp_4
X_69755_ _69755_/A _69770_/A sky130_fd_sc_hd__buf_2
X_54981_ _54985_/A _47561_/Y _54981_/Y sky130_fd_sc_hd__nand2_4
X_66967_ _87119_/Q _66868_/X _66919_/X _66966_/X _66967_/X sky130_fd_sc_hd__a211o_4
X_56720_ _56682_/X _56721_/A sky130_fd_sc_hd__inv_2
X_68706_ _68703_/X _68705_/X _68684_/X _68706_/X sky130_fd_sc_hd__a21o_4
X_87540_ _87824_/CLK _43204_/Y _87540_/Q sky130_fd_sc_hd__dfxtp_4
X_53932_ _53951_/A _53932_/B _53932_/Y sky130_fd_sc_hd__nand2_4
X_65918_ _65446_/A _66195_/B _65445_/X _65928_/A sky130_fd_sc_hd__nand3_4
X_84752_ _86665_/CLK _84752_/D _84752_/Q sky130_fd_sc_hd__dfxtp_4
X_69686_ _43137_/A _69645_/X _68613_/X _69685_/X _69686_/X sky130_fd_sc_hd__a211o_4
X_81964_ _87345_/CLK _81964_/D _81964_/Q sky130_fd_sc_hd__dfxtp_4
X_66898_ _69156_/A _66898_/X sky130_fd_sc_hd__buf_2
X_83703_ _83703_/CLK _70776_/Y _47087_/A sky130_fd_sc_hd__dfxtp_4
X_56651_ _83337_/Q _83336_/Q _56651_/Y sky130_fd_sc_hd__nand2_4
X_80915_ _81507_/CLK _80915_/D _80915_/Q sky130_fd_sc_hd__dfxtp_4
X_68637_ _68637_/A _69086_/A sky130_fd_sc_hd__buf_2
X_87471_ _87471_/CLK _43340_/X _87471_/Q sky130_fd_sc_hd__dfxtp_4
X_53863_ _53863_/A _53821_/B _53863_/Y sky130_fd_sc_hd__nand2_4
X_65849_ _65717_/X _85573_/Q _65718_/X _65848_/X _65849_/X sky130_fd_sc_hd__a211o_4
X_84683_ _84713_/CLK _59871_/Y _80277_/B sky130_fd_sc_hd__dfxtp_4
X_81895_ _82015_/CLK _81895_/D _77217_/B sky130_fd_sc_hd__dfxtp_4
X_55602_ _55601_/X _72641_/C sky130_fd_sc_hd__buf_2
X_86422_ _86422_/CLK _49264_/Y _86422_/Q sky130_fd_sc_hd__dfxtp_4
X_52814_ _85749_/Q _52792_/X _52813_/Y _52814_/Y sky130_fd_sc_hd__o21ai_4
X_59370_ _59368_/X _86051_/Q _59369_/X _59370_/Y sky130_fd_sc_hd__o21ai_4
X_83634_ _85514_/CLK _71009_/Y _83634_/Q sky130_fd_sc_hd__dfxtp_4
X_56582_ _56582_/A _55552_/X _55570_/D _72648_/C _56583_/B sky130_fd_sc_hd__nand4_4
X_80846_ _80792_/CLK _80878_/Q _74928_/B sky130_fd_sc_hd__dfxtp_4
X_68568_ _41914_/A _68069_/X _68439_/X _68567_/Y _68568_/X sky130_fd_sc_hd__a211o_4
X_53794_ _53825_/A _71970_/B _53794_/Y sky130_fd_sc_hd__nand2_4
X_58321_ _58310_/X _83455_/Q _58320_/Y _84879_/D sky130_fd_sc_hd__o21a_4
X_55533_ _55532_/X _55533_/X sky130_fd_sc_hd__buf_2
X_67519_ _67515_/X _67518_/X _67401_/X _67519_/Y sky130_fd_sc_hd__a21oi_4
X_86353_ _86353_/CLK _86353_/D _86353_/Q sky130_fd_sc_hd__dfxtp_4
X_52745_ _85762_/Q _52737_/X _52744_/Y _52745_/Y sky130_fd_sc_hd__o21ai_4
X_83565_ _83311_/CLK _71229_/Y _48671_/A sky130_fd_sc_hd__dfxtp_4
X_80777_ _80776_/CLK _75629_/X _80777_/Q sky130_fd_sc_hd__dfxtp_4
X_68499_ _87002_/Q _68394_/X _68421_/X _68498_/X _68499_/X sky130_fd_sc_hd__a211o_4
X_85304_ _85241_/CLK _56057_/Y _55915_/B sky130_fd_sc_hd__dfxtp_4
X_70530_ _71823_/A _70700_/A _70700_/B _70530_/Y sky130_fd_sc_hd__nand3_4
X_58252_ _58171_/X _83449_/Q _58251_/Y _58252_/X sky130_fd_sc_hd__o21a_4
X_82516_ _82532_/CLK _82516_/D _78582_/A sky130_fd_sc_hd__dfxtp_4
X_55464_ _55826_/A _85140_/Q _55464_/X sky130_fd_sc_hd__and2_4
X_86284_ _86282_/CLK _86284_/D _72377_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_563_0_CLK clkbuf_9_281_0_CLK/X _88121_/CLK sky130_fd_sc_hd__clkbuf_1
X_40690_ _40577_/X _82863_/Q _40689_/X _40691_/A sky130_fd_sc_hd__o21a_4
X_52676_ _52672_/Y _52673_/X _52675_/X _52676_/Y sky130_fd_sc_hd__a21oi_4
X_83496_ _83495_/CLK _83496_/D _58151_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_6_54_0_CLK clkbuf_6_55_0_CLK/A clkbuf_6_54_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_57203_ _57203_/A _85064_/D sky130_fd_sc_hd__inv_2
X_88023_ _87273_/CLK _42127_/X _88023_/Q sky130_fd_sc_hd__dfxtp_4
X_54415_ _54425_/A _52722_/B _54415_/Y sky130_fd_sc_hd__nand2_4
X_85235_ _85168_/CLK _85235_/D _55855_/B sky130_fd_sc_hd__dfxtp_4
X_51627_ _51627_/A _53153_/B _51627_/Y sky130_fd_sc_hd__nand2_4
X_70461_ _71462_/B _71483_/B sky130_fd_sc_hd__buf_2
X_58183_ _57665_/A _58184_/B sky130_fd_sc_hd__buf_2
X_82447_ _82822_/CLK _79139_/X _82447_/Q sky130_fd_sc_hd__dfxtp_4
X_55395_ _55296_/A _55293_/X _55162_/Y _55296_/B _55396_/B sky130_fd_sc_hd__and4_4
X_72200_ _59381_/X _85979_/Q _72199_/X _72200_/Y sky130_fd_sc_hd__o21ai_4
X_57134_ _57133_/X _57134_/Y sky130_fd_sc_hd__inv_2
X_42360_ _42360_/A _42360_/Y sky130_fd_sc_hd__inv_2
X_54346_ _54317_/A _54362_/C sky130_fd_sc_hd__buf_2
X_73180_ _73173_/Y _73174_/Y _73179_/X _73180_/Y sky130_fd_sc_hd__o21ai_4
X_85166_ _85198_/CLK _85166_/D _55814_/B sky130_fd_sc_hd__dfxtp_4
X_51558_ _51504_/A _51580_/B sky130_fd_sc_hd__buf_2
X_70392_ _70944_/A _70942_/A sky130_fd_sc_hd__buf_2
X_82378_ _86054_/CLK _82186_/Q _82378_/Q sky130_fd_sc_hd__dfxtp_4
X_41311_ _41290_/X _82908_/Q _41310_/X _41311_/Y sky130_fd_sc_hd__o21ai_4
X_72131_ _59346_/X _85344_/Q _72120_/X _72131_/X sky130_fd_sc_hd__o21a_4
X_84117_ _84111_/CLK _84117_/D _66469_/C sky130_fd_sc_hd__dfxtp_4
X_50509_ _86187_/Q _50506_/X _50508_/Y _50509_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_578_0_CLK clkbuf_9_289_0_CLK/X _80754_/CLK sky130_fd_sc_hd__clkbuf_1
X_81329_ _81492_/CLK _76375_/X _75976_/A sky130_fd_sc_hd__dfxtp_4
X_57065_ _56966_/X _57063_/Y _57064_/Y _57065_/X sky130_fd_sc_hd__a21o_4
X_42291_ _42259_/A _42291_/X sky130_fd_sc_hd__buf_2
X_54277_ _54288_/A _54277_/B _54277_/Y sky130_fd_sc_hd__nand2_4
X_85097_ _85096_/CLK _85097_/D _57039_/A sky130_fd_sc_hd__dfxtp_4
X_51489_ _51473_/A _51494_/B _51494_/C _53015_/D _51489_/X sky130_fd_sc_hd__and4_4
X_44030_ _57848_/A _72255_/A sky130_fd_sc_hd__buf_2
X_56016_ _56016_/A _56016_/X sky130_fd_sc_hd__buf_2
X_41242_ _41072_/X _41242_/X sky130_fd_sc_hd__buf_2
X_53228_ _85673_/Q _53225_/X _53227_/Y _53228_/Y sky130_fd_sc_hd__o21ai_4
X_72062_ _72040_/A _53886_/B _72062_/Y sky130_fd_sc_hd__nand2_4
X_84048_ _88116_/CLK _67947_/X _84048_/Q sky130_fd_sc_hd__dfxtp_4
X_71013_ _71013_/A _71013_/X sky130_fd_sc_hd__buf_2
X_53159_ _53139_/A _53159_/B _53143_/X _53159_/D _53159_/X sky130_fd_sc_hd__and4_4
X_41173_ _41136_/X _40654_/A _41172_/X _41173_/X sky130_fd_sc_hd__o21a_4
X_76870_ _76866_/Y _76854_/B _76869_/Y _76870_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_501_0_CLK clkbuf_9_250_0_CLK/X _85778_/CLK sky130_fd_sc_hd__clkbuf_1
X_75821_ _75821_/A _75821_/B _75823_/C sky130_fd_sc_hd__nor2_4
X_87807_ _87553_/CLK _42599_/Y _87807_/Q sky130_fd_sc_hd__dfxtp_4
X_45981_ _43756_/A _45981_/X sky130_fd_sc_hd__buf_2
X_57967_ _57966_/X _85712_/Q _57878_/X _57967_/X sky130_fd_sc_hd__o21a_4
X_85999_ _85712_/CLK _85999_/D _85999_/Q sky130_fd_sc_hd__dfxtp_4
X_47720_ _49379_/A _47758_/A sky130_fd_sc_hd__buf_2
X_59706_ _59705_/X _63001_/A sky130_fd_sc_hd__buf_2
X_78540_ _78503_/Y _78505_/X _78528_/X _78540_/X sky130_fd_sc_hd__a21bo_4
X_44932_ _44932_/A _45252_/A sky130_fd_sc_hd__buf_2
X_56918_ _56877_/X _57193_/D sky130_fd_sc_hd__buf_2
X_75752_ _75735_/A _75747_/A _75752_/X sky130_fd_sc_hd__and2_4
X_87738_ _88002_/CLK _42753_/X _68977_/B sky130_fd_sc_hd__dfxtp_4
X_72964_ _72816_/X _86522_/Q _72964_/X sky130_fd_sc_hd__and2_4
X_57898_ _86645_/Q _57845_/X _57898_/Y sky130_fd_sc_hd__nor2_4
X_74703_ _74642_/X _56917_/A _74702_/Y _74704_/A sky130_fd_sc_hd__o21ai_4
X_47651_ _47745_/A _47651_/X sky130_fd_sc_hd__buf_2
X_71915_ _71912_/Y _56922_/X _71914_/Y _71915_/X sky130_fd_sc_hd__a21o_4
X_59637_ _59637_/A _59648_/A _59806_/A _59638_/A sky130_fd_sc_hd__nor3_4
Xclkbuf_10_516_0_CLK clkbuf_9_258_0_CLK/X _83926_/CLK sky130_fd_sc_hd__clkbuf_1
X_78471_ _82798_/Q _78473_/A sky130_fd_sc_hd__inv_2
X_44863_ _44857_/X _44844_/X _41785_/X _68054_/B _44858_/X _44863_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56849_ _56676_/Y _56849_/X sky130_fd_sc_hd__buf_2
X_75683_ _80909_/Q _80781_/D _75682_/X _75684_/B sky130_fd_sc_hd__o21ai_4
X_87669_ _87671_/CLK _87669_/D _67294_/B sky130_fd_sc_hd__dfxtp_4
X_72895_ _72894_/X _72895_/X sky130_fd_sc_hd__buf_2
X_46602_ _54091_/A _51396_/A sky130_fd_sc_hd__buf_2
X_77422_ _77422_/A _77422_/Y sky130_fd_sc_hd__inv_2
X_43814_ _41093_/X _43801_/X _69523_/B _43802_/X _87255_/D sky130_fd_sc_hd__a2bb2o_4
X_74634_ _45952_/X _56570_/Y _45416_/A _74633_/X _83008_/D sky130_fd_sc_hd__a2bb2o_4
X_47582_ _47582_/A _53131_/B sky130_fd_sc_hd__buf_2
X_71846_ _71846_/A _70882_/Y _70500_/D _71846_/Y sky130_fd_sc_hd__nor3_4
X_59568_ _59546_/A _43998_/A _59560_/A _59568_/X sky130_fd_sc_hd__and3_4
X_44794_ _44794_/A _86952_/D sky130_fd_sc_hd__inv_2
X_49321_ _86410_/Q _49285_/X _49320_/Y _49321_/Y sky130_fd_sc_hd__o21ai_4
X_46533_ _83784_/Q _52545_/B sky130_fd_sc_hd__inv_2
X_58519_ _84829_/Q _58520_/A sky130_fd_sc_hd__buf_2
X_77353_ _77353_/A _82091_/D _77354_/B sky130_fd_sc_hd__xor2_4
X_43745_ _40913_/X _47846_/A _69932_/B _43607_/A _43745_/X sky130_fd_sc_hd__a2bb2o_4
X_74565_ _56050_/X _74625_/A _74564_/Y _83033_/D sky130_fd_sc_hd__a21boi_4
X_40957_ _82301_/Q _40970_/B _40957_/X sky130_fd_sc_hd__or2_4
X_71777_ _71779_/A _71777_/B _70986_/A _71777_/X sky130_fd_sc_hd__and3_4
X_59499_ _46179_/X _63424_/B _59498_/Y _84716_/D sky130_fd_sc_hd__o21a_4
X_76304_ _76300_/Y _76301_/Y _76303_/Y _76306_/A sky130_fd_sc_hd__or3_4
X_61530_ _61317_/A _61563_/C sky130_fd_sc_hd__buf_2
X_49252_ _86424_/Q _49222_/X _49251_/Y _49252_/Y sky130_fd_sc_hd__o21ai_4
X_73516_ _73516_/A _86467_/Q _73516_/X sky130_fd_sc_hd__and2_4
X_70728_ _52787_/B _70699_/A _70727_/Y _70728_/Y sky130_fd_sc_hd__o21ai_4
X_46464_ _83638_/Q _46464_/Y sky130_fd_sc_hd__inv_2
X_77284_ _77280_/X _77285_/C _77285_/A _77287_/A sky130_fd_sc_hd__a21oi_4
X_43676_ _40762_/A _43659_/X _69114_/B _43661_/X _43677_/A sky130_fd_sc_hd__a2bb2o_4
X_74496_ _83054_/Q _74474_/X _74495_/Y _74496_/Y sky130_fd_sc_hd__o21ai_4
X_40888_ _40888_/A _40623_/X _40888_/X sky130_fd_sc_hd__or2_4
X_48203_ _48169_/X _48203_/X sky130_fd_sc_hd__buf_2
X_79023_ _79014_/B _79023_/Y sky130_fd_sc_hd__inv_2
X_45415_ _45410_/X _45414_/X _45361_/X _45415_/X sky130_fd_sc_hd__a21o_4
X_76235_ _76234_/Y _76215_/A _76216_/Y _76235_/Y sky130_fd_sc_hd__o21ai_4
X_42627_ _42626_/X _52274_/A sky130_fd_sc_hd__buf_2
X_49183_ _49178_/Y _49138_/X _49182_/X _49183_/Y sky130_fd_sc_hd__a21oi_4
X_61461_ _58546_/A _61461_/X sky130_fd_sc_hd__buf_2
X_73447_ _73495_/A _85862_/Q _73447_/X sky130_fd_sc_hd__and2_4
X_46395_ _52484_/B _46396_/B sky130_fd_sc_hd__buf_2
X_70659_ _53050_/B _70631_/X _70658_/Y _70659_/Y sky130_fd_sc_hd__o21ai_4
X_63200_ _79343_/A _63189_/X _63199_/Y _63200_/X sky130_fd_sc_hd__a21o_4
X_48134_ _48914_/A _48134_/X sky130_fd_sc_hd__buf_2
X_60412_ _63060_/A _60412_/X sky130_fd_sc_hd__buf_2
X_45346_ _45272_/A _45381_/B sky130_fd_sc_hd__buf_2
X_64180_ _58210_/X _64192_/C _64180_/C _64192_/D _64181_/D sky130_fd_sc_hd__nand4_4
X_76166_ _76160_/X _76161_/Y _76165_/X _76166_/X sky130_fd_sc_hd__a21o_4
X_61392_ _61392_/A _61392_/Y sky130_fd_sc_hd__inv_2
X_42558_ _87821_/Q _42558_/Y sky130_fd_sc_hd__inv_2
X_73378_ _73378_/A _73378_/X sky130_fd_sc_hd__buf_2
X_63131_ _63010_/A _63131_/X sky130_fd_sc_hd__buf_2
X_75117_ _75117_/A _75117_/B _75117_/C _75120_/B sky130_fd_sc_hd__nand3_4
X_41509_ _81175_/Q _41523_/B _41509_/X sky130_fd_sc_hd__or2_4
X_72329_ _72327_/X _85968_/Q _72328_/X _72329_/Y sky130_fd_sc_hd__o21ai_4
X_48065_ _48065_/A _47915_/B _48065_/Y sky130_fd_sc_hd__nand2_4
X_60343_ _60344_/A _60331_/B _60268_/A _60343_/Y sky130_fd_sc_hd__nand3_4
X_45277_ _45350_/A _45277_/X sky130_fd_sc_hd__buf_2
X_76097_ _76096_/Y _76097_/B _76097_/Y sky130_fd_sc_hd__nand2_4
X_42489_ _42556_/A _42489_/X sky130_fd_sc_hd__buf_2
X_47016_ _47016_/A _52803_/B sky130_fd_sc_hd__buf_2
X_44228_ _44010_/A _44228_/X sky130_fd_sc_hd__buf_2
X_63062_ _60607_/A _63085_/D sky130_fd_sc_hd__buf_2
X_75048_ _75047_/A _75039_/X _75051_/B _75048_/Y sky130_fd_sc_hd__nand3_4
X_79925_ _79924_/B _79924_/C _79926_/A sky130_fd_sc_hd__nand2_4
X_60274_ _60239_/A _60274_/X sky130_fd_sc_hd__buf_2
X_62013_ _58258_/A _63585_/B sky130_fd_sc_hd__buf_2
X_67870_ _87389_/Q _67868_/X _67821_/X _67869_/X _67870_/X sky130_fd_sc_hd__a211o_4
X_44159_ _44151_/X _44153_/X _44157_/Y _44158_/Y _44159_/X sky130_fd_sc_hd__or4_4
X_79856_ _79853_/X _79856_/B _79855_/X _79856_/X sky130_fd_sc_hd__and3_4
X_66821_ _66818_/X _66820_/X _66726_/X _66821_/X sky130_fd_sc_hd__a21o_4
X_78807_ _78807_/A _82834_/Q _78807_/Y sky130_fd_sc_hd__nand2_4
X_48967_ _48967_/A _49009_/B _48967_/Y sky130_fd_sc_hd__nor2_4
X_79787_ _79786_/X _79793_/A sky130_fd_sc_hd__inv_2
X_76999_ _76999_/A _62254_/C _76999_/X sky130_fd_sc_hd__xor2_4
X_69540_ _69505_/X _69340_/X _69538_/Y _69539_/Y _69540_/X sky130_fd_sc_hd__a211o_4
X_47918_ _47918_/A _48790_/A sky130_fd_sc_hd__buf_2
X_66752_ _66728_/A _66752_/B _66752_/X sky130_fd_sc_hd__and2_4
X_78738_ _78770_/A _78737_/Y _78739_/A sky130_fd_sc_hd__and2_4
X_63964_ _64378_/B _64179_/B _64081_/C _60889_/X _63964_/Y sky130_fd_sc_hd__nand4_4
X_48898_ _48898_/A _48901_/A sky130_fd_sc_hd__buf_2
X_65703_ _65685_/X _86191_/Q _65701_/X _65702_/X _65703_/X sky130_fd_sc_hd__a211o_4
X_62915_ _60257_/X _61609_/X _62679_/X _60281_/A _84890_/Q _62916_/A
+ sky130_fd_sc_hd__a32o_4
X_69471_ _69467_/X _69470_/X _69346_/X _69471_/X sky130_fd_sc_hd__a21o_4
X_47849_ _82368_/Q _46579_/X _47849_/X sky130_fd_sc_hd__or2_4
X_78669_ _78667_/X _78669_/B _78669_/X sky130_fd_sc_hd__and2_4
X_66683_ _66683_/A _66683_/B _66683_/X sky130_fd_sc_hd__and2_4
X_63895_ _63831_/A _59392_/A _63862_/C _63895_/X sky130_fd_sc_hd__and3_4
X_80700_ _81084_/CLK _80732_/Q _80700_/Q sky130_fd_sc_hd__dfxtp_4
X_68422_ _69877_/A _88369_/Q _68422_/X sky130_fd_sc_hd__and2_4
X_65634_ _65634_/A _65397_/B _65634_/C _65634_/Y sky130_fd_sc_hd__nor3_4
X_50860_ _50845_/A _54071_/B _50860_/Y sky130_fd_sc_hd__nand2_4
X_62846_ _61522_/X _62834_/B _62801_/X _62889_/D _62846_/Y sky130_fd_sc_hd__nand4_4
X_81680_ _81680_/CLK _80078_/X _81680_/Q sky130_fd_sc_hd__dfxtp_4
X_49519_ _86372_/Q _49496_/X _49518_/Y _49519_/Y sky130_fd_sc_hd__o21ai_4
X_80631_ _80633_/C _80632_/B sky130_fd_sc_hd__inv_2
X_68353_ _69182_/A _68353_/X sky130_fd_sc_hd__buf_2
X_65565_ _65362_/X _85592_/Q _65363_/X _65564_/X _65565_/X sky130_fd_sc_hd__a211o_4
X_50791_ _86132_/Q _50775_/X _50790_/Y _50791_/Y sky130_fd_sc_hd__o21ai_4
X_62777_ _62731_/A _63127_/A _62744_/X _62789_/D _62777_/X sky130_fd_sc_hd__and4_4
X_67304_ _80899_/D _67211_/X _67303_/X _84075_/D sky130_fd_sc_hd__a21bo_4
X_52530_ _52518_/A _46500_/Y _52530_/Y sky130_fd_sc_hd__nand2_4
X_64516_ _58978_/Y _64249_/A _64515_/Y _64516_/Y sky130_fd_sc_hd__o21ai_4
X_83350_ _83480_/CLK _83350_/D _83350_/Q sky130_fd_sc_hd__dfxtp_4
X_61728_ _61728_/A _61728_/X sky130_fd_sc_hd__buf_2
X_80562_ _80554_/Y _80562_/B _80562_/Y sky130_fd_sc_hd__nand2_4
X_68284_ _67754_/X _67757_/X _68283_/X _68284_/Y sky130_fd_sc_hd__a21oi_4
X_65496_ _65399_/X _65494_/Y _65495_/Y _65496_/Y sky130_fd_sc_hd__o21ai_4
XPHY_109 sky130_fd_sc_hd__decap_3
X_82301_ _82301_/CLK _77194_/B _82301_/Q sky130_fd_sc_hd__dfxtp_4
X_67235_ _84078_/Q _67211_/X _67234_/X _67235_/X sky130_fd_sc_hd__a21bo_4
X_52461_ _85817_/Q _52438_/X _52460_/Y _52461_/Y sky130_fd_sc_hd__o21ai_4
X_64447_ _64494_/A _63238_/B _64207_/A _64447_/X sky130_fd_sc_hd__and3_4
X_83281_ _86303_/CLK _72127_/Y _83281_/Q sky130_fd_sc_hd__dfxtp_4
X_61659_ _61413_/A _61690_/A sky130_fd_sc_hd__buf_2
X_80493_ _80487_/Y _80492_/Y _80493_/X sky130_fd_sc_hd__xor2_4
X_54200_ _54196_/Y _54197_/X _54199_/X _54200_/Y sky130_fd_sc_hd__a21oi_4
X_85020_ _85050_/CLK _85020_/D _85020_/Q sky130_fd_sc_hd__dfxtp_4
X_51412_ _51409_/Y _51229_/X _51411_/X _86015_/D sky130_fd_sc_hd__a21oi_4
X_82232_ _81928_/CLK _82264_/Q _77549_/A sky130_fd_sc_hd__dfxtp_4
X_55180_ _55171_/X _83748_/Q _55178_/X _55181_/B sky130_fd_sc_hd__nand3_4
X_67166_ _66898_/X _67166_/X sky130_fd_sc_hd__buf_2
X_52392_ _52388_/Y _52390_/X _52391_/X _52392_/Y sky130_fd_sc_hd__a21oi_4
X_64378_ _64377_/X _64378_/B _64333_/X _64378_/X sky130_fd_sc_hd__and3_4
X_54131_ _85498_/Q _54113_/X _54130_/Y _54131_/Y sky130_fd_sc_hd__o21ai_4
X_66117_ _65595_/X _66117_/X sky130_fd_sc_hd__buf_2
X_51343_ _52524_/A _51266_/B _51352_/C _51343_/X sky130_fd_sc_hd__and3_4
X_63329_ _79183_/B _79184_/A sky130_fd_sc_hd__inv_2
X_82163_ _84161_/CLK _80481_/B _82163_/Q sky130_fd_sc_hd__dfxtp_4
X_67097_ _67023_/A _86784_/Q _67097_/X sky130_fd_sc_hd__and2_4
X_81114_ _81082_/CLK _79813_/X _75637_/A sky130_fd_sc_hd__dfxtp_4
X_54062_ _54059_/Y _54060_/X _54061_/Y _54062_/Y sky130_fd_sc_hd__a21boi_4
X_66048_ _66164_/A _65888_/B _66048_/C _66048_/Y sky130_fd_sc_hd__nor3_4
X_51274_ _51278_/A _46339_/A _51274_/X sky130_fd_sc_hd__and2_4
X_86971_ _87473_/CLK _44757_/X _86971_/Q sky130_fd_sc_hd__dfxtp_4
X_82094_ _82139_/CLK _82094_/D _82094_/Q sky130_fd_sc_hd__dfxtp_4
X_53013_ _85713_/Q _53010_/X _53012_/Y _53013_/Y sky130_fd_sc_hd__o21ai_4
X_50225_ _86240_/Q _50220_/X _50224_/Y _50225_/Y sky130_fd_sc_hd__o21ai_4
X_85922_ _85444_/CLK _51920_/Y _85922_/Q sky130_fd_sc_hd__dfxtp_4
X_81045_ _81117_/CLK _75357_/Y _81045_/Q sky130_fd_sc_hd__dfxtp_4
X_58870_ _58856_/Y _58857_/X _58863_/X _58869_/X _84794_/D sky130_fd_sc_hd__a22oi_4
X_57821_ _86651_/Q _57833_/B _57821_/Y sky130_fd_sc_hd__nor2_4
X_69807_ _44148_/A _69897_/A sky130_fd_sc_hd__buf_2
X_50156_ _52365_/A _51256_/B _50147_/C _50156_/X sky130_fd_sc_hd__and3_4
X_85853_ _83623_/CLK _85853_/D _64719_/B sky130_fd_sc_hd__dfxtp_4
X_67999_ _87959_/Q _67950_/X _67997_/X _67998_/X _67999_/X sky130_fd_sc_hd__a211o_4
X_84804_ _86713_/CLK _84804_/D _84804_/Q sky130_fd_sc_hd__dfxtp_4
X_57752_ _84950_/Q _57691_/X _57746_/X _57751_/X _84950_/D sky130_fd_sc_hd__a2bb2oi_4
X_69738_ _73108_/A _68467_/X _69371_/X _69737_/Y _69738_/X sky130_fd_sc_hd__a211o_4
X_54964_ _54964_/A _54955_/B _54255_/C _47540_/A _54964_/X sky130_fd_sc_hd__and4_4
X_50087_ _50085_/Y _50068_/X _50086_/X _86267_/D sky130_fd_sc_hd__a21oi_4
X_85784_ _82769_/CLK _85784_/D _85784_/Q sky130_fd_sc_hd__dfxtp_4
X_82996_ _85013_/CLK _74654_/X _45604_/A sky130_fd_sc_hd__dfxtp_4
X_56703_ _44253_/X _56703_/X sky130_fd_sc_hd__buf_2
X_87523_ _88034_/CLK _87523_/D _87523_/Q sky130_fd_sc_hd__dfxtp_4
X_53915_ _53902_/A _50183_/B _53915_/Y sky130_fd_sc_hd__nand2_4
X_84735_ _83402_/CLK _84735_/D _59430_/A sky130_fd_sc_hd__dfxtp_4
X_81947_ _82009_/CLK _78042_/Y _77609_/A sky130_fd_sc_hd__dfxtp_4
X_57683_ _84954_/Q _57683_/X sky130_fd_sc_hd__buf_2
X_69669_ _69238_/X _69241_/X _69575_/X _69669_/Y sky130_fd_sc_hd__a21oi_4
X_54895_ _85358_/Q _54892_/X _54894_/Y _54895_/Y sky130_fd_sc_hd__o21ai_4
X_71700_ _71338_/A _71685_/X _70476_/X _71700_/Y sky130_fd_sc_hd__nand3_4
X_59422_ _59417_/X _83482_/Q _59421_/Y _84738_/D sky130_fd_sc_hd__o21a_4
X_56634_ _56633_/X _56634_/X sky130_fd_sc_hd__buf_2
X_41860_ _40548_/X _48226_/A _88116_/Q _40599_/A _88116_/D sky130_fd_sc_hd__a2bb2o_4
X_87454_ _87708_/CLK _43374_/X _87454_/Q sky130_fd_sc_hd__dfxtp_4
X_53846_ _53846_/A _53846_/X sky130_fd_sc_hd__buf_2
X_72680_ _70221_/C _72672_/X _72679_/Y _72680_/X sky130_fd_sc_hd__a21bo_4
X_84666_ _84503_/CLK _84666_/D _80091_/A sky130_fd_sc_hd__dfxtp_4
X_81878_ _81883_/CLK _78069_/X _81846_/D sky130_fd_sc_hd__dfxtp_4
X_86405_ _83783_/CLK _86405_/D _65343_/B sky130_fd_sc_hd__dfxtp_4
X_40811_ _40810_/X _40793_/X _88330_/Q _40794_/X _40811_/X sky130_fd_sc_hd__a2bb2o_4
X_59353_ _84749_/Q _59339_/X _59343_/X _59352_/X _84749_/D sky130_fd_sc_hd__a2bb2oi_4
X_71631_ _71641_/A _71637_/C sky130_fd_sc_hd__buf_2
X_83617_ _85562_/CLK _71074_/Y _48962_/A sky130_fd_sc_hd__dfxtp_4
X_56565_ _56561_/X _56798_/B _56931_/A _56565_/Y sky130_fd_sc_hd__nand3_4
X_80829_ _81065_/CLK _83973_/Q _75669_/B sky130_fd_sc_hd__dfxtp_4
X_87385_ _87189_/CLK _43509_/X _87385_/Q sky130_fd_sc_hd__dfxtp_4
X_41791_ _41790_/X _41791_/X sky130_fd_sc_hd__buf_2
X_53777_ _85570_/Q _53722_/X _53776_/Y _53777_/Y sky130_fd_sc_hd__o21ai_4
X_84597_ _84333_/CLK _60575_/X _79137_/A sky130_fd_sc_hd__dfxtp_4
X_50989_ _50973_/X _50985_/B _50985_/C _52681_/D _50989_/X sky130_fd_sc_hd__and4_4
X_58304_ _64546_/C _63703_/B sky130_fd_sc_hd__buf_2
X_43530_ _43529_/Y _87374_/D sky130_fd_sc_hd__inv_2
X_55516_ _44112_/X _55516_/X sky130_fd_sc_hd__buf_2
X_86336_ _86655_/CLK _86336_/D _57721_/B sky130_fd_sc_hd__dfxtp_4
X_74350_ _83088_/Q _74340_/X _74349_/Y _74350_/X sky130_fd_sc_hd__a21bo_4
X_40742_ _40698_/X _82853_/Q _40741_/X _40742_/X sky130_fd_sc_hd__o21a_4
X_52728_ _52619_/A _52728_/X sky130_fd_sc_hd__buf_2
X_59284_ _59273_/X _85642_/Q _59196_/X _59284_/X sky130_fd_sc_hd__o21a_4
X_71562_ _71557_/X _83456_/Q _71561_/Y _83456_/D sky130_fd_sc_hd__a21o_4
X_83548_ _85354_/CLK _83548_/D _47725_/A sky130_fd_sc_hd__dfxtp_4
X_56496_ _56448_/X _56507_/B sky130_fd_sc_hd__buf_2
X_73301_ _73297_/X _73300_/X _73200_/X _73301_/X sky130_fd_sc_hd__a21o_4
XPHY_610 sky130_fd_sc_hd__decap_3
X_70513_ _71054_/A _70945_/B sky130_fd_sc_hd__buf_2
X_58235_ _46179_/X _58232_/X _58234_/Y _58235_/X sky130_fd_sc_hd__o21a_4
X_43461_ _43461_/A _87411_/D sky130_fd_sc_hd__inv_2
X_55447_ _55201_/Y _55299_/Y _55446_/X _55447_/Y sky130_fd_sc_hd__o21ai_4
X_74281_ _74279_/X _74268_/X _74281_/C _74281_/Y sky130_fd_sc_hd__nand3_4
X_86267_ _83305_/CLK _86267_/D _86267_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_621 sky130_fd_sc_hd__decap_3
X_52659_ _85778_/Q _52656_/X _52658_/Y _52659_/Y sky130_fd_sc_hd__o21ai_4
X_40673_ _40672_/Y _40673_/X sky130_fd_sc_hd__buf_2
X_71493_ _71487_/X _83480_/Q _71492_/X _83480_/D sky130_fd_sc_hd__a21o_4
X_83479_ _83415_/CLK _83479_/D _83479_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_632 sky130_fd_sc_hd__decap_3
XPHY_643 sky130_fd_sc_hd__decap_3
X_45200_ _44972_/X _45200_/X sky130_fd_sc_hd__buf_2
X_76020_ _81711_/D _76021_/B _76020_/Y sky130_fd_sc_hd__nor2_4
X_88006_ _88006_/CLK _88006_/D _88006_/Q sky130_fd_sc_hd__dfxtp_4
X_42412_ _42401_/X _42410_/X _40459_/X _87876_/Q _42411_/X _42412_/Y
+ sky130_fd_sc_hd__o32ai_4
XPHY_654 sky130_fd_sc_hd__decap_3
X_73232_ _87053_/Q _73129_/X _73231_/X _73232_/Y sky130_fd_sc_hd__o21ai_4
X_85218_ _85250_/CLK _85218_/D _55736_/B sky130_fd_sc_hd__dfxtp_4
X_70444_ _70426_/A _71650_/A sky130_fd_sc_hd__buf_2
X_46180_ _46120_/B _72527_/A _46179_/X _46112_/A _46111_/X _46180_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_58166_ _58166_/A _63069_/A sky130_fd_sc_hd__inv_2
XPHY_665 sky130_fd_sc_hd__decap_3
X_43392_ _41447_/X _43386_/X _87445_/Q _43388_/X _87445_/D sky130_fd_sc_hd__a2bb2o_4
X_55378_ _55322_/X _55324_/X _55378_/X sky130_fd_sc_hd__and2_4
X_86198_ _86196_/CLK _50452_/Y _86198_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_676 sky130_fd_sc_hd__decap_3
XPHY_687 sky130_fd_sc_hd__decap_3
XPHY_698 sky130_fd_sc_hd__decap_3
X_45131_ _45197_/A _45131_/X sky130_fd_sc_hd__buf_2
X_57117_ _56626_/X _57105_/Y _57116_/Y _85079_/D sky130_fd_sc_hd__a21oi_4
X_42343_ _42304_/X _42343_/X sky130_fd_sc_hd__buf_2
X_54329_ _54329_/A _54353_/B sky130_fd_sc_hd__buf_2
X_73163_ _73163_/A _73163_/X sky130_fd_sc_hd__buf_2
X_85149_ _85152_/CLK _56585_/X _55590_/B sky130_fd_sc_hd__dfxtp_4
X_70375_ _70366_/X _70374_/X _70375_/C _70375_/Y sky130_fd_sc_hd__nand3_4
X_58097_ _58097_/A _58136_/B _58097_/Y sky130_fd_sc_hd__nor2_4
X_72114_ _72111_/Y _72059_/X _72113_/X _72114_/Y sky130_fd_sc_hd__a21oi_4
X_45062_ _85207_/Q _45027_/X _45061_/X _45062_/Y sky130_fd_sc_hd__o21ai_4
X_57048_ _56551_/X _57049_/A sky130_fd_sc_hd__buf_2
X_42274_ _41511_/X _42271_/X _87945_/Q _42272_/X _42274_/X sky130_fd_sc_hd__a2bb2o_4
X_73094_ _72959_/X _85589_/Q _73092_/X _73093_/X _73094_/X sky130_fd_sc_hd__a211o_4
X_77971_ _81948_/D _77964_/A _77971_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_440_0_CLK clkbuf_9_220_0_CLK/X _84210_/CLK sky130_fd_sc_hd__clkbuf_1
X_44013_ _64806_/A _64629_/A sky130_fd_sc_hd__buf_2
X_79710_ _79699_/X _79710_/B _79710_/Y sky130_fd_sc_hd__nand2_4
X_41225_ _41224_/X _41225_/X sky130_fd_sc_hd__buf_2
X_72045_ _72041_/Y _71978_/X _72044_/X _72045_/Y sky130_fd_sc_hd__a21oi_4
X_76922_ _76914_/A _76914_/B _76921_/Y _76922_/Y sky130_fd_sc_hd__o21ai_4
X_49870_ _49924_/A _49870_/X sky130_fd_sc_hd__buf_2
X_48821_ _86476_/Q _48809_/X _48820_/Y _48821_/Y sky130_fd_sc_hd__o21ai_4
X_79641_ _79630_/X _79627_/Y _79642_/D sky130_fd_sc_hd__nand2_4
X_41156_ _41061_/X _81721_/Q _41155_/X _41157_/A sky130_fd_sc_hd__o21ai_4
X_76853_ _76837_/B _76850_/X _76852_/Y _76854_/B sky130_fd_sc_hd__a21oi_4
X_58999_ _58961_/X _85665_/Q _58900_/X _58999_/X sky130_fd_sc_hd__o21a_4
X_75804_ _75803_/C _75787_/A _75786_/X _75804_/Y sky130_fd_sc_hd__nand3_4
X_48752_ _48752_/A _48766_/B _48761_/C _48752_/X sky130_fd_sc_hd__and3_4
X_79572_ _65348_/C _83253_/Q _79572_/Y sky130_fd_sc_hd__nand2_4
X_45964_ _45964_/A _45964_/X sky130_fd_sc_hd__buf_2
X_41087_ _41086_/X _41087_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_455_0_CLK clkbuf_9_227_0_CLK/X _85692_/CLK sky130_fd_sc_hd__clkbuf_1
X_76784_ _81489_/Q _76784_/Y sky130_fd_sc_hd__inv_2
X_73996_ _72744_/X _85615_/Q _72857_/X _73995_/X _73996_/X sky130_fd_sc_hd__a211o_4
X_47703_ _47697_/Y _47698_/X _47702_/X _86607_/D sky130_fd_sc_hd__a21oi_4
X_78523_ _78524_/A _82673_/D _78526_/B sky130_fd_sc_hd__nor2_4
X_44915_ _56379_/C _44880_/X _44914_/X _44915_/Y sky130_fd_sc_hd__o21ai_4
X_75735_ _75735_/A _75735_/Y sky130_fd_sc_hd__inv_2
X_48683_ _48683_/A _48684_/B sky130_fd_sc_hd__buf_2
X_60961_ _59875_/A _60961_/X sky130_fd_sc_hd__buf_2
X_72947_ _72947_/A _72924_/B _72947_/Y sky130_fd_sc_hd__nor2_4
X_45895_ _45894_/X _86847_/D sky130_fd_sc_hd__inv_2
X_62700_ _62658_/A _84717_/Q _62676_/C _62657_/X _62700_/X sky130_fd_sc_hd__and4_4
X_47634_ _86614_/Q _47619_/X _47633_/Y _47634_/Y sky130_fd_sc_hd__o21ai_4
X_78454_ _82508_/Q _82764_/D _78454_/X sky130_fd_sc_hd__xor2_4
X_44846_ _44846_/A _86923_/D sky130_fd_sc_hd__inv_2
X_63680_ _63670_/A _63670_/B _80323_/B _63680_/Y sky130_fd_sc_hd__nor3_4
X_75666_ _75666_/A _75680_/A _75667_/B sky130_fd_sc_hd__xor2_4
X_60892_ _61293_/A _60861_/X _60844_/X _60857_/D _60892_/Y sky130_fd_sc_hd__a22oi_4
X_72878_ _72872_/X _72875_/X _72877_/X _72883_/A sky130_fd_sc_hd__a21o_4
X_77405_ _77406_/A _82094_/D _77405_/Y sky130_fd_sc_hd__nor2_4
X_62631_ _61695_/A _62631_/B _62631_/C _62631_/D _62634_/B sky130_fd_sc_hd__nand4_4
X_74617_ _74605_/X _74613_/X _56152_/Y _74614_/X _74617_/X sky130_fd_sc_hd__a211o_4
X_47565_ _47565_/A _47595_/C sky130_fd_sc_hd__buf_2
X_71829_ _71068_/B _71829_/X sky130_fd_sc_hd__buf_2
X_78385_ _78385_/A _82664_/D _78385_/Y sky130_fd_sc_hd__nand2_4
X_44777_ _41360_/Y _44774_/X _86961_/Q _44775_/X _44777_/X sky130_fd_sc_hd__a2bb2o_4
X_75597_ _80996_/Q _75597_/B _75597_/X sky130_fd_sc_hd__xor2_4
X_41989_ _41982_/X _41975_/X _40781_/X _41988_/Y _41984_/X _88080_/D
+ sky130_fd_sc_hd__o32ai_4
X_49304_ _51330_/A _49283_/B _49234_/X _49304_/X sky130_fd_sc_hd__and3_4
X_46516_ _51356_/B _49322_/B sky130_fd_sc_hd__buf_2
X_65350_ _64666_/A _65350_/X sky130_fd_sc_hd__buf_2
X_77336_ _77334_/Y _77335_/Y _82185_/D sky130_fd_sc_hd__xnor2_4
X_43728_ _87293_/Q _69862_/B sky130_fd_sc_hd__inv_2
X_62562_ _62556_/X _62558_/X _62561_/Y _58344_/A _62511_/X _62562_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74548_ _56019_/Y _74538_/Y _74547_/Y _74548_/Y sky130_fd_sc_hd__o21ai_4
X_47496_ _47492_/Y _47462_/X _47495_/X _47496_/Y sky130_fd_sc_hd__a21oi_4
X_64301_ _59388_/A _64301_/B _64301_/Y sky130_fd_sc_hd__nor2_4
X_49235_ _50755_/A _49113_/B _49234_/X _49235_/X sky130_fd_sc_hd__and3_4
X_61513_ _61513_/A _61468_/B _61467_/X _61512_/X _61513_/Y sky130_fd_sc_hd__nand4_4
X_46447_ _46505_/A _46447_/B _46447_/Y sky130_fd_sc_hd__nand2_4
X_65281_ _65281_/A _65280_/X _65281_/Y sky130_fd_sc_hd__nand2_4
X_77267_ _77264_/Y _82213_/Q _77265_/Y _77267_/Y sky130_fd_sc_hd__nand3_4
X_43659_ _47834_/A _43659_/X sky130_fd_sc_hd__buf_2
X_74479_ _74477_/Y _74463_/X _74478_/X _74479_/Y sky130_fd_sc_hd__a21oi_4
X_62493_ _62493_/A _62490_/Y _62493_/C _62492_/Y _62493_/Y sky130_fd_sc_hd__nand4_4
X_67020_ _87872_/Q _66994_/X _66926_/X _67019_/X _67020_/X sky130_fd_sc_hd__a211o_4
X_79006_ _78993_/A _79000_/A _79006_/X sky130_fd_sc_hd__and2_4
X_64232_ _79872_/B _63258_/X _64231_/X _64232_/X sky130_fd_sc_hd__a21o_4
X_76218_ _76215_/Y _76234_/A _76216_/Y _76221_/C sky130_fd_sc_hd__nand3_4
X_49166_ _83597_/Q _49166_/Y sky130_fd_sc_hd__inv_2
X_61444_ _61437_/Y _61439_/Y _61403_/X _61440_/Y _61443_/Y _61444_/X
+ sky130_fd_sc_hd__a41o_4
X_46378_ _46387_/A _50781_/B _46378_/Y sky130_fd_sc_hd__nand2_4
X_77198_ _77198_/A _77198_/B _77199_/B sky130_fd_sc_hd__xor2_4
X_48117_ _66298_/B _48103_/X _48116_/Y _48117_/Y sky130_fd_sc_hd__o21ai_4
X_45329_ _45325_/Y _45328_/Y _45287_/X _45329_/X sky130_fd_sc_hd__a21o_4
X_64163_ _64159_/X _63741_/X _64160_/Y _64161_/Y _64162_/X _64163_/X
+ sky130_fd_sc_hd__a41o_4
X_76149_ _76145_/A _76145_/B _76149_/C _76150_/B sky130_fd_sc_hd__nand3_4
X_49097_ _46495_/B _46348_/A _49097_/Y sky130_fd_sc_hd__nand2_4
X_61375_ _61375_/A _61375_/B _61375_/C _61375_/Y sky130_fd_sc_hd__nand3_4
X_63114_ _63231_/A _63114_/X sky130_fd_sc_hd__buf_2
X_60326_ _79700_/A _60323_/X _60306_/Y _60325_/Y _60326_/X sky130_fd_sc_hd__o22a_4
X_48048_ _48042_/Y _48007_/X _48047_/X _86573_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_408_0_CLK clkbuf_9_204_0_CLK/X _83515_/CLK sky130_fd_sc_hd__clkbuf_1
X_68971_ _87079_/Q _68948_/X _68875_/X _68970_/X _68971_/X sky130_fd_sc_hd__a211o_4
X_64094_ _64090_/Y _64094_/B _64094_/C _64094_/D _64094_/X sky130_fd_sc_hd__and4_4
X_67922_ _67664_/X _67911_/Y _67863_/X _67921_/Y _67922_/X sky130_fd_sc_hd__a211o_4
X_79908_ _60148_/C _79908_/B _79913_/B sky130_fd_sc_hd__nand2_4
X_63045_ _63042_/Y _63044_/X _61194_/X _63045_/Y sky130_fd_sc_hd__a21oi_4
X_60257_ _60199_/X _60179_/Y _60257_/X sky130_fd_sc_hd__and2_4
X_50010_ _50025_/A _49994_/X _50025_/C _53223_/D _50010_/X sky130_fd_sc_hd__and4_4
X_67853_ _67901_/A _87709_/Q _67853_/X sky130_fd_sc_hd__and2_4
X_79839_ _79835_/X _79854_/B _79839_/X sky130_fd_sc_hd__xor2_4
X_60188_ _60204_/A _60189_/A sky130_fd_sc_hd__buf_2
X_49999_ _49995_/A _49994_/X _50005_/C _53211_/D _49999_/X sky130_fd_sc_hd__and4_4
X_66804_ _66800_/X _66803_/X _66706_/X _66804_/Y sky130_fd_sc_hd__a21oi_4
X_82850_ _82563_/CLK _78083_/B _40927_/A sky130_fd_sc_hd__dfxtp_4
X_67784_ _87904_/Q _67713_/X _67761_/X _67783_/X _67784_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_8_82_0_CLK clkbuf_8_83_0_CLK/A clkbuf_8_82_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_64996_ _84219_/Q _64997_/C sky130_fd_sc_hd__inv_2
X_81801_ _81801_/CLK _81609_/Q _81801_/Q sky130_fd_sc_hd__dfxtp_4
X_69523_ _69383_/A _69523_/B _69523_/X sky130_fd_sc_hd__and2_4
X_66735_ _66534_/A _66760_/A sky130_fd_sc_hd__buf_2
X_51961_ _53199_/A _51961_/X sky130_fd_sc_hd__buf_2
X_63947_ _61492_/A _63947_/B _63947_/C _64025_/D _63947_/Y sky130_fd_sc_hd__nand4_4
X_82781_ _82973_/CLK _78725_/X _82781_/Q sky130_fd_sc_hd__dfxtp_4
X_53700_ _85585_/Q _53687_/X _53699_/Y _53700_/Y sky130_fd_sc_hd__o21ai_4
X_84520_ _84520_/CLK _61106_/Y _84520_/Q sky130_fd_sc_hd__dfxtp_4
X_50912_ _50932_/A _46662_/X _50912_/Y sky130_fd_sc_hd__nand2_4
X_81732_ _81169_/CLK _75938_/Y _41440_/A sky130_fd_sc_hd__dfxtp_4
X_69454_ _69454_/A _87260_/Q _69454_/X sky130_fd_sc_hd__and2_4
X_54680_ _54674_/A _54674_/B _54674_/C _47329_/A _54680_/X sky130_fd_sc_hd__and4_4
X_66666_ _87439_/Q _66642_/X _66643_/X _66665_/X _66666_/X sky130_fd_sc_hd__a211o_4
X_51892_ _52626_/A _51893_/C sky130_fd_sc_hd__buf_2
X_63878_ _63831_/A _59388_/A _63862_/C _63878_/X sky130_fd_sc_hd__and3_4
X_68405_ _68405_/A _87250_/Q _68405_/X sky130_fd_sc_hd__and2_4
X_65617_ _64599_/X _83069_/Q _65015_/X _65616_/X _65617_/X sky130_fd_sc_hd__a211o_4
X_53631_ _48388_/A _53658_/B _53620_/C _53631_/X sky130_fd_sc_hd__and3_4
X_84451_ _84454_/CLK _61836_/Y _78074_/B sky130_fd_sc_hd__dfxtp_4
X_50843_ _86122_/Q _50804_/X _50842_/Y _50843_/Y sky130_fd_sc_hd__o21ai_4
X_62829_ _62971_/A _84826_/Q _62819_/C _62782_/X _62829_/X sky130_fd_sc_hd__and4_4
Xclkbuf_8_97_0_CLK clkbuf_8_97_0_CLK/A clkbuf_8_97_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_81663_ _81269_/CLK _81695_/Q _76593_/A sky130_fd_sc_hd__dfxtp_4
X_69385_ _69678_/A _69385_/X sky130_fd_sc_hd__buf_2
X_66597_ _66597_/A _66596_/X _66597_/Y sky130_fd_sc_hd__nand2_4
X_83402_ _83402_/CLK _83402_/D _83402_/Q sky130_fd_sc_hd__dfxtp_4
X_56350_ _56350_/A _56350_/X sky130_fd_sc_hd__buf_2
X_80614_ _80614_/A _80614_/B _80614_/X sky130_fd_sc_hd__xor2_4
X_68336_ _68319_/X _68049_/Y _68326_/X _68335_/Y _68336_/X sky130_fd_sc_hd__a211o_4
X_87170_ _84534_/CLK _44314_/Y _44313_/B sky130_fd_sc_hd__dfxtp_4
X_53562_ _53559_/Y _53537_/X _53561_/X _85613_/D sky130_fd_sc_hd__a21oi_4
X_65548_ _64832_/X _65548_/B _64837_/X _65557_/A sky130_fd_sc_hd__nand3_4
X_84382_ _84520_/CLK _84382_/D _75912_/B sky130_fd_sc_hd__dfxtp_4
X_50774_ _50772_/Y _50768_/X _50773_/Y _86136_/D sky130_fd_sc_hd__a21boi_4
X_81594_ _81433_/CLK _65546_/C _76872_/A sky130_fd_sc_hd__dfxtp_4
X_55301_ _55300_/X _55301_/X sky130_fd_sc_hd__buf_2
X_86121_ _86121_/CLK _50851_/Y _86121_/Q sky130_fd_sc_hd__dfxtp_4
X_52513_ _52487_/X _50816_/B _52513_/Y sky130_fd_sc_hd__nand2_4
X_83333_ _83333_/CLK _83333_/D _83333_/Q sky130_fd_sc_hd__dfxtp_4
X_80545_ _84769_/Q _84161_/Q _80545_/Y sky130_fd_sc_hd__nand2_4
X_56281_ _56281_/A _56280_/Y _56281_/Y sky130_fd_sc_hd__nand2_4
X_68267_ _67388_/X _68447_/A sky130_fd_sc_hd__buf_2
X_53493_ _50270_/A _53474_/B _53492_/X _53493_/X sky130_fd_sc_hd__and3_4
X_65479_ _64682_/X _65647_/B _64685_/X _65479_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_8_20_0_CLK clkbuf_8_21_0_CLK/A clkbuf_8_20_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_58020_ _58020_/A _58020_/X sky130_fd_sc_hd__buf_2
X_55232_ _85028_/Q _55142_/A _80665_/Q _55231_/Y _55232_/X sky130_fd_sc_hd__a211o_4
X_67218_ _67149_/A _67218_/B _67218_/X sky130_fd_sc_hd__and2_4
X_86052_ _86054_/CLK _51221_/Y _86052_/Q sky130_fd_sc_hd__dfxtp_4
X_52444_ _52448_/A _46295_/A _52444_/Y sky130_fd_sc_hd__nand2_4
X_83264_ _81233_/CLK _83264_/D _72323_/A sky130_fd_sc_hd__dfxtp_4
X_80476_ _80476_/A _80476_/B _80489_/B sky130_fd_sc_hd__xnor2_4
X_68198_ _68196_/X _67220_/Y _68189_/X _68197_/Y _68198_/X sky130_fd_sc_hd__a211o_4
X_85003_ _85003_/CLK _57447_/Y _85003_/Q sky130_fd_sc_hd__dfxtp_4
X_82215_ _82084_/CLK _82247_/Q _77312_/A sky130_fd_sc_hd__dfxtp_4
X_55163_ _55296_/B _55162_/Y _55163_/Y sky130_fd_sc_hd__nand2_4
X_67149_ _67149_/A _88123_/Q _67149_/X sky130_fd_sc_hd__and2_4
X_52375_ _85835_/Q _52372_/X _52374_/Y _52375_/Y sky130_fd_sc_hd__o21ai_4
X_83195_ _83191_/CLK _72671_/X _83195_/Q sky130_fd_sc_hd__dfxtp_4
X_54114_ _54194_/A _54134_/A sky130_fd_sc_hd__buf_2
X_51326_ _51306_/X _51326_/B _51326_/X sky130_fd_sc_hd__and2_4
X_70160_ _70348_/A _70160_/X sky130_fd_sc_hd__buf_2
X_82146_ _82145_/CLK _84138_/Q _77728_/A sky130_fd_sc_hd__dfxtp_4
X_55094_ _85319_/Q _55072_/X _55093_/Y _55094_/Y sky130_fd_sc_hd__o21ai_4
X_59971_ _60042_/A _59971_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_35_0_CLK clkbuf_8_35_0_CLK/A clkbuf_9_71_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_54045_ _54037_/A _52526_/B _54045_/Y sky130_fd_sc_hd__nand2_4
X_58922_ _58635_/A _58923_/A sky130_fd_sc_hd__buf_2
X_51257_ _51254_/Y _51237_/X _51256_/X _51257_/Y sky130_fd_sc_hd__a21oi_4
X_70091_ _83852_/Q _70085_/X _70090_/X _70091_/X sky130_fd_sc_hd__a21bo_4
X_86954_ _88164_/CLK _86954_/D _86954_/Q sky130_fd_sc_hd__dfxtp_4
X_82077_ _81160_/CLK _84037_/Q _82077_/Q sky130_fd_sc_hd__dfxtp_4
X_41010_ _40999_/X _41000_/X _41009_/X _88294_/Q _40995_/X _41010_/Y
+ sky130_fd_sc_hd__o32ai_4
X_50208_ _86242_/Q _50185_/X _50207_/Y _50208_/Y sky130_fd_sc_hd__o21ai_4
X_85905_ _86541_/CLK _52018_/Y _66141_/B sky130_fd_sc_hd__dfxtp_4
X_81028_ _81933_/CLK _75107_/Y _81028_/Q sky130_fd_sc_hd__dfxtp_4
X_58853_ _58853_/A _59090_/B _58853_/Y sky130_fd_sc_hd__nor2_4
X_51188_ _51186_/Y _51175_/X _51187_/X _86058_/D sky130_fd_sc_hd__a21oi_4
X_86885_ _86873_/CLK _45310_/Y _45308_/A sky130_fd_sc_hd__dfxtp_4
X_57804_ _57804_/A _58697_/A sky130_fd_sc_hd__buf_2
X_50139_ _50153_/A _50649_/B _50139_/Y sky130_fd_sc_hd__nand2_4
X_85836_ _85837_/CLK _52371_/Y _65155_/B sky130_fd_sc_hd__dfxtp_4
X_73850_ _73355_/A _73850_/X sky130_fd_sc_hd__buf_2
X_58784_ _58784_/A _58785_/A sky130_fd_sc_hd__buf_2
X_55996_ _55995_/X _55863_/X _56073_/A _74317_/C _55996_/X sky130_fd_sc_hd__and4_4
X_72801_ _43117_/Y _72731_/X _72799_/X _72800_/Y _72801_/X sky130_fd_sc_hd__a211o_4
X_57735_ _46213_/X _57731_/Y _57734_/Y _57700_/X _57703_/X _57735_/X
+ sky130_fd_sc_hd__o32a_4
X_42961_ _40400_/X _42950_/X _87629_/Q _42951_/X _42961_/X sky130_fd_sc_hd__a2bb2o_4
X_54947_ _54945_/Y _54936_/X _54946_/X _85348_/D sky130_fd_sc_hd__a21oi_4
X_73781_ _73731_/X _86232_/Q _73683_/X _73780_/X _73781_/X sky130_fd_sc_hd__a211o_4
X_85767_ _85767_/CLK _52721_/Y _85767_/Q sky130_fd_sc_hd__dfxtp_4
X_70993_ _51324_/B _70983_/X _70992_/Y _83639_/D sky130_fd_sc_hd__o21ai_4
X_82979_ _82979_/CLK _74704_/Y _45861_/A sky130_fd_sc_hd__dfxtp_4
X_44700_ _44700_/A _44700_/Y sky130_fd_sc_hd__inv_2
X_75520_ _75516_/Y _75519_/C _75519_/A _75520_/Y sky130_fd_sc_hd__o21ai_4
X_87506_ _87766_/CLK _87506_/D _87506_/Q sky130_fd_sc_hd__dfxtp_4
X_41912_ _41912_/A _41912_/X sky130_fd_sc_hd__buf_2
X_72732_ _87315_/Q _72732_/B _72732_/Y sky130_fd_sc_hd__nor2_4
X_84718_ _84727_/CLK _59491_/Y _64248_/C sky130_fd_sc_hd__dfxtp_4
X_45680_ _85135_/Q _45556_/X _45651_/X _45680_/X sky130_fd_sc_hd__o21a_4
X_57666_ _57664_/X _57666_/B _57666_/Y sky130_fd_sc_hd__nor2_4
X_42892_ _41643_/X _42886_/X _67378_/B _42887_/X _87665_/D sky130_fd_sc_hd__a2bb2o_4
X_54878_ _54883_/A _54883_/B _54883_/C _53185_/D _54878_/X sky130_fd_sc_hd__and4_4
X_85698_ _85697_/CLK _85698_/D _85698_/Q sky130_fd_sc_hd__dfxtp_4
X_59405_ _84741_/Q _63150_/A sky130_fd_sc_hd__inv_2
X_44631_ _44631_/A _44631_/Y sky130_fd_sc_hd__inv_2
X_56617_ _56617_/A _72656_/C sky130_fd_sc_hd__buf_2
X_87437_ _87126_/CLK _43406_/Y _87437_/Q sky130_fd_sc_hd__dfxtp_4
X_75451_ _75466_/A _75450_/Y _75451_/Y sky130_fd_sc_hd__xnor2_4
X_41843_ _41843_/A _41843_/Y sky130_fd_sc_hd__inv_2
X_53829_ _53773_/A _53829_/X sky130_fd_sc_hd__buf_2
X_72663_ _83199_/Q _72658_/X _72662_/Y _83199_/D sky130_fd_sc_hd__a21bo_4
X_84649_ _84649_/CLK _84649_/D _60214_/C sky130_fd_sc_hd__dfxtp_4
X_57597_ _57597_/A _48297_/X _57597_/Y sky130_fd_sc_hd__nand2_4
X_74402_ _74399_/Y _74370_/X _74401_/X _74402_/Y sky130_fd_sc_hd__a21oi_4
X_47350_ _47346_/Y _47317_/X _47349_/X _86644_/D sky130_fd_sc_hd__a21oi_4
X_59336_ _59286_/X _86054_/Q _59335_/X _59336_/Y sky130_fd_sc_hd__o21ai_4
X_71614_ _71859_/A _70573_/B _71614_/C _71606_/X _71614_/Y sky130_fd_sc_hd__nor4_4
X_78170_ _78161_/A _82862_/D _78170_/Y sky130_fd_sc_hd__nand2_4
X_44562_ _44562_/A _44562_/Y sky130_fd_sc_hd__inv_2
X_56548_ _56547_/X _56548_/X sky130_fd_sc_hd__buf_2
X_75382_ _75382_/A _75383_/C sky130_fd_sc_hd__inv_2
X_87368_ _87373_/CLK _87368_/D _87368_/Q sky130_fd_sc_hd__dfxtp_4
X_41774_ _41753_/X _41754_/X _41773_/X _67992_/B _41736_/X _41775_/A
+ sky130_fd_sc_hd__o32ai_4
X_72594_ _72593_/X _72594_/Y sky130_fd_sc_hd__inv_2
X_46301_ _40365_/X _46301_/X sky130_fd_sc_hd__buf_2
X_77121_ _77126_/A _77111_/X _77120_/Y _77121_/Y sky130_fd_sc_hd__a21boi_4
X_43513_ _43513_/A _43513_/X sky130_fd_sc_hd__buf_2
X_74333_ _70318_/A _74327_/X _74332_/Y _74333_/X sky130_fd_sc_hd__a21bo_4
X_86319_ _86640_/CLK _49812_/Y _57971_/B sky130_fd_sc_hd__dfxtp_4
X_40725_ _40687_/X _40688_/X _40724_/X _88347_/Q _40683_/X _40726_/A
+ sky130_fd_sc_hd__o32ai_4
X_47281_ _47140_/A _47321_/C sky130_fd_sc_hd__buf_2
X_71545_ _71531_/X _83462_/Q _71544_/Y _83462_/D sky130_fd_sc_hd__a21o_4
X_59267_ _84756_/Q _59129_/X _59259_/X _59266_/X _84756_/D sky130_fd_sc_hd__a2bb2oi_4
X_44493_ _41230_/A _44474_/X _87081_/Q _44475_/X _87081_/D sky130_fd_sc_hd__a2bb2o_4
X_56479_ _56474_/X _56472_/B _85180_/Q _56479_/Y sky130_fd_sc_hd__nand3_4
X_87299_ _87553_/CLK _43712_/Y _87299_/Q sky130_fd_sc_hd__dfxtp_4
X_49020_ _49018_/X _48508_/A _49019_/Y _49021_/A sky130_fd_sc_hd__a21o_4
X_46232_ _46174_/X _46175_/Y _46158_/B _46232_/Y sky130_fd_sc_hd__o21ai_4
XPHY_440 sky130_fd_sc_hd__decap_3
X_58218_ _58171_/X _83401_/Q _58217_/Y _84905_/D sky130_fd_sc_hd__o21a_4
X_77052_ _77026_/Y _77051_/X _77052_/Y sky130_fd_sc_hd__nand2_4
X_43444_ _43443_/Y _43444_/Y sky130_fd_sc_hd__inv_2
X_74264_ _88084_/Q _73599_/B _74264_/Y sky130_fd_sc_hd__nor2_4
XPHY_451 sky130_fd_sc_hd__decap_3
X_40656_ _40656_/A _40656_/X sky130_fd_sc_hd__buf_2
X_59198_ _59121_/X _85425_/Q _59197_/X _59198_/Y sky130_fd_sc_hd__o21ai_4
X_71476_ _71827_/A _71479_/B _70782_/A _71476_/D _71476_/X sky130_fd_sc_hd__and4_4
XPHY_462 sky130_fd_sc_hd__decap_3
XPHY_473 sky130_fd_sc_hd__decap_3
X_76003_ _81517_/Q _81741_/D _76003_/X sky130_fd_sc_hd__xor2_4
X_73215_ _73239_/A _86512_/Q _73215_/X sky130_fd_sc_hd__and2_4
XPHY_484 sky130_fd_sc_hd__decap_3
X_70427_ _70984_/A _70940_/B sky130_fd_sc_hd__buf_2
X_46163_ _46162_/X _46166_/A sky130_fd_sc_hd__buf_2
X_58149_ _58149_/A _63022_/A sky130_fd_sc_hd__inv_2
XPHY_495 sky130_fd_sc_hd__decap_3
X_43375_ _43305_/A _43375_/X sky130_fd_sc_hd__buf_2
X_74195_ _74106_/X _85606_/Q _74107_/X _74194_/X _74195_/X sky130_fd_sc_hd__a211o_4
X_40587_ _40736_/A _40588_/B sky130_fd_sc_hd__buf_2
X_45114_ _85267_/Q _45073_/X _45113_/X _45114_/Y sky130_fd_sc_hd__o21ai_4
X_42326_ _42304_/X _42326_/X sky130_fd_sc_hd__buf_2
X_61160_ _61271_/A _61230_/C _61097_/X _64456_/C _60620_/Y _61160_/Y
+ sky130_fd_sc_hd__a41oi_4
X_73146_ _74139_/A _73339_/A sky130_fd_sc_hd__buf_2
X_46094_ _46094_/A _46094_/X sky130_fd_sc_hd__buf_2
X_70358_ HASH_ADDR[0] _70358_/X sky130_fd_sc_hd__buf_2
X_60111_ _65464_/A _60111_/X sky130_fd_sc_hd__buf_2
X_49922_ _49928_/A _53135_/B _49922_/Y sky130_fd_sc_hd__nand2_4
X_45045_ _55915_/B _45044_/X _45004_/X _45045_/X sky130_fd_sc_hd__o21a_4
X_42257_ _41461_/X _42248_/X _87955_/Q _42249_/X _87955_/D sky130_fd_sc_hd__a2bb2o_4
X_61091_ _61091_/A _61091_/Y sky130_fd_sc_hd__inv_2
X_73077_ _83166_/Q _72943_/X _73076_/Y _73077_/X sky130_fd_sc_hd__a21o_4
X_77954_ _77954_/A _77954_/B _77957_/A sky130_fd_sc_hd__xor2_4
X_70289_ _70238_/A _70289_/X sky130_fd_sc_hd__buf_2
X_41208_ _41136_/X _40689_/A _41207_/X _41209_/A sky130_fd_sc_hd__o21a_4
X_60042_ _60042_/A _60599_/A _60403_/C _60042_/D _60059_/A sky130_fd_sc_hd__and4_4
X_72028_ _83299_/Q _72016_/X _72027_/Y _72028_/Y sky130_fd_sc_hd__o21ai_4
X_76905_ _76905_/A _76904_/Y _76905_/Y sky130_fd_sc_hd__nand2_4
X_49853_ _49825_/A _49853_/X sky130_fd_sc_hd__buf_2
X_42188_ _42173_/X _42169_/X _41277_/X _87989_/Q _42170_/X _42189_/A
+ sky130_fd_sc_hd__o32ai_4
X_77885_ _77885_/A _77872_/Y _77885_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_394_0_CLK clkbuf_9_197_0_CLK/X _84469_/CLK sky130_fd_sc_hd__clkbuf_1
X_48804_ _86479_/Q _48781_/X _48803_/Y _48804_/Y sky130_fd_sc_hd__o21ai_4
X_79624_ _79624_/A _79624_/B _79624_/X sky130_fd_sc_hd__xor2_4
X_41139_ _41138_/X _41139_/X sky130_fd_sc_hd__buf_2
X_64850_ _64850_/A _64851_/A sky130_fd_sc_hd__buf_2
X_76836_ _76831_/Y _76818_/B _76835_/Y _76837_/B sky130_fd_sc_hd__o21ai_4
X_49784_ _49782_/Y _49759_/X _49783_/X _49784_/Y sky130_fd_sc_hd__a21oi_4
X_46996_ _59094_/A _46955_/X _46995_/Y _46996_/Y sky130_fd_sc_hd__o21ai_4
X_63801_ _63799_/X _63744_/X _63800_/Y _63801_/Y sky130_fd_sc_hd__a21oi_4
X_48735_ _48801_/A _48407_/A _48735_/X sky130_fd_sc_hd__and2_4
X_79555_ _79555_/A _79555_/B _79555_/C _79558_/A sky130_fd_sc_hd__nand3_4
X_45947_ _66517_/B _45947_/B _45947_/Y sky130_fd_sc_hd__nand2_4
X_64781_ _64678_/X _85531_/Q _64679_/X _64780_/X _64781_/X sky130_fd_sc_hd__a211o_4
X_76767_ _76765_/Y _76766_/Y _76770_/A sky130_fd_sc_hd__xor2_4
X_73979_ _48014_/Y _73979_/B _73979_/X sky130_fd_sc_hd__xor2_4
X_61993_ _63573_/A _59841_/X _61542_/A _61981_/X _61993_/X sky130_fd_sc_hd__a2bb2o_4
X_66520_ _79165_/B _64532_/X _66519_/X _84107_/D sky130_fd_sc_hd__o21ai_4
X_78506_ _78505_/B _78505_/C _78501_/Y _78510_/C sky130_fd_sc_hd__o21ai_4
X_75718_ _75707_/Y _80785_/D sky130_fd_sc_hd__inv_2
X_63732_ _63721_/Y _63726_/Y _63730_/Y _63731_/Y _63732_/X sky130_fd_sc_hd__and4_4
X_48666_ _48666_/A _48667_/A sky130_fd_sc_hd__buf_2
X_60944_ _64172_/D _60870_/X _63781_/B _60944_/Y sky130_fd_sc_hd__o21ai_4
X_79486_ _79483_/X _79486_/B _79486_/C _79487_/A sky130_fd_sc_hd__and3_4
X_45878_ _64190_/A _61695_/A sky130_fd_sc_hd__buf_2
X_76698_ _76688_/A _76687_/Y _76698_/Y sky130_fd_sc_hd__nor2_4
X_47617_ _47595_/A _47645_/B _47614_/X _53151_/D _47617_/X sky130_fd_sc_hd__and4_4
X_66451_ _66445_/A _66402_/B _66450_/Y _66451_/Y sky130_fd_sc_hd__nor3_4
X_78437_ _78439_/B _78439_/C _78436_/Y _78450_/A sky130_fd_sc_hd__a21boi_4
X_44829_ _41692_/Y _44817_/X _67605_/B _44818_/X _86932_/D sky130_fd_sc_hd__a2bb2o_4
X_63663_ _63670_/A _63670_/B _80357_/B _63663_/Y sky130_fd_sc_hd__nor3_4
X_75649_ _75649_/A _75649_/Y sky130_fd_sc_hd__inv_2
X_48597_ _81772_/Q _48959_/B _48597_/X sky130_fd_sc_hd__or2_4
X_60875_ _60870_/X _64172_/B _64172_/D _60881_/B sky130_fd_sc_hd__nand3_4
X_65402_ _65350_/X _86146_/Q _65400_/X _65401_/X _65402_/X sky130_fd_sc_hd__a211o_4
X_62614_ _62634_/A _62614_/B _62612_/Y _62613_/Y _62614_/Y sky130_fd_sc_hd__nand4_4
X_69170_ _87037_/Q _69153_/X _69168_/X _69169_/X _69170_/X sky130_fd_sc_hd__a211o_4
X_66382_ _64702_/X _66423_/B _64711_/X _66382_/Y sky130_fd_sc_hd__nand3_4
X_47548_ _47548_/A _53113_/D sky130_fd_sc_hd__buf_2
X_78368_ _78353_/A _78353_/C _78367_/Y _78369_/B sky130_fd_sc_hd__a21oi_4
X_63594_ _63471_/A _63595_/D sky130_fd_sc_hd__buf_2
Xclkbuf_10_332_0_CLK clkbuf_9_166_0_CLK/X _84746_/CLK sky130_fd_sc_hd__clkbuf_1
X_68121_ _67495_/X _68121_/X sky130_fd_sc_hd__buf_2
X_65333_ _65333_/A _65332_/X _65333_/Y sky130_fd_sc_hd__nand2_4
X_77319_ _77286_/A _77300_/A _77301_/A _77319_/X sky130_fd_sc_hd__a21o_4
X_62545_ _62544_/Y _59951_/C _84890_/Q _62196_/X _62545_/X sky130_fd_sc_hd__a2bb2o_4
X_47479_ _47525_/A _47517_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_962_0_CLK clkbuf_9_481_0_CLK/X _86238_/CLK sky130_fd_sc_hd__clkbuf_1
X_78299_ _82688_/Q _78299_/B _78299_/X sky130_fd_sc_hd__xor2_4
X_49218_ _49212_/A _50738_/B _49218_/Y sky130_fd_sc_hd__nand2_4
X_80330_ _80324_/A _80326_/X _80327_/Y _80330_/Y sky130_fd_sc_hd__nand3_4
X_68052_ _87893_/Q _68006_/X _67984_/X _68051_/X _68052_/X sky130_fd_sc_hd__a211o_4
X_65264_ _65289_/A _86408_/Q _65264_/X sky130_fd_sc_hd__and2_4
X_50490_ _86190_/Q _50464_/X _50489_/Y _50490_/Y sky130_fd_sc_hd__o21ai_4
X_62476_ _61549_/X _62492_/B _62449_/X _62475_/X _62476_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_9_453_0_CLK clkbuf_8_226_0_CLK/X clkbuf_9_453_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_67003_ _67028_/A _67003_/B _67003_/X sky130_fd_sc_hd__and2_4
X_64215_ _64490_/A _64490_/B _79883_/B _64215_/Y sky130_fd_sc_hd__nor3_4
X_61427_ _61375_/A _61427_/B _61398_/C _61427_/Y sky130_fd_sc_hd__nand3_4
X_49149_ _49128_/X _48654_/A _49148_/Y _52395_/B sky130_fd_sc_hd__a21o_4
X_80261_ _80261_/A _80261_/B _80261_/Y sky130_fd_sc_hd__nand2_4
X_65195_ _65529_/A _65195_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_347_0_CLK clkbuf_9_173_0_CLK/X _85428_/CLK sky130_fd_sc_hd__clkbuf_1
X_82000_ _82103_/CLK _82032_/Q _77114_/B sky130_fd_sc_hd__dfxtp_4
X_52160_ _51956_/X _52182_/C sky130_fd_sc_hd__buf_2
Xclkbuf_10_977_0_CLK clkbuf_9_488_0_CLK/X _86154_/CLK sky130_fd_sc_hd__clkbuf_1
X_64146_ _58198_/A _64158_/B _64158_/C _64045_/X _64146_/Y sky130_fd_sc_hd__nand4_4
X_61358_ _61358_/A _61367_/B _61367_/C _61367_/D _61358_/Y sky130_fd_sc_hd__nand4_4
X_80192_ _84947_/Q _65531_/C _80192_/Y sky130_fd_sc_hd__nand2_4
X_51111_ _51108_/Y _51093_/X _51110_/X _86072_/D sky130_fd_sc_hd__a21oi_4
X_60309_ _60170_/A _60253_/A _60309_/C _60309_/D _60309_/X sky130_fd_sc_hd__and4_4
X_52091_ _52100_/A _50389_/B _52091_/Y sky130_fd_sc_hd__nand2_4
X_68954_ _68586_/A _68954_/X sky130_fd_sc_hd__buf_2
X_64077_ _64076_/Y _64077_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_9_468_0_CLK clkbuf_9_469_0_CLK/A clkbuf_9_468_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_61289_ _72502_/A _72507_/A _72514_/A _61290_/A sky130_fd_sc_hd__and3_4
X_51042_ _51038_/Y _51039_/X _51041_/X _86085_/D sky130_fd_sc_hd__a21oi_4
X_67905_ _67902_/X _67904_/X _67858_/X _67905_/X sky130_fd_sc_hd__a21o_4
X_63028_ _60473_/C _63028_/X sky130_fd_sc_hd__buf_2
X_83951_ _81134_/CLK _83951_/D _83951_/Q sky130_fd_sc_hd__dfxtp_4
X_68885_ _87838_/Q _68886_/B sky130_fd_sc_hd__inv_2
Xclkbuf_10_900_0_CLK clkbuf_9_450_0_CLK/X _82536_/CLK sky130_fd_sc_hd__clkbuf_1
X_82902_ _81154_/CLK _78226_/B _82902_/Q sky130_fd_sc_hd__dfxtp_4
X_55850_ _55847_/X _55849_/X _44112_/X _55850_/X sky130_fd_sc_hd__a21o_4
X_67836_ _67739_/X _67836_/B _67836_/X sky130_fd_sc_hd__and2_4
X_86670_ _86351_/CLK _86670_/D _59240_/A sky130_fd_sc_hd__dfxtp_4
X_83882_ _82339_/CLK _83882_/D _83882_/Q sky130_fd_sc_hd__dfxtp_4
X_54801_ _85375_/Q _54784_/X _54800_/Y _54801_/Y sky130_fd_sc_hd__o21ai_4
X_85621_ _86554_/CLK _85621_/D _85621_/Q sky130_fd_sc_hd__dfxtp_4
X_82833_ _82833_/CLK _79348_/X _82833_/Q sky130_fd_sc_hd__dfxtp_4
X_67767_ _67790_/A _67767_/B _67767_/X sky130_fd_sc_hd__and2_4
X_55781_ _55778_/X _55780_/X _55781_/X sky130_fd_sc_hd__and2_4
X_52993_ _52997_/A _52997_/B _52997_/C _52993_/D _52993_/X sky130_fd_sc_hd__and4_4
X_64979_ _65607_/A _65056_/B sky130_fd_sc_hd__buf_2
X_57520_ _46401_/A _57531_/A sky130_fd_sc_hd__buf_2
X_69506_ _69315_/A _69506_/X sky130_fd_sc_hd__buf_2
X_88340_ _88327_/CLK _88340_/D _88340_/Q sky130_fd_sc_hd__dfxtp_4
X_54732_ _54731_/X _47420_/Y _54732_/Y sky130_fd_sc_hd__nand2_4
X_85552_ _83305_/CLK _53868_/Y _85552_/Q sky130_fd_sc_hd__dfxtp_4
X_66718_ _66669_/A _66718_/B _66718_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_915_0_CLK clkbuf_9_457_0_CLK/X _83141_/CLK sky130_fd_sc_hd__clkbuf_1
X_51944_ _52177_/A _52152_/A sky130_fd_sc_hd__buf_2
X_82764_ _82956_/CLK _82764_/D _82956_/D sky130_fd_sc_hd__dfxtp_4
X_67698_ _67698_/A _67698_/B _67698_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_4_0_CLK clkbuf_9_2_0_CLK/X _85168_/CLK sky130_fd_sc_hd__clkbuf_1
X_84503_ _84503_/CLK _84503_/D _84503_/Q sky130_fd_sc_hd__dfxtp_4
X_57451_ _57440_/X _57449_/X _57450_/Y _57452_/A sky130_fd_sc_hd__o21ai_4
X_81715_ _81514_/CLK _81339_/Q _81715_/Q sky130_fd_sc_hd__dfxtp_4
X_69437_ _81388_/D _69367_/X _69436_/X _83924_/D sky130_fd_sc_hd__a21bo_4
X_88271_ _88272_/CLK _41135_/X _68485_/B sky130_fd_sc_hd__dfxtp_4
X_54663_ _54661_/Y _54638_/X _54662_/X _85401_/D sky130_fd_sc_hd__a21oi_4
X_66649_ _88400_/Q _66593_/X _66594_/X _66648_/X _66649_/X sky130_fd_sc_hd__a211o_4
X_85483_ _84930_/CLK _85483_/D _85483_/Q sky130_fd_sc_hd__dfxtp_4
X_51875_ _51875_/A _51008_/B _51875_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_406_0_CLK clkbuf_9_407_0_CLK/A clkbuf_9_406_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_82695_ _82933_/CLK _78851_/X _78680_/B sky130_fd_sc_hd__dfxtp_4
X_56402_ _56055_/X _56394_/X _56401_/Y _85208_/D sky130_fd_sc_hd__o21ai_4
X_87222_ _87225_/CLK _87222_/D _87222_/Q sky130_fd_sc_hd__dfxtp_4
X_53614_ _50391_/A _53697_/B _53697_/C _53614_/Y sky130_fd_sc_hd__nand3_4
X_84434_ _81859_/CLK _62091_/Y _78057_/B sky130_fd_sc_hd__dfxtp_4
X_50826_ _50823_/Y _50801_/X _50825_/X _86126_/D sky130_fd_sc_hd__a21oi_4
X_81646_ _81296_/CLK _76907_/A _76314_/A sky130_fd_sc_hd__dfxtp_4
X_57382_ _44308_/X _57465_/A sky130_fd_sc_hd__inv_2
X_69368_ _69645_/A _69368_/X sky130_fd_sc_hd__buf_2
X_54594_ _54321_/A _54594_/X sky130_fd_sc_hd__buf_2
X_59121_ _59033_/A _59121_/X sky130_fd_sc_hd__buf_2
X_56333_ _56099_/X _56321_/X _56332_/Y _56333_/Y sky130_fd_sc_hd__o21ai_4
X_68319_ _68376_/A _68319_/X sky130_fd_sc_hd__buf_2
X_87153_ _87653_/CLK _87153_/D _87153_/Q sky130_fd_sc_hd__dfxtp_4
X_53545_ _53793_/A _53565_/A sky130_fd_sc_hd__buf_2
X_84365_ _84559_/CLK _62970_/Y _84365_/Q sky130_fd_sc_hd__dfxtp_4
X_50757_ _50771_/A _50757_/B _50757_/Y sky130_fd_sc_hd__nand2_4
X_81577_ _81344_/CLK _84177_/Q _76713_/A sky130_fd_sc_hd__dfxtp_4
X_69299_ _69065_/X _69299_/X sky130_fd_sc_hd__buf_2
X_86104_ _86104_/CLK _50935_/Y _86104_/Q sky130_fd_sc_hd__dfxtp_4
X_40510_ _40509_/X _40510_/X sky130_fd_sc_hd__buf_2
X_59052_ _59001_/X _86077_/Q _59051_/X _59052_/Y sky130_fd_sc_hd__o21ai_4
X_71330_ _50370_/B _71320_/X _71329_/Y _83534_/D sky130_fd_sc_hd__o21ai_4
X_83316_ _83316_/CLK _83316_/D _83316_/Q sky130_fd_sc_hd__dfxtp_4
X_56264_ _56153_/X _56255_/X _56263_/Y _85254_/D sky130_fd_sc_hd__o21ai_4
X_80528_ _80542_/A _80527_/Y _80551_/A sky130_fd_sc_hd__xor2_4
X_87084_ _88263_/CLK _44488_/Y _87084_/Q sky130_fd_sc_hd__dfxtp_4
X_53476_ _53448_/X _53476_/X sky130_fd_sc_hd__buf_2
X_41490_ _41490_/A _41490_/X sky130_fd_sc_hd__buf_2
X_84296_ _84671_/CLK _84296_/D _80241_/B sky130_fd_sc_hd__dfxtp_4
X_50688_ _50640_/A _72079_/B _50688_/Y sky130_fd_sc_hd__nand2_4
X_58003_ _58939_/A _58003_/X sky130_fd_sc_hd__buf_2
X_55215_ _55212_/X _55214_/X _55138_/A _72718_/C sky130_fd_sc_hd__a21o_4
X_86035_ _86424_/CLK _86035_/D _86035_/Q sky130_fd_sc_hd__dfxtp_4
X_40441_ _40437_/X _40364_/X _40440_/X _88391_/Q _40375_/X _40441_/Y
+ sky130_fd_sc_hd__o32ai_4
X_52427_ _52425_/Y _52415_/X _52426_/Y _85825_/D sky130_fd_sc_hd__a21oi_4
X_71261_ _71258_/A _71261_/B _71141_/B _71261_/Y sky130_fd_sc_hd__nand3_4
X_83247_ _84835_/CLK _83247_/D _62005_/A sky130_fd_sc_hd__dfxtp_4
X_80459_ _80445_/Y _80451_/B _80458_/X _80460_/B sky130_fd_sc_hd__o21ai_4
X_56195_ _56194_/X _56195_/X sky130_fd_sc_hd__buf_2
X_73000_ _87818_/Q _73000_/B _73000_/Y sky130_fd_sc_hd__nor2_4
X_70212_ _70214_/A _70214_/B _83195_/Q _70204_/X _70212_/X sky130_fd_sc_hd__and4_4
Xclkbuf_6_6_0_CLK clkbuf_6_7_0_CLK/A clkbuf_6_6_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_43160_ _43160_/A _43160_/Y sky130_fd_sc_hd__inv_2
X_55146_ _45745_/A _44059_/A _55140_/X _55145_/Y _55146_/X sky130_fd_sc_hd__a211o_4
X_40372_ _40344_/A _40361_/A _40372_/B1 _44624_/A sky130_fd_sc_hd__a21o_4
X_52358_ _65094_/B _52347_/X _52357_/Y _52358_/Y sky130_fd_sc_hd__o21ai_4
X_71192_ _71211_/A _71197_/A sky130_fd_sc_hd__buf_2
X_83178_ _81696_/CLK _72719_/X _83178_/Q sky130_fd_sc_hd__dfxtp_4
X_42111_ _42099_/X _42094_/X _41054_/X _88030_/Q _42096_/X _42112_/A
+ sky130_fd_sc_hd__o32ai_4
X_51309_ _51259_/A _51309_/X sky130_fd_sc_hd__buf_2
X_70143_ _83516_/Q _83164_/Q _83513_/Q _83161_/Q _70144_/D sky130_fd_sc_hd__a22oi_4
X_82129_ _81989_/CLK _82129_/D _77265_/B sky130_fd_sc_hd__dfxtp_4
X_59954_ _60422_/A _61587_/B sky130_fd_sc_hd__buf_2
X_43091_ _43085_/X _43086_/X _40716_/X _43089_/Y _43090_/X _87580_/D
+ sky130_fd_sc_hd__o32ai_4
X_55077_ _54973_/A _55083_/C sky130_fd_sc_hd__buf_2
X_52289_ _52262_/A _52289_/X sky130_fd_sc_hd__buf_2
X_87986_ _82906_/CLK _87986_/D _87986_/Q sky130_fd_sc_hd__dfxtp_4
X_42042_ _42035_/X _42010_/X _40890_/X _42041_/Y _42037_/X _88060_/D
+ sky130_fd_sc_hd__o32ai_4
X_58905_ _58904_/X _85767_/Q _58838_/X _58905_/X sky130_fd_sc_hd__o21a_4
X_54028_ _54020_/A _46455_/Y _54028_/Y sky130_fd_sc_hd__nand2_4
X_86937_ _87471_/CLK _86937_/D _86937_/Q sky130_fd_sc_hd__dfxtp_4
X_74951_ _81137_/D _80849_/Q _74961_/B sky130_fd_sc_hd__nand2_4
X_70074_ _68992_/X _68995_/X _69156_/X _70074_/Y sky130_fd_sc_hd__a21oi_4
X_59885_ _59532_/A _59520_/A _59535_/A _59885_/Y sky130_fd_sc_hd__nand3_4
X_73902_ _73850_/X _86227_/Q _73804_/X _73901_/X _73902_/X sky130_fd_sc_hd__a211o_4
X_46850_ _46850_/A _52713_/B sky130_fd_sc_hd__inv_2
X_58836_ _58730_/X _85932_/Q _58810_/X _58836_/X sky130_fd_sc_hd__o21a_4
X_77670_ _77662_/Y _77695_/B _82206_/D sky130_fd_sc_hd__xor2_4
X_74882_ _81127_/D _74875_/B _74882_/Y sky130_fd_sc_hd__nor2_4
X_86868_ _84408_/CLK _86868_/D _63137_/B sky130_fd_sc_hd__dfxtp_4
X_45801_ _45801_/A _45832_/B sky130_fd_sc_hd__buf_2
X_76621_ _76619_/Y _76620_/X _76621_/X sky130_fd_sc_hd__xor2_4
X_73833_ _73742_/A _73833_/B _73833_/X sky130_fd_sc_hd__and2_4
X_85819_ _85822_/CLK _52455_/Y _85819_/Q sky130_fd_sc_hd__dfxtp_4
X_46781_ _86704_/Q _46767_/X _46780_/Y _46781_/Y sky130_fd_sc_hd__o21ai_4
X_58767_ _58748_/X _58763_/Y _58764_/Y _58766_/X _58752_/X _58767_/X
+ sky130_fd_sc_hd__o32a_4
X_43993_ _43989_/Y _43955_/Y _43992_/Y _43994_/A sky130_fd_sc_hd__a21oi_4
X_55979_ _56379_/C _55690_/A _55611_/X _55978_/X _55979_/X sky130_fd_sc_hd__a211o_4
X_86799_ _87990_/CLK _86799_/D _86799_/Q sky130_fd_sc_hd__dfxtp_4
X_48520_ _48520_/A _48565_/B _48520_/Y sky130_fd_sc_hd__nand2_4
X_79340_ _84800_/Q _84120_/Q _79340_/Y sky130_fd_sc_hd__nand2_4
X_45732_ _45725_/X _45729_/Y _45731_/Y _45732_/Y sky130_fd_sc_hd__a21oi_4
X_57718_ _57718_/A _57718_/X sky130_fd_sc_hd__buf_2
X_76552_ _76552_/A _81545_/Q _76552_/Y sky130_fd_sc_hd__nand2_4
X_42944_ _42846_/X _42944_/X sky130_fd_sc_hd__buf_2
X_73764_ _73764_/A _73764_/B _73765_/B sky130_fd_sc_hd__nand2_4
X_70976_ _70976_/A _70954_/B _70969_/C _70976_/Y sky130_fd_sc_hd__nand3_4
X_58698_ _58698_/A _58699_/A sky130_fd_sc_hd__buf_2
X_75503_ _75503_/A _75503_/B _75503_/C _75503_/Y sky130_fd_sc_hd__nand3_4
X_48451_ _74406_/A _48752_/A sky130_fd_sc_hd__buf_2
X_72715_ _83180_/Q _72702_/X _72714_/Y _83180_/D sky130_fd_sc_hd__a21bo_4
X_79271_ _79270_/B _79257_/Y _79271_/Y sky130_fd_sc_hd__nand2_4
X_57649_ _57647_/Y _57627_/X _57648_/Y _84962_/D sky130_fd_sc_hd__a21boi_4
X_45663_ _57283_/B _45326_/X _45662_/X _45663_/Y sky130_fd_sc_hd__o21ai_4
X_76483_ _76482_/A _76463_/X _76461_/X _76483_/Y sky130_fd_sc_hd__a21oi_4
X_42875_ _42945_/A _42875_/X sky130_fd_sc_hd__buf_2
X_73695_ _73693_/X _73694_/Y _73546_/X _73695_/X sky130_fd_sc_hd__a21o_4
X_47402_ _83734_/Q _47403_/A sky130_fd_sc_hd__inv_2
X_78222_ _78220_/B _78203_/A _82492_/Q _78222_/Y sky130_fd_sc_hd__nand3_4
X_44614_ _44613_/Y _87032_/D sky130_fd_sc_hd__inv_2
X_75434_ _75433_/X _75466_/B sky130_fd_sc_hd__buf_2
X_41826_ _41824_/X _41825_/X _40446_/X _66892_/B _41821_/X _41826_/Y
+ sky130_fd_sc_hd__o32ai_4
X_48382_ _72817_/B _48350_/X _48381_/Y _48382_/Y sky130_fd_sc_hd__o21ai_4
X_60660_ _60660_/A _60660_/X sky130_fd_sc_hd__buf_2
X_72646_ _72687_/A _72656_/A sky130_fd_sc_hd__buf_2
X_45594_ _45587_/X _45590_/X _45593_/Y _45594_/Y sky130_fd_sc_hd__a21oi_4
X_47333_ _47147_/A _47333_/X sky130_fd_sc_hd__buf_2
X_59319_ _59273_/X _85639_/Q _59308_/X _59319_/X sky130_fd_sc_hd__o21a_4
X_78153_ _82668_/Q _78153_/B _78153_/X sky130_fd_sc_hd__xor2_4
X_44545_ _44496_/X _44497_/X _40826_/X _87059_/Q _44498_/X _44545_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75365_ _75364_/Y _75365_/Y sky130_fd_sc_hd__inv_2
X_41757_ _41756_/X _41757_/X sky130_fd_sc_hd__buf_2
X_60591_ _79132_/A _60132_/X _60551_/X _60590_/Y _60591_/X sky130_fd_sc_hd__a2bb2o_4
X_72577_ _72576_/Y _72577_/B _72569_/A _72577_/Y sky130_fd_sc_hd__nand3_4
X_77104_ _77105_/A _81913_/Q _77106_/A sky130_fd_sc_hd__or2_4
X_62330_ _62304_/A _57652_/X _62315_/C _62286_/X _62330_/X sky130_fd_sc_hd__and4_4
X_74316_ _74342_/A _74325_/B sky130_fd_sc_hd__buf_2
X_40708_ _40687_/X _40688_/X _40707_/X _68892_/B _40683_/X _40709_/A
+ sky130_fd_sc_hd__o32ai_4
X_47264_ _47264_/A _52948_/D sky130_fd_sc_hd__buf_2
X_71528_ _71527_/Y _71528_/X sky130_fd_sc_hd__buf_2
X_78084_ _82563_/Q _78091_/B _78084_/X sky130_fd_sc_hd__xor2_4
X_44476_ _41189_/A _44474_/X _87089_/Q _44475_/X _44476_/X sky130_fd_sc_hd__a2bb2o_4
X_75296_ _75294_/Y _75295_/X _81041_/D sky130_fd_sc_hd__xnor2_4
X_41688_ _41687_/X _41688_/X sky130_fd_sc_hd__buf_2
X_49003_ _49052_/A _49003_/X sky130_fd_sc_hd__buf_2
X_46215_ _46207_/Y _46215_/B _46215_/C _46216_/A sky130_fd_sc_hd__nand3_4
X_77035_ _77036_/A _77036_/B _77035_/Y sky130_fd_sc_hd__nand2_4
XPHY_270 sky130_fd_sc_hd__decap_3
X_43427_ _43422_/X _43426_/X _41545_/X _87427_/Q _43407_/X _43428_/A
+ sky130_fd_sc_hd__o32ai_4
X_62261_ _62249_/A _63396_/B _59987_/X _62261_/Y sky130_fd_sc_hd__nand3_4
X_74247_ _43107_/Y _72900_/X _73920_/X _74246_/Y _74247_/X sky130_fd_sc_hd__a211o_4
X_40639_ _40639_/A _40654_/B _40639_/X sky130_fd_sc_hd__or2_4
XPHY_281 sky130_fd_sc_hd__decap_3
X_47195_ _47195_/A _47195_/X sky130_fd_sc_hd__buf_2
X_71459_ _71444_/Y _83491_/Q _71458_/Y _71459_/X sky130_fd_sc_hd__a21o_4
XPHY_292 sky130_fd_sc_hd__decap_3
X_64000_ _61980_/A _64046_/B _64046_/C _64016_/D _64001_/D sky130_fd_sc_hd__nand4_4
X_61212_ _61254_/B _60296_/X _61238_/C _61212_/Y sky130_fd_sc_hd__nand3_4
X_46146_ _40591_/C _49793_/A sky130_fd_sc_hd__buf_2
X_43358_ _41352_/X _43356_/X _87463_/Q _43357_/X _87463_/D sky130_fd_sc_hd__a2bb2o_4
X_62192_ _62190_/Y _62166_/X _62191_/Y _62192_/Y sky130_fd_sc_hd__a21oi_4
X_74178_ _74155_/X _84967_/Q _74087_/X _74177_/X _74179_/B sky130_fd_sc_hd__a211o_4
Xpsn_inst_psn_buff_19 _56456_/A _56370_/C sky130_fd_sc_hd__buf_8
X_42309_ _42308_/Y _87929_/D sky130_fd_sc_hd__inv_2
X_61143_ _61140_/X _61179_/A _61172_/A _64250_/C _64210_/A sky130_fd_sc_hd__nand4_4
X_73129_ _72973_/B _73129_/X sky130_fd_sc_hd__buf_2
X_46077_ _46067_/X _43046_/A _41605_/X _86778_/Q _46068_/X _46077_/Y
+ sky130_fd_sc_hd__o32ai_4
X_43289_ _41165_/X _43287_/X _87497_/Q _43288_/X _43289_/X sky130_fd_sc_hd__a2bb2o_4
X_78986_ _78969_/A _78986_/B _78986_/X sky130_fd_sc_hd__and2_4
X_49905_ _49902_/Y _49897_/X _49904_/X _49905_/Y sky130_fd_sc_hd__a21oi_4
X_45028_ _56488_/C _44982_/X _44959_/X _45028_/X sky130_fd_sc_hd__o21a_4
X_65951_ _65896_/A _86558_/Q _65951_/X sky130_fd_sc_hd__and2_4
X_61074_ _61074_/A _61083_/B sky130_fd_sc_hd__buf_2
X_77937_ _77935_/Y _77946_/A _77941_/A sky130_fd_sc_hd__xor2_4
X_64902_ _64902_/A _64902_/X sky130_fd_sc_hd__buf_2
X_60025_ _59943_/X _60025_/X sky130_fd_sc_hd__buf_2
X_49836_ _49833_/Y _49815_/X _49835_/X _49836_/Y sky130_fd_sc_hd__a21oi_4
X_68670_ _73842_/A _68414_/X _68379_/X _68669_/Y _68670_/X sky130_fd_sc_hd__a211o_4
X_65882_ _65825_/A _86499_/Q _65882_/X sky130_fd_sc_hd__and2_4
X_77868_ _77851_/A _77866_/Y _77867_/Y _77868_/Y sky130_fd_sc_hd__a21oi_4
X_67621_ _67696_/A _88231_/Q _67621_/X sky130_fd_sc_hd__and2_4
X_79607_ _79607_/A _79607_/B _79609_/B sky130_fd_sc_hd__nand2_4
X_76819_ _76819_/A _76819_/B _76819_/X sky130_fd_sc_hd__xor2_4
X_64833_ _64731_/A _64834_/A sky130_fd_sc_hd__buf_2
X_49767_ _49764_/Y _49759_/X _49766_/X _49767_/Y sky130_fd_sc_hd__a21oi_4
X_46979_ _82395_/Q _46979_/Y sky130_fd_sc_hd__inv_2
X_77799_ _77787_/A _77786_/X _77799_/X sky130_fd_sc_hd__or2_4
X_48718_ _65441_/B _48150_/X _48717_/Y _48718_/Y sky130_fd_sc_hd__o21ai_4
X_67552_ _67312_/X _67552_/X sky130_fd_sc_hd__buf_2
X_79538_ _79538_/A _79538_/Y sky130_fd_sc_hd__inv_2
X_64764_ _64870_/A _64741_/B _64764_/C _64764_/Y sky130_fd_sc_hd__nor3_4
X_49698_ _49695_/Y _49677_/X _49697_/X _49698_/Y sky130_fd_sc_hd__a21oi_4
X_61976_ _61820_/A _62002_/B sky130_fd_sc_hd__buf_2
X_66503_ _65305_/X _66521_/B _65311_/X _66503_/Y sky130_fd_sc_hd__nand3_4
X_63715_ _60798_/X _63713_/Y _63358_/X _63714_/Y _63715_/X sky130_fd_sc_hd__a211o_4
X_60927_ _60844_/X _60857_/D _61293_/A _60861_/X _60928_/A sky130_fd_sc_hd__and4_4
X_48649_ _48661_/A _48847_/B _48649_/Y sky130_fd_sc_hd__nand2_4
X_79469_ _79484_/A _79484_/B _79480_/A sky130_fd_sc_hd__xor2_4
X_67483_ _87161_/Q _67432_/X _67433_/X _67482_/X _67483_/X sky130_fd_sc_hd__a211o_4
X_64695_ _64691_/X _86141_/Q _64692_/X _64694_/X _64695_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_271_0_CLK clkbuf_9_135_0_CLK/X _83491_/CLK sky130_fd_sc_hd__clkbuf_1
X_81500_ _84064_/CLK _81500_/D _81500_/Q sky130_fd_sc_hd__dfxtp_4
X_69222_ _69219_/X _69221_/X _69025_/X _69222_/X sky130_fd_sc_hd__a21o_4
X_66434_ _66432_/Y _66414_/X _66433_/X _84124_/D sky130_fd_sc_hd__a21o_4
X_51660_ _51671_/A _53183_/B _51660_/Y sky130_fd_sc_hd__nand2_4
X_63646_ _63670_/A _63670_/B _80379_/B _63646_/Y sky130_fd_sc_hd__nor3_4
X_82480_ _82563_/CLK _78520_/X _78125_/B sky130_fd_sc_hd__dfxtp_4
X_60858_ _60857_/X _60915_/A sky130_fd_sc_hd__buf_2
X_50611_ _50608_/Y _50609_/X _50610_/X _50611_/Y sky130_fd_sc_hd__a21oi_4
X_81431_ _81431_/CLK _81463_/Q _76070_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_53_0_CLK clkbuf_9_26_0_CLK/X _85128_/CLK sky130_fd_sc_hd__clkbuf_1
X_69153_ _68394_/A _69153_/X sky130_fd_sc_hd__buf_2
X_66365_ _66362_/Y _66343_/X _66364_/X _84137_/D sky130_fd_sc_hd__a21o_4
X_51591_ _85982_/Q _51566_/X _51590_/Y _51591_/Y sky130_fd_sc_hd__o21ai_4
X_63577_ _64328_/A _63578_/A sky130_fd_sc_hd__buf_2
X_60789_ _60792_/A _60761_/B _60789_/C _60789_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_9_392_0_CLK clkbuf_9_393_0_CLK/A clkbuf_9_392_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_68104_ _82078_/D _68101_/X _68103_/X _84038_/D sky130_fd_sc_hd__a21bo_4
X_53330_ _53330_/A _53330_/B _53330_/C _52811_/D _53330_/X sky130_fd_sc_hd__and4_4
X_65316_ _64696_/X _85542_/Q _64697_/X _65315_/X _65316_/X sky130_fd_sc_hd__a211o_4
X_84150_ _84150_/CLK _84150_/D _84150_/Q sky130_fd_sc_hd__dfxtp_4
X_50542_ _86181_/Q _50533_/X _50541_/Y _50542_/Y sky130_fd_sc_hd__o21ai_4
X_62528_ _62526_/Y _62467_/X _62527_/Y _62528_/Y sky130_fd_sc_hd__a21oi_4
X_81362_ _81362_/CLK _81362_/D _81362_/Q sky130_fd_sc_hd__dfxtp_4
X_69084_ _68907_/X _68882_/X _69075_/Y _69083_/Y _69084_/X sky130_fd_sc_hd__a211o_4
X_66296_ _66267_/X _66296_/B _66296_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_286_0_CLK clkbuf_9_143_0_CLK/X _82386_/CLK sky130_fd_sc_hd__clkbuf_1
X_83101_ _83846_/CLK _74318_/X _70301_/C sky130_fd_sc_hd__dfxtp_4
X_80313_ _80313_/A _80313_/Y sky130_fd_sc_hd__inv_2
X_68035_ _68371_/A _88214_/Q _68035_/X sky130_fd_sc_hd__and2_4
X_53261_ _53243_/X _51747_/A _53266_/C _53261_/D _53261_/X sky130_fd_sc_hd__and4_4
X_65247_ _65225_/A _65247_/B _65247_/X sky130_fd_sc_hd__and2_4
X_84081_ _83933_/CLK _67165_/X _84081_/Q sky130_fd_sc_hd__dfxtp_4
X_50473_ _50473_/A _50577_/A sky130_fd_sc_hd__buf_2
X_62459_ _62448_/A _58474_/A _62491_/C _62461_/C sky130_fd_sc_hd__nand3_4
X_81293_ _81260_/CLK _76981_/X _81261_/D sky130_fd_sc_hd__dfxtp_4
X_55000_ _55013_/A _54978_/X _55013_/C _47594_/A _55000_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_68_0_CLK clkbuf_9_34_0_CLK/X _86861_/CLK sky130_fd_sc_hd__clkbuf_1
X_52212_ _50511_/A _52198_/X _52218_/C _52212_/X sky130_fd_sc_hd__and3_4
X_83032_ _85180_/CLK _74567_/Y _45046_/A sky130_fd_sc_hd__dfxtp_4
X_80244_ _80244_/A _80244_/B _80244_/Y sky130_fd_sc_hd__nand2_4
X_53192_ _53188_/Y _53189_/X _53191_/X _53192_/Y sky130_fd_sc_hd__a21oi_4
X_65178_ _64809_/A _65178_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_214_0_CLK clkbuf_8_215_0_CLK/A clkbuf_9_429_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_52143_ _52127_/X _50440_/B _52143_/Y sky130_fd_sc_hd__nand2_4
X_64129_ _63912_/X _64129_/X sky130_fd_sc_hd__buf_2
X_87840_ _88104_/CLK _42510_/Y _74005_/A sky130_fd_sc_hd__dfxtp_4
X_80175_ _60021_/C _63864_/C _80175_/X sky130_fd_sc_hd__xor2_4
X_69986_ _69599_/Y _69916_/X _69984_/X _69985_/Y _69986_/X sky130_fd_sc_hd__a211o_4
X_52074_ _52126_/A _52438_/A sky130_fd_sc_hd__buf_2
X_56951_ _56940_/Y _56952_/A sky130_fd_sc_hd__inv_2
X_68937_ _68932_/X _68936_/X _68773_/X _68937_/X sky130_fd_sc_hd__a21o_4
X_87771_ _87273_/CLK _42684_/X _69466_/B sky130_fd_sc_hd__dfxtp_4
X_84983_ _86587_/CLK _84983_/D _84983_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_330_0_CLK clkbuf_9_331_0_CLK/A clkbuf_9_330_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_51025_ _51023_/Y _51011_/X _51024_/X _51025_/Y sky130_fd_sc_hd__a21oi_4
X_55902_ _55902_/A _55901_/X _55928_/B sky130_fd_sc_hd__and2_4
X_86722_ _86733_/CLK _86722_/D _86722_/Q sky130_fd_sc_hd__dfxtp_4
X_59670_ _64738_/A _66046_/A sky130_fd_sc_hd__buf_2
X_83934_ _81346_/CLK _83934_/D _81398_/D sky130_fd_sc_hd__dfxtp_4
X_56882_ _55654_/X _55672_/X _56881_/X _56885_/A sky130_fd_sc_hd__o21ai_4
X_68868_ _68779_/A _68868_/B _68868_/X sky130_fd_sc_hd__and2_4
Xclkbuf_8_229_0_CLK clkbuf_8_229_0_CLK/A clkbuf_9_459_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_224_0_CLK clkbuf_9_112_0_CLK/X _80696_/CLK sky130_fd_sc_hd__clkbuf_1
X_58621_ _58617_/Y _58620_/Y _58610_/X _58621_/X sky130_fd_sc_hd__a21o_4
X_55833_ _55836_/A _55833_/B _55833_/X sky130_fd_sc_hd__and2_4
X_67819_ _87903_/Q _67770_/X _67748_/X _67818_/X _67819_/X sky130_fd_sc_hd__a211o_4
X_86653_ _86651_/CLK _47266_/Y _57792_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_854_0_CLK clkbuf_9_427_0_CLK/X _86422_/CLK sky130_fd_sc_hd__clkbuf_1
X_83865_ _82541_/CLK _70043_/X _82545_/D sky130_fd_sc_hd__dfxtp_4
X_68799_ _66673_/X _69478_/A sky130_fd_sc_hd__buf_2
X_85604_ _86203_/CLK _85604_/D _85604_/Q sky130_fd_sc_hd__dfxtp_4
X_70830_ _70698_/A _70830_/B _70830_/Y sky130_fd_sc_hd__nor2_4
X_58552_ _58538_/X _83357_/Q _58551_/Y _84821_/D sky130_fd_sc_hd__o21a_4
X_82816_ _82740_/CLK _82848_/Q _82816_/Q sky130_fd_sc_hd__dfxtp_4
X_55764_ _55224_/A _55764_/B _55764_/X sky130_fd_sc_hd__and2_4
X_86584_ _86587_/CLK _86584_/D _66037_/B sky130_fd_sc_hd__dfxtp_4
X_52976_ _52893_/X _52997_/A sky130_fd_sc_hd__buf_2
X_40990_ _40986_/X _40987_/X _69279_/B _40989_/X _88297_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_9_345_0_CLK clkbuf_9_345_0_CLK/A clkbuf_9_345_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_83796_ _83787_/CLK _83796_/D _83796_/Q sky130_fd_sc_hd__dfxtp_4
X_57503_ _47819_/A _47863_/Y _57503_/Y sky130_fd_sc_hd__nand2_4
X_88323_ _88060_/CLK _88323_/D _88323_/Q sky130_fd_sc_hd__dfxtp_4
X_54715_ _85391_/Q _54703_/X _54714_/Y _54715_/Y sky130_fd_sc_hd__o21ai_4
X_85535_ _85535_/CLK _85535_/D _85535_/Q sky130_fd_sc_hd__dfxtp_4
X_51927_ _52398_/A _52126_/A sky130_fd_sc_hd__buf_2
X_70761_ _70761_/A _70761_/X sky130_fd_sc_hd__buf_2
X_82747_ _82748_/CLK _84131_/Q _82747_/Q sky130_fd_sc_hd__dfxtp_4
X_58483_ _58483_/A _58502_/B _58483_/Y sky130_fd_sc_hd__nor2_4
X_55695_ _55695_/A _85185_/Q _55695_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_239_0_CLK clkbuf_9_119_0_CLK/X _82220_/CLK sky130_fd_sc_hd__clkbuf_1
X_72500_ _64473_/A _72498_/B _72500_/Y sky130_fd_sc_hd__nand2_4
X_57434_ _57434_/A _57434_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_869_0_CLK clkbuf_9_434_0_CLK/X _85507_/CLK sky130_fd_sc_hd__clkbuf_1
X_88254_ _88006_/CLK _41227_/Y _88254_/Q sky130_fd_sc_hd__dfxtp_4
X_42660_ _42659_/Y _42660_/Y sky130_fd_sc_hd__inv_2
X_54646_ _54642_/Y _54638_/X _54645_/X _54646_/Y sky130_fd_sc_hd__a21oi_4
X_73480_ _73481_/B _73481_/C _73479_/X _73480_/X sky130_fd_sc_hd__a21o_4
X_85466_ _82961_/CLK _54308_/Y _85466_/Q sky130_fd_sc_hd__dfxtp_4
X_51858_ _85933_/Q _51846_/X _51857_/Y _51858_/Y sky130_fd_sc_hd__o21ai_4
X_70692_ _70692_/A _70692_/B _70692_/C _70692_/Y sky130_fd_sc_hd__nor3_4
X_82678_ _81216_/CLK _82678_/D _78226_/A sky130_fd_sc_hd__dfxtp_4
X_41611_ _41336_/X _41611_/X sky130_fd_sc_hd__buf_2
X_87205_ _87394_/CLK _43909_/X _67667_/B sky130_fd_sc_hd__dfxtp_4
X_72431_ _72419_/X _85351_/Q _72430_/X _72431_/Y sky130_fd_sc_hd__o21ai_4
X_84417_ _84414_/CLK _84417_/D _76993_/B sky130_fd_sc_hd__dfxtp_4
X_50809_ _50807_/Y _50792_/X _50808_/Y _50809_/Y sky130_fd_sc_hd__a21boi_4
X_57365_ _57261_/X _57362_/X _57364_/X _85028_/D sky130_fd_sc_hd__a21o_4
X_81629_ _81632_/CLK _76564_/X _81821_/D sky130_fd_sc_hd__dfxtp_4
X_88185_ _87417_/CLK _88185_/D _88185_/Q sky130_fd_sc_hd__dfxtp_4
X_42591_ _42429_/A _42592_/A sky130_fd_sc_hd__buf_2
X_54577_ _54574_/Y _54558_/X _54576_/X _54577_/Y sky130_fd_sc_hd__a21oi_4
X_85397_ _85492_/CLK _54686_/Y _85397_/Q sky130_fd_sc_hd__dfxtp_4
X_51789_ _51789_/A _51789_/X sky130_fd_sc_hd__buf_2
X_59104_ _58858_/X _85432_/Q _59103_/X _59104_/Y sky130_fd_sc_hd__o21ai_4
X_44330_ _44381_/A _44330_/X sky130_fd_sc_hd__buf_2
X_56316_ _56060_/X _56305_/X _56315_/Y _56316_/Y sky130_fd_sc_hd__o21ai_4
X_75150_ _80775_/Q _81031_/D _80743_/D sky130_fd_sc_hd__xor2_4
X_87136_ _87137_/CLK _44387_/Y _87136_/Q sky130_fd_sc_hd__dfxtp_4
X_41542_ _40413_/X _41604_/A sky130_fd_sc_hd__buf_2
X_53528_ _85619_/Q _53506_/X _53527_/Y _53528_/Y sky130_fd_sc_hd__o21ai_4
X_72362_ _64591_/X _72362_/X sky130_fd_sc_hd__buf_2
X_84348_ _83227_/CLK _63163_/X _79372_/A sky130_fd_sc_hd__dfxtp_4
X_57296_ _56766_/X _56782_/X _56735_/X _57319_/D _56733_/X _57296_/Y
+ sky130_fd_sc_hd__a41oi_4
X_74101_ _44727_/Y _73491_/X _74100_/Y _74102_/B sky130_fd_sc_hd__a21o_4
X_59035_ _59033_/X _85438_/Q _59034_/X _59035_/Y sky130_fd_sc_hd__o21ai_4
X_71313_ _70400_/A _71313_/X sky130_fd_sc_hd__buf_2
X_44261_ _64642_/A _44261_/X sky130_fd_sc_hd__buf_2
X_56247_ _56114_/X _56242_/X _56246_/Y _56247_/Y sky130_fd_sc_hd__o21ai_4
X_75081_ _80770_/Q _81026_/D _75081_/X sky130_fd_sc_hd__xor2_4
X_41473_ _41472_/X _41473_/X sky130_fd_sc_hd__buf_2
X_87067_ _88327_/CLK _87067_/D _87067_/Q sky130_fd_sc_hd__dfxtp_4
X_53459_ _53454_/Y _53455_/X _53458_/Y _53459_/Y sky130_fd_sc_hd__a21boi_4
X_72293_ _72289_/Y _72291_/Y _72292_/X _72293_/X sky130_fd_sc_hd__a21o_4
X_84279_ _84273_/CLK _84279_/D _64037_/C sky130_fd_sc_hd__dfxtp_4
X_46000_ _45999_/Y _86821_/D sky130_fd_sc_hd__inv_2
X_43212_ _43212_/A _43212_/X sky130_fd_sc_hd__buf_2
X_74032_ _68859_/B _73891_/X _73962_/X _74031_/Y _74032_/X sky130_fd_sc_hd__a211o_4
X_86018_ _85953_/CLK _51397_/Y _65413_/B sky130_fd_sc_hd__dfxtp_4
X_40424_ _82327_/Q _40907_/B _40424_/X sky130_fd_sc_hd__or2_4
X_71244_ _57489_/B _71239_/X _71243_/Y _71244_/Y sky130_fd_sc_hd__o21ai_4
X_44192_ _72838_/A _72745_/A sky130_fd_sc_hd__inv_2
X_56178_ _56175_/Y _56178_/B _56178_/Y sky130_fd_sc_hd__nand2_4
X_43143_ _43129_/X _43130_/X _40820_/X _43141_/Y _43142_/X _87560_/D
+ sky130_fd_sc_hd__o32ai_4
X_55129_ _55129_/A _55149_/A sky130_fd_sc_hd__buf_2
X_78840_ _78840_/A _78839_/X _78874_/A sky130_fd_sc_hd__xnor2_4
X_40355_ _40354_/X _40355_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_807_0_CLK clkbuf_9_403_0_CLK/X _82563_/CLK sky130_fd_sc_hd__clkbuf_1
X_71175_ _71175_/A _71173_/B _71181_/C _71178_/D _71175_/Y sky130_fd_sc_hd__nand4_4
X_70126_ _83505_/Q _83153_/Q _83145_/Q _83144_/Q _70125_/Y _70127_/D
+ sky130_fd_sc_hd__a2111oi_4
X_47951_ _53514_/B _48236_/B sky130_fd_sc_hd__buf_2
X_43074_ _43073_/Y _87586_/D sky130_fd_sc_hd__inv_2
X_59937_ _59936_/X _60042_/D sky130_fd_sc_hd__inv_2
X_78771_ _78771_/A _78772_/A sky130_fd_sc_hd__inv_2
X_75983_ _81707_/D _75991_/B _75986_/A sky130_fd_sc_hd__xor2_4
X_87969_ _87210_/CLK _87969_/D _87969_/Q sky130_fd_sc_hd__dfxtp_4
X_46902_ _46902_/A _46903_/A sky130_fd_sc_hd__buf_2
X_42025_ _42025_/A _42025_/X sky130_fd_sc_hd__buf_2
X_77722_ _82209_/D _77722_/B _77724_/A sky130_fd_sc_hd__nand2_4
X_74934_ _74942_/A _74933_/Y _74935_/B sky130_fd_sc_hd__xor2_4
X_70057_ _68863_/X _68866_/X _70044_/X _70057_/Y sky130_fd_sc_hd__a21oi_4
X_47882_ _47855_/A _51954_/B _47882_/Y sky130_fd_sc_hd__nand2_4
X_59868_ _63130_/A _59868_/X sky130_fd_sc_hd__buf_2
X_49621_ _49607_/X _52837_/B _49621_/Y sky130_fd_sc_hd__nand2_4
X_46833_ _52700_/B _51008_/B sky130_fd_sc_hd__buf_2
X_58819_ _86701_/Q _58873_/B _58819_/Y sky130_fd_sc_hd__nor2_4
X_77653_ _77652_/A _82110_/D _77653_/Y sky130_fd_sc_hd__nand2_4
X_74865_ _74865_/A _74865_/Y sky130_fd_sc_hd__inv_2
X_59799_ _59737_/A _59848_/B _80464_/A _59799_/Y sky130_fd_sc_hd__nor3_4
X_76604_ _76603_/X _76604_/Y sky130_fd_sc_hd__inv_2
X_49552_ _49416_/A _49580_/A sky130_fd_sc_hd__buf_2
X_61830_ _61398_/B _61795_/B _61795_/C _61778_/X _61830_/Y sky130_fd_sc_hd__nand4_4
X_73816_ _73814_/X _73815_/Y _73720_/X _73816_/X sky130_fd_sc_hd__a21o_4
X_46764_ _46737_/A _46784_/B _46784_/C _52661_/D _46764_/X sky130_fd_sc_hd__and4_4
X_77584_ _77584_/A _77584_/B _77584_/C _77584_/X sky130_fd_sc_hd__or3_4
X_43976_ _44072_/A _43944_/A _43945_/A _43975_/Y _43976_/X sky130_fd_sc_hd__a211o_4
X_74796_ _74796_/A _74796_/B _74796_/C _74769_/D _74796_/Y sky130_fd_sc_hd__nand4_4
X_48503_ _48503_/A _74428_/B sky130_fd_sc_hd__inv_2
X_79323_ _79336_/B _79322_/Y _79334_/A sky130_fd_sc_hd__xor2_4
X_45715_ _45710_/X _45713_/Y _45714_/X _45715_/Y sky130_fd_sc_hd__a21oi_4
X_76535_ _76531_/Y _76535_/B _76534_/Y _76535_/X sky130_fd_sc_hd__or3_4
X_42927_ _42916_/X _42917_/X _41735_/X _87647_/Q _42905_/X _42927_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49483_ _49467_/A _49500_/B _49467_/C _52698_/D _49483_/X sky130_fd_sc_hd__and4_4
X_61761_ _61354_/B _61795_/B _61761_/C _62130_/D _61761_/Y sky130_fd_sc_hd__nand4_4
X_73747_ _73745_/X _73727_/X _73730_/X _73747_/Y sky130_fd_sc_hd__nand3_4
X_46695_ _58672_/A _46672_/X _46694_/Y _46695_/Y sky130_fd_sc_hd__o21ai_4
X_70959_ _70506_/A _70959_/B _70959_/C _71115_/B _70959_/X sky130_fd_sc_hd__and4_4
X_63500_ _63488_/A _61909_/X _63500_/X sky130_fd_sc_hd__and2_4
X_48434_ _53651_/B _48435_/B sky130_fd_sc_hd__buf_2
X_60712_ _60722_/A _60712_/B _60711_/X _60820_/A sky130_fd_sc_hd__nand3_4
X_79254_ _79250_/Y _79253_/Y _82824_/D sky130_fd_sc_hd__xor2_4
X_45646_ _45643_/Y _45627_/X _45644_/X _45645_/Y _45646_/X sky130_fd_sc_hd__a211o_4
X_64480_ _64473_/Y _64477_/Y _64479_/Y _58465_/A _64213_/X _64480_/Y
+ sky130_fd_sc_hd__o32ai_4
X_76466_ _76429_/A _76430_/X _76440_/X _76482_/A sky130_fd_sc_hd__a21o_4
X_42858_ _42835_/X _42858_/X sky130_fd_sc_hd__buf_2
X_61692_ _61305_/A _61692_/B _61682_/C _61692_/Y sky130_fd_sc_hd__nand3_4
X_73678_ _68495_/B _73597_/X _73652_/X _73677_/Y _73678_/X sky130_fd_sc_hd__a211o_4
X_78205_ _78205_/A _78205_/B _78209_/A sky130_fd_sc_hd__nand2_4
X_63431_ _63368_/X _63424_/X _63425_/X _63429_/X _63430_/Y _63431_/Y
+ sky130_fd_sc_hd__o41ai_4
X_75417_ _75413_/X _75414_/Y _75416_/Y _75435_/B sky130_fd_sc_hd__a21o_4
X_41809_ _41808_/Y _88142_/D sky130_fd_sc_hd__inv_2
X_60643_ _59877_/X _59705_/X _60298_/C _60644_/C sky130_fd_sc_hd__a21boi_4
X_48365_ _53620_/A _48364_/X _48354_/X _48365_/X sky130_fd_sc_hd__and3_4
X_72629_ _72537_/Y _60123_/Y _72579_/Y _79158_/A _59868_/X _72629_/Y
+ sky130_fd_sc_hd__a32oi_4
X_79185_ _79185_/A _79185_/B _79185_/C _79188_/A sky130_fd_sc_hd__nand3_4
X_45577_ _45575_/Y _45576_/Y _44939_/B _45577_/X sky130_fd_sc_hd__o21a_4
X_76397_ _76392_/Y _76394_/Y _76398_/A sky130_fd_sc_hd__nor2_4
X_42789_ _41356_/X _42787_/X _87718_/Q _42788_/X _42789_/X sky130_fd_sc_hd__a2bb2o_4
X_47316_ _86647_/Q _47286_/X _47315_/Y _47316_/Y sky130_fd_sc_hd__o21ai_4
X_66150_ _66003_/A _66151_/B sky130_fd_sc_hd__buf_2
X_78136_ _78120_/C _78132_/Y _78135_/Y _78136_/X sky130_fd_sc_hd__o21a_4
X_44528_ _44528_/A _44529_/A sky130_fd_sc_hd__buf_2
X_63362_ _63357_/X _63363_/A sky130_fd_sc_hd__inv_2
X_75348_ _75348_/A _75348_/Y sky130_fd_sc_hd__inv_2
X_48296_ _66214_/B _48293_/X _48295_/Y _48296_/Y sky130_fd_sc_hd__o21ai_4
X_60574_ _60610_/A _60513_/B _79137_/A _60574_/X sky130_fd_sc_hd__or3_4
X_65101_ _65099_/X _83294_/Q _65028_/X _65100_/X _65102_/B sky130_fd_sc_hd__a211o_4
X_62313_ _62311_/Y _62253_/X _62312_/Y _84419_/D sky130_fd_sc_hd__a21oi_4
X_47247_ _81823_/Q _54630_/D sky130_fd_sc_hd__inv_2
X_66081_ _65615_/X _66195_/B _65617_/X _66081_/Y sky130_fd_sc_hd__nand3_4
X_78067_ _84572_/Q _78067_/B _78067_/X sky130_fd_sc_hd__xor2_4
X_44459_ _41133_/Y _44453_/X _87099_/Q _44454_/X _44459_/X sky130_fd_sc_hd__a2bb2o_4
X_63293_ _63287_/Y _63288_/X _63291_/X _63292_/X _63242_/X _63293_/Y
+ sky130_fd_sc_hd__o41ai_4
X_75279_ _75241_/Y _75279_/B _75279_/Y sky130_fd_sc_hd__nor2_4
X_65032_ _64929_/A _65032_/B _65032_/X sky130_fd_sc_hd__and2_4
X_77018_ _77018_/A _82277_/D _77021_/A sky130_fd_sc_hd__xnor2_4
X_62244_ _62194_/A _58225_/X _62244_/C _62244_/D _62244_/X sky130_fd_sc_hd__and4_4
X_47178_ _47130_/A _47181_/B sky130_fd_sc_hd__buf_2
X_46129_ _46129_/A _46164_/A sky130_fd_sc_hd__buf_2
X_69840_ _69836_/X _69839_/X _69768_/X _69840_/X sky130_fd_sc_hd__a21o_4
X_62175_ _62174_/X _62175_/B _61761_/C _62060_/X _62175_/Y sky130_fd_sc_hd__nand4_4
X_61126_ _61188_/B _61254_/B sky130_fd_sc_hd__buf_2
X_69771_ _44556_/A _69664_/X _69665_/X _69770_/X _69772_/B sky130_fd_sc_hd__a211o_4
Xclkbuf_7_60_0_CLK clkbuf_7_61_0_CLK/A clkbuf_7_60_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_66983_ _87938_/Q _66935_/X _66911_/X _66982_/X _66983_/X sky130_fd_sc_hd__a211o_4
X_78969_ _78969_/A _78979_/A sky130_fd_sc_hd__inv_2
X_68722_ _69956_/A _68938_/A sky130_fd_sc_hd__buf_2
X_65934_ _65158_/A _65934_/X sky130_fd_sc_hd__buf_2
X_61057_ _61055_/A _59771_/X _61057_/C _61057_/X sky130_fd_sc_hd__or3_4
X_81980_ _83905_/CLK _81980_/D _77814_/B sky130_fd_sc_hd__dfxtp_4
X_60008_ _59977_/A _60079_/B sky130_fd_sc_hd__buf_2
X_49819_ _49814_/Y _49815_/X _49818_/X _86318_/D sky130_fd_sc_hd__a21oi_4
X_68653_ _88008_/Q _68650_/X _68651_/X _68652_/X _68653_/X sky130_fd_sc_hd__a211o_4
X_80931_ _80931_/CLK _75082_/B _80931_/Q sky130_fd_sc_hd__dfxtp_4
X_65865_ _65768_/A _65865_/X sky130_fd_sc_hd__buf_2
X_67604_ _87912_/Q _67533_/X _67508_/X _67603_/X _67604_/X sky130_fd_sc_hd__a211o_4
X_52830_ _85747_/Q _52821_/X _52829_/Y _52830_/Y sky130_fd_sc_hd__o21ai_4
X_64816_ _64813_/Y _64814_/X _64815_/X _84226_/D sky130_fd_sc_hd__a21o_4
Xclkbuf_7_75_0_CLK clkbuf_7_74_0_CLK/A clkbuf_7_75_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_83650_ _85529_/CLK _70958_/Y _83650_/Q sky130_fd_sc_hd__dfxtp_4
X_80862_ _80961_/CLK _80894_/Q _75046_/B sky130_fd_sc_hd__dfxtp_4
X_68584_ _68516_/X _68574_/Y _68447_/X _68583_/Y _68584_/X sky130_fd_sc_hd__a211o_4
X_65796_ _65793_/X _65795_/X _65566_/X _65796_/X sky130_fd_sc_hd__a21o_4
X_82601_ _82924_/CLK _78869_/B _82569_/D sky130_fd_sc_hd__dfxtp_4
X_67535_ _87915_/Q _67533_/X _67508_/X _67534_/X _67535_/X sky130_fd_sc_hd__a211o_4
X_52761_ _85759_/Q _52737_/X _52760_/Y _52761_/Y sky130_fd_sc_hd__o21ai_4
X_64747_ _64744_/X _64746_/X _64629_/X _64747_/X sky130_fd_sc_hd__a21o_4
X_83581_ _83068_/CLK _71179_/Y _83581_/Q sky130_fd_sc_hd__dfxtp_4
X_61959_ _61645_/A _61959_/X sky130_fd_sc_hd__buf_2
X_80793_ _80968_/CLK _75789_/Y _80793_/Q sky130_fd_sc_hd__dfxtp_4
X_54500_ _54486_/X _47023_/Y _54500_/Y sky130_fd_sc_hd__nand2_4
X_85320_ _85351_/CLK _85320_/D _85320_/Q sky130_fd_sc_hd__dfxtp_4
X_51712_ _51717_/A _53236_/B _51712_/Y sky130_fd_sc_hd__nand2_4
X_82532_ _82532_/CLK _83852_/Q _82532_/Q sky130_fd_sc_hd__dfxtp_4
X_55480_ _85074_/Q _55481_/B sky130_fd_sc_hd__inv_2
X_67466_ _69751_/A _67466_/X sky130_fd_sc_hd__buf_2
X_52692_ _52706_/A _52692_/B _52692_/Y sky130_fd_sc_hd__nand2_4
X_64678_ _64678_/A _64678_/X sky130_fd_sc_hd__buf_2
X_69205_ _68384_/A _69205_/X sky130_fd_sc_hd__buf_2
X_54431_ _54376_/A _54431_/X sky130_fd_sc_hd__buf_2
X_66417_ _64876_/X _66417_/B _64879_/X _66417_/Y sky130_fd_sc_hd__nand3_4
X_85251_ _85186_/CLK _56271_/Y _56270_/C sky130_fd_sc_hd__dfxtp_4
X_51643_ _51627_/A _53167_/B _51643_/Y sky130_fd_sc_hd__nand2_4
X_63629_ _63657_/A _63629_/B _63629_/X sky130_fd_sc_hd__and2_4
X_82463_ _82463_/CLK _79155_/X _82463_/Q sky130_fd_sc_hd__dfxtp_4
X_67397_ _67393_/X _67396_/X _67322_/X _67397_/X sky130_fd_sc_hd__a21o_4
X_84202_ _85315_/CLK _84202_/D _65421_/C sky130_fd_sc_hd__dfxtp_4
X_57150_ _57149_/X _57141_/X _58981_/A _57150_/Y sky130_fd_sc_hd__a21oi_4
X_81414_ _82053_/CLK _81446_/Q _75952_/B sky130_fd_sc_hd__dfxtp_4
X_69136_ _69236_/A _87283_/Q _69136_/X sky130_fd_sc_hd__and2_4
X_54362_ _54362_/A _54362_/B _54362_/C _54362_/D _54362_/X sky130_fd_sc_hd__and4_4
X_66348_ _66266_/X _86210_/Q _66295_/X _66347_/X _66348_/X sky130_fd_sc_hd__a211o_4
X_85182_ _85248_/CLK _56476_/Y _55960_/B sky130_fd_sc_hd__dfxtp_4
X_51574_ _51629_/A _51580_/A sky130_fd_sc_hd__buf_2
X_82394_ _82394_/CLK _82202_/Q _82394_/Q sky130_fd_sc_hd__dfxtp_4
X_56101_ _56082_/X _56099_/X _56100_/Y _85296_/D sky130_fd_sc_hd__o21ai_4
X_53313_ _53310_/Y _53301_/X _53312_/X _85657_/D sky130_fd_sc_hd__a21oi_4
X_84133_ _82748_/CLK _84133_/D _84133_/Q sky130_fd_sc_hd__dfxtp_4
X_50525_ _50551_/A _50525_/X sky130_fd_sc_hd__buf_2
X_57081_ _56910_/X _56915_/Y _56982_/X _57081_/Y sky130_fd_sc_hd__a21oi_4
X_81345_ _83940_/CLK _76645_/Y _81721_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_13_0_CLK clkbuf_6_6_0_CLK/X clkbuf_8_27_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_69067_ _69067_/A _74226_/A _69067_/X sky130_fd_sc_hd__and2_4
X_54293_ _54289_/Y _54285_/X _54292_/X _54293_/Y sky130_fd_sc_hd__a21oi_4
X_66279_ _66003_/A _66319_/B sky130_fd_sc_hd__buf_2
Xclkbuf_8_153_0_CLK clkbuf_7_76_0_CLK/X clkbuf_9_307_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_68018_ _67972_/A _68018_/B _68018_/X sky130_fd_sc_hd__and2_4
X_56032_ _56023_/A _56017_/B _55943_/B _56032_/Y sky130_fd_sc_hd__nand3_4
X_53244_ _53243_/X _53244_/B _53222_/X _53244_/D _53244_/X sky130_fd_sc_hd__and4_4
X_84064_ _84064_/CLK _67567_/X _84064_/Q sky130_fd_sc_hd__dfxtp_4
X_50456_ _52161_/A _50456_/B _50462_/C _50456_/X sky130_fd_sc_hd__and3_4
X_81276_ _81627_/CLK _81276_/D _81276_/Q sky130_fd_sc_hd__dfxtp_4
X_83015_ _83013_/CLK _83015_/D _83015_/Q sky130_fd_sc_hd__dfxtp_4
X_80227_ _80189_/A _80221_/X _80226_/Y _80227_/Y sky130_fd_sc_hd__a21oi_4
X_53175_ _85683_/Q _53172_/X _53174_/Y _53175_/Y sky130_fd_sc_hd__o21ai_4
X_50387_ _50594_/A _50387_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_28_0_CLK clkbuf_7_28_0_CLK/A clkbuf_8_57_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_52126_ _52126_/A _52215_/A sky130_fd_sc_hd__buf_2
X_87823_ _87288_/CLK _42553_/Y _87823_/Q sky130_fd_sc_hd__dfxtp_4
X_80158_ _80142_/X _80145_/Y _80158_/X sky130_fd_sc_hd__or2_4
X_57983_ _58858_/A _57983_/X sky130_fd_sc_hd__buf_2
X_69969_ _68360_/X _69969_/B _69969_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_8_168_0_CLK clkbuf_7_84_0_CLK/X clkbuf_8_168_0_CLK/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_163_0_CLK clkbuf_9_81_0_CLK/X _81257_/CLK sky130_fd_sc_hd__clkbuf_1
X_59722_ _59722_/A _59722_/X sky130_fd_sc_hd__buf_2
X_56934_ _56933_/X _56934_/X sky130_fd_sc_hd__buf_2
X_52057_ _74127_/B _52041_/X _52056_/Y _52057_/Y sky130_fd_sc_hd__o21ai_4
X_87754_ _87757_/CLK _42715_/X _87754_/Q sky130_fd_sc_hd__dfxtp_4
X_72980_ _87307_/Q _72744_/X _72980_/Y sky130_fd_sc_hd__nor2_4
X_84966_ _86534_/CLK _84966_/D _84966_/Q sky130_fd_sc_hd__dfxtp_4
X_80089_ _57944_/Y _65683_/C _80088_/Y _80089_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_10_793_0_CLK clkbuf_9_396_0_CLK/X _82715_/CLK sky130_fd_sc_hd__clkbuf_1
X_51008_ _51003_/A _51008_/B _51008_/Y sky130_fd_sc_hd__nand2_4
X_86705_ _86384_/CLK _86705_/D _58776_/A sky130_fd_sc_hd__dfxtp_4
X_71931_ _71920_/Y _57170_/A _71930_/Y _71931_/X sky130_fd_sc_hd__a21o_4
X_59653_ _59961_/A _66064_/A sky130_fd_sc_hd__buf_2
X_83917_ _83918_/CLK _83917_/D _81381_/D sky130_fd_sc_hd__dfxtp_4
X_56865_ _58517_/A _55282_/B _56864_/X _56865_/Y sky130_fd_sc_hd__o21ai_4
X_87685_ _88128_/CLK _87685_/D _66900_/B sky130_fd_sc_hd__dfxtp_4
X_84897_ _84897_/CLK _58252_/X _61985_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_284_0_CLK clkbuf_9_285_0_CLK/A clkbuf_9_284_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_58604_ _58585_/X _58600_/Y _58601_/Y _58603_/X _58589_/X _58604_/X
+ sky130_fd_sc_hd__o32a_4
X_55816_ _55813_/X _55815_/X _55309_/X _55816_/X sky130_fd_sc_hd__a21o_4
X_43830_ _43830_/A _43830_/Y sky130_fd_sc_hd__inv_2
X_74650_ _74642_/X _45560_/A _74650_/Y sky130_fd_sc_hd__nand2_4
X_86636_ _86637_/CLK _86636_/D _86636_/Q sky130_fd_sc_hd__dfxtp_4
X_71862_ _71848_/X _83349_/Q _71861_/Y _83349_/D sky130_fd_sc_hd__a21o_4
X_83848_ _83843_/CLK _83848_/D _83848_/Q sky130_fd_sc_hd__dfxtp_4
X_59584_ _57686_/A _44003_/A _59584_/C _59585_/A sky130_fd_sc_hd__nor3_4
X_56796_ _72765_/A _56796_/B _56796_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_178_0_CLK clkbuf_9_89_0_CLK/X _81603_/CLK sky130_fd_sc_hd__clkbuf_1
X_73601_ _73596_/X _73600_/X _56549_/X _73601_/X sky130_fd_sc_hd__a21o_4
X_70813_ _52889_/B _70802_/X _70812_/Y _83695_/D sky130_fd_sc_hd__o21ai_4
X_58535_ _58535_/A _58535_/Y sky130_fd_sc_hd__inv_2
X_43761_ _43005_/X _43760_/X _40959_/X _87279_/Q _43756_/X _43762_/A
+ sky130_fd_sc_hd__o32ai_4
X_55747_ _55174_/X _55747_/X sky130_fd_sc_hd__buf_2
X_74581_ _45124_/A _74568_/X _74580_/X _74581_/Y sky130_fd_sc_hd__o21ai_4
X_86567_ _86213_/CLK _48113_/Y _66285_/B sky130_fd_sc_hd__dfxtp_4
X_40973_ _40944_/X _40946_/X _40972_/X _88300_/Q _40916_/X _40973_/Y
+ sky130_fd_sc_hd__o32ai_4
X_52959_ _52979_/A _52959_/B _52959_/Y sky130_fd_sc_hd__nand2_4
X_71793_ _58196_/Y _71784_/X _71792_/Y _71793_/Y sky130_fd_sc_hd__o21ai_4
X_83779_ _85953_/CLK _70403_/Y _83779_/Q sky130_fd_sc_hd__dfxtp_4
X_45500_ _45500_/A _45500_/Y sky130_fd_sc_hd__inv_2
X_76320_ _76299_/Y _76320_/Y sky130_fd_sc_hd__inv_2
X_42712_ _41147_/X _42710_/X _68528_/B _42711_/X _87757_/D sky130_fd_sc_hd__a2bb2o_4
X_88306_ _86989_/CLK _88306_/D _88306_/Q sky130_fd_sc_hd__dfxtp_4
X_73532_ _73528_/X _73531_/X _56549_/X _73532_/X sky130_fd_sc_hd__a21o_4
X_85518_ _86030_/CLK _54040_/Y _85518_/Q sky130_fd_sc_hd__dfxtp_4
X_70744_ _70755_/A _70753_/A sky130_fd_sc_hd__buf_2
X_46480_ _82925_/Q _48044_/B sky130_fd_sc_hd__inv_2
X_58466_ _58341_/X _58463_/Y _58465_/Y _58466_/Y sky130_fd_sc_hd__a21oi_4
X_43692_ _87305_/Q _69700_/B sky130_fd_sc_hd__inv_2
X_55678_ _55678_/A _55290_/A _55678_/X sky130_fd_sc_hd__and2_4
X_86498_ _86498_/CLK _48712_/Y _86498_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_299_0_CLK clkbuf_9_299_0_CLK/A clkbuf_9_299_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_8_106_0_CLK clkbuf_7_53_0_CLK/X clkbuf_8_106_0_CLK/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_101_0_CLK clkbuf_9_50_0_CLK/X _84538_/CLK sky130_fd_sc_hd__clkbuf_1
X_45431_ _83007_/Q _45401_/X _45430_/X _45431_/Y sky130_fd_sc_hd__o21ai_4
X_57417_ _57408_/X _57415_/X _57416_/Y _57417_/Y sky130_fd_sc_hd__o21ai_4
X_88237_ _88164_/CLK _88237_/D _88237_/Q sky130_fd_sc_hd__dfxtp_4
X_76251_ _76250_/Y _81641_/Q _76251_/C _76254_/B sky130_fd_sc_hd__nand3_4
X_42643_ _40964_/X _42631_/X _69203_/B _42634_/X _87790_/D sky130_fd_sc_hd__a2bb2o_4
X_54629_ _54521_/A _54645_/B sky130_fd_sc_hd__buf_2
X_85449_ _85770_/CLK _54403_/Y _85449_/Q sky130_fd_sc_hd__dfxtp_4
X_73463_ _69929_/Y _73224_/X _73393_/X _73462_/Y _73463_/X sky130_fd_sc_hd__a211o_4
X_70675_ _71857_/A _70676_/A sky130_fd_sc_hd__buf_2
X_58397_ _58396_/Y _58403_/B _58397_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_731_0_CLK clkbuf_9_365_0_CLK/X _87253_/CLK sky130_fd_sc_hd__clkbuf_1
X_75202_ _80682_/Q _80938_/D _75202_/Y sky130_fd_sc_hd__nand2_4
X_48150_ _48781_/A _48150_/X sky130_fd_sc_hd__buf_2
X_72414_ _59255_/A _72414_/X sky130_fd_sc_hd__buf_2
X_45362_ _45356_/Y _45359_/Y _45361_/X _45362_/X sky130_fd_sc_hd__a21o_4
X_57348_ _57346_/Y _56857_/X _46155_/A _57347_/Y _57348_/X sky130_fd_sc_hd__a211o_4
X_76182_ _76179_/Y _76182_/B _76182_/Y sky130_fd_sc_hd__nor2_4
X_88168_ _86934_/CLK _41694_/X _67608_/B sky130_fd_sc_hd__dfxtp_4
X_42574_ _42574_/A _42574_/X sky130_fd_sc_hd__buf_2
X_73394_ _73394_/A _73053_/B _73394_/Y sky130_fd_sc_hd__nor2_4
X_47101_ _59240_/A _47096_/X _47100_/Y _47101_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_222_0_CLK clkbuf_9_222_0_CLK/A clkbuf_9_222_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_44313_ _44313_/A _44313_/B _46228_/A _44313_/Y sky130_fd_sc_hd__nand3_4
X_75133_ _75130_/Y _75133_/B _75133_/Y sky130_fd_sc_hd__nor2_4
X_87119_ _87684_/CLK _87119_/D _87119_/Q sky130_fd_sc_hd__dfxtp_4
X_41525_ _41524_/Y _41525_/X sky130_fd_sc_hd__buf_2
X_72345_ _72341_/Y _72343_/Y _72344_/X _72345_/X sky130_fd_sc_hd__a21o_4
X_48081_ _83537_/Q _48081_/Y sky130_fd_sc_hd__inv_2
X_45293_ _64494_/B _61627_/B sky130_fd_sc_hd__buf_2
X_57279_ _56696_/A _44277_/X _57278_/Y _85041_/D sky130_fd_sc_hd__a21oi_4
X_88099_ _88104_/CLK _88099_/D _41941_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_116_0_CLK clkbuf_9_58_0_CLK/X _84905_/CLK sky130_fd_sc_hd__clkbuf_1
X_47032_ _53332_/B _52813_/B sky130_fd_sc_hd__buf_2
X_59018_ _58920_/A _86367_/Q _59018_/Y sky130_fd_sc_hd__nor2_4
X_44244_ _44244_/A _44245_/A sky130_fd_sc_hd__buf_2
X_75064_ _75062_/Y _75059_/B _75063_/Y _75067_/A sky130_fd_sc_hd__o21ai_4
X_79941_ _84925_/Q _65855_/C _79941_/Y sky130_fd_sc_hd__nand2_4
X_41456_ _40565_/Y _41457_/A sky130_fd_sc_hd__buf_2
X_60290_ _60259_/B _60350_/A _61286_/A _60290_/Y sky130_fd_sc_hd__a21oi_4
X_72276_ _72263_/Y _72237_/X _72269_/X _72275_/X _83269_/D sky130_fd_sc_hd__a22oi_4
Xclkbuf_10_746_0_CLK clkbuf_9_373_0_CLK/X _87484_/CLK sky130_fd_sc_hd__clkbuf_1
X_74015_ _74012_/X _86222_/Q _73948_/X _74014_/X _74015_/X sky130_fd_sc_hd__a211o_4
X_40407_ _40381_/X _81177_/Q _40406_/X _40407_/Y sky130_fd_sc_hd__o21ai_4
X_71227_ _48851_/B _71216_/X _71226_/Y _71227_/Y sky130_fd_sc_hd__o21ai_4
X_44175_ _44175_/A _64679_/A sky130_fd_sc_hd__buf_2
X_79872_ _79872_/A _79872_/B _79873_/B sky130_fd_sc_hd__xor2_4
X_41387_ _41387_/A _41387_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_237_0_CLK clkbuf_8_118_0_CLK/X clkbuf_9_237_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_43126_ _43126_/A _43126_/Y sky130_fd_sc_hd__inv_2
X_78823_ _79123_/B _78825_/A sky130_fd_sc_hd__inv_2
X_40338_ _40337_/X _46259_/A sky130_fd_sc_hd__buf_2
X_71158_ _52128_/B _71138_/A _71157_/Y _83587_/D sky130_fd_sc_hd__o21ai_4
X_48983_ _48964_/A _48982_/X _48983_/Y sky130_fd_sc_hd__nand2_4
X_70109_ _83126_/Q _70109_/Y sky130_fd_sc_hd__inv_2
X_47934_ _47857_/X _47946_/A sky130_fd_sc_hd__buf_2
X_43057_ _43057_/A _43057_/Y sky130_fd_sc_hd__inv_2
X_78754_ _78753_/B _78753_/C _78749_/Y _78758_/C sky130_fd_sc_hd__o21ai_4
X_63980_ _58533_/A _63934_/X _63949_/C _64027_/D _63980_/Y sky130_fd_sc_hd__nand4_4
X_71089_ _49025_/X _71070_/A _71088_/Y _71089_/Y sky130_fd_sc_hd__o21ai_4
X_75966_ _81512_/Q _81736_/D _75966_/X sky130_fd_sc_hd__xor2_4
X_42008_ _41960_/X _42006_/X _40814_/X _73033_/A _42007_/X _42009_/A
+ sky130_fd_sc_hd__o32ai_4
X_77705_ _77704_/Y _77702_/A _77710_/A sky130_fd_sc_hd__nand2_4
X_62931_ _62929_/Y _62893_/X _62930_/Y _84369_/D sky130_fd_sc_hd__a21oi_4
X_74917_ _74908_/Y _74915_/Y _74916_/Y _74917_/X sky130_fd_sc_hd__o21a_4
X_47865_ _47855_/A _51947_/B _47865_/Y sky130_fd_sc_hd__nand2_4
X_78685_ _78685_/A _78684_/X _78701_/A sky130_fd_sc_hd__xnor2_4
X_75897_ _61262_/C _84367_/Q _75897_/X sky130_fd_sc_hd__xor2_4
X_49604_ _49601_/Y _49596_/X _49603_/X _49604_/Y sky130_fd_sc_hd__a21oi_4
X_46816_ _52692_/B _50998_/B sky130_fd_sc_hd__buf_2
X_65650_ _84187_/Q _65651_/C sky130_fd_sc_hd__inv_2
X_77636_ _77635_/X _77636_/Y sky130_fd_sc_hd__inv_2
X_62862_ _62847_/X _63209_/A _62911_/C _62880_/D _62862_/X sky130_fd_sc_hd__and4_4
X_74848_ _81122_/D _74848_/B _74849_/B sky130_fd_sc_hd__xor2_4
X_47796_ _47790_/Y _47791_/X _47795_/X _47796_/Y sky130_fd_sc_hd__a21oi_4
X_64601_ _64601_/A _64602_/A sky130_fd_sc_hd__buf_2
X_49535_ _49546_/A _52748_/B _49535_/Y sky130_fd_sc_hd__nand2_4
X_61813_ _61811_/X _61765_/B _61846_/C _61846_/D _61813_/Y sky130_fd_sc_hd__nand4_4
X_46747_ _83675_/Q _52651_/B sky130_fd_sc_hd__inv_2
X_65581_ _65503_/X _85591_/Q _65504_/X _65580_/X _65581_/X sky130_fd_sc_hd__a211o_4
X_77567_ _77568_/A _82105_/D _77567_/Y sky130_fd_sc_hd__nor2_4
X_43959_ _43959_/A _43959_/B _59538_/D sky130_fd_sc_hd__and2_4
X_62793_ _62672_/A _62839_/B sky130_fd_sc_hd__buf_2
X_74779_ _70180_/Y _70692_/C _83830_/Q _74716_/X _74779_/X sky130_fd_sc_hd__a2bb2o_4
X_67320_ _67320_/A _86775_/Q _67320_/X sky130_fd_sc_hd__and2_4
X_79306_ _79303_/X _79306_/B _82829_/D sky130_fd_sc_hd__xor2_4
X_64532_ _72381_/A _64532_/X sky130_fd_sc_hd__buf_2
X_76518_ _76518_/A _76518_/B _76518_/X sky130_fd_sc_hd__xor2_4
X_61744_ _84728_/Q _61744_/X sky130_fd_sc_hd__buf_2
X_49466_ _49493_/A _49467_/C sky130_fd_sc_hd__buf_2
X_46678_ _58649_/A _46672_/X _46677_/Y _46678_/Y sky130_fd_sc_hd__o21ai_4
X_77498_ _77458_/X _77480_/Y _77478_/X _77498_/X sky130_fd_sc_hd__and3_4
X_48417_ _48557_/A _52123_/B _48417_/Y sky130_fd_sc_hd__nand2_4
X_67251_ _87415_/Q _67156_/X _67226_/X _67250_/X _67251_/X sky130_fd_sc_hd__a211o_4
X_79237_ _79213_/Y _79215_/X _79236_/Y _79239_/A sky130_fd_sc_hd__a21oi_4
X_45629_ _85074_/Q _45801_/A _45629_/Y sky130_fd_sc_hd__nor2_4
X_64463_ _64461_/Y _64186_/X _64462_/Y _64463_/Y sky130_fd_sc_hd__a21oi_4
X_76449_ _81366_/Q _76449_/B _76449_/X sky130_fd_sc_hd__xor2_4
X_49397_ _49397_/A _49420_/B _49408_/C _50919_/D _49397_/X sky130_fd_sc_hd__and4_4
X_61675_ _61292_/A _61675_/B _61675_/C _61675_/Y sky130_fd_sc_hd__nand3_4
X_66202_ _57761_/X _84973_/Q _65950_/X _66201_/X _66203_/C sky130_fd_sc_hd__a211o_4
X_63414_ _63400_/A _58232_/A _63463_/C _63414_/X sky130_fd_sc_hd__and3_4
X_48348_ _48348_/A _50385_/B _48348_/Y sky130_fd_sc_hd__nand2_4
X_60626_ _60626_/A _60628_/A sky130_fd_sc_hd__inv_2
X_67182_ _67062_/X _67183_/A sky130_fd_sc_hd__buf_2
X_79168_ _79168_/A _79169_/A sky130_fd_sc_hd__inv_2
X_64394_ _64380_/X _84818_/Q _64381_/X _64394_/Y sky130_fd_sc_hd__nand3_4
X_66133_ _66040_/X _84978_/Q _66027_/X _66132_/X _66133_/X sky130_fd_sc_hd__a211o_4
X_78119_ _78120_/A _78120_/C _78120_/B _78119_/X sky130_fd_sc_hd__a21o_4
X_63345_ _63343_/Y _63344_/X _63317_/X _63345_/X sky130_fd_sc_hd__a21o_4
X_48279_ _48244_/A _48024_/B _48279_/Y sky130_fd_sc_hd__nand2_4
X_60557_ _60556_/Y _60557_/Y sky130_fd_sc_hd__inv_2
X_79099_ _79099_/A _79099_/Y sky130_fd_sc_hd__inv_2
X_50310_ _50240_/A _50310_/B _50310_/Y sky130_fd_sc_hd__nand2_4
X_81130_ _81130_/CLK _81130_/D _40714_/A sky130_fd_sc_hd__dfxtp_4
X_66064_ _66064_/A _66065_/A sky130_fd_sc_hd__buf_2
X_51290_ _51298_/A _51290_/B _51290_/X sky130_fd_sc_hd__and2_4
X_63276_ _63285_/A _63285_/B _79267_/A _63276_/Y sky130_fd_sc_hd__nor3_4
X_60488_ _60488_/A _60488_/B _60488_/C _60488_/Y sky130_fd_sc_hd__nand3_4
X_65015_ _64600_/A _65015_/X sky130_fd_sc_hd__buf_2
X_50241_ _86238_/Q _50238_/X _50240_/Y _50241_/Y sky130_fd_sc_hd__o21ai_4
X_62227_ _62620_/A _62632_/A sky130_fd_sc_hd__buf_2
X_81061_ _81061_/CLK _81093_/Q _81061_/Q sky130_fd_sc_hd__dfxtp_4
X_80012_ _79988_/A _80011_/D _80011_/B _80012_/X sky130_fd_sc_hd__a21bo_4
X_69823_ _69908_/A _69823_/B _69823_/Y sky130_fd_sc_hd__nor2_4
X_50172_ _50170_/Y _50166_/X _50171_/X _86250_/D sky130_fd_sc_hd__a21oi_4
X_62158_ _59730_/A _62170_/B _62158_/C _63333_/B _62158_/X sky130_fd_sc_hd__and4_4
X_61109_ _61108_/Y _61109_/X sky130_fd_sc_hd__buf_2
X_84820_ _83451_/CLK _58555_/X _84820_/Q sky130_fd_sc_hd__dfxtp_4
X_69754_ _69750_/X _69753_/X _68697_/X _69758_/A sky130_fd_sc_hd__a21o_4
X_54980_ _54977_/Y _54971_/X _54979_/X _54980_/Y sky130_fd_sc_hd__a21oi_4
X_66966_ _66942_/A _66966_/B _66966_/X sky130_fd_sc_hd__and2_4
X_62089_ _62082_/X _62084_/X _62088_/Y _58465_/A _62048_/X _62089_/Y
+ sky130_fd_sc_hd__o32ai_4
X_68705_ _87494_/Q _68626_/X _68601_/X _68704_/X _68705_/X sky130_fd_sc_hd__a211o_4
X_53931_ _53928_/Y _53914_/X _53930_/Y _53931_/Y sky130_fd_sc_hd__a21boi_4
X_65917_ _65914_/Y _65915_/X _65916_/X _84169_/D sky130_fd_sc_hd__a21o_4
X_84751_ _84757_/CLK _59324_/Y _84751_/Q sky130_fd_sc_hd__dfxtp_4
X_81963_ _82299_/CLK _81963_/D _81963_/Q sky130_fd_sc_hd__dfxtp_4
X_69685_ _69685_/A _87306_/Q _69685_/X sky130_fd_sc_hd__and2_4
X_66897_ _69654_/A _69156_/A sky130_fd_sc_hd__buf_2
X_83702_ _83703_/CLK _83702_/D _83702_/Q sky130_fd_sc_hd__dfxtp_4
X_56650_ _56649_/X _56650_/B _56650_/Y sky130_fd_sc_hd__nor2_4
X_80914_ _81507_/CLK _80914_/D _80914_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_10_0_CLK clkbuf_3_5_1_CLK/X clkbuf_4_10_1_CLK/A sky130_fd_sc_hd__clkbuf_1
X_68636_ _69747_/A _68636_/X sky130_fd_sc_hd__buf_2
X_87470_ _86934_/CLK _87470_/D _87470_/Q sky130_fd_sc_hd__dfxtp_4
X_53862_ _53838_/A _53862_/X sky130_fd_sc_hd__buf_2
X_65848_ _65807_/A _86469_/Q _65848_/X sky130_fd_sc_hd__and2_4
X_84682_ _84713_/CLK _59874_/Y _80266_/B sky130_fd_sc_hd__dfxtp_4
X_81894_ _82139_/CLK _77291_/X _82302_/D sky130_fd_sc_hd__dfxtp_4
X_55601_ _55601_/A _55601_/B _55601_/X sky130_fd_sc_hd__and2_4
X_86421_ _86422_/CLK _49268_/Y _86421_/Q sky130_fd_sc_hd__dfxtp_4
X_52813_ _52803_/A _52813_/B _52813_/Y sky130_fd_sc_hd__nand2_4
X_83633_ _83275_/CLK _83633_/D _47597_/A sky130_fd_sc_hd__dfxtp_4
X_56581_ _56618_/B _56582_/A sky130_fd_sc_hd__inv_2
X_80845_ _80754_/CLK _80877_/Q _74921_/B sky130_fd_sc_hd__dfxtp_4
X_68567_ _66053_/A _68567_/B _68567_/Y sky130_fd_sc_hd__nor2_4
X_53793_ _53793_/A _53825_/A sky130_fd_sc_hd__buf_2
X_65779_ _65779_/A _86474_/Q _65779_/X sky130_fd_sc_hd__and2_4
X_58320_ _58320_/A _58326_/B _58320_/Y sky130_fd_sc_hd__nand2_4
X_55532_ _44097_/X _55532_/X sky130_fd_sc_hd__buf_2
X_67518_ _86968_/Q _67467_/X _67516_/X _67517_/X _67518_/X sky130_fd_sc_hd__a211o_4
X_86352_ _86353_/CLK _86352_/D _86352_/Q sky130_fd_sc_hd__dfxtp_4
X_52744_ _52744_/A _52744_/B _52744_/Y sky130_fd_sc_hd__nand2_4
X_83564_ _83564_/CLK _71231_/Y _48682_/A sky130_fd_sc_hd__dfxtp_4
X_80776_ _80776_/CLK _80776_/D _80776_/Q sky130_fd_sc_hd__dfxtp_4
X_68498_ _69877_/A _68498_/B _68498_/X sky130_fd_sc_hd__and2_4
X_85303_ _85269_/CLK _85303_/D _55900_/B sky130_fd_sc_hd__dfxtp_4
X_58251_ _58251_/A _58217_/B _58251_/Y sky130_fd_sc_hd__nand2_4
X_82515_ _82515_/CLK _82515_/D _82515_/Q sky130_fd_sc_hd__dfxtp_4
X_55463_ _55323_/A _55826_/A sky130_fd_sc_hd__buf_2
X_67449_ _67806_/A _67449_/X sky130_fd_sc_hd__buf_2
X_86283_ _85962_/CLK _86283_/D _86283_/Q sky130_fd_sc_hd__dfxtp_4
X_52675_ _52674_/X _52661_/B _52654_/C _46791_/X _52675_/X sky130_fd_sc_hd__and4_4
X_83495_ _83495_/CLK _83495_/D _83495_/Q sky130_fd_sc_hd__dfxtp_4
X_57202_ _57087_/X _57200_/Y _57201_/Y _57203_/A sky130_fd_sc_hd__o21ai_4
X_88022_ _87253_/CLK _88022_/D _88022_/Q sky130_fd_sc_hd__dfxtp_4
X_54414_ _54411_/Y _54394_/X _54413_/X _85447_/D sky130_fd_sc_hd__a21oi_4
X_85234_ _85167_/CLK _56329_/Y _55846_/B sky130_fd_sc_hd__dfxtp_4
X_51626_ _51624_/Y _51613_/X _51625_/X _51626_/Y sky130_fd_sc_hd__a21oi_4
X_70460_ _71337_/A _71323_/A sky130_fd_sc_hd__buf_2
X_58182_ _84913_/Q _58184_/A sky130_fd_sc_hd__buf_2
X_82446_ _82452_/CLK _79138_/X _82446_/Q sky130_fd_sc_hd__dfxtp_4
X_55394_ _55370_/X _55394_/B _55394_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_1003_0_CLK clkbuf_9_501_0_CLK/X _86490_/CLK sky130_fd_sc_hd__clkbuf_1
X_57133_ _57133_/A _56739_/A _57155_/D _56803_/A _57133_/X sky130_fd_sc_hd__and4_4
X_69119_ _86976_/Q _68864_/X _68891_/X _69118_/X _69119_/X sky130_fd_sc_hd__a211o_4
X_54345_ _54399_/A _54362_/A sky130_fd_sc_hd__buf_2
X_85165_ _85257_/CLK _85165_/D _56518_/C sky130_fd_sc_hd__dfxtp_4
X_51557_ _51557_/A _51557_/X sky130_fd_sc_hd__buf_2
X_70391_ _71003_/A _70944_/A sky130_fd_sc_hd__buf_2
X_82377_ _85635_/CLK _82185_/Q _82377_/Q sky130_fd_sc_hd__dfxtp_4
X_41310_ _41310_/A _41292_/B _41310_/X sky130_fd_sc_hd__or2_4
X_72130_ _59325_/X _72128_/Y _72129_/Y _59342_/X _59329_/X _72130_/X
+ sky130_fd_sc_hd__o32a_4
X_84116_ _84161_/CLK _84116_/D _84116_/Q sky130_fd_sc_hd__dfxtp_4
X_50508_ _50513_/A _50508_/B _50508_/Y sky130_fd_sc_hd__nand2_4
X_57064_ _56885_/A _56884_/Y _56982_/X _57064_/Y sky130_fd_sc_hd__a21oi_4
X_81328_ _81492_/CLK _76363_/X _81704_/D sky130_fd_sc_hd__dfxtp_4
X_54276_ _54273_/Y _54051_/X _54275_/X _85472_/D sky130_fd_sc_hd__a21oi_4
X_42290_ _42290_/A _42290_/X sky130_fd_sc_hd__buf_2
X_85096_ _85096_/CLK _85096_/D _85096_/Q sky130_fd_sc_hd__dfxtp_4
X_51488_ _86001_/Q _51485_/X _51487_/Y _51488_/Y sky130_fd_sc_hd__o21ai_4
X_56015_ _55975_/X _56015_/B _56016_/A sky130_fd_sc_hd__xor2_4
X_53227_ _53246_/A _53227_/B _53227_/Y sky130_fd_sc_hd__nand2_4
X_41241_ _41490_/A _41241_/X sky130_fd_sc_hd__buf_2
X_72061_ _72058_/Y _72059_/X _72060_/X _83293_/D sky130_fd_sc_hd__a21oi_4
X_84047_ _88116_/CLK _84047_/D _81479_/D sky130_fd_sc_hd__dfxtp_4
X_50439_ _50534_/A _50439_/X sky130_fd_sc_hd__buf_2
X_81259_ _81259_/CLK _81259_/D _81259_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_1018_0_CLK clkbuf_9_509_0_CLK/X _86506_/CLK sky130_fd_sc_hd__clkbuf_1
X_71012_ _71012_/A _71012_/B _71013_/A sky130_fd_sc_hd__nor2_4
X_41172_ _41002_/B _41223_/B _41172_/X sky130_fd_sc_hd__or2_4
X_53158_ _85686_/Q _53146_/X _53157_/Y _53158_/Y sky130_fd_sc_hd__o21ai_4
X_52109_ _48388_/A _52135_/B _52097_/X _52109_/X sky130_fd_sc_hd__and3_4
X_75820_ _75820_/A _75821_/B sky130_fd_sc_hd__inv_2
X_87806_ _87820_/CLK _42601_/Y _42600_/A sky130_fd_sc_hd__dfxtp_4
X_57966_ _58813_/A _57966_/X sky130_fd_sc_hd__buf_2
X_45980_ _45980_/A _45980_/X sky130_fd_sc_hd__buf_2
X_53089_ _53195_/A _53107_/C sky130_fd_sc_hd__buf_2
X_85998_ _85709_/CLK _85998_/D _85998_/Q sky130_fd_sc_hd__dfxtp_4
X_59705_ _59564_/B _59705_/X sky130_fd_sc_hd__buf_2
X_44931_ _44928_/Y _44930_/Y _44889_/X _44931_/X sky130_fd_sc_hd__a21o_4
X_56917_ _56917_/A _56798_/B _56917_/Y sky130_fd_sc_hd__nand2_4
X_75751_ _75751_/A _75750_/Y _75759_/A sky130_fd_sc_hd__xor2_4
X_87737_ _87993_/CLK _42754_/X _69008_/B sky130_fd_sc_hd__dfxtp_4
X_72963_ _73359_/A _72963_/X sky130_fd_sc_hd__buf_2
X_84949_ _85485_/CLK _84949_/D _84949_/Q sky130_fd_sc_hd__dfxtp_4
X_57897_ _57971_/A _57897_/B _57897_/Y sky130_fd_sc_hd__nor2_4
X_74702_ _74691_/A _74702_/B _74702_/Y sky130_fd_sc_hd__nand2_4
X_47650_ _86612_/Q _47619_/X _47649_/Y _47650_/Y sky130_fd_sc_hd__o21ai_4
X_71914_ _71576_/X _71930_/B _71536_/A _71914_/Y sky130_fd_sc_hd__nor3_4
X_59636_ _59635_/Y _59806_/A sky130_fd_sc_hd__buf_2
X_78470_ _78461_/A _78458_/Y _78460_/A _78474_/A sky130_fd_sc_hd__o21a_4
X_44862_ _41781_/Y _44848_/X _68020_/B _44849_/X _44862_/X sky130_fd_sc_hd__a2bb2o_4
X_56848_ _56700_/C _56848_/X sky130_fd_sc_hd__buf_2
X_75682_ _75670_/A _75669_/Y _75656_/A _80780_/D _75682_/X sky130_fd_sc_hd__a2bb2o_4
X_87668_ _88180_/CLK _87668_/D _87668_/Q sky130_fd_sc_hd__dfxtp_4
X_72894_ _72806_/A _72894_/X sky130_fd_sc_hd__buf_2
X_46601_ _46493_/X _48157_/B _46600_/Y _54091_/A sky130_fd_sc_hd__o21ai_4
X_77421_ _77421_/A _82191_/D _81903_/D sky130_fd_sc_hd__xor2_4
X_43813_ _43813_/A _43813_/Y sky130_fd_sc_hd__inv_2
X_74633_ _74691_/A _74633_/X sky130_fd_sc_hd__buf_2
X_86619_ _85981_/CLK _86619_/D _72193_/A sky130_fd_sc_hd__dfxtp_4
X_47581_ _83707_/Q _47582_/A sky130_fd_sc_hd__inv_2
X_71845_ _70886_/A _71846_/A sky130_fd_sc_hd__buf_2
X_59567_ _59661_/D _60599_/A _60380_/B _59633_/A sky130_fd_sc_hd__and3_4
X_44793_ _44512_/A _41887_/A _41407_/X _86952_/Q _44516_/A _44794_/A
+ sky130_fd_sc_hd__o32ai_4
X_56779_ _56567_/Y _56778_/Y _56779_/Y sky130_fd_sc_hd__nor2_4
X_87599_ _88111_/CLK _87599_/D _73653_/A sky130_fd_sc_hd__dfxtp_4
X_49320_ _49287_/A _49320_/B _49320_/Y sky130_fd_sc_hd__nand2_4
X_46532_ _46522_/Y _46523_/X _46531_/Y _46532_/Y sky130_fd_sc_hd__a21boi_4
X_58518_ _83421_/Q _58518_/Y sky130_fd_sc_hd__inv_2
X_77352_ _81930_/Q _82186_/D _81898_/D sky130_fd_sc_hd__xor2_4
X_43744_ _43744_/A _69932_/B sky130_fd_sc_hd__inv_2
X_74564_ _74541_/A _46228_/A _74564_/C _74564_/Y sky130_fd_sc_hd__nand3_4
X_40956_ _40955_/X _40941_/X _88304_/Q _40942_/X _88304_/D sky130_fd_sc_hd__a2bb2o_4
X_71776_ _71761_/Y _83380_/Q _71775_/X _71776_/X sky130_fd_sc_hd__a21o_4
X_59498_ _59498_/A _59497_/Y _59498_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_670_0_CLK clkbuf_9_335_0_CLK/X _88133_/CLK sky130_fd_sc_hd__clkbuf_1
X_76303_ _76302_/Y _76303_/Y sky130_fd_sc_hd__inv_2
X_49251_ _49241_/A _46356_/X _49251_/Y sky130_fd_sc_hd__nand2_4
X_73515_ _72721_/X _86179_/Q _73351_/X _73514_/X _73515_/X sky130_fd_sc_hd__a211o_4
X_46463_ _46458_/Y _46399_/X _46462_/Y _86735_/D sky130_fd_sc_hd__a21boi_4
X_70727_ _70727_/A _70779_/B _70727_/C _70769_/D _70727_/Y sky130_fd_sc_hd__nand4_4
X_58449_ _84845_/Q _63244_/A sky130_fd_sc_hd__inv_2
X_77283_ _77282_/Y _77285_/A sky130_fd_sc_hd__inv_2
X_43675_ _87316_/Q _69114_/B sky130_fd_sc_hd__inv_2
X_74495_ _74490_/A _48660_/A _74495_/Y sky130_fd_sc_hd__nand2_4
X_40887_ _40887_/A _40887_/Y sky130_fd_sc_hd__inv_2
X_48202_ _48199_/Y _48194_/X _48201_/X _48202_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_161_0_CLK clkbuf_8_80_0_CLK/X clkbuf_9_161_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_79022_ _79022_/A _79018_/A _79022_/Y sky130_fd_sc_hd__nand2_4
X_45414_ _55628_/B _45412_/X _45396_/X _45413_/Y _45414_/X sky130_fd_sc_hd__a211o_4
X_76234_ _76234_/A _76234_/Y sky130_fd_sc_hd__inv_2
X_42626_ _42626_/A _40591_/B _40591_/C _42626_/X sky130_fd_sc_hd__and3_4
X_49182_ _49173_/A _50714_/B _49182_/X sky130_fd_sc_hd__and2_4
X_73446_ _72905_/A _73446_/X sky130_fd_sc_hd__buf_2
X_61460_ _61437_/A _61460_/B _61459_/X _61460_/Y sky130_fd_sc_hd__nand3_4
X_46394_ _83644_/Q _52484_/B sky130_fd_sc_hd__inv_2
X_70658_ _70727_/A _70656_/B _70890_/C _70656_/D _70658_/Y sky130_fd_sc_hd__nand4_4
X_48133_ _74234_/B _48103_/X _48132_/Y _48133_/Y sky130_fd_sc_hd__o21ai_4
XPHY_90 sky130_fd_sc_hd__decap_3
X_60411_ _63118_/A _63060_/A sky130_fd_sc_hd__buf_2
X_45345_ _45345_/A _45347_/A sky130_fd_sc_hd__inv_2
X_76165_ _76163_/Y _81634_/Q _76164_/Y _76165_/X sky130_fd_sc_hd__a21bo_4
X_42557_ _42554_/X _40792_/A _42477_/X _42555_/Y _42556_/X _87822_/D
+ sky130_fd_sc_hd__o32ai_4
X_61391_ _64272_/A _61368_/B _61368_/C _61391_/D _61392_/A sky130_fd_sc_hd__nand4_4
X_73377_ _73370_/Y _73371_/Y _73376_/X _73377_/Y sky130_fd_sc_hd__o21ai_4
X_70589_ _70578_/A _70959_/C sky130_fd_sc_hd__buf_2
Xclkbuf_opt_4_CLK _83248_/CLK _84895_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_10_685_0_CLK clkbuf_9_342_0_CLK/X _87195_/CLK sky130_fd_sc_hd__clkbuf_1
X_63130_ _63130_/A _63130_/X sky130_fd_sc_hd__buf_2
X_75116_ _75117_/B _75117_/C _75117_/A _75116_/X sky130_fd_sc_hd__a21o_4
X_41508_ _41507_/X _41486_/X _88202_/Q _41487_/X _41508_/X sky130_fd_sc_hd__a2bb2o_4
X_48064_ _48064_/A _48065_/A sky130_fd_sc_hd__inv_2
X_60342_ _60275_/X _60285_/Y _60306_/Y _79649_/A _60341_/X _60342_/X
+ sky130_fd_sc_hd__o32a_4
X_72328_ _72240_/X _85680_/Q _72241_/X _72328_/X sky130_fd_sc_hd__o21a_4
X_45276_ _45270_/X _45273_/Y _45275_/X _45276_/Y sky130_fd_sc_hd__a21oi_4
X_76096_ _76096_/A _81720_/D _76075_/B _76096_/Y sky130_fd_sc_hd__nand3_4
X_42488_ _42488_/A _42556_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_176_0_CLK clkbuf_8_88_0_CLK/X clkbuf_9_176_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_47015_ _83047_/Q _47016_/A sky130_fd_sc_hd__inv_2
X_44227_ _44225_/Y _44227_/Y sky130_fd_sc_hd__inv_2
X_63061_ _58421_/A _63010_/X _63059_/X _59467_/Y _63060_/X _63061_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75047_ _75047_/A _75047_/B _75039_/X _75051_/B _75047_/Y sky130_fd_sc_hd__nand4_4
X_79924_ _79920_/Y _79924_/B _79924_/C _79927_/A sky130_fd_sc_hd__nand3_4
X_41439_ _40586_/A _41471_/B sky130_fd_sc_hd__buf_2
X_60273_ _60273_/A _60273_/X sky130_fd_sc_hd__buf_2
X_72259_ _72258_/X _85686_/Q _72146_/X _72259_/X sky130_fd_sc_hd__o21a_4
X_62012_ _61548_/B _61995_/X _62010_/X _62011_/X _62012_/Y sky130_fd_sc_hd__nand4_4
X_44158_ _60665_/C _44003_/X _44158_/Y sky130_fd_sc_hd__xnor2_4
X_79855_ _79854_/B _79835_/X _79840_/A _79827_/Y _79855_/X sky130_fd_sc_hd__a211o_4
X_43109_ _43105_/X _43106_/X _40753_/X _43107_/Y _43108_/X _43109_/Y
+ sky130_fd_sc_hd__o32ai_4
X_66820_ _87433_/Q _66797_/X _66747_/X _66819_/X _66820_/X sky130_fd_sc_hd__a211o_4
X_78806_ _82546_/Q _78807_/A sky130_fd_sc_hd__inv_2
X_48966_ _48904_/A _49009_/B sky130_fd_sc_hd__buf_2
X_44089_ _44052_/A _44090_/B sky130_fd_sc_hd__buf_2
X_79786_ _79782_/X _79785_/Y _79786_/X sky130_fd_sc_hd__xor2_4
X_76998_ _60931_/C _76998_/B _76998_/X sky130_fd_sc_hd__xor2_4
X_47917_ _47917_/A _50270_/A sky130_fd_sc_hd__buf_2
X_66751_ _66608_/A _66751_/X sky130_fd_sc_hd__buf_2
X_78737_ _78732_/X _78735_/Y _78733_/Y _78737_/Y sky130_fd_sc_hd__nand3_4
X_63963_ _60871_/Y _64179_/B sky130_fd_sc_hd__buf_2
X_75949_ _75949_/A _75948_/Y _81734_/D sky130_fd_sc_hd__xor2_4
X_48897_ _48897_/A _48898_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_623_0_CLK clkbuf_9_311_0_CLK/X _86758_/CLK sky130_fd_sc_hd__clkbuf_1
X_65702_ _65702_/A _85871_/Q _65702_/X sky130_fd_sc_hd__and2_4
X_62914_ _62912_/X _62893_/X _62913_/Y _84371_/D sky130_fd_sc_hd__a21oi_4
X_69470_ _87515_/Q _69468_/X _69343_/X _69469_/X _69470_/X sky130_fd_sc_hd__a211o_4
X_47848_ _51282_/A _47848_/X sky130_fd_sc_hd__buf_2
X_66682_ _57866_/A _66682_/X sky130_fd_sc_hd__buf_2
X_78668_ _78663_/X _78666_/Y _78664_/Y _78669_/B sky130_fd_sc_hd__nand3_4
X_63894_ _61438_/X _63877_/B _63894_/C _63877_/D _63894_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_9_114_0_CLK clkbuf_8_57_0_CLK/X clkbuf_9_114_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_68421_ _44245_/A _68421_/X sky130_fd_sc_hd__buf_2
X_65633_ _84188_/Q _65634_/C sky130_fd_sc_hd__inv_2
X_77619_ _77614_/X _77619_/B _77619_/C _77666_/A sky130_fd_sc_hd__nand3_4
Xclkbuf_9_41_0_CLK clkbuf_8_20_0_CLK/X clkbuf_9_41_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_62845_ _60274_/X _62889_/D sky130_fd_sc_hd__buf_2
X_47779_ _47779_/A _47780_/A sky130_fd_sc_hd__inv_2
X_78599_ _78623_/B _78623_/A _78599_/X sky130_fd_sc_hd__xor2_4
X_49518_ _49502_/A _51043_/B _49518_/Y sky130_fd_sc_hd__nand2_4
X_80630_ _80625_/X _80630_/B _80633_/C sky130_fd_sc_hd__xnor2_4
X_68352_ _68344_/X _68351_/X _58002_/A _68352_/X sky130_fd_sc_hd__a21o_4
X_65564_ _65779_/A _73012_/B _65564_/X sky130_fd_sc_hd__and2_4
X_50790_ _50777_/A _46396_/B _50790_/Y sky130_fd_sc_hd__nand2_4
X_62776_ _62717_/A _62789_/D sky130_fd_sc_hd__buf_2
Xclkbuf_10_638_0_CLK clkbuf_9_319_0_CLK/X _82288_/CLK sky130_fd_sc_hd__clkbuf_1
X_67303_ _67141_/X _67292_/Y _67269_/X _67302_/Y _67303_/X sky130_fd_sc_hd__a211o_4
X_64515_ _64515_/A _59433_/A _64515_/C _64515_/Y sky130_fd_sc_hd__nand3_4
X_49449_ _49454_/A _50971_/B _49449_/Y sky130_fd_sc_hd__nand2_4
X_61727_ _59824_/B _61728_/A sky130_fd_sc_hd__buf_2
X_80561_ _80557_/X _80561_/B _80561_/X sky130_fd_sc_hd__xor2_4
X_68283_ _68208_/X _68283_/X sky130_fd_sc_hd__buf_2
X_65495_ _64730_/X _65647_/B _64735_/X _65495_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_9_129_0_CLK clkbuf_8_64_0_CLK/X clkbuf_9_129_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_82300_ _82299_/CLK _82300_/D _40790_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_56_0_CLK clkbuf_9_57_0_CLK/A clkbuf_9_56_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_67234_ _67141_/X _67220_/Y _67152_/X _67233_/Y _67234_/X sky130_fd_sc_hd__a211o_4
X_52460_ _52466_/A _53980_/B _52460_/Y sky130_fd_sc_hd__nand2_4
X_64446_ _63611_/A _64419_/B _64446_/Y sky130_fd_sc_hd__nor2_4
X_83280_ _83711_/CLK _83280_/D _83280_/Q sky130_fd_sc_hd__dfxtp_4
X_61658_ _61649_/Y _61652_/Y _61594_/X _61655_/Y _61657_/Y _61658_/X
+ sky130_fd_sc_hd__a41o_4
X_80492_ _80471_/B _80488_/X _80491_/Y _80492_/Y sky130_fd_sc_hd__a21oi_4
X_51411_ _51410_/X _51230_/X _51225_/C _52938_/D _51411_/X sky130_fd_sc_hd__and4_4
X_82231_ _82515_/CLK _82263_/Q _77538_/B sky130_fd_sc_hd__dfxtp_4
X_60609_ _60399_/Y _60488_/C _60583_/Y _60608_/X _60609_/X sky130_fd_sc_hd__a211o_4
X_67165_ _84081_/Q _67092_/X _67164_/X _67165_/X sky130_fd_sc_hd__a21bo_4
X_52391_ _50693_/A _50693_/B _52295_/A _52391_/X sky130_fd_sc_hd__o21a_4
X_64377_ _64377_/A _64377_/X sky130_fd_sc_hd__buf_2
X_61589_ _72561_/C _61590_/C sky130_fd_sc_hd__buf_2
X_54130_ _54134_/A _54130_/B _54130_/Y sky130_fd_sc_hd__nand2_4
X_66116_ _66113_/X _66115_/X _65961_/X _66116_/X sky130_fd_sc_hd__a21o_4
X_51342_ _53671_/A _51352_/C sky130_fd_sc_hd__buf_2
X_63328_ _79198_/A _63310_/X _63327_/X _63328_/Y sky130_fd_sc_hd__o21ai_4
X_82162_ _82746_/CLK _66138_/A _82162_/Q sky130_fd_sc_hd__dfxtp_4
X_67096_ _87933_/Q _66994_/X _67046_/X _67095_/X _67096_/X sky130_fd_sc_hd__a211o_4
X_81113_ _80728_/CLK _79802_/X _81113_/Q sky130_fd_sc_hd__dfxtp_4
X_54061_ _54031_/A _50850_/B _54061_/Y sky130_fd_sc_hd__nand2_4
X_66047_ _84160_/Q _66048_/C sky130_fd_sc_hd__inv_2
X_51273_ _64794_/B _51259_/X _51272_/Y _51273_/Y sky130_fd_sc_hd__o21ai_4
X_63259_ _63010_/A _63259_/X sky130_fd_sc_hd__buf_2
X_86970_ _87472_/CLK _86970_/D _86970_/Q sky130_fd_sc_hd__dfxtp_4
X_82093_ _82139_/CLK _82093_/D _82093_/Q sky130_fd_sc_hd__dfxtp_4
X_53012_ _53025_/A _53012_/B _53012_/Y sky130_fd_sc_hd__nand2_4
X_50224_ _51737_/A _50224_/B _50224_/Y sky130_fd_sc_hd__nand2_4
X_85921_ _83161_/CLK _85921_/D _73561_/B sky130_fd_sc_hd__dfxtp_4
X_81044_ _81117_/CLK _75345_/X _81044_/Q sky130_fd_sc_hd__dfxtp_4
X_57820_ _57806_/X _57820_/B _57820_/Y sky130_fd_sc_hd__nor2_4
X_69806_ _73225_/A _69747_/X _69617_/X _69805_/Y _69806_/X sky130_fd_sc_hd__a211o_4
X_50155_ _48833_/A _51256_/B sky130_fd_sc_hd__buf_2
X_85852_ _85566_/CLK _52292_/Y _64753_/B sky130_fd_sc_hd__dfxtp_4
X_67998_ _67972_/A _87703_/Q _67998_/X sky130_fd_sc_hd__and2_4
X_84803_ _86713_/CLK _84803_/D _84803_/Q sky130_fd_sc_hd__dfxtp_4
X_57751_ _57748_/Y _57750_/Y _57718_/X _57751_/X sky130_fd_sc_hd__a21o_4
X_69737_ _69687_/A _69737_/B _69737_/Y sky130_fd_sc_hd__nor2_4
X_50086_ _50069_/A _71989_/B _50086_/X sky130_fd_sc_hd__and2_4
X_54963_ _54888_/A _54964_/A sky130_fd_sc_hd__buf_2
X_66949_ _87875_/Q _66875_/X _66926_/X _66948_/X _66949_/X sky130_fd_sc_hd__a211o_4
X_85783_ _82956_/CLK _85783_/D _85783_/Q sky130_fd_sc_hd__dfxtp_4
X_82995_ _85075_/CLK _82995_/D _82995_/Q sky130_fd_sc_hd__dfxtp_4
X_56702_ _56702_/A _56685_/B _56702_/X sky130_fd_sc_hd__and2_4
X_87522_ _88034_/CLK _87522_/D _87522_/Q sky130_fd_sc_hd__dfxtp_4
X_53914_ _53838_/A _53914_/X sky130_fd_sc_hd__buf_2
X_84734_ _83438_/CLK _84734_/D _59433_/A sky130_fd_sc_hd__dfxtp_4
X_57682_ _57682_/A _57682_/Y sky130_fd_sc_hd__inv_2
X_81946_ _81970_/CLK _77944_/B _81946_/Q sky130_fd_sc_hd__dfxtp_4
X_69668_ _69663_/X _69668_/B _69668_/Y sky130_fd_sc_hd__nand2_4
X_54894_ _54893_/X _54894_/B _54894_/Y sky130_fd_sc_hd__nand2_4
X_59421_ _59421_/A _59424_/B _59421_/Y sky130_fd_sc_hd__nand2_4
X_56633_ _55503_/D _56632_/Y _56633_/X sky130_fd_sc_hd__xor2_4
X_68619_ _88105_/Q _68467_/X _68617_/X _68618_/Y _68619_/X sky130_fd_sc_hd__a211o_4
X_87453_ _87446_/CLK _43377_/Y _87453_/Q sky130_fd_sc_hd__dfxtp_4
X_53845_ _53842_/Y _53838_/X _53844_/Y _53845_/Y sky130_fd_sc_hd__a21boi_4
X_84665_ _84508_/CLK _60082_/Y _80082_/A sky130_fd_sc_hd__dfxtp_4
X_81877_ _81872_/CLK _78068_/X _81877_/Q sky130_fd_sc_hd__dfxtp_4
X_69599_ _69596_/X _69598_/X _69599_/Y sky130_fd_sc_hd__nand2_4
X_86404_ _86404_/CLK _86404_/D _65367_/B sky130_fd_sc_hd__dfxtp_4
X_40810_ _40810_/A _40810_/X sky130_fd_sc_hd__buf_2
X_59352_ _59348_/Y _59350_/Y _59351_/X _59352_/X sky130_fd_sc_hd__a21o_4
X_71630_ _71655_/A _71641_/A sky130_fd_sc_hd__buf_2
X_83616_ _85558_/CLK _83616_/D _48972_/A sky130_fd_sc_hd__dfxtp_4
X_56564_ _56564_/A _56564_/B _56564_/C _56564_/D _56931_/A sky130_fd_sc_hd__nand4_4
X_80828_ _83944_/CLK _83972_/Q _75657_/B sky130_fd_sc_hd__dfxtp_4
X_87384_ _88215_/CLK _43511_/Y _87384_/Q sky130_fd_sc_hd__dfxtp_4
X_41790_ _40402_/A _41452_/A _41789_/X _41790_/X sky130_fd_sc_hd__o21a_4
X_53776_ _53791_/A _48704_/Y _53776_/Y sky130_fd_sc_hd__nand2_4
X_84596_ _82452_/CLK _84596_/D _79136_/A sky130_fd_sc_hd__dfxtp_4
X_50988_ _86094_/Q _50965_/X _50987_/Y _50988_/Y sky130_fd_sc_hd__o21ai_4
X_58303_ _58303_/A _58303_/Y sky130_fd_sc_hd__inv_2
X_55515_ _45567_/A _55511_/X _55513_/X _55514_/Y _55515_/X sky130_fd_sc_hd__a211o_4
X_86335_ _86655_/CLK _86335_/D _57731_/B sky130_fd_sc_hd__dfxtp_4
X_52727_ _85765_/Q _52711_/X _52726_/Y _52727_/Y sky130_fd_sc_hd__o21ai_4
X_40741_ _40741_/A _40760_/B _40741_/X sky130_fd_sc_hd__or2_4
X_71561_ _71586_/A _71553_/B _71558_/X _71561_/Y sky130_fd_sc_hd__nor3_4
X_59283_ _59253_/X _59281_/Y _59282_/Y _59271_/X _59258_/X _59283_/X
+ sky130_fd_sc_hd__o32a_4
X_83547_ _85354_/CLK _83547_/D _83547_/Q sky130_fd_sc_hd__dfxtp_4
X_56495_ _56064_/X _56483_/X _56494_/Y _56495_/Y sky130_fd_sc_hd__o21ai_4
X_80759_ _81134_/CLK _80759_/D _81135_/D sky130_fd_sc_hd__dfxtp_4
X_73300_ _43170_/Y _73298_/X _73251_/X _73299_/Y _73300_/X sky130_fd_sc_hd__a211o_4
X_70512_ _57655_/Y _70501_/X _70511_/Y _83760_/D sky130_fd_sc_hd__o21ai_4
XPHY_600 sky130_fd_sc_hd__decap_3
X_58234_ _58230_/A _58233_/Y _58234_/Y sky130_fd_sc_hd__nand2_4
X_43460_ _43449_/X _43452_/X _41631_/X _87411_/Q _43456_/X _43461_/A
+ sky130_fd_sc_hd__o32ai_4
X_55446_ _55446_/A _55328_/X _55446_/X sky130_fd_sc_hd__and2_4
X_74280_ _74268_/X _74281_/C _74279_/X _74280_/X sky130_fd_sc_hd__a21o_4
X_86266_ _85562_/CLK _50094_/Y _64804_/B sky130_fd_sc_hd__dfxtp_4
XPHY_611 sky130_fd_sc_hd__decap_3
X_40672_ _40670_/X _82866_/Q _40671_/X _40672_/Y sky130_fd_sc_hd__o21ai_4
X_52658_ _52657_/X _52658_/B _52658_/Y sky130_fd_sc_hd__nand2_4
X_71492_ _71488_/X _71297_/X _71496_/C _71492_/X sky130_fd_sc_hd__and3_4
X_83478_ _83415_/CLK _71497_/X _83478_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_622 sky130_fd_sc_hd__decap_3
XPHY_633 sky130_fd_sc_hd__decap_3
X_42411_ _41872_/A _42411_/X sky130_fd_sc_hd__buf_2
X_88005_ _88006_/CLK _88005_/D _88005_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_644 sky130_fd_sc_hd__decap_3
X_73231_ _88321_/Q _73086_/X _73202_/X _73231_/X sky130_fd_sc_hd__o21a_4
X_85217_ _85249_/CLK _85217_/D _85217_/Q sky130_fd_sc_hd__dfxtp_4
X_51609_ _51619_/A _51603_/B _51608_/X _53133_/D _51609_/X sky130_fd_sc_hd__and4_4
X_70443_ _50293_/B _70422_/X _70442_/Y _70443_/Y sky130_fd_sc_hd__o21ai_4
X_58165_ _58153_/X _83493_/Q _58164_/Y _58165_/X sky130_fd_sc_hd__o21a_4
XPHY_655 sky130_fd_sc_hd__decap_3
X_82429_ _84197_/CLK _82429_/D _78710_/A sky130_fd_sc_hd__dfxtp_4
X_55377_ _55374_/Y _55375_/A _55377_/Y sky130_fd_sc_hd__nand2_4
X_43391_ _43390_/Y _87446_/D sky130_fd_sc_hd__inv_2
X_86197_ _86191_/CLK _50457_/Y _86197_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_666 sky130_fd_sc_hd__decap_3
X_52589_ _52587_/Y _52532_/X _52588_/X _52589_/Y sky130_fd_sc_hd__a21oi_4
XPHY_677 sky130_fd_sc_hd__decap_3
XPHY_688 sky130_fd_sc_hd__decap_3
X_45130_ _45119_/X _45126_/Y _45129_/Y _45130_/Y sky130_fd_sc_hd__a21oi_4
X_57116_ _56960_/X _85079_/Q _57112_/X _57116_/Y sky130_fd_sc_hd__nor3_4
X_54328_ _85462_/Q _54320_/X _54327_/Y _54328_/Y sky130_fd_sc_hd__o21ai_4
X_42342_ _42290_/A _42342_/X sky130_fd_sc_hd__buf_2
X_73162_ _73159_/X _73161_/X _72877_/X _73168_/A sky130_fd_sc_hd__a21o_4
XPHY_699 sky130_fd_sc_hd__decap_3
X_85148_ _85114_/CLK _85148_/D _85148_/Q sky130_fd_sc_hd__dfxtp_4
X_70374_ _70809_/A _70374_/X sky130_fd_sc_hd__buf_2
X_58096_ _58576_/A _58096_/B _58096_/Y sky130_fd_sc_hd__nor2_4
X_72113_ _72113_/A _72113_/B _72048_/X _72113_/X sky130_fd_sc_hd__and3_4
X_45061_ _55896_/B _45060_/X _45040_/X _45061_/X sky130_fd_sc_hd__o21a_4
X_57047_ _56761_/X _57046_/Y _57038_/B _57047_/Y sky130_fd_sc_hd__o21ai_4
X_42273_ _41507_/X _42271_/X _87946_/Q _42272_/X _87946_/D sky130_fd_sc_hd__a2bb2o_4
X_54259_ _54255_/A _54246_/X _54255_/C _53090_/D _54259_/X sky130_fd_sc_hd__and4_4
X_73093_ _73093_/A _65612_/B _73093_/X sky130_fd_sc_hd__and2_4
X_77970_ _82172_/Q _77970_/B _77970_/X sky130_fd_sc_hd__xor2_4
X_85079_ _85013_/CLK _85079_/D _85079_/Q sky130_fd_sc_hd__dfxtp_4
X_44012_ _44012_/A _64806_/A sky130_fd_sc_hd__buf_2
X_41224_ _41136_/X _40705_/A _41223_/X _41224_/X sky130_fd_sc_hd__o21a_4
X_72044_ _49060_/A _72043_/X _71964_/X _72044_/X sky130_fd_sc_hd__and3_4
X_76921_ _76920_/Y _76921_/Y sky130_fd_sc_hd__inv_2
X_48820_ _48831_/A _48820_/B _48820_/Y sky130_fd_sc_hd__nand2_4
X_79640_ _79627_/Y _79630_/X _79642_/B sky130_fd_sc_hd__or2_4
X_41155_ _41159_/A _81145_/Q _41155_/X sky130_fd_sc_hd__or2_4
X_76852_ _76841_/A _76840_/Y _76851_/X _76852_/Y sky130_fd_sc_hd__a21oi_4
X_58998_ _58918_/X _58996_/Y _58997_/Y _58959_/X _58923_/X _58998_/X
+ sky130_fd_sc_hd__o32a_4
X_75803_ _75793_/B _75793_/A _75803_/C _75810_/A sky130_fd_sc_hd__nand3_4
X_48751_ _65551_/B _48730_/X _48750_/Y _48751_/Y sky130_fd_sc_hd__o21ai_4
X_79571_ _79571_/A _79573_/B sky130_fd_sc_hd__inv_2
X_45963_ _45962_/X _45963_/X sky130_fd_sc_hd__buf_2
X_41086_ _41073_/X _81702_/Q _41085_/X _41086_/X sky130_fd_sc_hd__o21a_4
X_57949_ _57947_/X _85713_/Q _57948_/X _57949_/X sky130_fd_sc_hd__o21a_4
X_76783_ _81584_/Q _76783_/B _81552_/D sky130_fd_sc_hd__xor2_4
X_73995_ _44126_/X _66168_/B _73995_/X sky130_fd_sc_hd__and2_4
X_47702_ _47692_/A _47739_/B _47692_/C _53196_/D _47702_/X sky130_fd_sc_hd__and4_4
X_78522_ _82801_/Q _78522_/Y sky130_fd_sc_hd__inv_2
X_44914_ _56469_/C _44882_/X _44884_/X _44914_/X sky130_fd_sc_hd__o21a_4
X_75734_ _75734_/A _75733_/Y _75735_/A sky130_fd_sc_hd__xor2_4
X_48682_ _48682_/A _48683_/A sky130_fd_sc_hd__inv_2
X_60960_ _60950_/Y _60881_/Y _60952_/X _60958_/X _60959_/X _84548_/D
+ sky130_fd_sc_hd__o41a_4
X_72946_ _41999_/Y _72921_/X _72944_/X _72945_/Y _72946_/X sky130_fd_sc_hd__a211o_4
X_45894_ _45884_/Y _45886_/X _58517_/A _45893_/Y _45894_/X sky130_fd_sc_hd__a211o_4
X_47633_ _47649_/A _53157_/B _47633_/Y sky130_fd_sc_hd__nand2_4
X_59619_ _60162_/A _60403_/C _59775_/A _61294_/D _59619_/X sky130_fd_sc_hd__and4_4
X_78453_ _78475_/B _78453_/B _82764_/D sky130_fd_sc_hd__xor2_4
X_44845_ _44832_/X _44844_/X _41734_/X _86923_/Q _44833_/X _44846_/A
+ sky130_fd_sc_hd__o32ai_4
X_75665_ _75665_/A _75665_/B _75680_/A sky130_fd_sc_hd__nand2_4
X_60891_ _60890_/X _60891_/Y sky130_fd_sc_hd__inv_2
X_72877_ _72877_/A _72877_/X sky130_fd_sc_hd__buf_2
X_77404_ _77404_/A _82190_/D _81902_/D sky130_fd_sc_hd__xor2_4
X_62630_ _62629_/Y _59945_/Y _62186_/X _59931_/A _62630_/X sky130_fd_sc_hd__a2bb2o_4
X_74616_ _45305_/Y _74612_/X _74615_/X _83015_/D sky130_fd_sc_hd__o21ai_4
X_47564_ _86621_/Q _47524_/X _47563_/Y _47564_/Y sky130_fd_sc_hd__o21ai_4
X_71828_ _71825_/X _83361_/Q _71827_/X _83361_/D sky130_fd_sc_hd__a21o_4
X_78384_ _78385_/A _82664_/D _78384_/Y sky130_fd_sc_hd__nor2_4
X_44776_ _41355_/Y _44774_/X _86962_/Q _44775_/X _86962_/D sky130_fd_sc_hd__a2bb2o_4
X_75596_ _75588_/Y _75596_/B _75597_/B sky130_fd_sc_hd__xor2_4
X_41988_ _88080_/Q _41988_/Y sky130_fd_sc_hd__inv_2
X_49303_ _65109_/B _49300_/X _49302_/Y _49303_/Y sky130_fd_sc_hd__o21ai_4
X_46515_ _46403_/X _49119_/A _46514_/X _51356_/B sky130_fd_sc_hd__o21ai_4
X_77335_ _77320_/Y _77316_/A _77316_/B _77335_/Y sky130_fd_sc_hd__a21boi_4
X_43727_ _40881_/X _43695_/X _73299_/A _43696_/X _87294_/D sky130_fd_sc_hd__a2bb2o_4
X_74547_ _74541_/A _46215_/B _74547_/C _74547_/Y sky130_fd_sc_hd__nand3_4
X_62561_ _62559_/Y _62561_/B _62560_/Y _62561_/Y sky130_fd_sc_hd__nand3_4
X_40939_ _40938_/Y _40939_/X sky130_fd_sc_hd__buf_2
X_47495_ _47513_/A _47463_/X _47513_/C _53078_/D _47495_/X sky130_fd_sc_hd__and4_4
X_71759_ _52965_/B _71736_/X _71758_/Y _83386_/D sky130_fd_sc_hd__o21ai_4
X_64300_ _79806_/B _64255_/X _64299_/X _84258_/D sky130_fd_sc_hd__a21o_4
X_49234_ _48623_/A _49234_/X sky130_fd_sc_hd__buf_2
X_61512_ _61342_/X _61512_/X sky130_fd_sc_hd__buf_2
X_46446_ _46446_/A _46447_/B sky130_fd_sc_hd__inv_2
X_65280_ _65252_/X _86727_/Q _65230_/X _65279_/X _65280_/X sky130_fd_sc_hd__a211o_4
X_77266_ _77264_/Y _77265_/Y _82213_/Q _77266_/X sky130_fd_sc_hd__a21o_4
X_43658_ _40716_/X _43656_/X _74097_/A _43657_/X _87324_/D sky130_fd_sc_hd__a2bb2o_4
X_62492_ _61560_/B _62492_/B _62449_/X _62475_/X _62492_/Y sky130_fd_sc_hd__nand4_4
X_74478_ _48621_/A _74478_/B _74478_/C _74478_/X sky130_fd_sc_hd__and3_4
X_79005_ _79022_/A _79010_/A sky130_fd_sc_hd__inv_2
X_64231_ _64219_/Y _64230_/X _72577_/B _64231_/X sky130_fd_sc_hd__o21a_4
X_76217_ _76215_/Y _76216_/Y _76234_/A _76217_/X sky130_fd_sc_hd__a21o_4
X_42609_ _42568_/X _42569_/X _40899_/X _69897_/B _42571_/X _87802_/D
+ sky130_fd_sc_hd__o32ai_4
X_49165_ _49160_/Y _49138_/X _49164_/X _86438_/D sky130_fd_sc_hd__a21oi_4
X_61443_ _61442_/Y _61443_/Y sky130_fd_sc_hd__inv_2
X_73429_ _73476_/A _86503_/Q _73429_/X sky130_fd_sc_hd__and2_4
X_46377_ _46376_/Y _50781_/B sky130_fd_sc_hd__buf_2
X_77197_ _77189_/Y _77202_/A _77196_/Y _77198_/B sky130_fd_sc_hd__a21boi_4
X_43589_ _43588_/X _47832_/A sky130_fd_sc_hd__buf_2
X_48116_ _48142_/A _50370_/B _48116_/Y sky130_fd_sc_hd__nand2_4
X_45328_ _56450_/C _45326_/X _45327_/X _45328_/Y sky130_fd_sc_hd__o21ai_4
X_76148_ _76145_/Y _76147_/Y _76150_/A sky130_fd_sc_hd__nand2_4
X_64162_ _64162_/A _58360_/A _64173_/C _64162_/X sky130_fd_sc_hd__and3_4
X_49096_ _65164_/B _49052_/X _49095_/Y _49096_/Y sky130_fd_sc_hd__o21ai_4
X_61374_ _61374_/A _61375_/A sky130_fd_sc_hd__buf_2
X_63113_ _59390_/Y _63113_/B _63103_/C _63092_/D _63113_/X sky130_fd_sc_hd__or4_4
X_48047_ _52039_/A _48069_/B _47919_/X _48047_/X sky130_fd_sc_hd__and3_4
X_60325_ _60267_/X _60325_/B _60325_/C _60367_/D _60325_/Y sky130_fd_sc_hd__nand4_4
X_45259_ _45256_/X _45258_/Y _45200_/X _45259_/Y sky130_fd_sc_hd__a21oi_4
X_68970_ _68994_/A _68970_/B _68970_/X sky130_fd_sc_hd__and2_4
X_64093_ _83243_/Q _64158_/B _64158_/C _64045_/X _64094_/D sky130_fd_sc_hd__nand4_4
X_76079_ _81719_/D _76070_/B _76079_/Y sky130_fd_sc_hd__nand2_4
X_67921_ _67918_/X _67920_/X _67875_/X _67921_/Y sky130_fd_sc_hd__a21oi_4
X_63044_ _63044_/A _63004_/B _63081_/C _63033_/D _63044_/X sky130_fd_sc_hd__or4_4
X_79907_ _79906_/Y _79907_/B _79913_/A sky130_fd_sc_hd__nand2_4
X_60256_ _60268_/C _60300_/B _60325_/C _60256_/X sky130_fd_sc_hd__o21a_4
X_67852_ _84052_/Q _67806_/X _67851_/X _84052_/D sky130_fd_sc_hd__a21bo_4
X_79838_ _79836_/X _79838_/B _79854_/B sky130_fd_sc_hd__xnor2_4
X_60187_ _60187_/A _60204_/A sky130_fd_sc_hd__buf_2
X_49998_ _72377_/B _49986_/X _49997_/Y _49998_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_562_0_CLK clkbuf_9_281_0_CLK/X _88116_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_53_0_CLK clkbuf_6_53_0_CLK/A clkbuf_6_53_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_66803_ _88394_/Q _66751_/X _66801_/X _66802_/X _66803_/X sky130_fd_sc_hd__a211o_4
X_48949_ _52295_/B _71989_/B sky130_fd_sc_hd__buf_2
X_67783_ _67690_/X _87648_/Q _67783_/X sky130_fd_sc_hd__and2_4
X_79769_ _79757_/A _79756_/Y _79768_/X _79769_/X sky130_fd_sc_hd__a21o_4
X_64995_ _64995_/A _64994_/Y _64995_/Y sky130_fd_sc_hd__nand2_4
X_81800_ _81684_/CLK _81800_/D _47464_/A sky130_fd_sc_hd__dfxtp_4
X_69522_ _88023_/Q _69368_/X _69478_/X _69521_/X _69522_/X sky130_fd_sc_hd__a211o_4
X_66734_ _66971_/A _66734_/X sky130_fd_sc_hd__buf_2
X_51960_ _51928_/X _51960_/X sky130_fd_sc_hd__buf_2
X_63946_ _63751_/X _64025_/D sky130_fd_sc_hd__buf_2
X_82780_ _83783_/CLK _82780_/D _82780_/Q sky130_fd_sc_hd__dfxtp_4
X_50911_ _50728_/A _50932_/A sky130_fd_sc_hd__buf_2
X_81731_ _84020_/CLK _75929_/B _41784_/B sky130_fd_sc_hd__dfxtp_4
X_69453_ _88028_/Q _69315_/X _69393_/X _69452_/X _69453_/X sky130_fd_sc_hd__a211o_4
X_66665_ _66664_/X _86802_/Q _66665_/X sky130_fd_sc_hd__and2_4
X_51891_ _52679_/A _52626_/A sky130_fd_sc_hd__buf_2
X_63877_ _61428_/X _63877_/B _63814_/C _63877_/D _63877_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_10_577_0_CLK clkbuf_9_288_0_CLK/X _80813_/CLK sky130_fd_sc_hd__clkbuf_1
X_68404_ _88018_/Q _68402_/X _68359_/X _68403_/X _68404_/X sky130_fd_sc_hd__a211o_4
X_53630_ _50724_/A _53658_/B sky130_fd_sc_hd__buf_2
X_65616_ _65753_/A _73096_/B _65616_/X sky130_fd_sc_hd__and2_4
X_84450_ _84449_/CLK _61850_/Y _78073_/B sky130_fd_sc_hd__dfxtp_4
X_50842_ _50806_/A _49320_/B _50842_/Y sky130_fd_sc_hd__nand2_4
X_62828_ _62979_/A _62971_/A sky130_fd_sc_hd__buf_2
X_81662_ _81680_/CLK _76755_/A _76572_/A sky130_fd_sc_hd__dfxtp_4
X_69384_ _87521_/Q _69356_/X _69371_/X _69383_/X _69384_/X sky130_fd_sc_hd__a211o_4
X_66596_ _87134_/Q _66593_/X _66594_/X _66595_/X _66596_/X sky130_fd_sc_hd__a211o_4
X_83401_ _84939_/CLK _83401_/D _83401_/Q sky130_fd_sc_hd__dfxtp_4
X_80613_ _84776_/Q _84168_/Q _80613_/X sky130_fd_sc_hd__xor2_4
X_68335_ _68056_/X _68061_/X _68327_/X _68335_/Y sky130_fd_sc_hd__a21oi_4
X_53561_ _52039_/A _53620_/B _53492_/X _53561_/X sky130_fd_sc_hd__and3_4
X_65547_ _65545_/Y _65529_/X _65546_/X _65547_/X sky130_fd_sc_hd__a21o_4
X_84381_ _84520_/CLK _84381_/D _62806_/C sky130_fd_sc_hd__dfxtp_4
X_50773_ _50764_/A _52468_/B _50773_/Y sky130_fd_sc_hd__nand2_4
X_62759_ _60211_/A _62759_/X sky130_fd_sc_hd__buf_2
X_81593_ _81428_/CLK _65559_/C _81593_/Q sky130_fd_sc_hd__dfxtp_4
X_55300_ _55168_/X _55300_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_500_0_CLK clkbuf_9_250_0_CLK/X _86096_/CLK sky130_fd_sc_hd__clkbuf_1
X_86120_ _86121_/CLK _86120_/D _86120_/Q sky130_fd_sc_hd__dfxtp_4
X_52512_ _65074_/B _52500_/X _52511_/Y _52512_/Y sky130_fd_sc_hd__o21ai_4
X_83332_ _83753_/CLK _71909_/Y _83332_/Q sky130_fd_sc_hd__dfxtp_4
X_56280_ _56280_/A _56177_/B _56280_/C _56280_/Y sky130_fd_sc_hd__nand3_4
X_80544_ _80551_/B _80544_/B _80544_/X sky130_fd_sc_hd__xor2_4
X_68266_ _83997_/Q _68259_/X _68265_/X _68266_/X sky130_fd_sc_hd__a21bo_4
X_53492_ _53671_/A _53492_/X sky130_fd_sc_hd__buf_2
X_65478_ _65984_/A _65647_/B sky130_fd_sc_hd__buf_2
X_55231_ _55125_/A _55231_/B _55231_/Y sky130_fd_sc_hd__nor2_4
X_67217_ _67214_/X _67216_/X _67147_/X _67220_/A sky130_fd_sc_hd__a21o_4
X_86051_ _85635_/CLK _86051_/D _86051_/Q sky130_fd_sc_hd__dfxtp_4
X_52443_ _52441_/Y _52430_/X _52442_/Y _52443_/Y sky130_fd_sc_hd__a21boi_4
X_64429_ _65296_/A _64429_/X sky130_fd_sc_hd__buf_2
X_83263_ _86289_/CLK _83263_/D _83263_/Q sky130_fd_sc_hd__dfxtp_4
X_80475_ _80475_/A _80475_/B _80476_/B sky130_fd_sc_hd__xor2_4
X_68197_ _67229_/X _67232_/X _68173_/X _68197_/Y sky130_fd_sc_hd__a21oi_4
X_85002_ _83335_/CLK _57452_/Y _57448_/A sky130_fd_sc_hd__dfxtp_4
X_82214_ _82220_/CLK _82246_/Q _82214_/Q sky130_fd_sc_hd__dfxtp_4
X_55162_ _55139_/X _83747_/Q _55146_/X _55162_/Y sky130_fd_sc_hd__nand3_4
X_67148_ _67143_/X _67146_/X _67147_/X _67148_/X sky130_fd_sc_hd__a21o_4
X_52374_ _52373_/X _50674_/B _52374_/Y sky130_fd_sc_hd__nand2_4
X_83194_ _83191_/CLK _72676_/X _83194_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_515_0_CLK clkbuf_9_257_0_CLK/X _81428_/CLK sky130_fd_sc_hd__clkbuf_1
X_54113_ _53351_/A _54113_/X sky130_fd_sc_hd__buf_2
X_51325_ _86031_/Q _51309_/X _51324_/Y _51325_/Y sky130_fd_sc_hd__o21ai_4
X_82145_ _82145_/CLK _82145_/D _82101_/D sky130_fd_sc_hd__dfxtp_4
X_55093_ _55093_/A _47771_/Y _55093_/Y sky130_fd_sc_hd__nand2_4
X_59970_ _59969_/X _60042_/A sky130_fd_sc_hd__inv_2
X_67079_ _67057_/A _67079_/B _67079_/X sky130_fd_sc_hd__and2_4
X_58921_ _58921_/A _58898_/B _58921_/Y sky130_fd_sc_hd__nor2_4
X_54044_ _54042_/Y _54015_/X _54043_/X _54044_/Y sky130_fd_sc_hd__a21oi_4
X_51256_ _51256_/A _51256_/B _51330_/C _51256_/X sky130_fd_sc_hd__and3_4
X_86953_ _88220_/CLK _86953_/D _86953_/Q sky130_fd_sc_hd__dfxtp_4
X_82076_ _81160_/CLK _82076_/D _77964_/A sky130_fd_sc_hd__dfxtp_4
X_70090_ _69603_/X _69951_/Y _70081_/X _70089_/Y _70090_/X sky130_fd_sc_hd__a211o_4
X_50207_ _50187_/X _50721_/B _50207_/Y sky130_fd_sc_hd__nand2_4
X_85904_ _86576_/CLK _85904_/D _66153_/B sky130_fd_sc_hd__dfxtp_4
X_81027_ _82786_/CLK _81027_/D _81027_/Q sky130_fd_sc_hd__dfxtp_4
X_58852_ _58721_/A _59090_/B sky130_fd_sc_hd__buf_2
X_51187_ _51177_/A _51192_/B _51192_/C _52879_/D _51187_/X sky130_fd_sc_hd__and4_4
X_86884_ _86869_/CLK _45323_/Y _63312_/B sky130_fd_sc_hd__dfxtp_4
X_57803_ _57803_/A _57804_/A sky130_fd_sc_hd__buf_2
X_50138_ _50064_/A _50153_/A sky130_fd_sc_hd__buf_2
X_85835_ _86155_/CLK _52378_/Y _85835_/Q sky130_fd_sc_hd__dfxtp_4
X_58783_ _58703_/X _85456_/Q _58782_/X _58783_/Y sky130_fd_sc_hd__o21ai_4
X_55995_ _55993_/Y _55994_/X _56083_/C _55854_/X _55995_/X sky130_fd_sc_hd__and4_4
X_72800_ _72800_/A _72924_/B _72800_/Y sky130_fd_sc_hd__nor2_4
X_57734_ _57734_/A _57833_/B _57734_/Y sky130_fd_sc_hd__nor2_4
X_42960_ _42960_/A _87630_/D sky130_fd_sc_hd__inv_2
X_50069_ _50069_/A _71970_/B _50069_/X sky130_fd_sc_hd__and2_4
X_54946_ _54955_/A _54942_/B _46617_/A _53253_/D _54946_/X sky130_fd_sc_hd__and4_4
X_73780_ _73733_/A _73780_/B _73780_/X sky130_fd_sc_hd__and2_4
X_85766_ _85767_/CLK _52725_/Y _85766_/Q sky130_fd_sc_hd__dfxtp_4
X_70992_ _70990_/A _70945_/B _70990_/C _70992_/Y sky130_fd_sc_hd__nand3_4
X_82978_ _82980_/CLK _74706_/X _45875_/A sky130_fd_sc_hd__dfxtp_4
X_41911_ _41911_/A _41912_/A sky130_fd_sc_hd__buf_2
X_87505_ _87520_/CLK _43275_/Y _87505_/Q sky130_fd_sc_hd__dfxtp_4
X_72731_ _72730_/X _72731_/X sky130_fd_sc_hd__buf_2
X_84717_ _84903_/CLK _84717_/D _84717_/Q sky130_fd_sc_hd__dfxtp_4
X_57665_ _57665_/A _57666_/B sky130_fd_sc_hd__buf_2
X_81929_ _82234_/CLK _77786_/X _81929_/Q sky130_fd_sc_hd__dfxtp_4
X_54877_ _85361_/Q _54865_/X _54876_/Y _54877_/Y sky130_fd_sc_hd__o21ai_4
X_42891_ _41636_/X _42886_/X _67356_/B _42887_/X _87666_/D sky130_fd_sc_hd__a2bb2o_4
X_85697_ _85697_/CLK _53104_/Y _85697_/Q sky130_fd_sc_hd__dfxtp_4
X_59404_ _59394_/X _83486_/Q _59403_/Y _84742_/D sky130_fd_sc_hd__o21a_4
X_56616_ _56616_/A _56616_/B _56617_/A sky130_fd_sc_hd__and2_4
X_44630_ _44622_/X _44623_/X _41009_/A _87026_/Q _44625_/X _44631_/A
+ sky130_fd_sc_hd__o32ai_4
X_75450_ _75438_/Y _75431_/X _75432_/Y _75450_/Y sky130_fd_sc_hd__a21boi_4
X_87436_ _87436_/CLK _43409_/Y _87436_/Q sky130_fd_sc_hd__dfxtp_4
X_53828_ _85560_/Q _53784_/X _53827_/Y _53828_/Y sky130_fd_sc_hd__o21ai_4
X_41842_ _41839_/X _41841_/X _40491_/X _88127_/Q _41835_/X _41843_/A
+ sky130_fd_sc_hd__o32ai_4
X_72662_ _72668_/A _72668_/B _72662_/C _72662_/Y sky130_fd_sc_hd__nand3_4
X_84648_ _84645_/CLK _60231_/Y _79872_/A sky130_fd_sc_hd__dfxtp_4
X_57596_ _84972_/Q _57550_/X _57595_/Y _57596_/Y sky130_fd_sc_hd__o21ai_4
X_74401_ _48440_/A _74395_/X _74421_/C _74401_/X sky130_fd_sc_hd__and3_4
X_59335_ _59311_/X _85734_/Q _59334_/X _59335_/X sky130_fd_sc_hd__o21a_4
X_71613_ _71604_/X _83439_/Q _71612_/Y _71613_/X sky130_fd_sc_hd__a21o_4
X_44561_ _44547_/X _44548_/X _40854_/X _87054_/Q _44549_/X _44562_/A
+ sky130_fd_sc_hd__o32ai_4
X_56547_ _72739_/A _56547_/X sky130_fd_sc_hd__buf_2
X_75381_ _75380_/Y _75381_/B _75382_/A sky130_fd_sc_hd__nand2_4
X_41773_ _41772_/X _41773_/X sky130_fd_sc_hd__buf_2
X_87367_ _86824_/CLK _43544_/Y _87367_/Q sky130_fd_sc_hd__dfxtp_4
X_53759_ _48667_/A _53774_/B _53748_/C _53759_/X sky130_fd_sc_hd__and3_4
X_72593_ _72546_/Y _59621_/X _72539_/Y _72510_/Y _72592_/Y _72593_/X
+ sky130_fd_sc_hd__a41o_4
X_84579_ _84454_/CLK _84579_/D _78074_/A sky130_fd_sc_hd__dfxtp_4
X_46300_ _72083_/A _46300_/X sky130_fd_sc_hd__buf_2
X_77120_ _77111_/A _82290_/D _77120_/Y sky130_fd_sc_hd__nand2_4
X_43512_ _41778_/X _43498_/X _87383_/Q _43499_/X _43512_/X sky130_fd_sc_hd__a2bb2o_4
X_74332_ _74338_/A _74338_/B _55994_/X _74332_/Y sky130_fd_sc_hd__nand3_4
X_86318_ _86637_/CLK _86318_/D _57991_/B sky130_fd_sc_hd__dfxtp_4
X_40724_ _40723_/X _40724_/X sky130_fd_sc_hd__buf_2
X_47280_ _86651_/Q _47240_/X _47279_/Y _47280_/Y sky130_fd_sc_hd__o21ai_4
X_59266_ _59262_/Y _59265_/Y _59140_/X _59266_/X sky130_fd_sc_hd__a21o_4
X_71544_ _70679_/A _71546_/B _71546_/C _71544_/Y sky130_fd_sc_hd__nor3_4
X_56478_ _56026_/X _56468_/X _56477_/Y _85181_/D sky130_fd_sc_hd__o21ai_4
X_44492_ _44491_/Y _87082_/D sky130_fd_sc_hd__inv_2
X_87298_ _87814_/CLK _43715_/Y _43713_/A sky130_fd_sc_hd__dfxtp_4
X_46231_ _46230_/X _86770_/Q _45909_/X _86756_/D sky130_fd_sc_hd__a21o_4
X_58217_ _63355_/A _58217_/B _58217_/Y sky130_fd_sc_hd__nand2_4
X_77051_ _77034_/B _77034_/C _77038_/X _77045_/X _77051_/X sky130_fd_sc_hd__and4_4
XPHY_430 sky130_fd_sc_hd__decap_3
X_43443_ _43422_/X _43426_/X _41596_/X _87417_/Q _43434_/X _43443_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74263_ _70134_/B _74003_/B _74262_/X _83115_/D sky130_fd_sc_hd__o21ai_4
X_55429_ _55429_/A _55429_/Y sky130_fd_sc_hd__inv_2
X_86249_ _83613_/CLK _50176_/Y _86249_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_441 sky130_fd_sc_hd__decap_3
X_40655_ _40577_/X _82869_/Q _40654_/X _40656_/A sky130_fd_sc_hd__o21a_4
X_59197_ _59135_/X _85649_/Q _59196_/X _59197_/X sky130_fd_sc_hd__o21a_4
X_71475_ _71068_/B _71827_/A sky130_fd_sc_hd__buf_2
XPHY_452 sky130_fd_sc_hd__decap_3
XPHY_463 sky130_fd_sc_hd__decap_3
X_76002_ _75999_/Y _76001_/Y _81741_/D sky130_fd_sc_hd__xor2_4
XPHY_474 sky130_fd_sc_hd__decap_3
X_73214_ _73359_/A _73214_/X sky130_fd_sc_hd__buf_2
X_46162_ _46162_/A _46162_/B _46162_/C _46162_/D _46162_/X sky130_fd_sc_hd__and4_4
X_70426_ _70426_/A _70442_/A sky130_fd_sc_hd__buf_2
X_58148_ _57677_/X _58145_/Y _58147_/Y _58148_/Y sky130_fd_sc_hd__a21oi_4
XPHY_485 sky130_fd_sc_hd__decap_3
X_43374_ _41397_/X _43371_/X _87454_/Q _43372_/X _43374_/X sky130_fd_sc_hd__a2bb2o_4
X_74194_ _74152_/A _66298_/B _74194_/X sky130_fd_sc_hd__and2_4
X_40586_ _40586_/A _40736_/A sky130_fd_sc_hd__buf_2
XPHY_496 sky130_fd_sc_hd__decap_3
X_45113_ _55855_/B _45056_/X _45087_/X _45113_/X sky130_fd_sc_hd__o21a_4
X_42325_ _42290_/A _42325_/X sky130_fd_sc_hd__buf_2
X_73145_ _83163_/Q _73079_/X _73144_/Y _73145_/X sky130_fd_sc_hd__a21o_4
X_58079_ _58696_/A _58079_/X sky130_fd_sc_hd__buf_2
X_70357_ _70356_/Y _70827_/C sky130_fd_sc_hd__buf_2
X_46093_ _80655_/Q _46121_/A sky130_fd_sc_hd__buf_2
X_60110_ _65607_/A _60110_/X sky130_fd_sc_hd__buf_2
X_49921_ _49919_/Y _49897_/X _49920_/X _49921_/Y sky130_fd_sc_hd__a21oi_4
X_45044_ _44895_/X _45044_/X sky130_fd_sc_hd__buf_2
X_42256_ _41454_/X _42248_/X _87956_/Q _42249_/X _87956_/D sky130_fd_sc_hd__a2bb2o_4
X_61090_ _61086_/X _72584_/C _60622_/D _61122_/B _61089_/Y _61091_/A
+ sky130_fd_sc_hd__a41o_4
X_73076_ _73074_/X _73075_/Y _72970_/X _73076_/Y sky130_fd_sc_hd__a21oi_4
X_77953_ _82251_/Q _81963_/Q _77954_/B sky130_fd_sc_hd__xnor2_4
X_70288_ _70269_/X _74722_/A _70287_/X _83810_/D sky130_fd_sc_hd__a21o_4
X_41207_ _41207_/A _41223_/B _41207_/X sky130_fd_sc_hd__or2_4
X_60041_ _60041_/A _60041_/Y sky130_fd_sc_hd__inv_2
X_72027_ _72017_/X _53852_/B _72027_/Y sky130_fd_sc_hd__nand2_4
X_76904_ _76904_/A _81597_/Q _76902_/B _76904_/Y sky130_fd_sc_hd__nand3_4
X_49852_ _49849_/Y _49844_/X _49851_/X _86312_/D sky130_fd_sc_hd__a21oi_4
X_42187_ _41272_/X _42183_/X _87990_/Q _42184_/X _42187_/X sky130_fd_sc_hd__a2bb2o_4
X_77884_ _77884_/A _77883_/Y _77887_/A sky130_fd_sc_hd__xor2_4
X_48803_ _48793_/A _48561_/B _48803_/Y sky130_fd_sc_hd__nand2_4
X_79623_ _79596_/Y _79621_/Y _79622_/Y _79624_/B sky130_fd_sc_hd__a21oi_4
X_41138_ _41136_/X _81148_/Q _41137_/X _41138_/X sky130_fd_sc_hd__o21a_4
X_76835_ _81493_/Q _76832_/Y _76834_/X _76835_/Y sky130_fd_sc_hd__o21ai_4
X_49783_ _49779_/A _49802_/B _49789_/C _52997_/D _49783_/X sky130_fd_sc_hd__and4_4
X_46995_ _46959_/A _52794_/B _46995_/Y sky130_fd_sc_hd__nand2_4
X_63800_ _63800_/A _63800_/B _63800_/C _63800_/Y sky130_fd_sc_hd__nor3_4
X_48734_ _48734_/A _48734_/X sky130_fd_sc_hd__buf_2
X_79554_ _79554_/A _79554_/B _79555_/C sky130_fd_sc_hd__nand2_4
X_45946_ _44207_/A _45947_/B sky130_fd_sc_hd__buf_2
X_41069_ _41061_/X _82281_/Q _41068_/X _41069_/Y sky130_fd_sc_hd__o21ai_4
X_64780_ _64680_/A _64780_/B _64780_/X sky130_fd_sc_hd__and2_4
X_76766_ _81695_/Q _76766_/B _76766_/Y sky130_fd_sc_hd__xnor2_4
X_61992_ _83248_/Q _63573_/A sky130_fd_sc_hd__inv_2
X_73978_ _73978_/A _73977_/X _73979_/B sky130_fd_sc_hd__nand2_4
X_78505_ _78501_/Y _78505_/B _78505_/C _78505_/X sky130_fd_sc_hd__or3_4
X_63731_ _62195_/A _64192_/B _64192_/C _63731_/D _63731_/Y sky130_fd_sc_hd__nand4_4
X_75717_ _75704_/B _75716_/X _75722_/A sky130_fd_sc_hd__nand2_4
X_48665_ _48652_/X _82342_/Q _48664_/Y _48666_/A sky130_fd_sc_hd__o21ai_4
X_60943_ _64067_/A _63781_/B sky130_fd_sc_hd__buf_2
X_72929_ _72929_/A _65519_/B _72929_/X sky130_fd_sc_hd__and2_4
X_79485_ _79484_/B _79484_/A _79470_/A _79470_/B _79486_/C sky130_fd_sc_hd__a211o_4
X_45877_ _45874_/X _45876_/Y _44972_/X _45877_/Y sky130_fd_sc_hd__a21oi_4
X_76697_ _76709_/B _76696_/X _76697_/Y sky130_fd_sc_hd__xnor2_4
X_47616_ _47616_/A _53151_/D sky130_fd_sc_hd__buf_2
X_66450_ _84121_/Q _66450_/Y sky130_fd_sc_hd__inv_2
X_78436_ _78418_/B _78418_/A _78435_/Y _78436_/Y sky130_fd_sc_hd__a21boi_4
X_44828_ _44827_/Y _86933_/D sky130_fd_sc_hd__inv_2
X_75648_ _81002_/Q _75648_/B _75648_/X sky130_fd_sc_hd__xor2_4
X_63662_ _63624_/X _63655_/X _63656_/X _63660_/X _63661_/Y _63662_/Y
+ sky130_fd_sc_hd__o41ai_4
X_48596_ _48904_/A _48959_/B sky130_fd_sc_hd__buf_2
X_60874_ _60865_/B _64172_/D sky130_fd_sc_hd__buf_2
X_65401_ _65401_/A _85826_/Q _65401_/X sky130_fd_sc_hd__and2_4
X_62613_ _61675_/B _62309_/B _62309_/C _62225_/X _62613_/Y sky130_fd_sc_hd__nand4_4
X_47547_ _47547_/A _47548_/A sky130_fd_sc_hd__inv_2
X_66381_ _65962_/X _65833_/B _65966_/X _66381_/Y sky130_fd_sc_hd__nand3_4
X_78367_ _78353_/B _78367_/Y sky130_fd_sc_hd__inv_2
X_44759_ _44740_/X _44741_/X _41316_/A _86969_/Q _44742_/X _44760_/A
+ sky130_fd_sc_hd__o32ai_4
X_63593_ _63589_/Y _63578_/X _63592_/Y _63593_/Y sky130_fd_sc_hd__a21oi_4
X_75579_ _81107_/Q _75579_/Y sky130_fd_sc_hd__inv_2
X_68120_ _68120_/A _68120_/X sky130_fd_sc_hd__buf_2
X_65332_ _65252_/X _83285_/Q _65230_/X _65331_/X _65332_/X sky130_fd_sc_hd__a211o_4
X_77318_ _77318_/A _77318_/B _77318_/Y sky130_fd_sc_hd__nand2_4
X_62544_ _62544_/A _62544_/Y sky130_fd_sc_hd__inv_2
X_47478_ _47619_/A _47478_/X sky130_fd_sc_hd__buf_2
X_78298_ _78298_/A _78298_/B _78299_/B sky130_fd_sc_hd__xor2_4
X_49217_ _49213_/Y _49214_/X _49216_/Y _49217_/Y sky130_fd_sc_hd__a21boi_4
X_68051_ _68403_/A _68051_/B _68051_/X sky130_fd_sc_hd__and2_4
X_46429_ _46422_/Y _46300_/X _46428_/X _46429_/Y sky130_fd_sc_hd__a21oi_4
X_65263_ _65782_/A _65289_/A sky130_fd_sc_hd__buf_2
X_77249_ _77249_/A _82084_/D _77250_/A sky130_fd_sc_hd__nor2_4
X_62475_ _62475_/A _62475_/X sky130_fd_sc_hd__buf_2
X_67002_ _66647_/A _67028_/A sky130_fd_sc_hd__buf_2
X_64214_ _64202_/Y _64210_/Y _64212_/Y _61323_/A _64213_/X _64214_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49148_ _49148_/A _49161_/B _49148_/Y sky130_fd_sc_hd__nor2_4
X_61426_ _61424_/X _61394_/X _61425_/Y _61426_/Y sky130_fd_sc_hd__a21oi_4
X_80260_ _80251_/A _80250_/X _80257_/Y _80261_/B sky130_fd_sc_hd__nand3_4
X_65194_ _65680_/A _65529_/A sky130_fd_sc_hd__buf_2
X_64145_ _63312_/B _64145_/B _64179_/C _64179_/D _64145_/Y sky130_fd_sc_hd__nand4_4
X_61357_ _61377_/A _61356_/X _61377_/C _61357_/Y sky130_fd_sc_hd__nand3_4
X_49079_ _49079_/A _53879_/B sky130_fd_sc_hd__buf_2
X_80191_ _80198_/B _80190_/X _80191_/Y sky130_fd_sc_hd__xnor2_4
X_51110_ _51115_/A _51115_/B _51110_/C _52801_/D _51110_/X sky130_fd_sc_hd__and4_4
X_60308_ _62737_/A _60309_/C sky130_fd_sc_hd__buf_2
X_52090_ _51922_/X _52100_/A sky130_fd_sc_hd__buf_2
X_68953_ _83954_/Q _68838_/X _68952_/X _83954_/D sky130_fd_sc_hd__a21bo_4
X_64076_ _60996_/Y _60934_/X _64184_/A _64184_/C _64076_/Y sky130_fd_sc_hd__a22oi_4
X_61288_ _61306_/A _72514_/A sky130_fd_sc_hd__inv_2
X_51041_ _51029_/A _51045_/B _51045_/C _52730_/D _51041_/X sky130_fd_sc_hd__and4_4
X_67904_ _87451_/Q _67834_/X _67835_/X _67903_/X _67904_/X sky130_fd_sc_hd__a211o_4
X_63027_ _60503_/X _63039_/A sky130_fd_sc_hd__buf_2
X_60239_ _60239_/A _60239_/B _60189_/A _60239_/X sky130_fd_sc_hd__and3_4
X_83950_ _81134_/CLK _83950_/D _80806_/D sky130_fd_sc_hd__dfxtp_4
X_68884_ _69088_/A _68884_/X sky130_fd_sc_hd__buf_2
X_82901_ _82896_/CLK _78218_/B _82901_/Q sky130_fd_sc_hd__dfxtp_4
X_67835_ _67359_/X _67835_/X sky130_fd_sc_hd__buf_2
X_83881_ _82558_/CLK _69980_/X _83881_/Q sky130_fd_sc_hd__dfxtp_4
X_54800_ _54790_/A _47543_/Y _54800_/Y sky130_fd_sc_hd__nand2_4
X_85620_ _86549_/CLK _53526_/Y _85620_/Q sky130_fd_sc_hd__dfxtp_4
X_82832_ _82833_/CLK _82832_/D _82800_/D sky130_fd_sc_hd__dfxtp_4
X_55780_ _45257_/A _55306_/X _55172_/X _55779_/X _55780_/X sky130_fd_sc_hd__a211o_4
X_67766_ _67763_/X _67765_/X _67742_/X _67766_/X sky130_fd_sc_hd__a21o_4
X_52992_ _85717_/Q _52984_/X _52991_/Y _52992_/Y sky130_fd_sc_hd__o21ai_4
X_64978_ _64975_/X _64977_/X _64574_/X _64978_/X sky130_fd_sc_hd__a21o_4
X_69505_ _69746_/A _69505_/X sky130_fd_sc_hd__buf_2
X_54731_ _54758_/A _54731_/X sky130_fd_sc_hd__buf_2
X_66717_ _66717_/A _66717_/X sky130_fd_sc_hd__buf_2
X_85551_ _86256_/CLK _53876_/Y _85551_/Q sky130_fd_sc_hd__dfxtp_4
X_51943_ _52322_/A _52177_/A sky130_fd_sc_hd__buf_2
X_63929_ _63849_/A _63960_/B sky130_fd_sc_hd__buf_2
X_82763_ _82769_/CLK _82763_/D _82955_/D sky130_fd_sc_hd__dfxtp_4
X_67697_ _87152_/Q _67670_/X _67671_/X _67696_/X _67698_/B sky130_fd_sc_hd__a211o_4
X_84502_ _84493_/CLK _61235_/Y _84502_/Q sky130_fd_sc_hd__dfxtp_4
X_81714_ _82053_/CLK _81714_/D _81714_/Q sky130_fd_sc_hd__dfxtp_4
X_57450_ _57188_/A _57445_/B _56818_/X _57450_/Y sky130_fd_sc_hd__nand3_4
X_69436_ _69423_/X _69340_/X _69434_/Y _69435_/Y _69436_/X sky130_fd_sc_hd__a211o_4
X_88270_ _88288_/CLK _41141_/Y _88270_/Q sky130_fd_sc_hd__dfxtp_4
X_54662_ _54667_/A _54674_/B _54644_/X _47302_/A _54662_/X sky130_fd_sc_hd__and4_4
X_66648_ _66669_/A _88144_/Q _66648_/X sky130_fd_sc_hd__and2_4
X_85482_ _84930_/CLK _54219_/Y _85482_/Q sky130_fd_sc_hd__dfxtp_4
X_51874_ _53269_/A _51875_/A sky130_fd_sc_hd__buf_2
X_82694_ _81190_/CLK _78845_/X _82694_/Q sky130_fd_sc_hd__dfxtp_4
X_56401_ _56397_/X _56399_/B _85208_/Q _56401_/Y sky130_fd_sc_hd__nand3_4
X_87221_ _87221_/CLK _87221_/D _69100_/B sky130_fd_sc_hd__dfxtp_4
X_53613_ _85602_/Q _53610_/X _53612_/Y _53613_/Y sky130_fd_sc_hd__o21ai_4
X_84433_ _81859_/CLK _62103_/Y _78056_/B sky130_fd_sc_hd__dfxtp_4
X_50825_ _51330_/A _50825_/B _50751_/C _50825_/X sky130_fd_sc_hd__and3_4
X_57381_ _56561_/X _57372_/X _56931_/X _45393_/A _57380_/X _85025_/D
+ sky130_fd_sc_hd__a32o_4
X_69367_ _69065_/X _69367_/X sky130_fd_sc_hd__buf_2
X_81645_ _81260_/CLK _81677_/Q _76300_/A sky130_fd_sc_hd__dfxtp_4
X_54593_ _54540_/A _54593_/X sky130_fd_sc_hd__buf_2
X_66579_ _69768_/A _66579_/X sky130_fd_sc_hd__buf_2
X_59120_ _59115_/X _59117_/Y _59118_/Y _59046_/X _59119_/X _59120_/X
+ sky130_fd_sc_hd__o32a_4
X_56332_ _56332_/A _56335_/B _55836_/B _56332_/Y sky130_fd_sc_hd__nand3_4
X_68318_ _68338_/A _68318_/X sky130_fd_sc_hd__buf_2
X_87152_ _88164_/CLK _87152_/D _87152_/Q sky130_fd_sc_hd__dfxtp_4
X_53544_ _53900_/A _53793_/A sky130_fd_sc_hd__buf_2
X_84364_ _84559_/CLK _62978_/Y _84364_/Q sky130_fd_sc_hd__dfxtp_4
X_50756_ _50754_/Y _50676_/X _50755_/X _50756_/Y sky130_fd_sc_hd__a21oi_4
X_81576_ _81575_/CLK _65817_/C _76706_/A sky130_fd_sc_hd__dfxtp_4
X_69298_ _81398_/D _69230_/X _69297_/X _83934_/D sky130_fd_sc_hd__a21bo_4
X_86103_ _82956_/CLK _50942_/Y _86103_/Q sky130_fd_sc_hd__dfxtp_4
X_59051_ _59013_/X _85757_/Q _59037_/X _59051_/X sky130_fd_sc_hd__o21a_4
X_83315_ _85003_/CLK _83315_/D _83315_/Q sky130_fd_sc_hd__dfxtp_4
X_56263_ _56263_/A _56263_/B _85254_/Q _56263_/Y sky130_fd_sc_hd__nand3_4
X_80527_ _80525_/X _80536_/B _80527_/Y sky130_fd_sc_hd__xnor2_4
X_68249_ _68246_/X _67532_/Y _68247_/X _68248_/Y _68249_/X sky130_fd_sc_hd__a211o_4
X_87083_ _87083_/CLK _44490_/Y _87083_/Q sky130_fd_sc_hd__dfxtp_4
X_53475_ _53469_/Y _53472_/X _53474_/X _85630_/D sky130_fd_sc_hd__a21oi_4
X_84295_ _84293_/CLK _84295_/D _63784_/C sky130_fd_sc_hd__dfxtp_4
X_50687_ _86153_/Q _50680_/X _50686_/Y _50687_/Y sky130_fd_sc_hd__o21ai_4
X_58002_ _58002_/A _58939_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_454_0_CLK clkbuf_9_227_0_CLK/X _85981_/CLK sky130_fd_sc_hd__clkbuf_1
X_55214_ _85026_/Q _55142_/A _80665_/Q _55213_/X _55214_/X sky130_fd_sc_hd__a211o_4
X_86034_ _85818_/CLK _51315_/Y _65002_/B sky130_fd_sc_hd__dfxtp_4
X_40440_ _40439_/X _40440_/X sky130_fd_sc_hd__buf_2
X_52426_ _50731_/A _51238_/B _53944_/C _52426_/Y sky130_fd_sc_hd__nor3_4
X_71260_ _71090_/A _71261_/B sky130_fd_sc_hd__buf_2
X_83246_ _83246_/CLK _83246_/D _62022_/A sky130_fd_sc_hd__dfxtp_4
X_56194_ _56186_/Y _56194_/X sky130_fd_sc_hd__buf_2
X_80458_ _80458_/A _80458_/B _80458_/X sky130_fd_sc_hd__or2_4
Xclkbuf_opt_27_CLK _86500_/CLK _85866_/CLK sky130_fd_sc_hd__clkbuf_16
X_70211_ _70209_/X _74763_/C _70210_/X _83836_/D sky130_fd_sc_hd__a21o_4
X_55145_ _55145_/A _55145_/B _55145_/Y sky130_fd_sc_hd__nor2_4
X_40371_ _40370_/X _40371_/X sky130_fd_sc_hd__buf_2
X_52357_ _52349_/A _49073_/X _52357_/Y sky130_fd_sc_hd__nand2_4
X_71191_ _71191_/A _71211_/A sky130_fd_sc_hd__inv_2
X_83177_ _83507_/CLK _83177_/D _83177_/Q sky130_fd_sc_hd__dfxtp_4
X_80389_ _80378_/X _80380_/B _80388_/Y _80406_/B sky130_fd_sc_hd__a21boi_4
X_42110_ _41050_/X _42103_/X _88031_/Q _42104_/X _88031_/D sky130_fd_sc_hd__a2bb2o_4
X_51308_ _51305_/Y _51289_/X _51307_/X _86035_/D sky130_fd_sc_hd__a21oi_4
X_70142_ _83528_/Q _83176_/Q _83510_/Q _83158_/Q _70144_/C sky130_fd_sc_hd__a22oi_4
X_82128_ _82084_/CLK _82128_/D _82084_/D sky130_fd_sc_hd__dfxtp_4
X_43090_ _43127_/A _43090_/X sky130_fd_sc_hd__buf_2
X_55076_ _55102_/A _55076_/X sky130_fd_sc_hd__buf_2
X_59953_ _59770_/A _60422_/A sky130_fd_sc_hd__buf_2
X_52288_ _64753_/B _52269_/X _52287_/Y _52288_/Y sky130_fd_sc_hd__o21ai_4
X_87985_ _87408_/CLK _87985_/D _87985_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_469_0_CLK clkbuf_9_234_0_CLK/X _85764_/CLK sky130_fd_sc_hd__clkbuf_1
X_42041_ _42041_/A _42041_/Y sky130_fd_sc_hd__inv_2
X_58904_ _58904_/A _58904_/X sky130_fd_sc_hd__buf_2
X_54027_ _54025_/Y _54015_/X _54026_/X _54027_/Y sky130_fd_sc_hd__a21oi_4
X_51239_ _51236_/Y _51237_/X _51238_/Y _51239_/Y sky130_fd_sc_hd__a21oi_4
X_74950_ _81137_/D _80849_/Q _74958_/B sky130_fd_sc_hd__or2_4
X_70073_ _82537_/D _70067_/X _70072_/X _83857_/D sky130_fd_sc_hd__a21bo_4
X_86936_ _86935_/CLK _86936_/D _86936_/Q sky130_fd_sc_hd__dfxtp_4
X_82059_ _84105_/CLK _82059_/D _82059_/Q sky130_fd_sc_hd__dfxtp_4
X_59884_ _59883_/Y _59884_/X sky130_fd_sc_hd__buf_2
X_73901_ _73949_/A _73901_/B _73901_/X sky130_fd_sc_hd__and2_4
X_58835_ _59033_/A _58835_/X sky130_fd_sc_hd__buf_2
X_74881_ _81127_/D _74875_/B _74881_/Y sky130_fd_sc_hd__nand2_4
X_86867_ _84409_/CLK _45594_/Y _63147_/B sky130_fd_sc_hd__dfxtp_4
X_45800_ _82983_/Q _74691_/B sky130_fd_sc_hd__inv_2
X_76620_ _76620_/A _81548_/Q _76620_/X sky130_fd_sc_hd__xor2_4
X_73832_ _73828_/X _73831_/X _73738_/X _73835_/A sky130_fd_sc_hd__a21o_4
X_85818_ _85818_/CLK _85818_/D _85818_/Q sky130_fd_sc_hd__dfxtp_4
X_46780_ _46806_/A _50976_/B _46780_/Y sky130_fd_sc_hd__nand2_4
X_58766_ _58766_/A _58766_/X sky130_fd_sc_hd__buf_2
X_55978_ _55695_/A _56469_/C _55978_/X sky130_fd_sc_hd__and2_4
X_43992_ _43990_/Y _43954_/X _43991_/Y _43992_/Y sky130_fd_sc_hd__a21oi_4
X_86798_ _87484_/CLK _86798_/D _66765_/B sky130_fd_sc_hd__dfxtp_4
X_57717_ _58882_/A _57718_/A sky130_fd_sc_hd__buf_2
X_45731_ _45668_/X _61582_/A _45685_/X _45731_/Y sky130_fd_sc_hd__o21ai_4
X_76551_ _76552_/A _81545_/Q _76554_/B sky130_fd_sc_hd__nor2_4
X_42943_ _41782_/X _42930_/X _68018_/B _42931_/X _87638_/D sky130_fd_sc_hd__a2bb2o_4
X_54929_ _54925_/Y _54909_/X _54928_/X _85352_/D sky130_fd_sc_hd__a21oi_4
X_73763_ _73665_/X _84985_/Q _73740_/X _73762_/X _73764_/B sky130_fd_sc_hd__a211o_4
X_85749_ _85751_/CLK _52819_/Y _85749_/Q sky130_fd_sc_hd__dfxtp_4
X_70975_ _46396_/B _70961_/A _70974_/Y _83644_/D sky130_fd_sc_hd__o21ai_4
X_58697_ _58697_/A _58698_/A sky130_fd_sc_hd__buf_2
X_75502_ _75503_/A _75503_/C _75503_/B _75536_/A sky130_fd_sc_hd__a21o_4
X_48450_ _48372_/X _47926_/A _48449_/Y _74406_/A sky130_fd_sc_hd__o21ai_4
X_72714_ _72714_/A _72714_/B _55656_/X _72714_/Y sky130_fd_sc_hd__nand3_4
X_79270_ _79257_/Y _79270_/B _79270_/X sky130_fd_sc_hd__or2_4
X_45662_ _57414_/A _45357_/X _45339_/X _45662_/X sky130_fd_sc_hd__o21a_4
X_57648_ _50391_/A _46620_/A _46428_/C _57648_/Y sky130_fd_sc_hd__nand3_4
X_76482_ _76482_/A _76482_/B _76482_/C _76463_/X _76482_/X sky130_fd_sc_hd__and4_4
X_42874_ _42846_/X _42874_/X sky130_fd_sc_hd__buf_2
X_73694_ _73692_/X _73694_/B _73694_/C _73694_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_407_0_CLK clkbuf_9_203_0_CLK/X _85338_/CLK sky130_fd_sc_hd__clkbuf_1
X_47401_ _47397_/Y _47364_/X _47400_/X _86639_/D sky130_fd_sc_hd__a21oi_4
X_78221_ _78210_/B _78221_/B _78221_/Y sky130_fd_sc_hd__nand2_4
X_44613_ _44588_/X _44589_/X _40972_/A _87032_/Q _44590_/X _44613_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75433_ _75431_/X _75432_/Y _75433_/X sky130_fd_sc_hd__and2_4
X_41825_ _41825_/A _41825_/X sky130_fd_sc_hd__buf_2
X_87419_ _81182_/CLK _87419_/D _87419_/Q sky130_fd_sc_hd__dfxtp_4
X_48381_ _48392_/A _48380_/X _48381_/Y sky130_fd_sc_hd__nand2_4
X_72645_ _72630_/X _72645_/X sky130_fd_sc_hd__buf_2
X_57579_ _84975_/Q _57550_/X _57578_/Y _57579_/Y sky130_fd_sc_hd__o21ai_4
X_45593_ _45591_/X _61483_/A _45530_/X _45593_/Y sky130_fd_sc_hd__o21ai_4
X_88399_ _86834_/CLK _40392_/X _88399_/Q sky130_fd_sc_hd__dfxtp_4
X_59318_ _59253_/X _59316_/Y _59317_/Y _59271_/X _59258_/X _59318_/X
+ sky130_fd_sc_hd__o32a_4
X_47332_ _47382_/A _47332_/X sky130_fd_sc_hd__buf_2
X_78152_ _78152_/A _78151_/Y _78153_/B sky130_fd_sc_hd__xor2_4
X_44544_ _44529_/X _44530_/X _40820_/A _44543_/Y _44533_/X _87060_/D
+ sky130_fd_sc_hd__o32ai_4
X_75364_ _75364_/A _75355_/X _75364_/Y sky130_fd_sc_hd__nor2_4
X_41756_ _41603_/X _82889_/Q _41755_/X _41756_/X sky130_fd_sc_hd__o21a_4
X_60590_ _63252_/B _60570_/C _63272_/A _60590_/Y sky130_fd_sc_hd__a21oi_4
X_72576_ _72576_/A _72576_/Y sky130_fd_sc_hd__inv_2
X_77103_ _82096_/Q _77103_/B _77103_/X sky130_fd_sc_hd__xor2_4
X_74315_ _72704_/A _74325_/A sky130_fd_sc_hd__buf_2
X_40707_ _40707_/A _40707_/X sky130_fd_sc_hd__buf_2
X_47263_ _81821_/Q _47264_/A sky130_fd_sc_hd__inv_2
X_59249_ _59199_/X _85741_/Q _59124_/X _59249_/X sky130_fd_sc_hd__o21a_4
X_71527_ _70933_/B _70694_/A _70700_/A _71527_/Y sky130_fd_sc_hd__nand3_4
X_78083_ _78083_/A _78083_/B _78085_/A sky130_fd_sc_hd__nand2_4
X_44475_ _44603_/A _44475_/X sky130_fd_sc_hd__buf_2
X_75295_ _75284_/A _75283_/Y _75276_/Y _75295_/X sky130_fd_sc_hd__o21a_4
X_41687_ _41603_/X _82903_/Q _41686_/X _41687_/X sky130_fd_sc_hd__o21a_4
X_49002_ _49002_/A _49052_/A sky130_fd_sc_hd__buf_2
X_46214_ _46213_/X _46098_/A _46214_/C _46214_/D _46215_/C sky130_fd_sc_hd__nand4_4
Xclkbuf_8_81_0_CLK clkbuf_8_81_0_CLK/A clkbuf_8_81_0_CLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_260 sky130_fd_sc_hd__decap_3
X_77034_ _77026_/Y _77034_/B _77034_/C _77041_/A sky130_fd_sc_hd__nand3_4
X_43426_ _43425_/X _43426_/X sky130_fd_sc_hd__buf_2
X_62260_ _61367_/A _62247_/X _62259_/X _62560_/D _62260_/Y sky130_fd_sc_hd__nand4_4
X_74246_ _87317_/Q _74246_/B _74246_/Y sky130_fd_sc_hd__nor2_4
XPHY_271 sky130_fd_sc_hd__decap_3
X_40638_ _40836_/A _40638_/X sky130_fd_sc_hd__buf_2
X_47194_ _47194_/A _47195_/A sky130_fd_sc_hd__inv_2
X_71458_ _70689_/A _71446_/X _71458_/C _71458_/Y sky130_fd_sc_hd__nor3_4
XPHY_282 sky130_fd_sc_hd__decap_3
XPHY_293 sky130_fd_sc_hd__decap_3
Xclkbuf_opt_18_CLK _83613_/CLK _86453_/CLK sky130_fd_sc_hd__clkbuf_16
X_61211_ _64457_/B _61238_/C sky130_fd_sc_hd__buf_2
X_70409_ MACRO_WR_SELECT _70609_/A sky130_fd_sc_hd__buf_2
X_46145_ _58547_/A _46150_/B sky130_fd_sc_hd__buf_2
X_43357_ _43302_/A _43357_/X sky130_fd_sc_hd__buf_2
X_62191_ _62181_/A _62181_/B _78049_/B _62191_/Y sky130_fd_sc_hd__nor3_4
X_74177_ _74237_/A _74177_/B _74177_/X sky130_fd_sc_hd__and2_4
X_40569_ _40550_/X _40556_/X _40560_/X _88371_/Q _40568_/X _40569_/Y
+ sky130_fd_sc_hd__o32ai_4
X_71389_ _71411_/A _71386_/B _71399_/C _71389_/Y sky130_fd_sc_hd__nor3_4
X_42308_ _42307_/X _42297_/X _41596_/X _87929_/Q _42298_/X _42308_/Y
+ sky130_fd_sc_hd__o32ai_4
X_61142_ _64323_/A _64250_/C sky130_fd_sc_hd__buf_2
X_73128_ _73125_/X _73127_/X _72951_/X _73128_/X sky130_fd_sc_hd__a21o_4
X_46076_ _41600_/Y _43586_/X _67227_/B _43593_/X _86779_/D sky130_fd_sc_hd__a2bb2o_4
X_43288_ _43218_/A _43288_/X sky130_fd_sc_hd__buf_2
X_78985_ _78998_/A _78998_/B _78993_/A sky130_fd_sc_hd__xor2_4
Xclkbuf_8_96_0_CLK clkbuf_8_97_0_CLK/A clkbuf_8_96_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_49904_ _49904_/A _49893_/B _49904_/C _53118_/D _49904_/X sky130_fd_sc_hd__and4_4
X_45027_ _45827_/B _45027_/X sky130_fd_sc_hd__buf_2
X_65950_ _65768_/A _65950_/X sky130_fd_sc_hd__buf_2
X_42239_ _42239_/A _87965_/D sky130_fd_sc_hd__inv_2
X_77936_ _82249_/Q _81961_/Q _77946_/A sky130_fd_sc_hd__xnor2_4
X_61073_ _61070_/X _61122_/C _61074_/A sky130_fd_sc_hd__and2_4
X_73059_ _72732_/B _73059_/X sky130_fd_sc_hd__buf_2
X_64901_ _64897_/X _64712_/B _64900_/X _64901_/Y sky130_fd_sc_hd__nand3_4
X_60024_ _62218_/A _62194_/D sky130_fd_sc_hd__buf_2
X_49835_ _49830_/A _49851_/B _49830_/C _53048_/D _49835_/X sky130_fd_sc_hd__and4_4
X_65881_ _65875_/X _65879_/X _65880_/X _65884_/A sky130_fd_sc_hd__a21o_4
X_77867_ _77855_/Y _77860_/B _77861_/A _77867_/Y sky130_fd_sc_hd__a21boi_4
X_67620_ _67614_/X _67617_/X _67619_/X _67623_/A sky130_fd_sc_hd__a21o_4
X_79606_ _79602_/X _79603_/Y _79607_/B sky130_fd_sc_hd__nand2_4
X_64832_ _64827_/X _64831_/X _64729_/X _64832_/X sky130_fd_sc_hd__a21o_4
X_76818_ _76818_/A _76818_/B _76819_/B sky130_fd_sc_hd__xor2_4
X_49766_ _49779_/A _49750_/X _49789_/C _52982_/D _49766_/X sky130_fd_sc_hd__and4_4
X_46978_ _59068_/A _46955_/X _46977_/Y _46978_/Y sky130_fd_sc_hd__o21ai_4
X_77798_ _77796_/Y _77798_/B _77798_/Y sky130_fd_sc_hd__nand2_4
X_48717_ _48725_/A _48368_/X _48717_/Y sky130_fd_sc_hd__nand2_4
X_67551_ _67550_/X _67551_/X sky130_fd_sc_hd__buf_2
X_79537_ _64542_/Y _79538_/A _79544_/A sky130_fd_sc_hd__nand2_4
X_45929_ _72745_/A _72905_/A sky130_fd_sc_hd__buf_2
X_64763_ _84228_/Q _64764_/C sky130_fd_sc_hd__inv_2
X_76749_ _76735_/Y _76749_/Y sky130_fd_sc_hd__inv_2
X_49697_ _49685_/A _49697_/B _49685_/C _51220_/D _49697_/X sky130_fd_sc_hd__and4_4
X_61975_ _61722_/A _62002_/A sky130_fd_sc_hd__buf_2
X_66502_ _66500_/Y _66483_/X _66501_/X _66502_/X sky130_fd_sc_hd__a21o_4
X_63714_ _59448_/A _63370_/A _63714_/Y sky130_fd_sc_hd__nor2_4
X_48648_ _48647_/Y _48847_/B sky130_fd_sc_hd__buf_2
X_60926_ _60853_/X _60926_/X sky130_fd_sc_hd__buf_2
X_67482_ _67575_/A _67482_/B _67482_/X sky130_fd_sc_hd__and2_4
X_79468_ _79466_/X _79468_/B _79484_/B sky130_fd_sc_hd__xnor2_4
X_64694_ _64694_/A _64694_/B _64694_/X sky130_fd_sc_hd__and2_4
Xclkbuf_8_34_0_CLK clkbuf_8_35_0_CLK/A clkbuf_9_69_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_69221_ _87533_/Q _69044_/X _68979_/X _69220_/X _69221_/X sky130_fd_sc_hd__a211o_4
X_66433_ _66433_/A _66419_/X _66433_/C _66433_/X sky130_fd_sc_hd__and3_4
X_78419_ _78418_/B _78418_/A _78423_/C sky130_fd_sc_hd__nand2_4
X_63645_ _63468_/A _63670_/B sky130_fd_sc_hd__buf_2
X_60857_ _60851_/X _60408_/A _59753_/B _60857_/D _60857_/X sky130_fd_sc_hd__and4_4
X_48579_ _52199_/A _48624_/B _48610_/C _48579_/X sky130_fd_sc_hd__and3_4
X_79399_ _79387_/A _79386_/Y _79398_/X _79399_/X sky130_fd_sc_hd__a21o_4
X_50610_ _48979_/A _50560_/X _50568_/C _50610_/X sky130_fd_sc_hd__and3_4
X_81430_ _84049_/CLK _81462_/Q _76062_/B sky130_fd_sc_hd__dfxtp_4
X_69152_ _69148_/X _69151_/X _69116_/X _69152_/X sky130_fd_sc_hd__a21o_4
X_66364_ _66318_/X _66415_/B _66364_/C _66364_/X sky130_fd_sc_hd__and3_4
X_51590_ _51590_/A _53115_/B _51590_/Y sky130_fd_sc_hd__nand2_4
X_63576_ _63556_/X _63569_/X _63570_/X _63574_/X _63575_/Y _63576_/Y
+ sky130_fd_sc_hd__o41ai_4
X_60788_ _60558_/X _60792_/A sky130_fd_sc_hd__buf_2
X_68103_ _68097_/X _66650_/Y _68089_/X _68102_/Y _68103_/X sky130_fd_sc_hd__a211o_4
X_65315_ _65836_/A _65315_/B _65315_/X sky130_fd_sc_hd__and2_4
X_50541_ _50541_/A _48673_/B _50541_/Y sky130_fd_sc_hd__nand2_4
X_62527_ _62483_/X _62541_/B _62527_/C _62527_/Y sky130_fd_sc_hd__nor3_4
X_81361_ _81361_/CLK _81361_/D _81361_/Q sky130_fd_sc_hd__dfxtp_4
X_69083_ _69080_/X _69082_/X _69017_/X _69083_/Y sky130_fd_sc_hd__a21oi_4
X_66295_ _66180_/A _66295_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_49_0_CLK clkbuf_8_49_0_CLK/A clkbuf_9_99_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_83100_ _83846_/CLK _83100_/D _70304_/C sky130_fd_sc_hd__dfxtp_4
X_80312_ _84749_/Q _66319_/C _80313_/A sky130_fd_sc_hd__nor2_4
X_68034_ _68029_/X _68032_/X _68033_/X _68034_/X sky130_fd_sc_hd__a21o_4
X_53260_ _85666_/Q _51929_/X _53259_/Y _53260_/Y sky130_fd_sc_hd__o21ai_4
X_65246_ _65243_/Y _65195_/X _65245_/X _65246_/X sky130_fd_sc_hd__a21o_4
X_84080_ _84079_/CLK _84080_/D _84080_/Q sky130_fd_sc_hd__dfxtp_4
X_50472_ _86194_/Q _50387_/X _50471_/Y _50472_/Y sky130_fd_sc_hd__o21ai_4
X_81292_ _81620_/CLK _76980_/X _81260_/D sky130_fd_sc_hd__dfxtp_4
X_62458_ _61542_/A _62472_/B _62490_/C _62431_/D _62458_/Y sky130_fd_sc_hd__nand4_4
X_52211_ _85867_/Q _52178_/X _52210_/Y _52211_/Y sky130_fd_sc_hd__o21ai_4
X_83031_ _85269_/CLK _83031_/D _83031_/Q sky130_fd_sc_hd__dfxtp_4
X_61409_ _64282_/A _61452_/B _61452_/C _61391_/D _61409_/Y sky130_fd_sc_hd__nand4_4
X_80243_ _80239_/Y _80242_/Y _80243_/X sky130_fd_sc_hd__xor2_4
X_53191_ _53211_/A _53181_/B _53169_/X _53191_/D _53191_/X sky130_fd_sc_hd__and4_4
X_65177_ _65174_/X _65176_/X _65161_/X _65177_/X sky130_fd_sc_hd__a21o_4
X_62389_ _62406_/A _62389_/B _62387_/Y _62389_/D _62389_/Y sky130_fd_sc_hd__nand4_4
X_52142_ _52138_/Y _52108_/X _52141_/X _85881_/D sky130_fd_sc_hd__a21oi_4
X_64128_ _64124_/X _64048_/X _64125_/Y _64126_/Y _64127_/X _64128_/X
+ sky130_fd_sc_hd__a41o_4
X_80174_ _84946_/Q _65546_/C _80176_/A sky130_fd_sc_hd__xor2_4
X_69985_ _68420_/X _68423_/X _69925_/X _69985_/Y sky130_fd_sc_hd__a21oi_4
X_52073_ _52071_/Y _52066_/X _52072_/Y _85894_/D sky130_fd_sc_hd__a21boi_4
X_56950_ _56949_/X _56589_/X _85116_/Q _56947_/X _85116_/D sky130_fd_sc_hd__a2bb2o_4
X_64059_ _84837_/Q _64091_/B _64091_/C _64091_/D _64059_/Y sky130_fd_sc_hd__nand4_4
X_87770_ _87525_/CLK _87770_/D _69480_/B sky130_fd_sc_hd__dfxtp_4
X_68936_ _74095_/A _68792_/X _68933_/X _68935_/Y _68936_/X sky130_fd_sc_hd__a211o_4
X_84982_ _86587_/CLK _57545_/Y _84982_/Q sky130_fd_sc_hd__dfxtp_4
X_51024_ _51018_/A _51029_/B _51029_/C _52716_/D _51024_/X sky130_fd_sc_hd__and4_4
X_55901_ _83031_/Q _55607_/A _44101_/A _55900_/X _55901_/X sky130_fd_sc_hd__a211o_4
X_86721_ _85471_/CLK _46621_/Y _86721_/Q sky130_fd_sc_hd__dfxtp_4
X_83933_ _83933_/CLK _69314_/X _83933_/Q sky130_fd_sc_hd__dfxtp_4
X_56881_ _55674_/A _46234_/Y _56881_/X sky130_fd_sc_hd__and2_4
X_68867_ _68863_/X _68866_/X _68846_/X _68867_/Y sky130_fd_sc_hd__a21oi_4
X_58620_ _58618_/X _86109_/Q _58619_/X _58620_/Y sky130_fd_sc_hd__o21ai_4
X_55832_ _85265_/Q _55475_/X _44048_/X _55831_/X _55832_/X sky130_fd_sc_hd__a211o_4
X_67818_ _67817_/X _87647_/Q _67818_/X sky130_fd_sc_hd__and2_4
X_86652_ _86651_/CLK _47276_/Y _86652_/Q sky130_fd_sc_hd__dfxtp_4
X_83864_ _82541_/CLK _70047_/X _82544_/D sky130_fd_sc_hd__dfxtp_4
X_68798_ _68795_/X _68798_/B _68798_/Y sky130_fd_sc_hd__nand2_4
X_85603_ _85599_/CLK _85603_/D _85603_/Q sky130_fd_sc_hd__dfxtp_4
X_82815_ _82152_/CLK _82847_/Q _78749_/A sky130_fd_sc_hd__dfxtp_4
X_58551_ _58551_/A _58557_/B _58551_/Y sky130_fd_sc_hd__nand2_4
X_55763_ _55760_/Y _44095_/X _55762_/X _56117_/C sky130_fd_sc_hd__a21boi_4
X_67749_ _67793_/A _87714_/Q _67749_/X sky130_fd_sc_hd__and2_4
X_86583_ _86554_/CLK _47947_/Y _66055_/B sky130_fd_sc_hd__dfxtp_4
X_52975_ _52892_/A _52975_/X sky130_fd_sc_hd__buf_2
X_83795_ _83819_/CLK _70329_/X _74742_/B sky130_fd_sc_hd__dfxtp_4
X_57502_ _57500_/Y _46576_/X _57501_/Y _84991_/D sky130_fd_sc_hd__a21boi_4
X_88322_ _88060_/CLK _88322_/D _88322_/Q sky130_fd_sc_hd__dfxtp_4
X_54714_ _54718_/A _47394_/Y _54714_/Y sky130_fd_sc_hd__nand2_4
X_85534_ _85535_/CLK _85534_/D _85534_/Q sky130_fd_sc_hd__dfxtp_4
X_51926_ _51926_/A _85921_/D sky130_fd_sc_hd__inv_2
X_70760_ _70698_/A _70760_/B _70761_/A sky130_fd_sc_hd__nor2_4
X_58482_ _58510_/A _58502_/B sky130_fd_sc_hd__buf_2
X_82746_ _82746_/CLK _79435_/B _82746_/Q sky130_fd_sc_hd__dfxtp_4
X_55694_ _55691_/A _55695_/A sky130_fd_sc_hd__buf_2
X_57433_ _57484_/A _57431_/Y _57432_/Y _57434_/A sky130_fd_sc_hd__a21o_4
X_69419_ _68874_/X _68877_/X _69418_/X _69419_/Y sky130_fd_sc_hd__a21oi_4
X_88253_ _87103_/CLK _88253_/D _68924_/B sky130_fd_sc_hd__dfxtp_4
X_54645_ _54667_/A _54645_/B _54644_/X _54645_/D _54645_/X sky130_fd_sc_hd__and4_4
X_85465_ _82768_/CLK _85465_/D _85465_/Q sky130_fd_sc_hd__dfxtp_4
X_51857_ _51853_/A _46805_/X _51857_/Y sky130_fd_sc_hd__nand2_4
X_70691_ _70570_/Y _70692_/A sky130_fd_sc_hd__buf_2
X_82677_ _82671_/CLK _82677_/D _82677_/Q sky130_fd_sc_hd__dfxtp_4
X_87204_ _87150_/CLK _43910_/X _87204_/Q sky130_fd_sc_hd__dfxtp_4
X_41610_ _41610_/A _41610_/Y sky130_fd_sc_hd__inv_2
X_72430_ _64758_/X _85319_/Q _72386_/X _72430_/X sky130_fd_sc_hd__o21a_4
X_84416_ _84403_/CLK _84416_/D _84416_/Q sky130_fd_sc_hd__dfxtp_4
X_50808_ _50787_/X _50808_/B _50808_/Y sky130_fd_sc_hd__nand2_4
X_57364_ _57222_/Y _56275_/X _73191_/B _57364_/D _57364_/X sky130_fd_sc_hd__and4_4
X_81628_ _81275_/CLK _76548_/X _81628_/Q sky130_fd_sc_hd__dfxtp_4
X_88184_ _87110_/CLK _88184_/D _67231_/B sky130_fd_sc_hd__dfxtp_4
X_42590_ _42590_/A _42590_/X sky130_fd_sc_hd__buf_2
X_54576_ _54565_/A _54585_/B _54565_/C _54576_/D _54576_/X sky130_fd_sc_hd__and4_4
X_85396_ _85492_/CLK _54690_/Y _85396_/Q sky130_fd_sc_hd__dfxtp_4
X_51788_ _51785_/Y _51767_/X _51787_/X _85946_/D sky130_fd_sc_hd__a21oi_4
X_59103_ _58934_/X _85656_/Q _59081_/X _59103_/X sky130_fd_sc_hd__o21a_4
X_56315_ _56309_/A _56312_/X _85239_/Q _56315_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_393_0_CLK clkbuf_9_196_0_CLK/X _84477_/CLK sky130_fd_sc_hd__clkbuf_1
X_41541_ _41490_/A _41541_/X sky130_fd_sc_hd__buf_2
X_87135_ _87484_/CLK _44388_/X _87135_/Q sky130_fd_sc_hd__dfxtp_4
X_53527_ _53509_/A _47978_/A _53527_/Y sky130_fd_sc_hd__nand2_4
X_72361_ _72155_/A _72361_/X sky130_fd_sc_hd__buf_2
X_84347_ _82263_/CLK _84347_/D _79363_/A sky130_fd_sc_hd__dfxtp_4
X_50739_ _86143_/Q _50706_/X _50738_/Y _50739_/Y sky130_fd_sc_hd__o21ai_4
X_57295_ _57295_/A _57295_/B _57295_/Y sky130_fd_sc_hd__nand2_4
X_81559_ _84049_/CLK _76845_/X _81515_/D sky130_fd_sc_hd__dfxtp_4
X_74100_ _88348_/Q _73153_/X _72901_/X _74100_/Y sky130_fd_sc_hd__o21ai_4
X_71312_ _50341_/B _71289_/Y _71311_/Y _83540_/D sky130_fd_sc_hd__o21ai_4
X_59034_ _58961_/X _85662_/Q _59010_/X _59034_/X sky130_fd_sc_hd__o21a_4
X_44260_ _44175_/A _64642_/A sky130_fd_sc_hd__buf_2
X_56246_ _56250_/A _56253_/B _56246_/C _56246_/Y sky130_fd_sc_hd__nand3_4
X_75080_ _81058_/Q _75080_/B _81026_/D sky130_fd_sc_hd__xor2_4
X_87066_ _87070_/CLK _87066_/D _87066_/Q sky130_fd_sc_hd__dfxtp_4
X_41472_ _41421_/X _82334_/Q _41471_/X _41472_/X sky130_fd_sc_hd__o21a_4
X_53458_ _53458_/A _48178_/X _53458_/Y sky130_fd_sc_hd__nand2_4
X_72292_ _59297_/A _72292_/X sky130_fd_sc_hd__buf_2
X_84278_ _84273_/CLK _64056_/Y _80049_/B sky130_fd_sc_hd__dfxtp_4
X_43211_ _43024_/A _43212_/A sky130_fd_sc_hd__buf_2
X_74031_ _74031_/A _73869_/X _74031_/Y sky130_fd_sc_hd__nor2_4
X_86017_ _83690_/CLK _51401_/Y _86017_/Q sky130_fd_sc_hd__dfxtp_4
X_40423_ _40947_/A _40907_/B sky130_fd_sc_hd__buf_2
X_52409_ _52400_/X _50712_/B _52409_/Y sky130_fd_sc_hd__nand2_4
X_71243_ _71252_/A _71217_/B _71248_/C _71243_/Y sky130_fd_sc_hd__nand3_4
X_83229_ _83229_/CLK _72578_/X _79385_/B sky130_fd_sc_hd__dfxtp_4
X_44191_ _44131_/A _72739_/A sky130_fd_sc_hd__buf_2
X_56177_ _56177_/A _56177_/B _55741_/B _56178_/B sky130_fd_sc_hd__nand3_4
X_53389_ _53387_/Y _53382_/X _53388_/X _85643_/D sky130_fd_sc_hd__a21oi_4
X_55128_ _55128_/A _55128_/X sky130_fd_sc_hd__buf_2
X_43142_ _43127_/A _43142_/X sky130_fd_sc_hd__buf_2
X_40354_ _40353_/Y _40354_/X sky130_fd_sc_hd__buf_2
X_71174_ _48763_/B _71165_/X _71173_/Y _71174_/Y sky130_fd_sc_hd__o21ai_4
X_70125_ _70125_/A _70122_/Y _70125_/C _70125_/D _70125_/Y sky130_fd_sc_hd__nand4_4
X_47950_ _83774_/Q _53514_/B sky130_fd_sc_hd__inv_2
X_43073_ _43072_/X _43050_/X _40682_/X _87586_/Q _43061_/X _43073_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55059_ _55054_/A _54894_/B _55059_/Y sky130_fd_sc_hd__nand2_4
X_59936_ _59935_/X _59936_/X sky130_fd_sc_hd__buf_2
X_78770_ _78770_/A _78770_/B _78737_/Y _78770_/D _78771_/A sky130_fd_sc_hd__and4_4
X_75982_ _81514_/Q _75982_/B _75982_/X sky130_fd_sc_hd__xor2_4
X_87968_ _87210_/CLK _87968_/D _87968_/Q sky130_fd_sc_hd__dfxtp_4
X_46901_ _58953_/A _46859_/X _46900_/Y _46901_/Y sky130_fd_sc_hd__o21ai_4
X_42024_ _42024_/A _42024_/X sky130_fd_sc_hd__buf_2
X_77721_ _77721_/A _77722_/B sky130_fd_sc_hd__inv_2
Xclkbuf_10_331_0_CLK clkbuf_9_165_0_CLK/X _86005_/CLK sky130_fd_sc_hd__clkbuf_1
X_74933_ _74930_/Y _74932_/X _74933_/Y sky130_fd_sc_hd__nand2_4
X_70056_ _70056_/A _70056_/X sky130_fd_sc_hd__buf_2
X_86919_ _87141_/CLK _86919_/D _67915_/B sky130_fd_sc_hd__dfxtp_4
X_47881_ _47880_/Y _51954_/B sky130_fd_sc_hd__buf_2
X_59867_ _57757_/A _63130_/A sky130_fd_sc_hd__buf_2
X_87899_ _87898_/CLK _87899_/D _87899_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_961_0_CLK clkbuf_9_480_0_CLK/X _86558_/CLK sky130_fd_sc_hd__clkbuf_1
X_49620_ _49618_/Y _49596_/X _49619_/X _86354_/D sky130_fd_sc_hd__a21oi_4
X_46832_ _83666_/Q _52700_/B sky130_fd_sc_hd__inv_2
X_58818_ _58699_/A _86381_/Q _58818_/Y sky130_fd_sc_hd__nor2_4
X_77652_ _77652_/A _82110_/D _77652_/Y sky130_fd_sc_hd__nor2_4
X_74864_ _81125_/D _74870_/B _74867_/A sky130_fd_sc_hd__xnor2_4
X_59798_ _59754_/C _59634_/A _59634_/B _59662_/B _59691_/X _59798_/Y
+ sky130_fd_sc_hd__a41oi_4
X_76603_ _76614_/B _76602_/Y _76603_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_452_0_CLK clkbuf_8_226_0_CLK/X clkbuf_9_452_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_49551_ _49496_/A _49551_/X sky130_fd_sc_hd__buf_2
X_73815_ _73813_/X _73815_/B _73815_/C _73815_/Y sky130_fd_sc_hd__nand3_4
X_46763_ _54353_/D _52661_/D sky130_fd_sc_hd__buf_2
X_58749_ _58749_/A _58763_/A sky130_fd_sc_hd__buf_2
X_77583_ _77583_/A _77584_/C sky130_fd_sc_hd__inv_2
X_43975_ _80667_/Q _43975_/B _43975_/Y sky130_fd_sc_hd__nor2_4
X_74795_ _74795_/A _74804_/C _74744_/X _74769_/D _74798_/B sky130_fd_sc_hd__nand4_4
Xclkbuf_10_346_0_CLK clkbuf_9_173_0_CLK/X _86353_/CLK sky130_fd_sc_hd__clkbuf_1
X_48502_ _48494_/Y _48459_/X _48501_/X _86517_/D sky130_fd_sc_hd__a21oi_4
X_79322_ _79320_/X _79322_/B _79322_/Y sky130_fd_sc_hd__xnor2_4
X_45714_ _45714_/A _45714_/X sky130_fd_sc_hd__buf_2
X_76534_ _76533_/Y _76534_/Y sky130_fd_sc_hd__inv_2
X_42926_ _41731_/X _42920_/X _87648_/Q _42922_/X _87648_/D sky130_fd_sc_hd__a2bb2o_4
X_61760_ _61842_/A _61795_/B sky130_fd_sc_hd__buf_2
X_49482_ _86379_/Q _49470_/X _49481_/Y _49482_/Y sky130_fd_sc_hd__o21ai_4
X_73746_ _73727_/X _73730_/X _73745_/X _73746_/X sky130_fd_sc_hd__a21o_4
X_70958_ _49241_/B _70936_/X _70957_/Y _70958_/Y sky130_fd_sc_hd__o21ai_4
X_46694_ _46712_/A _51791_/B _46694_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_976_0_CLK clkbuf_9_488_0_CLK/X _86155_/CLK sky130_fd_sc_hd__clkbuf_1
X_60711_ _60711_/A _60711_/X sky130_fd_sc_hd__buf_2
X_48433_ _83586_/Q _53651_/B sky130_fd_sc_hd__inv_2
X_79253_ _79225_/Y _79251_/Y _79252_/Y _79253_/Y sky130_fd_sc_hd__a21oi_4
X_45645_ _57137_/A _45801_/A _45645_/Y sky130_fd_sc_hd__nor2_4
X_76465_ _76440_/X _76437_/X _76482_/C sky130_fd_sc_hd__nand2_4
X_42857_ _42856_/Y _87684_/D sky130_fd_sc_hd__inv_2
X_61691_ _61689_/X _61645_/X _61690_/Y _84459_/D sky130_fd_sc_hd__a21oi_4
X_73677_ _73677_/A _73599_/B _73677_/Y sky130_fd_sc_hd__nor2_4
X_70889_ _50971_/B _70885_/X _70888_/Y _70889_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_467_0_CLK clkbuf_9_467_0_CLK/A clkbuf_9_467_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_78204_ _78204_/A _78204_/B _78205_/B sky130_fd_sc_hd__and2_4
X_63430_ _64272_/A _63465_/B _63418_/C _63465_/D _63430_/Y sky130_fd_sc_hd__nand4_4
X_75416_ _75416_/A _75416_/Y sky130_fd_sc_hd__inv_2
X_41808_ _41802_/X _41803_/X _40395_/X _66704_/B _41792_/X _41808_/Y
+ sky130_fd_sc_hd__o32ai_4
X_48364_ _46485_/X _48364_/X sky130_fd_sc_hd__buf_2
X_60642_ _60642_/A _60638_/Y _60642_/C _60662_/A sky130_fd_sc_hd__nand3_4
X_72628_ _79160_/B _79158_/A sky130_fd_sc_hd__inv_2
X_79184_ _79184_/A _79184_/B _79185_/C sky130_fd_sc_hd__nand2_4
X_45576_ _55529_/B _45464_/X _44964_/X _45576_/Y sky130_fd_sc_hd__o21ai_4
X_76396_ _76392_/Y _76394_/Y _76395_/Y _76396_/X sky130_fd_sc_hd__o21a_4
X_42788_ _42822_/A _42788_/X sky130_fd_sc_hd__buf_2
X_47315_ _47287_/X _52979_/B _47315_/Y sky130_fd_sc_hd__nand2_4
X_78135_ _82569_/Q _78124_/B _78134_/Y _78135_/Y sky130_fd_sc_hd__a21oi_4
X_44527_ _44512_/X _44513_/X _40792_/X _44526_/Y _44516_/X _87066_/D
+ sky130_fd_sc_hd__o32ai_4
X_63361_ _61315_/A _60654_/X _60667_/Y _60758_/X _59477_/A _63361_/X
+ sky130_fd_sc_hd__a32o_4
X_75347_ _75330_/Y _75331_/Y _75333_/A _75347_/X sky130_fd_sc_hd__o21a_4
X_41739_ _82892_/Q _41718_/X _41739_/X sky130_fd_sc_hd__or2_4
X_48295_ _48319_/A _50341_/B _48295_/Y sky130_fd_sc_hd__nand2_4
X_60573_ _59831_/X _60610_/A sky130_fd_sc_hd__buf_2
X_72559_ _60312_/Y _72579_/A _72556_/Y _72557_/Y _72558_/X _72559_/Y
+ sky130_fd_sc_hd__o41ai_4
X_65100_ _64924_/A _65100_/B _65100_/X sky130_fd_sc_hd__and2_4
X_62312_ _62267_/A _62267_/B _76995_/B _62312_/Y sky130_fd_sc_hd__nor3_4
X_47246_ _47198_/X _47246_/X sky130_fd_sc_hd__buf_2
X_66080_ _66077_/Y _66065_/X _66079_/X _84158_/D sky130_fd_sc_hd__a21o_4
X_78066_ _78066_/A _78066_/B _78066_/X sky130_fd_sc_hd__xor2_4
X_44458_ _41129_/Y _44453_/X _87100_/Q _44454_/X _87100_/D sky130_fd_sc_hd__a2bb2o_4
X_63292_ _63216_/X _63292_/B _63333_/C _63240_/X _63292_/X sky130_fd_sc_hd__and4_4
X_75278_ _75303_/B _75284_/A sky130_fd_sc_hd__inv_2
X_65031_ _65031_/A _65031_/B _65031_/Y sky130_fd_sc_hd__nand2_4
X_77017_ _77017_/A _77017_/B _82365_/D sky130_fd_sc_hd__xnor2_4
X_43409_ _43408_/Y _43409_/Y sky130_fd_sc_hd__inv_2
X_62243_ _62218_/A _62244_/C sky130_fd_sc_hd__buf_2
X_74229_ _88342_/Q _72865_/X _72982_/X _74229_/Y sky130_fd_sc_hd__o21ai_4
X_47177_ _47128_/A _47177_/X sky130_fd_sc_hd__buf_2
X_44389_ _41465_/X _44377_/X _87134_/Q _44379_/X _87134_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_10_914_0_CLK clkbuf_9_457_0_CLK/X _83139_/CLK sky130_fd_sc_hd__clkbuf_1
X_46128_ _46128_/A _46204_/D _46143_/A _46128_/D _46133_/A sky130_fd_sc_hd__and4_4
X_62174_ _58990_/A _62174_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_3_0_CLK clkbuf_9_1_0_CLK/X _85241_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_5_31_0_CLK clkbuf_5_30_0_CLK/A clkbuf_6_63_0_CLK/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_9_405_0_CLK clkbuf_8_202_0_CLK/X clkbuf_9_405_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_61125_ _61125_/A _64203_/B _64525_/B _61188_/B sky130_fd_sc_hd__nand3_4
X_46059_ _41552_/A _46043_/X _66985_/B _46044_/X _86789_/D sky130_fd_sc_hd__a2bb2o_4
X_69770_ _69770_/A _88324_/Q _69770_/X sky130_fd_sc_hd__and2_4
X_66982_ _67057_/A _66982_/B _66982_/X sky130_fd_sc_hd__and2_4
X_78968_ _78968_/A _78967_/Y _78969_/A sky130_fd_sc_hd__xor2_4
X_68721_ _68721_/A _69956_/A sky130_fd_sc_hd__buf_2
X_65933_ _65845_/X _86239_/Q _65904_/X _65932_/X _65933_/X sky130_fd_sc_hd__a211o_4
X_61056_ _60961_/X _60908_/X _63738_/B _60995_/Y _61055_/X _61056_/X
+ sky130_fd_sc_hd__o41a_4
X_77919_ _82247_/Q _77919_/B _77919_/Y sky130_fd_sc_hd__xnor2_4
Xclkbuf_10_929_0_CLK clkbuf_9_464_0_CLK/X _88108_/CLK sky130_fd_sc_hd__clkbuf_1
X_78899_ _78894_/Y _78898_/Y _78899_/Y sky130_fd_sc_hd__nand2_4
X_60007_ _60007_/A _84675_/D sky130_fd_sc_hd__inv_2
X_49818_ _49830_/A _49830_/B _49795_/X _53031_/D _49818_/X sky130_fd_sc_hd__and4_4
X_80930_ _81059_/CLK _75079_/B _80930_/Q sky130_fd_sc_hd__dfxtp_4
X_68652_ _68599_/A _87752_/Q _68652_/X sky130_fd_sc_hd__and2_4
X_65864_ _64683_/A _65868_/B sky130_fd_sc_hd__buf_2
X_67603_ _67675_/A _87656_/Q _67603_/X sky130_fd_sc_hd__and2_4
X_64815_ _64637_/X _64913_/B _84226_/Q _64815_/X sky130_fd_sc_hd__and3_4
X_49749_ _57832_/B _49742_/X _49748_/Y _49749_/Y sky130_fd_sc_hd__o21ai_4
X_68583_ _68579_/X _68582_/X _68512_/X _68583_/Y sky130_fd_sc_hd__a21oi_4
X_80861_ _80740_/CLK _80893_/Q _75040_/B sky130_fd_sc_hd__dfxtp_4
X_65795_ _65717_/X _85577_/Q _65718_/X _65794_/X _65795_/X sky130_fd_sc_hd__a211o_4
X_82600_ _82924_/CLK _78862_/B _82568_/D sky130_fd_sc_hd__dfxtp_4
X_67534_ _67460_/A _87659_/Q _67534_/X sky130_fd_sc_hd__and2_4
X_52760_ _52744_/A _52760_/B _52760_/Y sky130_fd_sc_hd__nand2_4
X_64746_ _64678_/X _85532_/Q _64679_/X _64745_/X _64746_/X sky130_fd_sc_hd__a211o_4
X_83580_ _83068_/CLK _71182_/Y _48503_/A sky130_fd_sc_hd__dfxtp_4
X_80792_ _80792_/CLK _75781_/Y _75408_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_6_5_0_CLK clkbuf_6_5_0_CLK/A clkbuf_6_5_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_61958_ _61947_/X _61950_/X _61957_/Y _84739_/Q _61895_/X _61958_/Y
+ sky130_fd_sc_hd__o32ai_4
X_51711_ _51708_/Y _51693_/X _51710_/X _85960_/D sky130_fd_sc_hd__a21oi_4
X_82531_ _82531_/CLK _82531_/D _78960_/B sky130_fd_sc_hd__dfxtp_4
X_60909_ _60909_/A _60909_/X sky130_fd_sc_hd__buf_2
X_67465_ _67461_/X _67464_/X _67442_/X _67465_/X sky130_fd_sc_hd__a21o_4
X_52691_ _52687_/Y _52673_/X _52690_/X _52691_/Y sky130_fd_sc_hd__a21oi_4
X_64677_ _64650_/X _86174_/Q _64583_/X _64676_/X _64677_/X sky130_fd_sc_hd__a211o_4
X_61889_ _61448_/X _61874_/B _61907_/C _61874_/D _61889_/Y sky130_fd_sc_hd__nand4_4
X_69204_ _88046_/Q _69162_/X _69202_/X _69203_/X _69204_/X sky130_fd_sc_hd__a211o_4
X_54430_ _54426_/Y _54422_/X _54429_/X _85444_/D sky130_fd_sc_hd__a21oi_4
X_66416_ _66413_/Y _66414_/X _66415_/X _66416_/X sky130_fd_sc_hd__a21o_4
X_85250_ _85250_/CLK _56281_/Y _56280_/C sky130_fd_sc_hd__dfxtp_4
X_51642_ _51638_/Y _51639_/X _51641_/X _85973_/D sky130_fd_sc_hd__a21oi_4
X_63628_ _58396_/Y _63626_/X _61597_/A _63627_/X _63628_/X sky130_fd_sc_hd__a2bb2o_4
X_82462_ _82462_/CLK _82462_/D _82462_/Q sky130_fd_sc_hd__dfxtp_4
X_67396_ _87473_/Q _67394_/X _67344_/X _67395_/X _67396_/X sky130_fd_sc_hd__a211o_4
X_84201_ _85315_/CLK _84201_/D _84201_/Q sky130_fd_sc_hd__dfxtp_4
X_81413_ _82053_/CLK _81445_/Q _75940_/B sky130_fd_sc_hd__dfxtp_4
X_69135_ _88051_/Q _69121_/X _69051_/X _69134_/X _69135_/X sky130_fd_sc_hd__a211o_4
X_54361_ _85456_/Q _54349_/X _54360_/Y _54361_/Y sky130_fd_sc_hd__o21ai_4
X_66347_ _66267_/X _85890_/Q _66347_/X sky130_fd_sc_hd__and2_4
X_85181_ _85180_/CLK _85181_/D _55949_/B sky130_fd_sc_hd__dfxtp_4
X_51573_ _85985_/Q _51566_/X _51572_/Y _51573_/Y sky130_fd_sc_hd__o21ai_4
X_63559_ _63372_/A _63559_/X sky130_fd_sc_hd__buf_2
X_82393_ _86104_/CLK _82393_/D _82393_/Q sky130_fd_sc_hd__dfxtp_4
X_56100_ _56100_/A _56115_/B _85296_/Q _56100_/Y sky130_fd_sc_hd__nand3_4
X_53312_ _53330_/A _53293_/B _53302_/X _52797_/D _53312_/X sky130_fd_sc_hd__and4_4
X_84132_ _82975_/CLK _84132_/D _79455_/B sky130_fd_sc_hd__dfxtp_4
X_50524_ _51010_/A _50551_/A sky130_fd_sc_hd__buf_2
X_57080_ _56976_/X _57318_/D _46178_/X _57080_/X sky130_fd_sc_hd__o21a_4
X_81344_ _81344_/CLK _76629_/Y _81720_/D sky130_fd_sc_hd__dfxtp_4
X_69066_ _69065_/X _69066_/X sky130_fd_sc_hd__buf_2
X_54292_ _54312_/A _54298_/B _54312_/C _46658_/A _54292_/X sky130_fd_sc_hd__and4_4
X_66278_ _66065_/A _66278_/X sky130_fd_sc_hd__buf_2
X_56031_ _56030_/X _56031_/X sky130_fd_sc_hd__buf_2
X_68017_ _81477_/D _67925_/X _68016_/X _84045_/D sky130_fd_sc_hd__a21bo_4
X_53243_ _53190_/A _53243_/X sky130_fd_sc_hd__buf_2
X_65229_ _65226_/X _65228_/X _65122_/X _65233_/A sky130_fd_sc_hd__a21o_4
X_84063_ _82648_/CLK _67590_/X _84063_/Q sky130_fd_sc_hd__dfxtp_4
X_50455_ _50491_/A _50455_/X sky130_fd_sc_hd__buf_2
X_81275_ _81275_/CLK _81275_/D _76522_/A sky130_fd_sc_hd__dfxtp_4
X_83014_ _86869_/CLK _83014_/D _83014_/Q sky130_fd_sc_hd__dfxtp_4
X_80226_ _80226_/A _80226_/Y sky130_fd_sc_hd__inv_2
X_53174_ _53187_/A _53174_/B _53174_/Y sky130_fd_sc_hd__nand2_4
X_50386_ _50384_/Y _50380_/X _50385_/Y _86211_/D sky130_fd_sc_hd__a21boi_4
X_52125_ _52152_/A _52125_/X sky130_fd_sc_hd__buf_2
X_87822_ _87821_/CLK _87822_/D _42555_/A sky130_fd_sc_hd__dfxtp_4
X_80157_ _80157_/A _80135_/X _80157_/X sky130_fd_sc_hd__and2_4
X_57982_ _57837_/A _58858_/A sky130_fd_sc_hd__buf_2
X_69968_ _87540_/Q _66529_/X _68436_/X _69967_/X _69968_/X sky130_fd_sc_hd__a211o_4
X_59721_ _59721_/A _59721_/X sky130_fd_sc_hd__buf_2
X_56933_ _72909_/A _56933_/X sky130_fd_sc_hd__buf_2
X_52056_ _52070_/A _48310_/B _52056_/Y sky130_fd_sc_hd__nand2_4
X_68919_ _87997_/Q _68895_/X _68916_/X _68918_/X _68919_/X sky130_fd_sc_hd__a211o_4
X_87753_ _87757_/CLK _87753_/D _68624_/B sky130_fd_sc_hd__dfxtp_4
X_84965_ _85895_/CLK _84965_/D _84965_/Q sky130_fd_sc_hd__dfxtp_4
X_80088_ _80081_/X _80088_/B _80088_/Y sky130_fd_sc_hd__nand2_4
X_69899_ _69896_/X _69898_/X _69624_/X _69902_/A sky130_fd_sc_hd__a21o_4
X_51007_ _51004_/Y _50983_/X _51006_/X _86091_/D sky130_fd_sc_hd__a21oi_4
X_86704_ _86384_/CLK _86704_/D _86704_/Q sky130_fd_sc_hd__dfxtp_4
X_71930_ _71570_/X _71930_/B _71377_/B _71930_/Y sky130_fd_sc_hd__nor3_4
X_83916_ _83918_/CLK _83916_/D _81380_/D sky130_fd_sc_hd__dfxtp_4
X_59652_ _80625_/A _59509_/X _59632_/X _59713_/A _59652_/X sky130_fd_sc_hd__o22a_4
X_56864_ _56857_/X _56862_/Y _56863_/X _56756_/X _56864_/X sky130_fd_sc_hd__a211o_4
X_87684_ _87684_/CLK _87684_/D _66927_/B sky130_fd_sc_hd__dfxtp_4
X_84896_ _84344_/CLK _58257_/X _58254_/A sky130_fd_sc_hd__dfxtp_4
X_58603_ _58603_/A _58603_/X sky130_fd_sc_hd__buf_2
X_55815_ _85198_/Q _55342_/X _55457_/X _55814_/X _55815_/X sky130_fd_sc_hd__a211o_4
X_86635_ _85993_/CLK _86635_/D _86635_/Q sky130_fd_sc_hd__dfxtp_4
X_71861_ _70558_/X _71857_/B _71851_/X _71857_/D _71861_/Y sky130_fd_sc_hd__nor4_4
X_59583_ _61071_/C _59615_/A sky130_fd_sc_hd__buf_2
X_83847_ _83843_/CLK _83847_/D _83847_/Q sky130_fd_sc_hd__dfxtp_4
X_56795_ _83324_/Q _56794_/Y _56796_/B sky130_fd_sc_hd__xor2_4
X_73600_ _68418_/B _73597_/X _73464_/X _73599_/Y _73600_/X sky130_fd_sc_hd__a211o_4
X_70812_ _70810_/A _70945_/B _70810_/C _70812_/Y sky130_fd_sc_hd__nand3_4
X_58534_ _58517_/X _58530_/Y _58533_/Y _84826_/D sky130_fd_sc_hd__a21oi_4
X_43760_ _43760_/A _43760_/X sky130_fd_sc_hd__buf_2
X_55746_ _56127_/B _56127_/C _56117_/A sky130_fd_sc_hd__nor2_4
X_86566_ _85895_/CLK _48121_/Y _66298_/B sky130_fd_sc_hd__dfxtp_4
X_74580_ _74575_/X _74569_/X _56079_/A _74570_/X _74580_/X sky130_fd_sc_hd__a211o_4
X_40972_ _40972_/A _40972_/X sky130_fd_sc_hd__buf_2
X_52958_ _52903_/X _52979_/A sky130_fd_sc_hd__buf_2
X_71792_ _71235_/A _71302_/X _71785_/X _71792_/Y sky130_fd_sc_hd__nand3_4
X_83778_ _85953_/CLK _83778_/D _83778_/Q sky130_fd_sc_hd__dfxtp_4
X_88305_ _87333_/CLK _88305_/D _88305_/Q sky130_fd_sc_hd__dfxtp_4
X_42711_ _42681_/A _42711_/X sky130_fd_sc_hd__buf_2
X_73531_ _43203_/Y _73529_/X _73464_/X _73530_/Y _73531_/X sky130_fd_sc_hd__a211o_4
X_85517_ _85516_/CLK _54044_/Y _85517_/Q sky130_fd_sc_hd__dfxtp_4
X_51909_ _51887_/A _51898_/B _51893_/C _52735_/D _51909_/X sky130_fd_sc_hd__and4_4
X_70743_ _53105_/B _70738_/X _70742_/Y _83712_/D sky130_fd_sc_hd__o21ai_4
X_58465_ _58465_/A _58474_/B _58465_/Y sky130_fd_sc_hd__nor2_4
X_82729_ _84111_/CLK _66490_/C _78869_/A sky130_fd_sc_hd__dfxtp_4
X_43691_ _40810_/X _43685_/X _87306_/Q _43686_/X _87306_/D sky130_fd_sc_hd__a2bb2o_4
X_55677_ _83321_/Q _55681_/A sky130_fd_sc_hd__inv_2
X_86497_ _85888_/CLK _48716_/Y _65425_/B sky130_fd_sc_hd__dfxtp_4
X_52889_ _52885_/A _52889_/B _52889_/Y sky130_fd_sc_hd__nand2_4
X_45430_ _55622_/B _44935_/X _45429_/X _45430_/X sky130_fd_sc_hd__o21a_4
X_57416_ _57416_/A _57400_/X _57416_/C _57416_/Y sky130_fd_sc_hd__nand3_4
X_76250_ _76245_/Y _76250_/Y sky130_fd_sc_hd__inv_2
X_88236_ _88220_/CLK _41323_/Y _88236_/Q sky130_fd_sc_hd__dfxtp_4
X_42642_ _42641_/Y _87791_/D sky130_fd_sc_hd__inv_2
X_54628_ _85407_/Q _54621_/X _54627_/Y _54628_/Y sky130_fd_sc_hd__o21ai_4
X_73462_ _73462_/A _73198_/B _73462_/Y sky130_fd_sc_hd__nor2_4
X_85448_ _85770_/CLK _85448_/D _85448_/Q sky130_fd_sc_hd__dfxtp_4
X_70674_ _70664_/X _47458_/A _70673_/Y _70674_/X sky130_fd_sc_hd__a21o_4
X_58396_ _84859_/Q _58396_/Y sky130_fd_sc_hd__inv_2
X_75201_ _75201_/A _75201_/B _75201_/Y sky130_fd_sc_hd__nand2_4
X_72413_ _59325_/A _72413_/X sky130_fd_sc_hd__buf_2
X_45361_ _45678_/A _45361_/X sky130_fd_sc_hd__buf_2
X_57347_ _57289_/B _56848_/X _56850_/X _57347_/Y sky130_fd_sc_hd__nor3_4
X_88167_ _86934_/CLK _88167_/D _67634_/B sky130_fd_sc_hd__dfxtp_4
X_76181_ _76181_/A _76182_/B sky130_fd_sc_hd__inv_2
X_42573_ _42610_/A _42573_/X sky130_fd_sc_hd__buf_2
X_54559_ _54538_/A _54559_/B _54538_/C _54559_/D _54559_/X sky130_fd_sc_hd__and4_4
X_73393_ _73343_/X _73393_/X sky130_fd_sc_hd__buf_2
X_85379_ _85379_/CLK _85379_/D _85379_/Q sky130_fd_sc_hd__dfxtp_4
X_47100_ _47109_/A _52855_/B _47100_/Y sky130_fd_sc_hd__nand2_4
X_44312_ _44139_/X _44141_/X _44142_/X _44300_/Y _44312_/Y sky130_fd_sc_hd__nand4_4
X_75132_ _75131_/Y _75133_/B sky130_fd_sc_hd__inv_2
X_87118_ _87686_/CLK _87118_/D _87118_/Q sky130_fd_sc_hd__dfxtp_4
X_41524_ _41481_/X _82324_/Q _41523_/X _41524_/Y sky130_fd_sc_hd__o21ai_4
X_48080_ _48074_/Y _48055_/X _48079_/X _86570_/D sky130_fd_sc_hd__a21oi_4
X_72344_ _72201_/A _72344_/X sky130_fd_sc_hd__buf_2
X_45292_ _45289_/X _45291_/Y _45275_/X _45292_/Y sky130_fd_sc_hd__a21oi_4
X_57278_ _57276_/X _57277_/Y _57322_/B _57278_/Y sky130_fd_sc_hd__a21oi_4
X_88098_ _88097_/CLK _41944_/Y _73963_/A sky130_fd_sc_hd__dfxtp_4
X_47031_ _47031_/A _53332_/B sky130_fd_sc_hd__inv_2
X_59017_ _84776_/Q _58956_/X _59009_/X _59016_/X _84776_/D sky130_fd_sc_hd__a2bb2oi_4
X_56229_ _56233_/A _56229_/B _85267_/Q _56229_/Y sky130_fd_sc_hd__nand3_4
X_44243_ _44241_/Y _44242_/Y _44256_/A _87178_/D sky130_fd_sc_hd__a21oi_4
X_75063_ _75062_/A _75062_/B _75063_/Y sky130_fd_sc_hd__nand2_4
X_79940_ _79939_/Y _79940_/Y sky130_fd_sc_hd__inv_2
X_87049_ _88326_/CLK _44576_/Y _87049_/Q sky130_fd_sc_hd__dfxtp_4
X_41455_ _41486_/A _41455_/X sky130_fd_sc_hd__buf_2
X_72275_ _72270_/X _72272_/Y _72273_/Y _72189_/X _72274_/X _72275_/X
+ sky130_fd_sc_hd__o32a_4
X_74014_ _74038_/A _85902_/Q _74014_/X sky130_fd_sc_hd__and2_4
X_40406_ _82329_/Q _40385_/B _40406_/X sky130_fd_sc_hd__or2_4
X_71226_ _71232_/A _71226_/B _71232_/C _71226_/Y sky130_fd_sc_hd__nand3_4
X_44174_ _44174_/A _44175_/A sky130_fd_sc_hd__buf_2
X_79871_ _81024_/D _83280_/Q _79871_/X sky130_fd_sc_hd__xor2_4
X_41386_ _41373_/X _41729_/A _41385_/X _41387_/A sky130_fd_sc_hd__o21a_4
X_43125_ _44530_/A _43125_/X sky130_fd_sc_hd__buf_2
X_78822_ _78810_/Y _78818_/Y _78816_/Y _78830_/A sky130_fd_sc_hd__a21oi_4
X_40337_ _40343_/A _40591_/B _43175_/B _40337_/X sky130_fd_sc_hd__and3_4
X_71157_ _71183_/A _71155_/B _71160_/C _71160_/D _71157_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_10_270_0_CLK clkbuf_9_135_0_CLK/X _83438_/CLK sky130_fd_sc_hd__clkbuf_1
X_48982_ _72007_/B _48982_/X sky130_fd_sc_hd__buf_2
X_70108_ _83127_/Q _70108_/Y sky130_fd_sc_hd__inv_2
X_47933_ _66037_/B _47897_/X _47932_/Y _47933_/Y sky130_fd_sc_hd__o21ai_4
X_59919_ _59918_/Y _62475_/A sky130_fd_sc_hd__buf_2
X_43056_ _43053_/X _43054_/X _40646_/X _43055_/Y _43034_/X _43056_/Y
+ sky130_fd_sc_hd__o32ai_4
X_78753_ _78749_/Y _78753_/B _78753_/C _78758_/A sky130_fd_sc_hd__or3_4
X_71088_ _71088_/A _71064_/B _71088_/C _71088_/Y sky130_fd_sc_hd__nand3_4
X_75965_ _75964_/X _81736_/D sky130_fd_sc_hd__buf_2
Xclkbuf_10_52_0_CLK clkbuf_9_26_0_CLK/X _85031_/CLK sky130_fd_sc_hd__clkbuf_1
X_42007_ _42025_/A _42007_/X sky130_fd_sc_hd__buf_2
X_77704_ _77695_/A _77695_/B _77703_/B _77704_/Y sky130_fd_sc_hd__o21ai_4
X_62930_ _62930_/A _62930_/B _84369_/Q _62930_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_9_391_0_CLK clkbuf_9_391_0_CLK/A clkbuf_9_391_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_74916_ _81131_/D _74916_/B _74916_/Y sky130_fd_sc_hd__nand2_4
X_70039_ _83866_/Q _70029_/X _70038_/X _83866_/D sky130_fd_sc_hd__a21bo_4
X_47864_ _47863_/Y _51947_/B sky130_fd_sc_hd__buf_2
X_78684_ _78684_/A _78684_/B _78684_/X sky130_fd_sc_hd__and2_4
X_75896_ _61265_/C _84366_/Q _75896_/X sky130_fd_sc_hd__xor2_4
X_49603_ _49610_/A _49592_/B _49615_/C _52818_/D _49603_/X sky130_fd_sc_hd__and4_4
X_46815_ _83668_/Q _52692_/B sky130_fd_sc_hd__inv_2
Xclkbuf_10_285_0_CLK clkbuf_9_142_0_CLK/X _83745_/CLK sky130_fd_sc_hd__clkbuf_1
X_77635_ _77614_/A _77614_/B _77612_/Y _77635_/X sky130_fd_sc_hd__o21a_4
X_62861_ _62667_/X _62911_/C sky130_fd_sc_hd__buf_2
X_74847_ _74846_/Y _80653_/D sky130_fd_sc_hd__inv_2
X_47795_ _47804_/A _49364_/B _47777_/C _53249_/D _47795_/X sky130_fd_sc_hd__and4_4
X_64600_ _64600_/A _64600_/X sky130_fd_sc_hd__buf_2
X_49534_ _49531_/Y _49514_/X _49533_/X _86370_/D sky130_fd_sc_hd__a21oi_4
X_61812_ _61747_/X _61846_/D sky130_fd_sc_hd__buf_2
X_46746_ _46742_/Y _46704_/X _46745_/X _86708_/D sky130_fd_sc_hd__a21oi_4
X_65580_ _65387_/A _73042_/B _65580_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_67_0_CLK clkbuf_9_33_0_CLK/X _86887_/CLK sky130_fd_sc_hd__clkbuf_1
X_77566_ _82233_/Q _77570_/A sky130_fd_sc_hd__inv_2
X_43958_ _44104_/A _43954_/X _43955_/Y _43957_/X _43959_/B sky130_fd_sc_hd__a211o_4
X_62792_ _62791_/X _62792_/X sky130_fd_sc_hd__buf_2
X_74778_ _74804_/A _74778_/B _74804_/C _74804_/D _74778_/X sky130_fd_sc_hd__and4_4
X_79305_ _79297_/A _79296_/Y _79304_/X _79306_/B sky130_fd_sc_hd__o21ai_4
X_64531_ _79554_/B _79552_/A sky130_fd_sc_hd__inv_2
Xclkbuf_8_213_0_CLK clkbuf_8_213_0_CLK/A clkbuf_9_427_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_76517_ _76517_/A _76516_/Y _76518_/B sky130_fd_sc_hd__xor2_4
X_42909_ _42895_/X _42896_/X _41688_/X _87657_/Q _42905_/X _42909_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49465_ _58804_/B _49443_/X _49464_/Y _49465_/Y sky130_fd_sc_hd__o21ai_4
X_61743_ _61329_/B _62149_/B _61761_/C _62130_/D _61743_/Y sky130_fd_sc_hd__nand4_4
X_73729_ _88364_/Q _73633_/X _73704_/X _73729_/Y sky130_fd_sc_hd__o21ai_4
X_46677_ _46712_/A _51779_/B _46677_/Y sky130_fd_sc_hd__nand2_4
X_77497_ _77497_/A _77502_/A sky130_fd_sc_hd__inv_2
X_43889_ _41312_/X _43886_/X _67453_/B _43887_/X _87214_/D sky130_fd_sc_hd__a2bb2o_4
X_48416_ _48416_/A _52123_/B sky130_fd_sc_hd__buf_2
X_67250_ _67250_/A _86778_/Q _67250_/X sky130_fd_sc_hd__and2_4
X_79236_ _79236_/A _79236_/Y sky130_fd_sc_hd__inv_2
X_45628_ _45281_/A _45801_/A sky130_fd_sc_hd__buf_2
X_64462_ _64490_/A _64490_/B _79658_/B _64462_/Y sky130_fd_sc_hd__nor3_4
X_76448_ _76441_/X _76448_/B _76449_/B sky130_fd_sc_hd__xor2_4
X_49396_ _49451_/A _49420_/B sky130_fd_sc_hd__buf_2
X_61674_ _84732_/Q _61675_/B sky130_fd_sc_hd__buf_2
X_66201_ _66011_/X _86541_/Q _66201_/X sky130_fd_sc_hd__and2_4
X_63413_ _63413_/A _63463_/C sky130_fd_sc_hd__buf_2
X_48347_ _48148_/B _50385_/B sky130_fd_sc_hd__buf_2
X_60625_ _60624_/X _60694_/C sky130_fd_sc_hd__buf_2
X_67181_ _67178_/X _67180_/X _67085_/X _67181_/X sky130_fd_sc_hd__a21o_4
X_79167_ _79165_/Y _79173_/A _79171_/A sky130_fd_sc_hd__nand2_4
X_45559_ _45272_/A _45654_/B sky130_fd_sc_hd__buf_2
X_64393_ _64344_/X _64379_/B _84826_/Q _64393_/X sky130_fd_sc_hd__and3_4
X_76379_ _76377_/Y _76379_/B _76379_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_8_228_0_CLK clkbuf_8_229_0_CLK/A clkbuf_8_228_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_66132_ _66226_/A _86546_/Q _66132_/X sky130_fd_sc_hd__and2_4
X_78118_ _78130_/C _78120_/B sky130_fd_sc_hd__inv_2
X_63344_ _63344_/A _63344_/B _60588_/X _63344_/D _63344_/X sky130_fd_sc_hd__or4_4
Xclkbuf_10_223_0_CLK clkbuf_9_111_0_CLK/X _84603_/CLK sky130_fd_sc_hd__clkbuf_1
X_48278_ _48272_/Y _48273_/X _48277_/Y _48278_/Y sky130_fd_sc_hd__a21boi_4
X_60556_ _60555_/Y _60556_/B _60556_/Y sky130_fd_sc_hd__nand2_4
X_79098_ _79095_/X _82752_/Q _79109_/A _79099_/A sky130_fd_sc_hd__nand3_4
Xclkbuf_10_853_0_CLK clkbuf_9_426_0_CLK/X _82774_/CLK sky130_fd_sc_hd__clkbuf_1
X_47229_ _47223_/Y _47224_/X _47228_/X _86657_/D sky130_fd_sc_hd__a21oi_4
X_66063_ _66020_/X _66061_/Y _66062_/Y _66063_/Y sky130_fd_sc_hd__o21ai_4
X_78049_ _78049_/A _78049_/B _78049_/X sky130_fd_sc_hd__xor2_4
X_63275_ _63248_/X _63270_/Y _63271_/X _63272_/Y _63274_/Y _63275_/X
+ sky130_fd_sc_hd__a41o_4
X_60487_ _79152_/A _60246_/X _60481_/X _60486_/Y _84612_/D sky130_fd_sc_hd__a2bb2oi_4
X_65014_ _65011_/X _65013_/X _64989_/X _65014_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_9_344_0_CLK clkbuf_9_345_0_CLK/A clkbuf_9_344_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_50240_ _50240_/A _51947_/B _50240_/Y sky130_fd_sc_hd__nand2_4
X_62226_ _61338_/A _62631_/B _62631_/C _62225_/X _62234_/B sky130_fd_sc_hd__nand4_4
X_81060_ _82084_/CLK _81092_/Q _75100_/A sky130_fd_sc_hd__dfxtp_4
X_80011_ _79988_/A _80011_/B _79988_/B _80011_/D _80011_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_10_238_0_CLK clkbuf_9_119_0_CLK/X _80679_/CLK sky130_fd_sc_hd__clkbuf_1
X_69822_ _73247_/A _44299_/A _68933_/X _69821_/Y _69822_/X sky130_fd_sc_hd__a211o_4
X_50171_ _50131_/A _53902_/B _50171_/X sky130_fd_sc_hd__and2_4
X_62157_ _62065_/B _62063_/X _63694_/B _62183_/D _62157_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_868_0_CLK clkbuf_9_434_0_CLK/X _86404_/CLK sky130_fd_sc_hd__clkbuf_1
X_61108_ _61122_/B _61122_/C _61082_/X _61108_/Y sky130_fd_sc_hd__a21boi_4
X_69753_ _73126_/A _69751_/X _68070_/X _69752_/Y _69753_/X sky130_fd_sc_hd__a211o_4
X_66965_ _66960_/X _66963_/X _66964_/X _66965_/X sky130_fd_sc_hd__a21o_4
X_62088_ _59794_/X _62088_/B _62086_/Y _62087_/Y _62088_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_9_359_0_CLK clkbuf_8_179_0_CLK/X clkbuf_9_359_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_68704_ _68604_/A _87238_/Q _68704_/X sky130_fd_sc_hd__and2_4
X_53930_ _53949_/A _50714_/B _53930_/Y sky130_fd_sc_hd__nand2_4
X_65916_ _65916_/A _65916_/B _65916_/C _65916_/X sky130_fd_sc_hd__and3_4
X_61039_ _60950_/Y _60940_/Y _60902_/Y _76980_/A _61020_/X _84532_/D
+ sky130_fd_sc_hd__o32a_4
X_84750_ _85718_/CLK _59338_/Y _84750_/Q sky130_fd_sc_hd__dfxtp_4
X_81962_ _82299_/CLK _81962_/D _81962_/Q sky130_fd_sc_hd__dfxtp_4
X_69684_ _83905_/Q _69632_/X _69683_/X _83905_/D sky130_fd_sc_hd__a21bo_4
X_66896_ _80916_/D _66850_/X _66895_/X _84092_/D sky130_fd_sc_hd__a21bo_4
X_83701_ _83699_/CLK _70785_/Y _83701_/Q sky130_fd_sc_hd__dfxtp_4
X_80913_ _83918_/CLK _80913_/D _80913_/Q sky130_fd_sc_hd__dfxtp_4
X_68635_ _83967_/Q _68586_/X _68634_/X _83967_/D sky130_fd_sc_hd__a21bo_4
X_53861_ _85553_/Q _53846_/X _53860_/Y _53861_/Y sky130_fd_sc_hd__o21ai_4
X_65847_ _65845_/X _86181_/Q _65790_/X _65846_/X _65847_/X sky130_fd_sc_hd__a211o_4
X_84681_ _84498_/CLK _59956_/X _84681_/Q sky130_fd_sc_hd__dfxtp_4
X_81893_ _82009_/CLK _81893_/D _77194_/B sky130_fd_sc_hd__dfxtp_4
X_55600_ _45448_/A _55617_/A _55533_/X _55599_/X _55601_/B sky130_fd_sc_hd__a211o_4
X_86420_ _86422_/CLK _49274_/Y _86420_/Q sky130_fd_sc_hd__dfxtp_4
X_52812_ _52808_/Y _52809_/X _52811_/X _52812_/Y sky130_fd_sc_hd__a21oi_4
X_83632_ _83275_/CLK _83632_/D _47609_/A sky130_fd_sc_hd__dfxtp_4
X_56580_ _55504_/Y _56580_/B _56618_/B sky130_fd_sc_hd__nand2_4
X_80844_ _80754_/CLK _80876_/Q _74912_/B sky130_fd_sc_hd__dfxtp_4
X_68566_ _87595_/Q _68066_/X _68517_/X _68565_/X _68566_/X sky130_fd_sc_hd__a211o_4
X_53792_ _85567_/Q _53722_/X _53791_/Y _53792_/Y sky130_fd_sc_hd__o21ai_4
X_65778_ _65623_/X _86186_/Q _65517_/X _65777_/X _65778_/X sky130_fd_sc_hd__a211o_4
X_55531_ _55505_/X _55531_/X sky130_fd_sc_hd__buf_2
X_67517_ _67517_/A _88236_/Q _67517_/X sky130_fd_sc_hd__and2_4
X_86351_ _86351_/CLK _49637_/Y _86351_/Q sky130_fd_sc_hd__dfxtp_4
X_52743_ _52740_/Y _52728_/X _52742_/X _85763_/D sky130_fd_sc_hd__a21oi_4
X_64729_ _64729_/A _64729_/X sky130_fd_sc_hd__buf_2
X_83563_ _83623_/CLK _71233_/Y _48693_/A sky130_fd_sc_hd__dfxtp_4
X_80775_ _81059_/CLK _80775_/D _80775_/Q sky130_fd_sc_hd__dfxtp_4
X_68497_ _68492_/X _68496_/X _68390_/X _68497_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_10_806_0_CLK clkbuf_9_403_0_CLK/X _82570_/CLK sky130_fd_sc_hd__clkbuf_1
X_85302_ _85270_/CLK _85302_/D _55889_/B sky130_fd_sc_hd__dfxtp_4
X_58250_ _61985_/A _58251_/A sky130_fd_sc_hd__inv_2
X_82514_ _82610_/CLK _79115_/Y _82514_/Q sky130_fd_sc_hd__dfxtp_4
X_55462_ _55453_/X _55462_/X sky130_fd_sc_hd__buf_2
X_86282_ _86282_/CLK _86282_/D _72400_/B sky130_fd_sc_hd__dfxtp_4
X_67448_ _84069_/Q _67331_/X _67447_/X _67448_/X sky130_fd_sc_hd__a21bo_4
X_52674_ _52648_/A _52674_/X sky130_fd_sc_hd__buf_2
X_83494_ _83495_/CLK _71453_/X _83494_/Q sky130_fd_sc_hd__dfxtp_4
X_57201_ _57050_/A _44239_/A _57201_/Y sky130_fd_sc_hd__nand2_4
X_88021_ _87253_/CLK _42129_/X _88021_/Q sky130_fd_sc_hd__dfxtp_4
X_54413_ _54399_/X _54417_/B _54402_/C _46866_/Y _54413_/X sky130_fd_sc_hd__and4_4
X_85233_ _85167_/CLK _85233_/D _85233_/Q sky130_fd_sc_hd__dfxtp_4
X_51625_ _51619_/A _51619_/B _51608_/X _53151_/D _51625_/X sky130_fd_sc_hd__and4_4
X_58181_ _83377_/Q _58181_/Y sky130_fd_sc_hd__inv_2
X_82445_ _82820_/CLK _79137_/X _82445_/Q sky130_fd_sc_hd__dfxtp_4
X_55393_ _55443_/A _55393_/B _55443_/C _55443_/D _55394_/B sky130_fd_sc_hd__nand4_4
X_67379_ _87921_/Q _67355_/X _67284_/X _67378_/X _67379_/X sky130_fd_sc_hd__a211o_4
X_57132_ _56739_/X _57133_/A _57155_/D _57170_/B _83329_/Q _57132_/Y
+ sky130_fd_sc_hd__a41oi_4
X_69118_ _69073_/A _88340_/Q _69118_/X sky130_fd_sc_hd__and2_4
X_54344_ _54344_/A _54399_/A sky130_fd_sc_hd__buf_2
X_85164_ _80671_/CLK _85164_/D _85164_/Q sky130_fd_sc_hd__dfxtp_4
X_51556_ _85988_/Q _51539_/X _51555_/Y _51556_/Y sky130_fd_sc_hd__o21ai_4
X_70390_ _51378_/B _70364_/X _70389_/Y _70390_/Y sky130_fd_sc_hd__o21ai_4
X_82376_ _86054_/CLK _82184_/Q _82376_/Q sky130_fd_sc_hd__dfxtp_4
X_84115_ _84115_/CLK _66480_/X _84115_/Q sky130_fd_sc_hd__dfxtp_4
X_50507_ _50534_/A _50513_/A sky130_fd_sc_hd__buf_2
X_81327_ _81333_/CLK _76343_/X _75957_/A sky130_fd_sc_hd__dfxtp_4
X_57063_ _58517_/A _45808_/Y _57062_/Y _57063_/Y sky130_fd_sc_hd__o21ai_4
X_69049_ _87075_/Q _68818_/X _68819_/X _69048_/X _69049_/X sky130_fd_sc_hd__a211o_4
X_54275_ _54286_/A _54298_/B _54286_/C _54275_/D _54275_/X sky130_fd_sc_hd__and4_4
X_85095_ _85128_/CLK _57060_/X _57058_/B sky130_fd_sc_hd__dfxtp_4
X_51487_ _51491_/A _53012_/B _51487_/Y sky130_fd_sc_hd__nand2_4
X_56014_ _56013_/Y _74297_/C _56003_/B _55966_/X _56015_/B sky130_fd_sc_hd__nand4_4
X_41240_ _40637_/A _41490_/A sky130_fd_sc_hd__buf_2
X_53226_ _53199_/A _53246_/A sky130_fd_sc_hd__buf_2
X_72060_ _49089_/A _72043_/X _72048_/X _72060_/X sky130_fd_sc_hd__and3_4
X_84046_ _88116_/CLK _67996_/X _81478_/D sky130_fd_sc_hd__dfxtp_4
X_50438_ _50655_/A _50534_/A sky130_fd_sc_hd__buf_2
X_81258_ _81275_/CLK _81258_/D _81258_/Q sky130_fd_sc_hd__dfxtp_4
X_71011_ _70886_/A _71010_/X _70735_/X _70758_/C _71012_/B sky130_fd_sc_hd__nand4_4
X_80209_ _80209_/A _80209_/B _80209_/X sky130_fd_sc_hd__or2_4
X_41171_ _41013_/A _41223_/B sky130_fd_sc_hd__buf_2
X_53157_ _53147_/X _53157_/B _53157_/Y sky130_fd_sc_hd__nand2_4
X_50369_ _50366_/Y _50351_/X _50368_/Y _50369_/Y sky130_fd_sc_hd__a21boi_4
X_81189_ _81190_/CLK _81189_/D _81189_/Q sky130_fd_sc_hd__dfxtp_4
X_52108_ _52203_/A _52108_/X sky130_fd_sc_hd__buf_2
X_87805_ _87553_/CLK _42603_/Y _69859_/A sky130_fd_sc_hd__dfxtp_4
X_57965_ _57965_/A _58813_/A sky130_fd_sc_hd__buf_2
X_53088_ _53221_/A _53195_/A sky130_fd_sc_hd__buf_2
X_85997_ _85709_/CLK _85997_/D _85997_/Q sky130_fd_sc_hd__dfxtp_4
X_59704_ _59649_/A _59628_/A _59648_/A _59790_/B sky130_fd_sc_hd__a21o_4
X_44930_ _56381_/C _44880_/X _44929_/X _44930_/Y sky130_fd_sc_hd__o21ai_4
X_52039_ _52039_/A _52098_/B _52033_/X _52039_/X sky130_fd_sc_hd__and3_4
X_56916_ _56910_/X _56915_/Y _56917_/A sky130_fd_sc_hd__nand2_4
X_75750_ _81094_/Q _75750_/B _75750_/Y sky130_fd_sc_hd__xnor2_4
X_87736_ _87993_/CLK _87736_/D _69031_/B sky130_fd_sc_hd__dfxtp_4
X_72962_ _72958_/X _72961_/X _72812_/X _72966_/A sky130_fd_sc_hd__a21o_4
X_84948_ _85404_/CLK _84948_/D _84948_/Q sky130_fd_sc_hd__dfxtp_4
X_57896_ _57896_/A _57896_/X sky130_fd_sc_hd__buf_2
X_74701_ _74630_/X _56903_/X _74700_/Y _82980_/D sky130_fd_sc_hd__o21a_4
X_71913_ _70554_/A _71930_/B sky130_fd_sc_hd__buf_2
X_59635_ _59624_/X _59635_/Y sky130_fd_sc_hd__inv_2
X_44861_ _41777_/Y _44848_/X _86915_/Q _44849_/X _44861_/X sky130_fd_sc_hd__a2bb2o_4
X_56847_ _56846_/Y _57050_/A sky130_fd_sc_hd__buf_2
X_87667_ _87671_/CLK _42890_/Y _87667_/Q sky130_fd_sc_hd__dfxtp_4
X_75681_ _75669_/Y _80781_/D sky130_fd_sc_hd__inv_2
X_72893_ _41994_/Y _72888_/X _72890_/X _72892_/Y _72893_/X sky130_fd_sc_hd__a211o_4
X_84879_ _84849_/CLK _84879_/D _58319_/A sky130_fd_sc_hd__dfxtp_4
X_46600_ _46505_/A _46600_/B _46600_/Y sky130_fd_sc_hd__nand2_4
X_77420_ _77416_/X _77419_/Y _82191_/D sky130_fd_sc_hd__xor2_4
X_43812_ _43810_/X _43797_/X _41087_/X _69509_/B _43811_/X _43813_/A
+ sky130_fd_sc_hd__o32ai_4
X_74632_ _74675_/A _74691_/A sky130_fd_sc_hd__buf_2
X_86618_ _85981_/CLK _86618_/D _86618_/Q sky130_fd_sc_hd__dfxtp_4
X_47580_ _47575_/Y _47555_/X _47579_/X _47580_/Y sky130_fd_sc_hd__a21oi_4
X_71844_ _71824_/Y _83354_/Q _71843_/X _71844_/X sky130_fd_sc_hd__a21o_4
X_59566_ _59751_/A _60122_/A _59752_/A _60122_/C _60380_/B sky130_fd_sc_hd__and4_4
X_44792_ _44791_/Y _86953_/D sky130_fd_sc_hd__inv_2
X_56778_ _72765_/A _56776_/X _56777_/Y _56778_/Y sky130_fd_sc_hd__a21boi_4
X_87598_ _88111_/CLK _87598_/D _73677_/A sky130_fd_sc_hd__dfxtp_4
X_46531_ _46531_/A _50850_/B _46531_/Y sky130_fd_sc_hd__nand2_4
X_58517_ _58517_/A _58517_/X sky130_fd_sc_hd__buf_2
X_77351_ _77371_/C _77351_/B _82186_/D sky130_fd_sc_hd__xnor2_4
X_55729_ _55711_/X _85285_/Q _55172_/A _55729_/Y sky130_fd_sc_hd__a21oi_4
X_43743_ _43743_/A _87288_/D sky130_fd_sc_hd__inv_2
X_74563_ _45020_/A _74551_/X _74562_/X _74563_/Y sky130_fd_sc_hd__o21ai_4
X_86549_ _86549_/CLK _86549_/D _66087_/B sky130_fd_sc_hd__dfxtp_4
X_40955_ _40954_/Y _40955_/X sky130_fd_sc_hd__buf_2
X_71775_ _71779_/A _71333_/C _70986_/A _71775_/X sky130_fd_sc_hd__and3_4
X_59497_ _83428_/Q _59497_/Y sky130_fd_sc_hd__inv_2
X_76302_ _76301_/A _81561_/Q _76302_/Y sky130_fd_sc_hd__nand2_4
X_49250_ _49246_/Y _49247_/X _49249_/Y _86425_/D sky130_fd_sc_hd__a21boi_4
X_73514_ _73353_/A _85859_/Q _73514_/X sky130_fd_sc_hd__and2_4
X_46462_ _46408_/A _50816_/B _46462_/Y sky130_fd_sc_hd__nand2_4
X_70726_ _70848_/A _70779_/B sky130_fd_sc_hd__buf_2
X_58448_ _58423_/A _58448_/X sky130_fd_sc_hd__buf_2
X_77282_ _77264_/Y _82213_/Q _77265_/Y _77282_/Y sky130_fd_sc_hd__a21boi_4
X_43674_ _40753_/X _43671_/X _87317_/Q _43673_/X _87317_/D sky130_fd_sc_hd__a2bb2o_4
X_74494_ _74491_/Y _74492_/X _74493_/X _83055_/D sky130_fd_sc_hd__a21oi_4
X_40886_ _40870_/X _40871_/X _40885_/X _69865_/B _40867_/X _40887_/A
+ sky130_fd_sc_hd__o32ai_4
X_48201_ _47886_/X _48201_/B _48195_/X _48201_/X sky130_fd_sc_hd__and3_4
X_79021_ _79021_/A _79021_/B _79027_/A sky130_fd_sc_hd__xor2_4
X_45413_ _45413_/A _45397_/X _45413_/Y sky130_fd_sc_hd__nor2_4
X_76233_ _76232_/Y _81640_/Q _76233_/C _76233_/Y sky130_fd_sc_hd__nand3_4
X_88219_ _87141_/CLK _88219_/D _67909_/B sky130_fd_sc_hd__dfxtp_4
X_42625_ _49210_/B _50731_/A _40929_/X _69969_/B _42612_/X _42625_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49181_ _49181_/A _50714_/B sky130_fd_sc_hd__buf_2
X_73445_ _73442_/X _73444_/Y _73445_/Y sky130_fd_sc_hd__nand2_4
X_46393_ _46388_/Y _46346_/X _46392_/Y _46393_/Y sky130_fd_sc_hd__a21boi_4
X_70657_ _53046_/B _70631_/X _70656_/Y _83731_/D sky130_fd_sc_hd__o21ai_4
X_58379_ _84864_/Q _58380_/A sky130_fd_sc_hd__inv_2
X_48132_ _48142_/A _50378_/B _48132_/Y sky130_fd_sc_hd__nand2_4
XPHY_80 sky130_fd_sc_hd__decap_3
X_60410_ _60472_/A _60410_/B _60482_/A _63118_/A sky130_fd_sc_hd__nand3_4
X_45344_ _56165_/C _45343_/X _45303_/X _45344_/X sky130_fd_sc_hd__o21a_4
XPHY_91 sky130_fd_sc_hd__decap_3
X_76164_ _76155_/A _76155_/B _76164_/Y sky130_fd_sc_hd__nand2_4
X_42556_ _42556_/A _42556_/X sky130_fd_sc_hd__buf_2
X_73376_ _73373_/X _73375_/X _72737_/A _73376_/X sky130_fd_sc_hd__a21o_4
X_61390_ _61390_/A _61367_/B _61367_/C _61390_/D _61390_/Y sky130_fd_sc_hd__nand4_4
X_70588_ _70588_/A _70613_/B sky130_fd_sc_hd__buf_2
X_75115_ _75115_/A _75117_/A sky130_fd_sc_hd__inv_2
X_41507_ _41506_/Y _41507_/X sky130_fd_sc_hd__buf_2
X_48063_ _74083_/B _48049_/X _48062_/Y _48063_/Y sky130_fd_sc_hd__o21ai_4
X_60341_ _60341_/A _60341_/X sky130_fd_sc_hd__buf_2
X_72327_ _59085_/A _72327_/X sky130_fd_sc_hd__buf_2
X_45275_ _45714_/A _45275_/X sky130_fd_sc_hd__buf_2
X_76095_ _76082_/A _76096_/A _76097_/B _76095_/X sky130_fd_sc_hd__and3_4
X_42487_ _73820_/A _68641_/B sky130_fd_sc_hd__inv_2
Xclkbuf_7_74_0_CLK clkbuf_7_74_0_CLK/A clkbuf_7_74_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_47014_ _47009_/Y _46987_/X _47013_/X _86680_/D sky130_fd_sc_hd__a21oi_4
X_44226_ _44006_/X _44164_/X _44225_/Y _44226_/Y sky130_fd_sc_hd__nand3_4
X_63060_ _63060_/A _63060_/X sky130_fd_sc_hd__buf_2
X_75046_ _81150_/D _75046_/B _75046_/X sky130_fd_sc_hd__xor2_4
X_79923_ _60145_/Y _79921_/A _79924_/C sky130_fd_sc_hd__nand2_4
X_41438_ _41437_/X _41418_/X _88215_/Q _41419_/X _88215_/D sky130_fd_sc_hd__a2bb2o_4
X_60272_ _60271_/X _60273_/A sky130_fd_sc_hd__buf_2
X_72258_ _72123_/A _72258_/X sky130_fd_sc_hd__buf_2
X_62011_ _59823_/X _62011_/X sky130_fd_sc_hd__buf_2
X_71209_ _70400_/A _71232_/B sky130_fd_sc_hd__buf_2
X_44157_ _66180_/A _57776_/A _44152_/A _44157_/Y sky130_fd_sc_hd__a21oi_4
X_79854_ _79835_/X _79854_/B _79856_/B sky130_fd_sc_hd__or2_4
X_41369_ _41369_/A _41325_/X _41369_/X sky130_fd_sc_hd__or2_4
X_72189_ _58766_/A _72189_/X sky130_fd_sc_hd__buf_2
X_43108_ _43127_/A _43108_/X sky130_fd_sc_hd__buf_2
X_78805_ _82722_/Q _78805_/B _78805_/X sky130_fd_sc_hd__xor2_4
X_48965_ _86457_/Q _48952_/X _48964_/Y _48965_/Y sky130_fd_sc_hd__o21ai_4
X_44088_ _44088_/A _43987_/A _44313_/B _44090_/A sky130_fd_sc_hd__nand3_4
Xclkbuf_7_89_0_CLK clkbuf_7_89_0_CLK/A clkbuf_7_89_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_79785_ _79794_/A _79794_/B _79785_/Y sky130_fd_sc_hd__xnor2_4
X_76997_ _60947_/C _84421_/Q _76997_/X sky130_fd_sc_hd__xor2_4
X_47916_ _47867_/X _46337_/A _47915_/Y _47917_/A sky130_fd_sc_hd__o21ai_4
X_43039_ _43038_/X _43017_/X _40610_/X _73677_/A _43025_/X _43040_/A
+ sky130_fd_sc_hd__o32ai_4
X_66750_ _66746_/X _66749_/X _66726_/X _66750_/X sky130_fd_sc_hd__a21o_4
X_78736_ _78732_/X _78733_/Y _78735_/Y _78770_/A sky130_fd_sc_hd__a21o_4
X_63962_ _64081_/C _64180_/C _60889_/X _84955_/Q _63962_/X sky130_fd_sc_hd__and4_4
X_75948_ _75946_/Y _75942_/Y _75947_/Y _75948_/Y sky130_fd_sc_hd__o21ai_4
X_48896_ _48612_/A _48896_/X sky130_fd_sc_hd__buf_2
X_65701_ _65400_/A _65701_/X sky130_fd_sc_hd__buf_2
X_62913_ _62930_/A _62930_/B _84371_/Q _62913_/Y sky130_fd_sc_hd__nor3_4
X_47847_ _48144_/A _51282_/A sky130_fd_sc_hd__buf_2
X_66681_ _66677_/X _66680_/X _66606_/X _66681_/X sky130_fd_sc_hd__a21o_4
X_78667_ _78663_/X _78664_/Y _78666_/Y _78667_/X sky130_fd_sc_hd__a21o_4
X_63893_ _63972_/A _63894_/C sky130_fd_sc_hd__buf_2
X_75879_ _75876_/A _81025_/Q _75876_/B _75880_/B sky130_fd_sc_hd__nand3_4
Xclkbuf_7_12_0_CLK clkbuf_6_6_0_CLK/X clkbuf_8_25_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_68420_ _68417_/X _68419_/X _68390_/X _68420_/X sky130_fd_sc_hd__a21o_4
X_65632_ _65516_/X _64953_/Y _65631_/Y _65632_/Y sky130_fd_sc_hd__o21ai_4
X_77618_ _77614_/X _77619_/C _77619_/B _77664_/C sky130_fd_sc_hd__a21o_4
X_62844_ _62869_/A _62812_/B _63561_/B _62844_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_8_152_0_CLK clkbuf_7_76_0_CLK/X clkbuf_8_152_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_47778_ _47774_/Y _47745_/X _47777_/X _86599_/D sky130_fd_sc_hd__a21oi_4
X_78598_ _78596_/Y _78597_/X _78623_/A sky130_fd_sc_hd__xor2_4
X_49517_ _49513_/Y _49514_/X _49516_/X _86373_/D sky130_fd_sc_hd__a21oi_4
X_68351_ _87507_/Q _68472_/A _68348_/X _68350_/X _68351_/X sky130_fd_sc_hd__a211o_4
X_46729_ _46737_/A _46717_/B _46717_/C _46728_/X _46729_/X sky130_fd_sc_hd__and4_4
X_65563_ _65158_/A _65779_/A sky130_fd_sc_hd__buf_2
X_77549_ _77549_/A _77553_/A sky130_fd_sc_hd__inv_2
X_62775_ _61448_/X _62743_/B _62742_/X _62729_/D _62775_/Y sky130_fd_sc_hd__nand4_4
X_67302_ _67298_/X _67301_/X _67255_/X _67302_/Y sky130_fd_sc_hd__a21oi_4
X_64514_ _64474_/A _64306_/A _84886_/Q _64514_/X sky130_fd_sc_hd__and3_4
X_49448_ _49446_/Y _49434_/X _49447_/X _86386_/D sky130_fd_sc_hd__a21oi_4
X_61726_ _61770_/A _61770_/B _63369_/B _61770_/D _61726_/X sky130_fd_sc_hd__and4_4
X_80560_ _80560_/A _80560_/B _80561_/B sky130_fd_sc_hd__xnor2_4
X_68282_ _83993_/Q _68279_/X _68281_/X _83993_/D sky130_fd_sc_hd__a21bo_4
X_65494_ _65491_/X _65494_/B _65494_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_7_27_0_CLK clkbuf_7_26_0_CLK/A clkbuf_8_55_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_67233_ _67229_/X _67232_/X _67015_/X _67233_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_8_167_0_CLK clkbuf_7_83_0_CLK/X clkbuf_9_335_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_79219_ _79202_/Y _79219_/Y sky130_fd_sc_hd__inv_2
X_64445_ _58452_/A _64511_/B _64445_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_162_0_CLK clkbuf_9_81_0_CLK/X _81697_/CLK sky130_fd_sc_hd__clkbuf_1
X_61657_ _61657_/A _61657_/Y sky130_fd_sc_hd__inv_2
X_49379_ _49379_/A _49397_/A sky130_fd_sc_hd__buf_2
X_80491_ _80478_/X _80489_/X _80490_/X _80491_/Y sky130_fd_sc_hd__a21oi_4
X_51410_ _51218_/X _51410_/X sky130_fd_sc_hd__buf_2
X_82230_ _82515_/CLK _82262_/Q _77517_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_792_0_CLK clkbuf_9_396_0_CLK/X _82503_/CLK sky130_fd_sc_hd__clkbuf_1
X_60608_ _60608_/A _60608_/X sky130_fd_sc_hd__buf_2
X_67164_ _67141_/X _67151_/Y _67152_/X _67163_/Y _67164_/X sky130_fd_sc_hd__a211o_4
X_52390_ _52496_/A _52390_/X sky130_fd_sc_hd__buf_2
X_64376_ _64363_/A _64363_/B _84955_/Q _61145_/X _64376_/X sky130_fd_sc_hd__and4_4
X_61588_ _59829_/X _61586_/Y _61587_/X _61588_/X sky130_fd_sc_hd__o21a_4
X_66115_ _64971_/X _85619_/Q _44261_/X _66114_/X _66115_/X sky130_fd_sc_hd__a211o_4
X_51341_ _51842_/A _53671_/A sky130_fd_sc_hd__buf_2
X_63327_ _63325_/Y _63326_/X _63317_/X _63327_/X sky130_fd_sc_hd__a21o_4
X_82161_ _84220_/CLK _84153_/Q _82161_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_283_0_CLK clkbuf_9_283_0_CLK/A clkbuf_9_283_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_60539_ _60459_/B _60541_/B sky130_fd_sc_hd__buf_2
X_67095_ _67095_/A _67095_/B _67095_/X sky130_fd_sc_hd__and2_4
X_81112_ _80696_/CLK _79793_/X _81112_/Q sky130_fd_sc_hd__dfxtp_4
X_54060_ _53982_/A _54060_/X sky130_fd_sc_hd__buf_2
X_66046_ _66046_/A _66164_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_177_0_CLK clkbuf_9_88_0_CLK/X _80721_/CLK sky130_fd_sc_hd__clkbuf_1
X_51272_ _51280_/A _49241_/B _51272_/Y sky130_fd_sc_hd__nand2_4
X_63258_ _64314_/A _63258_/X sky130_fd_sc_hd__buf_2
X_82092_ _82103_/CLK _77376_/B _82092_/Q sky130_fd_sc_hd__dfxtp_4
X_53011_ _52903_/X _53025_/A sky130_fd_sc_hd__buf_2
X_50223_ _50222_/X _51737_/A sky130_fd_sc_hd__buf_2
X_85920_ _85920_/CLK _85920_/D _73583_/B sky130_fd_sc_hd__dfxtp_4
X_81043_ _80719_/CLK _75328_/X _81043_/Q sky130_fd_sc_hd__dfxtp_4
X_62209_ _62522_/B _62560_/C sky130_fd_sc_hd__buf_2
X_63189_ _64314_/A _63189_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_298_0_CLK clkbuf_9_299_0_CLK/A clkbuf_9_298_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_69805_ _69791_/A _69804_/Y _69805_/Y sky130_fd_sc_hd__nor2_4
X_50154_ _86253_/Q _50137_/X _50153_/Y _50154_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_8_105_0_CLK clkbuf_7_52_0_CLK/X clkbuf_9_210_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_85851_ _83310_/CLK _52296_/Y _85851_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_100_0_CLK clkbuf_9_50_0_CLK/X _86878_/CLK sky130_fd_sc_hd__clkbuf_1
X_67997_ _67997_/A _67997_/X sky130_fd_sc_hd__buf_2
X_84802_ _84802_/CLK _84802_/D _84802_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_730_0_CLK clkbuf_9_365_0_CLK/X _87766_/CLK sky130_fd_sc_hd__clkbuf_1
X_57750_ _57726_/X _86014_/Q _57749_/X _57750_/Y sky130_fd_sc_hd__o21ai_4
X_69736_ _73106_/A _69645_/X _69478_/X _69735_/Y _69736_/X sky130_fd_sc_hd__a211o_4
X_50085_ _86267_/Q _50061_/X _50084_/Y _50085_/Y sky130_fd_sc_hd__o21ai_4
X_54962_ _85344_/Q _54249_/X _54961_/Y _54962_/Y sky130_fd_sc_hd__o21ai_4
X_66948_ _66851_/X _66948_/B _66948_/X sky130_fd_sc_hd__and2_4
X_85782_ _82956_/CLK _52640_/Y _85782_/Q sky130_fd_sc_hd__dfxtp_4
X_82994_ _82993_/CLK _74659_/Y _82994_/Q sky130_fd_sc_hd__dfxtp_4
X_56701_ _56700_/Y _83327_/Q _56682_/X _56674_/X _57270_/A _56702_/A
+ sky130_fd_sc_hd__a41o_4
X_87521_ _87525_/CLK _87521_/D _87521_/Q sky130_fd_sc_hd__dfxtp_4
X_53913_ _85543_/Q _53896_/X _53912_/Y _53913_/Y sky130_fd_sc_hd__o21ai_4
X_84733_ _84903_/CLK _59438_/Y _64526_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_221_0_CLK clkbuf_9_220_0_CLK/A clkbuf_9_221_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_57681_ _57677_/X _57678_/Y _57680_/Y _84955_/D sky130_fd_sc_hd__a21oi_4
X_81945_ _82133_/CLK _77946_/Y _81945_/Q sky130_fd_sc_hd__dfxtp_4
X_69667_ _87064_/Q _69664_/X _69665_/X _69666_/X _69668_/B sky130_fd_sc_hd__a211o_4
X_54893_ _54919_/A _54893_/X sky130_fd_sc_hd__buf_2
X_66879_ _66879_/A _66879_/X sky130_fd_sc_hd__buf_2
X_59420_ _59398_/A _59424_/B sky130_fd_sc_hd__buf_2
X_56632_ _56650_/B _55467_/X _55646_/X _56632_/Y sky130_fd_sc_hd__nand3_4
X_68618_ _57804_/A _68618_/B _68618_/Y sky130_fd_sc_hd__nor2_4
X_87452_ _87446_/CLK _87452_/D _87452_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_115_0_CLK clkbuf_9_57_0_CLK/X _84426_/CLK sky130_fd_sc_hd__clkbuf_1
X_53844_ _53844_/A _53844_/B _53844_/Y sky130_fd_sc_hd__nand2_4
X_84664_ _84671_/CLK _84664_/D _60089_/C sky130_fd_sc_hd__dfxtp_4
X_81876_ _81839_/CLK _78067_/X _81876_/Q sky130_fd_sc_hd__dfxtp_4
X_69598_ _87069_/Q _66550_/X _66552_/X _69597_/X _69598_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_745_0_CLK clkbuf_9_372_0_CLK/X _87993_/CLK sky130_fd_sc_hd__clkbuf_1
X_86403_ _86404_/CLK _86403_/D _65381_/B sky130_fd_sc_hd__dfxtp_4
X_83615_ _85562_/CLK _71079_/Y _83615_/Q sky130_fd_sc_hd__dfxtp_4
X_59351_ _72201_/A _59351_/X sky130_fd_sc_hd__buf_2
X_56563_ _56774_/C _56798_/B sky130_fd_sc_hd__buf_2
X_80827_ _81065_/CLK _80827_/D _75650_/B sky130_fd_sc_hd__dfxtp_4
X_68549_ _65381_/A _68549_/B _68549_/X sky130_fd_sc_hd__and2_4
X_87383_ _87189_/CLK _43512_/X _87383_/Q sky130_fd_sc_hd__dfxtp_4
X_53775_ _53771_/Y _53773_/X _53774_/X _53775_/Y sky130_fd_sc_hd__a21oi_4
X_84595_ _84469_/CLK _60582_/Y _79135_/A sky130_fd_sc_hd__dfxtp_4
X_50987_ _50971_/A _50987_/B _50987_/Y sky130_fd_sc_hd__nand2_4
X_58302_ _58282_/X _58298_/Y _58301_/Y _84884_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_236_0_CLK clkbuf_8_118_0_CLK/X clkbuf_9_236_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_55514_ _55507_/X _55514_/B _55514_/Y sky130_fd_sc_hd__nor2_4
X_86334_ _86655_/CLK _86334_/D _86334_/Q sky130_fd_sc_hd__dfxtp_4
X_40740_ _40739_/X _40719_/X _88344_/Q _40720_/X _40740_/X sky130_fd_sc_hd__a2bb2o_4
X_52726_ _52718_/A _52726_/B _52726_/Y sky130_fd_sc_hd__nand2_4
X_59282_ _86666_/Q _59282_/B _59282_/Y sky130_fd_sc_hd__nor2_4
X_71560_ _71557_/X _83457_/Q _71559_/Y _83457_/D sky130_fd_sc_hd__a21o_4
X_83546_ _85354_/CLK _71286_/Y _83546_/Q sky130_fd_sc_hd__dfxtp_4
X_56494_ _56487_/X _56484_/X _56494_/C _56494_/Y sky130_fd_sc_hd__nand3_4
X_80758_ _81134_/CLK _80758_/D _81134_/D sky130_fd_sc_hd__dfxtp_4
X_70511_ _70511_/A _70374_/X _70508_/X _70511_/Y sky130_fd_sc_hd__nand3_4
X_58233_ _83397_/Q _58233_/Y sky130_fd_sc_hd__inv_2
X_55445_ _55445_/A _55445_/B _55445_/C _55445_/D _55446_/A sky130_fd_sc_hd__and4_4
X_86265_ _85562_/CLK _86265_/D _86265_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_601 sky130_fd_sc_hd__decap_3
X_40671_ _40671_/A _40588_/B _40671_/X sky130_fd_sc_hd__or2_4
X_52657_ _52657_/A _52657_/X sky130_fd_sc_hd__buf_2
X_71491_ _71483_/B _71496_/C sky130_fd_sc_hd__buf_2
X_83477_ _83414_/CLK _83477_/D _83477_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_612 sky130_fd_sc_hd__decap_3
X_80689_ _81074_/CLK _80721_/Q _75288_/A sky130_fd_sc_hd__dfxtp_4
XPHY_623 sky130_fd_sc_hd__decap_3
X_88004_ _87249_/CLK _88004_/D _88004_/Q sky130_fd_sc_hd__dfxtp_4
X_42410_ _42397_/A _42410_/X sky130_fd_sc_hd__buf_2
XPHY_634 sky130_fd_sc_hd__decap_3
X_73230_ _73226_/X _73229_/X _73200_/X _73230_/X sky130_fd_sc_hd__a21o_4
X_85216_ _85184_/CLK _56380_/Y _56379_/C sky130_fd_sc_hd__dfxtp_4
X_51608_ _51608_/A _51608_/X sky130_fd_sc_hd__buf_2
X_70442_ _70442_/A _70949_/B _71194_/C _70442_/Y sky130_fd_sc_hd__nand3_4
X_82428_ _82692_/CLK _82428_/D _78691_/A sky130_fd_sc_hd__dfxtp_4
X_58164_ _64257_/A _58160_/B _58164_/Y sky130_fd_sc_hd__nand2_4
XPHY_645 sky130_fd_sc_hd__decap_3
X_43390_ _43367_/X _43375_/X _41442_/X _87446_/Q _43378_/X _43390_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55376_ _55375_/Y _55383_/A sky130_fd_sc_hd__inv_2
X_86196_ _86196_/CLK _50463_/Y _86196_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_656 sky130_fd_sc_hd__decap_3
X_52588_ _52588_/A _52594_/B _51919_/C _51761_/D _52588_/X sky130_fd_sc_hd__and4_4
XPHY_667 sky130_fd_sc_hd__decap_3
XPHY_678 sky130_fd_sc_hd__decap_3
X_57115_ _57109_/X _56619_/X _85080_/Q _57110_/X _85080_/D sky130_fd_sc_hd__a2bb2o_4
X_42341_ _41693_/X _42325_/X _87912_/Q _42326_/X _42341_/X sky130_fd_sc_hd__a2bb2o_4
X_54327_ _54332_/A _52637_/B _54327_/Y sky130_fd_sc_hd__nand2_4
XPHY_689 sky130_fd_sc_hd__decap_3
X_73161_ _72908_/X _85586_/Q _72909_/X _73160_/X _73161_/X sky130_fd_sc_hd__a211o_4
X_85147_ _85057_/CLK _56605_/Y _56604_/B sky130_fd_sc_hd__dfxtp_4
X_51539_ _51539_/A _51539_/X sky130_fd_sc_hd__buf_2
X_58095_ _58599_/A _58095_/X sky130_fd_sc_hd__buf_2
X_70373_ DATA_TO_HASH[6] _70809_/A sky130_fd_sc_hd__buf_2
X_82359_ _82349_/CLK _77208_/X _82359_/Q sky130_fd_sc_hd__dfxtp_4
X_72112_ _74453_/A _72113_/B sky130_fd_sc_hd__buf_2
X_45060_ _45284_/A _45060_/X sky130_fd_sc_hd__buf_2
X_57046_ _56848_/X _56850_/X _56976_/X _57046_/Y sky130_fd_sc_hd__nor3_4
X_42272_ _42259_/A _42272_/X sky130_fd_sc_hd__buf_2
X_54258_ _85475_/Q _54249_/X _54257_/Y _54258_/Y sky130_fd_sc_hd__o21ai_4
X_73092_ _73092_/A _73092_/X sky130_fd_sc_hd__buf_2
X_85078_ _85083_/CLK _85078_/D _85078_/Q sky130_fd_sc_hd__dfxtp_4
X_44011_ _44152_/A _44024_/A sky130_fd_sc_hd__inv_2
X_41223_ _41223_/A _41223_/B _41223_/X sky130_fd_sc_hd__or2_4
X_53209_ _53219_/A _53209_/B _53209_/Y sky130_fd_sc_hd__nand2_4
X_72043_ _74453_/A _72043_/X sky130_fd_sc_hd__buf_2
X_76920_ _76906_/Y _76934_/A _76920_/Y sky130_fd_sc_hd__nor2_4
X_84029_ _81160_/CLK _84029_/D _82069_/D sky130_fd_sc_hd__dfxtp_4
X_54189_ _85487_/Q _54167_/X _54188_/Y _54189_/Y sky130_fd_sc_hd__o21ai_4
X_41154_ _41151_/X _41152_/X _68549_/B _41153_/X _41154_/X sky130_fd_sc_hd__a2bb2o_4
X_76851_ _76829_/A _76828_/Y _76841_/A _76840_/Y _76851_/X sky130_fd_sc_hd__o22a_4
X_58997_ _58997_/A _58898_/B _58997_/Y sky130_fd_sc_hd__nor2_4
X_75802_ _75796_/Y _75802_/B _75803_/C sky130_fd_sc_hd__nand2_4
X_48750_ _48737_/A _52137_/B _48750_/Y sky130_fd_sc_hd__nand2_4
X_79570_ _65348_/C _83253_/Q _79571_/A sky130_fd_sc_hd__nor2_4
X_45962_ _51337_/A _45962_/X sky130_fd_sc_hd__buf_2
X_41085_ _41085_/A _41079_/X _41085_/X sky130_fd_sc_hd__or2_4
X_57948_ _58126_/A _57948_/X sky130_fd_sc_hd__buf_2
X_76782_ _76774_/X _76781_/Y _76783_/B sky130_fd_sc_hd__xor2_4
X_73994_ _72894_/X _86223_/Q _45896_/X _73993_/X _73994_/X sky130_fd_sc_hd__a211o_4
X_47701_ _47701_/A _53196_/D sky130_fd_sc_hd__buf_2
X_78521_ _78501_/Y _78505_/B _78503_/Y _78521_/X sky130_fd_sc_hd__o21a_4
X_44913_ _56196_/C _44911_/X _44912_/X _44913_/Y sky130_fd_sc_hd__o21ai_4
X_75733_ _81092_/Q _75733_/B _75733_/Y sky130_fd_sc_hd__xnor2_4
X_87719_ _88232_/CLK _42786_/X _67613_/B sky130_fd_sc_hd__dfxtp_4
X_48681_ _48674_/Y _48651_/X _48680_/X _48681_/Y sky130_fd_sc_hd__a21oi_4
X_72945_ _72945_/A _73000_/B _72945_/Y sky130_fd_sc_hd__nor2_4
X_45893_ _41869_/A _45893_/B _45893_/C _45893_/Y sky130_fd_sc_hd__nor3_4
X_57879_ _57852_/X _85719_/Q _57878_/X _57879_/X sky130_fd_sc_hd__o21a_4
X_47632_ _47632_/A _53157_/B sky130_fd_sc_hd__buf_2
X_59618_ _59905_/B _61294_/D sky130_fd_sc_hd__inv_2
X_78452_ _78429_/Y _78450_/Y _78451_/Y _78453_/B sky130_fd_sc_hd__a21oi_4
X_44844_ _46001_/A _44844_/X sky130_fd_sc_hd__buf_2
X_75664_ _75649_/A _75661_/Y _75663_/X _75665_/B sky130_fd_sc_hd__o21ai_4
X_72876_ _44131_/A _72877_/A sky130_fd_sc_hd__buf_2
X_60890_ _64191_/B _60997_/A _60888_/Y _60889_/X _60890_/X sky130_fd_sc_hd__and4_4
X_77403_ _77434_/B _77403_/B _82190_/D sky130_fd_sc_hd__xnor2_4
X_74615_ _74605_/X _74613_/X _56148_/A _74614_/X _74615_/X sky130_fd_sc_hd__a211o_4
X_47563_ _47553_/A _53122_/B _47563_/Y sky130_fd_sc_hd__nand2_4
X_71827_ _71827_/A _71716_/B _70763_/A _71826_/X _71827_/X sky130_fd_sc_hd__and4_4
X_59549_ _59609_/D _59581_/C sky130_fd_sc_hd__buf_2
X_78383_ _78383_/A _82759_/D _82471_/D sky130_fd_sc_hd__xor2_4
X_44775_ _44650_/A _44775_/X sky130_fd_sc_hd__buf_2
X_75595_ _75595_/A _75594_/Y _75596_/B sky130_fd_sc_hd__nand2_4
X_41987_ _41982_/X _41975_/X _40776_/X _41986_/Y _41984_/X _41987_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49302_ _49302_/A _51328_/B _49302_/Y sky130_fd_sc_hd__nand2_4
X_46514_ _82922_/Q _46459_/B _46514_/X sky130_fd_sc_hd__or2_4
X_77334_ _77334_/A _77334_/B _77334_/Y sky130_fd_sc_hd__nor2_4
X_43726_ _43726_/A _43726_/Y sky130_fd_sc_hd__inv_2
X_62560_ _61618_/X _62560_/B _62560_/C _62560_/D _62560_/Y sky130_fd_sc_hd__nand4_4
X_74546_ _56016_/A _74538_/Y _74545_/Y _74546_/Y sky130_fd_sc_hd__o21ai_4
X_40938_ _40504_/X _82304_/Q _40937_/X _40938_/Y sky130_fd_sc_hd__o21ai_4
X_47494_ _47494_/A _53078_/D sky130_fd_sc_hd__buf_2
X_71758_ _71041_/X _70635_/A _71755_/X _71753_/D _71758_/Y sky130_fd_sc_hd__nand4_4
X_61511_ _61482_/A _61510_/X _61482_/C _61511_/Y sky130_fd_sc_hd__nand3_4
X_49233_ _64749_/B _49204_/X _49232_/Y _49233_/Y sky130_fd_sc_hd__o21ai_4
X_70709_ _52748_/B _70699_/X _70708_/Y _70709_/Y sky130_fd_sc_hd__o21ai_4
X_46445_ _72083_/A _46445_/X sky130_fd_sc_hd__buf_2
X_77265_ _77265_/A _77265_/B _77265_/Y sky130_fd_sc_hd__nand2_4
X_43657_ _43607_/A _43657_/X sky130_fd_sc_hd__buf_2
X_62491_ _62533_/A _58483_/A _62491_/C _62493_/C sky130_fd_sc_hd__nand3_4
X_74477_ _83058_/Q _74474_/X _74476_/Y _74477_/Y sky130_fd_sc_hd__o21ai_4
X_40869_ _40869_/A _40869_/Y sky130_fd_sc_hd__inv_2
X_71689_ _71682_/Y _83410_/Q _71688_/Y _83410_/D sky130_fd_sc_hd__a21o_4
X_79004_ _79002_/Y _79003_/Y _79022_/A sky130_fd_sc_hd__xor2_4
X_64230_ _64222_/X _64223_/X _64225_/X _64228_/Y _64229_/X _64230_/X
+ sky130_fd_sc_hd__o41a_4
X_76216_ _81255_/Q _81511_/D _76216_/Y sky130_fd_sc_hd__nand2_4
X_42608_ _73394_/A _69897_/B sky130_fd_sc_hd__inv_2
X_49164_ _49080_/A _53919_/B _49164_/X sky130_fd_sc_hd__and2_4
X_61442_ _59392_/A _61452_/B _61452_/C _61452_/D _61442_/Y sky130_fd_sc_hd__nand4_4
X_73428_ _73425_/X _73427_/X _72949_/X _73428_/X sky130_fd_sc_hd__a21o_4
X_46376_ _83646_/Q _46376_/Y sky130_fd_sc_hd__inv_2
X_77196_ _82012_/Q _82300_/D _77196_/Y sky130_fd_sc_hd__nand2_4
X_43588_ _42447_/A _41869_/B _42447_/B _42447_/D _43588_/X sky130_fd_sc_hd__and4_4
X_48115_ _53593_/B _50370_/B sky130_fd_sc_hd__buf_2
X_45327_ _55732_/B _45284_/X _45265_/X _45327_/X sky130_fd_sc_hd__o21a_4
X_64161_ _61665_/B _64161_/B _64172_/C _64161_/D _64161_/Y sky130_fd_sc_hd__nand4_4
X_76147_ _76149_/C _76147_/Y sky130_fd_sc_hd__inv_2
X_42539_ _42536_/X _42527_/X _40753_/X _69089_/B _42538_/X _87829_/D
+ sky130_fd_sc_hd__o32ai_4
X_61373_ _61290_/X _61374_/A sky130_fd_sc_hd__buf_2
X_49095_ _49056_/A _52367_/B _49095_/Y sky130_fd_sc_hd__nand2_4
X_73359_ _73359_/A _73359_/X sky130_fd_sc_hd__buf_2
X_63112_ _63053_/A _63113_/B sky130_fd_sc_hd__buf_2
X_48046_ _48046_/A _52039_/A sky130_fd_sc_hd__buf_2
X_60324_ _60324_/A _60324_/B _60324_/C _60367_/D sky130_fd_sc_hd__nand3_4
X_45258_ _45257_/Y _45199_/B _45258_/Y sky130_fd_sc_hd__nand2_4
X_64092_ _64466_/B _64145_/B _64029_/C _64029_/D _64094_/C sky130_fd_sc_hd__nand4_4
X_76078_ _81719_/D _76070_/B _76078_/Y sky130_fd_sc_hd__nor2_4
X_44209_ _44153_/X _45950_/A sky130_fd_sc_hd__buf_2
X_67920_ _87143_/Q _67825_/X _67872_/X _67919_/X _67920_/X sky130_fd_sc_hd__a211o_4
X_63043_ _60489_/X _63081_/C sky130_fd_sc_hd__buf_2
X_75029_ _75042_/A _75042_/B _75047_/A sky130_fd_sc_hd__xor2_4
X_79906_ _79908_/B _79906_/Y sky130_fd_sc_hd__inv_2
X_60255_ _60255_/A _60255_/B _60324_/B _60325_/C sky130_fd_sc_hd__nand3_4
X_45189_ _45265_/A _45189_/X sky130_fd_sc_hd__buf_2
X_67851_ _67782_/X _67842_/Y _67747_/X _67850_/Y _67851_/X sky130_fd_sc_hd__a211o_4
X_79837_ _79837_/A _79837_/B _79838_/B sky130_fd_sc_hd__xor2_4
X_60186_ _60185_/X _60166_/X _60187_/A sky130_fd_sc_hd__and2_4
X_49997_ _50001_/A _53209_/B _49997_/Y sky130_fd_sc_hd__nand2_4
X_66802_ _66728_/A _66802_/B _66802_/X sky130_fd_sc_hd__and2_4
X_48948_ _48946_/X _48426_/Y _48947_/Y _52295_/B sky130_fd_sc_hd__a21o_4
X_67782_ _67495_/X _67782_/X sky130_fd_sc_hd__buf_2
X_79768_ _79740_/X _79743_/Y _79757_/A _79756_/Y _79768_/X sky130_fd_sc_hd__o22a_4
X_64994_ _64990_/X _64888_/B _64993_/X _64994_/Y sky130_fd_sc_hd__nand3_4
X_69521_ _69605_/A _69521_/B _69521_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_1002_0_CLK clkbuf_9_501_0_CLK/X _86203_/CLK sky130_fd_sc_hd__clkbuf_1
X_66733_ _59816_/A _66971_/A sky130_fd_sc_hd__buf_2
X_78719_ _78717_/X _78718_/Y _78720_/A sky130_fd_sc_hd__and2_4
X_63945_ _63943_/X _63913_/X _63944_/Y _84285_/D sky130_fd_sc_hd__a21oi_4
X_48879_ _86465_/Q _48669_/X _48878_/Y _48879_/Y sky130_fd_sc_hd__o21ai_4
X_79699_ _84216_/Q _72323_/A _79699_/X sky130_fd_sc_hd__xor2_4
X_50910_ _50819_/X _50910_/X sky130_fd_sc_hd__buf_2
X_81730_ _80928_/CLK _75925_/B _41452_/A sky130_fd_sc_hd__dfxtp_4
X_69452_ _69286_/A _69452_/B _69452_/X sky130_fd_sc_hd__and2_4
X_66664_ _68614_/A _66664_/X sky130_fd_sc_hd__buf_2
X_51890_ _85927_/Q _51873_/X _51889_/Y _51890_/Y sky130_fd_sc_hd__o21ai_4
X_63876_ _61861_/X _63876_/B _63860_/C _63860_/D _63876_/Y sky130_fd_sc_hd__nand4_4
X_68403_ _68403_/A _68403_/B _68403_/X sky130_fd_sc_hd__and2_4
X_65615_ _65610_/X _65613_/X _65614_/X _65615_/X sky130_fd_sc_hd__a21o_4
X_50841_ _50837_/Y _50839_/X _50840_/X _86123_/D sky130_fd_sc_hd__a21oi_4
X_62827_ _60288_/C _62827_/X sky130_fd_sc_hd__buf_2
X_81661_ _81680_/CLK _81693_/Q _81661_/Q sky130_fd_sc_hd__dfxtp_4
X_69383_ _69383_/A _87265_/Q _69383_/X sky130_fd_sc_hd__and2_4
X_66595_ _69853_/A _88210_/Q _66595_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_1017_0_CLK clkbuf_9_508_0_CLK/X _86193_/CLK sky130_fd_sc_hd__clkbuf_1
X_83400_ _84939_/CLK _83400_/D _83400_/Q sky130_fd_sc_hd__dfxtp_4
X_80612_ _80606_/A _80606_/B _80611_/Y _80623_/A sky130_fd_sc_hd__a21boi_4
X_68334_ _82628_/D _68318_/X _68333_/X _83980_/D sky130_fd_sc_hd__a21bo_4
X_53560_ _50724_/A _53620_/B sky130_fd_sc_hd__buf_2
X_65546_ _65559_/A _65546_/B _65546_/C _65546_/X sky130_fd_sc_hd__and3_4
X_84380_ _84375_/CLK _62817_/Y _62816_/C sky130_fd_sc_hd__dfxtp_4
X_50772_ _86136_/Q _50742_/X _50771_/Y _50772_/Y sky130_fd_sc_hd__o21ai_4
X_62758_ _62756_/X _62721_/X _62757_/Y _62758_/Y sky130_fd_sc_hd__a21oi_4
X_81592_ _81428_/CLK _84192_/Q _76855_/A sky130_fd_sc_hd__dfxtp_4
X_52511_ _52501_/X _46455_/Y _52511_/Y sky130_fd_sc_hd__nand2_4
X_83331_ _83337_/CLK _83331_/D _83331_/Q sky130_fd_sc_hd__dfxtp_4
X_61709_ _61708_/X _62187_/C sky130_fd_sc_hd__buf_2
X_80543_ _80529_/Y _80534_/Y _80542_/X _80544_/B sky130_fd_sc_hd__o21ai_4
X_68265_ _68246_/X _67623_/Y _68247_/X _68264_/Y _68265_/X sky130_fd_sc_hd__a211o_4
X_53491_ _85626_/Q _53466_/X _53490_/Y _53491_/Y sky130_fd_sc_hd__o21ai_4
X_65477_ _65473_/X _65477_/B _65477_/Y sky130_fd_sc_hd__nand2_4
X_62689_ _60217_/A _62689_/X sky130_fd_sc_hd__buf_2
X_55230_ _85092_/Q _55142_/A _55133_/X _55229_/X _55230_/X sky130_fd_sc_hd__a211o_4
X_67216_ _87352_/Q _67121_/X _67122_/X _67215_/X _67216_/X sky130_fd_sc_hd__a211o_4
X_86050_ _83690_/CLK _86050_/D _86050_/Q sky130_fd_sc_hd__dfxtp_4
X_52442_ _52436_/A _53959_/B _52442_/Y sky130_fd_sc_hd__nand2_4
X_64428_ _79691_/B _64373_/X _64427_/X _84247_/D sky130_fd_sc_hd__a21o_4
X_83262_ _86289_/CLK _83262_/D _83262_/Q sky130_fd_sc_hd__dfxtp_4
X_80474_ _84763_/Q _80481_/B _80476_/A sky130_fd_sc_hd__xor2_4
X_68196_ _68097_/A _68196_/X sky130_fd_sc_hd__buf_2
X_85001_ _83335_/CLK _85001_/D _85001_/Q sky130_fd_sc_hd__dfxtp_4
X_82213_ _82220_/CLK _82245_/Q _82213_/Q sky130_fd_sc_hd__dfxtp_4
X_55161_ _55156_/X _83746_/Q _55160_/X _55296_/B sky130_fd_sc_hd__nand3_4
X_67147_ _67025_/X _67147_/X sky130_fd_sc_hd__buf_2
X_52373_ _52271_/A _52373_/X sky130_fd_sc_hd__buf_2
X_64359_ _79755_/B _64314_/X _64358_/X _64359_/X sky130_fd_sc_hd__a21o_4
X_83193_ _83191_/CLK _83193_/D _70219_/C sky130_fd_sc_hd__dfxtp_4
X_54112_ _54107_/Y _53437_/X _54111_/X _54112_/Y sky130_fd_sc_hd__a21oi_4
X_51324_ _51310_/X _51324_/B _51324_/Y sky130_fd_sc_hd__nand2_4
X_82144_ _82575_/CLK _82144_/D _77488_/B sky130_fd_sc_hd__dfxtp_4
X_55092_ _55090_/Y _55076_/X _55091_/X _85320_/D sky130_fd_sc_hd__a21oi_4
X_67078_ _67078_/A _67078_/B _67078_/Y sky130_fd_sc_hd__nand2_4
X_58920_ _58920_/A _58920_/B _58920_/Y sky130_fd_sc_hd__nor2_4
X_54043_ _54043_/A _54043_/B _53969_/C _54043_/X sky130_fd_sc_hd__and3_4
X_66029_ _65824_/X _84985_/Q _66027_/X _66028_/X _66029_/X sky130_fd_sc_hd__a211o_4
X_51255_ _48853_/A _51330_/C sky130_fd_sc_hd__buf_2
X_86952_ _88220_/CLK _86952_/D _86952_/Q sky130_fd_sc_hd__dfxtp_4
X_82075_ _81160_/CLK _84035_/Q _77952_/A sky130_fd_sc_hd__dfxtp_4
X_50206_ _50204_/Y _50191_/X _50205_/X _50206_/Y sky130_fd_sc_hd__a21oi_4
X_81026_ _85317_/CLK _81026_/D _81026_/Q sky130_fd_sc_hd__dfxtp_4
X_85903_ _86576_/CLK _52030_/Y _66166_/B sky130_fd_sc_hd__dfxtp_4
X_58851_ _58763_/A _86379_/Q _58851_/Y sky130_fd_sc_hd__nor2_4
X_51186_ _86058_/Q _51183_/X _51185_/Y _51186_/Y sky130_fd_sc_hd__o21ai_4
X_86883_ _86869_/CLK _45336_/Y _64524_/B sky130_fd_sc_hd__dfxtp_4
X_57802_ _44147_/A _57803_/A sky130_fd_sc_hd__buf_2
X_50137_ _50113_/A _50137_/X sky130_fd_sc_hd__buf_2
X_85834_ _86155_/CLK _85834_/D _85834_/Q sky130_fd_sc_hd__dfxtp_4
X_58782_ _58730_/X _85936_/Q _58679_/X _58782_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_9_160_0_CLK clkbuf_8_80_0_CLK/X clkbuf_9_160_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_55994_ _55828_/X _55994_/X sky130_fd_sc_hd__buf_2
X_57733_ _59286_/A _57833_/B sky130_fd_sc_hd__buf_2
X_69719_ _68587_/X _69719_/B _69719_/Y sky130_fd_sc_hd__nor2_4
X_50068_ _50092_/A _50068_/X sky130_fd_sc_hd__buf_2
X_54945_ _85348_/Q _53449_/X _54944_/Y _54945_/Y sky130_fd_sc_hd__o21ai_4
X_85765_ _85767_/CLK _52731_/Y _85765_/Q sky130_fd_sc_hd__dfxtp_4
X_70991_ _51320_/B _70983_/X _70990_/Y _83640_/D sky130_fd_sc_hd__o21ai_4
X_82977_ _83783_/CLK _82785_/Q _82977_/Q sky130_fd_sc_hd__dfxtp_4
X_87504_ _87766_/CLK _43276_/X _87504_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_684_0_CLK clkbuf_9_342_0_CLK/X _87644_/CLK sky130_fd_sc_hd__clkbuf_1
X_41910_ _41909_/Y _41911_/A sky130_fd_sc_hd__buf_2
X_72730_ _73163_/A _72730_/X sky130_fd_sc_hd__buf_2
X_84716_ _84716_/CLK _84716_/D _64276_/C sky130_fd_sc_hd__dfxtp_4
X_57664_ _57664_/A _57664_/X sky130_fd_sc_hd__buf_2
X_81928_ _81928_/CLK _81928_/D _81928_/Q sky130_fd_sc_hd__dfxtp_4
X_42890_ _42889_/Y _42890_/Y sky130_fd_sc_hd__inv_2
X_54876_ _54885_/A _47679_/A _54876_/Y sky130_fd_sc_hd__nand2_4
X_85696_ _85697_/CLK _85696_/D _85696_/Q sky130_fd_sc_hd__dfxtp_4
X_59403_ _59403_/A _59399_/B _59403_/Y sky130_fd_sc_hd__nand2_4
X_56615_ _56613_/X _56553_/Y _56614_/Y _85145_/D sky130_fd_sc_hd__a21oi_4
X_87435_ _87484_/CLK _87435_/D _87435_/Q sky130_fd_sc_hd__dfxtp_4
X_41841_ _42465_/A _41841_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_175_0_CLK clkbuf_8_87_0_CLK/X clkbuf_9_175_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_53827_ _53786_/A _48973_/A _53827_/Y sky130_fd_sc_hd__nand2_4
X_72661_ _72688_/A _72668_/B sky130_fd_sc_hd__buf_2
X_84647_ _84645_/CLK _60245_/Y _79863_/A sky130_fd_sc_hd__dfxtp_4
X_57595_ _57552_/X _48051_/Y _57595_/Y sky130_fd_sc_hd__nand2_4
X_81859_ _81859_/CLK _81859_/D _81827_/D sky130_fd_sc_hd__dfxtp_4
X_74400_ _71964_/A _74421_/C sky130_fd_sc_hd__buf_2
X_59334_ _59037_/A _59334_/X sky130_fd_sc_hd__buf_2
X_71612_ _71857_/A _70573_/B _71614_/C _71606_/X _71612_/Y sky130_fd_sc_hd__nor4_4
X_56546_ _56546_/A _56545_/Y _85154_/D sky130_fd_sc_hd__nand2_4
X_44560_ _44560_/A _87055_/D sky130_fd_sc_hd__inv_2
X_75380_ _75375_/Y _75377_/Y _75380_/Y sky130_fd_sc_hd__nor2_4
X_87366_ _86824_/CLK _43548_/Y _87366_/Q sky130_fd_sc_hd__dfxtp_4
X_41772_ _40402_/A _81734_/Q _41771_/X _41772_/X sky130_fd_sc_hd__o21a_4
X_53758_ _53733_/A _53774_/B sky130_fd_sc_hd__buf_2
X_84578_ _84458_/CLK _60734_/Y _84578_/Q sky130_fd_sc_hd__dfxtp_4
X_72592_ _72592_/A _61414_/A _79330_/B _72592_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_10_699_0_CLK clkbuf_9_349_0_CLK/X _87952_/CLK sky130_fd_sc_hd__clkbuf_1
X_43511_ _43511_/A _43511_/Y sky130_fd_sc_hd__inv_2
X_86317_ _86317_/CLK _86317_/D _86317_/Q sky130_fd_sc_hd__dfxtp_4
X_74331_ _70315_/C _74327_/X _74330_/Y _83096_/D sky130_fd_sc_hd__a21bo_4
X_40723_ _40698_/X _82857_/Q _40722_/X _40723_/X sky130_fd_sc_hd__o21a_4
X_52709_ _52704_/A _52694_/B _52708_/X _52709_/D _52709_/X sky130_fd_sc_hd__and4_4
X_59265_ _59177_/X _86060_/Q _59264_/X _59265_/Y sky130_fd_sc_hd__o21ai_4
X_83529_ _83526_/CLK _83529_/D _83529_/Q sky130_fd_sc_hd__dfxtp_4
X_71543_ _71531_/X _59457_/B _71542_/Y _83463_/D sky130_fd_sc_hd__a21o_4
X_44491_ _44481_/X _44482_/X _41224_/X _87082_/Q _44484_/X _44491_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56477_ _56474_/X _56472_/B _55949_/B _56477_/Y sky130_fd_sc_hd__nand3_4
X_87297_ _87814_/CLK _43720_/Y _43717_/A sky130_fd_sc_hd__dfxtp_4
X_53689_ _53713_/A _48514_/A _53689_/Y sky130_fd_sc_hd__nand2_4
X_46230_ _45893_/B _42447_/D _45893_/C _46230_/X sky130_fd_sc_hd__or3_4
X_58216_ _84905_/Q _63355_/A sky130_fd_sc_hd__inv_2
XPHY_420 sky130_fd_sc_hd__decap_3
X_77050_ _77050_/A _81906_/Q _77067_/A sky130_fd_sc_hd__xor2_4
X_43442_ _41592_/X _43431_/X _87418_/Q _43432_/X _43442_/X sky130_fd_sc_hd__a2bb2o_4
X_55428_ _55421_/Y _55423_/Y _55428_/C _55427_/Y _55429_/A sky130_fd_sc_hd__nand4_4
X_74262_ _74260_/X _74261_/Y _73982_/X _74262_/X sky130_fd_sc_hd__a21o_4
X_86248_ _86154_/CLK _50180_/Y _65249_/B sky130_fd_sc_hd__dfxtp_4
XPHY_431 sky130_fd_sc_hd__decap_3
X_40654_ _40654_/A _40654_/B _40654_/X sky130_fd_sc_hd__or2_4
X_59196_ _58810_/A _59196_/X sky130_fd_sc_hd__buf_2
X_71474_ _71464_/X _83486_/Q _71473_/X _83486_/D sky130_fd_sc_hd__a21o_4
XPHY_442 sky130_fd_sc_hd__decap_3
XPHY_453 sky130_fd_sc_hd__decap_3
X_76001_ _75994_/Y _76005_/A _76000_/Y _76001_/Y sky130_fd_sc_hd__a21boi_4
X_73213_ _73208_/X _73212_/X _73067_/X _73217_/A sky130_fd_sc_hd__a21o_4
XPHY_464 sky130_fd_sc_hd__decap_3
X_70425_ _70424_/X _70426_/A sky130_fd_sc_hd__buf_2
X_46161_ _46099_/X _74846_/B _46162_/D sky130_fd_sc_hd__nor2_4
Xclkbuf_10_622_0_CLK clkbuf_9_311_0_CLK/X _82335_/CLK sky130_fd_sc_hd__clkbuf_1
X_58147_ _58147_/A _57666_/B _58147_/Y sky130_fd_sc_hd__nor2_4
XPHY_475 sky130_fd_sc_hd__decap_3
X_43373_ _41393_/X _43371_/X _87455_/Q _43372_/X _87455_/D sky130_fd_sc_hd__a2bb2o_4
X_55359_ _55352_/A _55352_/C _55360_/A sky130_fd_sc_hd__and2_4
X_86179_ _86500_/CLK _50553_/Y _86179_/Q sky130_fd_sc_hd__dfxtp_4
X_74193_ _45931_/X _86214_/Q _74103_/X _74192_/X _74193_/X sky130_fd_sc_hd__a211o_4
XPHY_486 sky130_fd_sc_hd__decap_3
X_40585_ _40585_/A _40585_/X sky130_fd_sc_hd__buf_2
XPHY_497 sky130_fd_sc_hd__decap_3
X_45112_ _45105_/X _45109_/Y _45111_/Y _45112_/Y sky130_fd_sc_hd__a21oi_4
X_42324_ _41643_/X _42303_/X _87921_/Q _42305_/X _87921_/D sky130_fd_sc_hd__a2bb2o_4
X_73144_ _73142_/X _73143_/Y _72970_/X _73144_/Y sky130_fd_sc_hd__a21oi_4
X_46092_ _80656_/Q _46092_/X sky130_fd_sc_hd__buf_2
X_58078_ _84927_/Q _58025_/X _58072_/X _58077_/X _84927_/D sky130_fd_sc_hd__a2bb2oi_4
X_70356_ HASH_ADDR[2] _70356_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_9_113_0_CLK clkbuf_8_56_0_CLK/X clkbuf_9_113_0_CLK/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_9_40_0_CLK clkbuf_8_20_0_CLK/X clkbuf_9_40_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_49920_ _49904_/A _49915_/X _49904_/C _53133_/D _49920_/X sky130_fd_sc_hd__and4_4
X_45043_ _45039_/Y _45042_/Y _44986_/X _45043_/X sky130_fd_sc_hd__a21o_4
X_57029_ _57029_/A _57043_/B _56812_/X _57029_/Y sky130_fd_sc_hd__nand3_4
X_42255_ _41447_/X _42248_/X _87957_/Q _42249_/X _87957_/D sky130_fd_sc_hd__a2bb2o_4
X_73075_ _73073_/X _73058_/X _73075_/C _73075_/Y sky130_fd_sc_hd__nand3_4
X_77952_ _77952_/A _77954_/A sky130_fd_sc_hd__inv_2
X_70287_ _70292_/A _70292_/B _83106_/Q _70292_/D _70287_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_637_0_CLK clkbuf_9_318_0_CLK/X _82008_/CLK sky130_fd_sc_hd__clkbuf_1
X_41206_ _40946_/A _41206_/X sky130_fd_sc_hd__buf_2
X_72026_ _72023_/Y _72009_/X _72025_/Y _72026_/Y sky130_fd_sc_hd__a21boi_4
X_76903_ _76904_/A _76902_/B _81597_/Q _76905_/A sky130_fd_sc_hd__a21o_4
X_60040_ _64689_/A _72604_/B _80153_/A _60038_/Y _60049_/A _60041_/A
+ sky130_fd_sc_hd__o32ai_4
X_49851_ _49851_/A _49851_/B _49862_/C _53063_/D _49851_/X sky130_fd_sc_hd__and4_4
X_42186_ _41268_/X _42183_/X _87991_/Q _42184_/X _87991_/D sky130_fd_sc_hd__a2bb2o_4
X_77883_ _82243_/Q _77883_/B _77883_/Y sky130_fd_sc_hd__xnor2_4
X_48802_ _48800_/Y _48785_/X _48801_/X _48802_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_128_0_CLK clkbuf_8_64_0_CLK/X clkbuf_9_128_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_79622_ _79611_/A _79594_/Y _79611_/B _79622_/Y sky130_fd_sc_hd__a21boi_4
X_41137_ _81724_/Q _41079_/X _41137_/X sky130_fd_sc_hd__or2_4
X_76834_ _76822_/A _76821_/Y _76810_/A _81364_/D _76834_/X sky130_fd_sc_hd__a2bb2o_4
X_49782_ _57918_/B _49768_/X _49781_/Y _49782_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_55_0_CLK clkbuf_9_55_0_CLK/A clkbuf_9_55_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_46994_ _53309_/B _52794_/B sky130_fd_sc_hd__buf_2
X_48733_ _65489_/B _48730_/X _48732_/Y _48733_/Y sky130_fd_sc_hd__o21ai_4
X_79553_ _79553_/A _79554_/A sky130_fd_sc_hd__inv_2
X_45945_ _60150_/A _66517_/B sky130_fd_sc_hd__buf_2
X_41068_ _40937_/A _41068_/B _41068_/X sky130_fd_sc_hd__or2_4
X_76765_ _81487_/Q _76765_/Y sky130_fd_sc_hd__inv_2
X_61991_ _61962_/X _61945_/X _58474_/A _61947_/D _61991_/X sky130_fd_sc_hd__and4_4
X_73977_ _73907_/X _84976_/Q _73859_/X _73976_/X _73977_/X sky130_fd_sc_hd__a211o_4
X_78504_ _78503_/Y _78505_/C sky130_fd_sc_hd__inv_2
X_63730_ _84721_/Q _64191_/B _63731_/D _64190_/D _63730_/Y sky130_fd_sc_hd__nand4_4
X_75716_ _75696_/X _75711_/A _75716_/X sky130_fd_sc_hd__and2_4
X_48664_ _48664_/A _48632_/B _48664_/Y sky130_fd_sc_hd__nand2_4
X_60942_ _61003_/A _64067_/A sky130_fd_sc_hd__buf_2
X_72928_ _44531_/Y _72775_/X _72927_/Y _72928_/X sky130_fd_sc_hd__a21o_4
X_79484_ _79484_/A _79484_/B _79486_/B sky130_fd_sc_hd__or2_4
X_45876_ _45876_/A _45876_/B _45876_/Y sky130_fd_sc_hd__nand2_4
X_76696_ _81688_/Q _76696_/B _76696_/X sky130_fd_sc_hd__xor2_4
X_47615_ _81240_/Q _47616_/A sky130_fd_sc_hd__inv_2
X_78435_ _78417_/A _82710_/Q _78435_/Y sky130_fd_sc_hd__nand2_4
X_44827_ _44807_/X _44821_/X _41687_/X _86933_/Q _44808_/X _44827_/Y
+ sky130_fd_sc_hd__o32ai_4
X_63661_ _58348_/A _63600_/X _63661_/C _63661_/D _63661_/Y sky130_fd_sc_hd__nand4_4
X_75647_ _75659_/A _75660_/A _75648_/B sky130_fd_sc_hd__xor2_4
X_60873_ _61003_/A _64172_/B sky130_fd_sc_hd__buf_2
X_48595_ _73310_/B _48548_/X _48594_/Y _48595_/Y sky130_fd_sc_hd__o21ai_4
X_72859_ _72859_/A _74095_/B _72859_/Y sky130_fd_sc_hd__nor2_4
X_65400_ _65400_/A _65400_/X sky130_fd_sc_hd__buf_2
X_62612_ _62632_/A _63694_/B _62632_/C _62612_/Y sky130_fd_sc_hd__nand3_4
X_47546_ _86623_/Q _47524_/X _47545_/Y _47546_/Y sky130_fd_sc_hd__o21ai_4
X_66380_ _66376_/Y _66377_/X _66379_/X _84134_/D sky130_fd_sc_hd__a21o_4
X_78366_ _78363_/Y _78365_/Y _78369_/A sky130_fd_sc_hd__nor2_4
X_44758_ _41311_/Y _44754_/X _86970_/Q _44755_/X _86970_/D sky130_fd_sc_hd__a2bb2o_4
X_63592_ _63615_/A _63615_/B _84311_/Q _63592_/Y sky130_fd_sc_hd__nor3_4
X_75578_ _75577_/Y _81107_/Q _75888_/A sky130_fd_sc_hd__nand2_4
X_65331_ _65408_/A _86437_/Q _65331_/X sky130_fd_sc_hd__and2_4
X_77317_ _77317_/A _77317_/X sky130_fd_sc_hd__buf_2
X_43709_ _40845_/X _43695_/X _73149_/A _43696_/X _43709_/X sky130_fd_sc_hd__a2bb2o_4
X_62543_ _62556_/A _61611_/A _59977_/A _62548_/D _62543_/X sky130_fd_sc_hd__and4_4
X_74529_ _74529_/A _74531_/B _74531_/C _74531_/D _74529_/Y sky130_fd_sc_hd__nand4_4
X_47477_ _47003_/A _47619_/A sky130_fd_sc_hd__buf_2
X_78297_ _78295_/Y _78291_/Y _78296_/Y _78298_/B sky130_fd_sc_hd__o21ai_4
X_44689_ _44533_/A _44689_/X sky130_fd_sc_hd__buf_2
X_49216_ _49220_/A _53949_/B _49216_/Y sky130_fd_sc_hd__nand2_4
X_68050_ _68479_/A _68403_/A sky130_fd_sc_hd__buf_2
X_46428_ _50802_/A _46428_/B _46428_/C _46428_/X sky130_fd_sc_hd__and3_4
X_65262_ _65259_/X _65261_/X _65161_/X _65262_/X sky130_fd_sc_hd__a21o_4
X_77248_ _81923_/Q _82179_/D _81891_/D sky130_fd_sc_hd__xor2_4
X_62474_ _62533_/A _58478_/A _62491_/C _62477_/C sky130_fd_sc_hd__nand3_4
X_67001_ _66996_/X _67000_/X _66905_/X _67001_/X sky130_fd_sc_hd__a21o_4
X_64213_ _64457_/C _64213_/X sky130_fd_sc_hd__buf_2
X_49147_ _46349_/A _49161_/B sky130_fd_sc_hd__buf_2
X_61425_ _61434_/A _61434_/B _79150_/B _61425_/Y sky130_fd_sc_hd__nor3_4
X_46359_ _82936_/Q _46380_/B _46359_/X sky130_fd_sc_hd__or2_4
X_65193_ _65181_/Y _65192_/Y _65193_/Y sky130_fd_sc_hd__nand2_4
X_77179_ _82011_/Q _82299_/D _77184_/A sky130_fd_sc_hd__xor2_4
X_64144_ _63672_/B _64190_/B _64178_/C _64091_/D _64144_/Y sky130_fd_sc_hd__nand4_4
X_49078_ _49018_/X _48576_/A _49077_/Y _49079_/A sky130_fd_sc_hd__a21o_4
X_61356_ _84855_/Q _61356_/X sky130_fd_sc_hd__buf_2
X_80190_ _80173_/Y _80176_/Y _80189_/Y _80190_/X sky130_fd_sc_hd__o21a_4
X_48029_ _48025_/Y _48007_/X _48028_/X _48029_/Y sky130_fd_sc_hd__a21oi_4
X_60307_ _60305_/Y _60306_/Y _60286_/X _79764_/A _59814_/X _60307_/X
+ sky130_fd_sc_hd__o32a_4
X_68952_ _68929_/X _68940_/Y _68824_/X _68951_/Y _68952_/X sky130_fd_sc_hd__a211o_4
X_64075_ _64072_/X _64073_/X _64074_/Y _64075_/Y sky130_fd_sc_hd__a21oi_4
X_61287_ _61287_/A _61284_/Y _72621_/B _61287_/D _61306_/A sky130_fd_sc_hd__nand4_4
X_51040_ _51013_/A _51045_/B sky130_fd_sc_hd__buf_2
X_67903_ _67955_/A _87195_/Q _67903_/X sky130_fd_sc_hd__and2_4
X_63026_ _60562_/B _64235_/B _63347_/C _60541_/B _63026_/X sky130_fd_sc_hd__and4_4
X_60238_ _60233_/Y _60324_/A _60259_/B _60350_/A _60238_/Y sky130_fd_sc_hd__a22oi_4
X_68883_ _68377_/A _68883_/X sky130_fd_sc_hd__buf_2
X_82900_ _82284_/CLK _78211_/B _82900_/Q sky130_fd_sc_hd__dfxtp_4
X_67834_ _68640_/A _67834_/X sky130_fd_sc_hd__buf_2
X_60169_ _60239_/A _60170_/A sky130_fd_sc_hd__inv_2
X_83880_ _82557_/CLK _69983_/X _82560_/D sky130_fd_sc_hd__dfxtp_4
X_82831_ _84119_/CLK _82831_/D _82831_/Q sky130_fd_sc_hd__dfxtp_4
X_67765_ _87457_/Q _67717_/X _67718_/X _67764_/X _67765_/X sky130_fd_sc_hd__a211o_4
X_52991_ _52999_/A _52991_/B _52991_/Y sky130_fd_sc_hd__nand2_4
X_64977_ _44149_/X _85523_/Q _64571_/X _64976_/X _64977_/X sky130_fd_sc_hd__a211o_4
X_69504_ _69696_/A _69504_/X sky130_fd_sc_hd__buf_2
X_54730_ _54321_/A _54758_/A sky130_fd_sc_hd__buf_2
X_66716_ _64706_/A _66717_/A sky130_fd_sc_hd__buf_2
X_85550_ _85535_/CLK _85550_/D _85550_/Q sky130_fd_sc_hd__dfxtp_4
X_51942_ _51940_/Y _51934_/X _51941_/Y _51942_/Y sky130_fd_sc_hd__a21boi_4
X_63928_ _63644_/A _63960_/A sky130_fd_sc_hd__buf_2
X_82762_ _82768_/CLK _82762_/D _82954_/D sky130_fd_sc_hd__dfxtp_4
X_67696_ _67696_/A _88164_/Q _67696_/X sky130_fd_sc_hd__and2_4
X_84501_ _84501_/CLK _84501_/D _75903_/A sky130_fd_sc_hd__dfxtp_4
X_81713_ _81749_/CLK _81713_/D _81713_/Q sky130_fd_sc_hd__dfxtp_4
X_69435_ _68900_/X _68903_/X _69418_/X _69435_/Y sky130_fd_sc_hd__a21oi_4
X_54661_ _85401_/Q _54648_/X _54660_/Y _54661_/Y sky130_fd_sc_hd__o21ai_4
X_66647_ _66647_/A _66669_/A sky130_fd_sc_hd__buf_2
X_85481_ _84926_/CLK _85481_/D _85481_/Q sky130_fd_sc_hd__dfxtp_4
X_51873_ _51900_/A _51873_/X sky130_fd_sc_hd__buf_2
X_63859_ _63853_/Y _63859_/B _63857_/Y _63859_/D _63859_/X sky130_fd_sc_hd__and4_4
X_82693_ _82923_/CLK _78838_/X _82681_/D sky130_fd_sc_hd__dfxtp_4
X_56400_ _56372_/X _56050_/X _56399_/Y _85209_/D sky130_fd_sc_hd__o21ai_4
X_87220_ _87141_/CLK _43881_/X _69125_/B sky130_fd_sc_hd__dfxtp_4
X_53612_ _53611_/X _48153_/A _53612_/Y sky130_fd_sc_hd__nand2_4
X_84432_ _84430_/CLK _84432_/D _62122_/C sky130_fd_sc_hd__dfxtp_4
X_50824_ _50724_/A _50825_/B sky130_fd_sc_hd__buf_2
X_57380_ _57379_/Y _57380_/X sky130_fd_sc_hd__buf_2
X_81644_ _81620_/CLK _81676_/Q _81644_/Q sky130_fd_sc_hd__dfxtp_4
X_69366_ _81393_/D _69299_/X _69365_/X _83929_/D sky130_fd_sc_hd__a21bo_4
X_54592_ _54588_/Y _54584_/X _54591_/X _85414_/D sky130_fd_sc_hd__a21oi_4
X_66578_ _87379_/Q _66571_/X _66574_/X _66577_/X _66578_/X sky130_fd_sc_hd__a211o_4
X_56331_ _56368_/A _56094_/X _56330_/Y _85233_/D sky130_fd_sc_hd__o21ai_4
X_68317_ _82632_/D _68299_/X _68316_/X _83984_/D sky130_fd_sc_hd__a21bo_4
X_87151_ _87150_/CLK _87151_/D _87151_/Q sky130_fd_sc_hd__dfxtp_4
X_53543_ _85616_/Q _53540_/X _53542_/Y _53543_/Y sky130_fd_sc_hd__o21ai_4
X_65529_ _65529_/A _65529_/X sky130_fd_sc_hd__buf_2
X_84363_ _84559_/CLK _62989_/Y _62988_/C sky130_fd_sc_hd__dfxtp_4
X_50755_ _50755_/A _50751_/B _50751_/C _50755_/X sky130_fd_sc_hd__and3_4
X_81575_ _81575_/CLK _84175_/Q _76695_/A sky130_fd_sc_hd__dfxtp_4
X_69297_ _69216_/X _69293_/Y _69231_/X _69296_/Y _69297_/X sky130_fd_sc_hd__a211o_4
X_86102_ _82956_/CLK _50949_/Y _86102_/Q sky130_fd_sc_hd__dfxtp_4
X_59050_ _59033_/X _85437_/Q _59049_/X _59050_/Y sky130_fd_sc_hd__o21ai_4
X_83314_ _83325_/CLK _71956_/X _83314_/Q sky130_fd_sc_hd__dfxtp_4
X_80526_ _80526_/A _80526_/B _80536_/B sky130_fd_sc_hd__xor2_4
X_56262_ _56148_/X _56255_/X _56261_/Y _85255_/D sky130_fd_sc_hd__o21ai_4
X_68248_ _67538_/X _67541_/X _68216_/X _68248_/Y sky130_fd_sc_hd__a21oi_4
X_87082_ _87083_/CLK _87082_/D _87082_/Q sky130_fd_sc_hd__dfxtp_4
X_53474_ _48196_/A _53474_/B _51352_/C _53474_/X sky130_fd_sc_hd__and3_4
X_84294_ _84671_/CLK _63801_/Y _63800_/C sky130_fd_sc_hd__dfxtp_4
X_50686_ _50682_/A _49125_/X _50686_/Y sky130_fd_sc_hd__nand2_4
X_58001_ _57926_/X _85997_/Q _58000_/X _58001_/Y sky130_fd_sc_hd__o21ai_4
X_55213_ _55149_/A _84994_/Q _55213_/X sky130_fd_sc_hd__and2_4
X_86033_ _86040_/CLK _51319_/Y _65025_/B sky130_fd_sc_hd__dfxtp_4
X_52425_ _85825_/Q _52422_/X _52424_/Y _52425_/Y sky130_fd_sc_hd__o21ai_4
X_83245_ _84892_/CLK _72495_/X _83245_/Q sky130_fd_sc_hd__dfxtp_4
X_56193_ _56188_/X _55987_/X _56192_/Y _85281_/D sky130_fd_sc_hd__o21ai_4
X_80457_ _80457_/A _80456_/Y _80457_/X sky130_fd_sc_hd__xor2_4
X_68179_ _82059_/D _68160_/X _68178_/X _68179_/X sky130_fd_sc_hd__a21bo_4
X_70210_ _70214_/A _70214_/B _70210_/C _70204_/X _70210_/X sky130_fd_sc_hd__and4_4
X_55144_ _85131_/Q _55145_/B sky130_fd_sc_hd__inv_2
X_52356_ _52354_/Y _52340_/X _52355_/X _85839_/D sky130_fd_sc_hd__a21oi_4
X_40370_ _41061_/A _82335_/Q _40369_/X _40370_/X sky130_fd_sc_hd__o21a_4
X_71190_ _71190_/A _71190_/X sky130_fd_sc_hd__buf_2
X_83176_ _83508_/CLK _72793_/X _83176_/Q sky130_fd_sc_hd__dfxtp_4
X_80388_ _84754_/Q _66247_/C _80388_/Y sky130_fd_sc_hd__nand2_4
X_51307_ _51306_/X _46416_/A _51307_/X sky130_fd_sc_hd__and2_4
X_70141_ _83517_/Q _83165_/Q _83501_/Q _83149_/Q _70144_/B sky130_fd_sc_hd__a22oi_4
X_82127_ _83905_/CLK _77850_/X _82083_/D sky130_fd_sc_hd__dfxtp_4
X_55075_ _85323_/Q _55072_/X _55074_/Y _55075_/Y sky130_fd_sc_hd__o21ai_4
X_59952_ _59831_/X _60513_/A sky130_fd_sc_hd__buf_2
X_52287_ _52293_/A _52287_/B _52287_/Y sky130_fd_sc_hd__nand2_4
X_87984_ _87472_/CLK _87984_/D _87984_/Q sky130_fd_sc_hd__dfxtp_4
X_42040_ _42040_/A _42040_/Y sky130_fd_sc_hd__inv_2
X_58903_ _57965_/A _58904_/A sky130_fd_sc_hd__buf_2
X_54026_ _46449_/A _53964_/B _53969_/C _54026_/X sky130_fd_sc_hd__and3_4
X_51238_ _53944_/A _51238_/B _53944_/C _51238_/Y sky130_fd_sc_hd__nor3_4
X_70072_ _70040_/X _69890_/Y _70056_/X _70071_/Y _70072_/X sky130_fd_sc_hd__a211o_4
X_86935_ _86935_/CLK _86935_/D _67536_/B sky130_fd_sc_hd__dfxtp_4
X_82058_ _84020_/CLK _84018_/Q _82058_/Q sky130_fd_sc_hd__dfxtp_4
X_59883_ _59905_/B _59882_/X _59570_/A _60626_/A _59883_/Y sky130_fd_sc_hd__nor4_4
X_73900_ _86993_/Q _73776_/X _73899_/X _73913_/C sky130_fd_sc_hd__o21ai_4
X_81009_ _84223_/CLK _84217_/Q _81009_/Q sky130_fd_sc_hd__dfxtp_4
X_58834_ _58834_/A _59033_/A sky130_fd_sc_hd__buf_2
X_51169_ _51033_/A _51170_/A sky130_fd_sc_hd__buf_2
X_74880_ _74872_/Y _74897_/A _74897_/B _74887_/A sky130_fd_sc_hd__nand3_4
X_86866_ _86770_/CLK _86866_/D _63158_/B sky130_fd_sc_hd__dfxtp_4
X_85817_ _85529_/CLK _52465_/Y _85817_/Q sky130_fd_sc_hd__dfxtp_4
X_73831_ _73735_/X _85622_/Q _73782_/X _73830_/X _73831_/X sky130_fd_sc_hd__a211o_4
X_58765_ _44315_/A _58766_/A sky130_fd_sc_hd__buf_2
X_43991_ _87187_/Q _43954_/X _80669_/Q _43991_/Y sky130_fd_sc_hd__o21ai_4
X_55977_ _56196_/C _55690_/A _44052_/X _55976_/X _55977_/X sky130_fd_sc_hd__a211o_4
X_86797_ _87487_/CLK _86797_/D _66785_/B sky130_fd_sc_hd__dfxtp_4
X_45730_ _62057_/D _61582_/A sky130_fd_sc_hd__buf_2
X_57716_ _57716_/A _58882_/A sky130_fd_sc_hd__buf_2
X_76550_ _81661_/Q _76550_/Y sky130_fd_sc_hd__inv_2
X_42942_ _41778_/X _42930_/X _87639_/Q _42931_/X _87639_/D sky130_fd_sc_hd__a2bb2o_4
X_54928_ _54932_/A _54942_/B _54932_/C _53234_/D _54928_/X sky130_fd_sc_hd__and4_4
X_73762_ _73742_/A _66028_/B _73762_/X sky130_fd_sc_hd__and2_4
X_85748_ _85748_/CLK _52828_/Y _85748_/Q sky130_fd_sc_hd__dfxtp_4
X_70974_ _70976_/A _70952_/B _70969_/C _70974_/Y sky130_fd_sc_hd__nand3_4
X_58696_ _58696_/A _58696_/X sky130_fd_sc_hd__buf_2
X_75501_ _75500_/X _75503_/B sky130_fd_sc_hd__inv_2
X_72713_ _83181_/Q _72709_/X _72712_/X _72713_/X sky130_fd_sc_hd__a21o_4
X_45661_ _45659_/Y _45596_/X _45644_/X _45660_/Y _45661_/X sky130_fd_sc_hd__a211o_4
X_57647_ _84962_/Q _57635_/X _57646_/Y _57647_/Y sky130_fd_sc_hd__o21ai_4
X_76481_ _76481_/A _76485_/A sky130_fd_sc_hd__inv_2
X_42873_ _41592_/X _42866_/X _87674_/Q _42867_/X _42873_/X sky130_fd_sc_hd__a2bb2o_4
X_54859_ _54850_/A _54859_/B _54859_/Y sky130_fd_sc_hd__nand2_4
X_85679_ _85679_/CLK _85679_/D _85679_/Q sky130_fd_sc_hd__dfxtp_4
X_73693_ _73694_/B _73694_/C _73692_/X _73693_/X sky130_fd_sc_hd__a21o_4
X_47400_ _47418_/A _47408_/B _47377_/X _53023_/D _47400_/X sky130_fd_sc_hd__and4_4
X_78220_ _78220_/A _78220_/B _78220_/C _78221_/B sky130_fd_sc_hd__and3_4
X_44612_ _40968_/A _44602_/X _87033_/Q _44603_/X _44612_/X sky130_fd_sc_hd__a2bb2o_4
X_87418_ _82317_/CLK _43442_/X _87418_/Q sky130_fd_sc_hd__dfxtp_4
X_75432_ _75427_/X _75430_/Y _75432_/C _75432_/Y sky130_fd_sc_hd__nand3_4
X_41824_ _41802_/A _41824_/X sky130_fd_sc_hd__buf_2
X_48380_ _74373_/B _48380_/X sky130_fd_sc_hd__buf_2
X_72644_ _70183_/C _72631_/X _72643_/Y _83205_/D sky130_fd_sc_hd__a21bo_4
X_45592_ _63147_/B _61483_/A sky130_fd_sc_hd__buf_2
X_57578_ _57552_/X _48022_/Y _57578_/Y sky130_fd_sc_hd__nand2_4
X_88398_ _88398_/CLK _40397_/Y _88398_/Q sky130_fd_sc_hd__dfxtp_4
X_47331_ _47326_/Y _47317_/X _47330_/X _86646_/D sky130_fd_sc_hd__a21oi_4
X_59317_ _86663_/Q _59306_/B _59317_/Y sky130_fd_sc_hd__nor2_4
X_78151_ _78147_/Y _78150_/X _78151_/Y sky130_fd_sc_hd__nand2_4
X_44543_ _44543_/A _44543_/Y sky130_fd_sc_hd__inv_2
X_56529_ _56533_/A _56533_/B _85161_/Q _56529_/Y sky130_fd_sc_hd__nand3_4
X_75363_ _75359_/X _75362_/X _75370_/A sky130_fd_sc_hd__xor2_4
X_41755_ _40414_/X _41414_/A _41755_/X sky130_fd_sc_hd__or2_4
X_87349_ _86807_/CLK _43579_/X _87349_/Q sky130_fd_sc_hd__dfxtp_4
X_72575_ _72575_/A _72516_/A _72576_/A sky130_fd_sc_hd__nor2_4
X_77102_ _77112_/A _77113_/A _77103_/B sky130_fd_sc_hd__xor2_4
X_74314_ _72686_/A _74314_/X sky130_fd_sc_hd__buf_2
X_40706_ _40698_/X _82860_/Q _40705_/X _40707_/A sky130_fd_sc_hd__o21a_4
X_47262_ _57792_/A _47240_/X _47261_/Y _47262_/Y sky130_fd_sc_hd__o21ai_4
X_71526_ _53259_/B _71512_/A _71525_/Y _83466_/D sky130_fd_sc_hd__o21ai_4
X_59248_ _59121_/X _85421_/Q _59247_/X _59248_/Y sky130_fd_sc_hd__o21ai_4
X_78082_ _78082_/A _78082_/B _82939_/D sky130_fd_sc_hd__xor2_4
Xclkbuf_10_561_0_CLK clkbuf_9_280_0_CLK/X _81475_/CLK sky130_fd_sc_hd__clkbuf_1
X_44474_ _44602_/A _44474_/X sky130_fd_sc_hd__buf_2
X_75294_ _75294_/A _75293_/X _75294_/Y sky130_fd_sc_hd__xnor2_4
Xclkbuf_6_52_0_CLK clkbuf_6_53_0_CLK/A clkbuf_6_52_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_41686_ _41604_/A _41686_/B _41686_/X sky130_fd_sc_hd__or2_4
X_49001_ _48186_/A _49002_/A sky130_fd_sc_hd__buf_2
X_46213_ _59325_/A _46213_/X sky130_fd_sc_hd__buf_2
XPHY_250 sky130_fd_sc_hd__decap_3
X_77033_ _82087_/Q _77033_/B _82368_/D sky130_fd_sc_hd__xor2_4
X_43425_ _43166_/A _43425_/X sky130_fd_sc_hd__buf_2
X_74245_ _41976_/Y _56182_/X _73962_/X _74244_/Y _74245_/X sky130_fd_sc_hd__a211o_4
XPHY_261 sky130_fd_sc_hd__decap_3
X_40637_ _40637_/A _40836_/A sky130_fd_sc_hd__buf_2
X_47193_ _47147_/A _47196_/A sky130_fd_sc_hd__buf_2
X_59179_ _59177_/X _86067_/Q _59178_/X _59179_/Y sky130_fd_sc_hd__o21ai_4
X_71457_ _71445_/X _83492_/Q _71456_/Y _71457_/X sky130_fd_sc_hd__a21o_4
XPHY_272 sky130_fd_sc_hd__decap_3
XPHY_283 sky130_fd_sc_hd__decap_3
XPHY_294 sky130_fd_sc_hd__decap_3
X_61210_ _61107_/A _61083_/C _64234_/B _64457_/B sky130_fd_sc_hd__nand3_4
X_46144_ _46138_/A _46119_/A _46143_/Y _46134_/A _46144_/X sky130_fd_sc_hd__a211o_4
X_70408_ _51394_/B _70364_/A _70407_/Y _83778_/D sky130_fd_sc_hd__o21ai_4
X_43356_ _43287_/A _43356_/X sky130_fd_sc_hd__buf_2
X_74176_ _74173_/X _74175_/X _74085_/X _74176_/X sky130_fd_sc_hd__a21o_4
X_62190_ _62183_/X _62188_/Y _62189_/X _58374_/A _61782_/A _62190_/Y
+ sky130_fd_sc_hd__o32ai_4
X_40568_ _40568_/A _40568_/X sky130_fd_sc_hd__buf_2
X_71388_ _71458_/C _71399_/C sky130_fd_sc_hd__buf_2
X_42307_ _42204_/X _42307_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_576_0_CLK clkbuf_9_288_0_CLK/X _80849_/CLK sky130_fd_sc_hd__clkbuf_1
X_61141_ _61083_/B _61179_/A sky130_fd_sc_hd__inv_2
X_73127_ _69752_/B _57377_/X _73055_/X _73126_/Y _73127_/X sky130_fd_sc_hd__a211o_4
X_46075_ _46075_/A _46075_/Y sky130_fd_sc_hd__inv_2
X_70339_ _70337_/X _74795_/A _70338_/X _83792_/D sky130_fd_sc_hd__a21o_4
X_43287_ _43287_/A _43287_/X sky130_fd_sc_hd__buf_2
X_78984_ _82822_/Q _82534_/Q _78998_/B sky130_fd_sc_hd__xnor2_4
X_40499_ _82315_/Q _40471_/X _40499_/X sky130_fd_sc_hd__or2_4
X_49903_ _49794_/X _49904_/C sky130_fd_sc_hd__buf_2
X_45026_ _85273_/Q _44998_/X _45025_/X _45026_/Y sky130_fd_sc_hd__o21ai_4
X_42238_ _42231_/X _42226_/X _41403_/X _87965_/Q _42228_/X _42239_/A
+ sky130_fd_sc_hd__o32ai_4
X_61072_ _61071_/X _61122_/C sky130_fd_sc_hd__buf_2
X_77935_ _82073_/Q _77935_/Y sky130_fd_sc_hd__inv_2
X_73058_ _73054_/X _73057_/X _72951_/X _73058_/X sky130_fd_sc_hd__a21o_4
X_64900_ _64704_/X _86742_/Q _64707_/X _64899_/X _64900_/X sky130_fd_sc_hd__a211o_4
X_60023_ _59935_/A _62218_/A sky130_fd_sc_hd__buf_2
X_72009_ _72009_/A _72009_/X sky130_fd_sc_hd__buf_2
X_49834_ _49861_/A _49851_/B sky130_fd_sc_hd__buf_2
X_42169_ _42077_/A _42169_/X sky130_fd_sc_hd__buf_2
X_65880_ _65880_/A _65880_/X sky130_fd_sc_hd__buf_2
X_77866_ _77852_/Y _77866_/Y sky130_fd_sc_hd__inv_2
X_79605_ _79605_/A _79605_/B _79607_/A sky130_fd_sc_hd__xnor2_4
X_64831_ _64828_/X _85561_/Q _64829_/X _64830_/X _64831_/X sky130_fd_sc_hd__a211o_4
X_76817_ _76801_/B _76814_/X _76816_/Y _76818_/B sky130_fd_sc_hd__a21oi_4
X_49765_ _49657_/A _49789_/C sky130_fd_sc_hd__buf_2
X_46977_ _46959_/A _52781_/B _46977_/Y sky130_fd_sc_hd__nand2_4
X_77797_ _77763_/Y _77773_/A _77798_/B sky130_fd_sc_hd__nor2_4
X_48716_ _48714_/Y _48156_/X _48715_/X _48716_/Y sky130_fd_sc_hd__a21oi_4
X_67550_ _68342_/A _67550_/X sky130_fd_sc_hd__buf_2
X_79536_ _79534_/Y _79542_/A _79536_/Y sky130_fd_sc_hd__nand2_4
X_45928_ _43990_/Y _45927_/X _45928_/X sky130_fd_sc_hd__or2_4
X_64762_ _64751_/Y _64761_/Y _64762_/Y sky130_fd_sc_hd__nand2_4
X_76748_ _76746_/Y _76747_/Y _76757_/B sky130_fd_sc_hd__xor2_4
X_61974_ _61963_/X _61965_/X _61972_/Y _84738_/Q _61973_/X _61974_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49696_ _49641_/A _49697_/B sky130_fd_sc_hd__buf_2
X_66501_ _66501_/A _66501_/B _84111_/Q _66501_/X sky130_fd_sc_hd__and3_4
X_63713_ _63713_/A _60642_/A _60638_/Y _60642_/C _63713_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_10_514_0_CLK clkbuf_9_257_0_CLK/X _81333_/CLK sky130_fd_sc_hd__clkbuf_1
X_48647_ _83567_/Q _48647_/Y sky130_fd_sc_hd__inv_2
X_60925_ _60905_/Y _60913_/Y _60988_/A _60923_/Y _60924_/Y _84551_/D
+ sky130_fd_sc_hd__a41oi_4
X_67481_ _67126_/X _67575_/A sky130_fd_sc_hd__buf_2
X_79467_ _79467_/A _79467_/B _79468_/B sky130_fd_sc_hd__xor2_4
X_45859_ _45855_/X _45858_/X _44898_/X _45859_/X sky130_fd_sc_hd__a21o_4
X_64693_ _64601_/A _64694_/A sky130_fd_sc_hd__buf_2
X_76679_ _76672_/Y _76679_/Y sky130_fd_sc_hd__inv_2
X_69220_ _69179_/A _87277_/Q _69220_/X sky130_fd_sc_hd__and2_4
X_66432_ _66411_/X _66103_/Y _66431_/Y _66432_/Y sky130_fd_sc_hd__o21ai_4
X_78418_ _78418_/A _78418_/B _78423_/A sky130_fd_sc_hd__or2_4
X_63644_ _63644_/A _63670_/A sky130_fd_sc_hd__buf_2
X_48578_ _48578_/A _52199_/A sky130_fd_sc_hd__buf_2
X_60856_ _60855_/X _60865_/B sky130_fd_sc_hd__buf_2
X_79398_ _79374_/A _79373_/Y _79387_/A _79386_/Y _79398_/X sky130_fd_sc_hd__o22a_4
X_69151_ _87538_/Q _68958_/X _69113_/X _69150_/X _69151_/X sky130_fd_sc_hd__a211o_4
X_47529_ _86625_/Q _47524_/X _47528_/Y _47529_/Y sky130_fd_sc_hd__o21ai_4
X_66363_ _66003_/A _66415_/B sky130_fd_sc_hd__buf_2
X_78349_ _78345_/X _78346_/Y _78350_/A _78353_/C sky130_fd_sc_hd__a21o_4
X_63575_ _58438_/A _63541_/B _63575_/C _63541_/D _63575_/Y sky130_fd_sc_hd__nand4_4
X_60787_ _60778_/Y _60782_/Y _60708_/Y _60785_/Y _60786_/Y _60787_/Y
+ sky130_fd_sc_hd__a41oi_4
X_68102_ _66655_/X _66657_/X _68062_/X _68102_/Y sky130_fd_sc_hd__a21oi_4
X_65314_ _64691_/X _86150_/Q _64972_/X _65313_/X _65314_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_529_0_CLK clkbuf_9_264_0_CLK/X _81351_/CLK sky130_fd_sc_hd__clkbuf_1
X_50540_ _50536_/Y _50525_/X _50539_/X _86182_/D sky130_fd_sc_hd__a21oi_4
X_62526_ _62516_/X _62521_/Y _62525_/X _58457_/A _62511_/X _62526_/Y
+ sky130_fd_sc_hd__o32ai_4
X_81360_ _81361_/CLK _81360_/D _81360_/Q sky130_fd_sc_hd__dfxtp_4
X_69082_ _87074_/Q _69058_/X _68993_/X _69081_/X _69082_/X sky130_fd_sc_hd__a211o_4
X_66294_ _66366_/A _66294_/X sky130_fd_sc_hd__buf_2
X_68033_ _68429_/A _68033_/X sky130_fd_sc_hd__buf_2
X_80311_ _80308_/Y _80310_/Y _80315_/A sky130_fd_sc_hd__nand2_4
X_65245_ _65268_/A _65268_/B _84209_/Q _65245_/X sky130_fd_sc_hd__and3_4
X_50471_ _50481_/A _48788_/B _50471_/Y sky130_fd_sc_hd__nand2_4
X_62457_ _62415_/X _83248_/Q _62618_/D _62194_/D _62457_/X sky130_fd_sc_hd__and4_4
X_81291_ _81631_/CLK _76979_/X _81259_/D sky130_fd_sc_hd__dfxtp_4
X_52210_ _52210_/A _50508_/B _52210_/Y sky130_fd_sc_hd__nand2_4
X_83030_ _85269_/CLK _83030_/D _45081_/A sky130_fd_sc_hd__dfxtp_4
X_61408_ _61317_/X _61452_/C sky130_fd_sc_hd__buf_2
X_80242_ _80242_/A _80241_/X _80242_/Y sky130_fd_sc_hd__xnor2_4
X_53190_ _53190_/A _53211_/A sky130_fd_sc_hd__buf_2
X_65176_ _65035_/X _85515_/Q _65036_/X _65175_/X _65176_/X sky130_fd_sc_hd__a211o_4
X_62388_ _61481_/X _62420_/B _62420_/C _62334_/D _62389_/D sky130_fd_sc_hd__nand4_4
X_52141_ _48752_/A _52140_/X _52156_/C _52141_/X sky130_fd_sc_hd__and3_4
X_64127_ _64162_/A _58348_/A _64173_/C _64127_/X sky130_fd_sc_hd__and3_4
X_61339_ _72507_/A _61340_/A sky130_fd_sc_hd__buf_2
X_80173_ _80167_/A _80166_/X _80172_/Y _80173_/Y sky130_fd_sc_hd__a21boi_4
X_69984_ _70012_/A _69984_/X sky130_fd_sc_hd__buf_2
X_52072_ _52083_/A _50372_/B _52072_/Y sky130_fd_sc_hd__nand2_4
X_64058_ _63241_/B _64118_/B _64155_/C _64142_/D _64058_/Y sky130_fd_sc_hd__nand4_4
X_68935_ _68934_/X _42518_/Y _68935_/Y sky130_fd_sc_hd__nor2_4
X_84981_ _84981_/CLK _84981_/D _84981_/Q sky130_fd_sc_hd__dfxtp_4
X_55900_ _55949_/A _55900_/B _55900_/X sky130_fd_sc_hd__and2_4
X_51023_ _86088_/Q _51020_/X _51022_/Y _51023_/Y sky130_fd_sc_hd__o21ai_4
X_63009_ _60447_/B _63010_/A sky130_fd_sc_hd__buf_2
X_86720_ _86400_/CLK _86720_/D _58577_/A sky130_fd_sc_hd__dfxtp_4
X_83932_ _83932_/CLK _83932_/D _81396_/D sky130_fd_sc_hd__dfxtp_4
X_56880_ _56878_/Y _56880_/B _44134_/X _56880_/X sky130_fd_sc_hd__or3_4
X_68866_ _86987_/Q _68864_/X _68421_/X _68865_/X _68866_/X sky130_fd_sc_hd__a211o_4
X_55831_ _55836_/A _85233_/Q _55831_/X sky130_fd_sc_hd__and2_4
X_67817_ _68479_/A _67817_/X sky130_fd_sc_hd__buf_2
X_86651_ _86651_/CLK _86651_/D _86651_/Q sky130_fd_sc_hd__dfxtp_4
X_83863_ _82553_/CLK _70051_/X _82543_/D sky130_fd_sc_hd__dfxtp_4
X_68797_ _87086_/Q _68353_/X _68354_/X _68796_/X _68798_/B sky130_fd_sc_hd__a211o_4
X_85602_ _86210_/CLK _85602_/D _85602_/Q sky130_fd_sc_hd__dfxtp_4
X_58550_ _84821_/Q _58551_/A sky130_fd_sc_hd__inv_2
X_82814_ _81019_/CLK _82814_/D _78728_/A sky130_fd_sc_hd__dfxtp_4
X_67748_ _67270_/X _67748_/X sky130_fd_sc_hd__buf_2
X_55762_ _83015_/Q _44059_/X _55172_/X _55761_/X _55762_/X sky130_fd_sc_hd__a211o_4
X_86582_ _86582_/CLK _86582_/D _73830_/B sky130_fd_sc_hd__dfxtp_4
X_52974_ _85720_/Q _52957_/X _52973_/Y _52974_/Y sky130_fd_sc_hd__o21ai_4
X_83794_ _81620_/CLK _83794_/D _83794_/Q sky130_fd_sc_hd__dfxtp_4
X_57501_ _57497_/A _50234_/B _57501_/Y sky130_fd_sc_hd__nand2_4
X_88321_ _88062_/CLK _40863_/Y _88321_/Q sky130_fd_sc_hd__dfxtp_4
X_54713_ _54710_/Y _54694_/X _54712_/X _85392_/D sky130_fd_sc_hd__a21oi_4
X_85533_ _86246_/CLK _85533_/D _85533_/Q sky130_fd_sc_hd__dfxtp_4
X_51925_ _73561_/B _42612_/X _51924_/X _51926_/A sky130_fd_sc_hd__o21ai_4
X_58481_ _84838_/Q _58483_/A sky130_fd_sc_hd__buf_2
X_82745_ _84175_/CLK _84129_/Q _82745_/Q sky130_fd_sc_hd__dfxtp_4
X_55693_ _56192_/C _55690_/X _44052_/X _55692_/X _55693_/X sky130_fd_sc_hd__a211o_4
X_67679_ _67678_/X _67679_/B _67679_/X sky130_fd_sc_hd__and2_4
X_57432_ _57465_/A _57007_/X _57432_/Y sky130_fd_sc_hd__nor2_4
X_69418_ _69575_/A _69418_/X sky130_fd_sc_hd__buf_2
X_88252_ _87073_/CLK _88252_/D _88252_/Q sky130_fd_sc_hd__dfxtp_4
X_54644_ _54537_/A _54644_/X sky130_fd_sc_hd__buf_2
X_85464_ _82768_/CLK _85464_/D _85464_/Q sky130_fd_sc_hd__dfxtp_4
X_51856_ _51854_/Y _51850_/X _51855_/X _51856_/Y sky130_fd_sc_hd__a21oi_4
X_70690_ _70664_/A _47505_/A _70689_/Y _83723_/D sky130_fd_sc_hd__a21o_4
X_82676_ _81198_/CLK _82720_/Q _82676_/Q sky130_fd_sc_hd__dfxtp_4
X_87203_ _87394_/CLK _87203_/D _67729_/B sky130_fd_sc_hd__dfxtp_4
X_84415_ _84421_/CLK _84415_/D _84415_/Q sky130_fd_sc_hd__dfxtp_4
X_50807_ _86129_/Q _50804_/X _50806_/Y _50807_/Y sky130_fd_sc_hd__o21ai_4
X_81627_ _81627_/CLK _81627_/D _81819_/D sky130_fd_sc_hd__dfxtp_4
X_57363_ _56688_/X _73191_/B sky130_fd_sc_hd__buf_2
X_69349_ _87024_/Q _69153_/X _69168_/X _69348_/X _69349_/X sky130_fd_sc_hd__a211o_4
X_88183_ _87417_/CLK _41610_/Y _88183_/Q sky130_fd_sc_hd__dfxtp_4
X_54575_ _54521_/A _54585_/B sky130_fd_sc_hd__buf_2
X_85395_ _85491_/CLK _54696_/Y _85395_/Q sky130_fd_sc_hd__dfxtp_4
X_51787_ _51794_/A _51794_/B _51794_/C _51787_/D _51787_/X sky130_fd_sc_hd__and4_4
X_59102_ _84768_/Q _59102_/Y sky130_fd_sc_hd__inv_2
X_56314_ _56055_/X _56305_/X _56313_/Y _85240_/D sky130_fd_sc_hd__o21ai_4
X_87134_ _87888_/CLK _87134_/D _87134_/Q sky130_fd_sc_hd__dfxtp_4
X_41540_ _41336_/X _41540_/X sky130_fd_sc_hd__buf_2
X_53526_ _53523_/Y _53524_/X _53525_/Y _53526_/Y sky130_fd_sc_hd__a21boi_4
X_72360_ _72264_/X _85357_/Q _72359_/X _72360_/Y sky130_fd_sc_hd__o21ai_4
X_84346_ _82253_/CLK _84346_/D _84346_/Q sky130_fd_sc_hd__dfxtp_4
X_50738_ _50738_/A _50738_/B _50738_/Y sky130_fd_sc_hd__nand2_4
X_57294_ _57292_/Y _57293_/Y _57249_/X _57295_/B sky130_fd_sc_hd__a21o_4
X_81558_ _81330_/CLK _81558_/D _81514_/D sky130_fd_sc_hd__dfxtp_4
X_59033_ _59033_/A _59033_/X sky130_fd_sc_hd__buf_2
X_71311_ _71500_/A _71314_/B _71333_/C _71311_/Y sky130_fd_sc_hd__nand3_4
X_56245_ _56245_/A _56253_/B sky130_fd_sc_hd__buf_2
X_80509_ _80487_/A _80502_/A _80509_/Y sky130_fd_sc_hd__nand2_4
X_87065_ _87063_/CLK _87065_/D _44531_/A sky130_fd_sc_hd__dfxtp_4
X_53457_ _53821_/B _53458_/A sky130_fd_sc_hd__buf_2
X_41471_ _81182_/Q _41471_/B _41471_/X sky130_fd_sc_hd__or2_4
X_72291_ _72228_/X _85971_/Q _72290_/X _72291_/Y sky130_fd_sc_hd__o21ai_4
X_84277_ _84273_/CLK _64075_/Y _80040_/B sky130_fd_sc_hd__dfxtp_4
X_50669_ _50667_/Y _50609_/X _50668_/X _50669_/Y sky130_fd_sc_hd__a21oi_4
X_81489_ _81492_/CLK _84057_/Q _81489_/Q sky130_fd_sc_hd__dfxtp_4
X_43210_ _40955_/X _43180_/X _87536_/Q _43185_/X _43210_/X sky130_fd_sc_hd__a2bb2o_4
X_74030_ _70109_/Y _73939_/X _74029_/X _83126_/D sky130_fd_sc_hd__o21ai_4
X_86016_ _85727_/CLK _86016_/D _86016_/Q sky130_fd_sc_hd__dfxtp_4
X_40422_ _40321_/A _40947_/A sky130_fd_sc_hd__buf_2
X_52408_ _52406_/Y _52390_/X _52407_/X _52408_/Y sky130_fd_sc_hd__a21oi_4
X_71242_ _71225_/A _71248_/C sky130_fd_sc_hd__buf_2
X_83228_ _83231_/CLK _72582_/Y _79372_/B sky130_fd_sc_hd__dfxtp_4
X_44190_ _44189_/X _72899_/A sky130_fd_sc_hd__buf_2
X_56176_ _44907_/A _56177_/B sky130_fd_sc_hd__buf_2
X_53388_ _53371_/A _53388_/B _53388_/C _52872_/D _53388_/X sky130_fd_sc_hd__and4_4
X_43141_ _43141_/A _43141_/Y sky130_fd_sc_hd__inv_2
X_55127_ _80665_/Q _55128_/A sky130_fd_sc_hd__buf_2
X_40353_ _46725_/A _74458_/A _46290_/A _40353_/Y sky130_fd_sc_hd__a21oi_4
X_52339_ _85842_/Q _52324_/X _52338_/Y _52339_/Y sky130_fd_sc_hd__o21ai_4
X_71173_ _71173_/A _71173_/B _71181_/C _71178_/D _71173_/Y sky130_fd_sc_hd__nand4_4
X_83159_ _85895_/CLK _83159_/D _83159_/Q sky130_fd_sc_hd__dfxtp_4
X_70124_ _83140_/Q _70125_/D sky130_fd_sc_hd__inv_2
X_55058_ _55055_/Y _55050_/X _55057_/X _85327_/D sky130_fd_sc_hd__a21oi_4
X_59935_ _59935_/A _62237_/A _59973_/A _59943_/A _59935_/X sky130_fd_sc_hd__and4_4
X_43072_ _43146_/A _43072_/X sky130_fd_sc_hd__buf_2
X_75981_ _75981_/A _75980_/Y _75982_/B sky130_fd_sc_hd__xor2_4
X_87967_ _87720_/CLK _42236_/X _87967_/Q sky130_fd_sc_hd__dfxtp_4
X_46900_ _46860_/X _46899_/X _46900_/Y sky130_fd_sc_hd__nand2_4
X_42023_ _42023_/A _42023_/Y sky130_fd_sc_hd__inv_2
X_54009_ _53991_/A _46411_/A _54009_/Y sky130_fd_sc_hd__nand2_4
X_77720_ _77723_/A _77723_/C _82209_/D sky130_fd_sc_hd__nand2_4
X_86918_ _87141_/CLK _86918_/D _67929_/B sky130_fd_sc_hd__dfxtp_4
X_74932_ _74931_/Y _74923_/B _74932_/X sky130_fd_sc_hd__and2_4
X_70055_ _83862_/Q _70048_/X _70054_/Y _83862_/D sky130_fd_sc_hd__a21bo_4
X_47880_ _47880_/A _47880_/Y sky130_fd_sc_hd__inv_2
X_59866_ _80294_/B _59866_/Y sky130_fd_sc_hd__inv_2
X_87898_ _87898_/CLK _42367_/Y _87898_/Q sky130_fd_sc_hd__dfxtp_4
X_46831_ _46827_/Y _46798_/X _46830_/X _86699_/D sky130_fd_sc_hd__a21oi_4
X_58817_ _84798_/Q _58725_/X _58808_/X _58816_/X _84798_/D sky130_fd_sc_hd__a2bb2oi_4
X_77651_ _82238_/Q _77655_/A sky130_fd_sc_hd__inv_2
X_74863_ _80932_/Q _74863_/B _81213_/D sky130_fd_sc_hd__xnor2_4
X_86849_ _84420_/CLK _45866_/Y _63342_/B sky130_fd_sc_hd__dfxtp_4
X_59797_ _59797_/A _59797_/B _59797_/Y sky130_fd_sc_hd__nor2_4
X_76602_ _76597_/X _76602_/B _76598_/Y _76602_/Y sky130_fd_sc_hd__nand3_4
X_49550_ _49547_/Y _49541_/X _49549_/X _86367_/D sky130_fd_sc_hd__a21oi_4
X_73814_ _73815_/B _73815_/C _73813_/X _73814_/X sky130_fd_sc_hd__a21o_4
X_46762_ _46762_/A _54353_/D sky130_fd_sc_hd__inv_2
X_58748_ _58864_/A _58748_/X sky130_fd_sc_hd__buf_2
X_77582_ _77582_/A _82118_/Q _77583_/A sky130_fd_sc_hd__nand2_4
X_43974_ _87169_/Q _43975_/B sky130_fd_sc_hd__inv_2
X_74794_ _74723_/X _74794_/B _74780_/D _74794_/Y sky130_fd_sc_hd__nand3_4
X_48501_ _52161_/A _48500_/X _48533_/C _48501_/X sky130_fd_sc_hd__and3_4
X_79321_ _79321_/A _79321_/B _79322_/B sky130_fd_sc_hd__xor2_4
X_45713_ _45713_/A _45746_/B _45713_/Y sky130_fd_sc_hd__nand2_4
X_76533_ _81276_/Q _76533_/B _76533_/Y sky130_fd_sc_hd__nand2_4
X_42925_ _41727_/X _42920_/X _87649_/Q _42922_/X _87649_/D sky130_fd_sc_hd__a2bb2o_4
X_49481_ _49481_/A _51003_/B _49481_/Y sky130_fd_sc_hd__nand2_4
X_73745_ _57523_/B _73745_/B _73745_/X sky130_fd_sc_hd__xor2_4
X_46693_ _54309_/B _51791_/B sky130_fd_sc_hd__buf_2
X_58679_ _58679_/A _58679_/X sky130_fd_sc_hd__buf_2
X_70957_ _70969_/A _71066_/B _70954_/C _70957_/Y sky130_fd_sc_hd__nand3_4
X_48432_ _48425_/Y _48383_/X _48431_/X _48432_/Y sky130_fd_sc_hd__a21oi_4
X_60710_ _60713_/A _60659_/A _60722_/A sky130_fd_sc_hd__nor2_4
X_79252_ _79224_/B _79240_/Y _79238_/Y _79252_/Y sky130_fd_sc_hd__a21boi_4
X_45644_ _45720_/A _45644_/X sky130_fd_sc_hd__buf_2
X_76464_ _76482_/B _76463_/X _76464_/Y sky130_fd_sc_hd__nand2_4
X_42856_ _42847_/X _42849_/X _41536_/X _66927_/B _42836_/X _42856_/Y
+ sky130_fd_sc_hd__o32ai_4
X_61690_ _61690_/A _61690_/B _61690_/C _61690_/Y sky130_fd_sc_hd__nor3_4
X_73676_ _68491_/B _73674_/X _73344_/X _73675_/Y _73676_/X sky130_fd_sc_hd__a211o_4
X_70888_ _70860_/A _70890_/B _70890_/C _70890_/D _70888_/Y sky130_fd_sc_hd__nand4_4
X_78203_ _78203_/A _82492_/Q _78220_/A sky130_fd_sc_hd__xor2_4
X_75415_ _75396_/A _75393_/Y _75394_/Y _75416_/A sky130_fd_sc_hd__o21a_4
X_41807_ _40391_/X _41799_/X _66683_/B _41800_/X _88143_/D sky130_fd_sc_hd__a2bb2o_4
X_48363_ _74366_/A _53620_/A sky130_fd_sc_hd__buf_2
X_60641_ _60641_/A _60642_/C sky130_fd_sc_hd__inv_2
X_72627_ _60069_/Y _72583_/Y _72625_/X _61079_/Y _72626_/Y _72627_/Y
+ sky130_fd_sc_hd__a41oi_4
X_79183_ _79183_/A _79183_/B _79185_/B sky130_fd_sc_hd__nand2_4
X_45575_ _45575_/A _45604_/B _45575_/Y sky130_fd_sc_hd__nor2_4
X_76395_ _81651_/Q _76395_/Y sky130_fd_sc_hd__inv_2
X_42787_ _42745_/A _42787_/X sky130_fd_sc_hd__buf_2
X_47314_ _47313_/Y _52979_/B sky130_fd_sc_hd__buf_2
X_78134_ _78125_/Y _78134_/B _78134_/Y sky130_fd_sc_hd__nor2_4
X_44526_ _87066_/Q _44526_/Y sky130_fd_sc_hd__inv_2
X_63360_ _60798_/X _63355_/Y _63358_/X _63359_/Y _63360_/X sky130_fd_sc_hd__a211o_4
X_75346_ _75346_/A _75345_/X _80756_/D sky130_fd_sc_hd__xor2_4
X_41738_ _41737_/Y _88159_/D sky130_fd_sc_hd__inv_2
X_48294_ _49223_/A _48319_/A sky130_fd_sc_hd__buf_2
X_60572_ _60572_/A _60572_/B _60572_/C _60572_/X sky130_fd_sc_hd__and3_4
X_72558_ _64561_/A _57872_/A _79436_/B _72558_/X sky130_fd_sc_hd__or3_4
X_62311_ _62304_/X _62306_/X _62310_/Y _84915_/Q _62300_/X _62311_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47245_ _57734_/A _47240_/X _47244_/Y _47245_/Y sky130_fd_sc_hd__o21ai_4
X_71509_ _71525_/A _71512_/A sky130_fd_sc_hd__buf_2
X_78065_ _84570_/Q _78065_/B _78065_/X sky130_fd_sc_hd__xor2_4
X_44457_ _44457_/A _44457_/Y sky130_fd_sc_hd__inv_2
X_75277_ _75277_/A _75276_/Y _75303_/B sky130_fd_sc_hd__and2_4
X_63291_ _63289_/X _84888_/Q _63341_/C _63332_/D _63291_/X sky130_fd_sc_hd__and4_4
X_41669_ _41611_/X _41613_/X _41667_/X _88172_/Q _41668_/X _41670_/A
+ sky130_fd_sc_hd__o32ai_4
X_72489_ _72484_/X _83384_/Q _72488_/Y _83248_/D sky130_fd_sc_hd__o21a_4
X_65030_ _64797_/X _86737_/Q _65028_/X _65029_/X _65031_/B sky130_fd_sc_hd__a211o_4
X_77016_ _77017_/B _77016_/Y sky130_fd_sc_hd__inv_2
X_43408_ _43399_/X _43404_/X _41498_/X _87436_/Q _43407_/X _43408_/Y
+ sky130_fd_sc_hd__o32ai_4
X_62242_ _62240_/Y _62166_/X _62241_/Y _84424_/D sky130_fd_sc_hd__a21oi_4
X_74228_ _74225_/X _74227_/X _73602_/X _74228_/X sky130_fd_sc_hd__a21o_4
X_47176_ _86662_/Q _47145_/X _47175_/Y _47176_/Y sky130_fd_sc_hd__o21ai_4
X_44388_ _41461_/X _44377_/X _87135_/Q _44379_/X _44388_/X sky130_fd_sc_hd__a2bb2o_4
X_46127_ _46094_/X _46128_/D sky130_fd_sc_hd__inv_2
X_43339_ _41302_/X _43336_/X _87472_/Q _43337_/X _87472_/D sky130_fd_sc_hd__a2bb2o_4
X_62173_ _61682_/B _62161_/B _62187_/C _61706_/X _62173_/Y sky130_fd_sc_hd__nand4_4
X_74159_ _74154_/X _74158_/X _74160_/B sky130_fd_sc_hd__nand2_4
X_61124_ _64306_/A _64525_/B sky130_fd_sc_hd__buf_2
X_46058_ _46058_/A _86790_/D sky130_fd_sc_hd__inv_2
X_66981_ _66625_/A _67057_/A sky130_fd_sc_hd__buf_2
X_78967_ _82820_/Q _82532_/Q _78967_/Y sky130_fd_sc_hd__xnor2_4
X_45009_ _64284_/B _61398_/B sky130_fd_sc_hd__buf_2
X_68720_ _68717_/X _68719_/X _58002_/A _68720_/X sky130_fd_sc_hd__a21o_4
X_65932_ _65932_/A _65932_/B _65932_/X sky130_fd_sc_hd__and2_4
X_61055_ _61055_/A _61000_/X _61055_/C _61055_/X sky130_fd_sc_hd__or3_4
X_77918_ _82071_/Q _77920_/A sky130_fd_sc_hd__inv_2
X_78898_ _82635_/Q _82507_/D _78897_/X _78898_/Y sky130_fd_sc_hd__o21ai_4
X_60006_ _80186_/A _59787_/X _60003_/Y _60005_/Y _60007_/A sky130_fd_sc_hd__a2bb2o_4
X_49817_ _49925_/A _49830_/A sky130_fd_sc_hd__buf_2
X_68651_ _68651_/A _68651_/X sky130_fd_sc_hd__buf_2
X_65863_ _65858_/X _65862_/X _65809_/X _65863_/X sky130_fd_sc_hd__a21o_4
X_77849_ _77849_/A _77849_/B _77850_/B sky130_fd_sc_hd__xnor2_4
X_67602_ _67602_/A _67602_/B _67602_/Y sky130_fd_sc_hd__nand2_4
X_64814_ _64939_/A _64814_/X sky130_fd_sc_hd__buf_2
X_49748_ _49757_/A _52965_/B _49748_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_453_0_CLK clkbuf_9_226_0_CLK/X _85697_/CLK sky130_fd_sc_hd__clkbuf_1
X_68582_ _87095_/Q _68580_/X _68509_/X _68581_/X _68582_/X sky130_fd_sc_hd__a211o_4
X_80860_ _80740_/CLK _80892_/Q _75042_/B sky130_fd_sc_hd__dfxtp_4
X_65794_ _65779_/A _86473_/Q _65794_/X sky130_fd_sc_hd__and2_4
X_67533_ _67055_/X _67533_/X sky130_fd_sc_hd__buf_2
X_79519_ _79519_/A _79520_/B sky130_fd_sc_hd__inv_2
X_64745_ _64680_/A _64745_/B _64745_/X sky130_fd_sc_hd__and2_4
X_49679_ _49678_/X _49685_/A sky130_fd_sc_hd__buf_2
X_61957_ _61957_/A _61952_/Y _61953_/Y _61956_/Y _61957_/Y sky130_fd_sc_hd__nand4_4
X_80791_ _83973_/CLK _80791_/D _80791_/Q sky130_fd_sc_hd__dfxtp_4
X_51710_ _51709_/X _51715_/B _51695_/C _53234_/D _51710_/X sky130_fd_sc_hd__and4_4
X_82530_ _82786_/CLK _82530_/D _78949_/B sky130_fd_sc_hd__dfxtp_4
X_60908_ _60908_/A _60908_/X sky130_fd_sc_hd__buf_2
X_67464_ _87406_/Q _67394_/X _67462_/X _67463_/X _67464_/X sky130_fd_sc_hd__a211o_4
X_52690_ _52674_/X _52694_/B _52694_/C _46810_/X _52690_/X sky130_fd_sc_hd__and4_4
X_64676_ _64676_/A _85854_/Q _64676_/X sky130_fd_sc_hd__and2_4
X_61888_ _59668_/B _61907_/C sky130_fd_sc_hd__buf_2
X_69203_ _69067_/A _69203_/B _69203_/X sky130_fd_sc_hd__and2_4
X_66415_ _66433_/A _66415_/B _66415_/C _66415_/X sky130_fd_sc_hd__and3_4
Xclkbuf_10_468_0_CLK clkbuf_9_234_0_CLK/X _85444_/CLK sky130_fd_sc_hd__clkbuf_1
X_51641_ _51629_/X _51651_/B _51651_/C _53165_/D _51641_/X sky130_fd_sc_hd__and4_4
X_63627_ _63372_/A _63627_/X sky130_fd_sc_hd__buf_2
X_82461_ _83514_/CLK _79153_/X _82429_/D sky130_fd_sc_hd__dfxtp_4
X_60839_ _60826_/A _60838_/X _78049_/A _60839_/Y sky130_fd_sc_hd__nor3_4
X_67395_ _67320_/A _67395_/B _67395_/X sky130_fd_sc_hd__and2_4
X_84200_ _85315_/CLK _84200_/D _65449_/C sky130_fd_sc_hd__dfxtp_4
X_81412_ _81412_/CLK _81412_/D _75930_/B sky130_fd_sc_hd__dfxtp_4
X_69134_ _69134_/A _87795_/Q _69134_/X sky130_fd_sc_hd__and2_4
X_54360_ _54355_/A _52667_/B _54360_/Y sky130_fd_sc_hd__nand2_4
X_66346_ _66342_/Y _66343_/X _66345_/Y _84139_/D sky130_fd_sc_hd__a21o_4
X_85180_ _85180_/CLK _85180_/D _85180_/Q sky130_fd_sc_hd__dfxtp_4
X_51572_ _51590_/A _53101_/B _51572_/Y sky130_fd_sc_hd__nand2_4
X_63558_ _63436_/A _63558_/X sky130_fd_sc_hd__buf_2
X_82392_ _83681_/CLK _82392_/D _82392_/Q sky130_fd_sc_hd__dfxtp_4
X_53311_ _53311_/A _53330_/A sky130_fd_sc_hd__buf_2
X_84131_ _82975_/CLK _84131_/D _84131_/Q sky130_fd_sc_hd__dfxtp_4
X_50523_ _50523_/A _51010_/A sky130_fd_sc_hd__buf_2
X_62509_ _62570_/A _63610_/B _62601_/C _62463_/X _62509_/X sky130_fd_sc_hd__and4_4
X_81343_ _83926_/CLK _81343_/D _81719_/D sky130_fd_sc_hd__dfxtp_4
X_69065_ _70009_/A _69065_/X sky130_fd_sc_hd__buf_2
X_54291_ _54317_/A _54312_/C sky130_fd_sc_hd__buf_2
X_66277_ _66179_/X _66275_/Y _66276_/Y _66277_/Y sky130_fd_sc_hd__o21ai_4
X_63489_ _63463_/A _84959_/Q _63476_/C _63489_/X sky130_fd_sc_hd__and3_4
X_56030_ _74297_/C _56030_/B _56030_/X sky130_fd_sc_hd__xor2_4
X_68016_ _67948_/X _68005_/Y _67983_/X _68015_/Y _68016_/X sky130_fd_sc_hd__a211o_4
X_53242_ _53189_/A _53242_/X sky130_fd_sc_hd__buf_2
X_65228_ _65118_/X _85545_/Q _65146_/X _65227_/X _65228_/X sky130_fd_sc_hd__a211o_4
X_84062_ _82648_/CLK _84062_/D _81494_/D sky130_fd_sc_hd__dfxtp_4
X_50454_ _86197_/Q _50437_/X _50453_/Y _50454_/Y sky130_fd_sc_hd__o21ai_4
X_81274_ _81279_/CLK _81306_/Q _76503_/A sky130_fd_sc_hd__dfxtp_4
X_83013_ _83013_/CLK _83013_/D _45331_/A sky130_fd_sc_hd__dfxtp_4
X_80225_ _80222_/X _80225_/B _80224_/X _80226_/A sky130_fd_sc_hd__and3_4
X_53173_ _53199_/A _53187_/A sky130_fd_sc_hd__buf_2
X_65159_ _65159_/A _86252_/Q _65159_/X sky130_fd_sc_hd__and2_4
X_50385_ _50381_/A _50385_/B _50385_/Y sky130_fd_sc_hd__nand2_4
X_52124_ _52122_/Y _52117_/X _52123_/Y _85884_/D sky130_fd_sc_hd__a21boi_4
X_87821_ _87821_/CLK _42559_/Y _87821_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_406_0_CLK clkbuf_9_203_0_CLK/X _83278_/CLK sky130_fd_sc_hd__clkbuf_1
X_80156_ _80178_/A _80156_/Y sky130_fd_sc_hd__inv_2
X_57981_ _58857_/A _57981_/X sky130_fd_sc_hd__buf_2
X_69967_ _69633_/A _69967_/B _69967_/X sky130_fd_sc_hd__and2_4
X_59720_ _59642_/X _59721_/A sky130_fd_sc_hd__buf_2
X_56932_ _72838_/A _72909_/A sky130_fd_sc_hd__buf_2
X_52055_ _52053_/Y _52022_/X _52054_/Y _85898_/D sky130_fd_sc_hd__a21boi_4
X_68918_ _68987_/A _68918_/B _68918_/X sky130_fd_sc_hd__and2_4
X_87752_ _88006_/CLK _87752_/D _87752_/Q sky130_fd_sc_hd__dfxtp_4
X_84964_ _86203_/CLK _84964_/D _84964_/Q sky130_fd_sc_hd__dfxtp_4
X_80087_ _80084_/X _80087_/B _81681_/D sky130_fd_sc_hd__xor2_4
X_69898_ _88058_/Q _69837_/X _69088_/X _69897_/Y _69898_/X sky130_fd_sc_hd__a211o_4
X_51006_ _51018_/A _50985_/B _51029_/C _52698_/D _51006_/X sky130_fd_sc_hd__and4_4
X_86703_ _86384_/CLK _86703_/D _86703_/Q sky130_fd_sc_hd__dfxtp_4
X_59651_ _59651_/A _59651_/B _59651_/C _59713_/A sky130_fd_sc_hd__nand3_4
X_83915_ _80784_/CLK _69552_/X _83915_/Q sky130_fd_sc_hd__dfxtp_4
X_56863_ _56995_/A _56863_/X sky130_fd_sc_hd__buf_2
X_68849_ _88000_/Q _68778_/X _68800_/X _68848_/X _68849_/X sky130_fd_sc_hd__a211o_4
X_87683_ _87686_/CLK _42860_/Y _66959_/B sky130_fd_sc_hd__dfxtp_4
X_84895_ _84895_/CLK _84895_/D _58258_/A sky130_fd_sc_hd__dfxtp_4
X_58602_ _58602_/A _58603_/A sky130_fd_sc_hd__buf_2
X_55814_ _44077_/X _55814_/B _55814_/X sky130_fd_sc_hd__and2_4
X_86634_ _85993_/CLK _86634_/D _86634_/Q sky130_fd_sc_hd__dfxtp_4
X_71860_ _71848_/X _83350_/Q _71859_/Y _83350_/D sky130_fd_sc_hd__a21o_4
X_59582_ _59582_/A _59582_/B _61071_/C sky130_fd_sc_hd__and2_4
X_83846_ _83846_/CLK _70182_/Y _83846_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_80_0_CLK clkbuf_8_81_0_CLK/A clkbuf_8_80_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_56794_ _56653_/Y _56651_/Y _56721_/D _56794_/Y sky130_fd_sc_hd__nor3_4
X_70811_ _52885_/B _70802_/X _70810_/Y _70811_/Y sky130_fd_sc_hd__o21ai_4
X_58533_ _58533_/A _58532_/X _58533_/Y sky130_fd_sc_hd__nor2_4
X_55745_ _56167_/B _56163_/A _56158_/A _55745_/D _56127_/C sky130_fd_sc_hd__nand4_4
X_86565_ _86213_/CLK _86565_/D _66310_/B sky130_fd_sc_hd__dfxtp_4
X_52957_ _53065_/A _52957_/X sky130_fd_sc_hd__buf_2
X_40971_ _40512_/X _41149_/A _40970_/X _40972_/A sky130_fd_sc_hd__o21a_4
X_71791_ _58192_/Y _71784_/X _71790_/Y _71791_/Y sky130_fd_sc_hd__o21ai_4
X_83777_ _86553_/CLK _70432_/Y _83777_/Q sky130_fd_sc_hd__dfxtp_4
X_80989_ _80968_/CLK _80989_/D _80945_/D sky130_fd_sc_hd__dfxtp_4
X_88304_ _86989_/CLK _88304_/D _88304_/Q sky130_fd_sc_hd__dfxtp_4
X_42710_ _42651_/X _42710_/X sky130_fd_sc_hd__buf_2
X_73530_ _69967_/B _73530_/B _73530_/Y sky130_fd_sc_hd__nor2_4
X_85516_ _85516_/CLK _85516_/D _85516_/Q sky130_fd_sc_hd__dfxtp_4
X_51908_ _85924_/Q _51900_/X _51907_/Y _51908_/Y sky130_fd_sc_hd__o21ai_4
X_70742_ _70740_/A _70710_/A _70742_/Y sky130_fd_sc_hd__nand2_4
X_82728_ _84111_/CLK _66495_/C _78862_/A sky130_fd_sc_hd__dfxtp_4
X_58464_ _84842_/Q _58465_/A sky130_fd_sc_hd__buf_2
X_43690_ _40806_/X _43685_/X _87307_/Q _43686_/X _87307_/D sky130_fd_sc_hd__a2bb2o_4
X_55676_ _55676_/A _55676_/B _55676_/C _55675_/X _55683_/B sky130_fd_sc_hd__and4_4
X_86496_ _86490_/CLK _86496_/D _65441_/B sky130_fd_sc_hd__dfxtp_4
X_52888_ _52886_/Y _52865_/X _52887_/X _52888_/Y sky130_fd_sc_hd__a21oi_4
X_57415_ _57275_/X _57270_/X _57414_/X _57415_/X sky130_fd_sc_hd__o21a_4
X_88235_ _86934_/CLK _88235_/D _88235_/Q sky130_fd_sc_hd__dfxtp_4
X_42641_ _42614_/X _42615_/X _40959_/X _87791_/Q _42637_/X _42641_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54627_ _54636_/A _54102_/B _54627_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_95_0_CLK clkbuf_8_95_0_CLK/A clkbuf_8_95_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_73461_ _83150_/Q _73437_/X _73460_/Y _83150_/D sky130_fd_sc_hd__a21o_4
X_85447_ _85447_/CLK _85447_/D _85447_/Q sky130_fd_sc_hd__dfxtp_4
X_51839_ _51836_/Y _51823_/X _51838_/X _51839_/Y sky130_fd_sc_hd__a21oi_4
X_70673_ _70673_/A _70676_/B _70676_/C _70673_/Y sky130_fd_sc_hd__nor3_4
X_58395_ _58388_/X _83348_/Q _58394_/Y _58395_/X sky130_fd_sc_hd__o21a_4
X_82659_ _82665_/CLK _82659_/D _82659_/Q sky130_fd_sc_hd__dfxtp_4
X_75200_ _75201_/B _75201_/A _75207_/B sky130_fd_sc_hd__or2_4
X_72412_ _83257_/Q _72381_/X _72406_/X _72411_/X _83257_/D sky130_fd_sc_hd__a2bb2oi_4
X_45360_ _44887_/X _45678_/A sky130_fd_sc_hd__buf_2
X_57346_ _57318_/D _56894_/Y _57346_/C _57346_/Y sky130_fd_sc_hd__nand3_4
X_76180_ _76178_/Y _76177_/Y _76174_/Y _76181_/A sky130_fd_sc_hd__nand3_4
X_88166_ _86930_/CLK _88166_/D _67659_/B sky130_fd_sc_hd__dfxtp_4
X_54558_ _54558_/A _54558_/X sky130_fd_sc_hd__buf_2
X_42572_ _42568_/X _42569_/X _40820_/X _69710_/B _42571_/X _42572_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73392_ _83153_/Q _73318_/X _73391_/Y _83153_/D sky130_fd_sc_hd__a21o_4
X_85378_ _85378_/CLK _54789_/Y _85378_/Q sky130_fd_sc_hd__dfxtp_4
X_44311_ _44301_/Y _44304_/Y _44318_/A _44311_/Y sky130_fd_sc_hd__a21oi_4
X_75131_ _75129_/Y _75126_/X _75143_/A _75131_/Y sky130_fd_sc_hd__nand3_4
X_87117_ _82888_/CLK _44420_/X _87117_/Q sky130_fd_sc_hd__dfxtp_4
X_41523_ _41523_/A _41523_/B _41523_/X sky130_fd_sc_hd__or2_4
X_72343_ _72209_/X _85967_/Q _72342_/X _72343_/Y sky130_fd_sc_hd__o21ai_4
X_53509_ _53509_/A _57537_/B _53509_/Y sky130_fd_sc_hd__nand2_4
X_84329_ _84329_/CLK _63366_/Y _63365_/C sky130_fd_sc_hd__dfxtp_4
X_45291_ _45290_/Y _45272_/X _45291_/Y sky130_fd_sc_hd__nand2_4
X_57277_ _45647_/Y _56671_/X _57277_/Y sky130_fd_sc_hd__nand2_4
X_88097_ _88097_/CLK _41946_/Y _73987_/A sky130_fd_sc_hd__dfxtp_4
X_54489_ _54483_/A _54471_/B _54483_/C _46999_/A _54489_/X sky130_fd_sc_hd__and4_4
X_47030_ _47026_/Y _46987_/X _47029_/X _86678_/D sky130_fd_sc_hd__a21oi_4
X_59016_ _59012_/Y _59015_/Y _58966_/X _59016_/X sky130_fd_sc_hd__a21o_4
X_44242_ _44227_/Y _87178_/Q _44242_/C _44242_/Y sky130_fd_sc_hd__nand3_4
X_56228_ _56074_/X _56225_/X _56227_/Y _85268_/D sky130_fd_sc_hd__o21ai_4
X_75062_ _75062_/A _75062_/B _75062_/Y sky130_fd_sc_hd__nor2_4
X_41454_ _41453_/Y _41454_/X sky130_fd_sc_hd__buf_2
X_87048_ _87045_/CLK _87048_/D _87048_/Q sky130_fd_sc_hd__dfxtp_4
X_72274_ _72176_/A _72274_/X sky130_fd_sc_hd__buf_2
X_74013_ _73709_/X _74038_/A sky130_fd_sc_hd__buf_2
X_40405_ _40404_/X _40342_/X _88396_/Q _40355_/X _40405_/X sky130_fd_sc_hd__a2bb2o_4
X_71225_ _71225_/A _71232_/C sky130_fd_sc_hd__buf_2
X_44173_ _44315_/A _44173_/X sky130_fd_sc_hd__buf_2
X_79870_ _79862_/X _79864_/B _79869_/Y _79870_/Y sky130_fd_sc_hd__a21boi_4
X_56159_ _56159_/A _56159_/X sky130_fd_sc_hd__buf_2
X_41385_ _81742_/Q _41379_/X _41385_/X sky130_fd_sc_hd__or2_4
X_43124_ _42059_/A _44530_/A sky130_fd_sc_hd__buf_2
X_78821_ _82723_/Q _78821_/B _78821_/X sky130_fd_sc_hd__xor2_4
X_40336_ _43175_/A _40591_/B sky130_fd_sc_hd__buf_2
X_71156_ _52121_/B _71138_/A _71155_/Y _71156_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_8_33_0_CLK clkbuf_7_16_0_CLK/X clkbuf_9_67_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_48981_ _83615_/Q _72007_/B sky130_fd_sc_hd__inv_2
X_70107_ _70107_/A _70107_/B _70107_/C _70106_/Y _70107_/Y sky130_fd_sc_hd__nand4_4
X_47932_ _47912_/A _47932_/B _47932_/Y sky130_fd_sc_hd__nand2_4
X_43055_ _87593_/Q _43055_/Y sky130_fd_sc_hd__inv_2
X_59918_ _59917_/X _59918_/Y sky130_fd_sc_hd__inv_2
X_78752_ _78752_/A _78753_/C sky130_fd_sc_hd__inv_2
X_71087_ _49015_/X _71070_/A _71086_/Y _71087_/Y sky130_fd_sc_hd__o21ai_4
X_75964_ _75964_/A _75963_/Y _75964_/X sky130_fd_sc_hd__and2_4
X_42006_ _42024_/A _42006_/X sky130_fd_sc_hd__buf_2
X_77703_ _77703_/A _77703_/B _77703_/C _77703_/Y sky130_fd_sc_hd__nand3_4
X_74915_ _81131_/D _74916_/B _74915_/Y sky130_fd_sc_hd__nor2_4
X_70038_ _69520_/X _69772_/Y _70033_/X _70037_/Y _70038_/X sky130_fd_sc_hd__a211o_4
X_47863_ _83558_/Q _47863_/Y sky130_fd_sc_hd__inv_2
X_59849_ _59634_/B _59790_/X _59745_/X _59847_/Y _59848_/Y _84689_/D
+ sky130_fd_sc_hd__a41oi_4
X_78683_ _78682_/B _78682_/C _78682_/A _78684_/B sky130_fd_sc_hd__o21ai_4
X_75895_ _84493_/Q _84365_/Q _75895_/X sky130_fd_sc_hd__xor2_4
X_49602_ _49548_/A _49615_/C sky130_fd_sc_hd__buf_2
X_46814_ _46720_/A _46817_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_48_0_CLK clkbuf_8_49_0_CLK/A clkbuf_9_97_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_77634_ _77633_/B _77632_/Y _77629_/Y _77634_/Y sky130_fd_sc_hd__o21ai_4
X_62860_ _61541_/B _62858_/X _62859_/X _62889_/D _62860_/Y sky130_fd_sc_hd__nand4_4
X_74846_ _58153_/X _74846_/B _74846_/Y sky130_fd_sc_hd__nand2_4
X_47794_ _47794_/A _53249_/D sky130_fd_sc_hd__buf_2
X_49533_ _49537_/A _49537_/B _49522_/C _52746_/D _49533_/X sky130_fd_sc_hd__and4_4
X_61811_ _84724_/Q _61811_/X sky130_fd_sc_hd__buf_2
X_46745_ _46737_/A _46717_/B _46717_/C _46744_/X _46745_/X sky130_fd_sc_hd__and4_4
X_77565_ _81944_/Q _82200_/D _81912_/D sky130_fd_sc_hd__xor2_4
X_43957_ _43957_/A _43957_/B _43957_/X sky130_fd_sc_hd__and2_4
X_74777_ _74741_/X _74777_/B _74776_/Y _74777_/Y sky130_fd_sc_hd__nand3_4
X_62791_ _44173_/X _62791_/X sky130_fd_sc_hd__buf_2
X_71989_ _71970_/A _71989_/B _71989_/Y sky130_fd_sc_hd__nand2_4
X_79304_ _79286_/X _79304_/B _79304_/X sky130_fd_sc_hd__or2_4
X_76516_ _76514_/Y _76484_/Y _76515_/X _76516_/Y sky130_fd_sc_hd__o21ai_4
X_64530_ _79566_/A _63310_/X _64529_/Y _84237_/D sky130_fd_sc_hd__o21ai_4
X_42908_ _41681_/X _42900_/X _67556_/B _42901_/X _42908_/X sky130_fd_sc_hd__a2bb2o_4
X_49464_ _49454_/A _50987_/B _49464_/Y sky130_fd_sc_hd__nand2_4
X_61742_ _59766_/X _62130_/D sky130_fd_sc_hd__buf_2
X_73728_ _72723_/X _73728_/X sky130_fd_sc_hd__buf_2
X_46676_ _46676_/A _51779_/B sky130_fd_sc_hd__buf_2
X_77496_ _77496_/A _77495_/Y _77497_/A sky130_fd_sc_hd__and2_4
X_43888_ _41306_/X _43886_/X _67440_/B _43887_/X _43888_/X sky130_fd_sc_hd__a2bb2o_4
X_48415_ _48134_/X _47893_/A _48414_/X _48416_/A sky130_fd_sc_hd__o21ai_4
X_79235_ _79248_/C _79235_/B _79238_/A sky130_fd_sc_hd__nand2_4
X_45627_ _45734_/A _45627_/X sky130_fd_sc_hd__buf_2
X_64461_ _64454_/Y _64457_/Y _64460_/X _84844_/Q _64213_/X _64461_/Y
+ sky130_fd_sc_hd__o32ai_4
X_76447_ _76443_/Y _76422_/Y _76446_/X _76448_/B sky130_fd_sc_hd__o21ai_4
X_42839_ _42816_/X _42817_/X _41498_/X _66745_/B _42836_/X _42839_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49395_ _86395_/Q _49388_/X _49394_/Y _49395_/Y sky130_fd_sc_hd__o21ai_4
X_61673_ _61636_/A _61673_/B _61682_/C _61673_/Y sky130_fd_sc_hd__nand3_4
X_73659_ _73607_/A _85917_/Q _73659_/X sky130_fd_sc_hd__and2_4
X_66200_ _66197_/X _66199_/X _65304_/X _66200_/X sky130_fd_sc_hd__a21o_4
X_63412_ _63427_/A _61796_/X _63412_/X sky130_fd_sc_hd__and2_4
X_60624_ _60624_/A _60624_/X sky130_fd_sc_hd__buf_2
X_48346_ _86531_/Q _48333_/X _48345_/Y _48346_/Y sky130_fd_sc_hd__o21ai_4
X_67180_ _87354_/Q _67156_/X _67106_/X _67179_/X _67180_/X sky130_fd_sc_hd__a211o_4
X_79166_ _84787_/Q _82723_/D _79173_/A sky130_fd_sc_hd__nand2_4
X_45558_ _45558_/A _45560_/A sky130_fd_sc_hd__inv_2
X_76378_ _81266_/Q _81522_/D _76379_/B sky130_fd_sc_hd__xor2_4
X_64392_ _64377_/X _64392_/B _64391_/X _64392_/X sky130_fd_sc_hd__and3_4
X_66131_ _66128_/X _66130_/X _66057_/X _66134_/A sky130_fd_sc_hd__a21o_4
X_78117_ _82568_/Q _78125_/B _78130_/C sky130_fd_sc_hd__xor2_4
X_44509_ _44509_/A _44509_/Y sky130_fd_sc_hd__inv_2
X_63343_ _63339_/Y _63340_/X _63341_/X _63342_/X _63020_/A _63343_/Y
+ sky130_fd_sc_hd__o41ai_4
X_75329_ _75329_/A _75328_/X _80755_/D sky130_fd_sc_hd__xor2_4
X_48277_ _48275_/X _50322_/B _48277_/Y sky130_fd_sc_hd__nand2_4
X_60555_ _60555_/A _60555_/Y sky130_fd_sc_hd__inv_2
X_79097_ _79095_/X _79109_/A _82752_/Q _79097_/Y sky130_fd_sc_hd__a21oi_4
X_45489_ _44891_/X _45489_/X sky130_fd_sc_hd__buf_2
X_47228_ _47210_/A _47228_/B _47210_/C _52927_/D _47228_/X sky130_fd_sc_hd__and4_4
X_66062_ _65582_/X _66062_/B _65585_/X _66062_/Y sky130_fd_sc_hd__nand3_4
X_78048_ _77756_/Y _78048_/Y sky130_fd_sc_hd__inv_2
X_63274_ _63273_/X _63274_/Y sky130_fd_sc_hd__inv_2
X_60486_ _60488_/A _60488_/C _59691_/X _60414_/Y _60427_/A _60486_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_65013_ _64828_/X _85554_/Q _64829_/X _65012_/X _65013_/X sky130_fd_sc_hd__a211o_4
X_62225_ _60084_/A _62225_/X sky130_fd_sc_hd__buf_2
X_47159_ _47150_/A _52885_/B _47159_/Y sky130_fd_sc_hd__nand2_4
X_80010_ _79999_/X _80000_/A _80011_/D sky130_fd_sc_hd__nand2_4
X_69821_ _64696_/A _69820_/Y _69821_/Y sky130_fd_sc_hd__nor2_4
X_50170_ _86250_/Q _50162_/X _50169_/Y _50170_/Y sky130_fd_sc_hd__o21ai_4
X_62156_ _62154_/Y _62101_/X _62155_/Y _62156_/Y sky130_fd_sc_hd__a21oi_4
X_79999_ _79997_/X _80003_/B _79999_/X sky130_fd_sc_hd__xor2_4
X_61107_ _61107_/A _61107_/X sky130_fd_sc_hd__buf_2
X_69752_ _69766_/A _69752_/B _69752_/Y sky130_fd_sc_hd__nor2_4
X_66964_ _66606_/A _66964_/X sky130_fd_sc_hd__buf_2
X_62087_ _84834_/Q _62065_/B _62063_/X _62130_/D _62087_/Y sky130_fd_sc_hd__nand4_4
X_68703_ _88006_/Q _68650_/X _68651_/X _68702_/X _68703_/X sky130_fd_sc_hd__a211o_4
X_65915_ _65757_/A _65915_/X sky130_fd_sc_hd__buf_2
X_61038_ _61035_/X _61025_/X _61037_/Y _76981_/A _61020_/X _84533_/D
+ sky130_fd_sc_hd__o32a_4
X_81961_ _87345_/CLK _83889_/Q _81961_/Q sky130_fd_sc_hd__dfxtp_4
X_69683_ _69255_/Y _69644_/X _69672_/X _69682_/Y _69683_/X sky130_fd_sc_hd__a211o_4
X_66895_ _66757_/X _66886_/Y _66793_/X _66894_/Y _66895_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_392_0_CLK clkbuf_9_196_0_CLK/X _84606_/CLK sky130_fd_sc_hd__clkbuf_1
X_83700_ _85645_/CLK _70788_/Y _47115_/A sky130_fd_sc_hd__dfxtp_4
X_80912_ _80912_/CLK _84088_/Q _75694_/A sky130_fd_sc_hd__dfxtp_4
X_68634_ _68376_/X _68612_/X _68623_/Y _68633_/Y _68634_/X sky130_fd_sc_hd__a211o_4
X_53860_ _53848_/A _53860_/B _53860_/Y sky130_fd_sc_hd__nand2_4
X_65846_ _65804_/A _85861_/Q _65846_/X sky130_fd_sc_hd__and2_4
X_84680_ _84430_/CLK _59964_/Y _80241_/A sky130_fd_sc_hd__dfxtp_4
X_81892_ _82009_/CLK _77262_/X _82300_/D sky130_fd_sc_hd__dfxtp_4
X_52811_ _52818_/A _52818_/B _52789_/X _52811_/D _52811_/X sky130_fd_sc_hd__and4_4
X_83631_ _83630_/CLK _83631_/D _47622_/A sky130_fd_sc_hd__dfxtp_4
X_80843_ _80754_/CLK _80875_/Q _74916_/B sky130_fd_sc_hd__dfxtp_4
X_68565_ _68437_/A _73752_/A _68565_/X sky130_fd_sc_hd__and2_4
X_53791_ _53791_/A _48899_/Y _53791_/Y sky130_fd_sc_hd__nand2_4
X_65777_ _65777_/A _85866_/Q _65777_/X sky130_fd_sc_hd__and2_4
X_62989_ _62984_/X _62987_/X _62988_/Y _62989_/Y sky130_fd_sc_hd__a21oi_4
X_55530_ _45575_/A _55527_/X _44098_/X _55529_/X _55536_/C sky130_fd_sc_hd__a211o_4
X_67516_ _67039_/X _67516_/X sky130_fd_sc_hd__buf_2
X_86350_ _83703_/CLK _49643_/Y _86350_/Q sky130_fd_sc_hd__dfxtp_4
X_52742_ _52729_/X _52746_/B _52746_/C _52742_/D _52742_/X sky130_fd_sc_hd__and4_4
X_64728_ _64806_/A _64729_/A sky130_fd_sc_hd__buf_2
X_83562_ _83562_/CLK _71236_/Y _48704_/A sky130_fd_sc_hd__dfxtp_4
X_80774_ _80962_/CLK _80774_/D _80774_/Q sky130_fd_sc_hd__dfxtp_4
X_68496_ _73677_/A _68493_/X _68494_/X _68495_/Y _68496_/X sky130_fd_sc_hd__a211o_4
X_85301_ _85270_/CLK _56072_/Y _55879_/B sky130_fd_sc_hd__dfxtp_4
X_82513_ _82580_/CLK _82513_/D _82513_/Q sky130_fd_sc_hd__dfxtp_4
X_55461_ _55456_/X _55460_/X _44111_/X _55461_/X sky130_fd_sc_hd__a21o_4
X_67447_ _67305_/X _67436_/Y _67390_/X _67446_/Y _67447_/X sky130_fd_sc_hd__a211o_4
X_86281_ _86600_/CLK _86281_/D _86281_/Q sky130_fd_sc_hd__dfxtp_4
X_52673_ _52619_/A _52673_/X sky130_fd_sc_hd__buf_2
X_64659_ _64657_/X _83311_/Q _64600_/X _64658_/X _64659_/X sky130_fd_sc_hd__a211o_4
X_83493_ _83495_/CLK _71455_/X _83493_/Q sky130_fd_sc_hd__dfxtp_4
X_57200_ _57198_/X _56703_/X _57199_/Y _57200_/Y sky130_fd_sc_hd__a21oi_4
X_88020_ _87253_/CLK _88020_/D _88020_/Q sky130_fd_sc_hd__dfxtp_4
X_54412_ _54385_/A _54417_/B sky130_fd_sc_hd__buf_2
X_85232_ _85167_/CLK _56333_/Y _55836_/B sky130_fd_sc_hd__dfxtp_4
X_51624_ _85976_/Q _51621_/X _51623_/Y _51624_/Y sky130_fd_sc_hd__o21ai_4
X_58180_ _58171_/X _83490_/Q _58179_/Y _84914_/D sky130_fd_sc_hd__o21a_4
X_82444_ _82820_/CLK _79136_/X _82444_/Q sky130_fd_sc_hd__dfxtp_4
X_55392_ _55392_/A _55392_/B _55443_/D sky130_fd_sc_hd__xor2_4
X_67378_ _67333_/A _67378_/B _67378_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_330_0_CLK clkbuf_9_165_0_CLK/X _86322_/CLK sky130_fd_sc_hd__clkbuf_1
X_57131_ _57131_/A _57155_/D sky130_fd_sc_hd__inv_2
X_69117_ _69112_/X _69115_/X _69116_/X _69117_/X sky130_fd_sc_hd__a21o_4
X_54343_ _53097_/A _54344_/A sky130_fd_sc_hd__buf_2
X_66329_ _65863_/X _66276_/B _65867_/X _66329_/Y sky130_fd_sc_hd__nand3_4
X_85163_ _80671_/CLK _56524_/Y _56523_/C sky130_fd_sc_hd__dfxtp_4
X_51555_ _51545_/A _53080_/B _51555_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_960_0_CLK clkbuf_9_480_0_CLK/X _86554_/CLK sky130_fd_sc_hd__clkbuf_1
X_82375_ _85407_/CLK _82183_/Q _82375_/Q sky130_fd_sc_hd__dfxtp_4
X_84114_ _84115_/CLK _84114_/D _84114_/Q sky130_fd_sc_hd__dfxtp_4
X_50506_ _50506_/A _50506_/X sky130_fd_sc_hd__buf_2
X_57062_ _57056_/Y _57673_/A _57061_/Y _57062_/Y sky130_fd_sc_hd__nand3_4
X_81326_ _81492_/CLK _76326_/X _81702_/D sky130_fd_sc_hd__dfxtp_4
X_69048_ _69027_/A _69048_/B _69048_/X sky130_fd_sc_hd__and2_4
X_54274_ _54329_/A _54298_/B sky130_fd_sc_hd__buf_2
X_85094_ _85096_/CLK _57065_/X _45808_/A sky130_fd_sc_hd__dfxtp_4
X_51486_ _51211_/A _51491_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_451_0_CLK clkbuf_9_451_0_CLK/A clkbuf_9_451_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_56013_ _56030_/B _56013_/Y sky130_fd_sc_hd__inv_2
X_53225_ _51928_/X _53225_/X sky130_fd_sc_hd__buf_2
X_84045_ _88116_/CLK _84045_/D _81477_/D sky130_fd_sc_hd__dfxtp_4
X_50437_ _50464_/A _50437_/X sky130_fd_sc_hd__buf_2
X_81257_ _81257_/CLK _81257_/D _81257_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_345_0_CLK clkbuf_9_172_0_CLK/X _83703_/CLK sky130_fd_sc_hd__clkbuf_1
X_71010_ _71266_/A _71010_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_975_0_CLK clkbuf_9_487_0_CLK/X _83313_/CLK sky130_fd_sc_hd__clkbuf_1
X_80208_ _80204_/Y _80207_/Y _80208_/X sky130_fd_sc_hd__xor2_4
X_41170_ _41169_/X _41152_/X _68658_/B _41153_/X _41170_/X sky130_fd_sc_hd__a2bb2o_4
X_53156_ _53154_/Y _53137_/X _53155_/X _85687_/D sky130_fd_sc_hd__a21oi_4
X_50368_ _50381_/A _50368_/B _50368_/Y sky130_fd_sc_hd__nand2_4
X_81188_ _82692_/CLK _81188_/D _49179_/A sky130_fd_sc_hd__dfxtp_4
X_52107_ _52618_/A _52203_/A sky130_fd_sc_hd__buf_2
X_87804_ _88062_/CLK _87804_/D _73345_/A sky130_fd_sc_hd__dfxtp_4
X_80139_ _80136_/Y _80119_/Y _80138_/X _80139_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_466_0_CLK clkbuf_9_467_0_CLK/A clkbuf_9_466_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_53087_ _85699_/Q _53065_/X _53086_/Y _53087_/Y sky130_fd_sc_hd__o21ai_4
X_57964_ _57875_/X _85392_/Q _57963_/X _57964_/Y sky130_fd_sc_hd__o21ai_4
X_50299_ _50227_/A _50299_/X sky130_fd_sc_hd__buf_2
X_85996_ _85709_/CLK _85996_/D _85996_/Q sky130_fd_sc_hd__dfxtp_4
X_59703_ _59655_/X _59700_/Y _59680_/Y _59689_/Y _59702_/Y _59703_/Y
+ sky130_fd_sc_hd__a41oi_4
X_52038_ _51265_/A _52098_/B sky130_fd_sc_hd__buf_2
X_56915_ _56609_/X _56914_/Y _56915_/Y sky130_fd_sc_hd__nand2_4
X_87735_ _88002_/CLK _42756_/X _69042_/B sky130_fd_sc_hd__dfxtp_4
X_72961_ _72959_/X _85594_/Q _72839_/X _72960_/X _72961_/X sky130_fd_sc_hd__a211o_4
X_84947_ _83745_/CLK _57831_/Y _84947_/Q sky130_fd_sc_hd__dfxtp_4
X_57895_ _57883_/Y _57758_/X _57890_/X _57894_/X _57895_/Y sky130_fd_sc_hd__a22oi_4
X_74700_ _74673_/A _74700_/B _74700_/Y sky130_fd_sc_hd__nand2_4
X_71912_ _71891_/Y _71912_/Y sky130_fd_sc_hd__inv_2
X_59634_ _59634_/A _59634_/B _59662_/B _59648_/A sky130_fd_sc_hd__nand3_4
X_44860_ _44860_/A _86916_/D sky130_fd_sc_hd__inv_2
X_56846_ _56691_/A _56836_/Y _56843_/Y _56844_/X _56845_/Y _56846_/Y
+ sky130_fd_sc_hd__a32oi_4
X_75680_ _75680_/A _75679_/X _75684_/A sky130_fd_sc_hd__nand2_4
X_87666_ _81783_/CLK _87666_/D _67356_/B sky130_fd_sc_hd__dfxtp_4
X_72892_ _42555_/A _72892_/B _72892_/Y sky130_fd_sc_hd__nor2_4
X_84878_ _84849_/CLK _84878_/D _58322_/A sky130_fd_sc_hd__dfxtp_4
X_43811_ _43776_/A _43811_/X sky130_fd_sc_hd__buf_2
X_74631_ _56560_/X _45935_/X _56931_/X _83009_/Q _74630_/X _83009_/D
+ sky130_fd_sc_hd__a32o_4
X_86617_ _85974_/CLK _86617_/D _86617_/Q sky130_fd_sc_hd__dfxtp_4
X_71843_ _71072_/A _71714_/Y _71439_/C _70721_/A _71843_/X sky130_fd_sc_hd__and4_4
X_83829_ _83188_/CLK _83829_/D _83829_/Q sky130_fd_sc_hd__dfxtp_4
X_59565_ _59564_/A _59890_/B _59544_/D _60122_/C sky130_fd_sc_hd__nand3_4
X_44791_ _44512_/A _41887_/A _41402_/X _86953_/Q _44516_/A _44791_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56777_ _56777_/A _56777_/B _56777_/Y sky130_fd_sc_hd__nand2_4
X_87597_ _87070_/CLK _87597_/D _87597_/Q sky130_fd_sc_hd__dfxtp_4
X_53989_ _53921_/A _53989_/X sky130_fd_sc_hd__buf_2
X_46530_ _51360_/B _50850_/B sky130_fd_sc_hd__buf_2
X_58516_ _58492_/X _58513_/Y _58515_/Y _58516_/Y sky130_fd_sc_hd__a21oi_4
X_77350_ _77346_/Y _77290_/B _77349_/X _77351_/B sky130_fd_sc_hd__o21ai_4
X_43742_ _40908_/X _47846_/A _43741_/Y _43607_/A _43743_/A sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_10_913_0_CLK clkbuf_9_456_0_CLK/X _83133_/CLK sky130_fd_sc_hd__clkbuf_1
X_55728_ _45331_/A _55145_/A _55728_/Y sky130_fd_sc_hd__nand2_4
X_74562_ _74559_/X _74553_/X _56039_/Y _74554_/X _74562_/X sky130_fd_sc_hd__a211o_4
X_86548_ _86549_/CLK _86548_/D _66101_/B sky130_fd_sc_hd__dfxtp_4
X_40954_ _40931_/X _81726_/Q _40953_/X _40954_/Y sky130_fd_sc_hd__o21ai_4
X_71774_ _70502_/Y _71779_/A sky130_fd_sc_hd__buf_2
X_59496_ _64276_/C _63424_/B sky130_fd_sc_hd__buf_2
X_76301_ _76301_/A _81561_/Q _76301_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_2_0_CLK clkbuf_9_1_0_CLK/X _85269_/CLK sky130_fd_sc_hd__clkbuf_1
X_73513_ _44598_/Y _73420_/X _73512_/Y _73524_/C sky130_fd_sc_hd__a21o_4
X_70725_ _52781_/B _70699_/A _70724_/Y _70725_/Y sky130_fd_sc_hd__o21ai_4
X_46461_ _51326_/B _50816_/B sky130_fd_sc_hd__buf_2
X_58447_ _58423_/X _83478_/Q _58446_/Y _58447_/X sky130_fd_sc_hd__o21a_4
X_77281_ _77278_/X _82214_/Q _77279_/Y _77285_/C sky130_fd_sc_hd__nand3_4
Xclkbuf_5_30_0_CLK clkbuf_5_30_0_CLK/A clkbuf_6_61_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_43673_ _43673_/A _43673_/X sky130_fd_sc_hd__buf_2
X_55659_ _55656_/X _55657_/Y _55658_/Y _55659_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_404_0_CLK clkbuf_8_202_0_CLK/X clkbuf_9_404_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_74493_ _48656_/A _74501_/B _74501_/C _74493_/X sky130_fd_sc_hd__and3_4
X_86479_ _86191_/CLK _86479_/D _86479_/Q sky130_fd_sc_hd__dfxtp_4
X_40885_ _40885_/A _40885_/X sky130_fd_sc_hd__buf_2
X_48200_ _46485_/X _48201_/B sky130_fd_sc_hd__buf_2
X_79020_ _82826_/Q _79020_/B _79021_/B sky130_fd_sc_hd__xor2_4
X_45412_ _44891_/X _45412_/X sky130_fd_sc_hd__buf_2
X_76232_ _76232_/A _76232_/Y sky130_fd_sc_hd__inv_2
X_88218_ _88208_/CLK _88218_/D _88218_/Q sky130_fd_sc_hd__dfxtp_4
X_42624_ _73527_/A _69969_/B sky130_fd_sc_hd__inv_2
X_49180_ _49128_/X _48687_/A _49179_/Y _49181_/A sky130_fd_sc_hd__a21o_4
X_73444_ _87044_/Q _57092_/X _73443_/X _73444_/Y sky130_fd_sc_hd__o21ai_4
X_46392_ _46362_/A _52482_/B _46392_/Y sky130_fd_sc_hd__nand2_4
X_70656_ _70724_/A _70656_/B _70890_/C _70656_/D _70656_/Y sky130_fd_sc_hd__nand4_4
X_58378_ _58366_/X _83353_/Q _58377_/Y _84865_/D sky130_fd_sc_hd__o21a_4
X_48131_ _57637_/B _50378_/B sky130_fd_sc_hd__buf_2
XPHY_70 sky130_fd_sc_hd__decap_3
Xclkbuf_10_928_0_CLK clkbuf_9_464_0_CLK/X _88327_/CLK sky130_fd_sc_hd__clkbuf_1
X_45343_ _45709_/A _45343_/X sky130_fd_sc_hd__buf_2
X_57329_ _57280_/X _57325_/Y _57326_/Y _57328_/Y _57330_/A sky130_fd_sc_hd__a211o_4
XPHY_81 sky130_fd_sc_hd__decap_3
X_76163_ _76162_/Y _76163_/Y sky130_fd_sc_hd__inv_2
X_88149_ _88208_/CLK _41788_/Y _88149_/Q sky130_fd_sc_hd__dfxtp_4
X_42555_ _42555_/A _42555_/Y sky130_fd_sc_hd__inv_2
X_73375_ _69885_/B _44235_/X _72798_/X _73374_/Y _73375_/X sky130_fd_sc_hd__a211o_4
XPHY_92 sky130_fd_sc_hd__decap_3
X_70587_ _70586_/X _70588_/A sky130_fd_sc_hd__buf_2
X_75114_ _75100_/Y _75096_/A _75099_/A _75115_/A sky130_fd_sc_hd__o21a_4
X_41506_ _41481_/X _82328_/Q _41505_/X _41506_/Y sky130_fd_sc_hd__o21ai_4
X_60340_ _60249_/X _60325_/C _60367_/C _60229_/Y _60339_/Y _84628_/D
+ sky130_fd_sc_hd__a41oi_4
Xclkbuf_9_419_0_CLK clkbuf_9_419_0_CLK/A clkbuf_9_419_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_72326_ _72264_/X _85360_/Q _72325_/X _72326_/Y sky130_fd_sc_hd__o21ai_4
X_48062_ _48092_/A _52047_/B _48062_/Y sky130_fd_sc_hd__nand2_4
X_45274_ _44972_/A _45714_/A sky130_fd_sc_hd__buf_2
X_76094_ _76094_/A _76093_/Y _76099_/A sky130_fd_sc_hd__nor2_4
X_42486_ _42554_/A _42486_/X sky130_fd_sc_hd__buf_2
X_47013_ _47029_/A _47029_/B _47029_/C _52801_/D _47013_/X sky130_fd_sc_hd__and4_4
X_44225_ _65614_/A _44225_/B _57736_/A _44265_/D _44225_/Y sky130_fd_sc_hd__nor4_4
X_75045_ _75045_/A _75045_/B _75045_/X sky130_fd_sc_hd__xor2_4
X_79922_ _79922_/A _60145_/A _79924_/B sky130_fd_sc_hd__nand2_4
X_41437_ _41436_/Y _41437_/X sky130_fd_sc_hd__buf_2
X_60271_ _60271_/A _60271_/X sky130_fd_sc_hd__buf_2
X_72257_ _72143_/X _85366_/Q _72256_/X _72257_/Y sky130_fd_sc_hd__o21ai_4
X_62010_ _61708_/X _62010_/X sky130_fd_sc_hd__buf_2
Xclkbuf_6_4_0_CLK clkbuf_6_5_0_CLK/A clkbuf_6_4_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_71208_ _48820_/B _71190_/A _71207_/Y _71208_/Y sky130_fd_sc_hd__o21ai_4
X_44156_ _44012_/A _57776_/A sky130_fd_sc_hd__buf_2
X_79853_ _79819_/A _79818_/Y _79830_/X _79828_/Y _79850_/Y _79853_/X
+ sky130_fd_sc_hd__a2111o_4
X_41368_ _41367_/X _41362_/X _67707_/B _41363_/X _88228_/D sky130_fd_sc_hd__a2bb2o_4
X_72188_ _72188_/A _72162_/B _72188_/Y sky130_fd_sc_hd__nor2_4
X_43107_ _87573_/Q _43107_/Y sky130_fd_sc_hd__inv_2
X_78804_ _78802_/Y _78804_/B _78805_/B sky130_fd_sc_hd__xor2_4
X_71139_ _71145_/A _71141_/B sky130_fd_sc_hd__buf_2
X_48964_ _48964_/A _48963_/X _48964_/Y sky130_fd_sc_hd__nand2_4
X_44087_ _43950_/A _44087_/B _43975_/B _44088_/A sky130_fd_sc_hd__nor3_4
X_79784_ _79784_/A _79784_/B _79794_/B sky130_fd_sc_hd__xor2_4
X_41299_ _41298_/X _41283_/X _67399_/B _41284_/X _88241_/D sky130_fd_sc_hd__a2bb2o_4
X_76996_ _60959_/C _62302_/C _76996_/X sky130_fd_sc_hd__xor2_4
X_47915_ _48438_/B _47915_/B _47915_/Y sky130_fd_sc_hd__nand2_4
X_43038_ _43146_/A _43038_/X sky130_fd_sc_hd__buf_2
X_78735_ _78735_/A _78735_/Y sky130_fd_sc_hd__inv_2
X_63961_ _63959_/X _63913_/X _63960_/Y _84284_/D sky130_fd_sc_hd__a21oi_4
X_75947_ _81701_/D _75940_/B _75947_/Y sky130_fd_sc_hd__nand2_4
X_48895_ _48890_/Y _48880_/X _48894_/X _48895_/Y sky130_fd_sc_hd__a21oi_4
X_65700_ _65198_/A _65700_/X sky130_fd_sc_hd__buf_2
X_62912_ _62906_/X _62886_/X _62907_/Y _62909_/Y _62911_/X _62912_/X
+ sky130_fd_sc_hd__a41o_4
X_47846_ _47846_/A _47846_/X sky130_fd_sc_hd__buf_2
X_66680_ _87375_/Q _66678_/X _66629_/X _66679_/X _66680_/X sky130_fd_sc_hd__a211o_4
X_78666_ _78665_/X _78666_/Y sky130_fd_sc_hd__inv_2
X_63892_ _61876_/X _63876_/B _63860_/C _63892_/D _63892_/Y sky130_fd_sc_hd__nand4_4
X_75878_ _80897_/D _75878_/B _75880_/A sky130_fd_sc_hd__nand2_4
X_65631_ _65628_/X _65631_/B _65630_/X _65631_/Y sky130_fd_sc_hd__nand3_4
X_77617_ _77616_/X _77619_/B sky130_fd_sc_hd__inv_2
X_62843_ _63562_/A _60337_/D _62842_/Y _62843_/X sky130_fd_sc_hd__o21a_4
X_74829_ _74829_/A _46141_/A _74829_/Y sky130_fd_sc_hd__nand2_4
X_47777_ _47804_/A _47777_/B _47777_/C _53238_/D _47777_/X sky130_fd_sc_hd__and4_4
X_78597_ _78608_/A _82678_/D _78597_/X sky130_fd_sc_hd__xor2_4
X_44989_ _44989_/A _44990_/A sky130_fd_sc_hd__inv_2
X_49516_ _49537_/A _49516_/B _49493_/X _52730_/D _49516_/X sky130_fd_sc_hd__and4_4
X_68350_ _69906_/A _87251_/Q _68350_/X sky130_fd_sc_hd__and2_4
X_46728_ _46727_/Y _46728_/X sky130_fd_sc_hd__buf_2
X_65562_ _65334_/X _86200_/Q _65517_/X _65561_/X _65562_/X sky130_fd_sc_hd__a211o_4
X_77548_ _81943_/Q _82199_/D _81911_/D sky130_fd_sc_hd__xor2_4
X_62774_ _62773_/X _62762_/B _61891_/X _62774_/Y sky130_fd_sc_hd__nand3_4
X_67301_ _87105_/Q _67230_/X _67278_/X _67300_/X _67301_/X sky130_fd_sc_hd__a211o_4
X_64513_ _64494_/A _63312_/B _64207_/A _64513_/X sky130_fd_sc_hd__and3_4
X_61725_ _61720_/Y _61699_/X _61724_/Y _84457_/D sky130_fd_sc_hd__a21oi_4
X_49447_ _49447_/A _49447_/B _49447_/C _52661_/D _49447_/X sky130_fd_sc_hd__and4_4
X_68281_ _68254_/X _67726_/Y _68268_/X _68280_/Y _68281_/X sky130_fd_sc_hd__a211o_4
X_46659_ _46670_/A _46682_/B _46659_/C _51772_/D _46659_/X sky130_fd_sc_hd__and4_4
X_65493_ _65428_/X _83077_/Q _65407_/X _65492_/X _65494_/B sky130_fd_sc_hd__a211o_4
X_77479_ _77478_/B _77477_/Y _77478_/A _77479_/X sky130_fd_sc_hd__o21a_4
X_79218_ _79215_/X _79236_/A _79213_/Y _79218_/X sky130_fd_sc_hd__a21o_4
X_67232_ _87108_/Q _67230_/X _67160_/X _67231_/X _67232_/X sky130_fd_sc_hd__a211o_4
X_64444_ _84246_/Q _64429_/X _64443_/X _64444_/X sky130_fd_sc_hd__a21o_4
X_49378_ _49405_/A _49378_/X sky130_fd_sc_hd__buf_2
X_61656_ _61656_/A _61598_/X _61677_/C _61563_/D _61657_/A sky130_fd_sc_hd__nand4_4
X_80490_ _80489_/B _80489_/A _80490_/X sky130_fd_sc_hd__and2_4
X_48329_ _48329_/A _50372_/B sky130_fd_sc_hd__buf_2
X_60607_ _60607_/A _60606_/X _60420_/A _60430_/Y _60608_/A sky130_fd_sc_hd__and4_4
X_67163_ _67159_/X _67162_/X _67015_/X _67163_/Y sky130_fd_sc_hd__a21oi_4
X_79149_ _79149_/A _61434_/C _79149_/X sky130_fd_sc_hd__xor2_4
X_64375_ _59415_/A _64418_/B _64375_/Y sky130_fd_sc_hd__nor2_4
X_61587_ _59834_/A _61587_/B _79136_/B _61587_/X sky130_fd_sc_hd__or3_4
X_66114_ _57788_/X _73904_/B _66114_/X sky130_fd_sc_hd__and2_4
X_51340_ _51340_/A _51842_/A sky130_fd_sc_hd__buf_2
X_63326_ _63326_/A _63344_/B _60588_/X _63344_/D _63326_/X sky130_fd_sc_hd__or4_4
X_82160_ _81224_/CLK _84152_/Q _82160_/Q sky130_fd_sc_hd__dfxtp_4
X_60538_ _60588_/A _63301_/C sky130_fd_sc_hd__buf_2
X_67094_ _67093_/X _67095_/A sky130_fd_sc_hd__buf_2
X_81111_ _81111_/CLK _79780_/Y _81111_/Q sky130_fd_sc_hd__dfxtp_4
X_66045_ _66020_/X _66043_/Y _66044_/Y _66045_/Y sky130_fd_sc_hd__o21ai_4
X_51271_ _51269_/Y _51263_/X _51270_/X _51271_/Y sky130_fd_sc_hd__a21oi_4
X_63257_ _63255_/X _62987_/X _63256_/Y _84340_/D sky130_fd_sc_hd__a21oi_4
X_82091_ _82008_/CLK _82091_/D _77065_/A sky130_fd_sc_hd__dfxtp_4
X_60469_ _60472_/A _60469_/X sky130_fd_sc_hd__buf_2
X_53010_ _53065_/A _53010_/X sky130_fd_sc_hd__buf_2
X_50222_ _51074_/A _50222_/X sky130_fd_sc_hd__buf_2
X_62208_ _62237_/A _62522_/B sky130_fd_sc_hd__buf_2
X_81042_ _81070_/CLK _81042_/D _81042_/Q sky130_fd_sc_hd__dfxtp_4
X_63188_ _57757_/A _64314_/A sky130_fd_sc_hd__buf_2
X_69804_ _69804_/A _69804_/Y sky130_fd_sc_hd__inv_2
X_50153_ _50153_/A _50153_/B _50153_/Y sky130_fd_sc_hd__nand2_4
X_62139_ _61649_/B _62161_/B _62128_/C _61706_/X _62139_/Y sky130_fd_sc_hd__nand4_4
X_85850_ _85558_/CLK _52302_/Y _85850_/Q sky130_fd_sc_hd__dfxtp_4
X_67996_ _81478_/D _67925_/X _67995_/X _67996_/X sky130_fd_sc_hd__a21bo_4
X_84801_ _86713_/CLK _84801_/D _84801_/Q sky130_fd_sc_hd__dfxtp_4
X_69735_ _69735_/A _69734_/Y _69735_/Y sky130_fd_sc_hd__nor2_4
X_50084_ _50084_/A _48944_/B _50084_/Y sky130_fd_sc_hd__nand2_4
X_54961_ _54961_/A _47536_/A _54961_/Y sky130_fd_sc_hd__nand2_4
X_66947_ _64608_/A _66947_/X sky130_fd_sc_hd__buf_2
X_85781_ _82956_/CLK _85781_/D _85781_/Q sky130_fd_sc_hd__dfxtp_4
X_82993_ _82993_/CLK _82993_/D _82993_/Q sky130_fd_sc_hd__dfxtp_4
X_56700_ _56698_/Y _56842_/A _56700_/C _56676_/Y _56700_/Y sky130_fd_sc_hd__nor4_4
X_87520_ _87520_/CLK _43246_/Y _87520_/Q sky130_fd_sc_hd__dfxtp_4
X_53912_ _53898_/A _49144_/A _53912_/Y sky130_fd_sc_hd__nand2_4
X_84732_ _84732_/CLK _59441_/X _84732_/Q sky130_fd_sc_hd__dfxtp_4
X_81944_ _82133_/CLK _81944_/D _81944_/Q sky130_fd_sc_hd__dfxtp_4
X_57680_ _57680_/A _57666_/B _57680_/Y sky130_fd_sc_hd__nor2_4
X_69666_ _69092_/A _88332_/Q _69666_/X sky130_fd_sc_hd__and2_4
X_54892_ _54892_/A _54892_/X sky130_fd_sc_hd__buf_2
X_66878_ _66642_/A _66878_/X sky130_fd_sc_hd__buf_2
X_56631_ _56587_/X _56630_/X _55529_/B _56590_/X _85142_/D sky130_fd_sc_hd__a2bb2o_4
X_68617_ _68617_/A _68617_/X sky130_fd_sc_hd__buf_2
X_87451_ _87446_/CLK _43381_/X _87451_/Q sky130_fd_sc_hd__dfxtp_4
X_53843_ _53793_/A _53844_/A sky130_fd_sc_hd__buf_2
X_65829_ _65700_/X _65827_/Y _65828_/Y _65829_/Y sky130_fd_sc_hd__o21ai_4
X_84663_ _84672_/CLK _60093_/X _84663_/Q sky130_fd_sc_hd__dfxtp_4
X_81875_ _81857_/CLK _78066_/X _81875_/Q sky130_fd_sc_hd__dfxtp_4
X_69597_ _69586_/A _69597_/B _69597_/X sky130_fd_sc_hd__and2_4
X_86402_ _86733_/CLK _86402_/D _86402_/Q sky130_fd_sc_hd__dfxtp_4
X_59350_ _59286_/X _86053_/Q _59349_/X _59350_/Y sky130_fd_sc_hd__o21ai_4
X_83614_ _85558_/CLK _71081_/Y _83614_/Q sky130_fd_sc_hd__dfxtp_4
X_56562_ _44135_/X _56774_/C sky130_fd_sc_hd__buf_2
X_68548_ _68544_/X _68547_/X _58002_/A _68548_/X sky130_fd_sc_hd__a21o_4
X_80826_ _81065_/CLK _80826_/D _80826_/Q sky130_fd_sc_hd__dfxtp_4
X_87382_ _87382_/CLK _87382_/D _87382_/Q sky130_fd_sc_hd__dfxtp_4
X_53774_ _48702_/A _53774_/B _53774_/C _53774_/X sky130_fd_sc_hd__and3_4
X_84594_ _84606_/CLK _60585_/X _79134_/A sky130_fd_sc_hd__dfxtp_4
X_50986_ _50982_/Y _50983_/X _50985_/X _86095_/D sky130_fd_sc_hd__a21oi_4
X_58301_ _63694_/B _58344_/B _58301_/Y sky130_fd_sc_hd__nor2_4
X_55513_ _55512_/X _55513_/X sky130_fd_sc_hd__buf_2
X_86333_ _86651_/CLK _49735_/Y _86333_/Q sky130_fd_sc_hd__dfxtp_4
X_52725_ _52723_/Y _52702_/X _52724_/X _52725_/Y sky130_fd_sc_hd__a21oi_4
X_59281_ _59256_/A _86346_/Q _59281_/Y sky130_fd_sc_hd__nor2_4
X_83545_ _85630_/CLK _83545_/D _83545_/Q sky130_fd_sc_hd__dfxtp_4
X_56493_ _56060_/X _56483_/X _56492_/Y _85175_/D sky130_fd_sc_hd__o21ai_4
X_80757_ _80804_/CLK _75358_/X _80757_/Q sky130_fd_sc_hd__dfxtp_4
X_68479_ _68479_/A _68553_/A sky130_fd_sc_hd__buf_2
X_70510_ _57651_/Y _70501_/X _70509_/Y _83761_/D sky130_fd_sc_hd__o21ai_4
X_58232_ _58232_/A _58232_/X sky130_fd_sc_hd__buf_2
X_55444_ _55430_/Y _55435_/X _55443_/Y _55444_/Y sky130_fd_sc_hd__a21oi_4
X_86264_ _85558_/CLK _50102_/Y _86264_/Q sky130_fd_sc_hd__dfxtp_4
X_40670_ _40585_/A _40670_/X sky130_fd_sc_hd__buf_2
X_52656_ _52515_/X _52656_/X sky130_fd_sc_hd__buf_2
X_71490_ _71487_/X _83481_/Q _71489_/X _71490_/X sky130_fd_sc_hd__a21o_4
X_83476_ _83476_/CLK _83476_/D _83476_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_602 sky130_fd_sc_hd__decap_3
X_80688_ _81038_/CLK _80688_/D _75269_/A sky130_fd_sc_hd__dfxtp_4
XPHY_613 sky130_fd_sc_hd__decap_3
X_88003_ _88002_/CLK _88003_/D _88003_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_624 sky130_fd_sc_hd__decap_3
Xclkbuf_10_51_0_CLK clkbuf_9_25_0_CLK/X _85039_/CLK sky130_fd_sc_hd__clkbuf_1
X_85215_ _85249_/CLK _85215_/D _56381_/C sky130_fd_sc_hd__dfxtp_4
X_51607_ _51033_/A _51608_/A sky130_fd_sc_hd__buf_2
X_70441_ _71196_/A _71194_/C sky130_fd_sc_hd__buf_2
X_58163_ _63054_/A _64257_/A sky130_fd_sc_hd__buf_2
XPHY_635 sky130_fd_sc_hd__decap_3
X_82427_ _83507_/CLK _82427_/D _78680_/A sky130_fd_sc_hd__dfxtp_4
X_55375_ _55375_/A _55374_/Y _55375_/Y sky130_fd_sc_hd__nor2_4
X_86195_ _86191_/CLK _86195_/D _86195_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_646 sky130_fd_sc_hd__decap_3
X_52587_ _85791_/Q _52575_/X _52586_/Y _52587_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_390_0_CLK clkbuf_9_391_0_CLK/A clkbuf_9_390_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_657 sky130_fd_sc_hd__decap_3
XPHY_668 sky130_fd_sc_hd__decap_3
X_57114_ _56613_/X _57106_/X _57113_/Y _85081_/D sky130_fd_sc_hd__a21oi_4
X_42340_ _42340_/A _42340_/Y sky130_fd_sc_hd__inv_2
X_54326_ _54324_/Y _54311_/X _54325_/X _85463_/D sky130_fd_sc_hd__a21oi_4
XPHY_679 sky130_fd_sc_hd__decap_3
X_73160_ _73381_/A _86482_/Q _73160_/X sky130_fd_sc_hd__and2_4
X_85146_ _85144_/CLK _85146_/D _85146_/Q sky130_fd_sc_hd__dfxtp_4
X_51538_ _51536_/Y _51531_/X _51537_/X _85992_/D sky130_fd_sc_hd__a21oi_4
X_70372_ _51358_/B _70364_/X _70371_/Y _70372_/Y sky130_fd_sc_hd__o21ai_4
X_58094_ _58094_/A _58599_/A sky130_fd_sc_hd__buf_2
X_82358_ _84981_/CLK _77199_/X _47955_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_284_0_CLK clkbuf_9_142_0_CLK/X _84945_/CLK sky130_fd_sc_hd__clkbuf_1
X_72111_ _83282_/Q _72066_/X _72110_/Y _72111_/Y sky130_fd_sc_hd__o21ai_4
X_57045_ _57044_/Y _85097_/D sky130_fd_sc_hd__inv_2
X_81309_ _81627_/CLK _76997_/X _81277_/D sky130_fd_sc_hd__dfxtp_4
X_42271_ _42258_/A _42271_/X sky130_fd_sc_hd__buf_2
X_54257_ _54961_/A _53086_/B _54257_/Y sky130_fd_sc_hd__nand2_4
X_73091_ _73062_/X _86197_/Q _72955_/X _73090_/X _73091_/X sky130_fd_sc_hd__a211o_4
X_85077_ _85042_/CLK _85077_/D _85077_/Q sky130_fd_sc_hd__dfxtp_4
X_51469_ _51481_/A _52995_/B _51469_/Y sky130_fd_sc_hd__nand2_4
X_82289_ _82339_/CLK _81913_/Q _41026_/A sky130_fd_sc_hd__dfxtp_4
X_44010_ _44010_/A _44247_/A _44152_/A sky130_fd_sc_hd__nand2_4
Xclkbuf_10_66_0_CLK clkbuf_9_33_0_CLK/X _83016_/CLK sky130_fd_sc_hd__clkbuf_1
X_53208_ _53206_/Y _53189_/X _53207_/X _85677_/D sky130_fd_sc_hd__a21oi_4
X_41222_ _41221_/Y _41222_/Y sky130_fd_sc_hd__inv_2
X_72042_ _46610_/A _74453_/A sky130_fd_sc_hd__buf_2
X_84028_ _86807_/CLK _84028_/D _84028_/Q sky130_fd_sc_hd__dfxtp_4
X_54188_ _54184_/A _47394_/Y _54188_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_212_0_CLK clkbuf_8_213_0_CLK/A clkbuf_9_424_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_41153_ _40989_/A _41153_/X sky130_fd_sc_hd__buf_2
X_53139_ _53139_/A _53133_/B _53133_/C _53139_/D _53139_/X sky130_fd_sc_hd__and4_4
X_76850_ _76837_/A _76844_/A _76850_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_299_0_CLK clkbuf_9_149_0_CLK/X _84329_/CLK sky130_fd_sc_hd__clkbuf_1
X_58996_ _58920_/A _86369_/Q _58996_/Y sky130_fd_sc_hd__nor2_4
X_75801_ _81019_/Q _80891_/D _80987_/D sky130_fd_sc_hd__xor2_4
X_57947_ _57947_/A _57947_/X sky130_fd_sc_hd__buf_2
X_45961_ _45961_/A _45961_/Y sky130_fd_sc_hd__inv_2
X_41084_ _41084_/A _41084_/Y sky130_fd_sc_hd__inv_2
X_76781_ _76776_/Y _76780_/Y _76781_/Y sky130_fd_sc_hd__nand2_4
X_73993_ _44126_/X _66166_/B _73993_/X sky130_fd_sc_hd__and2_4
X_85979_ _85692_/CLK _51610_/Y _85979_/Q sky130_fd_sc_hd__dfxtp_4
X_47700_ _81231_/Q _47701_/A sky130_fd_sc_hd__inv_2
X_78520_ _82512_/Q _82768_/D _78520_/X sky130_fd_sc_hd__xor2_4
X_44912_ _55976_/B _44874_/X _44875_/X _44912_/X sky130_fd_sc_hd__o21a_4
X_75732_ _75732_/A _75734_/A sky130_fd_sc_hd__inv_2
X_87718_ _87150_/CLK _42789_/X _87718_/Q sky130_fd_sc_hd__dfxtp_4
X_48680_ _48680_/A _48657_/B _48894_/C _48680_/X sky130_fd_sc_hd__and3_4
X_72944_ _72725_/A _72944_/X sky130_fd_sc_hd__buf_2
X_45892_ _45891_/X _45893_/C sky130_fd_sc_hd__buf_2
Xclkbuf_8_227_0_CLK clkbuf_8_227_0_CLK/A clkbuf_9_455_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_57878_ _58020_/A _57878_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_222_0_CLK clkbuf_9_111_0_CLK/X _84559_/CLK sky130_fd_sc_hd__clkbuf_1
X_47631_ _47631_/A _47632_/A sky130_fd_sc_hd__inv_2
X_59617_ _59893_/C _59905_/B sky130_fd_sc_hd__buf_2
X_78451_ _78439_/Y _78423_/Y _78450_/A _78451_/Y sky130_fd_sc_hd__a21oi_4
X_44843_ _41730_/Y _44838_/X _86924_/Q _44839_/X _86924_/D sky130_fd_sc_hd__a2bb2o_4
X_56829_ _56738_/X _56828_/Y _45888_/A _56829_/X sky130_fd_sc_hd__o21a_4
X_75663_ _75649_/Y _75650_/Y _80906_/Q _75662_/Y _75663_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_10_852_0_CLK clkbuf_9_426_0_CLK/X _82961_/CLK sky130_fd_sc_hd__clkbuf_1
X_87649_ _87646_/CLK _87649_/D _87649_/Q sky130_fd_sc_hd__dfxtp_4
X_72875_ _45931_/X _85597_/Q _56933_/X _72874_/X _72875_/X sky130_fd_sc_hd__a211o_4
X_77402_ _77397_/Y _77374_/B _77401_/X _77403_/B sky130_fd_sc_hd__o21ai_4
X_74614_ _74614_/A _74614_/X sky130_fd_sc_hd__buf_2
X_47562_ _47561_/Y _53122_/B sky130_fd_sc_hd__buf_2
X_71826_ _70773_/A _71826_/X sky130_fd_sc_hd__buf_2
X_59548_ _60183_/A _59552_/C sky130_fd_sc_hd__buf_2
X_78382_ _78397_/B _78382_/B _82759_/D sky130_fd_sc_hd__xor2_4
X_44774_ _44618_/A _44774_/X sky130_fd_sc_hd__buf_2
X_75594_ _75590_/X _75594_/B _75591_/Y _75594_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_9_343_0_CLK clkbuf_9_343_0_CLK/A clkbuf_9_343_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_41986_ _88081_/Q _41986_/Y sky130_fd_sc_hd__inv_2
X_49301_ _49205_/A _49302_/A sky130_fd_sc_hd__buf_2
X_46513_ _86730_/Q _46430_/X _46512_/Y _46513_/Y sky130_fd_sc_hd__o21ai_4
X_77333_ _77333_/A _77334_/B sky130_fd_sc_hd__inv_2
X_43725_ _40873_/X _43716_/X _69838_/B _43718_/X _43726_/A sky130_fd_sc_hd__a2bb2o_4
X_74545_ _74541_/A _46215_/B _74545_/C _74545_/Y sky130_fd_sc_hd__nand3_4
X_40937_ _40937_/A _41119_/A _40937_/X sky130_fd_sc_hd__or2_4
X_47493_ _47493_/A _47494_/A sky130_fd_sc_hd__inv_2
X_71757_ _52959_/B _71736_/X _71756_/Y _83387_/D sky130_fd_sc_hd__o21ai_4
X_59479_ _59462_/X _83433_/Q _59478_/Y _84721_/D sky130_fd_sc_hd__o21a_4
Xclkbuf_10_237_0_CLK clkbuf_9_118_0_CLK/X _81834_/CLK sky130_fd_sc_hd__clkbuf_1
X_49232_ _49232_/A _51261_/B _49232_/Y sky130_fd_sc_hd__nand2_4
X_61510_ _84818_/Q _61510_/X sky130_fd_sc_hd__buf_2
X_46444_ _86736_/Q _46292_/X _46443_/Y _46444_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_867_0_CLK clkbuf_9_433_0_CLK/X _86560_/CLK sky130_fd_sc_hd__clkbuf_1
X_70708_ _70585_/X _70703_/X _70710_/C _70710_/D _70708_/Y sky130_fd_sc_hd__nand4_4
X_77264_ _77264_/A _77264_/Y sky130_fd_sc_hd__inv_2
X_43656_ _43685_/A _43656_/X sky130_fd_sc_hd__buf_2
X_62490_ _61561_/A _62566_/B _62490_/C _62566_/D _62490_/Y sky130_fd_sc_hd__nand4_4
X_74476_ _74490_/A _48615_/A _74476_/Y sky130_fd_sc_hd__nand2_4
X_40868_ _40835_/X _40836_/X _40866_/X _69826_/B _40867_/X _40869_/A
+ sky130_fd_sc_hd__o32ai_4
X_71688_ _71576_/X _71626_/B _71289_/B _71688_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_10_19_0_CLK clkbuf_9_9_0_CLK/X _83022_/CLK sky130_fd_sc_hd__clkbuf_1
X_79003_ _82824_/Q _82536_/Q _79003_/Y sky130_fd_sc_hd__xnor2_4
X_76215_ _76215_/A _76215_/Y sky130_fd_sc_hd__inv_2
X_42607_ _42607_/A _42607_/Y sky130_fd_sc_hd__inv_2
X_61441_ _61380_/A _61452_/D sky130_fd_sc_hd__buf_2
X_73427_ _73355_/X _85575_/Q _73284_/X _73426_/X _73427_/X sky130_fd_sc_hd__a211o_4
X_49163_ _49163_/A _53919_/B sky130_fd_sc_hd__buf_2
X_46375_ _46370_/Y _46346_/X _46374_/Y _46375_/Y sky130_fd_sc_hd__a21boi_4
X_70639_ _70585_/X _70639_/B _70620_/C _70638_/X _70639_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_9_358_0_CLK clkbuf_8_179_0_CLK/X clkbuf_9_358_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_77195_ _77202_/B _77202_/C _77198_/A sky130_fd_sc_hd__nand2_4
X_43587_ _43587_/A _43587_/Y sky130_fd_sc_hd__inv_2
X_40799_ _40798_/X _40793_/X _88333_/Q _40794_/X _88333_/D sky130_fd_sc_hd__a2bb2o_4
X_48114_ _83534_/Q _53593_/B sky130_fd_sc_hd__inv_2
X_45326_ _45252_/A _45326_/X sky130_fd_sc_hd__buf_2
X_64160_ _62151_/X _64182_/B _64095_/C _64182_/D _64160_/Y sky130_fd_sc_hd__nand4_4
X_76146_ _81729_/D _76146_/B _76149_/C sky130_fd_sc_hd__xnor2_4
X_42538_ _42556_/A _42538_/X sky130_fd_sc_hd__buf_2
X_49094_ _53886_/B _52367_/B sky130_fd_sc_hd__buf_2
X_61372_ _61370_/X _61349_/X _61371_/Y _84486_/D sky130_fd_sc_hd__a21oi_4
X_73358_ _73354_/X _73357_/X _73262_/X _73362_/A sky130_fd_sc_hd__a21o_4
X_63111_ _63106_/Y _63108_/X _63109_/X _63110_/X _63067_/X _63111_/Y
+ sky130_fd_sc_hd__o41ai_4
X_48045_ _48043_/X _82349_/Q _48044_/Y _48046_/A sky130_fd_sc_hd__o21ai_4
X_60323_ _59756_/A _60323_/X sky130_fd_sc_hd__buf_2
X_72309_ _72258_/X _85682_/Q _72308_/X _72309_/X sky130_fd_sc_hd__o21a_4
X_45257_ _45257_/A _45257_/Y sky130_fd_sc_hd__inv_2
X_64091_ _64467_/C _64091_/B _64091_/C _64091_/D _64094_/B sky130_fd_sc_hd__nand4_4
X_76077_ _76067_/Y _76076_/X _76077_/Y sky130_fd_sc_hd__nand2_4
X_42469_ _42468_/Y _87855_/D sky130_fd_sc_hd__inv_2
X_73289_ _73214_/X _83061_/Q _73238_/X _73288_/X _73290_/B sky130_fd_sc_hd__a211o_4
X_44208_ _44204_/Y _44067_/B _58547_/A _44208_/X sky130_fd_sc_hd__and3_4
X_75028_ _80955_/Q _75028_/B _75028_/X sky130_fd_sc_hd__xor2_4
X_79905_ _79903_/Y _79911_/A _79909_/A sky130_fd_sc_hd__nand2_4
X_63042_ _63036_/Y _63038_/X _63039_/X _63041_/X _63020_/X _63042_/Y
+ sky130_fd_sc_hd__o41ai_4
X_60254_ _60159_/A _60254_/B _60255_/A sky130_fd_sc_hd__nor2_4
X_45188_ _56243_/C _45147_/X _45187_/X _45188_/Y sky130_fd_sc_hd__o21ai_4
X_44139_ _44024_/A _44139_/X sky130_fd_sc_hd__buf_2
X_67850_ _67847_/X _67849_/X _67709_/X _67850_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_805_0_CLK clkbuf_9_402_0_CLK/X _82498_/CLK sky130_fd_sc_hd__clkbuf_1
X_79836_ _79836_/A _72165_/A _79836_/X sky130_fd_sc_hd__xor2_4
X_60185_ _59613_/Y _60172_/A _60182_/Y _61278_/B _60185_/X sky130_fd_sc_hd__and4_4
X_49996_ _49993_/Y _49977_/X _49995_/X _86285_/D sky130_fd_sc_hd__a21oi_4
X_66801_ _57866_/A _66801_/X sky130_fd_sc_hd__buf_2
X_48947_ _48947_/A _48976_/A _48947_/Y sky130_fd_sc_hd__nor2_4
X_79767_ _79745_/A _79767_/B _79767_/Y sky130_fd_sc_hd__nand2_4
X_67781_ _84055_/Q _67688_/X _67780_/X _84055_/D sky130_fd_sc_hd__a21bo_4
X_64993_ _64934_/X _83299_/Q _64991_/X _64992_/X _64993_/X sky130_fd_sc_hd__a211o_4
X_76979_ _84531_/Q _62541_/C _76979_/X sky130_fd_sc_hd__xor2_4
X_69520_ _68300_/X _69520_/X sky130_fd_sc_hd__buf_2
X_78718_ _78713_/X _78716_/Y _78718_/C _78718_/Y sky130_fd_sc_hd__nand3_4
X_66732_ _80923_/D _66614_/X _66731_/X _66732_/X sky130_fd_sc_hd__a21bo_4
X_63944_ _63960_/A _63960_/B _63944_/C _63944_/Y sky130_fd_sc_hd__nor3_4
X_48878_ _48695_/A _48878_/B _48878_/Y sky130_fd_sc_hd__nand2_4
X_79698_ _79692_/A _79692_/B _79697_/Y _79702_/A sky130_fd_sc_hd__a21boi_4
X_69451_ _83923_/Q _69439_/X _69450_/X _83923_/D sky130_fd_sc_hd__a21bo_4
X_47829_ _47829_/A _57491_/C sky130_fd_sc_hd__buf_2
X_66663_ _87951_/Q _66639_/X _66531_/X _66662_/X _66663_/X sky130_fd_sc_hd__a211o_4
X_78649_ _78645_/Y _78649_/B _78648_/Y _78654_/A sky130_fd_sc_hd__or3_4
X_63875_ _64032_/A _63876_/B sky130_fd_sc_hd__buf_2
X_68402_ _68402_/A _68402_/X sky130_fd_sc_hd__buf_2
X_65614_ _65614_/A _65614_/X sky130_fd_sc_hd__buf_2
X_50840_ _52533_/A _50825_/B _50830_/C _50840_/X sky130_fd_sc_hd__and3_4
X_62826_ _62824_/X _62779_/X _62825_/Y _84379_/D sky130_fd_sc_hd__a21oi_4
X_81660_ _81660_/CLK _81692_/Q _81660_/Q sky130_fd_sc_hd__dfxtp_4
X_69382_ _88033_/Q _69368_/X _69232_/X _69381_/X _69382_/X sky130_fd_sc_hd__a211o_4
X_66594_ _69183_/A _66594_/X sky130_fd_sc_hd__buf_2
X_80611_ _84775_/Q _84167_/Q _80611_/Y sky130_fd_sc_hd__nand2_4
X_68333_ _68301_/X _68027_/Y _68326_/X _68332_/Y _68333_/X sky130_fd_sc_hd__a211o_4
X_65545_ _65533_/X _65543_/Y _65544_/Y _65545_/Y sky130_fd_sc_hd__o21ai_4
X_50771_ _50771_/A _46356_/X _50771_/Y sky130_fd_sc_hd__nand2_4
X_62757_ _62766_/A _62766_/B _75915_/B _62757_/Y sky130_fd_sc_hd__nor3_4
X_81591_ _81482_/CLK _84191_/Q _76845_/A sky130_fd_sc_hd__dfxtp_4
X_52510_ _52507_/Y _52496_/X _52509_/X _85808_/D sky130_fd_sc_hd__a21oi_4
X_83330_ _83753_/CLK _71915_/X _83330_/Q sky130_fd_sc_hd__dfxtp_4
X_61708_ _59664_/C _61708_/X sky130_fd_sc_hd__buf_2
X_80542_ _80542_/A _80527_/Y _80542_/X sky130_fd_sc_hd__or2_4
X_68264_ _67631_/X _67635_/X _68260_/X _68264_/Y sky130_fd_sc_hd__a21oi_4
X_65476_ _65428_/X _83078_/Q _65407_/X _65475_/X _65477_/B sky130_fd_sc_hd__a211o_4
X_53490_ _53468_/A _57523_/B _53490_/Y sky130_fd_sc_hd__nand2_4
X_62688_ _62686_/X _62652_/X _62687_/Y _62688_/Y sky130_fd_sc_hd__a21oi_4
X_67215_ _67241_/A _67215_/B _67215_/X sky130_fd_sc_hd__and2_4
X_52441_ _85822_/Q _52438_/X _52440_/Y _52441_/Y sky130_fd_sc_hd__o21ai_4
X_64427_ _64418_/Y _64426_/X _64386_/X _64427_/X sky130_fd_sc_hd__o21a_4
X_83261_ _81227_/CLK _83261_/D _72357_/A sky130_fd_sc_hd__dfxtp_4
X_61639_ _61342_/X _61639_/X sky130_fd_sc_hd__buf_2
X_80473_ _59182_/Y _66138_/Y _80472_/Y _80489_/A sky130_fd_sc_hd__o21a_4
X_68195_ _82055_/D _68180_/X _68194_/X _68195_/X sky130_fd_sc_hd__a21bo_4
X_85000_ _83335_/CLK _85000_/D _55248_/B sky130_fd_sc_hd__dfxtp_4
X_82212_ _81834_/CLK _82244_/Q _77254_/A sky130_fd_sc_hd__dfxtp_4
X_55160_ _82986_/Q _55157_/X _55172_/A _55159_/X _55160_/X sky130_fd_sc_hd__a211o_4
X_67146_ _87355_/Q _67121_/X _67122_/X _67145_/X _67146_/X sky130_fd_sc_hd__a211o_4
X_52372_ _52324_/A _52372_/X sky130_fd_sc_hd__buf_2
X_64358_ _64351_/Y _64357_/X _64328_/X _64358_/X sky130_fd_sc_hd__o21a_4
X_83192_ _83191_/CLK _72680_/X _70221_/C sky130_fd_sc_hd__dfxtp_4
X_54111_ _54123_/A _54123_/B _54111_/C _52942_/D _54111_/X sky130_fd_sc_hd__and4_4
X_51323_ _51321_/Y _51313_/X _51322_/X _86032_/D sky130_fd_sc_hd__a21oi_4
X_63309_ _79211_/B _79212_/A sky130_fd_sc_hd__inv_2
X_82143_ _82575_/CLK _78007_/Y _77471_/B sky130_fd_sc_hd__dfxtp_4
X_55091_ _55083_/A _55104_/B _55083_/C _47768_/A _55091_/X sky130_fd_sc_hd__and4_4
X_67077_ _88382_/Q _67074_/X _67075_/X _67076_/X _67078_/B sky130_fd_sc_hd__a211o_4
X_64289_ _64283_/X _64284_/X _64286_/X _64288_/Y _64267_/X _64289_/X
+ sky130_fd_sc_hd__o41a_4
X_54042_ _85517_/Q _54035_/X _54041_/Y _54042_/Y sky130_fd_sc_hd__o21ai_4
X_66028_ _65980_/X _66028_/B _66028_/X sky130_fd_sc_hd__and2_4
X_51254_ _86045_/Q _51233_/X _51253_/Y _51254_/Y sky130_fd_sc_hd__o21ai_4
X_86951_ _87141_/CLK _86951_/D _86951_/Q sky130_fd_sc_hd__dfxtp_4
X_82074_ _81970_/CLK _82074_/D _77961_/B sky130_fd_sc_hd__dfxtp_4
X_50205_ _51242_/A _50719_/B _50205_/X sky130_fd_sc_hd__and2_4
X_85902_ _86530_/CLK _85902_/D _85902_/Q sky130_fd_sc_hd__dfxtp_4
X_81025_ _84175_/CLK _84233_/Q _81025_/Q sky130_fd_sc_hd__dfxtp_4
X_58850_ _58845_/Y _58849_/Y _58761_/X _58850_/X sky130_fd_sc_hd__a21o_4
X_51185_ _51184_/X _52876_/B _51185_/Y sky130_fd_sc_hd__nand2_4
X_86882_ _86882_/CLK _45353_/Y _64535_/B sky130_fd_sc_hd__dfxtp_4
X_57801_ _57800_/X _57801_/X sky130_fd_sc_hd__buf_2
X_50136_ _50134_/Y _50117_/X _50135_/X _86257_/D sky130_fd_sc_hd__a21oi_4
X_85833_ _86154_/CLK _52386_/Y _65225_/B sky130_fd_sc_hd__dfxtp_4
X_58781_ _58696_/X _58779_/Y _58780_/Y _58728_/X _58701_/X _58781_/X
+ sky130_fd_sc_hd__o32a_4
X_55993_ _56102_/B _55993_/Y sky130_fd_sc_hd__inv_2
X_67979_ _68025_/A _88216_/Q _67979_/X sky130_fd_sc_hd__and2_4
X_57732_ _58805_/A _59286_/A sky130_fd_sc_hd__buf_2
X_69718_ _87815_/Q _69719_/B sky130_fd_sc_hd__inv_2
X_50067_ _48759_/A _50092_/A sky130_fd_sc_hd__buf_2
X_54944_ _53460_/A _47798_/A _54944_/Y sky130_fd_sc_hd__nand2_4
X_85764_ _85764_/CLK _52736_/Y _85764_/Q sky130_fd_sc_hd__dfxtp_4
X_70990_ _70990_/A _70942_/B _70990_/C _70990_/Y sky130_fd_sc_hd__nand3_4
X_82976_ _82973_/CLK _82784_/Q _46629_/A sky130_fd_sc_hd__dfxtp_4
X_87503_ _87260_/CLK _87503_/D _87503_/Q sky130_fd_sc_hd__dfxtp_4
X_84715_ _84903_/CLK _59503_/Y _64286_/C sky130_fd_sc_hd__dfxtp_4
X_57663_ _83758_/Q _57663_/Y sky130_fd_sc_hd__inv_2
X_81927_ _82124_/CLK _81927_/D _81927_/Q sky130_fd_sc_hd__dfxtp_4
X_69649_ _41996_/A _69607_/X _68555_/X _69648_/Y _69649_/X sky130_fd_sc_hd__a211o_4
X_54875_ _54872_/Y _54856_/X _54874_/X _54875_/Y sky130_fd_sc_hd__a21oi_4
X_85695_ _85697_/CLK _85695_/D _85695_/Q sky130_fd_sc_hd__dfxtp_4
X_59402_ _63139_/A _59403_/A sky130_fd_sc_hd__buf_2
X_56614_ _56602_/X _56614_/B _56696_/B _56614_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_7_73_0_CLK clkbuf_6_36_0_CLK/X clkbuf_7_73_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_87434_ _87484_/CLK _43411_/X _87434_/Q sky130_fd_sc_hd__dfxtp_4
X_41840_ _40637_/A _42465_/A sky130_fd_sc_hd__buf_2
X_53826_ _53824_/Y _53799_/X _53825_/Y _85561_/D sky130_fd_sc_hd__a21boi_4
X_72660_ _44290_/X _72688_/A sky130_fd_sc_hd__buf_2
X_84646_ _83218_/CLK _60248_/Y _79846_/A sky130_fd_sc_hd__dfxtp_4
X_57594_ _57591_/Y _57592_/X _57593_/X _57594_/Y sky130_fd_sc_hd__a21oi_4
X_81858_ _82211_/CLK _78049_/X _81858_/Q sky130_fd_sc_hd__dfxtp_4
X_59333_ _59331_/X _85414_/Q _59332_/X _59333_/Y sky130_fd_sc_hd__o21ai_4
X_71611_ _71215_/C _71614_/C sky130_fd_sc_hd__buf_2
X_56545_ _56545_/A _56177_/B _55738_/B _56545_/Y sky130_fd_sc_hd__nand3_4
X_80809_ _81134_/CLK _80809_/D _80809_/Q sky130_fd_sc_hd__dfxtp_4
X_41771_ _82886_/Q _48946_/A _41771_/X sky130_fd_sc_hd__or2_4
X_87365_ _86824_/CLK _43551_/Y _87365_/Q sky130_fd_sc_hd__dfxtp_4
X_53757_ _85574_/Q _53754_/X _53756_/Y _53757_/Y sky130_fd_sc_hd__o21ai_4
X_72591_ _79343_/B _72590_/X _61178_/Y _72562_/A _72591_/X sky130_fd_sc_hd__o22a_4
X_84577_ _84562_/CLK _84577_/D _60744_/C sky130_fd_sc_hd__dfxtp_4
X_50969_ _50963_/A _50963_/B _50963_/C _52661_/D _50969_/X sky130_fd_sc_hd__and4_4
X_81789_ _86753_/CLK _75939_/Y _48405_/A sky130_fd_sc_hd__dfxtp_4
X_43510_ _43495_/X _43503_/X _41773_/X _87384_/Q _43506_/X _43511_/A
+ sky130_fd_sc_hd__o32ai_4
X_74330_ _74338_/A _74338_/B _56098_/A _74330_/Y sky130_fd_sc_hd__nand3_4
X_86316_ _86637_/CLK _49831_/Y _58012_/B sky130_fd_sc_hd__dfxtp_4
X_52708_ _52708_/A _52708_/X sky130_fd_sc_hd__buf_2
X_40722_ _40722_/A _40760_/B _40722_/X sky130_fd_sc_hd__or2_4
X_59264_ _59199_/X _85740_/Q _59263_/X _59264_/X sky130_fd_sc_hd__o21a_4
X_71542_ _70676_/A _71546_/B _71546_/C _71542_/Y sky130_fd_sc_hd__nor3_4
X_83528_ _83526_/CLK _83528_/D _83528_/Q sky130_fd_sc_hd__dfxtp_4
X_44490_ _44489_/Y _44490_/Y sky130_fd_sc_hd__inv_2
X_56476_ _56020_/X _56468_/X _56475_/Y _56476_/Y sky130_fd_sc_hd__o21ai_4
X_87296_ _87813_/CLK _43723_/Y _87296_/Q sky130_fd_sc_hd__dfxtp_4
X_53688_ _53755_/A _53713_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_88_0_CLK clkbuf_7_89_0_CLK/A clkbuf_7_88_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_58215_ _58171_/X _83370_/Q _58214_/Y _84906_/D sky130_fd_sc_hd__o21a_4
XPHY_410 sky130_fd_sc_hd__decap_3
X_43441_ _41586_/X _43431_/X _87419_/Q _43432_/X _87419_/D sky130_fd_sc_hd__a2bb2o_4
X_55427_ _57186_/B _55426_/X _55427_/Y sky130_fd_sc_hd__nand2_4
X_86247_ _86154_/CLK _50184_/Y _65285_/B sky130_fd_sc_hd__dfxtp_4
X_74261_ _74259_/X _74248_/X _74250_/X _74261_/Y sky130_fd_sc_hd__nand3_4
X_40653_ _40650_/X _40651_/X _68645_/B _40652_/X _40653_/X sky130_fd_sc_hd__a2bb2o_4
XPHY_421 sky130_fd_sc_hd__decap_3
X_52639_ _52643_/A _52654_/B _52643_/C _46728_/X _52639_/X sky130_fd_sc_hd__and4_4
X_59195_ _59115_/X _59192_/Y _59194_/Y _59133_/X _59119_/X _59195_/X
+ sky130_fd_sc_hd__o32a_4
X_71473_ _70880_/B _71479_/B _70778_/A _71476_/D _71473_/X sky130_fd_sc_hd__and4_4
X_83459_ _83495_/CLK _83459_/D _83459_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_432 sky130_fd_sc_hd__decap_3
XPHY_443 sky130_fd_sc_hd__decap_3
X_76000_ _81708_/D _81420_/Q _76000_/Y sky130_fd_sc_hd__nand2_4
XPHY_454 sky130_fd_sc_hd__decap_3
X_73212_ _73210_/X _85584_/Q _73092_/X _73211_/X _73212_/X sky130_fd_sc_hd__a211o_4
X_46160_ _46087_/A _46121_/A _46162_/C sky130_fd_sc_hd__nor2_4
X_70424_ _71162_/B _70423_/X _70495_/A _70609_/A _70424_/X sky130_fd_sc_hd__and4_4
X_58146_ _61323_/A _58147_/A sky130_fd_sc_hd__buf_2
XPHY_465 sky130_fd_sc_hd__decap_3
X_43372_ _43302_/A _43372_/X sky130_fd_sc_hd__buf_2
X_55358_ _55369_/A _55369_/B _56689_/A sky130_fd_sc_hd__nand2_4
X_74192_ _74232_/A _66296_/B _74192_/X sky130_fd_sc_hd__and2_4
X_86178_ _83307_/CLK _50557_/Y _86178_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_476 sky130_fd_sc_hd__decap_3
X_40584_ _40878_/A _40585_/A sky130_fd_sc_hd__buf_2
XPHY_487 sky130_fd_sc_hd__decap_3
X_45111_ _45052_/X _61489_/B _45070_/X _45111_/Y sky130_fd_sc_hd__o21ai_4
XPHY_498 sky130_fd_sc_hd__decap_3
X_54309_ _54314_/A _54309_/B _54309_/Y sky130_fd_sc_hd__nand2_4
X_42323_ _41636_/X _42303_/X _87922_/Q _42305_/X _87922_/D sky130_fd_sc_hd__a2bb2o_4
X_73143_ _73141_/X _73128_/X _73131_/Y _73143_/Y sky130_fd_sc_hd__nand3_4
X_85129_ _85031_/CLK _85129_/D _85129_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_11_0_CLK clkbuf_6_5_0_CLK/X clkbuf_8_23_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_70355_ _70355_/A _71003_/A sky130_fd_sc_hd__buf_2
X_46091_ _46111_/A _46091_/Y sky130_fd_sc_hd__inv_2
X_58077_ _58074_/Y _58076_/Y _58035_/X _58077_/X sky130_fd_sc_hd__a21o_4
X_55289_ _55674_/B _55286_/Y _55284_/X _55289_/X sky130_fd_sc_hd__a21bo_4
Xclkbuf_8_151_0_CLK clkbuf_7_75_0_CLK/X clkbuf_9_303_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_45042_ _85208_/Q _45027_/X _45041_/X _45042_/Y sky130_fd_sc_hd__o21ai_4
X_57028_ _57025_/X _46178_/X _57027_/Y _57028_/Y sky130_fd_sc_hd__a21oi_4
X_42254_ _42254_/A _42254_/Y sky130_fd_sc_hd__inv_2
X_73074_ _73058_/X _73075_/C _73073_/X _73074_/X sky130_fd_sc_hd__a21o_4
X_77951_ _82170_/Q _77951_/B _82138_/D sky130_fd_sc_hd__xor2_4
X_70286_ _70269_/X _74756_/B _70285_/X _70286_/X sky130_fd_sc_hd__a21o_4
X_41205_ _40999_/A _41205_/X sky130_fd_sc_hd__buf_2
X_72025_ _72025_/A _72025_/B _72025_/Y sky130_fd_sc_hd__nand2_4
X_76902_ _76904_/A _76902_/B _76902_/Y sky130_fd_sc_hd__nand2_4
X_49850_ _49794_/X _49862_/C sky130_fd_sc_hd__buf_2
X_42185_ _41264_/X _42183_/X _87992_/Q _42184_/X _42185_/X sky130_fd_sc_hd__a2bb2o_4
X_77882_ _82067_/Q _77884_/A sky130_fd_sc_hd__inv_2
X_48801_ _48801_/A _48801_/B _48801_/X sky130_fd_sc_hd__and2_4
Xclkbuf_7_26_0_CLK clkbuf_7_26_0_CLK/A clkbuf_8_53_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_79621_ _79597_/A _79611_/Y _79621_/Y sky130_fd_sc_hd__nor2_4
X_41136_ _41072_/X _41136_/X sky130_fd_sc_hd__buf_2
X_76833_ _76811_/Y _81364_/D sky130_fd_sc_hd__inv_2
X_49781_ _49769_/X _52995_/B _49781_/Y sky130_fd_sc_hd__nand2_4
X_46993_ _83049_/Q _53309_/B sky130_fd_sc_hd__inv_2
X_58979_ _58978_/Y _58973_/B _58979_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_166_0_CLK clkbuf_7_83_0_CLK/X clkbuf_8_166_0_CLK/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_161_0_CLK clkbuf_9_80_0_CLK/X _85003_/CLK sky130_fd_sc_hd__clkbuf_1
X_48732_ _48737_/A _48401_/B _48732_/Y sky130_fd_sc_hd__nand2_4
X_79552_ _79552_/A _79553_/A _79555_/B sky130_fd_sc_hd__nand2_4
X_45944_ _64961_/A _60150_/A sky130_fd_sc_hd__buf_2
X_41067_ _41064_/X _41065_/X _88284_/Q _41066_/X _88284_/D sky130_fd_sc_hd__a2bb2o_4
X_76764_ _81582_/Q _76764_/B _81550_/D sky130_fd_sc_hd__xor2_4
X_61990_ _61988_/Y _61959_/X _61989_/Y _61990_/Y sky130_fd_sc_hd__a21oi_4
X_73976_ _73954_/A _66159_/B _73976_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_791_0_CLK clkbuf_9_395_0_CLK/X _81019_/CLK sky130_fd_sc_hd__clkbuf_1
X_78503_ _78503_/A _82672_/D _78503_/Y sky130_fd_sc_hd__nand2_4
X_75715_ _75715_/A _75714_/Y _75723_/A sky130_fd_sc_hd__xor2_4
X_60941_ _60940_/Y _61024_/B sky130_fd_sc_hd__inv_2
X_72927_ _88333_/Q _72803_/X _72776_/X _72927_/Y sky130_fd_sc_hd__o21ai_4
X_48663_ _81766_/Q _48664_/A sky130_fd_sc_hd__inv_2
X_79483_ _79449_/A _79448_/Y _79460_/X _79481_/A _79480_/Y _79483_/X
+ sky130_fd_sc_hd__a2111o_4
X_45875_ _45875_/A _45876_/A sky130_fd_sc_hd__inv_2
X_76695_ _76695_/A _81447_/D _81543_/D sky130_fd_sc_hd__xor2_4
Xclkbuf_9_282_0_CLK clkbuf_9_283_0_CLK/A clkbuf_9_282_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_47614_ _47661_/A _47614_/X sky130_fd_sc_hd__buf_2
X_78434_ _78434_/A _78434_/B _78439_/C sky130_fd_sc_hd__nand2_4
X_44826_ _41680_/Y _44817_/X _67559_/B _44818_/X _44826_/X sky130_fd_sc_hd__a2bb2o_4
X_63660_ _61627_/B _63609_/X _63657_/X _63659_/X _63660_/X sky130_fd_sc_hd__a211o_4
X_75646_ _75641_/Y _75609_/Y _75645_/Y _75660_/A sky130_fd_sc_hd__o21ai_4
X_48594_ _49212_/A _48820_/B _48594_/Y sky130_fd_sc_hd__nand2_4
X_60872_ _60871_/Y _61003_/A sky130_fd_sc_hd__buf_2
X_72858_ _72857_/X _72858_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_176_0_CLK clkbuf_9_88_0_CLK/X _83316_/CLK sky130_fd_sc_hd__clkbuf_1
X_62611_ _61676_/A _62631_/B _62259_/X _62631_/D _62614_/B sky130_fd_sc_hd__nand4_4
X_47545_ _47553_/A _53109_/B _47545_/Y sky130_fd_sc_hd__nand2_4
X_71809_ _71805_/X _83368_/Q _71808_/X _83368_/D sky130_fd_sc_hd__a21o_4
X_78365_ _78365_/A _78365_/Y sky130_fd_sc_hd__inv_2
X_44757_ _41305_/Y _44754_/X _86971_/Q _44755_/X _44757_/X sky130_fd_sc_hd__a2bb2o_4
X_63591_ _63468_/A _63615_/B sky130_fd_sc_hd__buf_2
X_75577_ _80819_/Q _75577_/Y sky130_fd_sc_hd__inv_2
X_41969_ _88088_/Q _41969_/Y sky130_fd_sc_hd__inv_2
X_72789_ _48367_/Y _72789_/B _72789_/X sky130_fd_sc_hd__xor2_4
X_65330_ _65673_/A _65408_/A sky130_fd_sc_hd__buf_2
X_77316_ _77316_/A _77316_/B _77317_/A sky130_fd_sc_hd__and2_4
X_62542_ _62539_/Y _62540_/X _62541_/Y _84403_/D sky130_fd_sc_hd__a21oi_4
X_43708_ _43707_/X _87301_/D sky130_fd_sc_hd__inv_2
X_74528_ _52813_/B _74517_/X _74527_/Y _74528_/Y sky130_fd_sc_hd__o21ai_4
X_47476_ _47471_/Y _47462_/X _47475_/X _86631_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_297_0_CLK clkbuf_9_296_0_CLK/A clkbuf_9_297_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_78296_ _78296_/A _78296_/B _78296_/Y sky130_fd_sc_hd__nand2_4
X_44688_ _44688_/A _44688_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_104_0_CLK clkbuf_7_52_0_CLK/X clkbuf_8_104_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_49215_ _49215_/A _49220_/A sky130_fd_sc_hd__buf_2
X_46427_ _46427_/A _50802_/A sky130_fd_sc_hd__buf_2
X_65261_ _65211_/X _85512_/Q _65212_/X _65260_/X _65261_/X sky130_fd_sc_hd__a211o_4
X_77247_ _77246_/X _82179_/D sky130_fd_sc_hd__buf_2
X_43639_ _40673_/X _43624_/X _73921_/A _43625_/X _87332_/D sky130_fd_sc_hd__a2bb2o_4
X_62473_ _62203_/Y _62533_/A sky130_fd_sc_hd__buf_2
X_74459_ _48578_/A _74478_/B _74478_/C _74459_/X sky130_fd_sc_hd__and3_4
X_67000_ _87361_/Q _66997_/X _66998_/X _66999_/X _67000_/X sky130_fd_sc_hd__a211o_4
X_64212_ _63355_/A _61226_/X _64211_/Y _64212_/Y sky130_fd_sc_hd__o21ai_4
X_49146_ _65289_/B _49104_/X _49145_/Y _49146_/Y sky130_fd_sc_hd__o21ai_4
X_61424_ _61417_/Y _61420_/Y _61403_/X _61421_/Y _61423_/Y _61424_/X
+ sky130_fd_sc_hd__a41o_4
X_46358_ _86744_/Q _46279_/X _46357_/Y _46358_/Y sky130_fd_sc_hd__o21ai_4
X_65192_ _65188_/X _65192_/B _65191_/X _65192_/Y sky130_fd_sc_hd__nand3_4
X_77178_ _82106_/Q _77178_/B _77178_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_9_220_0_CLK clkbuf_9_220_0_CLK/A clkbuf_9_220_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_45309_ _45277_/X _61636_/B _45294_/X _45309_/Y sky130_fd_sc_hd__o21ai_4
X_76129_ _76122_/X _76129_/B _76130_/B sky130_fd_sc_hd__xor2_4
X_64143_ _64026_/A _64190_/B sky130_fd_sc_hd__buf_2
X_49077_ _49077_/A _49029_/B _49077_/Y sky130_fd_sc_hd__nor2_4
X_61355_ _61355_/A _61377_/A sky130_fd_sc_hd__buf_2
X_46289_ _46284_/Y _46258_/X _46288_/Y _46289_/Y sky130_fd_sc_hd__a21boi_4
Xclkbuf_8_119_0_CLK clkbuf_7_59_0_CLK/X clkbuf_9_239_0_CLK/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_114_0_CLK clkbuf_9_57_0_CLK/X _84424_/CLK sky130_fd_sc_hd__clkbuf_1
X_48028_ _47981_/X _48028_/B _48028_/X sky130_fd_sc_hd__and2_4
X_60306_ _60263_/A _60367_/C _60241_/A _60306_/Y sky130_fd_sc_hd__o21ai_4
X_68951_ _68946_/X _68950_/X _68878_/X _68951_/Y sky130_fd_sc_hd__a21oi_4
X_64074_ _64074_/A _64074_/B _80040_/B _64074_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_10_744_0_CLK clkbuf_9_372_0_CLK/X _87995_/CLK sky130_fd_sc_hd__clkbuf_1
X_61286_ _61286_/A _61286_/B _61287_/D sky130_fd_sc_hd__nor2_4
X_67902_ _87963_/Q _67831_/X _67879_/X _67901_/X _67902_/X sky130_fd_sc_hd__a211o_4
X_63025_ _58412_/A _63010_/X _60523_/X _59456_/Y _60412_/X _63025_/Y
+ sky130_fd_sc_hd__o32ai_4
X_60237_ _60254_/B _60255_/B _60350_/A sky130_fd_sc_hd__nor2_4
X_68882_ _60111_/X _68882_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_235_0_CLK clkbuf_9_235_0_CLK/A clkbuf_9_235_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_79819_ _79819_/A _79818_/Y _79829_/B sky130_fd_sc_hd__xor2_4
X_67833_ _87902_/Q _67831_/X _67761_/X _67832_/X _67833_/X sky130_fd_sc_hd__a211o_4
X_60168_ _60168_/A _60239_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_129_0_CLK clkbuf_9_64_0_CLK/X _83819_/CLK sky130_fd_sc_hd__clkbuf_1
X_49979_ _49995_/A _49973_/B _49973_/C _53191_/D _49979_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_759_0_CLK clkbuf_9_379_0_CLK/X _88087_/CLK sky130_fd_sc_hd__clkbuf_1
X_82830_ _82425_/CLK _82830_/D _82830_/Q sky130_fd_sc_hd__dfxtp_4
X_67764_ _67739_/X _87201_/Q _67764_/X sky130_fd_sc_hd__and2_4
X_64976_ _58785_/A _86035_/Q _64976_/X sky130_fd_sc_hd__and2_4
X_52990_ _52987_/Y _52975_/X _52989_/X _52990_/Y sky130_fd_sc_hd__a21oi_4
X_60099_ _60042_/D _59951_/B _60087_/Y _60099_/X sky130_fd_sc_hd__and3_4
X_69503_ _81383_/D _69439_/X _69502_/X _83919_/D sky130_fd_sc_hd__a21bo_4
X_66715_ _69457_/A _66715_/X sky130_fd_sc_hd__buf_2
X_51941_ _51941_/A _50234_/B _51941_/Y sky130_fd_sc_hd__nand2_4
X_63927_ _63922_/X _63890_/X _63923_/Y _63924_/Y _63926_/X _63927_/X
+ sky130_fd_sc_hd__a41o_4
X_82761_ _82774_/CLK _82761_/D _82953_/D sky130_fd_sc_hd__dfxtp_4
X_67695_ _67692_/X _67694_/X _67619_/X _67698_/A sky130_fd_sc_hd__a21o_4
X_84500_ _84501_/CLK _61242_/Y _75902_/A sky130_fd_sc_hd__dfxtp_4
X_81712_ _81749_/CLK _81712_/D _81712_/Q sky130_fd_sc_hd__dfxtp_4
X_69434_ _69429_/X _69432_/X _69433_/X _69434_/Y sky130_fd_sc_hd__a21oi_4
X_54660_ _54649_/X _47297_/Y _54660_/Y sky130_fd_sc_hd__nand2_4
X_66646_ _66641_/X _66645_/X _66547_/X _66646_/X sky130_fd_sc_hd__a21o_4
X_85480_ _84926_/CLK _54233_/Y _85480_/Q sky130_fd_sc_hd__dfxtp_4
X_51872_ _48808_/A _51900_/A sky130_fd_sc_hd__buf_2
X_63858_ _58248_/A _63858_/B _63858_/C _63793_/D _63859_/D sky130_fd_sc_hd__nand4_4
X_82692_ _82692_/CLK _78831_/X _82692_/Q sky130_fd_sc_hd__dfxtp_4
X_53611_ _53723_/A _53611_/X sky130_fd_sc_hd__buf_2
X_84431_ _84430_/CLK _84431_/D _78054_/B sky130_fd_sc_hd__dfxtp_4
X_50823_ _86126_/Q _50820_/X _50822_/Y _50823_/Y sky130_fd_sc_hd__o21ai_4
X_62809_ _62819_/A _84828_/Q _62819_/C _62782_/X _62809_/X sky130_fd_sc_hd__and4_4
X_81643_ _81660_/CLK _76874_/A _81643_/Q sky130_fd_sc_hd__dfxtp_4
X_69365_ _69329_/X _68777_/Y _69325_/X _69364_/Y _69365_/X sky130_fd_sc_hd__a211o_4
X_54591_ _54589_/X _54585_/B _54591_/C _47180_/A _54591_/X sky130_fd_sc_hd__and4_4
X_66577_ _69223_/A _66577_/B _66577_/X sky130_fd_sc_hd__and2_4
X_63789_ _63396_/B _63820_/B _63753_/C _63820_/D _63789_/Y sky130_fd_sc_hd__nand4_4
X_56330_ _56332_/A _56335_/B _85233_/Q _56330_/Y sky130_fd_sc_hd__nand3_4
X_68316_ _68301_/X _67934_/Y _68308_/X _68315_/Y _68316_/X sky130_fd_sc_hd__a211o_4
X_87150_ _87150_/CLK _44357_/X _87150_/Q sky130_fd_sc_hd__dfxtp_4
X_53542_ _53548_/A _48014_/Y _53542_/Y sky130_fd_sc_hd__nand2_4
X_65528_ _65516_/X _64775_/Y _65527_/Y _65528_/Y sky130_fd_sc_hd__o21ai_4
X_84362_ _83216_/CLK _84362_/D _62995_/C sky130_fd_sc_hd__dfxtp_4
X_50754_ _86140_/Q _50727_/X _50753_/Y _50754_/Y sky130_fd_sc_hd__o21ai_4
X_81574_ _81412_/CLK _84174_/Q _76689_/A sky130_fd_sc_hd__dfxtp_4
X_69296_ _68656_/X _68659_/X _69295_/X _69296_/Y sky130_fd_sc_hd__a21oi_4
X_86101_ _86104_/CLK _86101_/D _86101_/Q sky130_fd_sc_hd__dfxtp_4
X_83313_ _83313_/CLK _71961_/Y _83313_/Q sky130_fd_sc_hd__dfxtp_4
X_56261_ _56263_/A _56263_/B _85255_/Q _56261_/Y sky130_fd_sc_hd__nand3_4
X_80525_ _84768_/Q _84160_/Q _80525_/X sky130_fd_sc_hd__xor2_4
X_68247_ _68168_/A _68247_/X sky130_fd_sc_hd__buf_2
X_87081_ _87086_/CLK _87081_/D _87081_/Q sky130_fd_sc_hd__dfxtp_4
X_53473_ _50724_/A _53474_/B sky130_fd_sc_hd__buf_2
X_65459_ _65408_/A _72817_/B _65459_/X sky130_fd_sc_hd__and2_4
X_84293_ _84293_/CLK _84293_/D _80206_/B sky130_fd_sc_hd__dfxtp_4
X_50685_ _50683_/Y _50644_/X _50684_/Y _50685_/Y sky130_fd_sc_hd__a21boi_4
X_58000_ _57947_/X _85709_/Q _57948_/X _58000_/X sky130_fd_sc_hd__o21a_4
X_55212_ _85090_/Q _55152_/A _55133_/X _55211_/X _55212_/X sky130_fd_sc_hd__a211o_4
X_86032_ _86030_/CLK _86032_/D _65051_/B sky130_fd_sc_hd__dfxtp_4
X_52424_ _52448_/A _51235_/B _52424_/Y sky130_fd_sc_hd__nand2_4
X_83244_ _84555_/CLK _72497_/X _62055_/B sky130_fd_sc_hd__dfxtp_4
X_80456_ _80456_/A _80456_/B _80456_/Y sky130_fd_sc_hd__xnor2_4
X_56192_ _56280_/A _56192_/B _56192_/C _56192_/Y sky130_fd_sc_hd__nand3_4
X_68178_ _68144_/X _67102_/Y _68168_/X _68177_/Y _68178_/X sky130_fd_sc_hd__a211o_4
X_55143_ _55278_/A _55145_/A sky130_fd_sc_hd__buf_2
X_67129_ _87112_/Q _67074_/X _67075_/X _67128_/X _67129_/X sky130_fd_sc_hd__a211o_4
X_52355_ _52355_/A _52310_/B _52291_/C _52355_/X sky130_fd_sc_hd__and3_4
X_83175_ _83161_/CLK _83175_/D _83175_/Q sky130_fd_sc_hd__dfxtp_4
X_80387_ _80404_/B _80386_/Y _80387_/X sky130_fd_sc_hd__xor2_4
X_51306_ _51282_/A _51306_/X sky130_fd_sc_hd__buf_2
X_70140_ _83518_/Q _83166_/Q _83515_/Q _83163_/Q _70144_/A sky130_fd_sc_hd__a22oi_4
X_82126_ _83906_/CLK _77843_/X _82082_/D sky130_fd_sc_hd__dfxtp_4
X_55074_ _55093_/A _54907_/B _55074_/Y sky130_fd_sc_hd__nand2_4
X_59951_ _60042_/D _59951_/B _59951_/C _59951_/D _59951_/Y sky130_fd_sc_hd__nand4_4
X_52286_ _52284_/Y _52262_/X _52285_/X _85853_/D sky130_fd_sc_hd__a21oi_4
X_87983_ _87471_/CLK _87983_/D _87983_/Q sky130_fd_sc_hd__dfxtp_4
X_58902_ _58835_/X _85447_/Q _58901_/X _58902_/Y sky130_fd_sc_hd__o21ai_4
X_54025_ _85520_/Q _53940_/X _54024_/Y _54025_/Y sky130_fd_sc_hd__o21ai_4
X_51237_ _51263_/A _51237_/X sky130_fd_sc_hd__buf_2
X_86934_ _86934_/CLK _44826_/X _67559_/B sky130_fd_sc_hd__dfxtp_4
X_82057_ _84014_/CLK _82057_/D _77787_/A sky130_fd_sc_hd__dfxtp_4
X_70071_ _68961_/X _68963_/X _70044_/X _70071_/Y sky130_fd_sc_hd__a21oi_4
X_59882_ _59741_/A _59544_/B _59581_/C _59882_/X sky130_fd_sc_hd__and3_4
X_81008_ _84228_/CLK _84216_/Q _81008_/Q sky130_fd_sc_hd__dfxtp_4
X_58833_ _58828_/X _58830_/Y _58831_/Y _58728_/X _58832_/X _58833_/X
+ sky130_fd_sc_hd__o32a_4
X_51168_ _86061_/Q _51156_/X _51167_/Y _51168_/Y sky130_fd_sc_hd__o21ai_4
X_86865_ _84408_/CLK _86865_/D _63168_/B sky130_fd_sc_hd__dfxtp_4
X_50119_ _50116_/Y _50117_/X _50118_/X _86261_/D sky130_fd_sc_hd__a21oi_4
X_73830_ _73829_/X _73830_/B _73830_/X sky130_fd_sc_hd__and2_4
X_85816_ _85529_/CLK _52469_/Y _85816_/Q sky130_fd_sc_hd__dfxtp_4
X_58764_ _86706_/Q _58764_/B _58764_/Y sky130_fd_sc_hd__nor2_4
X_43990_ _86842_/Q _43990_/Y sky130_fd_sc_hd__inv_2
X_51099_ _51084_/A _51115_/B _51110_/C _52790_/D _51099_/X sky130_fd_sc_hd__and4_4
X_55976_ _55695_/A _55976_/B _55976_/X sky130_fd_sc_hd__and2_4
X_86796_ _86796_/CLK _86796_/D _66819_/B sky130_fd_sc_hd__dfxtp_4
X_57715_ _64850_/A _57716_/A sky130_fd_sc_hd__buf_2
X_42941_ _42940_/Y _42941_/Y sky130_fd_sc_hd__inv_2
X_54927_ _54927_/A _54942_/B sky130_fd_sc_hd__buf_2
X_85747_ _85748_/CLK _52832_/Y _85747_/Q sky130_fd_sc_hd__dfxtp_4
X_73761_ _73758_/X _73760_/X _73738_/X _73764_/A sky130_fd_sc_hd__a21o_4
X_70973_ _49265_/B _70961_/X _70972_/Y _83645_/D sky130_fd_sc_hd__o21ai_4
X_58695_ _84807_/Q _58599_/X _58689_/X _58694_/X _58695_/Y sky130_fd_sc_hd__a2bb2oi_4
X_82959_ _82769_/CLK _82767_/Q _46790_/A sky130_fd_sc_hd__dfxtp_4
X_75500_ _75477_/A _75477_/B _75475_/Y _75500_/X sky130_fd_sc_hd__o21a_4
X_72712_ _72710_/A _44907_/A _72712_/C _55209_/X _72712_/X sky130_fd_sc_hd__and4_4
X_45660_ _56989_/B _45793_/B _45660_/Y sky130_fd_sc_hd__nor2_4
X_57646_ _71972_/A _48153_/A _57646_/Y sky130_fd_sc_hd__nand2_4
X_76480_ _76478_/X _76513_/C _76481_/A sky130_fd_sc_hd__and2_4
X_42872_ _41586_/X _42866_/X _87675_/Q _42867_/X _87675_/D sky130_fd_sc_hd__a2bb2o_4
X_54858_ _54855_/Y _54856_/X _54857_/X _54858_/Y sky130_fd_sc_hd__a21oi_4
X_73692_ _73692_/A _73692_/B _73692_/X sky130_fd_sc_hd__xor2_4
X_85678_ _84802_/CLK _85678_/D _85678_/Q sky130_fd_sc_hd__dfxtp_4
X_44611_ _40964_/A _44602_/X _87034_/Q _44603_/X _87034_/D sky130_fd_sc_hd__a2bb2o_4
X_75431_ _75427_/X _75432_/C _75430_/Y _75431_/X sky130_fd_sc_hd__a21o_4
X_87417_ _87417_/CLK _43444_/Y _87417_/Q sky130_fd_sc_hd__dfxtp_4
X_53809_ _85564_/Q _53784_/X _53808_/Y _53809_/Y sky130_fd_sc_hd__o21ai_4
X_41823_ _41822_/Y _88135_/D sky130_fd_sc_hd__inv_2
X_72643_ _72633_/X _72643_/B _72643_/C _72643_/Y sky130_fd_sc_hd__nand3_4
X_84629_ _84590_/CLK _60338_/X _79671_/A sky130_fd_sc_hd__dfxtp_4
X_45591_ _45668_/A _45591_/X sky130_fd_sc_hd__buf_2
X_57577_ _57575_/Y _57543_/X _57576_/Y _57577_/Y sky130_fd_sc_hd__a21boi_4
X_88397_ _86834_/CLK _88397_/D _88397_/Q sky130_fd_sc_hd__dfxtp_4
X_54789_ _54787_/Y _54774_/X _54788_/X _54789_/Y sky130_fd_sc_hd__a21oi_4
X_47330_ _47330_/A _47349_/B _47370_/C _52989_/D _47330_/X sky130_fd_sc_hd__and4_4
X_59316_ _59256_/A _86343_/Q _59316_/Y sky130_fd_sc_hd__nor2_4
X_78150_ _78141_/Y _78148_/Y _78149_/Y _78150_/X sky130_fd_sc_hd__o21a_4
X_44542_ _44542_/A _44542_/Y sky130_fd_sc_hd__inv_2
X_56528_ _56528_/A _56528_/X sky130_fd_sc_hd__buf_2
X_75362_ _75362_/A _75362_/B _75362_/X sky130_fd_sc_hd__xor2_4
X_41754_ _41825_/A _41754_/X sky130_fd_sc_hd__buf_2
X_87348_ _87348_/CLK _87348_/D _87348_/Q sky130_fd_sc_hd__dfxtp_4
X_72574_ _72517_/B _72546_/Y _72572_/X _72537_/Y _72573_/Y _72574_/Y
+ sky130_fd_sc_hd__a41oi_4
X_77101_ _77097_/Y _77100_/X _77113_/A sky130_fd_sc_hd__nand2_4
X_74313_ _83102_/Q _74301_/X _74312_/Y _83102_/D sky130_fd_sc_hd__a21bo_4
X_40705_ _40705_/A _40760_/B _40705_/X sky130_fd_sc_hd__or2_4
X_47261_ _47241_/X _52944_/B _47261_/Y sky130_fd_sc_hd__nand2_4
X_59247_ _59135_/X _85645_/Q _59196_/X _59247_/X sky130_fd_sc_hd__o21a_4
X_71525_ _71525_/A _70727_/A _71525_/Y sky130_fd_sc_hd__nand2_4
X_78081_ _78083_/A _78083_/B _78082_/B sky130_fd_sc_hd__xor2_4
X_56459_ _56459_/A _56458_/Y _56459_/Y sky130_fd_sc_hd__nand2_4
X_44473_ _41178_/Y _44464_/X _87090_/Q _44466_/X _44473_/X sky130_fd_sc_hd__a2bb2o_4
X_75293_ _75291_/X _75292_/Y _75293_/X sky130_fd_sc_hd__and2_4
X_87279_ _88056_/CLK _43762_/Y _87279_/Q sky130_fd_sc_hd__dfxtp_4
X_41685_ _41681_/X _41682_/X _67563_/B _41684_/X _88170_/D sky130_fd_sc_hd__a2bb2o_4
X_49000_ _48994_/Y _48985_/X _48999_/X _49000_/Y sky130_fd_sc_hd__a21oi_4
X_46212_ _46212_/A _59325_/A sky130_fd_sc_hd__buf_2
XPHY_240 sky130_fd_sc_hd__decap_3
X_77032_ _77034_/C _77031_/Y _77033_/B sky130_fd_sc_hd__xnor2_4
X_43424_ _43424_/A _87428_/D sky130_fd_sc_hd__inv_2
X_74244_ _87829_/Q _74244_/B _74244_/Y sky130_fd_sc_hd__nor2_4
XPHY_251 sky130_fd_sc_hd__decap_3
X_40636_ _40636_/A _40637_/A sky130_fd_sc_hd__buf_2
X_47192_ _47004_/A _47192_/X sky130_fd_sc_hd__buf_2
X_59178_ _59073_/X _85747_/Q _59124_/X _59178_/X sky130_fd_sc_hd__o21a_4
X_71456_ _71411_/A _71446_/X _71458_/C _71456_/Y sky130_fd_sc_hd__nor3_4
XPHY_262 sky130_fd_sc_hd__decap_3
Xclkbuf_10_1001_0_CLK clkbuf_9_500_0_CLK/X _85599_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_273 sky130_fd_sc_hd__decap_3
XPHY_284 sky130_fd_sc_hd__decap_3
X_46143_ _46143_/A _46143_/B _46121_/Y _46143_/D _46143_/Y sky130_fd_sc_hd__nand4_4
X_70407_ _70942_/A _74533_/A _70407_/C _70407_/Y sky130_fd_sc_hd__nand3_4
X_58129_ _58122_/Y _58128_/Y _58003_/X _58129_/X sky130_fd_sc_hd__a21o_4
XPHY_295 sky130_fd_sc_hd__decap_3
X_43355_ _43355_/A _87464_/D sky130_fd_sc_hd__inv_2
X_74175_ _74106_/X _85607_/Q _74107_/X _74174_/X _74175_/X sky130_fd_sc_hd__a211o_4
X_40567_ _40567_/A _40568_/A sky130_fd_sc_hd__buf_2
X_71387_ _71373_/X _83517_/Q _71386_/Y _83517_/D sky130_fd_sc_hd__a21o_4
X_42306_ _41592_/X _42303_/X _87930_/Q _42305_/X _87930_/D sky130_fd_sc_hd__a2bb2o_4
X_61140_ _64243_/A _61140_/X sky130_fd_sc_hd__buf_2
X_73126_ _73126_/A _73198_/B _73126_/Y sky130_fd_sc_hd__nor2_4
X_70338_ _70338_/A _70333_/B _83088_/Q _70332_/X _70338_/X sky130_fd_sc_hd__and4_4
X_46074_ _46067_/X _46054_/X _41595_/X _86780_/Q _46068_/X _46075_/A
+ sky130_fd_sc_hd__o32ai_4
X_43286_ _43178_/X _43287_/A sky130_fd_sc_hd__buf_2
X_78983_ _82646_/Q _78998_/A sky130_fd_sc_hd__inv_2
X_40498_ _40497_/X _40410_/X _88382_/Q _40411_/X _40498_/X sky130_fd_sc_hd__a2bb2o_4
X_49902_ _72160_/B _49880_/X _49901_/Y _49902_/Y sky130_fd_sc_hd__o21ai_4
X_45025_ _85241_/Q _44979_/X _45012_/X _45025_/X sky130_fd_sc_hd__o21a_4
X_42237_ _41397_/X _42222_/X _87966_/Q _42224_/X _42237_/X sky130_fd_sc_hd__a2bb2o_4
X_77934_ _82168_/Q _77934_/B _82136_/D sky130_fd_sc_hd__xor2_4
X_61071_ _61071_/A _59602_/A _61071_/C _59532_/A _61071_/X sky130_fd_sc_hd__and4_4
X_73057_ _43141_/Y _72830_/X _73055_/X _73056_/Y _73057_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_1016_0_CLK clkbuf_9_508_0_CLK/X _86191_/CLK sky130_fd_sc_hd__clkbuf_1
X_70269_ _70238_/A _70269_/X sky130_fd_sc_hd__buf_2
X_60022_ _60009_/Y _60015_/Y _60019_/Y _59998_/B _60021_/Y _84674_/D
+ sky130_fd_sc_hd__a41oi_4
X_72008_ _83303_/Q _71985_/X _72007_/Y _72008_/Y sky130_fd_sc_hd__o21ai_4
X_49833_ _58026_/B _49825_/X _49832_/Y _49833_/Y sky130_fd_sc_hd__o21ai_4
X_42168_ _42167_/Y _88000_/D sky130_fd_sc_hd__inv_2
X_77865_ _77863_/Y _77864_/Y _77869_/A sky130_fd_sc_hd__xor2_4
X_79604_ _79601_/X _79602_/X _79603_/Y _79609_/A sky130_fd_sc_hd__nand3_4
X_41119_ _41119_/A _41102_/B _41119_/X sky130_fd_sc_hd__or2_4
X_64830_ _64883_/A _86265_/Q _64830_/X sky130_fd_sc_hd__and2_4
X_76816_ _76805_/A _76804_/Y _76815_/X _76816_/Y sky130_fd_sc_hd__a21oi_4
X_49764_ _57870_/B _49742_/X _49763_/Y _49764_/Y sky130_fd_sc_hd__o21ai_4
X_46976_ _54473_/B _52781_/B sky130_fd_sc_hd__buf_2
X_42099_ _42083_/A _42099_/X sky130_fd_sc_hd__buf_2
X_77796_ _77796_/A _77796_/B _77796_/Y sky130_fd_sc_hd__nor2_4
X_48715_ _53620_/A _48099_/X _48723_/C _48715_/X sky130_fd_sc_hd__and3_4
X_79535_ _84203_/Q _72465_/A _79542_/A sky130_fd_sc_hd__nand2_4
X_45927_ _45922_/X _45923_/X _65880_/A _45926_/X _44184_/A _45927_/X
+ sky130_fd_sc_hd__a41o_4
X_64761_ _64757_/X _64761_/B _64760_/X _64761_/Y sky130_fd_sc_hd__nand3_4
X_76747_ _81693_/Q _76747_/B _76747_/Y sky130_fd_sc_hd__xnor2_4
X_49695_ _59360_/B _49687_/X _49694_/Y _49695_/Y sky130_fd_sc_hd__o21ai_4
X_61973_ _61719_/A _61973_/X sky130_fd_sc_hd__buf_2
X_73959_ _73957_/X _73945_/X _73947_/X _73959_/Y sky130_fd_sc_hd__nand3_4
X_66500_ _60110_/X _65281_/Y _66499_/Y _66500_/Y sky130_fd_sc_hd__o21ai_4
X_63712_ _58993_/Y _60748_/X _60654_/X _62629_/Y _60671_/B _63712_/Y
+ sky130_fd_sc_hd__o32ai_4
X_48646_ _48641_/Y _48585_/X _48645_/X _48646_/Y sky130_fd_sc_hd__a21oi_4
X_60924_ _60826_/A _60838_/X _76999_/A _60924_/Y sky130_fd_sc_hd__nor3_4
X_67480_ _67475_/X _67479_/X _67383_/X _67484_/A sky130_fd_sc_hd__a21o_4
X_79466_ _84813_/Q _84133_/Q _79466_/X sky130_fd_sc_hd__xor2_4
X_45858_ _45856_/Y _44968_/X _44875_/X _45857_/Y _45858_/X sky130_fd_sc_hd__a211o_4
X_64692_ _64766_/A _64692_/X sky130_fd_sc_hd__buf_2
X_76678_ _76686_/A _76969_/A _76678_/X sky130_fd_sc_hd__xor2_4
X_66431_ _64960_/X _66417_/B _64964_/X _66431_/Y sky130_fd_sc_hd__nand3_4
X_78417_ _78417_/A _82710_/Q _78418_/B sky130_fd_sc_hd__xor2_4
X_44809_ _44807_/X _43924_/X _41630_/X _86943_/Q _44808_/X _44810_/A
+ sky130_fd_sc_hd__o32ai_4
X_75629_ _81113_/Q _80825_/Q _75629_/X sky130_fd_sc_hd__xor2_4
X_63643_ _44173_/X _63644_/A sky130_fd_sc_hd__buf_2
X_48577_ _48563_/X _82350_/Q _48576_/Y _48578_/A sky130_fd_sc_hd__o21ai_4
X_60855_ _60854_/Y _60855_/X sky130_fd_sc_hd__buf_2
X_79397_ _79374_/X _79387_/X _79397_/Y sky130_fd_sc_hd__nand2_4
X_45789_ _63292_/B _61630_/A sky130_fd_sc_hd__buf_2
X_69150_ _69755_/A _87282_/Q _69150_/X sky130_fd_sc_hd__and2_4
X_47528_ _47553_/A _53101_/B _47528_/Y sky130_fd_sc_hd__nand2_4
X_66362_ _66294_/X _64582_/Y _66361_/Y _66362_/Y sky130_fd_sc_hd__o21ai_4
X_78348_ _78347_/X _78350_/A sky130_fd_sc_hd__inv_2
X_63574_ _61538_/B _63548_/X _63571_/X _63573_/Y _63574_/X sky130_fd_sc_hd__a211o_4
X_60786_ _60761_/A _60761_/B _84568_/Q _60786_/Y sky130_fd_sc_hd__nor3_4
X_68101_ _68120_/A _68101_/X sky130_fd_sc_hd__buf_2
X_65313_ _57788_/X _65313_/B _65313_/X sky130_fd_sc_hd__and2_4
X_62525_ _60085_/A _61582_/A _62522_/X _62524_/X _62525_/X sky130_fd_sc_hd__a211o_4
X_69081_ _69059_/A _88246_/Q _69081_/X sky130_fd_sc_hd__and2_4
X_47459_ _47459_/A _53060_/B sky130_fd_sc_hd__buf_2
X_66293_ _66291_/Y _66278_/X _66292_/X _84143_/D sky130_fd_sc_hd__a21o_4
X_78279_ _82590_/Q _78290_/B _78279_/X sky130_fd_sc_hd__xor2_4
X_68032_ _87446_/Q _67987_/X _67938_/X _68031_/X _68032_/X sky130_fd_sc_hd__a211o_4
X_80310_ _80309_/Y _80310_/B _80310_/Y sky130_fd_sc_hd__nand2_4
X_65244_ _64967_/X _65268_/A sky130_fd_sc_hd__buf_2
X_50470_ _50467_/Y _50455_/X _50469_/X _86195_/D sky130_fd_sc_hd__a21oi_4
X_62456_ _62454_/Y _62396_/X _62455_/Y _84409_/D sky130_fd_sc_hd__a21oi_4
X_81290_ _81275_/CLK _76978_/X _81258_/D sky130_fd_sc_hd__dfxtp_4
X_49129_ _49129_/A _49029_/B _49129_/Y sky130_fd_sc_hd__nor2_4
X_61407_ _61340_/A _61452_/B sky130_fd_sc_hd__buf_2
X_80241_ _80241_/A _80241_/B _80241_/X sky130_fd_sc_hd__xor2_4
X_65175_ _65159_/A _86027_/Q _65175_/X sky130_fd_sc_hd__and2_4
X_62387_ _62319_/A _58520_/A _62375_/C _62387_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_683_0_CLK clkbuf_9_341_0_CLK/X _87210_/CLK sky130_fd_sc_hd__clkbuf_1
X_52140_ _52198_/A _52140_/X sky130_fd_sc_hd__buf_2
X_64126_ _61629_/B _64161_/B _64150_/C _64161_/D _64126_/Y sky130_fd_sc_hd__nand4_4
X_61338_ _61338_/A _61367_/B _61367_/C _61367_/D _61338_/Y sky130_fd_sc_hd__nand4_4
X_80172_ _84945_/Q _65559_/C _80172_/Y sky130_fd_sc_hd__nand2_4
X_69983_ _82560_/D _69955_/X _69982_/X _69983_/X sky130_fd_sc_hd__a21bo_4
Xclkbuf_9_174_0_CLK clkbuf_8_87_0_CLK/X clkbuf_9_174_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_52071_ _66296_/B _52041_/X _52070_/Y _52071_/Y sky130_fd_sc_hd__o21ai_4
X_64057_ _60855_/X _64155_/C sky130_fd_sc_hd__buf_2
X_68934_ _65117_/A _68934_/X sky130_fd_sc_hd__buf_2
X_61269_ _61190_/X _61170_/Y _61267_/Y _64210_/A _61268_/Y _61269_/Y
+ sky130_fd_sc_hd__a41oi_4
X_84980_ _84980_/CLK _84980_/D _84980_/Q sky130_fd_sc_hd__dfxtp_4
X_51022_ _51022_/A _51022_/B _51022_/Y sky130_fd_sc_hd__nand2_4
X_63008_ _63130_/A _63008_/X sky130_fd_sc_hd__buf_2
X_83931_ _83932_/CLK _69339_/X _83931_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_698_0_CLK clkbuf_9_349_0_CLK/X _87221_/CLK sky130_fd_sc_hd__clkbuf_1
X_68865_ _68750_/A _88351_/Q _68865_/X sky130_fd_sc_hd__and2_4
X_55830_ _55830_/A _55830_/X sky130_fd_sc_hd__buf_2
X_67816_ _67816_/A _68479_/A sky130_fd_sc_hd__buf_2
X_86650_ _86647_/CLK _86650_/D _86650_/Q sky130_fd_sc_hd__dfxtp_4
X_83862_ _82553_/CLK _83862_/D _83862_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_189_0_CLK clkbuf_8_94_0_CLK/X clkbuf_9_189_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_68796_ _68938_/A _68796_/B _68796_/X sky130_fd_sc_hd__and2_4
X_85601_ _85601_/CLK _53621_/Y _85601_/Q sky130_fd_sc_hd__dfxtp_4
X_82813_ _81019_/CLK _82845_/Q _82813_/Q sky130_fd_sc_hd__dfxtp_4
X_55761_ _55761_/A _55761_/B _55761_/X sky130_fd_sc_hd__and2_4
X_67747_ _67863_/A _67747_/X sky130_fd_sc_hd__buf_2
X_86581_ _86582_/CLK _47966_/Y _66084_/B sky130_fd_sc_hd__dfxtp_4
X_52973_ _52979_/A _52973_/B _52973_/Y sky130_fd_sc_hd__nand2_4
X_64959_ _64807_/A _64959_/X sky130_fd_sc_hd__buf_2
X_83793_ _81620_/CLK _83793_/D _83793_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_621_0_CLK clkbuf_9_310_0_CLK/X _83974_/CLK sky130_fd_sc_hd__clkbuf_1
X_57500_ _84991_/Q _57493_/X _57499_/Y _57500_/Y sky130_fd_sc_hd__o21ai_4
X_88320_ _87813_/CLK _40869_/Y _69826_/B sky130_fd_sc_hd__dfxtp_4
X_54712_ _54699_/X _54734_/B _54721_/C _47391_/A _54712_/X sky130_fd_sc_hd__and4_4
X_85532_ _86045_/CLK _53970_/Y _85532_/Q sky130_fd_sc_hd__dfxtp_4
X_51924_ _52021_/A _57491_/C _51923_/Y _51924_/X sky130_fd_sc_hd__o21a_4
X_58480_ _58480_/A _58480_/Y sky130_fd_sc_hd__inv_2
X_82744_ _82152_/CLK _66415_/C _79011_/A sky130_fd_sc_hd__dfxtp_4
X_55692_ _55698_/A _56287_/C _55692_/X sky130_fd_sc_hd__and2_4
X_67678_ _68451_/A _67678_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_112_0_CLK clkbuf_8_56_0_CLK/X clkbuf_9_112_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_57431_ _44292_/A _57010_/A _57430_/X _57431_/Y sky130_fd_sc_hd__o21ai_4
X_69417_ _69413_/X _69416_/X _69171_/X _69417_/Y sky130_fd_sc_hd__a21oi_4
X_88251_ _87073_/CLK _41247_/Y _68970_/B sky130_fd_sc_hd__dfxtp_4
X_54643_ _54616_/X _54667_/A sky130_fd_sc_hd__buf_2
X_66629_ _66628_/X _66629_/X sky130_fd_sc_hd__buf_2
X_85463_ _82769_/CLK _85463_/D _85463_/Q sky130_fd_sc_hd__dfxtp_4
X_51855_ _51851_/A _51851_/B _51851_/C _52681_/D _51855_/X sky130_fd_sc_hd__and4_4
X_82675_ _82675_/CLK _82675_/D _78202_/A sky130_fd_sc_hd__dfxtp_4
X_87202_ _87720_/CLK _87202_/D _67752_/B sky130_fd_sc_hd__dfxtp_4
X_84414_ _84414_/CLK _84414_/D _84414_/Q sky130_fd_sc_hd__dfxtp_4
X_50806_ _50806_/A _51316_/B _50806_/Y sky130_fd_sc_hd__nand2_4
X_57362_ _56900_/X _56703_/X _57361_/Y _57362_/X sky130_fd_sc_hd__a21bo_4
X_81626_ _81279_/CLK _76518_/B _81626_/Q sky130_fd_sc_hd__dfxtp_4
X_69348_ _69309_/A _88292_/Q _69348_/X sky130_fd_sc_hd__and2_4
X_88182_ _87926_/CLK _88182_/D _67279_/B sky130_fd_sc_hd__dfxtp_4
X_54574_ _85417_/Q _54567_/X _54573_/Y _54574_/Y sky130_fd_sc_hd__o21ai_4
X_85394_ _85491_/CLK _85394_/D _85394_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_636_0_CLK clkbuf_9_318_0_CLK/X _82005_/CLK sky130_fd_sc_hd__clkbuf_1
X_51786_ _51814_/A _51794_/B sky130_fd_sc_hd__buf_2
X_59101_ _84769_/Q _59043_/X _59095_/X _59100_/X _84769_/D sky130_fd_sc_hd__a2bb2oi_4
X_56313_ _56309_/A _56312_/X _55908_/B _56313_/Y sky130_fd_sc_hd__nand3_4
X_87133_ _87484_/CLK _44390_/X _87133_/Q sky130_fd_sc_hd__dfxtp_4
X_53525_ _53503_/X _50300_/B _53525_/Y sky130_fd_sc_hd__nand2_4
X_84345_ _84849_/CLK _63200_/X _79343_/A sky130_fd_sc_hd__dfxtp_4
X_50737_ _50734_/Y _50735_/X _50736_/Y _50737_/Y sky130_fd_sc_hd__a21boi_4
X_57293_ _56824_/X _85039_/Q _57293_/Y sky130_fd_sc_hd__nand2_4
X_81557_ _84087_/CLK _76826_/X _81513_/D sky130_fd_sc_hd__dfxtp_4
X_69279_ _69253_/A _69279_/B _69279_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_127_0_CLK clkbuf_8_63_0_CLK/X clkbuf_9_127_0_CLK/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_9_54_0_CLK clkbuf_9_55_0_CLK/A clkbuf_9_54_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_59032_ _59027_/X _59029_/Y _59030_/Y _58959_/X _59031_/X _59032_/X
+ sky130_fd_sc_hd__o32a_4
X_71310_ _70819_/A _71333_/C sky130_fd_sc_hd__buf_2
X_80508_ _80504_/X _80520_/B _80513_/A sky130_fd_sc_hd__xor2_4
X_56244_ _56109_/X _56242_/X _56243_/Y _85262_/D sky130_fd_sc_hd__o21ai_4
X_41470_ _41469_/X _41455_/X _66634_/B _41457_/X _41470_/X sky130_fd_sc_hd__a2bb2o_4
X_87064_ _87063_/CLK _44536_/Y _87064_/Q sky130_fd_sc_hd__dfxtp_4
X_53456_ _53900_/A _53821_/B sky130_fd_sc_hd__buf_2
X_72290_ _72240_/X _85683_/Q _72241_/X _72290_/X sky130_fd_sc_hd__o21a_4
X_84276_ _84276_/CLK _84276_/D _64088_/C sky130_fd_sc_hd__dfxtp_4
X_50668_ _52365_/A _50651_/X _50668_/C _50668_/X sky130_fd_sc_hd__and3_4
X_81488_ _81361_/CLK _84056_/Q _81488_/Q sky130_fd_sc_hd__dfxtp_4
X_86015_ _85727_/CLK _86015_/D _86015_/Q sky130_fd_sc_hd__dfxtp_4
X_40421_ _47867_/A _40421_/X sky130_fd_sc_hd__buf_2
X_52407_ _52407_/A _49172_/A _52407_/X sky130_fd_sc_hd__and2_4
X_71241_ _71241_/A _71252_/A sky130_fd_sc_hd__buf_2
X_83227_ _83227_/CLK _72586_/Y _79363_/B sky130_fd_sc_hd__dfxtp_4
X_56175_ _56175_/A _56175_/B _56174_/X _56175_/Y sky130_fd_sc_hd__nand3_4
X_80439_ _80432_/X _80434_/B _80439_/Y sky130_fd_sc_hd__nand2_4
X_53387_ _85643_/Q _53378_/X _53386_/Y _53387_/Y sky130_fd_sc_hd__o21ai_4
X_50599_ _50599_/A _50599_/B _50599_/X sky130_fd_sc_hd__or2_4
X_43140_ _43140_/A _43140_/Y sky130_fd_sc_hd__inv_2
X_55126_ _55126_/A _55126_/X sky130_fd_sc_hd__buf_2
X_40352_ _40352_/A _46290_/A sky130_fd_sc_hd__buf_2
X_52338_ _52334_/A _52338_/B _52338_/Y sky130_fd_sc_hd__nand2_4
X_71172_ _50440_/B _71165_/X _71171_/Y _83584_/D sky130_fd_sc_hd__o21ai_4
X_83158_ _83158_/CLK _73272_/X _83158_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_69_0_CLK clkbuf_9_69_0_CLK/A clkbuf_9_69_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_70123_ _70123_/A _70125_/C sky130_fd_sc_hd__inv_2
X_82109_ _82860_/CLK _82109_/D _82109_/Q sky130_fd_sc_hd__dfxtp_4
X_43071_ _43053_/X _43054_/X _40678_/X _43070_/Y _43058_/X _87587_/D
+ sky130_fd_sc_hd__o32ai_4
X_55057_ _55043_/X _55056_/X _55070_/C _47701_/A _55057_/X sky130_fd_sc_hd__and4_4
X_59934_ _59917_/X _59943_/A sky130_fd_sc_hd__buf_2
X_52269_ _52214_/A _52269_/X sky130_fd_sc_hd__buf_2
X_75980_ _75980_/A _75980_/B _75980_/Y sky130_fd_sc_hd__nand2_4
X_83089_ _81627_/CLK _83089_/D _83089_/Q sky130_fd_sc_hd__dfxtp_4
X_87966_ _87720_/CLK _42237_/X _87966_/Q sky130_fd_sc_hd__dfxtp_4
X_42022_ _42013_/X _42006_/X _40849_/X _73175_/A _42007_/X _42023_/A
+ sky130_fd_sc_hd__o32ai_4
X_54008_ _54005_/Y _54006_/X _54007_/Y _54008_/Y sky130_fd_sc_hd__a21boi_4
X_74931_ _74923_/A _81132_/D _74912_/B _74931_/Y sky130_fd_sc_hd__nand3_4
X_70054_ _70054_/A _70053_/X _70021_/C _70054_/Y sky130_fd_sc_hd__nand3_4
X_86917_ _86914_/CLK _86917_/D _67964_/B sky130_fd_sc_hd__dfxtp_4
X_59865_ _59811_/Y _59758_/X _59862_/X _59783_/Y _59864_/Y _59865_/Y
+ sky130_fd_sc_hd__a41oi_4
X_87897_ _87195_/CLK _87897_/D _87897_/Q sky130_fd_sc_hd__dfxtp_4
X_46830_ _46830_/A _46830_/B _46830_/C _52698_/D _46830_/X sky130_fd_sc_hd__and4_4
X_58816_ _58812_/Y _58815_/Y _58735_/X _58816_/X sky130_fd_sc_hd__a21o_4
X_77650_ _77650_/A _77650_/B _77650_/Y sky130_fd_sc_hd__nor2_4
X_74862_ _74863_/B _81156_/D sky130_fd_sc_hd__inv_2
X_86848_ _84420_/CLK _45880_/Y _64190_/A sky130_fd_sc_hd__dfxtp_4
X_59796_ _59727_/X _59790_/X _59745_/X _59794_/X _59795_/Y _84699_/D
+ sky130_fd_sc_hd__a41oi_4
X_76601_ _76597_/X _76598_/Y _76602_/B _76614_/B sky130_fd_sc_hd__a21o_4
X_73813_ _57537_/B _73813_/B _73813_/X sky130_fd_sc_hd__xor2_4
X_46761_ _46667_/A _46784_/C sky130_fd_sc_hd__buf_2
X_58747_ _64600_/A _58864_/A sky130_fd_sc_hd__buf_2
X_77581_ _77582_/A _82118_/Q _77584_/B sky130_fd_sc_hd__nor2_4
X_43973_ _44067_/B _43944_/A _43945_/Y _43972_/Y _43973_/X sky130_fd_sc_hd__a211o_4
X_55959_ _85278_/Q _55689_/A _44052_/X _55958_/X _55959_/X sky130_fd_sc_hd__a211o_4
X_74793_ _83807_/Q _74738_/A _74787_/Y _74788_/Y _74792_/X _74793_/X
+ sky130_fd_sc_hd__a2111o_4
X_86779_ _81182_/CLK _86779_/D _67227_/B sky130_fd_sc_hd__dfxtp_4
X_48500_ _48635_/A _48500_/X sky130_fd_sc_hd__buf_2
X_79320_ _84799_/Q _82735_/D _79320_/X sky130_fd_sc_hd__xor2_4
X_45712_ _45272_/A _45746_/B sky130_fd_sc_hd__buf_2
X_76532_ _81276_/Q _76533_/B _76535_/B sky130_fd_sc_hd__nor2_4
X_42924_ _41721_/X _42920_/X _87650_/Q _42922_/X _87650_/D sky130_fd_sc_hd__a2bb2o_4
X_49480_ _49477_/Y _49460_/X _49479_/X _49480_/Y sky130_fd_sc_hd__a21oi_4
X_73744_ _73739_/X _73743_/X _73745_/B sky130_fd_sc_hd__nand2_4
X_46692_ _83681_/Q _54309_/B sky130_fd_sc_hd__inv_2
X_70956_ _70944_/A _70969_/A sky130_fd_sc_hd__buf_2
X_58678_ _58585_/X _58675_/Y _58677_/Y _58603_/X _58589_/X _58678_/X
+ sky130_fd_sc_hd__o32a_4
X_48431_ _48744_/A _48364_/X _48476_/C _48431_/X sky130_fd_sc_hd__and3_4
X_79251_ _79251_/A _79251_/B _79251_/Y sky130_fd_sc_hd__nor2_4
X_45643_ _85105_/Q _45643_/Y sky130_fd_sc_hd__inv_2
X_57629_ _57626_/Y _57627_/X _57628_/Y _84966_/D sky130_fd_sc_hd__a21boi_4
X_76463_ _76458_/Y _76459_/Y _76454_/X _76457_/Y _76463_/X sky130_fd_sc_hd__a211o_4
X_42855_ _41529_/X _42852_/X _66900_/B _42853_/X _87685_/D sky130_fd_sc_hd__a2bb2o_4
X_73675_ _73675_/A _73649_/X _73675_/Y sky130_fd_sc_hd__nor2_4
X_70887_ _70905_/D _70890_/D sky130_fd_sc_hd__buf_2
X_78202_ _78202_/A _78202_/B _78202_/X sky130_fd_sc_hd__xor2_4
X_75414_ _75413_/B _75413_/C _75413_/A _75414_/Y sky130_fd_sc_hd__o21ai_4
X_41806_ _40387_/X _41799_/X _88144_/Q _41800_/X _88144_/D sky130_fd_sc_hd__a2bb2o_4
X_48362_ _48043_/X _81793_/Q _48361_/Y _74366_/A sky130_fd_sc_hd__o21ai_4
X_60640_ _59613_/Y _60183_/A _61075_/C _60641_/A sky130_fd_sc_hd__nand3_4
X_72626_ _72581_/A _72604_/B _79168_/A _72626_/Y sky130_fd_sc_hd__nor3_4
X_79182_ _79180_/Y _79181_/Y _79185_/A sky130_fd_sc_hd__nand2_4
X_45574_ _45568_/X _45573_/X _45523_/X _45574_/X sky130_fd_sc_hd__a21o_4
X_76394_ _76394_/A _76394_/Y sky130_fd_sc_hd__inv_2
X_42786_ _41352_/X _42767_/X _67613_/B _42768_/X _42786_/X sky130_fd_sc_hd__a2bb2o_4
X_47313_ _47313_/A _47313_/Y sky130_fd_sc_hd__inv_2
X_78133_ _82569_/Q _78124_/B _78134_/B sky130_fd_sc_hd__nor2_4
X_44525_ _44524_/Y _87067_/D sky130_fd_sc_hd__inv_2
X_75345_ _75364_/A _75345_/B _75345_/X sky130_fd_sc_hd__xor2_4
X_41737_ _41672_/X _41673_/X _41735_/X _67826_/B _41736_/X _41737_/Y
+ sky130_fd_sc_hd__o32ai_4
X_48293_ _48169_/X _48293_/X sky130_fd_sc_hd__buf_2
X_60571_ _60413_/X _60571_/B _60571_/Y sky130_fd_sc_hd__nand2_4
X_72557_ _72517_/A _72557_/Y sky130_fd_sc_hd__inv_2
X_62310_ _62634_/A _62307_/Y _62310_/C _62310_/D _62310_/Y sky130_fd_sc_hd__nand4_4
X_47244_ _47241_/X _52936_/B _47244_/Y sky130_fd_sc_hd__nand2_4
X_71508_ _71525_/A _71508_/X sky130_fd_sc_hd__buf_2
X_78064_ _78064_/A _78064_/B _78064_/X sky130_fd_sc_hd__xor2_4
X_44456_ _44447_/X _44448_/X _41124_/X _87101_/Q _44449_/X _44457_/A
+ sky130_fd_sc_hd__o32ai_4
X_63290_ _60606_/X _63341_/C sky130_fd_sc_hd__buf_2
X_75276_ _75271_/X _75274_/Y _75272_/Y _75276_/Y sky130_fd_sc_hd__nand3_4
X_41668_ _41607_/X _41668_/X sky130_fd_sc_hd__buf_2
X_72488_ _63573_/A _72488_/B _72488_/Y sky130_fd_sc_hd__nand2_4
X_77015_ _77015_/A _77014_/Y _77017_/B sky130_fd_sc_hd__xnor2_4
X_43407_ _43329_/X _43407_/X sky130_fd_sc_hd__buf_2
X_62241_ _62181_/A _62181_/B _84424_/Q _62241_/Y sky130_fd_sc_hd__nor3_4
X_74227_ _43103_/Y _56273_/X _73035_/X _74226_/Y _74227_/X sky130_fd_sc_hd__a211o_4
X_40619_ _40413_/X _48461_/A sky130_fd_sc_hd__buf_2
X_47175_ _47150_/A _47174_/X _47175_/Y sky130_fd_sc_hd__nand2_4
X_71439_ _70370_/A _71435_/B _71439_/C _71432_/D _71439_/X sky130_fd_sc_hd__and4_4
X_44387_ _44387_/A _44387_/Y sky130_fd_sc_hd__inv_2
X_41599_ _41358_/X _82310_/Q _41599_/X sky130_fd_sc_hd__or2_4
X_46126_ _46092_/X _46121_/A _46128_/A sky130_fd_sc_hd__nor2_4
X_43338_ _41298_/X _43336_/X _87473_/Q _43337_/X _87473_/D sky130_fd_sc_hd__a2bb2o_4
X_62172_ _61683_/X _62149_/B _61765_/C _61749_/B _62172_/Y sky130_fd_sc_hd__nand4_4
X_74158_ _74155_/X _84968_/Q _74087_/X _74157_/X _74158_/X sky130_fd_sc_hd__a211o_4
X_61123_ _64421_/A _64306_/A sky130_fd_sc_hd__buf_2
X_73109_ _69737_/B _73227_/A _72979_/X _73108_/Y _73109_/X sky130_fd_sc_hd__a211o_4
X_46057_ _46046_/X _46054_/X _41544_/X _66962_/B _46047_/X _46058_/A
+ sky130_fd_sc_hd__o32ai_4
X_43269_ _43167_/A _43269_/X sky130_fd_sc_hd__buf_2
X_66980_ _66977_/X _66979_/X _66980_/Y sky130_fd_sc_hd__nand2_4
X_74089_ _73566_/X _84971_/Q _74087_/X _74088_/X _74090_/B sky130_fd_sc_hd__a211o_4
X_78966_ _78966_/A _78968_/A sky130_fd_sc_hd__inv_2
X_45008_ _45005_/X _45007_/Y _44973_/X _45008_/Y sky130_fd_sc_hd__a21oi_4
X_65931_ _65928_/Y _65915_/X _65930_/X _84168_/D sky130_fd_sc_hd__a21o_4
X_61054_ _60599_/A _61051_/Y _60403_/B _60980_/Y _61053_/Y _84527_/D
+ sky130_fd_sc_hd__a41oi_4
X_77917_ _82166_/Q _82038_/D _82134_/D sky130_fd_sc_hd__xor2_4
X_78897_ _78885_/A _78885_/B _78870_/A _82506_/D _78897_/X sky130_fd_sc_hd__a2bb2o_4
X_60005_ _59913_/X _59985_/X _59881_/X _59884_/X _65842_/A _60005_/Y
+ sky130_fd_sc_hd__a41oi_4
X_49816_ _48499_/A _49925_/A sky130_fd_sc_hd__buf_2
X_68650_ _69007_/A _68650_/X sky130_fd_sc_hd__buf_2
X_65862_ _65859_/X _85572_/Q _65860_/X _65861_/X _65862_/X sky130_fd_sc_hd__a211o_4
X_77848_ _77841_/Y _77842_/A _77847_/Y _77849_/B sky130_fd_sc_hd__a21oi_4
X_67601_ _86964_/Q _67551_/X _67552_/X _67600_/X _67602_/B sky130_fd_sc_hd__a211o_4
X_64813_ _64561_/X _64800_/Y _64812_/Y _64813_/Y sky130_fd_sc_hd__o21ai_4
X_49747_ _49745_/Y _49732_/X _49746_/X _86331_/D sky130_fd_sc_hd__a21oi_4
X_68581_ _68560_/A _88267_/Q _68581_/X sky130_fd_sc_hd__and2_4
X_46959_ _46959_/A _52773_/B _46959_/Y sky130_fd_sc_hd__nand2_4
X_65793_ _65623_/X _86185_/Q _65790_/X _65792_/X _65793_/X sky130_fd_sc_hd__a211o_4
X_77779_ _77771_/Y _77779_/Y sky130_fd_sc_hd__inv_2
X_67532_ _67532_/A _67531_/X _67532_/Y sky130_fd_sc_hd__nand2_4
X_79518_ _79513_/X _79518_/B _79519_/A sky130_fd_sc_hd__xnor2_4
X_64744_ _64650_/X _86140_/Q _64583_/X _64743_/X _64744_/X sky130_fd_sc_hd__a211o_4
X_49678_ _49406_/A _49678_/X sky130_fd_sc_hd__buf_2
X_61956_ _61954_/X _61924_/B _61971_/C _61910_/D _61956_/Y sky130_fd_sc_hd__nand4_4
X_80790_ _80931_/CLK _75883_/Y _75371_/A sky130_fd_sc_hd__dfxtp_4
X_48629_ _86505_/Q _48612_/X _48628_/Y _48629_/Y sky130_fd_sc_hd__o21ai_4
X_60907_ _60906_/X _60908_/A sky130_fd_sc_hd__buf_2
X_67463_ _67513_/A _86938_/Q _67463_/X sky130_fd_sc_hd__and2_4
X_79449_ _79449_/A _79448_/Y _79459_/B sky130_fd_sc_hd__xor2_4
X_64675_ _64672_/X _64674_/X _64675_/Y sky130_fd_sc_hd__nand2_4
X_61887_ _57660_/X _61824_/X _61838_/X _61870_/X _61886_/X _61887_/X
+ sky130_fd_sc_hd__a41o_4
X_69202_ _69088_/A _69202_/X sky130_fd_sc_hd__buf_2
X_66414_ _66377_/A _66414_/X sky130_fd_sc_hd__buf_2
X_51640_ _51694_/A _51651_/B sky130_fd_sc_hd__buf_2
X_63626_ _63436_/A _63626_/X sky130_fd_sc_hd__buf_2
X_82460_ _84187_/CLK _79152_/X _82428_/D sky130_fd_sc_hd__dfxtp_4
X_60838_ _60715_/X _60838_/X sky130_fd_sc_hd__buf_2
X_67394_ _66915_/A _67394_/X sky130_fd_sc_hd__buf_2
X_81411_ _84014_/CLK _81443_/Q _75927_/B sky130_fd_sc_hd__dfxtp_4
X_69133_ _80802_/D _69066_/X _69132_/X _83946_/D sky130_fd_sc_hd__a21bo_4
X_66345_ _66177_/A _66389_/B _66345_/C _66345_/Y sky130_fd_sc_hd__nor3_4
X_51571_ _51569_/Y _51557_/X _51570_/X _51571_/Y sky130_fd_sc_hd__a21oi_4
X_63557_ _63546_/A _63557_/B _63520_/C _63546_/D _63557_/X sky130_fd_sc_hd__and4_4
X_82391_ _82390_/CLK _82391_/D _82391_/Q sky130_fd_sc_hd__dfxtp_4
X_60769_ _60376_/X _60765_/Y _60767_/X _60690_/X _60768_/X _60769_/X
+ sky130_fd_sc_hd__o41a_4
X_53310_ _85657_/Q _53295_/X _53309_/Y _53310_/Y sky130_fd_sc_hd__o21ai_4
X_84130_ _84175_/CLK _84130_/D _79435_/B sky130_fd_sc_hd__dfxtp_4
X_50522_ _86184_/Q _50506_/X _50521_/Y _50522_/Y sky130_fd_sc_hd__o21ai_4
X_62508_ _62276_/X _62601_/C sky130_fd_sc_hd__buf_2
X_81342_ _81473_/CLK _76592_/X _81718_/D sky130_fd_sc_hd__dfxtp_4
X_69064_ _83949_/Q _68954_/X _69063_/X _83949_/D sky130_fd_sc_hd__a21bo_4
X_54290_ _54316_/A _54312_/A sky130_fd_sc_hd__buf_2
X_66276_ _65810_/X _66276_/B _65813_/X _66276_/Y sky130_fd_sc_hd__nand3_4
X_63488_ _63488_/A _61891_/X _63488_/X sky130_fd_sc_hd__and2_4
X_68015_ _68011_/X _68014_/X _67875_/X _68015_/Y sky130_fd_sc_hd__a21oi_4
X_65227_ _65227_/A _86249_/Q _65227_/X sky130_fd_sc_hd__and2_4
X_53241_ _85670_/Q _53225_/X _53240_/Y _53241_/Y sky130_fd_sc_hd__o21ai_4
X_84061_ _82648_/CLK _84061_/D _84061_/Q sky130_fd_sc_hd__dfxtp_4
X_50453_ _50439_/X _52158_/B _50453_/Y sky130_fd_sc_hd__nand2_4
X_62439_ _61509_/B _62390_/X _62436_/X _62407_/X _62438_/X _62439_/X
+ sky130_fd_sc_hd__a41o_4
X_81273_ _81304_/CLK _81305_/Q _76489_/A sky130_fd_sc_hd__dfxtp_4
X_83012_ _83012_/CLK _83012_/D _45345_/A sky130_fd_sc_hd__dfxtp_4
X_80224_ _80207_/Y _80204_/Y _80209_/A _80209_/B _80224_/X sky130_fd_sc_hd__a211o_4
X_53172_ _53172_/A _53172_/X sky130_fd_sc_hd__buf_2
X_65158_ _65158_/A _65159_/A sky130_fd_sc_hd__buf_2
X_50384_ _86211_/Q _50363_/X _50383_/Y _50384_/Y sky130_fd_sc_hd__o21ai_4
X_52123_ _52188_/A _52123_/B _52123_/Y sky130_fd_sc_hd__nand2_4
X_64109_ _64107_/Y _64073_/X _64108_/Y _84274_/D sky130_fd_sc_hd__a21oi_4
X_87820_ _87820_/CLK _87820_/D _72945_/A sky130_fd_sc_hd__dfxtp_4
X_80155_ _80151_/Y _80169_/B _80178_/A sky130_fd_sc_hd__xor2_4
X_65089_ _65086_/X _65192_/B _65088_/X _65089_/Y sky130_fd_sc_hd__nand3_4
X_57980_ _84934_/Q _57980_/Y sky130_fd_sc_hd__inv_2
X_69966_ _83883_/Q _69955_/X _69965_/X _83883_/D sky130_fd_sc_hd__a21bo_4
X_52054_ _52058_/A _57609_/B _52054_/Y sky130_fd_sc_hd__nand2_4
X_56931_ _56931_/A _56931_/X sky130_fd_sc_hd__buf_2
X_68917_ _69233_/A _68987_/A sky130_fd_sc_hd__buf_2
X_87751_ _87758_/CLK _42725_/Y _87751_/Q sky130_fd_sc_hd__dfxtp_4
X_84963_ _85599_/CLK _57645_/Y _84963_/Q sky130_fd_sc_hd__dfxtp_4
X_80086_ _80072_/Y _80077_/Y _80085_/X _80087_/B sky130_fd_sc_hd__o21ai_4
X_69897_ _69897_/A _69897_/B _69897_/Y sky130_fd_sc_hd__nor2_4
X_51005_ _50952_/A _51029_/C sky130_fd_sc_hd__buf_2
X_86702_ _86381_/CLK _86702_/D _58807_/A sky130_fd_sc_hd__dfxtp_4
X_59650_ _59649_/Y _59651_/C sky130_fd_sc_hd__inv_2
X_83914_ _83914_/CLK _83914_/D _83914_/Q sky130_fd_sc_hd__dfxtp_4
X_56862_ _57346_/C _56860_/X _56893_/B _56862_/Y sky130_fd_sc_hd__nand3_4
X_68848_ _68779_/A _68848_/B _68848_/X sky130_fd_sc_hd__and2_4
X_87682_ _88128_/CLK _42861_/X _66982_/B sky130_fd_sc_hd__dfxtp_4
X_84894_ _84894_/CLK _84894_/D _62027_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_560_0_CLK clkbuf_9_280_0_CLK/X _81703_/CLK sky130_fd_sc_hd__clkbuf_1
X_58601_ _58601_/A _58614_/B _58601_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_6_51_0_CLK clkbuf_6_51_0_CLK/A clkbuf_6_51_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_55813_ _56243_/C _55311_/X _44046_/X _55812_/X _55813_/X sky130_fd_sc_hd__a211o_4
X_86633_ _85993_/CLK _47457_/Y _86633_/Q sky130_fd_sc_hd__dfxtp_4
X_83845_ _83843_/CLK _83845_/D _83845_/Q sky130_fd_sc_hd__dfxtp_4
X_59581_ _59546_/A _59563_/A _59581_/C _59582_/B sky130_fd_sc_hd__nand3_4
X_56793_ _55399_/X _56707_/X _55409_/Y _56797_/A sky130_fd_sc_hd__nand3_4
X_68779_ _68779_/A _87331_/Q _68779_/X sky130_fd_sc_hd__and2_4
X_70810_ _70810_/A _70942_/B _70810_/C _70810_/Y sky130_fd_sc_hd__nand3_4
X_58532_ _57673_/A _58532_/X sky130_fd_sc_hd__buf_2
X_55744_ _55740_/Y _44095_/A _55743_/Y _55745_/D sky130_fd_sc_hd__a21oi_4
X_86564_ _86490_/CLK _86564_/D _74234_/B sky130_fd_sc_hd__dfxtp_4
X_40970_ _40800_/B _40970_/B _40970_/X sky130_fd_sc_hd__or2_4
X_52956_ _52515_/A _53065_/A sky130_fd_sc_hd__buf_2
X_71790_ _71235_/A _70472_/X _71785_/X _71790_/Y sky130_fd_sc_hd__nand3_4
X_83776_ _86553_/CLK _83776_/D _83776_/Q sky130_fd_sc_hd__dfxtp_4
X_80988_ _80849_/CLK _80988_/D _80944_/D sky130_fd_sc_hd__dfxtp_4
X_88303_ _88097_/CLK _88303_/D _88303_/Q sky130_fd_sc_hd__dfxtp_4
X_85515_ _86029_/CLK _54053_/Y _85515_/Q sky130_fd_sc_hd__dfxtp_4
X_51907_ _51902_/A _51043_/B _51907_/Y sky130_fd_sc_hd__nand2_4
X_70741_ _53101_/B _70738_/X _70740_/Y _70741_/Y sky130_fd_sc_hd__o21ai_4
X_58463_ _83474_/Q _58463_/Y sky130_fd_sc_hd__inv_2
X_82727_ _81190_/CLK _84111_/Q _82727_/Q sky130_fd_sc_hd__dfxtp_4
X_55675_ _55671_/Y _55675_/B _55675_/X sky130_fd_sc_hd__xor2_4
X_86495_ _85888_/CLK _86495_/D _65455_/B sky130_fd_sc_hd__dfxtp_4
X_52887_ _52867_/A _52879_/B _52872_/C _52887_/D _52887_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_575_0_CLK clkbuf_9_287_0_CLK/X _82886_/CLK sky130_fd_sc_hd__clkbuf_1
X_57414_ _57414_/A _57413_/X _57414_/X sky130_fd_sc_hd__or2_4
X_88234_ _88164_/CLK _88234_/D _67553_/B sky130_fd_sc_hd__dfxtp_4
X_54626_ _54624_/Y _54611_/X _54625_/X _85408_/D sky130_fd_sc_hd__a21oi_4
X_42640_ _40955_/X _42631_/X _69176_/B _42634_/X _42640_/X sky130_fd_sc_hd__a2bb2o_4
X_73460_ _73339_/A _73460_/B _73460_/Y sky130_fd_sc_hd__nor2_4
X_85446_ _85447_/CLK _85446_/D _85446_/Q sky130_fd_sc_hd__dfxtp_4
X_51838_ _51851_/A _51815_/B _51851_/C _46775_/X _51838_/X sky130_fd_sc_hd__and4_4
X_70672_ _70543_/Y _70673_/A sky130_fd_sc_hd__buf_2
X_82658_ _82498_/CLK _82658_/D _78082_/A sky130_fd_sc_hd__dfxtp_4
X_58394_ _58393_/Y _58403_/B _58394_/Y sky130_fd_sc_hd__nand2_4
X_72411_ _72408_/Y _72410_/Y _72344_/X _72411_/X sky130_fd_sc_hd__a21o_4
X_81609_ _81801_/CLK _76258_/Y _81609_/Q sky130_fd_sc_hd__dfxtp_4
X_57345_ _56873_/X _57322_/B _57351_/A sky130_fd_sc_hd__nand2_4
X_88165_ _87915_/CLK _88165_/D _67683_/B sky130_fd_sc_hd__dfxtp_4
X_42571_ _42556_/A _42571_/X sky130_fd_sc_hd__buf_2
X_54557_ _54284_/A _54558_/A sky130_fd_sc_hd__buf_2
X_73391_ _73339_/A _73391_/B _73391_/Y sky130_fd_sc_hd__nor2_4
X_85377_ _83711_/CLK _85377_/D _85377_/Q sky130_fd_sc_hd__dfxtp_4
X_51769_ _51766_/Y _51767_/X _51768_/X _51769_/Y sky130_fd_sc_hd__a21oi_4
X_82589_ _82589_/CLK _82621_/Q _78273_/A sky130_fd_sc_hd__dfxtp_4
X_44310_ _57470_/B _44318_/A sky130_fd_sc_hd__buf_2
X_75130_ _75126_/X _75143_/A _75129_/Y _75130_/Y sky130_fd_sc_hd__a21oi_4
X_41522_ _41522_/A _41522_/Y sky130_fd_sc_hd__inv_2
X_87116_ _87116_/CLK _87116_/D _87116_/Q sky130_fd_sc_hd__dfxtp_4
X_53508_ _53723_/A _53509_/A sky130_fd_sc_hd__buf_2
X_72342_ _72258_/X _85679_/Q _72308_/X _72342_/X sky130_fd_sc_hd__o21a_4
X_84328_ _84355_/CLK _84328_/D _80614_/B sky130_fd_sc_hd__dfxtp_4
X_57276_ _57271_/Y _57274_/Y _57275_/X _57276_/X sky130_fd_sc_hd__a21o_4
X_45290_ _45290_/A _45290_/Y sky130_fd_sc_hd__inv_2
X_88096_ _88104_/CLK _41948_/Y _88096_/Q sky130_fd_sc_hd__dfxtp_4
X_54488_ _85433_/Q _54485_/X _54487_/Y _54488_/Y sky130_fd_sc_hd__o21ai_4
X_59015_ _59001_/X _86080_/Q _59014_/X _59015_/Y sky130_fd_sc_hd__o21ai_4
X_44241_ _44139_/X _44141_/X _44142_/X _44225_/Y _44241_/Y sky130_fd_sc_hd__nand4_4
X_56227_ _56233_/A _56229_/B _85268_/Q _56227_/Y sky130_fd_sc_hd__nand3_4
X_75061_ _80744_/Q _75061_/B _75067_/B sky130_fd_sc_hd__xor2_4
X_87047_ _88326_/CLK _87047_/D _73370_/A sky130_fd_sc_hd__dfxtp_4
X_41453_ _41449_/X _82882_/Q _41452_/X _41453_/Y sky130_fd_sc_hd__o21ai_4
X_53439_ _53420_/A _53428_/X _54111_/C _47218_/D _53439_/X sky130_fd_sc_hd__and4_4
X_72273_ _86613_/Q _72332_/B _72273_/Y sky130_fd_sc_hd__nor2_4
X_84259_ _84314_/CLK _64291_/X _79817_/B sky130_fd_sc_hd__dfxtp_4
X_74012_ _74012_/A _74012_/X sky130_fd_sc_hd__buf_2
X_40404_ _40403_/Y _40404_/X sky130_fd_sc_hd__buf_2
X_71224_ _48847_/B _71216_/X _71223_/Y _71224_/Y sky130_fd_sc_hd__o21ai_4
X_44172_ _44247_/A _44315_/A sky130_fd_sc_hd__buf_2
X_56158_ _56158_/A _56157_/Y _56159_/A sky130_fd_sc_hd__xor2_4
X_41384_ _41383_/Y _88225_/D sky130_fd_sc_hd__inv_2
Xclkbuf_10_513_0_CLK clkbuf_9_256_0_CLK/X _81461_/CLK sky130_fd_sc_hd__clkbuf_1
X_43123_ _43123_/A _43123_/Y sky130_fd_sc_hd__inv_2
X_55109_ _55107_/Y _55102_/X _55108_/X _55109_/Y sky130_fd_sc_hd__a21oi_4
X_78820_ _78810_/Y _78820_/B _78821_/B sky130_fd_sc_hd__xnor2_4
X_40335_ _40321_/A _40335_/B _43175_/A sky130_fd_sc_hd__nand2_4
X_71155_ _71181_/A _71155_/B _71160_/C _71160_/D _71155_/Y sky130_fd_sc_hd__nand4_4
X_48980_ _48975_/Y _48935_/X _48979_/X _48980_/Y sky130_fd_sc_hd__a21oi_4
X_56089_ _55845_/B _55844_/X _56089_/X sky130_fd_sc_hd__and2_4
X_70106_ _83136_/Q _70106_/Y sky130_fd_sc_hd__inv_2
X_47931_ _53501_/B _47932_/B sky130_fd_sc_hd__buf_2
X_43054_ _43046_/A _43054_/X sky130_fd_sc_hd__buf_2
X_59917_ _59917_/A _59904_/B _60155_/C _59917_/X sky130_fd_sc_hd__and3_4
X_78751_ _78750_/A _82687_/D _78752_/A sky130_fd_sc_hd__nand2_4
X_71086_ _71088_/A _71230_/B _71088_/C _71086_/Y sky130_fd_sc_hd__nand3_4
X_75963_ _75956_/Y _75961_/Y _75963_/C _75963_/Y sky130_fd_sc_hd__nand3_4
X_87949_ _87952_/CLK _87949_/D _87949_/Q sky130_fd_sc_hd__dfxtp_4
X_42005_ _41998_/X _41993_/X _40810_/X _42004_/Y _42000_/X _88074_/D
+ sky130_fd_sc_hd__o32ai_4
X_77702_ _77702_/A _77703_/C sky130_fd_sc_hd__inv_2
X_74914_ _74904_/Y _74914_/B _74914_/Y sky130_fd_sc_hd__nand2_4
X_70037_ _68749_/X _68751_/X _70005_/X _70037_/Y sky130_fd_sc_hd__a21oi_4
X_47862_ _47856_/Y _47846_/X _47861_/X _47862_/Y sky130_fd_sc_hd__a21oi_4
X_59848_ _59855_/A _59848_/B _80371_/A _59848_/Y sky130_fd_sc_hd__nor3_4
X_78682_ _78682_/A _78682_/B _78682_/C _78684_/A sky130_fd_sc_hd__or3_4
Xclkbuf_10_528_0_CLK clkbuf_9_264_0_CLK/X _83940_/CLK sky130_fd_sc_hd__clkbuf_1
X_75894_ _84492_/Q _84364_/Q _80708_/D sky130_fd_sc_hd__xor2_4
Xclkbuf_6_19_0_CLK clkbuf_5_9_0_CLK/X clkbuf_7_39_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_49601_ _86357_/Q _49579_/X _49600_/Y _49601_/Y sky130_fd_sc_hd__o21ai_4
X_46813_ _46767_/A _46813_/X sky130_fd_sc_hd__buf_2
X_77633_ _77629_/Y _77633_/B _77632_/Y _77633_/X sky130_fd_sc_hd__or3_4
X_74845_ _74844_/Y _80652_/D sky130_fd_sc_hd__inv_2
X_47793_ _81221_/Q _47794_/A sky130_fd_sc_hd__inv_2
X_59779_ _59758_/X _59775_/X _59724_/Y _59744_/Y _59778_/Y _59780_/A
+ sky130_fd_sc_hd__a41o_4
X_49532_ _49614_/A _49537_/B sky130_fd_sc_hd__buf_2
X_61810_ _61386_/B _61795_/B _61795_/C _61778_/X _61810_/Y sky130_fd_sc_hd__nand4_4
X_46744_ _46743_/Y _46744_/X sky130_fd_sc_hd__buf_2
X_77564_ _77560_/Y _77564_/B _82200_/D sky130_fd_sc_hd__xor2_4
X_43956_ _80667_/Q _43957_/A sky130_fd_sc_hd__inv_2
X_62790_ _62784_/Y _62772_/X _62785_/Y _62787_/Y _62789_/X _62790_/X
+ sky130_fd_sc_hd__a41o_4
X_74776_ _83845_/Q _74735_/X _74773_/X _74774_/X _74775_/X _74776_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_71988_ _83307_/Q _71985_/X _71987_/Y _71988_/Y sky130_fd_sc_hd__o21ai_4
X_79303_ _79303_/A _79302_/Y _79303_/X sky130_fd_sc_hd__xor2_4
X_76515_ _76513_/C _76513_/D _76513_/B _76515_/X sky130_fd_sc_hd__a21bo_4
X_42907_ _42907_/A _87659_/D sky130_fd_sc_hd__inv_2
X_49463_ _49459_/Y _49460_/X _49462_/X _86383_/D sky130_fd_sc_hd__a21oi_4
X_61741_ _61777_/A _61761_/C sky130_fd_sc_hd__buf_2
X_73727_ _73724_/X _73726_/X _73679_/X _73727_/X sky130_fd_sc_hd__a21o_4
X_70939_ _70939_/A _70947_/C sky130_fd_sc_hd__buf_2
X_46675_ _83683_/Q _46676_/A sky130_fd_sc_hd__inv_2
X_77495_ _77495_/A _77493_/Y _77491_/Y _77495_/Y sky130_fd_sc_hd__nand3_4
X_43887_ _43869_/X _43887_/X sky130_fd_sc_hd__buf_2
X_48414_ _81788_/Q _48136_/B _48414_/X sky130_fd_sc_hd__or2_4
X_79234_ _79232_/B _79230_/Y _79235_/B sky130_fd_sc_hd__nand2_4
X_45626_ _85106_/Q _45626_/Y sky130_fd_sc_hd__inv_2
X_76446_ _76425_/X _76444_/Y _76445_/Y _76446_/X sky130_fd_sc_hd__a21bo_4
X_64460_ _61135_/X _84836_/Q _64458_/X _64459_/Y _64460_/X sky130_fd_sc_hd__a211o_4
X_42838_ _42837_/Y _87693_/D sky130_fd_sc_hd__inv_2
X_49394_ _49410_/A _51779_/B _49394_/Y sky130_fd_sc_hd__nand2_4
X_61672_ _61670_/X _61645_/X _61671_/Y _61672_/Y sky130_fd_sc_hd__a21oi_4
X_73658_ _87003_/Q _56550_/X _73657_/X _73658_/Y sky130_fd_sc_hd__o21ai_4
X_63411_ _58418_/A _63370_/X _61378_/A _63372_/X _63411_/X sky130_fd_sc_hd__a2bb2o_4
X_48345_ _48401_/A _50383_/B _48345_/Y sky130_fd_sc_hd__nand2_4
X_60623_ _60655_/A _60624_/A sky130_fd_sc_hd__inv_2
X_72609_ _79267_/B _72590_/X _72606_/X _72608_/Y _83218_/D sky130_fd_sc_hd__o22a_4
X_79165_ _58946_/Y _79165_/B _79165_/Y sky130_fd_sc_hd__nand2_4
X_45557_ _56627_/B _45556_/X _45378_/X _45557_/X sky130_fd_sc_hd__o21a_4
X_64391_ _64274_/A _64391_/X sky130_fd_sc_hd__buf_2
X_76377_ _81650_/Q _76377_/Y sky130_fd_sc_hd__inv_2
X_42769_ _41302_/X _42767_/X _67406_/B _42768_/X _87728_/D sky130_fd_sc_hd__a2bb2o_4
X_73589_ _73566_/X _84992_/Q _73385_/X _73588_/X _73589_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_opt_7_CLK _83248_/CLK _84837_/CLK sky130_fd_sc_hd__clkbuf_16
X_66130_ _66053_/X _85618_/Q _66096_/X _66129_/X _66130_/X sky130_fd_sc_hd__a211o_4
X_78116_ _78109_/Y _78114_/Y _78115_/Y _78120_/C sky130_fd_sc_hd__a21o_4
X_44508_ _44496_/X _44497_/X _41276_/X _87073_/Q _44498_/X _44509_/A
+ sky130_fd_sc_hd__o32ai_4
X_63342_ _60433_/A _63342_/B _63342_/C _60484_/A _63342_/X sky130_fd_sc_hd__and4_4
X_75328_ _75325_/Y _75328_/B _75328_/X sky130_fd_sc_hd__xor2_4
X_60554_ _60443_/A _60588_/A _60607_/A _60555_/A sky130_fd_sc_hd__nor3_4
X_48276_ _48020_/B _50322_/B sky130_fd_sc_hd__buf_2
X_79096_ _79095_/B _79095_/A _79109_/A sky130_fd_sc_hd__nand2_4
X_45488_ _57392_/B _45488_/Y sky130_fd_sc_hd__inv_2
X_47227_ _47227_/A _52927_/D sky130_fd_sc_hd__buf_2
X_66061_ _66061_/A _66061_/B _66061_/Y sky130_fd_sc_hd__nand2_4
X_78047_ _78046_/Y _78047_/Y sky130_fd_sc_hd__inv_2
X_44439_ _44425_/X _44427_/X _41606_/X _87107_/Q _44428_/X _44439_/Y
+ sky130_fd_sc_hd__o32ai_4
X_63273_ _84842_/Q _63281_/B _63301_/C _63281_/D _63273_/X sky130_fd_sc_hd__or4_4
X_75259_ _75258_/B _75258_/C _75254_/Y _75259_/Y sky130_fd_sc_hd__o21ai_4
X_60485_ _63280_/C _60488_/C sky130_fd_sc_hd__buf_2
X_65012_ _65012_/A _65012_/B _65012_/X sky130_fd_sc_hd__and2_4
X_62224_ _62501_/A _62631_/C sky130_fd_sc_hd__buf_2
X_47158_ _54578_/B _52885_/B sky130_fd_sc_hd__buf_2
X_46109_ _46109_/A _46108_/X _46109_/Y sky130_fd_sc_hd__nand2_4
X_69820_ _87808_/Q _69820_/Y sky130_fd_sc_hd__inv_2
X_62155_ _62144_/A _62121_/X _78052_/B _62155_/Y sky130_fd_sc_hd__nor3_4
X_47089_ _47063_/A _52850_/B _47089_/Y sky130_fd_sc_hd__nand2_4
X_79998_ _79998_/A _79998_/B _80003_/B sky130_fd_sc_hd__xor2_4
X_61106_ _84520_/Q _60979_/X _61104_/Y _61105_/X _61106_/Y sky130_fd_sc_hd__a2bb2oi_4
X_69751_ _69751_/A _69751_/X sky130_fd_sc_hd__buf_2
X_66963_ _87427_/Q _66915_/X _66863_/X _66962_/X _66963_/X sky130_fd_sc_hd__a211o_4
X_62086_ _84890_/Q _62128_/B _62128_/C _62060_/X _62086_/Y sky130_fd_sc_hd__nand4_4
X_78949_ _82818_/Q _78949_/B _79115_/A sky130_fd_sc_hd__xnor2_4
X_68702_ _68599_/A _87750_/Q _68702_/X sky130_fd_sc_hd__and2_4
X_65914_ _65903_/X _65431_/Y _65913_/Y _65914_/Y sky130_fd_sc_hd__o21ai_4
X_61037_ _61037_/A _61037_/Y sky130_fd_sc_hd__inv_2
X_81960_ _82339_/CLK _83888_/Q _81960_/Q sky130_fd_sc_hd__dfxtp_4
X_69682_ _69679_/X _69681_/X _69655_/X _69682_/Y sky130_fd_sc_hd__a21oi_4
X_66894_ _66891_/X _66893_/X _66871_/X _66894_/Y sky130_fd_sc_hd__a21oi_4
X_80911_ _83918_/CLK _80911_/D _75687_/A sky130_fd_sc_hd__dfxtp_4
X_68633_ _68629_/X _68632_/X _68512_/X _68633_/Y sky130_fd_sc_hd__a21oi_4
X_65845_ _64752_/A _65845_/X sky130_fd_sc_hd__buf_2
X_81891_ _82145_/CLK _81891_/D _82299_/D sky130_fd_sc_hd__dfxtp_4
X_52810_ _52757_/A _52818_/A sky130_fd_sc_hd__buf_2
X_83630_ _83630_/CLK _71031_/Y _47631_/A sky130_fd_sc_hd__dfxtp_4
X_80842_ _80754_/CLK _80874_/Q _80842_/Q sky130_fd_sc_hd__dfxtp_4
X_68564_ _80826_/D _68462_/X _68563_/X _83970_/D sky130_fd_sc_hd__a21bo_4
X_53790_ _53787_/Y _53773_/X _53789_/X _53790_/Y sky130_fd_sc_hd__a21oi_4
X_65776_ _65772_/Y _65757_/X _65775_/X _84179_/D sky130_fd_sc_hd__a21o_4
X_62988_ _62988_/A _62988_/B _62988_/C _62988_/Y sky130_fd_sc_hd__nor3_4
X_67515_ _67510_/X _67514_/X _67442_/X _67515_/X sky130_fd_sc_hd__a21o_4
X_52741_ _52770_/A _52746_/B sky130_fd_sc_hd__buf_2
X_64727_ _64722_/X _85565_/Q _64724_/X _64726_/X _64727_/X sky130_fd_sc_hd__a211o_4
X_83561_ _83561_/CLK _71244_/Y _83561_/Q sky130_fd_sc_hd__dfxtp_4
X_61939_ _58329_/A _61939_/X sky130_fd_sc_hd__buf_2
X_80773_ _81990_/CLK _80773_/D _80773_/Q sky130_fd_sc_hd__dfxtp_4
X_68495_ _69001_/A _68495_/B _68495_/Y sky130_fd_sc_hd__nor2_4
X_85300_ _85270_/CLK _85300_/D _55870_/B sky130_fd_sc_hd__dfxtp_4
X_82512_ _82580_/CLK _82512_/D _82512_/Q sky130_fd_sc_hd__dfxtp_4
X_55460_ _45600_/A _55453_/X _55458_/X _55459_/Y _55460_/X sky130_fd_sc_hd__a211o_4
X_67446_ _67443_/X _67445_/X _67401_/X _67446_/Y sky130_fd_sc_hd__a21oi_4
X_86280_ _86600_/CLK _86280_/D _72415_/B sky130_fd_sc_hd__dfxtp_4
X_52672_ _85775_/Q _52656_/X _52671_/Y _52672_/Y sky130_fd_sc_hd__o21ai_4
X_64658_ _64684_/A _64658_/B _64658_/X sky130_fd_sc_hd__and2_4
X_83492_ _83495_/CLK _71457_/X _83492_/Q sky130_fd_sc_hd__dfxtp_4
X_54411_ _85447_/Q _54404_/X _54410_/Y _54411_/Y sky130_fd_sc_hd__o21ai_4
X_85231_ _85167_/CLK _56336_/Y _55821_/B sky130_fd_sc_hd__dfxtp_4
X_51623_ _51627_/A _53148_/B _51623_/Y sky130_fd_sc_hd__nand2_4
X_63609_ _63487_/A _63609_/X sky130_fd_sc_hd__buf_2
X_82443_ _82443_/CLK _79135_/X _82411_/D sky130_fd_sc_hd__dfxtp_4
X_55391_ _55380_/Y _55389_/Y _55441_/C _55393_/B sky130_fd_sc_hd__o21a_4
X_67377_ _81504_/D _67331_/X _67376_/X _84072_/D sky130_fd_sc_hd__a21bo_4
X_64589_ _64678_/A _64589_/X sky130_fd_sc_hd__buf_2
X_57130_ _56700_/Y _56808_/A _56816_/A _57129_/Y _57133_/A sky130_fd_sc_hd__and4_4
X_69116_ _64806_/A _69116_/X sky130_fd_sc_hd__buf_2
X_54342_ _85459_/Q _54320_/X _54341_/Y _54342_/Y sky130_fd_sc_hd__o21ai_4
X_66328_ _66325_/X _66328_/B _66328_/Y sky130_fd_sc_hd__nand2_4
X_85162_ _80671_/CLK _85162_/D _85162_/Q sky130_fd_sc_hd__dfxtp_4
X_51554_ _51551_/Y _51531_/X _51553_/X _85989_/D sky130_fd_sc_hd__a21oi_4
X_82374_ _86655_/CLK _82374_/D _82374_/Q sky130_fd_sc_hd__dfxtp_4
X_84113_ _84111_/CLK _84113_/D _66490_/C sky130_fd_sc_hd__dfxtp_4
X_50505_ _50505_/A _50506_/A sky130_fd_sc_hd__buf_2
X_57061_ _56850_/X _56976_/X _57055_/A _57061_/Y sky130_fd_sc_hd__o21ai_4
X_81325_ _81431_/CLK _76312_/X _81701_/D sky130_fd_sc_hd__dfxtp_4
X_69047_ _69043_/X _69046_/X _69025_/X _69047_/X sky130_fd_sc_hd__a21o_4
X_54273_ _85472_/Q _54266_/X _54272_/Y _54273_/Y sky130_fd_sc_hd__o21ai_4
X_66259_ _66104_/A _66276_/B sky130_fd_sc_hd__buf_2
X_85093_ _85128_/CLK _85093_/D _57071_/B sky130_fd_sc_hd__dfxtp_4
X_51485_ _51539_/A _51485_/X sky130_fd_sc_hd__buf_2
X_56012_ _56054_/B _55928_/C _55927_/X _55956_/B _56030_/B sky130_fd_sc_hd__nand4_4
X_53224_ _53220_/Y _53215_/X _53223_/X _53224_/Y sky130_fd_sc_hd__a21oi_4
X_84044_ _88116_/CLK _84044_/D _84044_/Q sky130_fd_sc_hd__dfxtp_4
X_50436_ _50433_/Y _50429_/X _50435_/X _86201_/D sky130_fd_sc_hd__a21oi_4
X_81256_ _81288_/CLK _81256_/D _81256_/Q sky130_fd_sc_hd__dfxtp_4
X_80207_ _80205_/X _80207_/B _80207_/Y sky130_fd_sc_hd__xnor2_4
X_53155_ _53139_/A _53159_/B _53143_/X _53155_/D _53155_/X sky130_fd_sc_hd__and4_4
X_50367_ _50572_/A _50381_/A sky130_fd_sc_hd__buf_2
X_81187_ _80821_/CLK _74906_/X _49190_/A sky130_fd_sc_hd__dfxtp_4
X_52106_ _65451_/B _52089_/X _52105_/Y _52106_/Y sky130_fd_sc_hd__o21ai_4
X_87803_ _87813_/CLK _42607_/Y _69882_/A sky130_fd_sc_hd__dfxtp_4
X_80138_ _80122_/X _80125_/Y _80137_/X _80138_/X sky130_fd_sc_hd__a21o_4
X_53086_ _53080_/A _53086_/B _53086_/Y sky130_fd_sc_hd__nand2_4
X_57963_ _57903_/X _85488_/Q _57962_/X _57963_/X sky130_fd_sc_hd__o21a_4
X_69949_ _69900_/A _88310_/Q _69949_/X sky130_fd_sc_hd__and2_4
X_50298_ _86228_/Q _50282_/X _50297_/Y _50298_/Y sky130_fd_sc_hd__o21ai_4
X_85995_ _85709_/CLK _51523_/Y _85995_/Q sky130_fd_sc_hd__dfxtp_4
X_59702_ _59696_/A _59711_/B _80588_/A _59702_/Y sky130_fd_sc_hd__nor3_4
X_52037_ _85901_/Q _52013_/X _52036_/Y _52037_/Y sky130_fd_sc_hd__o21ai_4
X_56914_ _56985_/D _57319_/D _56914_/Y sky130_fd_sc_hd__nor2_4
X_87734_ _87990_/CLK _87734_/D _69076_/B sky130_fd_sc_hd__dfxtp_4
X_72960_ _73093_/A _72960_/B _72960_/X sky130_fd_sc_hd__and2_4
X_84946_ _84945_/CLK _84946_/D _84946_/Q sky130_fd_sc_hd__dfxtp_4
X_80069_ _60089_/C _64022_/C _80069_/X sky130_fd_sc_hd__xor2_4
X_57894_ _57781_/X _57891_/Y _57892_/Y _57893_/X _57795_/X _57894_/X
+ sky130_fd_sc_hd__o32a_4
X_71911_ _56878_/Y _71891_/Y _71910_/Y _83331_/D sky130_fd_sc_hd__o21ai_4
X_59633_ _59633_/A _59634_/A sky130_fd_sc_hd__inv_2
X_56845_ _46233_/Y _55680_/B _56845_/Y sky130_fd_sc_hd__nor2_4
X_87665_ _81783_/CLK _87665_/D _67378_/B sky130_fd_sc_hd__dfxtp_4
X_72891_ _44270_/X _72892_/B sky130_fd_sc_hd__buf_2
X_84877_ _84877_/CLK _84877_/D _84877_/Q sky130_fd_sc_hd__dfxtp_4
X_43810_ _43810_/A _43810_/X sky130_fd_sc_hd__buf_2
X_74630_ _74694_/A _74630_/X sky130_fd_sc_hd__buf_2
X_86616_ _85974_/CLK _86616_/D _86616_/Q sky130_fd_sc_hd__dfxtp_4
X_71842_ _71824_/Y _83355_/Q _71841_/X _83355_/D sky130_fd_sc_hd__a21o_4
X_59564_ _59564_/A _59564_/B _59890_/C _59752_/A sky130_fd_sc_hd__nand3_4
X_83828_ _83188_/CLK _70235_/X _83828_/Q sky130_fd_sc_hd__dfxtp_4
X_44790_ _41397_/A _44788_/X _86954_/Q _44789_/X _86954_/D sky130_fd_sc_hd__a2bb2o_4
X_56776_ _83325_/Q _56776_/B _56776_/X sky130_fd_sc_hd__xor2_4
X_87596_ _87045_/CLK _87596_/D _43043_/A sky130_fd_sc_hd__dfxtp_4
X_53988_ _53986_/Y _53982_/X _53987_/Y _85528_/D sky130_fd_sc_hd__a21boi_4
X_58515_ _63496_/B _58510_/X _58515_/Y sky130_fd_sc_hd__nor2_4
X_43741_ _87288_/Q _43741_/Y sky130_fd_sc_hd__inv_2
X_74561_ _45007_/A _74551_/X _74560_/X _83035_/D sky130_fd_sc_hd__o21ai_4
X_55727_ _55719_/Y _55721_/Y _55726_/Y _56163_/A sky130_fd_sc_hd__a21oi_4
X_86547_ _86549_/CLK _48258_/Y _66119_/B sky130_fd_sc_hd__dfxtp_4
X_40953_ _82302_/Q _40932_/X _40953_/X sky130_fd_sc_hd__or2_4
X_52939_ _52937_/Y _52920_/X _52938_/X _52939_/Y sky130_fd_sc_hd__a21oi_4
X_83759_ _84945_/CLK _83759_/D _83759_/Q sky130_fd_sc_hd__dfxtp_4
X_71773_ _71762_/X _83381_/Q _71772_/X _71773_/X sky130_fd_sc_hd__a21o_4
X_59495_ _46179_/X _63410_/B _59494_/Y _84717_/D sky130_fd_sc_hd__o21a_4
Xclkbuf_4_9_1_CLK clkbuf_4_9_0_CLK/X clkbuf_4_9_1_CLK/X sky130_fd_sc_hd__clkbuf_1
X_76300_ _76300_/A _76300_/Y sky130_fd_sc_hd__inv_2
X_73512_ _69961_/B _73026_/X _73421_/X _73512_/Y sky130_fd_sc_hd__o21ai_4
X_46460_ _46403_/X _81199_/Q _46459_/X _51326_/B sky130_fd_sc_hd__o21ai_4
X_70724_ _70724_/A _70713_/X _70727_/C _70769_/D _70724_/Y sky130_fd_sc_hd__nand4_4
X_58446_ _58446_/A _58426_/X _58446_/Y sky130_fd_sc_hd__nand2_4
X_77280_ _77278_/X _77279_/Y _82214_/Q _77280_/X sky130_fd_sc_hd__a21o_4
X_43672_ _43606_/A _43673_/A sky130_fd_sc_hd__buf_2
X_55658_ _83315_/Q _83314_/Q _55658_/Y sky130_fd_sc_hd__nor2_4
X_74492_ _74492_/A _74492_/X sky130_fd_sc_hd__buf_2
X_86478_ _86506_/CLK _48815_/Y _86478_/Q sky130_fd_sc_hd__dfxtp_4
X_40884_ _40857_/X _41057_/A _40883_/X _40885_/A sky130_fd_sc_hd__o21a_4
X_45411_ _85024_/Q _55628_/B sky130_fd_sc_hd__inv_2
X_76231_ _76232_/A _76229_/Y _76230_/Y _76231_/Y sky130_fd_sc_hd__o21ai_4
X_88217_ _88215_/CLK _41430_/X _88217_/Q sky130_fd_sc_hd__dfxtp_4
X_42623_ _49210_/B _42569_/X _40925_/X _69958_/B _42612_/X _87797_/D
+ sky130_fd_sc_hd__o32ai_4
X_54609_ _54600_/A _47212_/Y _54609_/Y sky130_fd_sc_hd__nand2_4
X_73443_ _69923_/B _72865_/X _72866_/X _73443_/X sky130_fd_sc_hd__o21a_4
X_85429_ _83046_/CLK _54510_/Y _85429_/Q sky130_fd_sc_hd__dfxtp_4
X_46391_ _46391_/A _52482_/B sky130_fd_sc_hd__buf_2
X_70655_ _70925_/A _70890_/C sky130_fd_sc_hd__buf_2
X_58377_ _58377_/A _58369_/X _58377_/Y sky130_fd_sc_hd__nand2_4
X_55589_ _55843_/A _55908_/A sky130_fd_sc_hd__buf_2
XPHY_60 sky130_fd_sc_hd__decap_3
X_48130_ _48130_/A _57637_/B sky130_fd_sc_hd__inv_2
X_45342_ _45338_/Y _45341_/Y _45287_/X _45342_/X sky130_fd_sc_hd__a21o_4
XPHY_71 sky130_fd_sc_hd__decap_3
X_57328_ _57328_/A _57328_/Y sky130_fd_sc_hd__inv_2
X_88148_ _88208_/CLK _41794_/Y _88148_/Q sky130_fd_sc_hd__dfxtp_4
X_76162_ _76155_/A _76155_/B _76162_/Y sky130_fd_sc_hd__nor2_4
X_42554_ _42554_/A _42554_/X sky130_fd_sc_hd__buf_2
X_73374_ _73374_/A _73372_/B _73374_/Y sky130_fd_sc_hd__nor2_4
XPHY_82 sky130_fd_sc_hd__decap_3
X_70586_ _70576_/X _70586_/X sky130_fd_sc_hd__buf_2
XPHY_93 sky130_fd_sc_hd__decap_3
X_75113_ _75113_/A _81061_/Q _75113_/C _75117_/C sky130_fd_sc_hd__nand3_4
X_41505_ _81176_/Q _41523_/B _41505_/X sky130_fd_sc_hd__or2_4
X_48061_ _53567_/B _52047_/B sky130_fd_sc_hd__buf_2
X_72325_ _72287_/X _85328_/Q _72324_/X _72325_/X sky130_fd_sc_hd__o21a_4
X_45273_ _45273_/A _45272_/X _45273_/Y sky130_fd_sc_hd__nand2_4
X_57259_ _57243_/X _56630_/X _45567_/A _57245_/X _57259_/X sky130_fd_sc_hd__a2bb2o_4
X_76093_ _76093_/A _76093_/Y sky130_fd_sc_hd__inv_2
X_88079_ _87288_/CLK _41991_/Y _72855_/A sky130_fd_sc_hd__dfxtp_4
X_42485_ _42465_/A _42554_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_452_0_CLK clkbuf_9_226_0_CLK/X _84922_/CLK sky130_fd_sc_hd__clkbuf_1
X_47012_ _54494_/D _52801_/D sky130_fd_sc_hd__buf_2
X_44224_ _66608_/A _44225_/B sky130_fd_sc_hd__buf_2
X_75044_ _75041_/Y _75043_/Y _75045_/B sky130_fd_sc_hd__xor2_4
X_79921_ _79921_/A _79922_/A sky130_fd_sc_hd__inv_2
X_41436_ _41412_/X _82885_/Q _41435_/X _41436_/Y sky130_fd_sc_hd__o21ai_4
X_72256_ _72196_/X _85334_/Q _72255_/X _72256_/X sky130_fd_sc_hd__o21a_4
X_60270_ _60156_/Y _60204_/A _60271_/A sky130_fd_sc_hd__and2_4
X_71207_ _71211_/A _71230_/B _71197_/C _71207_/Y sky130_fd_sc_hd__nand3_4
X_44155_ _66563_/A _66180_/A sky130_fd_sc_hd__buf_2
X_79852_ _79851_/Y _79852_/B _79852_/X sky130_fd_sc_hd__and2_4
X_41367_ _41366_/Y _41367_/X sky130_fd_sc_hd__buf_2
X_72187_ _72220_/A _72187_/B _72187_/Y sky130_fd_sc_hd__nor2_4
X_43106_ _43189_/A _43106_/X sky130_fd_sc_hd__buf_2
X_78803_ _82834_/Q _82546_/Q _78804_/B sky130_fd_sc_hd__xnor2_4
X_71138_ _71138_/A _71138_/X sky130_fd_sc_hd__buf_2
X_48963_ _71996_/B _48963_/X sky130_fd_sc_hd__buf_2
X_44086_ _44086_/A _44087_/B sky130_fd_sc_hd__buf_2
X_79783_ _84224_/Q _72224_/A _79794_/A sky130_fd_sc_hd__xor2_4
X_41298_ _41298_/A _41298_/X sky130_fd_sc_hd__buf_2
X_76995_ _60970_/C _76995_/B _76995_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_10_467_0_CLK clkbuf_9_233_0_CLK/X _83663_/CLK sky130_fd_sc_hd__clkbuf_1
X_47914_ _82362_/Q _48438_/B sky130_fd_sc_hd__inv_2
X_43037_ _43036_/Y _87599_/D sky130_fd_sc_hd__inv_2
X_78734_ _78709_/Y _78713_/B _78712_/A _78735_/A sky130_fd_sc_hd__o21a_4
X_75946_ _81701_/D _75940_/B _75946_/Y sky130_fd_sc_hd__nor2_4
X_63960_ _63960_/A _63960_/B _80111_/B _63960_/Y sky130_fd_sc_hd__nor3_4
X_71069_ _71069_/A _71070_/A sky130_fd_sc_hd__buf_2
X_48894_ _48894_/A _48894_/B _48894_/C _48894_/X sky130_fd_sc_hd__and3_4
X_62911_ _62967_/A _58459_/Y _62911_/C _62967_/D _62911_/X sky130_fd_sc_hd__and4_4
X_47845_ _65921_/B _47840_/X _47844_/Y _47845_/Y sky130_fd_sc_hd__o21ai_4
X_78665_ _78645_/Y _78649_/B _78648_/A _78665_/X sky130_fd_sc_hd__o21a_4
X_63891_ _60984_/A _63892_/D sky130_fd_sc_hd__buf_2
X_75877_ _81025_/Q _75878_/B sky130_fd_sc_hd__inv_2
X_65630_ _65524_/X _83068_/Q _65568_/X _65629_/X _65630_/X sky130_fd_sc_hd__a211o_4
X_77616_ _77603_/A _77600_/Y _77601_/Y _77616_/X sky130_fd_sc_hd__o21a_4
X_62842_ _63557_/B _62841_/X _60309_/C _60254_/B _62842_/Y sky130_fd_sc_hd__nand4_4
X_74828_ _74828_/A _74828_/Y sky130_fd_sc_hd__inv_2
X_47776_ _47776_/A _53238_/D sky130_fd_sc_hd__buf_2
X_78596_ _82806_/Q _78596_/Y sky130_fd_sc_hd__inv_2
X_44988_ _55943_/B _44963_/X _44964_/X _44988_/X sky130_fd_sc_hd__o21a_4
X_49515_ _49407_/A _49537_/A sky130_fd_sc_hd__buf_2
X_46727_ _46727_/A _46727_/Y sky130_fd_sc_hd__inv_2
X_65561_ _65777_/A _85880_/Q _65561_/X sky130_fd_sc_hd__and2_4
X_77547_ _77547_/A _77547_/B _82199_/D sky130_fd_sc_hd__xor2_4
X_43939_ _43927_/X _43939_/X sky130_fd_sc_hd__buf_2
X_62773_ _60362_/A _62773_/X sky130_fd_sc_hd__buf_2
X_74759_ _70735_/X _74780_/D sky130_fd_sc_hd__buf_2
Xclkbuf_9_511_0_CLK clkbuf_9_510_0_CLK/A clkbuf_9_511_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_67300_ _67324_/A _88181_/Q _67300_/X sky130_fd_sc_hd__and2_4
X_64512_ _64363_/A _64363_/B _84910_/Q _61145_/X _64512_/X sky130_fd_sc_hd__and4_4
X_49446_ _58763_/B _49443_/X _49445_/Y _49446_/Y sky130_fd_sc_hd__o21ai_4
X_61724_ _61752_/A _61723_/X _78080_/B _61724_/Y sky130_fd_sc_hd__nor3_4
X_68280_ _67731_/X _67733_/X _68239_/X _68280_/Y sky130_fd_sc_hd__a21oi_4
X_46658_ _46658_/A _51772_/D sky130_fd_sc_hd__buf_2
X_65492_ _65474_/X _86525_/Q _65492_/X sky130_fd_sc_hd__and2_4
X_77478_ _77478_/A _77478_/B _77477_/Y _77478_/X sky130_fd_sc_hd__or3_4
Xclkbuf_10_405_0_CLK clkbuf_9_202_0_CLK/X _85375_/CLK sky130_fd_sc_hd__clkbuf_1
X_67231_ _67183_/A _67231_/B _67231_/X sky130_fd_sc_hd__and2_4
X_79217_ _79213_/Y _79215_/X _79236_/A _79217_/Y sky130_fd_sc_hd__nand3_4
X_45609_ _45591_/X _61492_/A _45608_/X _45609_/Y sky130_fd_sc_hd__o21ai_4
X_64443_ _64431_/Y _64441_/X _64442_/X _64443_/X sky130_fd_sc_hd__o21a_4
X_76429_ _76429_/A _76430_/C sky130_fd_sc_hd__inv_2
X_49377_ _86398_/Q _49360_/X _49376_/Y _49377_/Y sky130_fd_sc_hd__o21ai_4
X_61655_ _61655_/A _61653_/X _61654_/X _61639_/X _61655_/Y sky130_fd_sc_hd__nand4_4
X_46589_ _82915_/Q _46579_/X _46589_/X sky130_fd_sc_hd__or2_4
X_48328_ _66301_/B _48293_/X _48327_/Y _48328_/Y sky130_fd_sc_hd__o21ai_4
X_60606_ _60606_/A _60606_/X sky130_fd_sc_hd__buf_2
X_67162_ _87111_/Q _67110_/X _67160_/X _67161_/X _67162_/X sky130_fd_sc_hd__a211o_4
X_79148_ _79148_/A _79148_/B _82456_/D sky130_fd_sc_hd__xor2_4
X_64374_ _64315_/A _64418_/B sky130_fd_sc_hd__buf_2
X_61586_ _61579_/Y _61581_/Y _61582_/Y _61583_/Y _61585_/Y _61586_/Y
+ sky130_fd_sc_hd__a41oi_4
X_66113_ _72155_/A _86227_/Q _64692_/X _66112_/X _66113_/X sky130_fd_sc_hd__a211o_4
X_63325_ _63321_/Y _63322_/X _63323_/X _63324_/X _63242_/X _63325_/Y
+ sky130_fd_sc_hd__o41ai_4
X_48259_ _48190_/A _50306_/B _48259_/Y sky130_fd_sc_hd__nand2_4
X_60537_ _60536_/X _60537_/Y sky130_fd_sc_hd__inv_2
X_67093_ _66565_/A _67093_/X sky130_fd_sc_hd__buf_2
X_79079_ _79075_/Y _79078_/Y _79080_/A sky130_fd_sc_hd__xor2_4
X_81110_ _80708_/CLK _79771_/X _81110_/Q sky130_fd_sc_hd__dfxtp_4
X_66044_ _66044_/A _66062_/B _65570_/X _66044_/Y sky130_fd_sc_hd__nand3_4
X_51270_ _51278_/A _46330_/A _51270_/X sky130_fd_sc_hd__and2_4
X_63256_ _63285_/A _63285_/B _79288_/A _63256_/Y sky130_fd_sc_hd__nor3_4
X_82090_ _82009_/CLK _77338_/B _77060_/A sky130_fd_sc_hd__dfxtp_4
X_60468_ _60399_/B _60570_/B sky130_fd_sc_hd__buf_2
X_50221_ _50221_/A _51074_/A sky130_fd_sc_hd__buf_2
X_62207_ _59896_/X _62560_/B sky130_fd_sc_hd__buf_2
X_81041_ _81041_/CLK _81041_/D _81041_/Q sky130_fd_sc_hd__dfxtp_4
X_63187_ _84346_/Q _63130_/X _63186_/Y _84346_/D sky130_fd_sc_hd__a21o_4
X_60399_ _60515_/C _60399_/B _60570_/A _60399_/Y sky130_fd_sc_hd__nor3_4
X_69803_ _81968_/D _69763_/X _69802_/X _83896_/D sky130_fd_sc_hd__a21bo_4
X_50152_ _50150_/Y _50141_/X _50151_/X _50152_/Y sky130_fd_sc_hd__a21oi_4
X_62138_ _61652_/B _62149_/B _62149_/C _61749_/B _62138_/Y sky130_fd_sc_hd__nand4_4
X_67995_ _67948_/X _67981_/Y _67983_/X _67994_/Y _67995_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_8_94_0_CLK clkbuf_8_95_0_CLK/A clkbuf_8_94_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_84800_ _86713_/CLK _84800_/D _84800_/Q sky130_fd_sc_hd__dfxtp_4
X_69734_ _69734_/A _69734_/Y sky130_fd_sc_hd__inv_2
X_50083_ _50081_/Y _50068_/X _50082_/X _50083_/Y sky130_fd_sc_hd__a21oi_4
X_54960_ _54958_/Y _54253_/X _54959_/X _85345_/D sky130_fd_sc_hd__a21oi_4
X_66946_ _80914_/D _66850_/X _66945_/X _66946_/X sky130_fd_sc_hd__a21bo_4
X_62069_ _62067_/Y _62033_/X _62068_/Y _62069_/Y sky130_fd_sc_hd__a21oi_4
X_85780_ _82956_/CLK _52650_/Y _85780_/Q sky130_fd_sc_hd__dfxtp_4
X_82992_ _85039_/CLK _74664_/Y _82992_/Q sky130_fd_sc_hd__dfxtp_4
X_53911_ _53909_/Y _53862_/X _53910_/Y _85544_/D sky130_fd_sc_hd__a21boi_4
X_84731_ _84732_/CLK _84731_/D _59443_/A sky130_fd_sc_hd__dfxtp_4
X_81943_ _82133_/CLK _81943_/D _81943_/Q sky130_fd_sc_hd__dfxtp_4
X_69665_ _69797_/A _69665_/X sky130_fd_sc_hd__buf_2
X_54891_ _54886_/Y _54882_/X _54890_/X _54891_/Y sky130_fd_sc_hd__a21oi_4
X_66877_ _87942_/Q _66875_/X _66807_/X _66876_/X _66877_/X sky130_fd_sc_hd__a211o_4
X_56630_ _56630_/A _56630_/X sky130_fd_sc_hd__buf_2
X_68616_ _87593_/Q _68463_/X _68613_/X _68615_/X _68616_/X sky130_fd_sc_hd__a211o_4
X_87450_ _87446_/CLK _87450_/D _87450_/Q sky130_fd_sc_hd__dfxtp_4
X_53842_ _85557_/Q _53816_/X _53841_/Y _53842_/Y sky130_fd_sc_hd__o21ai_4
X_65828_ _65288_/X _65828_/B _65290_/X _65828_/Y sky130_fd_sc_hd__nand3_4
X_84662_ _84660_/CLK _84662_/D _60097_/C sky130_fd_sc_hd__dfxtp_4
X_81874_ _81857_/CLK _78065_/X _81842_/D sky130_fd_sc_hd__dfxtp_4
X_69596_ _69593_/X _69595_/X _69570_/X _69596_/X sky130_fd_sc_hd__a21o_4
X_86401_ _84815_/CLK _49365_/Y _86401_/Q sky130_fd_sc_hd__dfxtp_4
X_83613_ _83613_/CLK _71083_/Y _49005_/A sky130_fd_sc_hd__dfxtp_4
X_56561_ _56560_/X _56561_/X sky130_fd_sc_hd__buf_2
X_68547_ _87500_/Q _68472_/A _68545_/X _68546_/X _68547_/X sky130_fd_sc_hd__a211o_4
X_80825_ _80931_/CLK _80825_/D _80825_/Q sky130_fd_sc_hd__dfxtp_4
X_87381_ _86914_/CLK _87381_/D _87381_/Q sky130_fd_sc_hd__dfxtp_4
X_53773_ _53773_/A _53773_/X sky130_fd_sc_hd__buf_2
X_65759_ _65756_/Y _65757_/X _65758_/X _84180_/D sky130_fd_sc_hd__a21o_4
X_84593_ _82452_/CLK _60587_/Y _79133_/A sky130_fd_sc_hd__dfxtp_4
X_50985_ _50973_/X _50985_/B _50985_/C _46791_/X _50985_/X sky130_fd_sc_hd__and4_4
X_58300_ _58510_/A _58344_/B sky130_fd_sc_hd__buf_2
X_55512_ _55458_/X _55512_/X sky130_fd_sc_hd__buf_2
X_86332_ _86651_/CLK _86332_/D _86332_/Q sky130_fd_sc_hd__dfxtp_4
X_52724_ _52704_/A _52724_/B _52708_/X _52724_/D _52724_/X sky130_fd_sc_hd__and4_4
X_59280_ _84755_/Q _59268_/X _59272_/X _59279_/X _84755_/D sky130_fd_sc_hd__a2bb2oi_4
X_83544_ _83544_/CLK _83544_/D _83544_/Q sky130_fd_sc_hd__dfxtp_4
X_56492_ _56487_/X _56484_/X _55896_/B _56492_/Y sky130_fd_sc_hd__nand3_4
X_80756_ _80804_/CLK _80756_/D _81132_/D sky130_fd_sc_hd__dfxtp_4
X_68478_ _68471_/X _68476_/X _68477_/X _68478_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_8_32_0_CLK clkbuf_7_16_0_CLK/X clkbuf_9_65_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_58231_ _46179_/X _58228_/X _58230_/Y _84902_/D sky130_fd_sc_hd__o21a_4
X_55443_ _55443_/A _55442_/Y _55443_/C _55443_/D _55443_/Y sky130_fd_sc_hd__nand4_4
X_67429_ _67381_/A _67429_/B _67429_/X sky130_fd_sc_hd__and2_4
X_86263_ _83305_/CLK _86263_/D _86263_/Q sky130_fd_sc_hd__dfxtp_4
X_52655_ _52652_/Y _52647_/X _52654_/X _85779_/D sky130_fd_sc_hd__a21oi_4
X_83475_ _83763_/CLK _71503_/X _83475_/Q sky130_fd_sc_hd__dfxtp_4
X_80687_ _80719_/CLK _80687_/D _75255_/A sky130_fd_sc_hd__dfxtp_4
XPHY_603 sky130_fd_sc_hd__decap_3
X_88002_ _88002_/CLK _88002_/D _88002_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_614 sky130_fd_sc_hd__decap_3
X_85214_ _83001_/CLK _56387_/Y _56386_/C sky130_fd_sc_hd__dfxtp_4
X_51606_ _85979_/Q _51594_/X _51605_/Y _51606_/Y sky130_fd_sc_hd__o21ai_4
X_70440_ _70997_/A _70949_/B sky130_fd_sc_hd__buf_2
X_58162_ _58162_/A _63054_/A sky130_fd_sc_hd__inv_2
XPHY_625 sky130_fd_sc_hd__decap_3
X_82426_ _82833_/CLK _82458_/Q _78661_/A sky130_fd_sc_hd__dfxtp_4
X_55374_ _55373_/Y _55298_/X _55201_/Y _55374_/Y sky130_fd_sc_hd__a21oi_4
X_86194_ _83313_/CLK _50476_/Y _86194_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_636 sky130_fd_sc_hd__decap_3
X_52586_ _52590_/A _54277_/B _52586_/Y sky130_fd_sc_hd__nand2_4
XPHY_647 sky130_fd_sc_hd__decap_3
XPHY_658 sky130_fd_sc_hd__decap_3
X_57113_ _56960_/X _57113_/B _57112_/X _57113_/Y sky130_fd_sc_hd__nor3_4
X_54325_ _54325_/A _54325_/B _54317_/X _54325_/D _54325_/X sky130_fd_sc_hd__and4_4
XPHY_669 sky130_fd_sc_hd__decap_3
X_85145_ _85057_/CLK _85145_/D _56614_/B sky130_fd_sc_hd__dfxtp_4
X_51537_ _51521_/X _51553_/B _51533_/C _53063_/D _51537_/X sky130_fd_sc_hd__and4_4
X_70371_ _70366_/X _70368_/X _70375_/C _70371_/Y sky130_fd_sc_hd__nand3_4
X_58093_ _84926_/Q _58025_/X _58084_/X _58092_/X _84926_/D sky130_fd_sc_hd__a2bb2oi_4
X_82357_ _84981_/CLK _77191_/X _47963_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_47_0_CLK clkbuf_8_47_0_CLK/A clkbuf_9_94_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_72110_ _72068_/A _53936_/B _72110_/Y sky130_fd_sc_hd__nand2_4
X_81308_ _81632_/CLK _76996_/X _81276_/D sky130_fd_sc_hd__dfxtp_4
X_57044_ _56930_/X _57040_/Y _57043_/Y _57044_/Y sky130_fd_sc_hd__o21ai_4
X_42270_ _41503_/X _42258_/X _87947_/Q _42259_/X _87947_/D sky130_fd_sc_hd__a2bb2o_4
X_54256_ _54252_/Y _54253_/X _54255_/X _54256_/Y sky130_fd_sc_hd__a21oi_4
X_73090_ _73132_/A _85877_/Q _73090_/X sky130_fd_sc_hd__and2_4
X_85076_ _85042_/CLK _85076_/D _45595_/A sky130_fd_sc_hd__dfxtp_4
X_51468_ _51465_/Y _51448_/X _51467_/X _86005_/D sky130_fd_sc_hd__a21oi_4
X_82288_ _82288_/CLK _82288_/D _40852_/B sky130_fd_sc_hd__dfxtp_4
X_41221_ _41205_/X _41206_/X _41220_/X _88255_/Q _41194_/X _41221_/Y
+ sky130_fd_sc_hd__o32ai_4
X_53207_ _53211_/A _53211_/B _53195_/X _53207_/D _53207_/X sky130_fd_sc_hd__and4_4
X_72041_ _83296_/Q _72001_/X _72040_/Y _72041_/Y sky130_fd_sc_hd__o21ai_4
X_84027_ _82067_/CLK _68147_/X _82067_/D sky130_fd_sc_hd__dfxtp_4
X_50419_ _50481_/A _52121_/B _50419_/Y sky130_fd_sc_hd__nand2_4
X_81239_ _85335_/CLK _81047_/Q _81239_/Q sky130_fd_sc_hd__dfxtp_4
X_54187_ _54185_/Y _54171_/X _54186_/X _54187_/Y sky130_fd_sc_hd__a21oi_4
X_51399_ _86017_/Q _51209_/X _51398_/Y _51399_/Y sky130_fd_sc_hd__o21ai_4
X_53138_ _53112_/A _53139_/A sky130_fd_sc_hd__buf_2
X_41152_ _40941_/A _41152_/X sky130_fd_sc_hd__buf_2
X_58995_ _58334_/X _58993_/Y _58994_/Y _58995_/Y sky130_fd_sc_hd__a21oi_4
X_75800_ _75800_/A _75800_/B _80891_/D sky130_fd_sc_hd__xnor2_4
X_45960_ _45954_/X _74831_/A _45933_/Y _45958_/X _45959_/X _45961_/A
+ sky130_fd_sc_hd__a32o_4
X_41083_ _41040_/X _41041_/X _41082_/X _88281_/Q _41037_/X _41084_/A
+ sky130_fd_sc_hd__o32ai_4
X_53069_ _53069_/A _53069_/X sky130_fd_sc_hd__buf_2
X_57946_ _57760_/X _85393_/Q _57945_/X _57946_/Y sky130_fd_sc_hd__o21ai_4
X_76780_ _81487_/Q _81359_/D _76779_/X _76780_/Y sky130_fd_sc_hd__o21ai_4
X_73992_ _73985_/Y _73986_/Y _73991_/X _73992_/Y sky130_fd_sc_hd__o21ai_4
X_85978_ _85974_/CLK _85978_/D _85978_/Q sky130_fd_sc_hd__dfxtp_4
X_44911_ _45824_/B _44911_/X sky130_fd_sc_hd__buf_2
X_75731_ _81011_/Q _75731_/B _75731_/X sky130_fd_sc_hd__xor2_4
X_87717_ _87394_/CLK _42790_/X _87717_/Q sky130_fd_sc_hd__dfxtp_4
X_72943_ _72943_/A _72943_/X sky130_fd_sc_hd__buf_2
X_84929_ _85379_/CLK _84929_/D _84929_/Q sky130_fd_sc_hd__dfxtp_4
X_57877_ _57875_/X _85399_/Q _57876_/X _57877_/Y sky130_fd_sc_hd__o21ai_4
X_45891_ _45890_/X _45891_/X sky130_fd_sc_hd__buf_2
X_47630_ _47625_/Y _47602_/X _47629_/X _47630_/Y sky130_fd_sc_hd__a21oi_4
X_59616_ _44008_/A _61078_/B _59893_/C sky130_fd_sc_hd__nor2_4
X_78450_ _78450_/A _78450_/B _78450_/C _78450_/Y sky130_fd_sc_hd__nor3_4
X_44842_ _41727_/A _44838_/X _67773_/B _44839_/X _44842_/X sky130_fd_sc_hd__a2bb2o_4
X_56828_ _56756_/X _56788_/X _56732_/X _56828_/Y sky130_fd_sc_hd__a21oi_4
X_87648_ _87646_/CLK _87648_/D _87648_/Q sky130_fd_sc_hd__dfxtp_4
X_75662_ _75637_/Y _75662_/Y sky130_fd_sc_hd__inv_2
X_72874_ _72874_/A _65489_/B _72874_/X sky130_fd_sc_hd__and2_4
X_77401_ _77387_/X _77399_/Y _77400_/Y _77401_/X sky130_fd_sc_hd__a21o_4
X_74613_ _74552_/X _74613_/X sky130_fd_sc_hd__buf_2
X_47561_ _47561_/A _47561_/Y sky130_fd_sc_hd__inv_2
X_71825_ _71824_/Y _71825_/X sky130_fd_sc_hd__buf_2
X_59547_ _59564_/A _59562_/B _59741_/C _60183_/A sky130_fd_sc_hd__nand3_4
X_78381_ _78363_/Y _78369_/B _78365_/A _78382_/B sky130_fd_sc_hd__o21ai_4
X_44773_ _41351_/Y _44754_/X _86963_/Q _44755_/X _86963_/D sky130_fd_sc_hd__a2bb2o_4
X_56759_ _83336_/Q _56759_/X sky130_fd_sc_hd__buf_2
X_75593_ _75590_/X _75591_/Y _75594_/B _75595_/A sky130_fd_sc_hd__a21o_4
X_87579_ _88108_/CLK _87579_/D _74123_/A sky130_fd_sc_hd__dfxtp_4
X_41985_ _41982_/X _41975_/X _40771_/X _41983_/Y _41984_/X _41985_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49300_ _49415_/A _49300_/X sky130_fd_sc_hd__buf_2
X_46512_ _46434_/A _49320_/B _46512_/Y sky130_fd_sc_hd__nand2_4
X_77332_ _77327_/Y _77329_/Y _77332_/C _77333_/A sky130_fd_sc_hd__nand3_4
X_43724_ _43724_/A _69838_/B sky130_fd_sc_hd__inv_2
X_74544_ _56004_/X _74538_/Y _74543_/Y _83040_/D sky130_fd_sc_hd__o21ai_4
X_40936_ _40935_/X _40904_/X _88307_/Q _40905_/X _40936_/X sky130_fd_sc_hd__a2bb2o_4
X_47492_ _58097_/A _47478_/X _47491_/Y _47492_/Y sky130_fd_sc_hd__o21ai_4
X_71756_ _71183_/A _71753_/B _71755_/X _71753_/D _71756_/Y sky130_fd_sc_hd__nand4_4
X_59478_ _59478_/A _59478_/B _59478_/Y sky130_fd_sc_hd__nand2_4
X_49231_ _49229_/Y _49189_/X _49230_/X _86429_/D sky130_fd_sc_hd__a21oi_4
X_70707_ _70721_/A _70710_/D sky130_fd_sc_hd__buf_2
X_46443_ _46421_/A _51320_/B _46443_/Y sky130_fd_sc_hd__nand2_4
X_58429_ _84850_/Q _58429_/Y sky130_fd_sc_hd__inv_2
X_77263_ _77265_/A _77265_/B _77264_/A sky130_fd_sc_hd__nor2_4
X_43655_ _43602_/X _43685_/A sky130_fd_sc_hd__buf_2
X_74475_ _46280_/A _74490_/A sky130_fd_sc_hd__buf_2
X_40867_ _40832_/A _40867_/X sky130_fd_sc_hd__buf_2
X_71687_ _58493_/Y _71669_/A _71686_/Y _83411_/D sky130_fd_sc_hd__o21ai_4
X_79002_ _82648_/Q _79002_/Y sky130_fd_sc_hd__inv_2
X_76214_ _81255_/Q _81511_/D _76215_/A sky130_fd_sc_hd__nor2_4
X_42606_ _42590_/X _42592_/X _40894_/X _69882_/A _42597_/X _42607_/A
+ sky130_fd_sc_hd__o32ai_4
X_49162_ _49128_/X _48664_/A _49161_/Y _49163_/A sky130_fd_sc_hd__a21o_4
X_61440_ _61440_/A _61404_/X _61406_/C _61390_/D _61440_/Y sky130_fd_sc_hd__nand4_4
X_73426_ _73426_/A _86471_/Q _73426_/X sky130_fd_sc_hd__and2_4
X_46374_ _46362_/A _53993_/B _46374_/Y sky130_fd_sc_hd__nand2_4
X_70638_ _70638_/A _70638_/X sky130_fd_sc_hd__buf_2
X_77194_ _77194_/A _77194_/B _77202_/C sky130_fd_sc_hd__nand2_4
X_43586_ _43585_/X _43586_/X sky130_fd_sc_hd__buf_2
X_40798_ _40798_/A _40798_/X sky130_fd_sc_hd__buf_2
X_48113_ _48108_/Y _48109_/X _48112_/X _48113_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_391_0_CLK clkbuf_9_195_0_CLK/X _83229_/CLK sky130_fd_sc_hd__clkbuf_1
X_45325_ _85253_/Q _45297_/X _45324_/X _45325_/Y sky130_fd_sc_hd__o21ai_4
X_76145_ _76145_/A _76145_/B _76145_/Y sky130_fd_sc_hd__nand2_4
X_42537_ _87829_/Q _69089_/B sky130_fd_sc_hd__inv_2
X_73357_ _73355_/X _85578_/Q _73284_/X _73356_/X _73357_/X sky130_fd_sc_hd__a211o_4
X_49093_ _49093_/A _53886_/B sky130_fd_sc_hd__inv_2
X_61371_ _61384_/A _61384_/B _79154_/B _61371_/Y sky130_fd_sc_hd__nor3_4
X_70569_ _70532_/Y _83747_/Q _70568_/Y _83747_/D sky130_fd_sc_hd__a21o_4
X_63110_ _63100_/A _63110_/B _63079_/C _63066_/D _63110_/X sky130_fd_sc_hd__and4_4
X_48044_ _48044_/A _48044_/B _48044_/Y sky130_fd_sc_hd__nand2_4
X_60322_ _60268_/Y _60350_/A _79713_/A _59868_/X _60322_/X sky130_fd_sc_hd__a2bb2o_4
X_72308_ _58126_/A _72308_/X sky130_fd_sc_hd__buf_2
X_45256_ _85290_/Q _45194_/X _45229_/X _45256_/X sky130_fd_sc_hd__o21a_4
X_64090_ _63265_/B _64118_/B _64155_/C _64142_/D _64090_/Y sky130_fd_sc_hd__nand4_4
X_76076_ _76068_/A _76073_/A _76076_/X sky130_fd_sc_hd__and2_4
X_42468_ _42466_/X _42467_/X _40605_/X _87855_/Q _42453_/X _42468_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73288_ _73407_/A _86509_/Q _73288_/X sky130_fd_sc_hd__and2_4
X_44207_ _44207_/A _58547_/A sky130_fd_sc_hd__buf_2
X_63041_ _63041_/A _63041_/B _63030_/C _60541_/C _63041_/X sky130_fd_sc_hd__and4_4
X_75027_ _75030_/A _75026_/Y _75028_/B sky130_fd_sc_hd__xor2_4
X_79904_ _84923_/Q _84171_/Q _79911_/A sky130_fd_sc_hd__nand2_4
X_41419_ _41253_/A _41419_/X sky130_fd_sc_hd__buf_2
X_60253_ _60253_/A _60268_/C sky130_fd_sc_hd__buf_2
X_72239_ _72166_/X _85367_/Q _72238_/X _72239_/Y sky130_fd_sc_hd__o21ai_4
X_45187_ _56339_/C _45131_/X _45161_/X _45187_/X sky130_fd_sc_hd__o21a_4
X_42399_ _42378_/X _42397_/X _40426_/X _87881_/Q _42398_/X _42400_/A
+ sky130_fd_sc_hd__o32ai_4
X_44138_ _44026_/Y _44041_/Y _44163_/B _44138_/Y sky130_fd_sc_hd__a21oi_4
X_79835_ _64764_/C _72179_/Y _79834_/Y _79835_/X sky130_fd_sc_hd__o21a_4
X_60184_ _60184_/A _61278_/B sky130_fd_sc_hd__buf_2
X_49995_ _49995_/A _49994_/X _50005_/C _53207_/D _49995_/X sky130_fd_sc_hd__and4_4
X_66800_ _66796_/X _66799_/X _66726_/X _66800_/X sky130_fd_sc_hd__a21o_4
X_48946_ _48946_/A _48946_/X sky130_fd_sc_hd__buf_2
X_44069_ _44086_/A _44070_/B sky130_fd_sc_hd__buf_2
X_67780_ _67664_/X _67769_/Y _67747_/X _67779_/Y _67780_/X sky130_fd_sc_hd__a211o_4
X_79766_ _79762_/X _79766_/B _79766_/X sky130_fd_sc_hd__xor2_4
X_64992_ _64877_/X _64992_/B _64992_/X sky130_fd_sc_hd__and2_4
X_76978_ _84530_/Q _84402_/Q _76978_/X sky130_fd_sc_hd__xor2_4
X_66731_ _66526_/X _66720_/Y _66672_/X _66730_/Y _66731_/X sky130_fd_sc_hd__a211o_4
X_78717_ _78713_/X _78718_/C _78716_/Y _78717_/X sky130_fd_sc_hd__a21o_4
X_63943_ _63939_/X _63890_/X _63940_/Y _63941_/Y _63942_/X _63943_/X
+ sky130_fd_sc_hd__a41o_4
X_75929_ _75929_/A _75929_/B _81788_/D sky130_fd_sc_hd__xor2_4
X_48877_ _48876_/Y _48878_/B sky130_fd_sc_hd__buf_2
X_79697_ _84215_/Q _83263_/Q _79697_/Y sky130_fd_sc_hd__nand2_4
X_69450_ _69423_/X _69448_/Y _69405_/X _69449_/Y _69450_/X sky130_fd_sc_hd__a211o_4
X_47828_ _48914_/A _82945_/Q _47827_/Y _47829_/A sky130_fd_sc_hd__o21a_4
X_66662_ _66689_/A _87695_/Q _66662_/X sky130_fd_sc_hd__and2_4
X_78648_ _78648_/A _78648_/Y sky130_fd_sc_hd__inv_2
X_63874_ _63867_/Y _63869_/Y _63871_/Y _63873_/Y _63874_/X sky130_fd_sc_hd__and4_4
X_68401_ _68391_/X _68398_/X _68400_/X _68401_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_450_0_CLK clkbuf_9_451_0_CLK/A clkbuf_9_450_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_65613_ _65503_/X _85589_/Q _65504_/X _65612_/X _65613_/X sky130_fd_sc_hd__a211o_4
X_62825_ _62792_/X _62839_/B _62825_/C _62825_/Y sky130_fd_sc_hd__nor3_4
X_69381_ _69234_/A _69381_/B _69381_/X sky130_fd_sc_hd__and2_4
X_47759_ _47754_/Y _47745_/X _47758_/X _86601_/D sky130_fd_sc_hd__a21oi_4
X_66593_ _69457_/A _66593_/X sky130_fd_sc_hd__buf_2
X_78579_ _78578_/X _78560_/A _78558_/X _78579_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_344_0_CLK clkbuf_9_172_0_CLK/X _86351_/CLK sky130_fd_sc_hd__clkbuf_1
X_80610_ _80607_/X _80610_/B _82271_/D sky130_fd_sc_hd__xor2_4
X_68332_ _68034_/X _68036_/X _68331_/X _68332_/Y sky130_fd_sc_hd__a21oi_4
X_65544_ _64808_/X _65647_/B _64811_/X _65544_/Y sky130_fd_sc_hd__nand3_4
X_50770_ _50767_/Y _50768_/X _50769_/Y _50770_/Y sky130_fd_sc_hd__a21boi_4
X_62756_ _62751_/Y _62713_/X _62753_/Y _62754_/Y _62755_/X _62756_/X
+ sky130_fd_sc_hd__a41o_4
X_81590_ _81330_/CLK _84190_/Q _81590_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_974_0_CLK clkbuf_9_487_0_CLK/X _86525_/CLK sky130_fd_sc_hd__clkbuf_1
X_49429_ _49420_/A _49447_/B _49420_/C _46736_/X _49429_/X sky130_fd_sc_hd__and4_4
X_61707_ _63355_/A _61706_/X _59763_/A _61715_/B sky130_fd_sc_hd__a21o_4
X_80541_ _80537_/X _80541_/B _80551_/B sky130_fd_sc_hd__xor2_4
X_68263_ _83998_/Q _68259_/X _68262_/X _68263_/X sky130_fd_sc_hd__a21bo_4
X_65475_ _65474_/X _72843_/B _65475_/X sky130_fd_sc_hd__and2_4
X_62687_ _62673_/A _62673_/B _84391_/Q _62687_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_9_465_0_CLK clkbuf_8_232_0_CLK/X clkbuf_9_465_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_67214_ _87864_/Q _67117_/X _67167_/X _67213_/X _67214_/X sky130_fd_sc_hd__a211o_4
X_52440_ _52466_/A _52440_/B _52440_/Y sky130_fd_sc_hd__nand2_4
X_64426_ _64419_/Y _64420_/X _64422_/X _64425_/Y _64384_/X _64426_/X
+ sky130_fd_sc_hd__o41a_4
X_83260_ _81227_/CLK _83260_/D _83260_/Q sky130_fd_sc_hd__dfxtp_4
X_61638_ _61608_/X _61637_/X _61619_/C _61638_/Y sky130_fd_sc_hd__nand3_4
X_80472_ _80472_/A _80472_/B _80472_/Y sky130_fd_sc_hd__nand2_4
X_68194_ _68188_/X _67197_/Y _68189_/X _68193_/Y _68194_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_359_0_CLK clkbuf_9_179_0_CLK/X _82390_/CLK sky130_fd_sc_hd__clkbuf_1
X_82211_ _82211_/CLK _82243_/Q _77239_/B sky130_fd_sc_hd__dfxtp_4
X_67145_ _67241_/A _86814_/Q _67145_/X sky130_fd_sc_hd__and2_4
X_52371_ _52368_/Y _52364_/X _52370_/X _52371_/Y sky130_fd_sc_hd__a21oi_4
X_64357_ _64352_/X _64353_/X _64354_/X _64356_/Y _64326_/X _64357_/X
+ sky130_fd_sc_hd__o41a_4
X_83191_ _83191_/CLK _72682_/X _70225_/C sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_989_0_CLK clkbuf_9_494_0_CLK/X _85558_/CLK sky130_fd_sc_hd__clkbuf_1
X_61569_ _84861_/Q _61570_/B sky130_fd_sc_hd__buf_2
X_54110_ _54217_/A _54123_/B sky130_fd_sc_hd__buf_2
X_51322_ _50812_/A _51266_/B _51330_/C _51322_/X sky130_fd_sc_hd__and3_4
X_63308_ _63303_/X _63284_/X _63307_/Y _63308_/Y sky130_fd_sc_hd__a21oi_4
X_82142_ _82575_/CLK _82142_/D _77468_/B sky130_fd_sc_hd__dfxtp_4
X_55090_ _85320_/Q _55072_/X _55089_/Y _55090_/Y sky130_fd_sc_hd__o21ai_4
X_67076_ _67028_/A _88126_/Q _67076_/X sky130_fd_sc_hd__and2_4
X_64288_ _59471_/A _64249_/X _64287_/Y _64288_/Y sky130_fd_sc_hd__o21ai_4
X_54041_ _54037_/A _52522_/B _54041_/Y sky130_fd_sc_hd__nand2_4
X_66027_ _65407_/A _66027_/X sky130_fd_sc_hd__buf_2
X_51253_ _51240_/A _46295_/X _51253_/Y sky130_fd_sc_hd__nand2_4
X_63239_ _63203_/X _84837_/Q _63204_/X _63239_/D _63239_/X sky130_fd_sc_hd__and4_4
X_86950_ _88208_/CLK _44797_/Y _86950_/Q sky130_fd_sc_hd__dfxtp_4
X_82073_ _81154_/CLK _82073_/D _82073_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_912_0_CLK clkbuf_9_456_0_CLK/X _82553_/CLK sky130_fd_sc_hd__clkbuf_1
X_50204_ _86243_/Q _50185_/X _50203_/Y _50204_/Y sky130_fd_sc_hd__o21ai_4
X_85901_ _86530_/CLK _85901_/D _85901_/Q sky130_fd_sc_hd__dfxtp_4
X_81024_ _84175_/CLK _81024_/D _81024_/Q sky130_fd_sc_hd__dfxtp_4
X_51184_ _51129_/A _51184_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_1_0_CLK clkbuf_9_0_0_CLK/X _86900_/CLK sky130_fd_sc_hd__clkbuf_1
X_86881_ _86882_/CLK _45372_/Y _64545_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_403_0_CLK clkbuf_9_402_0_CLK/A clkbuf_9_403_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_57800_ _57800_/A _57800_/X sky130_fd_sc_hd__buf_2
X_50135_ _50645_/A _50645_/B _47848_/X _50135_/X sky130_fd_sc_hd__o21a_4
X_85832_ _86154_/CLK _52392_/Y _65247_/B sky130_fd_sc_hd__dfxtp_4
X_58780_ _86704_/Q _58688_/B _58780_/Y sky130_fd_sc_hd__nor2_4
X_55992_ _55802_/X _55811_/X _56108_/A _56102_/B sky130_fd_sc_hd__nand3_4
X_67978_ _67973_/X _67976_/X _67977_/X _67978_/X sky130_fd_sc_hd__a21o_4
X_57731_ _44151_/X _57731_/B _57731_/Y sky130_fd_sc_hd__nor2_4
X_69717_ _83902_/Q _69696_/X _69716_/X _83902_/D sky130_fd_sc_hd__a21bo_4
X_50066_ _86271_/Q _50061_/X _50065_/Y _50066_/Y sky130_fd_sc_hd__o21ai_4
X_54943_ _54940_/Y _54936_/X _54942_/X _54943_/Y sky130_fd_sc_hd__a21oi_4
X_66929_ _66902_/X _86791_/Q _66929_/X sky130_fd_sc_hd__and2_4
X_85763_ _85764_/CLK _85763_/D _85763_/Q sky130_fd_sc_hd__dfxtp_4
X_82975_ _82975_/CLK _82783_/Q _46637_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_927_0_CLK clkbuf_9_463_0_CLK/X _86570_/CLK sky130_fd_sc_hd__clkbuf_1
X_87502_ _87520_/CLK _87502_/D _87502_/Q sky130_fd_sc_hd__dfxtp_4
X_84714_ _84714_/CLK _59507_/Y _64295_/C sky130_fd_sc_hd__dfxtp_4
X_57662_ _57650_/X _57659_/Y _57661_/Y _84959_/D sky130_fd_sc_hd__a21oi_4
X_81926_ _82124_/CLK _81926_/D _81926_/Q sky130_fd_sc_hd__dfxtp_4
X_69648_ _69648_/A _42558_/Y _69648_/Y sky130_fd_sc_hd__nor2_4
X_54874_ _54883_/A _54883_/B _54883_/C _53181_/D _54874_/X sky130_fd_sc_hd__and4_4
X_85694_ _85692_/CLK _85694_/D _85694_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_418_0_CLK clkbuf_9_419_0_CLK/A clkbuf_9_418_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_59401_ _84742_/Q _63139_/A sky130_fd_sc_hd__inv_2
X_56613_ _56613_/A _56613_/X sky130_fd_sc_hd__buf_2
X_87433_ _86796_/CLK _87433_/D _87433_/Q sky130_fd_sc_hd__dfxtp_4
X_53825_ _53825_/A _71998_/B _53825_/Y sky130_fd_sc_hd__nand2_4
X_84645_ _84645_/CLK _60261_/Y _79837_/A sky130_fd_sc_hd__dfxtp_4
X_57593_ _48046_/A _57619_/B _71960_/C _57593_/X sky130_fd_sc_hd__and3_4
X_69579_ _69746_/A _69579_/X sky130_fd_sc_hd__buf_2
X_81857_ _81857_/CLK _81857_/D _77715_/A sky130_fd_sc_hd__dfxtp_4
X_71610_ _71604_/X _83440_/Q _71609_/Y _83440_/D sky130_fd_sc_hd__a21o_4
X_59332_ _59273_/X _85638_/Q _59308_/X _59332_/X sky130_fd_sc_hd__o21a_4
X_56544_ _56175_/A _57364_/D _56174_/X _56546_/A sky130_fd_sc_hd__nand3_4
X_80808_ _80776_/CLK _80808_/D _80808_/Q sky130_fd_sc_hd__dfxtp_4
X_87364_ _86824_/CLK _87364_/D _87364_/Q sky130_fd_sc_hd__dfxtp_4
X_41770_ _48135_/A _48946_/A sky130_fd_sc_hd__buf_2
X_53756_ _53766_/A _48660_/A _53756_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_6_3_0_CLK clkbuf_6_3_0_CLK/A clkbuf_7_6_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_72590_ _72590_/A _72590_/X sky130_fd_sc_hd__buf_2
X_84576_ _84562_/CLK _60747_/Y _60746_/C sky130_fd_sc_hd__dfxtp_4
X_50968_ _86098_/Q _50965_/X _50967_/Y _50968_/Y sky130_fd_sc_hd__o21ai_4
X_81788_ _86753_/CLK _81788_/D _81788_/Q sky130_fd_sc_hd__dfxtp_4
X_86315_ _86312_/CLK _49836_/Y _58026_/B sky130_fd_sc_hd__dfxtp_4
X_40721_ _40716_/X _40719_/X _88348_/Q _40720_/X _40721_/X sky130_fd_sc_hd__a2bb2o_4
X_52707_ _85769_/Q _52684_/X _52706_/Y _52707_/Y sky130_fd_sc_hd__o21ai_4
X_59263_ _59037_/A _59263_/X sky130_fd_sc_hd__buf_2
X_71541_ _71585_/A _71546_/B sky130_fd_sc_hd__buf_2
X_83527_ _83498_/CLK _71358_/X _83527_/Q sky130_fd_sc_hd__dfxtp_4
X_56475_ _56474_/X _56472_/B _55960_/B _56475_/Y sky130_fd_sc_hd__nand3_4
X_80739_ _80740_/CLK _75094_/X _81147_/D sky130_fd_sc_hd__dfxtp_4
X_87295_ _87814_/CLK _43726_/Y _43724_/A sky130_fd_sc_hd__dfxtp_4
X_53687_ _53687_/A _53687_/X sky130_fd_sc_hd__buf_2
X_50899_ _50894_/Y _50839_/X _50898_/X _50899_/Y sky130_fd_sc_hd__a21oi_4
X_58214_ _63713_/A _58217_/B _58214_/Y sky130_fd_sc_hd__nand2_4
XPHY_400 sky130_fd_sc_hd__decap_3
X_55426_ _55156_/X _55160_/X _55426_/X sky130_fd_sc_hd__and2_4
X_43440_ _41580_/X _43431_/X _87420_/Q _43432_/X _43440_/X sky130_fd_sc_hd__a2bb2o_4
X_74260_ _74248_/X _74250_/X _74259_/X _74260_/X sky130_fd_sc_hd__a21o_4
X_86246_ _86246_/CLK _86246_/D _65315_/B sky130_fd_sc_hd__dfxtp_4
XPHY_411 sky130_fd_sc_hd__decap_3
X_52638_ _85782_/Q _52629_/X _52637_/Y _52638_/Y sky130_fd_sc_hd__o21ai_4
X_40652_ _40599_/A _40652_/X sky130_fd_sc_hd__buf_2
X_71472_ _71464_/X _83487_/Q _71471_/X _71472_/X sky130_fd_sc_hd__a21o_4
X_59194_ _86673_/Q _59282_/B _59194_/Y sky130_fd_sc_hd__nor2_4
X_83458_ _83495_/CLK _83458_/D _83458_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_422 sky130_fd_sc_hd__decap_3
XPHY_433 sky130_fd_sc_hd__decap_3
X_73211_ _73260_/A _86480_/Q _73211_/X sky130_fd_sc_hd__and2_4
XPHY_444 sky130_fd_sc_hd__decap_3
X_70423_ HASH_ADDR[0] _70423_/X sky130_fd_sc_hd__buf_2
X_58145_ _83497_/Q _58145_/Y sky130_fd_sc_hd__inv_2
X_82409_ _82820_/CLK _82409_/D _78403_/A sky130_fd_sc_hd__dfxtp_4
XPHY_455 sky130_fd_sc_hd__decap_3
X_43371_ _43396_/A _43371_/X sky130_fd_sc_hd__buf_2
X_55357_ _56708_/A _55445_/D _55353_/X _55369_/B sky130_fd_sc_hd__a21bo_4
X_74191_ _74188_/X _74190_/X _74191_/Y sky130_fd_sc_hd__nand2_4
X_86177_ _83311_/CLK _86177_/D _86177_/Q sky130_fd_sc_hd__dfxtp_4
X_40583_ _40583_/A _40583_/Y sky130_fd_sc_hd__inv_2
X_52569_ _52280_/X _54087_/B _52569_/Y sky130_fd_sc_hd__nand2_4
XPHY_466 sky130_fd_sc_hd__decap_3
X_83389_ _85499_/CLK _71752_/Y _47259_/A sky130_fd_sc_hd__dfxtp_4
XPHY_477 sky130_fd_sc_hd__decap_3
XPHY_488 sky130_fd_sc_hd__decap_3
X_45110_ _64364_/B _61489_/B sky130_fd_sc_hd__buf_2
X_42322_ _42321_/Y _42322_/Y sky130_fd_sc_hd__inv_2
X_54308_ _54306_/Y _54285_/X _54307_/X _54308_/Y sky130_fd_sc_hd__a21oi_4
XPHY_499 sky130_fd_sc_hd__decap_3
X_73142_ _73128_/X _73131_/Y _73141_/X _73142_/X sky130_fd_sc_hd__a21o_4
X_85128_ _85128_/CLK _56855_/Y _85128_/Q sky130_fd_sc_hd__dfxtp_4
X_46090_ _46112_/A _46090_/Y sky130_fd_sc_hd__inv_2
X_58076_ _58043_/X _85991_/Q _58075_/X _58076_/Y sky130_fd_sc_hd__o21ai_4
X_70354_ _70496_/A _70412_/A HASH_ADDR[4] MACRO_WR_SELECT _70355_/A
+ sky130_fd_sc_hd__and4_4
X_55288_ _55288_/A _55288_/B _55288_/C _55287_/X _55288_/Y sky130_fd_sc_hd__nand4_4
X_45041_ _85176_/Q _44982_/X _45040_/X _45041_/X sky130_fd_sc_hd__o21a_4
X_57027_ _57027_/A _57026_/X _57027_/Y sky130_fd_sc_hd__nor2_4
X_42253_ _42252_/X _42243_/X _41442_/X _87958_/Q _42244_/X _42254_/A
+ sky130_fd_sc_hd__o32ai_4
X_73073_ _73073_/A _73073_/B _73073_/X sky130_fd_sc_hd__xor2_4
X_54239_ _54230_/A _53072_/B _54239_/Y sky130_fd_sc_hd__nand2_4
X_77950_ _77950_/A _77950_/B _77951_/B sky130_fd_sc_hd__xor2_4
X_85059_ _85005_/CLK _85059_/D _85059_/Q sky130_fd_sc_hd__dfxtp_4
X_70285_ _70292_/A _70292_/B _70285_/C _70292_/D _70285_/X sky130_fd_sc_hd__and4_4
X_41204_ _41203_/X _41181_/X _68796_/B _41182_/X _41204_/X sky130_fd_sc_hd__a2bb2o_4
X_72024_ _71993_/A _72025_/A sky130_fd_sc_hd__buf_2
X_76901_ _76901_/A _76893_/Y _76899_/Y _76902_/B sky130_fd_sc_hd__nand3_4
X_42184_ _42162_/A _42184_/X sky130_fd_sc_hd__buf_2
X_77881_ _82162_/Q _77880_/X _82130_/D sky130_fd_sc_hd__xor2_4
X_48800_ _86480_/Q _48781_/X _48799_/Y _48800_/Y sky130_fd_sc_hd__o21ai_4
X_79620_ _79620_/A _79624_/A sky130_fd_sc_hd__inv_2
X_41135_ _41134_/X _41109_/X _68485_/B _41110_/X _41135_/X sky130_fd_sc_hd__a2bb2o_4
X_76832_ _76821_/Y _76832_/Y sky130_fd_sc_hd__inv_2
X_49780_ _49775_/Y _49759_/X _49779_/X _86325_/D sky130_fd_sc_hd__a21oi_4
X_46992_ _46986_/Y _46987_/X _46991_/X _86682_/D sky130_fd_sc_hd__a21oi_4
X_58978_ _84782_/Q _58978_/Y sky130_fd_sc_hd__inv_2
X_48731_ _48731_/A _48737_/A sky130_fd_sc_hd__buf_2
X_79551_ _79549_/Y _79550_/Y _79555_/A sky130_fd_sc_hd__nand2_4
X_45943_ _45943_/A _64961_/A sky130_fd_sc_hd__buf_2
X_41066_ _40989_/A _41066_/X sky130_fd_sc_hd__buf_2
X_57929_ _57925_/Y _57928_/Y _57889_/X _57929_/X sky130_fd_sc_hd__a21o_4
X_76763_ _76763_/A _76762_/Y _76764_/B sky130_fd_sc_hd__xor2_4
X_73975_ _73971_/X _73974_/X _73857_/X _73978_/A sky130_fd_sc_hd__a21o_4
X_78502_ _78503_/A _82672_/D _78505_/B sky130_fd_sc_hd__nor2_4
X_75714_ _81090_/Q _75714_/B _75714_/Y sky130_fd_sc_hd__xnor2_4
X_48662_ _86502_/Q _48612_/X _48661_/Y _48662_/Y sky130_fd_sc_hd__o21ai_4
X_60940_ _60901_/A _64172_/D _60957_/B _60940_/Y sky130_fd_sc_hd__nor3_4
X_72926_ _72923_/X _72925_/X _72737_/X _72926_/X sky130_fd_sc_hd__a21o_4
X_79482_ _79481_/Y _79482_/B _79482_/X sky130_fd_sc_hd__and2_4
X_45874_ _85122_/Q _45627_/X _44889_/A _45874_/X sky130_fd_sc_hd__o21a_4
X_76694_ _76694_/A _76694_/B _81447_/D sky130_fd_sc_hd__xnor2_4
X_47613_ _46902_/A _47661_/A sky130_fd_sc_hd__buf_2
X_78433_ _78434_/B _78434_/A _78439_/B sky130_fd_sc_hd__or2_4
X_44825_ _44825_/A _86935_/D sky130_fd_sc_hd__inv_2
X_75645_ _75625_/Y _75641_/A _75644_/X _75645_/Y sky130_fd_sc_hd__a21oi_4
X_48593_ _48593_/A _48820_/B sky130_fd_sc_hd__buf_2
X_72857_ _73092_/A _72857_/X sky130_fd_sc_hd__buf_2
X_60871_ _60857_/D _60844_/X _60863_/X _60871_/Y sky130_fd_sc_hd__a21boi_4
X_62610_ _62196_/X _62162_/X _62609_/X _62610_/X sky130_fd_sc_hd__a21o_4
X_47544_ _47543_/Y _53109_/B sky130_fd_sc_hd__buf_2
X_71808_ _71779_/A _71424_/C _70852_/C _71808_/X sky130_fd_sc_hd__and3_4
X_78364_ _78362_/Y _78359_/X _78364_/C _78365_/A sky130_fd_sc_hd__nand3_4
X_44756_ _41301_/Y _44754_/X _86972_/Q _44755_/X _44756_/X sky130_fd_sc_hd__a2bb2o_4
X_63590_ _63528_/A _63615_/A sky130_fd_sc_hd__buf_2
X_75576_ _75573_/Y _75575_/Y _75570_/A _75586_/A sky130_fd_sc_hd__a21oi_4
X_41968_ _41965_/X _41956_/X _40734_/X _41966_/Y _41967_/X _88089_/D
+ sky130_fd_sc_hd__o32ai_4
X_72788_ _72783_/X _72788_/B _72789_/B sky130_fd_sc_hd__nand2_4
X_77315_ _77315_/A _77315_/B _77315_/C _77316_/B sky130_fd_sc_hd__nand3_4
X_43707_ _40839_/A _43698_/X _69752_/B _43700_/X _43707_/X sky130_fd_sc_hd__a2bb2o_4
X_62541_ _62483_/X _62541_/B _62541_/C _62541_/Y sky130_fd_sc_hd__nor3_4
X_74527_ _74527_/A _74531_/B _74531_/C _74531_/D _74527_/Y sky130_fd_sc_hd__nand4_4
X_40919_ _46469_/B _40919_/B _40919_/X sky130_fd_sc_hd__or2_4
X_47475_ _47437_/X _47463_/X _47513_/C _53070_/D _47475_/X sky130_fd_sc_hd__and4_4
X_71739_ _71738_/X _71753_/D sky130_fd_sc_hd__buf_2
X_78295_ _78296_/A _78296_/B _78295_/Y sky130_fd_sc_hd__nor2_4
X_44687_ _43047_/A _44687_/X sky130_fd_sc_hd__buf_2
X_41899_ _88109_/Q _41899_/Y sky130_fd_sc_hd__inv_2
X_49214_ _49247_/A _49214_/X sky130_fd_sc_hd__buf_2
X_46426_ _46423_/X _49039_/A _46425_/Y _46427_/A sky130_fd_sc_hd__o21ai_4
X_65260_ _65159_/A _65260_/B _65260_/X sky130_fd_sc_hd__and2_4
X_77246_ _77244_/X _77261_/A _77246_/X sky130_fd_sc_hd__and2_4
X_43638_ _43637_/X _87333_/D sky130_fd_sc_hd__inv_2
X_74458_ _74458_/A _74478_/C sky130_fd_sc_hd__buf_2
X_62472_ _61551_/A _62472_/B _62490_/C _62566_/D _62472_/Y sky130_fd_sc_hd__nand4_4
X_64211_ _61182_/X _61301_/X _64211_/C _64211_/Y sky130_fd_sc_hd__nand3_4
X_49145_ _49117_/A _49144_/X _49145_/Y sky130_fd_sc_hd__nand2_4
X_61423_ _61422_/Y _61423_/Y sky130_fd_sc_hd__inv_2
X_73409_ _73409_/A _73408_/X _73409_/Y sky130_fd_sc_hd__nand2_4
X_46357_ _46326_/A _46356_/X _46357_/Y sky130_fd_sc_hd__nand2_4
X_65191_ _64835_/X _83291_/Q _65015_/X _65190_/X _65191_/X sky130_fd_sc_hd__a211o_4
X_77177_ _77177_/A _77177_/B _77178_/B sky130_fd_sc_hd__xnor2_4
X_43569_ _40507_/X _43560_/X _87356_/Q _43561_/X _43569_/X sky130_fd_sc_hd__a2bb2o_4
X_74389_ _74466_/A _74389_/B _74389_/Y sky130_fd_sc_hd__nand2_4
X_45308_ _45308_/A _61636_/B sky130_fd_sc_hd__buf_2
X_64142_ _61655_/A _64177_/B _64155_/C _64142_/D _64142_/Y sky130_fd_sc_hd__nand4_4
X_76128_ _76123_/Y _76099_/B _76127_/X _76129_/B sky130_fd_sc_hd__o21ai_4
X_61354_ _61329_/A _61354_/B _61375_/C _61354_/Y sky130_fd_sc_hd__nand3_4
X_49076_ _48995_/A _49080_/A sky130_fd_sc_hd__buf_2
X_46288_ _46288_/A _53959_/B _46288_/Y sky130_fd_sc_hd__nand2_4
X_60305_ _60268_/C _60300_/B _60337_/C _60305_/Y sky130_fd_sc_hd__o21ai_4
X_48027_ _47971_/X _46459_/A _48026_/X _48028_/B sky130_fd_sc_hd__o21ai_4
X_45239_ _56250_/C _45222_/X _45238_/X _45239_/Y sky130_fd_sc_hd__o21ai_4
X_68950_ _87080_/Q _68948_/X _68875_/X _68949_/X _68950_/X sky130_fd_sc_hd__a211o_4
X_64073_ _63912_/X _64073_/X sky130_fd_sc_hd__buf_2
X_76059_ _76052_/Y _76063_/A _76058_/Y _76060_/B sky130_fd_sc_hd__a21boi_4
X_61285_ _59536_/A _60122_/A _61285_/C _60122_/C _72621_/B sky130_fd_sc_hd__and4_4
X_63024_ _79502_/A _63008_/X _63023_/Y _84360_/D sky130_fd_sc_hd__a21o_4
X_67901_ _67901_/A _67901_/B _67901_/X sky130_fd_sc_hd__and2_4
X_60236_ _60227_/A _60254_/B sky130_fd_sc_hd__buf_2
X_68881_ _83957_/Q _68838_/X _68880_/X _68881_/X sky130_fd_sc_hd__a21bo_4
X_67832_ _67901_/A _67832_/B _67832_/X sky130_fd_sc_hd__and2_4
X_79818_ _79816_/X _79817_/X _79818_/Y sky130_fd_sc_hd__xnor2_4
X_60167_ _60387_/A _60164_/Y _60166_/X _60168_/A sky130_fd_sc_hd__and3_4
X_49978_ _46308_/A _49995_/A sky130_fd_sc_hd__buf_2
X_48929_ _48923_/Y _48880_/X _48928_/X _86461_/D sky130_fd_sc_hd__a21oi_4
X_67763_ _87969_/Q _67713_/X _67761_/X _67762_/X _67763_/X sky130_fd_sc_hd__a211o_4
X_79749_ _79736_/X _79747_/X _79748_/X _79749_/Y sky130_fd_sc_hd__a21oi_4
X_64975_ _64971_/X _86131_/Q _64972_/X _64974_/X _64975_/X sky130_fd_sc_hd__a211o_4
X_60098_ _60078_/X _60092_/B _60045_/Y _60096_/Y _60097_/Y _84662_/D
+ sky130_fd_sc_hd__a41oi_4
Xclkbuf_10_50_0_CLK clkbuf_9_25_0_CLK/X _85042_/CLK sky130_fd_sc_hd__clkbuf_1
X_69502_ _69423_/X _69499_/Y _69405_/X _69501_/Y _69502_/X sky130_fd_sc_hd__a211o_4
X_66714_ _66711_/X _66713_/X _66667_/X _66720_/A sky130_fd_sc_hd__a21o_4
X_51940_ _65932_/B _51929_/X _51939_/Y _51940_/Y sky130_fd_sc_hd__o21ai_4
X_63926_ _63942_/A _59403_/A _63958_/C _63926_/X sky130_fd_sc_hd__and3_4
X_82760_ _82961_/CLK _82760_/D _82760_/Q sky130_fd_sc_hd__dfxtp_4
X_67694_ _87396_/Q _67594_/X _67595_/X _67693_/X _67694_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_283_0_CLK clkbuf_9_141_0_CLK/X _83756_/CLK sky130_fd_sc_hd__clkbuf_1
X_81711_ _87348_/CLK _81711_/D _41207_/A sky130_fd_sc_hd__dfxtp_4
X_69433_ _69156_/A _69433_/X sky130_fd_sc_hd__buf_2
X_66645_ _87376_/Q _66642_/X _66643_/X _66644_/X _66645_/X sky130_fd_sc_hd__a211o_4
X_51871_ _51868_/Y _51850_/X _51870_/X _51871_/Y sky130_fd_sc_hd__a21oi_4
X_63857_ _64294_/B _63790_/X _63840_/C _63920_/D _63857_/Y sky130_fd_sc_hd__nand4_4
X_82691_ _82147_/CLK _78821_/X _82679_/D sky130_fd_sc_hd__dfxtp_4
X_53610_ _53846_/A _53610_/X sky130_fd_sc_hd__buf_2
X_84430_ _84430_/CLK _62145_/Y _78053_/B sky130_fd_sc_hd__dfxtp_4
X_50822_ _50822_/A _51328_/B _50822_/Y sky130_fd_sc_hd__nand2_4
X_62808_ _60217_/A _62808_/X sky130_fd_sc_hd__buf_2
X_81642_ _81275_/CLK _81674_/Q _81642_/Q sky130_fd_sc_hd__dfxtp_4
X_69364_ _69360_/X _69363_/X _69142_/X _69364_/Y sky130_fd_sc_hd__a21oi_4
X_54590_ _54537_/A _54591_/C sky130_fd_sc_hd__buf_2
Xclkbuf_10_65_0_CLK clkbuf_9_32_0_CLK/X _80670_/CLK sky130_fd_sc_hd__clkbuf_1
X_66576_ _68742_/A _69223_/A sky130_fd_sc_hd__buf_2
X_63788_ _63751_/X _63820_/D sky130_fd_sc_hd__buf_2
X_68315_ _67941_/X _67944_/X _68283_/X _68315_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_8_211_0_CLK clkbuf_8_211_0_CLK/A clkbuf_9_423_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_53541_ _53723_/A _53548_/A sky130_fd_sc_hd__buf_2
X_65527_ _65523_/X _65631_/B _65526_/X _65527_/Y sky130_fd_sc_hd__nand3_4
X_84361_ _83216_/CLK _84361_/D _79513_/A sky130_fd_sc_hd__dfxtp_4
X_50753_ _50799_/A _51261_/B _50753_/Y sky130_fd_sc_hd__nand2_4
X_62739_ _58248_/A _62689_/X _62708_/X _62699_/X _62738_/X _62739_/Y
+ sky130_fd_sc_hd__a41oi_4
X_81573_ _84079_/CLK _65855_/C _76682_/A sky130_fd_sc_hd__dfxtp_4
X_69295_ _69575_/A _69295_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_298_0_CLK clkbuf_9_149_0_CLK/X _84713_/CLK sky130_fd_sc_hd__clkbuf_1
X_86100_ _86100_/CLK _86100_/D _86100_/Q sky130_fd_sc_hd__dfxtp_4
X_83312_ _85547_/CLK _83312_/D _83312_/Q sky130_fd_sc_hd__dfxtp_4
X_80524_ _80518_/A _80518_/B _80523_/Y _80542_/A sky130_fd_sc_hd__a21boi_4
X_56260_ _56144_/X _56255_/X _56259_/Y _85256_/D sky130_fd_sc_hd__o21ai_4
X_68246_ _68376_/A _68246_/X sky130_fd_sc_hd__buf_2
X_87080_ _87083_/CLK _87080_/D _87080_/Q sky130_fd_sc_hd__dfxtp_4
X_53472_ _53982_/A _53472_/X sky130_fd_sc_hd__buf_2
X_65458_ _65452_/X _65456_/X _65457_/X _65458_/X sky130_fd_sc_hd__a21o_4
X_84292_ _84292_/CLK _63835_/Y _84292_/Q sky130_fd_sc_hd__dfxtp_4
X_50684_ _50640_/A _53902_/B _50684_/Y sky130_fd_sc_hd__nand2_4
X_55211_ _55149_/A _55211_/B _55211_/X sky130_fd_sc_hd__and2_4
X_86031_ _86424_/CLK _51327_/Y _86031_/Q sky130_fd_sc_hd__dfxtp_4
X_52423_ _52602_/A _52448_/A sky130_fd_sc_hd__buf_2
X_64409_ _58438_/A _64418_/B _64409_/Y sky130_fd_sc_hd__nor2_4
X_83243_ _84835_/CLK _83243_/D _83243_/Q sky130_fd_sc_hd__dfxtp_4
X_56191_ _56123_/A _56192_/B sky130_fd_sc_hd__buf_2
X_80455_ _80455_/A _80455_/B _80456_/B sky130_fd_sc_hd__xor2_4
X_68177_ _67109_/X _67112_/X _68169_/X _68177_/Y sky130_fd_sc_hd__a21oi_4
X_65389_ _64729_/A _65389_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_226_0_CLK clkbuf_8_227_0_CLK/A clkbuf_8_226_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_55142_ _55142_/A _55278_/A sky130_fd_sc_hd__buf_2
X_67128_ _67149_/A _67128_/B _67128_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_221_0_CLK clkbuf_9_110_0_CLK/X _84624_/CLK sky130_fd_sc_hd__clkbuf_1
X_52354_ _85839_/Q _52347_/X _52353_/Y _52354_/Y sky130_fd_sc_hd__o21ai_4
X_83174_ _83161_/CLK _83174_/D _83174_/Q sky130_fd_sc_hd__dfxtp_4
X_80386_ _80384_/Y _80366_/B _80385_/X _80386_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_851_0_CLK clkbuf_9_425_0_CLK/X _85471_/CLK sky130_fd_sc_hd__clkbuf_1
X_51305_ _86035_/Q _51285_/X _51304_/Y _51305_/Y sky130_fd_sc_hd__o21ai_4
X_82125_ _82485_/CLK _77831_/X _82125_/Q sky130_fd_sc_hd__dfxtp_4
X_55073_ _47838_/X _55093_/A sky130_fd_sc_hd__buf_2
X_59950_ _59913_/A _59950_/B _59950_/C _59973_/A _59951_/D sky130_fd_sc_hd__nand4_4
X_67059_ _66961_/X _86818_/Q _67059_/X sky130_fd_sc_hd__and2_4
X_52285_ _48928_/A _52267_/B _52267_/C _52285_/X sky130_fd_sc_hd__and3_4
X_87982_ _87472_/CLK _42198_/X _87982_/Q sky130_fd_sc_hd__dfxtp_4
X_58901_ _58877_/X _85927_/Q _58900_/X _58901_/X sky130_fd_sc_hd__o21a_4
X_54024_ _53942_/A _46441_/Y _54024_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_342_0_CLK clkbuf_9_343_0_CLK/A clkbuf_9_342_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_51236_ _64572_/B _51233_/X _51235_/Y _51236_/Y sky130_fd_sc_hd__o21ai_4
X_70070_ _82538_/D _70067_/X _70069_/X _83858_/D sky130_fd_sc_hd__a21bo_4
X_86933_ _87188_/CLK _86933_/D _86933_/Q sky130_fd_sc_hd__dfxtp_4
X_82056_ _84014_/CLK _84016_/Q _77776_/A sky130_fd_sc_hd__dfxtp_4
X_59881_ _59880_/X _59881_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_236_0_CLK clkbuf_9_118_0_CLK/X _81104_/CLK sky130_fd_sc_hd__clkbuf_1
X_81007_ _84177_/CLK _84215_/Q _81007_/Q sky130_fd_sc_hd__dfxtp_4
X_58832_ _58701_/A _58832_/X sky130_fd_sc_hd__buf_2
X_51167_ _51167_/A _52859_/B _51167_/Y sky130_fd_sc_hd__nand2_4
X_86864_ _86770_/CLK _45642_/Y _63182_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_866_0_CLK clkbuf_9_433_0_CLK/X _85915_/CLK sky130_fd_sc_hd__clkbuf_1
X_50118_ _50106_/A _53844_/B _50118_/X sky130_fd_sc_hd__and2_4
X_85815_ _85815_/CLK _52475_/Y _85815_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_18_0_CLK clkbuf_9_9_0_CLK/X _83025_/CLK sky130_fd_sc_hd__clkbuf_1
X_58763_ _58763_/A _58763_/B _58763_/Y sky130_fd_sc_hd__nor2_4
X_51098_ _86074_/Q _51073_/X _51097_/Y _51098_/Y sky130_fd_sc_hd__o21ai_4
X_55975_ _55975_/A _55975_/X sky130_fd_sc_hd__buf_2
X_86795_ _88245_/CLK _86795_/D _66830_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_357_0_CLK clkbuf_8_178_0_CLK/X clkbuf_9_357_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_57714_ _57709_/X _86017_/Q _57713_/X _57714_/Y sky130_fd_sc_hd__o21ai_4
X_42940_ _42916_/X _42917_/X _41773_/X _67985_/B _42934_/X _42940_/Y
+ sky130_fd_sc_hd__o32ai_4
X_50049_ _72475_/B _48170_/X _50048_/Y _50049_/Y sky130_fd_sc_hd__o21ai_4
X_54926_ _51340_/A _54927_/A sky130_fd_sc_hd__buf_2
X_73760_ _73735_/X _85625_/Q _73661_/X _73759_/X _73760_/X sky130_fd_sc_hd__a211o_4
X_85746_ _85748_/CLK _52836_/Y _85746_/Q sky130_fd_sc_hd__dfxtp_4
X_70972_ _70976_/A _70949_/B _70969_/C _70972_/Y sky130_fd_sc_hd__nand3_4
X_82958_ _85778_/CLK _82766_/Q _82958_/Q sky130_fd_sc_hd__dfxtp_4
X_58694_ _58691_/Y _58693_/Y _58610_/X _58694_/X sky130_fd_sc_hd__a21o_4
X_72711_ _83182_/Q _72709_/X _72710_/X _83182_/D sky130_fd_sc_hd__a21o_4
X_57645_ _57643_/Y _57627_/X _57644_/Y _57645_/Y sky130_fd_sc_hd__a21boi_4
X_81909_ _82133_/CLK _81909_/D _82285_/D sky130_fd_sc_hd__dfxtp_4
X_42871_ _41580_/X _42866_/X _67118_/B _42867_/X _42871_/X sky130_fd_sc_hd__a2bb2o_4
X_54857_ _54857_/A _54857_/B _54857_/C _53165_/D _54857_/X sky130_fd_sc_hd__and4_4
X_73691_ _73688_/X _73690_/X _73692_/B sky130_fd_sc_hd__nand2_4
X_85677_ _84802_/CLK _85677_/D _85677_/Q sky130_fd_sc_hd__dfxtp_4
X_82889_ _82317_/CLK _78128_/B _82889_/Q sky130_fd_sc_hd__dfxtp_4
X_44610_ _44609_/Y _87035_/D sky130_fd_sc_hd__inv_2
X_75430_ _75430_/A _75430_/Y sky130_fd_sc_hd__inv_2
X_87416_ _87416_/CLK _43448_/X _87416_/Q sky130_fd_sc_hd__dfxtp_4
X_41822_ _41802_/X _41803_/X _40440_/X _88135_/Q _41821_/X _41822_/Y
+ sky130_fd_sc_hd__o32ai_4
X_53808_ _53786_/A _48931_/A _53808_/Y sky130_fd_sc_hd__nand2_4
X_72642_ _70181_/A _72631_/X _72641_/Y _83206_/D sky130_fd_sc_hd__a21bo_4
X_84628_ _84645_/CLK _84628_/D _79658_/A sky130_fd_sc_hd__dfxtp_4
X_45590_ _45589_/Y _45590_/B _45590_/X sky130_fd_sc_hd__and2_4
X_57576_ _57597_/A _50322_/B _57576_/Y sky130_fd_sc_hd__nand2_4
X_88396_ _86834_/CLK _40405_/X _88396_/Q sky130_fd_sc_hd__dfxtp_4
X_54788_ _54798_/A _54788_/B _54798_/C _47521_/A _54788_/X sky130_fd_sc_hd__and4_4
X_59315_ _84752_/Q _59268_/X _59307_/X _59314_/X _84752_/D sky130_fd_sc_hd__a2bb2oi_4
X_56527_ _56134_/X _56515_/X _56526_/Y _85162_/D sky130_fd_sc_hd__o21ai_4
X_44541_ _44496_/X _44497_/X _40814_/X _73024_/A _44498_/X _44542_/A
+ sky130_fd_sc_hd__o32ai_4
X_75361_ _80694_/Q _80950_/D _75362_/B sky130_fd_sc_hd__xor2_4
X_87347_ _87345_/CLK _87347_/D _43587_/A sky130_fd_sc_hd__dfxtp_4
X_41753_ _41802_/A _41753_/X sky130_fd_sc_hd__buf_2
X_53739_ _52218_/A _53748_/B _53748_/C _53739_/X sky130_fd_sc_hd__and3_4
X_72573_ _72573_/A _72573_/B _79394_/B _72573_/Y sky130_fd_sc_hd__nor3_4
X_84559_ _84559_/CLK _84559_/D _60817_/C sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_804_0_CLK clkbuf_9_402_0_CLK/X _82595_/CLK sky130_fd_sc_hd__clkbuf_1
X_77100_ _77091_/Y _77098_/Y _77099_/Y _77100_/X sky130_fd_sc_hd__o21a_4
X_74312_ _74302_/X _74310_/B _74312_/C _74312_/Y sky130_fd_sc_hd__nand3_4
X_40704_ _40703_/Y _40704_/Y sky130_fd_sc_hd__inv_2
X_47260_ _47260_/A _52944_/B sky130_fd_sc_hd__buf_2
X_59246_ _59115_/X _59244_/Y _59245_/Y _59133_/X _59119_/X _59246_/X
+ sky130_fd_sc_hd__o32a_4
X_71524_ _53255_/B _71512_/A _71523_/Y _83467_/D sky130_fd_sc_hd__o21ai_4
X_78080_ _78080_/A _78080_/B _78080_/X sky130_fd_sc_hd__xor2_4
X_44472_ _44472_/A _87091_/D sky130_fd_sc_hd__inv_2
X_56458_ _56458_/A _56177_/B _56458_/C _56458_/Y sky130_fd_sc_hd__nand3_4
X_75292_ _75288_/Y _75291_/C _75287_/Y _75292_/Y sky130_fd_sc_hd__o21ai_4
X_41684_ _41814_/A _41684_/X sky130_fd_sc_hd__buf_2
X_87278_ _88084_/CLK _87278_/D _69206_/B sky130_fd_sc_hd__dfxtp_4
X_46211_ _69611_/A _46212_/A sky130_fd_sc_hd__buf_2
XPHY_230 sky130_fd_sc_hd__decap_3
X_77031_ _77026_/Y _77034_/B _77030_/Y _77031_/Y sky130_fd_sc_hd__a21boi_4
X_43423_ _43422_/X _43404_/X _41536_/X _87428_/Q _43407_/X _43424_/A
+ sky130_fd_sc_hd__o32ai_4
X_55409_ _55409_/A _55398_/Y _55397_/Y _55409_/Y sky130_fd_sc_hd__nand3_4
X_74243_ _70130_/B _74139_/X _74242_/Y _74243_/X sky130_fd_sc_hd__a21o_4
X_86229_ _86578_/CLK _86229_/D _86229_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_241 sky130_fd_sc_hd__decap_3
X_40635_ _44733_/A _40635_/X sky130_fd_sc_hd__buf_2
X_59177_ _59061_/A _59177_/X sky130_fd_sc_hd__buf_2
X_47191_ _47186_/Y _47177_/X _47190_/X _47191_/Y sky130_fd_sc_hd__a21oi_4
X_71455_ _71445_/X _83493_/Q _71454_/Y _71455_/X sky130_fd_sc_hd__a21o_4
X_56389_ _56026_/X _56378_/X _56388_/Y _56389_/Y sky130_fd_sc_hd__o21ai_4
XPHY_252 sky130_fd_sc_hd__decap_3
XPHY_263 sky130_fd_sc_hd__decap_3
XPHY_274 sky130_fd_sc_hd__decap_3
X_70406_ _70824_/A _74533_/A sky130_fd_sc_hd__buf_2
X_58128_ _58112_/X _85987_/Q _58127_/X _58128_/Y sky130_fd_sc_hd__o21ai_4
X_46142_ _46099_/X _46143_/D sky130_fd_sc_hd__inv_2
XPHY_285 sky130_fd_sc_hd__decap_3
X_43354_ _43347_/X _43350_/X _41347_/X _87464_/Q _43353_/X _43355_/A
+ sky130_fd_sc_hd__o32ai_4
X_74174_ _74152_/A _66285_/B _74174_/X sky130_fd_sc_hd__and2_4
X_40566_ _40565_/Y _40567_/A sky130_fd_sc_hd__inv_2
XPHY_296 sky130_fd_sc_hd__decap_3
X_71386_ _70682_/A _71386_/B _71377_/C _71386_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_10_819_0_CLK clkbuf_9_409_0_CLK/X _81198_/CLK sky130_fd_sc_hd__clkbuf_1
X_42305_ _42304_/X _42305_/X sky130_fd_sc_hd__buf_2
X_73125_ _69749_/B _73104_/B _72944_/X _73124_/Y _73125_/X sky130_fd_sc_hd__a211o_4
X_46073_ _41591_/Y _46061_/X _86781_/Q _46062_/X _46073_/X sky130_fd_sc_hd__a2bb2o_4
X_58059_ _58676_/A _58136_/B sky130_fd_sc_hd__buf_2
X_70337_ _70337_/A _70337_/X sky130_fd_sc_hd__buf_2
X_43285_ _41161_/X _43277_/X _87498_/Q _43278_/X _43285_/X sky130_fd_sc_hd__a2bb2o_4
X_78982_ _82741_/Q _78982_/B _82709_/D sky130_fd_sc_hd__xor2_4
X_40497_ _40496_/Y _40497_/X sky130_fd_sc_hd__buf_2
X_49901_ _49901_/A _53115_/B _49901_/Y sky130_fd_sc_hd__nand2_4
X_45024_ _45017_/X _45021_/Y _45023_/Y _45024_/Y sky130_fd_sc_hd__a21oi_4
X_42236_ _41393_/X _42222_/X _87967_/Q _42224_/X _42236_/X sky130_fd_sc_hd__a2bb2o_4
X_61070_ _59613_/Y _61070_/B _61070_/C _59552_/C _61070_/X sky130_fd_sc_hd__and4_4
X_77933_ _77933_/A _77933_/B _77934_/B sky130_fd_sc_hd__xor2_4
X_73056_ _73056_/A _73003_/B _73056_/Y sky130_fd_sc_hd__nor2_4
X_70268_ _70255_/X _74807_/A _70267_/X _83817_/D sky130_fd_sc_hd__a21o_4
X_60021_ _60064_/A _59873_/B _60021_/C _60021_/Y sky130_fd_sc_hd__nor3_4
X_72007_ _72007_/A _72007_/B _72007_/Y sky130_fd_sc_hd__nand2_4
X_49832_ _49827_/X _53046_/B _49832_/Y sky130_fd_sc_hd__nand2_4
X_42167_ _42154_/X _42141_/X _41214_/X _88000_/Q _42142_/X _42167_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77864_ _82273_/Q _81985_/Q _77864_/Y sky130_fd_sc_hd__xnor2_4
X_70199_ _70195_/X _74799_/C _70198_/X _70199_/X sky130_fd_sc_hd__a21o_4
X_79603_ _65294_/C _83255_/Q _79603_/Y sky130_fd_sc_hd__nand2_4
X_41118_ _41118_/A _88275_/D sky130_fd_sc_hd__inv_2
X_76815_ _76806_/A _76792_/Y _76805_/A _76804_/Y _76815_/X sky130_fd_sc_hd__o22a_4
X_49763_ _49757_/A _52979_/B _49763_/Y sky130_fd_sc_hd__nand2_4
X_46975_ _46975_/A _54473_/B sky130_fd_sc_hd__inv_2
X_42098_ _42097_/Y _88037_/D sky130_fd_sc_hd__inv_2
X_77795_ _77809_/A _77819_/A _77795_/X sky130_fd_sc_hd__xor2_4
X_48714_ _65425_/B _48150_/X _48713_/Y _48714_/Y sky130_fd_sc_hd__o21ai_4
X_79534_ _65397_/C _72465_/Y _79534_/Y sky130_fd_sc_hd__nand2_4
X_64760_ _64758_/X _83308_/Q _44171_/X _64759_/X _64760_/X sky130_fd_sc_hd__a211o_4
X_45926_ _64656_/A _45926_/X sky130_fd_sc_hd__buf_2
X_41049_ _41024_/X _81709_/Q _41048_/X _41050_/A sky130_fd_sc_hd__o21ai_4
X_76746_ _76746_/A _76746_/Y sky130_fd_sc_hd__inv_2
X_49694_ _49699_/A _47195_/X _49694_/Y sky130_fd_sc_hd__nand2_4
X_73958_ _73945_/X _73947_/X _73957_/X _73958_/X sky130_fd_sc_hd__a21o_4
X_61972_ _61957_/A _61967_/Y _61968_/Y _61971_/Y _61972_/Y sky130_fd_sc_hd__nand4_4
X_63711_ _63709_/Y _63679_/X _63710_/Y _63711_/Y sky130_fd_sc_hd__a21oi_4
X_48645_ _48845_/A _48657_/B _48657_/C _48645_/X sky130_fd_sc_hd__and3_4
X_60923_ _60918_/X _60921_/X _60994_/B _60923_/Y sky130_fd_sc_hd__o21ai_4
X_72909_ _72909_/A _72909_/X sky130_fd_sc_hd__buf_2
X_79465_ _58623_/Y _66389_/C _79464_/Y _79484_/A sky130_fd_sc_hd__o21a_4
X_45857_ _55219_/B _45740_/B _45857_/Y sky130_fd_sc_hd__nor2_4
X_64691_ _58124_/A _64691_/X sky130_fd_sc_hd__buf_2
X_76677_ _81685_/Q _81397_/Q _76969_/A sky130_fd_sc_hd__xnor2_4
X_73889_ _73887_/X _73888_/Y _73839_/X _73889_/X sky130_fd_sc_hd__a21o_4
X_66430_ _66427_/Y _66414_/X _66429_/Y _84125_/D sky130_fd_sc_hd__a21o_4
X_78416_ _78416_/A _82761_/D _82473_/D sky130_fd_sc_hd__xor2_4
X_44808_ _43896_/X _44808_/X sky130_fd_sc_hd__buf_2
X_63642_ _63638_/Y _63639_/Y _63641_/X _58465_/A _63363_/X _63642_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75628_ _75628_/A _75628_/B _80968_/D sky130_fd_sc_hd__xor2_4
X_48576_ _48576_/A _48565_/B _48576_/Y sky130_fd_sc_hd__nand2_4
X_60854_ _60853_/X _60854_/Y sky130_fd_sc_hd__inv_2
X_79396_ _79392_/X _79396_/B _79418_/B sky130_fd_sc_hd__xor2_4
X_45788_ _45785_/X _45787_/Y _45714_/X _45788_/Y sky130_fd_sc_hd__a21oi_4
X_47527_ _47526_/Y _53101_/B sky130_fd_sc_hd__buf_2
X_66361_ _65910_/X _66367_/B _65912_/X _66361_/Y sky130_fd_sc_hd__nand3_4
X_78347_ _78333_/Y _78329_/A _78332_/A _78347_/X sky130_fd_sc_hd__o21a_4
X_44739_ _49210_/A _50731_/B _40739_/A _44738_/Y _44736_/X _86980_/D
+ sky130_fd_sc_hd__o32ai_4
X_75559_ _80961_/D _75559_/B _75559_/X sky130_fd_sc_hd__xor2_4
X_63573_ _63573_/A _60712_/B _63630_/C _63573_/Y sky130_fd_sc_hd__nor3_4
X_60785_ _63384_/C _63384_/D _60694_/C _60660_/A _60785_/Y sky130_fd_sc_hd__nand4_4
X_68100_ _82079_/D _68040_/X _68099_/X _84039_/D sky130_fd_sc_hd__a21bo_4
X_65312_ _65305_/X _65833_/B _65311_/X _65312_/Y sky130_fd_sc_hd__nand3_4
X_62524_ _62623_/A _84892_/Q _62623_/C _62623_/D _62524_/X sky130_fd_sc_hd__and4_4
X_69080_ _69077_/X _69079_/X _69035_/X _69080_/X sky130_fd_sc_hd__a21o_4
X_47458_ _47458_/A _47459_/A sky130_fd_sc_hd__inv_2
X_66292_ _66231_/X _66319_/B _84143_/Q _66292_/X sky130_fd_sc_hd__and3_4
X_78278_ _78278_/A _78278_/B _78278_/X sky130_fd_sc_hd__xor2_4
X_68031_ _68405_/A _87190_/Q _68031_/X sky130_fd_sc_hd__and2_4
X_46409_ _46397_/Y _46399_/X _46408_/Y _46409_/Y sky130_fd_sc_hd__a21boi_4
X_65243_ _65198_/X _65233_/Y _65242_/Y _65243_/Y sky130_fd_sc_hd__o21ai_4
X_77229_ _77230_/A _77230_/C _77230_/B _77229_/Y sky130_fd_sc_hd__a21oi_4
X_62455_ _62411_/X _62412_/X _76985_/B _62455_/Y sky130_fd_sc_hd__nor3_4
X_47389_ _47198_/X _47418_/A sky130_fd_sc_hd__buf_2
X_61406_ _61406_/A _61404_/X _61406_/C _61390_/D _61406_/Y sky130_fd_sc_hd__nand4_4
X_49128_ _48946_/A _49128_/X sky130_fd_sc_hd__buf_2
X_80240_ _84952_/Q _65449_/C _80242_/A sky130_fd_sc_hd__xor2_4
X_65174_ _65172_/X _86123_/Q _65127_/X _65173_/X _65174_/X sky130_fd_sc_hd__a211o_4
X_62386_ _61483_/A _62332_/B _62386_/C _62332_/D _62389_/B sky130_fd_sc_hd__nand4_4
X_64125_ _62113_/X _64095_/B _64095_/C _64095_/D _64125_/Y sky130_fd_sc_hd__nand4_4
X_49059_ _48881_/X _81776_/Q _49058_/Y _49060_/A sky130_fd_sc_hd__o21ai_4
X_61337_ _72550_/C _61367_/D sky130_fd_sc_hd__buf_2
X_80171_ _80178_/B _80171_/B _80171_/X sky130_fd_sc_hd__xor2_4
X_69982_ _69588_/Y _69916_/X _69938_/X _69981_/Y _69982_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_7_72_0_CLK clkbuf_6_36_0_CLK/X clkbuf_7_72_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_52070_ _52070_/A _50370_/B _52070_/Y sky130_fd_sc_hd__nand2_4
X_64056_ _64054_/X _63994_/X _64055_/Y _64056_/Y sky130_fd_sc_hd__a21oi_4
X_68933_ _69567_/A _68933_/X sky130_fd_sc_hd__buf_2
X_61268_ _61262_/A _72544_/B _84493_/Q _61268_/Y sky130_fd_sc_hd__nor3_4
X_51021_ _51021_/A _51022_/A sky130_fd_sc_hd__buf_2
X_63007_ _63005_/Y _62987_/X _63006_/Y _84361_/D sky130_fd_sc_hd__a21oi_4
X_60219_ _60288_/C _60220_/A sky130_fd_sc_hd__buf_2
X_83930_ _83932_/CLK _69353_/X _83930_/Q sky130_fd_sc_hd__dfxtp_4
X_68864_ _68394_/A _68864_/X sky130_fd_sc_hd__buf_2
X_61199_ _72296_/A _66518_/B sky130_fd_sc_hd__buf_2
X_67815_ _67812_/X _67814_/X _67815_/Y sky130_fd_sc_hd__nand2_4
X_83861_ _82541_/CLK _70059_/X _82541_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_87_0_CLK clkbuf_7_87_0_CLK/A clkbuf_7_87_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_68795_ _68791_/X _68794_/X _68773_/X _68795_/X sky130_fd_sc_hd__a21o_4
X_85600_ _85601_/CLK _53625_/Y _85600_/Q sky130_fd_sc_hd__dfxtp_4
X_82812_ _84115_/CLK _82844_/Q _78689_/A sky130_fd_sc_hd__dfxtp_4
X_55760_ _55757_/X _55759_/X _55760_/Y sky130_fd_sc_hd__nand2_4
X_86580_ _86578_/CLK _47976_/Y _66097_/B sky130_fd_sc_hd__dfxtp_4
X_67746_ _67743_/X _67745_/X _67746_/Y sky130_fd_sc_hd__nand2_4
X_52972_ _52970_/Y _52946_/X _52971_/X _52972_/Y sky130_fd_sc_hd__a21oi_4
X_64958_ _64858_/X _85524_/Q _64859_/X _64957_/X _64958_/X sky130_fd_sc_hd__a211o_4
X_83792_ _81631_/CLK _83792_/D _74795_/A sky130_fd_sc_hd__dfxtp_4
X_54711_ _54656_/X _54734_/B sky130_fd_sc_hd__buf_2
X_85531_ _85822_/CLK _85531_/D _85531_/Q sky130_fd_sc_hd__dfxtp_4
X_51923_ _52021_/A _47830_/Y _51922_/X _51923_/Y sky130_fd_sc_hd__nand3_4
X_63909_ _64184_/A _63942_/A sky130_fd_sc_hd__buf_2
X_82743_ _82743_/CLK _66420_/C _79001_/A sky130_fd_sc_hd__dfxtp_4
X_55691_ _55691_/A _55698_/A sky130_fd_sc_hd__buf_2
X_67677_ _44020_/A _68451_/A sky130_fd_sc_hd__buf_2
X_64889_ _64880_/Y _64888_/Y _64889_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_7_10_0_CLK clkbuf_6_5_0_CLK/X clkbuf_8_21_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_57430_ _57430_/A _57413_/X _57430_/X sky130_fd_sc_hd__or2_4
X_69416_ _87019_/Q _69414_/X _69168_/X _69415_/X _69416_/X sky130_fd_sc_hd__a211o_4
X_88250_ _88247_/CLK _88250_/D _68984_/B sky130_fd_sc_hd__dfxtp_4
X_54642_ _85404_/Q _54621_/X _54641_/Y _54642_/Y sky130_fd_sc_hd__o21ai_4
X_66628_ _66572_/X _66628_/X sky130_fd_sc_hd__buf_2
X_85462_ _82769_/CLK _85462_/D _85462_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_150_0_CLK clkbuf_7_75_0_CLK/X clkbuf_8_150_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_51854_ _85934_/Q _51846_/X _51853_/Y _51854_/Y sky130_fd_sc_hd__o21ai_4
X_82674_ _81190_/CLK _82674_/D _78197_/A sky130_fd_sc_hd__dfxtp_4
X_87201_ _87720_/CLK _43915_/Y _87201_/Q sky130_fd_sc_hd__dfxtp_4
X_84413_ _84421_/CLK _84413_/D _62397_/C sky130_fd_sc_hd__dfxtp_4
X_50805_ _50505_/A _50806_/A sky130_fd_sc_hd__buf_2
X_57361_ _44231_/A _85028_/Q _57361_/Y sky130_fd_sc_hd__nand2_4
X_81625_ _81689_/CLK _76499_/X _81625_/Q sky130_fd_sc_hd__dfxtp_4
X_69347_ _69342_/X _69345_/X _69346_/X _69347_/X sky130_fd_sc_hd__a21o_4
X_88181_ _87926_/CLK _41623_/Y _88181_/Q sky130_fd_sc_hd__dfxtp_4
X_54573_ _54578_/A _53395_/B _54573_/Y sky130_fd_sc_hd__nand2_4
X_66559_ _66548_/X _66559_/B _66559_/Y sky130_fd_sc_hd__nand2_4
X_85393_ _85489_/CLK _54708_/Y _85393_/Q sky130_fd_sc_hd__dfxtp_4
X_51785_ _85946_/Q _51763_/X _51784_/Y _51785_/Y sky130_fd_sc_hd__o21ai_4
X_59100_ _59097_/Y _59099_/Y _59053_/X _59100_/X sky130_fd_sc_hd__a21o_4
X_56312_ _56351_/A _56312_/X sky130_fd_sc_hd__buf_2
X_87132_ _88215_/CLK _87132_/D _87132_/Q sky130_fd_sc_hd__dfxtp_4
X_53524_ _53696_/A _53524_/X sky130_fd_sc_hd__buf_2
X_84344_ _84344_/CLK _63211_/X _79330_/A sky130_fd_sc_hd__dfxtp_4
X_50736_ _50740_/A _53949_/B _50736_/Y sky130_fd_sc_hd__nand2_4
X_57292_ _56727_/X _57290_/X _57291_/Y _57292_/Y sky130_fd_sc_hd__o21ai_4
X_81556_ _84087_/CLK _76819_/X _81512_/D sky130_fd_sc_hd__dfxtp_4
X_69278_ _69183_/A _69278_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_25_0_CLK clkbuf_6_12_0_CLK/X clkbuf_8_51_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_59031_ _58923_/A _59031_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_165_0_CLK clkbuf_7_82_0_CLK/X clkbuf_9_331_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_56243_ _56250_/A _56243_/B _56243_/C _56243_/Y sky130_fd_sc_hd__nand3_4
X_80507_ _80505_/X _80506_/X _80520_/B sky130_fd_sc_hd__xnor2_4
X_68229_ _67419_/X _67422_/X _68216_/X _68229_/Y sky130_fd_sc_hd__a21oi_4
X_87063_ _87063_/CLK _44538_/Y _72973_/A sky130_fd_sc_hd__dfxtp_4
X_53455_ _53455_/A _53455_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_160_0_CLK clkbuf_9_80_0_CLK/X _81801_/CLK sky130_fd_sc_hd__clkbuf_1
X_84275_ _84273_/CLK _64101_/Y _64100_/C sky130_fd_sc_hd__dfxtp_4
X_50667_ _86157_/Q _50654_/X _50666_/Y _50667_/Y sky130_fd_sc_hd__o21ai_4
X_81487_ _81333_/CLK _84055_/Q _81487_/Q sky130_fd_sc_hd__dfxtp_4
X_86014_ _85727_/CLK _86014_/D _86014_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_790_0_CLK clkbuf_9_395_0_CLK/X _82147_/CLK sky130_fd_sc_hd__clkbuf_1
X_40420_ _40420_/A _47867_/A sky130_fd_sc_hd__buf_2
X_52406_ _65324_/B _52397_/X _52405_/Y _52406_/Y sky130_fd_sc_hd__o21ai_4
X_71240_ _71238_/B _71241_/A sky130_fd_sc_hd__inv_2
X_83226_ _83227_/CLK _83226_/D _79352_/B sky130_fd_sc_hd__dfxtp_4
X_56174_ _56173_/Y _56174_/X sky130_fd_sc_hd__buf_2
X_80438_ _80435_/X _80437_/Y _80438_/Y sky130_fd_sc_hd__xnor2_4
X_53386_ _53386_/A _53386_/B _53386_/Y sky130_fd_sc_hd__nand2_4
X_50598_ _86170_/Q _50594_/X _50597_/Y _50598_/Y sky130_fd_sc_hd__o21ai_4
X_55125_ _55125_/A _55126_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_281_0_CLK clkbuf_9_281_0_CLK/A clkbuf_9_281_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_40351_ _42447_/C _42447_/A _41869_/C _40351_/Y sky130_fd_sc_hd__nor3_4
X_52337_ _52335_/Y _52314_/X _52336_/X _52337_/Y sky130_fd_sc_hd__a21oi_4
X_71171_ _71171_/A _71173_/B _71181_/C _71178_/D _71171_/Y sky130_fd_sc_hd__nand4_4
X_83157_ _85895_/CLK _73295_/X _83157_/Q sky130_fd_sc_hd__dfxtp_4
X_80369_ _80368_/Y _80383_/B sky130_fd_sc_hd__inv_2
X_70122_ _83142_/Q _70122_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_175_0_CLK clkbuf_9_87_0_CLK/X _80784_/CLK sky130_fd_sc_hd__clkbuf_1
X_82108_ _82015_/CLK _82108_/D _82108_/Q sky130_fd_sc_hd__dfxtp_4
X_43070_ _43070_/A _43070_/Y sky130_fd_sc_hd__inv_2
X_55056_ _47918_/A _55056_/X sky130_fd_sc_hd__buf_2
X_59933_ _59927_/A _59973_/A sky130_fd_sc_hd__buf_2
X_52268_ _52266_/Y _52262_/X _52267_/X _52268_/Y sky130_fd_sc_hd__a21oi_4
X_87965_ _87644_/CLK _87965_/D _87965_/Q sky130_fd_sc_hd__dfxtp_4
X_83088_ _83187_/CLK _74350_/X _83088_/Q sky130_fd_sc_hd__dfxtp_4
X_42021_ _41998_/X _42010_/X _40845_/X _42020_/Y _42000_/X _42021_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54007_ _53998_/A _46407_/X _54007_/Y sky130_fd_sc_hd__nand2_4
X_51219_ _51218_/X _51220_/A sky130_fd_sc_hd__buf_2
X_74930_ _74930_/A _74929_/X _74930_/Y sky130_fd_sc_hd__nand2_4
X_70053_ _69825_/X _69827_/X _69994_/X _70053_/X sky130_fd_sc_hd__a21o_4
X_86916_ _88215_/CLK _86916_/D _67988_/B sky130_fd_sc_hd__dfxtp_4
X_82039_ _82008_/CLK _82039_/D _82007_/D sky130_fd_sc_hd__dfxtp_4
X_59864_ _59873_/A _59855_/B _80308_/B _59864_/Y sky130_fd_sc_hd__nor3_4
X_52199_ _52199_/A _52198_/X _52218_/C _52199_/X sky130_fd_sc_hd__and3_4
X_87896_ _86914_/CLK _87896_/D _87896_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_296_0_CLK clkbuf_9_296_0_CLK/A clkbuf_9_296_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_58815_ _58787_/X _86094_/Q _58814_/X _58815_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_8_103_0_CLK clkbuf_7_51_0_CLK/X clkbuf_9_206_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_74861_ _74857_/Y _74860_/Y _74863_/B sky130_fd_sc_hd__xnor2_4
X_86847_ _81117_/CLK _86847_/D _41869_/A sky130_fd_sc_hd__dfxtp_4
X_59795_ _59737_/A _59848_/B _80475_/A _59795_/Y sky130_fd_sc_hd__nor3_4
X_76600_ _76599_/X _76602_/B sky130_fd_sc_hd__inv_2
X_73812_ _73812_/A _73812_/B _73813_/B sky130_fd_sc_hd__nand2_4
X_46760_ _86706_/Q _46719_/X _46759_/Y _46760_/Y sky130_fd_sc_hd__o21ai_4
X_58746_ _44170_/A _64600_/A sky130_fd_sc_hd__buf_2
X_77580_ _77580_/A _77584_/A sky130_fd_sc_hd__inv_2
X_43972_ _80667_/Q _43972_/B _43972_/Y sky130_fd_sc_hd__nor2_4
X_55958_ _55695_/A _55958_/B _55958_/X sky130_fd_sc_hd__and2_4
X_74792_ _74734_/Y _83847_/Q _74789_/X _74790_/X _74791_/X _74792_/X
+ sky130_fd_sc_hd__a2111o_4
X_86778_ _86814_/CLK _46078_/Y _86778_/Q sky130_fd_sc_hd__dfxtp_4
X_45711_ _82989_/Q _45713_/A sky130_fd_sc_hd__inv_2
X_76531_ _81660_/Q _76531_/Y sky130_fd_sc_hd__inv_2
X_42923_ _41715_/X _42920_/X _67714_/B _42922_/X _87651_/D sky130_fd_sc_hd__a2bb2o_4
X_54909_ _54882_/A _54909_/X sky130_fd_sc_hd__buf_2
X_73743_ _73665_/X _84986_/Q _73740_/X _73742_/X _73743_/X sky130_fd_sc_hd__a211o_4
X_85729_ _83690_/CLK _85729_/D _85729_/Q sky130_fd_sc_hd__dfxtp_4
X_70955_ _50757_/B _70936_/X _70954_/Y _70955_/Y sky130_fd_sc_hd__o21ai_4
X_58677_ _58677_/A _58688_/B _58677_/Y sky130_fd_sc_hd__nor2_4
X_46691_ _46687_/Y _46654_/X _46690_/X _86714_/D sky130_fd_sc_hd__a21oi_4
X_55889_ _55903_/A _55889_/B _55889_/X sky130_fd_sc_hd__and2_4
Xclkbuf_8_118_0_CLK clkbuf_7_59_0_CLK/X clkbuf_8_118_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_48430_ _48545_/A _48476_/C sky130_fd_sc_hd__buf_2
X_79250_ _79250_/A _79250_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_113_0_CLK clkbuf_9_56_0_CLK/X _83242_/CLK sky130_fd_sc_hd__clkbuf_1
X_57628_ _57608_/X _50372_/B _57628_/Y sky130_fd_sc_hd__nand2_4
X_45642_ _45635_/X _45639_/Y _45641_/Y _45642_/Y sky130_fd_sc_hd__a21oi_4
X_76462_ _76461_/X _76482_/B sky130_fd_sc_hd__inv_2
X_42854_ _41525_/X _42852_/X _66876_/B _42853_/X _87686_/D sky130_fd_sc_hd__a2bb2o_4
X_73674_ _73250_/A _73674_/X sky130_fd_sc_hd__buf_2
X_70886_ _70886_/A _70882_/Y _70905_/D sky130_fd_sc_hd__nor2_4
Xclkbuf_10_743_0_CLK clkbuf_9_371_0_CLK/X _87235_/CLK sky130_fd_sc_hd__clkbuf_1
X_78201_ _78204_/B _78200_/Y _78202_/B sky130_fd_sc_hd__xnor2_4
X_75413_ _75413_/A _75413_/B _75413_/C _75413_/X sky130_fd_sc_hd__or3_4
X_41805_ _41805_/A _41805_/Y sky130_fd_sc_hd__inv_2
X_48361_ _48044_/A _48361_/B _48361_/Y sky130_fd_sc_hd__nand2_4
X_72625_ _72625_/A _72625_/B _72625_/X sky130_fd_sc_hd__and2_4
X_79181_ _84788_/Q _84108_/Q _79181_/Y sky130_fd_sc_hd__nand2_4
X_45573_ _55508_/B _45570_/X _45571_/X _45572_/Y _45573_/X sky130_fd_sc_hd__a211o_4
X_57559_ _84979_/Q _57550_/X _57558_/Y _57559_/Y sky130_fd_sc_hd__o21ai_4
X_76393_ _76393_/A _81567_/Q _76394_/A sky130_fd_sc_hd__nand2_4
X_88379_ _87417_/CLK _88379_/D _88379_/Q sky130_fd_sc_hd__dfxtp_4
X_42785_ _42785_/A _87720_/D sky130_fd_sc_hd__inv_2
X_47312_ _47308_/Y _47271_/X _47311_/X _86648_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_234_0_CLK clkbuf_9_235_0_CLK/A clkbuf_9_234_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_78132_ _78130_/C _78130_/D _78132_/Y sky130_fd_sc_hd__nand2_4
X_44524_ _44496_/X _44497_/X _40787_/X _87067_/Q _44498_/X _44524_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75344_ _75308_/Y _75342_/X _75343_/Y _75345_/B sky130_fd_sc_hd__a21oi_4
X_41736_ _41607_/X _41736_/X sky130_fd_sc_hd__buf_2
X_60570_ _60570_/A _60570_/B _60570_/C _60570_/X sky130_fd_sc_hd__and3_4
X_48292_ _48290_/Y _48233_/X _48291_/X _86541_/D sky130_fd_sc_hd__a21oi_4
X_72556_ _72572_/A _72556_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_128_0_CLK clkbuf_9_64_0_CLK/X _81807_/CLK sky130_fd_sc_hd__clkbuf_1
X_47243_ _54102_/B _52936_/B sky130_fd_sc_hd__buf_2
X_71507_ _71507_/A _71507_/B _71525_/A sky130_fd_sc_hd__nor2_4
X_59229_ _59229_/A _59229_/Y sky130_fd_sc_hd__inv_2
X_78063_ _84568_/Q _78063_/B _78063_/X sky130_fd_sc_hd__xor2_4
X_44455_ _41121_/A _44453_/X _87102_/Q _44454_/X _44455_/X sky130_fd_sc_hd__a2bb2o_4
X_75275_ _75271_/X _75272_/Y _75274_/Y _75277_/A sky130_fd_sc_hd__a21o_4
X_41667_ _41666_/X _41667_/X sky130_fd_sc_hd__buf_2
X_72487_ _72484_/X _83385_/Q _72486_/Y _83249_/D sky130_fd_sc_hd__o21a_4
Xclkbuf_10_758_0_CLK clkbuf_9_379_0_CLK/X _87533_/CLK sky130_fd_sc_hd__clkbuf_1
X_77014_ _77004_/Y _77012_/Y _77013_/Y _77014_/Y sky130_fd_sc_hd__o21ai_4
X_43406_ _43405_/Y _43406_/Y sky130_fd_sc_hd__inv_2
X_62240_ _62220_/X _62234_/Y _62239_/X _58149_/A _62214_/X _62240_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74226_ _74226_/A _74073_/X _74226_/Y sky130_fd_sc_hd__nor2_4
X_40618_ _40617_/X _40596_/X _88365_/Q _40599_/X _40618_/X sky130_fd_sc_hd__a2bb2o_4
X_47174_ _54587_/B _47174_/X sky130_fd_sc_hd__buf_2
X_71438_ _71419_/Y _83499_/Q _71437_/X _71438_/X sky130_fd_sc_hd__a21o_4
X_44386_ _44381_/X _44382_/X _41791_/X _87136_/Q _44383_/X _44387_/A
+ sky130_fd_sc_hd__o32ai_4
X_41598_ _41597_/Y _88185_/D sky130_fd_sc_hd__inv_2
Xclkbuf_9_249_0_CLK clkbuf_8_124_0_CLK/X clkbuf_9_249_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_46125_ _46125_/A _46195_/A sky130_fd_sc_hd__buf_2
X_43337_ _43302_/A _43337_/X sky130_fd_sc_hd__buf_2
X_62171_ _58210_/X _62105_/X _62065_/D _62055_/A _62170_/X _62171_/X
+ sky130_fd_sc_hd__a41o_4
X_74157_ _74237_/A _86536_/Q _74157_/X sky130_fd_sc_hd__and2_4
X_40549_ _40548_/X _40543_/X _88372_/Q _40544_/X _40549_/X sky130_fd_sc_hd__a2bb2o_4
X_71369_ _71366_/A _70939_/A _71439_/C _71365_/X _71369_/X sky130_fd_sc_hd__and4_4
X_61122_ _61122_/A _61122_/B _61122_/C _64421_/A sky130_fd_sc_hd__and3_4
X_73108_ _73108_/A _44127_/X _73108_/Y sky130_fd_sc_hd__nor2_4
X_46056_ _46055_/Y _86791_/D sky130_fd_sc_hd__inv_2
X_43268_ _41108_/X _43264_/X _87508_/Q _43265_/X _43268_/X sky130_fd_sc_hd__a2bb2o_4
X_74088_ _73588_/A _86539_/Q _74088_/X sky130_fd_sc_hd__and2_4
X_78965_ _78965_/A _78965_/B _78965_/X sky130_fd_sc_hd__xor2_4
X_45007_ _45007_/A _45033_/B _45007_/Y sky130_fd_sc_hd__nand2_4
X_42219_ _41356_/X _42209_/X _87974_/Q _42210_/X _87974_/D sky130_fd_sc_hd__a2bb2o_4
X_65930_ _65916_/A _65970_/B _84168_/Q _65930_/X sky130_fd_sc_hd__and3_4
X_61053_ _60946_/X _61138_/B _76975_/A _61053_/Y sky130_fd_sc_hd__nor3_4
X_77916_ _77916_/A _77916_/B _82038_/D sky130_fd_sc_hd__xor2_4
X_73039_ _73024_/Y _73029_/Y _73038_/X _73039_/Y sky130_fd_sc_hd__o21ai_4
X_43199_ _43199_/A _43199_/Y sky130_fd_sc_hd__inv_2
X_78896_ _78896_/A _82506_/D sky130_fd_sc_hd__inv_2
X_60004_ _63055_/A _65842_/A sky130_fd_sc_hd__buf_2
X_49815_ _49787_/A _49815_/X sky130_fd_sc_hd__buf_2
X_65861_ _65807_/A _86468_/Q _65861_/X sky130_fd_sc_hd__and2_4
X_77847_ _77847_/A _77833_/Y _77847_/Y sky130_fd_sc_hd__nor2_4
X_67600_ _67696_/A _67600_/B _67600_/X sky130_fd_sc_hd__and2_4
X_64812_ _64808_/X _64937_/B _64811_/X _64812_/Y sky130_fd_sc_hd__nand3_4
X_49746_ _49751_/A _49724_/B _49761_/C _52963_/D _49746_/X sky130_fd_sc_hd__and4_4
X_68580_ _68059_/A _68580_/X sky130_fd_sc_hd__buf_2
X_46958_ _54464_/B _52773_/B sky130_fd_sc_hd__buf_2
X_65792_ _65804_/A _85865_/Q _65792_/X sky130_fd_sc_hd__and2_4
X_77778_ _77780_/B _81927_/D _77778_/X sky130_fd_sc_hd__or2_4
X_67531_ _86967_/Q _67432_/X _67433_/X _67530_/X _67531_/X sky130_fd_sc_hd__a211o_4
X_79517_ _79517_/A _79517_/B _79518_/B sky130_fd_sc_hd__xor2_4
X_45909_ _45909_/A _45909_/X sky130_fd_sc_hd__buf_2
X_64743_ _64676_/A _64743_/B _64743_/X sky130_fd_sc_hd__and2_4
X_76729_ _76727_/Y _76728_/Y _76732_/A sky130_fd_sc_hd__xor2_4
X_61955_ _61777_/A _61971_/C sky130_fd_sc_hd__buf_2
X_49677_ _49570_/A _49677_/X sky130_fd_sc_hd__buf_2
X_46889_ _58942_/A _46859_/X _46888_/Y _46889_/Y sky130_fd_sc_hd__o21ai_4
X_60906_ _60892_/Y _60906_/X sky130_fd_sc_hd__buf_2
X_48628_ _48661_/A _48628_/B _48628_/Y sky130_fd_sc_hd__nand2_4
X_79448_ _79446_/X _79453_/B _79448_/Y sky130_fd_sc_hd__xnor2_4
X_67462_ _67226_/A _67462_/X sky130_fd_sc_hd__buf_2
X_64674_ _64577_/X _86750_/Q _64579_/X _64673_/X _64674_/X sky130_fd_sc_hd__a211o_4
X_61886_ _61871_/A _61839_/B _61839_/C _63124_/B _61886_/X sky130_fd_sc_hd__and4_4
X_69201_ _81405_/D _69161_/X _69200_/X _83941_/D sky130_fd_sc_hd__a21bo_4
X_66413_ _66411_/X _66043_/Y _66412_/Y _66413_/Y sky130_fd_sc_hd__o21ai_4
X_63625_ _63655_/A _58495_/A _63581_/X _63595_/D _63625_/X sky130_fd_sc_hd__and4_4
X_48559_ _48559_/A _48559_/Y sky130_fd_sc_hd__inv_2
X_60837_ _60376_/X _60834_/X _60804_/Y _60799_/X _60836_/X _84555_/D
+ sky130_fd_sc_hd__o41a_4
X_67393_ _87985_/Q _67293_/X _67391_/X _67392_/X _67393_/X sky130_fd_sc_hd__a211o_4
X_79379_ _79366_/X _79377_/X _79378_/X _79379_/Y sky130_fd_sc_hd__a21oi_4
X_81410_ _84079_/CLK _81442_/Q _75924_/B sky130_fd_sc_hd__dfxtp_4
X_69132_ _68907_/X _69109_/X _69120_/Y _69131_/Y _69132_/X sky130_fd_sc_hd__a211o_4
X_66344_ _84139_/Q _66345_/C sky130_fd_sc_hd__inv_2
X_51570_ _51553_/A _51580_/B _51553_/C _53099_/D _51570_/X sky130_fd_sc_hd__and4_4
X_63556_ _63368_/A _63556_/X sky130_fd_sc_hd__buf_2
X_82390_ _82390_/CLK _82390_/D _82390_/Q sky130_fd_sc_hd__dfxtp_4
X_60768_ _60610_/A _60513_/B _78066_/A _60768_/X sky130_fd_sc_hd__or3_4
X_50521_ _50513_/A _48843_/B _50521_/Y sky130_fd_sc_hd__nand2_4
X_81341_ _81330_/CLK _81341_/D _81717_/D sky130_fd_sc_hd__dfxtp_4
X_62507_ _59950_/C _62507_/X sky130_fd_sc_hd__buf_2
X_69063_ _69050_/Y _68823_/X _68824_/X _69062_/Y _69063_/X sky130_fd_sc_hd__a211o_4
X_66275_ _66272_/X _66274_/X _66275_/Y sky130_fd_sc_hd__nand2_4
X_63487_ _63487_/A _63487_/X sky130_fd_sc_hd__buf_2
X_60699_ _60558_/X _60700_/A sky130_fd_sc_hd__buf_2
X_68014_ _87139_/Q _67942_/X _67991_/X _68013_/X _68014_/X sky130_fd_sc_hd__a211o_4
X_53240_ _53246_/A _53240_/B _53240_/Y sky130_fd_sc_hd__nand2_4
X_65226_ _65199_/X _86153_/Q _65224_/X _65225_/X _65226_/X sky130_fd_sc_hd__a211o_4
X_84060_ _81749_/CLK _67663_/X _81492_/D sky130_fd_sc_hd__dfxtp_4
X_50452_ _50450_/Y _50429_/X _50451_/X _50452_/Y sky130_fd_sc_hd__a21oi_4
X_62438_ _62479_/A _61969_/X _62479_/C _62392_/D _62438_/X sky130_fd_sc_hd__and4_4
X_81272_ _81697_/CLK _81304_/Q _81272_/Q sky130_fd_sc_hd__dfxtp_4
X_83011_ _83012_/CLK _74624_/Y _83011_/Q sky130_fd_sc_hd__dfxtp_4
X_80223_ _80204_/Y _80207_/Y _80225_/B sky130_fd_sc_hd__or2_4
X_53171_ _53168_/Y _53163_/X _53170_/X _85684_/D sky130_fd_sc_hd__a21oi_4
X_65157_ _64717_/A _65158_/A sky130_fd_sc_hd__buf_2
X_50383_ _50383_/A _50383_/B _50383_/Y sky130_fd_sc_hd__nand2_4
X_62369_ _62342_/A _62341_/X _84415_/Q _62369_/Y sky130_fd_sc_hd__nor3_4
X_52122_ _65501_/B _52075_/X _52121_/Y _52122_/Y sky130_fd_sc_hd__o21ai_4
X_64108_ _64116_/A _64087_/X _64108_/C _64108_/Y sky130_fd_sc_hd__nor3_4
X_80154_ _80154_/A _80153_/X _80169_/B sky130_fd_sc_hd__xnor2_4
X_65088_ _65065_/X _83295_/Q _64991_/X _65087_/X _65088_/X sky130_fd_sc_hd__a211o_4
X_69965_ _69943_/X _46199_/X _69963_/Y _69964_/Y _69965_/X sky130_fd_sc_hd__a211o_4
X_52053_ _74104_/B _52041_/X _52052_/Y _52053_/Y sky130_fd_sc_hd__o21ai_4
X_56930_ _56953_/A _56930_/X sky130_fd_sc_hd__buf_2
X_68916_ _69478_/A _68916_/X sky130_fd_sc_hd__buf_2
X_64039_ _63751_/X _64142_/D sky130_fd_sc_hd__buf_2
X_87750_ _88006_/CLK _87750_/D _87750_/Q sky130_fd_sc_hd__dfxtp_4
X_84962_ _86210_/CLK _84962_/D _84962_/Q sky130_fd_sc_hd__dfxtp_4
X_80085_ _80071_/A _80070_/Y _80085_/X sky130_fd_sc_hd__or2_4
X_69896_ _43190_/A _69833_/X _68348_/X _69895_/X _69896_/X sky130_fd_sc_hd__a211o_4
X_51004_ _86091_/Q _50992_/X _51003_/Y _51004_/Y sky130_fd_sc_hd__o21ai_4
X_86701_ _86701_/CLK _86701_/D _86701_/Q sky130_fd_sc_hd__dfxtp_4
X_83913_ _81985_/CLK _83913_/D _81985_/D sky130_fd_sc_hd__dfxtp_4
X_56861_ _56675_/X _56893_/B sky130_fd_sc_hd__buf_2
X_68847_ _68843_/X _68845_/X _68846_/X _68847_/Y sky130_fd_sc_hd__a21oi_4
X_87681_ _82888_/CLK _42862_/X _87681_/Q sky130_fd_sc_hd__dfxtp_4
X_84893_ _84250_/CLK _84893_/D _58264_/A sky130_fd_sc_hd__dfxtp_4
X_58600_ _58687_/A _86398_/Q _58600_/Y sky130_fd_sc_hd__nor2_4
X_55812_ _44077_/X _56339_/C _55812_/X sky130_fd_sc_hd__and2_4
X_86632_ _85993_/CLK _47467_/Y _86632_/Q sky130_fd_sc_hd__dfxtp_4
X_59580_ _59557_/A _59516_/A _59581_/C _59582_/A sky130_fd_sc_hd__nand3_4
X_83844_ _83835_/CLK _83844_/D _83844_/Q sky130_fd_sc_hd__dfxtp_4
X_56792_ _46159_/A _55176_/Y _56791_/Y _56792_/X sky130_fd_sc_hd__o21a_4
X_68778_ _69007_/A _68778_/X sky130_fd_sc_hd__buf_2
X_58531_ _84826_/Q _58533_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_1000_0_CLK clkbuf_9_500_0_CLK/X _85888_/CLK sky130_fd_sc_hd__clkbuf_1
X_55743_ _55742_/X _55743_/Y sky130_fd_sc_hd__inv_2
X_67729_ _67678_/X _67729_/B _67729_/X sky130_fd_sc_hd__and2_4
X_86563_ _85888_/CLK _86563_/D _86563_/Q sky130_fd_sc_hd__dfxtp_4
X_52955_ _52951_/Y _52946_/X _52954_/X _85724_/D sky130_fd_sc_hd__a21oi_4
X_83775_ _86553_/CLK _83775_/D _83775_/Q sky130_fd_sc_hd__dfxtp_4
X_80987_ _80818_/CLK _80987_/D _80943_/D sky130_fd_sc_hd__dfxtp_4
X_88302_ _86989_/CLK _88302_/D _69209_/B sky130_fd_sc_hd__dfxtp_4
X_85514_ _85514_/CLK _85514_/D _85514_/Q sky130_fd_sc_hd__dfxtp_4
X_51906_ _51903_/Y _51904_/X _51905_/X _51906_/Y sky130_fd_sc_hd__a21oi_4
X_70740_ _70740_/A _70585_/X _70740_/Y sky130_fd_sc_hd__nand2_4
X_58462_ _58448_/X _83475_/Q _58461_/Y _84843_/D sky130_fd_sc_hd__o21a_4
X_82726_ _81190_/CLK _84110_/Q _82726_/Q sky130_fd_sc_hd__dfxtp_4
X_55674_ _55674_/A _55674_/B _55675_/B sky130_fd_sc_hd__nand2_4
X_86494_ _86203_/CLK _86494_/D _72840_/B sky130_fd_sc_hd__dfxtp_4
X_52886_ _85736_/Q _52874_/X _52885_/Y _52886_/Y sky130_fd_sc_hd__o21ai_4
X_57413_ _44037_/X _57413_/X sky130_fd_sc_hd__buf_2
X_88233_ _88224_/CLK _41343_/Y _88233_/Q sky130_fd_sc_hd__dfxtp_4
X_54625_ _54625_/A _54607_/B _54618_/X _47236_/A _54625_/X sky130_fd_sc_hd__and4_4
X_85445_ _85767_/CLK _54424_/Y _85445_/Q sky130_fd_sc_hd__dfxtp_4
X_51837_ _51781_/A _51851_/C sky130_fd_sc_hd__buf_2
X_70671_ _70664_/X _83729_/Q _70670_/Y _70671_/X sky130_fd_sc_hd__a21o_4
X_58393_ _84860_/Q _58393_/Y sky130_fd_sc_hd__inv_2
X_82657_ _84014_/CLK _82657_/D _82657_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_1015_0_CLK clkbuf_9_507_0_CLK/X _85571_/CLK sky130_fd_sc_hd__clkbuf_1
X_72410_ _72352_/X _85961_/Q _72409_/X _72410_/Y sky130_fd_sc_hd__o21ai_4
X_57344_ _57344_/A _57344_/Y sky130_fd_sc_hd__inv_2
X_81608_ _81582_/CLK _81608_/D _81800_/D sky130_fd_sc_hd__dfxtp_4
X_88164_ _88164_/CLK _41712_/Y _88164_/Q sky130_fd_sc_hd__dfxtp_4
X_42570_ _87816_/Q _69710_/B sky130_fd_sc_hd__inv_2
X_54556_ _85420_/Q _54540_/X _54555_/Y _54556_/Y sky130_fd_sc_hd__o21ai_4
X_85376_ _83711_/CLK _54799_/Y _85376_/Q sky130_fd_sc_hd__dfxtp_4
X_73390_ _73377_/Y _73389_/X _73391_/B sky130_fd_sc_hd__xnor2_4
X_51768_ _51768_/A _51782_/B _51755_/X _51768_/D _51768_/X sky130_fd_sc_hd__and4_4
X_82588_ _82589_/CLK _82620_/Q _78262_/A sky130_fd_sc_hd__dfxtp_4
X_87115_ _87684_/CLK _87115_/D _87115_/Q sky130_fd_sc_hd__dfxtp_4
X_41521_ _41489_/X _41490_/X _41520_/X _66857_/B _41474_/X _41522_/A
+ sky130_fd_sc_hd__o32ai_4
X_53507_ _53817_/A _53723_/A sky130_fd_sc_hd__buf_2
X_72341_ _72305_/X _85359_/Q _72340_/X _72341_/Y sky130_fd_sc_hd__o21ai_4
X_84327_ _84355_/CLK _63393_/Y _63392_/C sky130_fd_sc_hd__dfxtp_4
X_50719_ _50740_/A _50719_/B _50719_/Y sky130_fd_sc_hd__nand2_4
X_57275_ _44207_/A _57275_/X sky130_fd_sc_hd__buf_2
X_81539_ _81351_/CLK _81539_/D _81539_/Q sky130_fd_sc_hd__dfxtp_4
X_88095_ _88111_/CLK _41950_/Y _74031_/A sky130_fd_sc_hd__dfxtp_4
X_54487_ _54486_/X _53309_/B _54487_/Y sky130_fd_sc_hd__nand2_4
X_51699_ _51695_/A _51715_/B _51695_/C _53223_/D _51699_/X sky130_fd_sc_hd__and4_4
X_59014_ _59013_/X _85760_/Q _58928_/X _59014_/X sky130_fd_sc_hd__o21a_4
X_44240_ _44226_/Y _44232_/Y _44256_/A _87179_/D sky130_fd_sc_hd__a21oi_4
X_56226_ _56252_/A _56233_/A sky130_fd_sc_hd__buf_2
X_75060_ _80959_/Q _75059_/X _75060_/X sky130_fd_sc_hd__xor2_4
X_41452_ _41452_/A _41459_/B _41452_/X sky130_fd_sc_hd__or2_4
X_87046_ _87285_/CLK _87046_/D _87046_/Q sky130_fd_sc_hd__dfxtp_4
X_53438_ _53357_/A _54111_/C sky130_fd_sc_hd__buf_2
X_72272_ _72366_/A _86293_/Q _72272_/Y sky130_fd_sc_hd__nor2_4
X_84258_ _83402_/CLK _84258_/D _79806_/B sky130_fd_sc_hd__dfxtp_4
X_74011_ _44719_/Y _56183_/X _74010_/Y _74028_/C sky130_fd_sc_hd__a21o_4
X_40403_ _40325_/X _82330_/Q _40402_/X _40403_/Y sky130_fd_sc_hd__o21ai_4
X_71223_ _71232_/A _71223_/B _71219_/C _71223_/Y sky130_fd_sc_hd__nand3_4
X_83209_ _83095_/CLK _72636_/X _70165_/A sky130_fd_sc_hd__dfxtp_4
X_44171_ _65768_/A _44171_/X sky130_fd_sc_hd__buf_2
X_56157_ _56163_/A _56167_/B _56167_/A _56157_/Y sky130_fd_sc_hd__nand3_4
X_41383_ _41337_/X _41338_/X _41382_/X _67767_/B _41333_/X _41383_/Y
+ sky130_fd_sc_hd__o32ai_4
X_53369_ _53353_/A _53369_/B _53369_/Y sky130_fd_sc_hd__nand2_4
X_84189_ _84192_/CLK _84189_/D _84189_/Q sky130_fd_sc_hd__dfxtp_4
X_43122_ _43100_/X _43110_/X _40787_/X _72859_/A _43121_/X _43123_/A
+ sky130_fd_sc_hd__o32ai_4
X_55108_ _55112_/A _47877_/A _55120_/C _47794_/A _55108_/X sky130_fd_sc_hd__and4_4
X_40334_ _86757_/Q _40335_/B sky130_fd_sc_hd__inv_2
X_71154_ _70716_/A _71160_/C sky130_fd_sc_hd__buf_2
X_56088_ _56088_/A _55842_/X _56088_/X sky130_fd_sc_hd__and2_4
X_70105_ _83137_/Q _70107_/C sky130_fd_sc_hd__inv_2
X_47930_ _83776_/Q _53501_/B sky130_fd_sc_hd__inv_2
X_55039_ _55017_/X _55030_/X _55026_/C _47675_/A _55039_/X sky130_fd_sc_hd__and4_4
X_59916_ _59660_/C _60620_/C _59660_/D _60620_/B _60155_/C sky130_fd_sc_hd__and4_4
X_43053_ _43129_/A _43053_/X sky130_fd_sc_hd__buf_2
X_78750_ _78750_/A _82687_/D _78753_/B sky130_fd_sc_hd__nor2_4
X_71085_ _70819_/A _71230_/B sky130_fd_sc_hd__buf_2
X_75962_ _75956_/Y _75963_/C _75961_/Y _75964_/A sky130_fd_sc_hd__a21o_4
X_87948_ _87952_/CLK _42269_/Y _87948_/Q sky130_fd_sc_hd__dfxtp_4
X_42004_ _88074_/Q _42004_/Y sky130_fd_sc_hd__inv_2
X_77701_ _77701_/A _77700_/X _77702_/A sky130_fd_sc_hd__xor2_4
X_74913_ _74905_/A _74910_/A _74914_/B sky130_fd_sc_hd__and2_4
X_70036_ _82547_/D _70029_/X _70035_/X _70036_/X sky130_fd_sc_hd__a21bo_4
X_47861_ _47887_/A _47861_/B _47861_/X sky130_fd_sc_hd__and2_4
X_59847_ _43969_/A _59741_/A _59581_/C _43969_/B _59846_/X _59847_/Y
+ sky130_fd_sc_hd__a41oi_4
X_78681_ _78680_/Y _78682_/C sky130_fd_sc_hd__inv_2
X_75893_ _84491_/Q _62988_/C _75893_/X sky130_fd_sc_hd__xor2_4
X_87879_ _87883_/CLK _42405_/Y _87879_/Q sky130_fd_sc_hd__dfxtp_4
X_49600_ _49580_/X _52813_/B _49600_/Y sky130_fd_sc_hd__nand2_4
X_46812_ _46807_/Y _46798_/X _46811_/X _86701_/D sky130_fd_sc_hd__a21oi_4
X_77632_ _77632_/A _77632_/Y sky130_fd_sc_hd__inv_2
X_74844_ _74844_/A _46099_/X _74844_/Y sky130_fd_sc_hd__nand2_4
X_47792_ _47792_/A _49364_/B sky130_fd_sc_hd__buf_2
X_59778_ _59772_/A _59837_/B _80506_/A _59778_/Y sky130_fd_sc_hd__nor3_4
X_49531_ _58957_/B _49524_/X _49530_/Y _49531_/Y sky130_fd_sc_hd__o21ai_4
X_46743_ _82964_/Q _46743_/Y sky130_fd_sc_hd__inv_2
X_58729_ _58696_/X _58726_/Y _58727_/Y _58728_/X _58701_/X _58729_/X
+ sky130_fd_sc_hd__o32a_4
X_77563_ _77526_/Y _77561_/X _77562_/Y _77564_/B sky130_fd_sc_hd__a21oi_4
X_43955_ _80669_/Q _43955_/Y sky130_fd_sc_hd__inv_2
X_74775_ _74775_/A _74775_/B _71846_/A _70500_/B _74775_/X sky130_fd_sc_hd__and4_4
X_71987_ _72007_/A _71987_/B _71987_/Y sky130_fd_sc_hd__nand2_4
X_79302_ _79302_/A _79301_/X _79302_/Y sky130_fd_sc_hd__xnor2_4
Xclkbuf_10_682_0_CLK clkbuf_9_341_0_CLK/X _87720_/CLK sky130_fd_sc_hd__clkbuf_1
X_76514_ _76514_/A _76514_/Y sky130_fd_sc_hd__inv_2
X_42906_ _42895_/X _42896_/X _41676_/X _87659_/Q _42905_/X _42907_/A
+ sky130_fd_sc_hd__o32ai_4
X_49462_ _49467_/A _49456_/B _49447_/C _46791_/X _49462_/X sky130_fd_sc_hd__and4_4
X_61740_ _59664_/C _61777_/A sky130_fd_sc_hd__buf_2
X_73726_ _43043_/Y _73627_/X _73652_/X _73725_/Y _73726_/X sky130_fd_sc_hd__a211o_4
X_46674_ _46720_/A _46712_/A sky130_fd_sc_hd__buf_2
X_70938_ _70935_/A _70939_/A sky130_fd_sc_hd__buf_2
X_77494_ _77495_/A _77491_/Y _77493_/Y _77496_/A sky130_fd_sc_hd__a21o_4
X_43886_ _43842_/A _43886_/X sky130_fd_sc_hd__buf_2
X_48413_ _86524_/Q _48333_/X _48412_/Y _48413_/Y sky130_fd_sc_hd__o21ai_4
X_79233_ _79233_/A _79248_/C sky130_fd_sc_hd__buf_2
X_45625_ _45619_/X _45622_/X _45624_/Y _86865_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_173_0_CLK clkbuf_8_86_0_CLK/X clkbuf_9_173_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_76445_ _76425_/X _76444_/Y _76417_/Y _76445_/Y sky130_fd_sc_hd__o21ai_4
X_42837_ _42816_/X _42817_/X _41493_/X _66710_/B _42836_/X _42837_/Y
+ sky130_fd_sc_hd__o32ai_4
X_61671_ _61690_/A _61690_/B _79129_/B _61671_/Y sky130_fd_sc_hd__nor3_4
X_49393_ _49391_/Y _49378_/X _49392_/X _86396_/D sky130_fd_sc_hd__a21oi_4
X_73657_ _88367_/Q _73279_/X _73656_/X _73657_/X sky130_fd_sc_hd__o21a_4
X_70869_ _70869_/A _70869_/B _70869_/C _70869_/D _70869_/Y sky130_fd_sc_hd__nand4_4
X_63410_ _63410_/A _63410_/B _63410_/C _63410_/D _63410_/X sky130_fd_sc_hd__and4_4
X_48344_ _48341_/Y _48322_/X _48343_/Y _86532_/D sky130_fd_sc_hd__a21boi_4
X_60622_ _60622_/A _60616_/Y _60622_/C _60622_/D _60655_/A sky130_fd_sc_hd__and4_4
X_72608_ _72607_/Y _72572_/A _72572_/B _72608_/Y sky130_fd_sc_hd__nand3_4
X_79164_ _79161_/Y _79524_/A _79163_/Y _79164_/Y sky130_fd_sc_hd__a21boi_4
X_45556_ _45709_/A _45556_/X sky130_fd_sc_hd__buf_2
X_64390_ _64363_/A _64363_/B _84954_/Q _61145_/X _64390_/X sky130_fd_sc_hd__and4_4
X_76376_ _76369_/A _76369_/B _76368_/A _76376_/X sky130_fd_sc_hd__o21a_4
X_42768_ _42822_/A _42768_/X sky130_fd_sc_hd__buf_2
X_73588_ _73588_/A _73588_/B _73588_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_697_0_CLK clkbuf_9_348_0_CLK/X _87382_/CLK sky130_fd_sc_hd__clkbuf_1
X_78115_ _82567_/Q _78108_/B _78115_/Y sky130_fd_sc_hd__nor2_4
X_44507_ _41271_/Y _44502_/X _87074_/Q _44503_/X _87074_/D sky130_fd_sc_hd__a2bb2o_4
X_63341_ _63289_/X _64546_/C _63341_/C _60383_/A _63341_/X sky130_fd_sc_hd__and4_4
X_75327_ _75308_/Y _75309_/A _75326_/X _75328_/B sky130_fd_sc_hd__a21boi_4
X_41719_ _41719_/A _41718_/X _41719_/X sky130_fd_sc_hd__or2_4
X_48275_ _49215_/A _48275_/X sky130_fd_sc_hd__buf_2
X_60553_ _60459_/B _60607_/A sky130_fd_sc_hd__buf_2
X_72539_ _72535_/Y _72539_/B _72539_/Y sky130_fd_sc_hd__nand2_4
X_79095_ _79095_/A _79095_/B _79095_/X sky130_fd_sc_hd__or2_4
X_45487_ _45485_/Y _45439_/X _45471_/X _45486_/Y _45487_/X sky130_fd_sc_hd__a211o_4
X_42699_ _42579_/A _42700_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_188_0_CLK clkbuf_8_94_0_CLK/X clkbuf_9_188_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_47226_ _47226_/A _47227_/A sky130_fd_sc_hd__inv_2
X_66060_ _66040_/X _84983_/Q _66027_/X _66059_/X _66061_/B sky130_fd_sc_hd__a211o_4
X_78046_ _82260_/Q _81972_/Q _78046_/Y sky130_fd_sc_hd__xnor2_4
X_44438_ _41601_/X _44431_/X _87108_/Q _44432_/X _87108_/D sky130_fd_sc_hd__a2bb2o_4
X_63272_ _63272_/A _61611_/A _60488_/C _63272_/Y sky130_fd_sc_hd__nand3_4
X_75258_ _75254_/Y _75258_/B _75258_/C _75258_/X sky130_fd_sc_hd__or3_4
X_60484_ _60484_/A _63280_/C sky130_fd_sc_hd__buf_2
X_65011_ _65009_/X _86162_/Q _64902_/X _65010_/X _65011_/X sky130_fd_sc_hd__a211o_4
X_62223_ _62236_/A _62631_/B sky130_fd_sc_hd__buf_2
X_74209_ _88343_/Q _72769_/B _73007_/A _74209_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_10_620_0_CLK clkbuf_9_310_0_CLK/X _81195_/CLK sky130_fd_sc_hd__clkbuf_1
X_47157_ _47157_/A _54578_/B sky130_fd_sc_hd__inv_2
X_44369_ _44350_/X _44351_/X _41757_/X _87143_/Q _44353_/X _44370_/A
+ sky130_fd_sc_hd__o32ai_4
X_75189_ _75190_/A _75190_/C _75190_/B _75189_/X sky130_fd_sc_hd__a21o_4
X_46108_ _46214_/D _72484_/A _46214_/C _46108_/D _46108_/X sky130_fd_sc_hd__and4_4
X_62154_ _62146_/X _62148_/X _62153_/Y _84869_/Q _62117_/X _62154_/Y
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_9_111_0_CLK clkbuf_8_55_0_CLK/X clkbuf_9_111_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_47088_ _53364_/B _52850_/B sky130_fd_sc_hd__buf_2
X_79997_ _84929_/Q _84177_/Q _79997_/X sky130_fd_sc_hd__xor2_4
X_61105_ _61172_/A _61082_/X _61096_/X _61153_/A _61105_/X sky130_fd_sc_hd__a211o_4
X_46039_ _46013_/X _46032_/X _41497_/X _86799_/Q _46014_/X _46039_/Y
+ sky130_fd_sc_hd__o32ai_4
X_69750_ _73124_/A _69747_/X _68691_/X _69749_/Y _69750_/X sky130_fd_sc_hd__a211o_4
X_66962_ _66961_/X _66962_/B _66962_/X sky130_fd_sc_hd__and2_4
X_62085_ _61708_/X _62128_/C sky130_fd_sc_hd__buf_2
X_78948_ _78948_/A _78948_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_635_0_CLK clkbuf_9_317_0_CLK/X _82284_/CLK sky130_fd_sc_hd__clkbuf_1
X_68701_ _68698_/X _68700_/X _68701_/Y sky130_fd_sc_hd__nand2_4
X_65913_ _65910_/X _65868_/B _65912_/X _65913_/Y sky130_fd_sc_hd__nand3_4
X_61036_ _61028_/X _61018_/Y _61036_/C _61037_/A sky130_fd_sc_hd__nor3_4
X_69681_ _72973_/A _69485_/X _69611_/X _69680_/X _69681_/X sky130_fd_sc_hd__a211o_4
X_66893_ _88390_/Q _66868_/X _66801_/X _66892_/X _66893_/X sky130_fd_sc_hd__a211o_4
X_78879_ _78859_/Y _78873_/Y _78878_/X _78879_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_126_0_CLK clkbuf_8_63_0_CLK/X clkbuf_9_126_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_80910_ _83918_/CLK _80910_/D _80910_/Q sky130_fd_sc_hd__dfxtp_4
X_68632_ _87093_/Q _68580_/X _68630_/X _68631_/X _68632_/X sky130_fd_sc_hd__a211o_4
X_65844_ _84174_/Q _65296_/X _65843_/Y _84174_/D sky130_fd_sc_hd__a21o_4
Xclkbuf_9_53_0_CLK clkbuf_9_53_0_CLK/A clkbuf_9_53_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_81890_ _82015_/CLK _77235_/X _77170_/B sky130_fd_sc_hd__dfxtp_4
X_49729_ _49727_/Y _49706_/X _49728_/X _86334_/D sky130_fd_sc_hd__a21oi_4
X_80841_ _80746_/CLK _80873_/Q _74891_/B sky130_fd_sc_hd__dfxtp_4
X_68563_ _68551_/Y _68358_/X _68447_/X _68562_/Y _68563_/X sky130_fd_sc_hd__a211o_4
X_65775_ _65855_/A _65775_/B _84179_/Q _65775_/X sky130_fd_sc_hd__and3_4
X_62987_ _63516_/A _62987_/X sky130_fd_sc_hd__buf_2
X_67514_ _87468_/Q _67512_/X _67462_/X _67513_/X _67514_/X sky130_fd_sc_hd__a211o_4
X_52740_ _85763_/Q _52737_/X _52739_/Y _52740_/Y sky130_fd_sc_hd__o21ai_4
X_64726_ _64883_/A _86269_/Q _64726_/X sky130_fd_sc_hd__and2_4
X_83560_ _86592_/CLK _71247_/Y _47842_/A sky130_fd_sc_hd__dfxtp_4
X_61938_ _61489_/B _61953_/B _61953_/C _61937_/X _61938_/Y sky130_fd_sc_hd__nand4_4
X_80772_ _83967_/CLK _75890_/Y _75108_/A sky130_fd_sc_hd__dfxtp_4
X_68494_ _68385_/A _68494_/X sky130_fd_sc_hd__buf_2
X_82511_ _82711_/CLK _82511_/D _82511_/Q sky130_fd_sc_hd__dfxtp_4
X_67445_ _86971_/Q _67348_/X _67398_/X _67444_/X _67445_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_9_68_0_CLK clkbuf_9_69_0_CLK/A clkbuf_9_68_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_52671_ _52657_/X _54364_/B _52671_/Y sky130_fd_sc_hd__nand2_4
X_64657_ _64809_/A _64657_/X sky130_fd_sc_hd__buf_2
X_83491_ _83491_/CLK _71459_/X _83491_/Q sky130_fd_sc_hd__dfxtp_4
X_61869_ _61823_/A _61915_/B _58506_/A _61915_/D _61869_/X sky130_fd_sc_hd__and4_4
X_54410_ _54425_/A _52718_/B _54410_/Y sky130_fd_sc_hd__nand2_4
X_85230_ _85257_/CLK _85230_/D _56339_/C sky130_fd_sc_hd__dfxtp_4
X_51622_ _51622_/A _51627_/A sky130_fd_sc_hd__buf_2
X_63608_ _58391_/A _63558_/X _61572_/A _63559_/X _63608_/X sky130_fd_sc_hd__a2bb2o_4
X_82442_ _82443_/CLK _79134_/X _82410_/D sky130_fd_sc_hd__dfxtp_4
X_55390_ _56719_/A _56719_/B _55388_/Y _55441_/C sky130_fd_sc_hd__nand3_4
X_67376_ _67305_/X _67367_/Y _67269_/X _67375_/Y _67376_/X sky130_fd_sc_hd__a211o_4
X_64588_ _59345_/X _86177_/Q _64583_/X _64587_/X _64588_/X sky130_fd_sc_hd__a211o_4
X_69115_ _74266_/A _68958_/X _69113_/X _69114_/Y _69115_/X sky130_fd_sc_hd__a211o_4
X_54341_ _54332_/A _52651_/B _54341_/Y sky130_fd_sc_hd__nand2_4
X_66327_ _66117_/X _84964_/Q _66118_/X _66326_/X _66328_/B sky130_fd_sc_hd__a211o_4
X_85161_ _83016_/CLK _85161_/D _85161_/Q sky130_fd_sc_hd__dfxtp_4
X_51553_ _51553_/A _51553_/B _51553_/C _53078_/D _51553_/X sky130_fd_sc_hd__and4_4
X_63539_ _63478_/A _63541_/B sky130_fd_sc_hd__buf_2
X_82373_ _83690_/CLK _82181_/Q _82373_/Q sky130_fd_sc_hd__dfxtp_4
X_84112_ _84161_/CLK _84112_/D _66495_/C sky130_fd_sc_hd__dfxtp_4
X_50504_ _50502_/Y _50474_/X _50503_/Y _86188_/D sky130_fd_sc_hd__a21boi_4
X_81324_ _84049_/CLK _76297_/X _81700_/D sky130_fd_sc_hd__dfxtp_4
X_57060_ _56873_/X _44220_/B _57059_/Y _57060_/X sky130_fd_sc_hd__a21o_4
X_69046_ _87479_/Q _69044_/X _68979_/X _69045_/X _69046_/X sky130_fd_sc_hd__a211o_4
X_54272_ _54288_/A _46624_/Y _54272_/Y sky130_fd_sc_hd__nand2_4
X_66258_ _66254_/X _66257_/X _66258_/Y sky130_fd_sc_hd__nand2_4
X_85092_ _85041_/CLK _85092_/D _85092_/Q sky130_fd_sc_hd__dfxtp_4
X_51484_ _51482_/Y _51477_/X _51483_/X _86002_/D sky130_fd_sc_hd__a21oi_4
X_56011_ _56010_/X _56054_/B sky130_fd_sc_hd__buf_2
X_53223_ _53217_/A _53211_/B _53222_/X _53223_/D _53223_/X sky130_fd_sc_hd__and4_4
X_65209_ _65155_/A _65209_/B _65209_/X sky130_fd_sc_hd__and2_4
X_84043_ _81475_/CLK _68065_/X _81475_/D sky130_fd_sc_hd__dfxtp_4
X_50435_ _48752_/A _50456_/B _50435_/C _50435_/X sky130_fd_sc_hd__and3_4
X_81255_ _81671_/CLK _81255_/D _81255_/Q sky130_fd_sc_hd__dfxtp_4
X_66189_ _66185_/X _66188_/X _66189_/Y sky130_fd_sc_hd__nand2_4
X_80206_ _59992_/C _80206_/B _80207_/B sky130_fd_sc_hd__xor2_4
X_53154_ _85687_/Q _53146_/X _53153_/Y _53154_/Y sky130_fd_sc_hd__o21ai_4
X_50366_ _86215_/Q _50363_/X _50365_/Y _50366_/Y sky130_fd_sc_hd__o21ai_4
X_81186_ _81211_/CLK _81186_/D _81186_/Q sky130_fd_sc_hd__dfxtp_4
X_52105_ _52100_/A _48380_/X _52105_/Y sky130_fd_sc_hd__nand2_4
X_87802_ _88062_/CLK _87802_/D _73394_/A sky130_fd_sc_hd__dfxtp_4
X_80137_ _80109_/X _80112_/Y _80122_/X _80125_/Y _80137_/X sky130_fd_sc_hd__o22a_4
X_53085_ _53081_/Y _53082_/X _53084_/X _85700_/D sky130_fd_sc_hd__a21oi_4
X_57962_ _58679_/A _57962_/X sky130_fd_sc_hd__buf_2
X_69948_ _69945_/X _69947_/X _69624_/X _69948_/X sky130_fd_sc_hd__a21o_4
X_50297_ _50285_/A _47969_/B _50297_/Y sky130_fd_sc_hd__nand2_4
X_85994_ _85704_/CLK _51528_/Y _85994_/Q sky130_fd_sc_hd__dfxtp_4
X_59701_ _66262_/A _59711_/B sky130_fd_sc_hd__buf_2
X_52036_ _52014_/X _52036_/B _52036_/Y sky130_fd_sc_hd__nand2_4
X_56913_ _57272_/D _57319_/D sky130_fd_sc_hd__buf_2
X_87733_ _87487_/CLK _42762_/Y _87733_/Q sky130_fd_sc_hd__dfxtp_4
X_84945_ _84945_/CLK _57856_/Y _84945_/Q sky130_fd_sc_hd__dfxtp_4
X_80068_ _84936_/Q _65698_/C _80068_/X sky130_fd_sc_hd__xor2_4
X_57893_ _58007_/A _57893_/X sky130_fd_sc_hd__buf_2
X_69879_ _69876_/X _69878_/X _69742_/X _69879_/Y sky130_fd_sc_hd__a21oi_4
X_71910_ _74531_/A _70710_/C _71902_/X _71928_/D _71910_/Y sky130_fd_sc_hd__nand4_4
X_59632_ _59512_/X _59689_/A _59631_/Y _59632_/X sky130_fd_sc_hd__o21a_4
X_56844_ _55290_/A _55678_/A _55670_/B _56844_/X sky130_fd_sc_hd__a21bo_4
X_87664_ _87408_/CLK _87664_/D _67415_/B sky130_fd_sc_hd__dfxtp_4
X_84876_ _84823_/CLK _84876_/D _58329_/A sky130_fd_sc_hd__dfxtp_4
X_72890_ _72889_/X _72890_/X sky130_fd_sc_hd__buf_2
X_86615_ _85969_/CLK _47630_/Y _72247_/A sky130_fd_sc_hd__dfxtp_4
X_71841_ _71072_/A _71714_/Y _70790_/A _70721_/A _71841_/X sky130_fd_sc_hd__and4_4
X_83827_ _83188_/CLK _83827_/D _74755_/B sky130_fd_sc_hd__dfxtp_4
X_59563_ _59563_/A _59564_/B sky130_fd_sc_hd__buf_2
X_56775_ _56775_/A _83324_/Q _56768_/Y _56776_/B sky130_fd_sc_hd__nand3_4
X_87595_ _87595_/CLK _43049_/Y _87595_/Q sky130_fd_sc_hd__dfxtp_4
X_53987_ _53978_/A _52468_/B _53987_/Y sky130_fd_sc_hd__nand2_4
X_58514_ _84830_/Q _63496_/B sky130_fd_sc_hd__buf_2
X_43740_ _48759_/A _47846_/A sky130_fd_sc_hd__buf_2
X_55726_ _55723_/X _55725_/X _55138_/A _55726_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_9_0_CLK clkbuf_8_4_0_CLK/X clkbuf_9_9_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_74560_ _74559_/X _74553_/X _56035_/A _74554_/X _74560_/X sky130_fd_sc_hd__a211o_4
X_86546_ _86554_/CLK _86546_/D _86546_/Q sky130_fd_sc_hd__dfxtp_4
X_40952_ _40952_/A _88305_/D sky130_fd_sc_hd__inv_2
X_52938_ _52922_/A _52954_/B _52926_/X _52938_/D _52938_/X sky130_fd_sc_hd__and4_4
X_71772_ _71763_/X _71815_/B _70986_/A _71772_/X sky130_fd_sc_hd__and3_4
X_59494_ _58230_/A _59493_/Y _59494_/Y sky130_fd_sc_hd__nand2_4
X_83758_ _83761_/CLK _83758_/D _83758_/Q sky130_fd_sc_hd__dfxtp_4
X_73511_ _73508_/X _73510_/X _73347_/X _73524_/B sky130_fd_sc_hd__a21o_4
X_70723_ _52777_/B _70699_/A _70722_/Y _70723_/Y sky130_fd_sc_hd__o21ai_4
X_58445_ _63230_/A _58446_/A sky130_fd_sc_hd__buf_2
X_82709_ _82665_/CLK _82709_/D _82709_/Q sky130_fd_sc_hd__dfxtp_4
X_43671_ _43685_/A _43671_/X sky130_fd_sc_hd__buf_2
X_55657_ _55241_/B _55228_/Y _55657_/Y sky130_fd_sc_hd__xnor2_4
X_86477_ _86499_/CLK _86477_/D _86477_/Q sky130_fd_sc_hd__dfxtp_4
X_74491_ _83055_/Q _74474_/X _74490_/Y _74491_/Y sky130_fd_sc_hd__o21ai_4
X_40883_ _40883_/A _40883_/B _40883_/X sky130_fd_sc_hd__or2_4
X_52869_ _52850_/A _52869_/B _52869_/Y sky130_fd_sc_hd__nand2_4
X_83689_ _83685_/CLK _83689_/D _83689_/Q sky130_fd_sc_hd__dfxtp_4
X_45410_ _55625_/B _45388_/X _45390_/X _45409_/Y _45410_/X sky130_fd_sc_hd__a211o_4
X_88216_ _88215_/CLK _41434_/X _88216_/Q sky130_fd_sc_hd__dfxtp_4
X_76230_ _81640_/Q _76230_/Y sky130_fd_sc_hd__inv_2
X_42622_ _73507_/A _69958_/B sky130_fd_sc_hd__inv_2
X_54608_ _54606_/Y _54584_/X _54607_/X _54608_/Y sky130_fd_sc_hd__a21oi_4
X_73442_ _73439_/X _73441_/X _72862_/X _73442_/X sky130_fd_sc_hd__a21o_4
X_85428_ _85428_/CLK _54517_/Y _85428_/Q sky130_fd_sc_hd__dfxtp_4
X_46390_ _46348_/X _49009_/A _46389_/X _46391_/A sky130_fd_sc_hd__o21ai_4
X_70654_ _53041_/B _70631_/X _70653_/Y _83732_/D sky130_fd_sc_hd__o21ai_4
X_58376_ _84865_/Q _58377_/A sky130_fd_sc_hd__inv_2
X_55588_ _55527_/X _55617_/A sky130_fd_sc_hd__buf_2
XPHY_50 sky130_fd_sc_hd__decap_3
X_45341_ _56452_/C _45326_/X _45340_/X _45341_/Y sky130_fd_sc_hd__o21ai_4
X_57327_ _57188_/A _57327_/B _56818_/X _57328_/A sky130_fd_sc_hd__nand3_4
XPHY_61 sky130_fd_sc_hd__decap_3
X_76161_ _76158_/X _81635_/Q _76159_/Y _76161_/Y sky130_fd_sc_hd__nand3_4
X_88147_ _87436_/CLK _88147_/D _66583_/B sky130_fd_sc_hd__dfxtp_4
X_54539_ _54534_/Y _54530_/X _54538_/X _85424_/D sky130_fd_sc_hd__a21oi_4
X_42553_ _42553_/A _42553_/Y sky130_fd_sc_hd__inv_2
X_73373_ _69883_/B _44235_/X _73031_/X _73372_/Y _73373_/X sky130_fd_sc_hd__a211o_4
X_85359_ _86289_/CLK _54891_/Y _85359_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_72 sky130_fd_sc_hd__decap_3
X_70585_ _70984_/A _70585_/X sky130_fd_sc_hd__buf_2
XPHY_83 sky130_fd_sc_hd__decap_3
XPHY_94 sky130_fd_sc_hd__decap_3
X_75112_ _75113_/A _75113_/C _81061_/Q _75117_/B sky130_fd_sc_hd__a21o_4
X_41504_ _41503_/X _41486_/X _88203_/Q _41487_/X _88203_/D sky130_fd_sc_hd__a2bb2o_4
X_72324_ _59081_/A _72324_/X sky130_fd_sc_hd__buf_2
X_48060_ _48060_/A _53567_/B sky130_fd_sc_hd__inv_2
X_45272_ _45272_/A _45272_/X sky130_fd_sc_hd__buf_2
X_57258_ _56626_/X _57247_/Y _57257_/Y _57258_/Y sky130_fd_sc_hd__a21oi_4
X_76092_ _81722_/D _76092_/B _76093_/A sky130_fd_sc_hd__nand2_4
X_42484_ _42460_/X _42472_/X _40646_/X _68618_/B _42463_/X _87849_/D
+ sky130_fd_sc_hd__o32ai_4
X_88078_ _88081_/CLK _88078_/D _88078_/Q sky130_fd_sc_hd__dfxtp_4
X_47011_ _82392_/Q _54494_/D sky130_fd_sc_hd__inv_2
X_44223_ _69751_/A _66608_/A sky130_fd_sc_hd__buf_2
X_56209_ _56035_/X _56195_/X _56208_/Y _85275_/D sky130_fd_sc_hd__o21ai_4
X_75043_ _75035_/Y _75047_/A _75042_/Y _75043_/Y sky130_fd_sc_hd__a21boi_4
X_79920_ _79918_/Y _79919_/Y _79920_/Y sky130_fd_sc_hd__nand2_4
X_41435_ _41435_/A _41435_/B _41435_/X sky130_fd_sc_hd__or2_4
X_87029_ _88301_/CLK _87029_/D _87029_/Q sky130_fd_sc_hd__dfxtp_4
X_72255_ _72255_/A _72255_/X sky130_fd_sc_hd__buf_2
X_57189_ _57087_/X _57185_/Y _57188_/Y _57189_/Y sky130_fd_sc_hd__o21ai_4
X_71206_ _48816_/B _71190_/X _71205_/Y _83573_/D sky130_fd_sc_hd__o21ai_4
X_44154_ _45920_/A _66563_/A sky130_fd_sc_hd__buf_2
X_79851_ _79828_/Y _79850_/Y _79851_/Y sky130_fd_sc_hd__nor2_4
X_41366_ _41261_/X _81746_/Q _41365_/X _41366_/Y sky130_fd_sc_hd__o21ai_4
X_72186_ _72182_/Y _72184_/Y _72185_/X _72186_/X sky130_fd_sc_hd__a21o_4
X_43105_ _43129_/A _43105_/X sky130_fd_sc_hd__buf_2
X_78802_ _82626_/Q _78802_/Y sky130_fd_sc_hd__inv_2
X_71137_ _71137_/A _71137_/B _71138_/A sky130_fd_sc_hd__nor2_4
X_48962_ _48962_/A _71996_/B sky130_fd_sc_hd__inv_2
X_44085_ _44072_/Y _44293_/B _44085_/C _44085_/D _44085_/Y sky130_fd_sc_hd__nor4_4
X_79782_ _64891_/C _72236_/Y _79781_/Y _79782_/X sky130_fd_sc_hd__o21a_4
X_41297_ _41290_/X _82911_/Q _41296_/X _41298_/A sky130_fd_sc_hd__o21ai_4
X_76994_ _84546_/Q _62328_/C _76994_/X sky130_fd_sc_hd__xor2_4
X_47913_ _66008_/B _47897_/X _47912_/Y _47913_/Y sky130_fd_sc_hd__o21ai_4
X_43036_ _42439_/X _43017_/X _40605_/X _73653_/A _43025_/X _43036_/Y
+ sky130_fd_sc_hd__o32ai_4
X_78733_ _78732_/B _78732_/C _78732_/A _78733_/Y sky130_fd_sc_hd__o21ai_4
X_71068_ _70355_/A _71068_/B _71069_/A sky130_fd_sc_hd__and2_4
X_75945_ _81702_/D _75952_/B _75949_/A sky130_fd_sc_hd__xor2_4
X_48893_ _48893_/A _48894_/A sky130_fd_sc_hd__buf_2
X_62910_ _62910_/A _62967_/A sky130_fd_sc_hd__buf_2
X_70019_ _68620_/X _68622_/X _69992_/X _70021_/A sky130_fd_sc_hd__a21o_4
X_47844_ _47855_/A _50224_/B _47844_/Y sky130_fd_sc_hd__nand2_4
X_78664_ _78663_/B _78663_/C _78663_/A _78664_/Y sky130_fd_sc_hd__o21ai_4
X_63890_ _63741_/A _63890_/X sky130_fd_sc_hd__buf_2
X_75876_ _75876_/A _75876_/B _80897_/D sky130_fd_sc_hd__nand2_4
X_77615_ _77614_/B _77614_/C _77614_/A _77619_/C sky130_fd_sc_hd__o21ai_4
X_62841_ _62979_/A _62841_/X sky130_fd_sc_hd__buf_2
X_74827_ _74829_/A _46188_/A _74828_/A sky130_fd_sc_hd__nand2_4
X_47775_ _81223_/Q _47776_/A sky130_fd_sc_hd__inv_2
X_78595_ _78584_/Y _78585_/Y _78586_/Y _78623_/B sky130_fd_sc_hd__o21a_4
X_44987_ _44981_/Y _44984_/Y _44986_/X _44987_/X sky130_fd_sc_hd__a21o_4
X_49514_ _49434_/A _49514_/X sky130_fd_sc_hd__buf_2
X_46726_ _46915_/A _46737_/A sky130_fd_sc_hd__buf_2
X_65560_ _65557_/Y _65529_/X _65559_/X _84193_/D sky130_fd_sc_hd__a21o_4
X_77546_ _77526_/Y _77561_/B _77561_/A _77547_/B sky130_fd_sc_hd__a21boi_4
X_43938_ _41447_/X _43928_/X _68044_/B _43929_/X _43938_/X sky130_fd_sc_hd__a2bb2o_4
X_62772_ _62949_/B _62772_/X sky130_fd_sc_hd__buf_2
X_74758_ _74741_/X _74758_/B _74758_/C _80644_/A sky130_fd_sc_hd__nand3_4
X_64511_ _61656_/A _64511_/B _64511_/Y sky130_fd_sc_hd__nor2_4
X_49445_ _49454_/A _46758_/X _49445_/Y sky130_fd_sc_hd__nand2_4
X_73709_ _44124_/A _73709_/X sky130_fd_sc_hd__buf_2
X_61723_ _61476_/A _61723_/X sky130_fd_sc_hd__buf_2
X_46657_ _82973_/Q _46658_/A sky130_fd_sc_hd__inv_2
X_65491_ _65488_/X _65490_/X _65457_/X _65491_/X sky130_fd_sc_hd__a21o_4
X_77477_ _77476_/Y _77477_/Y sky130_fd_sc_hd__inv_2
X_43869_ _43605_/A _43869_/X sky130_fd_sc_hd__buf_2
X_74689_ _57050_/A _74656_/X _74688_/Y _74689_/X sky130_fd_sc_hd__a21bo_4
X_67230_ _66868_/A _67230_/X sky130_fd_sc_hd__buf_2
X_79216_ _84790_/Q _84110_/Q _79236_/A sky130_fd_sc_hd__nand2_4
X_45608_ _45452_/A _45608_/X sky130_fd_sc_hd__buf_2
X_64442_ _64386_/A _64442_/X sky130_fd_sc_hd__buf_2
X_76428_ _81269_/Q _81525_/D _76429_/A sky130_fd_sc_hd__nand2_4
X_49376_ _49382_/A _51765_/B _49376_/Y sky130_fd_sc_hd__nand2_4
X_61654_ _61340_/A _61654_/X sky130_fd_sc_hd__buf_2
X_46588_ _86723_/Q _46543_/X _46587_/Y _46588_/Y sky130_fd_sc_hd__o21ai_4
X_48327_ _48319_/A _50370_/B _48327_/Y sky130_fd_sc_hd__nand2_4
X_60605_ _79128_/A _60577_/X _60491_/X _60572_/B _84588_/D sky130_fd_sc_hd__a2bb2oi_4
X_67161_ _67087_/A _67161_/B _67161_/X sky130_fd_sc_hd__and2_4
X_79147_ _79147_/A _84479_/Q _79147_/X sky130_fd_sc_hd__xor2_4
X_45539_ _55539_/B _45489_/X _45520_/X _45538_/Y _45539_/X sky130_fd_sc_hd__a211o_4
X_64373_ _64314_/A _64373_/X sky130_fd_sc_hd__buf_2
X_76359_ _76336_/A _76336_/B _76338_/A _76359_/Y sky130_fd_sc_hd__a21boi_4
X_61585_ _61584_/X _61585_/Y sky130_fd_sc_hd__inv_2
X_66112_ _57694_/X _73901_/B _66112_/X sky130_fd_sc_hd__and2_4
X_63324_ _60433_/A _63324_/B _63333_/C _63240_/X _63324_/X sky130_fd_sc_hd__and4_4
X_48258_ _48255_/Y _48226_/X _48257_/Y _48258_/Y sky130_fd_sc_hd__a21boi_4
X_60536_ _60481_/A _60532_/Y _60586_/A _60534_/Y _60535_/Y _60536_/X
+ sky130_fd_sc_hd__a41o_4
X_67092_ _66971_/A _67092_/X sky130_fd_sc_hd__buf_2
X_79078_ _79065_/Y _79070_/B _79077_/Y _79078_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_6_50_0_CLK clkbuf_6_51_0_CLK/A clkbuf_6_50_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_47209_ _47208_/Y _51225_/D sky130_fd_sc_hd__buf_2
X_66043_ _66043_/A _66042_/X _66043_/Y sky130_fd_sc_hd__nand2_4
X_78029_ _82081_/Q _78028_/X _78030_/A sky130_fd_sc_hd__xor2_4
X_63255_ _63248_/X _63249_/Y _63251_/X _63252_/Y _63254_/Y _63255_/X
+ sky130_fd_sc_hd__a41o_4
X_60467_ _60466_/X _63347_/C sky130_fd_sc_hd__buf_2
X_48189_ _48163_/X _48190_/A sky130_fd_sc_hd__buf_2
X_50220_ _50219_/X _50220_/X sky130_fd_sc_hd__buf_2
X_62206_ _62249_/A _59477_/A _59987_/X _62206_/Y sky130_fd_sc_hd__nand3_4
X_81040_ _81040_/CLK _75284_/X _81040_/Q sky130_fd_sc_hd__dfxtp_4
X_63186_ _63184_/Y _63185_/X _63172_/X _63186_/Y sky130_fd_sc_hd__a21oi_4
X_60398_ _60473_/B _60570_/A sky130_fd_sc_hd__buf_2
X_69802_ _69746_/X _69800_/Y _69733_/X _69801_/Y _69802_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_574_0_CLK clkbuf_9_287_0_CLK/X _87675_/CLK sky130_fd_sc_hd__clkbuf_1
X_50151_ _50131_/A _53879_/B _50151_/X sky130_fd_sc_hd__and2_4
X_62137_ _58198_/A _62105_/X _62065_/D _61948_/X _62136_/X _62137_/X
+ sky130_fd_sc_hd__a41o_4
X_67994_ _67990_/X _67993_/X _67875_/X _67994_/Y sky130_fd_sc_hd__a21oi_4
X_69733_ _69733_/A _69733_/X sky130_fd_sc_hd__buf_2
X_50082_ _52291_/A _50082_/B _50059_/C _50082_/X sky130_fd_sc_hd__and3_4
X_66945_ _66899_/X _66934_/Y _66910_/X _66944_/Y _66945_/X sky130_fd_sc_hd__a211o_4
X_62068_ _62050_/X _62090_/B _78059_/B _62068_/Y sky130_fd_sc_hd__nor3_4
X_82991_ _85134_/CLK _82991_/D _45681_/A sky130_fd_sc_hd__dfxtp_4
X_53910_ _53910_/A _53821_/B _53910_/Y sky130_fd_sc_hd__nand2_4
X_61019_ _60954_/X _60994_/B _60996_/Y _61019_/X sky130_fd_sc_hd__a21o_4
X_84730_ _83464_/CLK _59449_/X _84730_/Q sky130_fd_sc_hd__dfxtp_4
X_81942_ _82005_/CLK _81942_/D _77528_/A sky130_fd_sc_hd__dfxtp_4
X_69664_ _69796_/A _69664_/X sky130_fd_sc_hd__buf_2
X_54890_ _54910_/A _54883_/B _54910_/C _53196_/D _54890_/X sky130_fd_sc_hd__and4_4
X_66876_ _66851_/X _66876_/B _66876_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_589_0_CLK clkbuf_9_294_0_CLK/X _80776_/CLK sky130_fd_sc_hd__clkbuf_1
X_68615_ _69685_/A _73797_/A _68615_/X sky130_fd_sc_hd__and2_4
X_53841_ _53819_/A _53841_/B _53841_/Y sky130_fd_sc_hd__nand2_4
X_65827_ _65827_/A _65827_/B _65827_/Y sky130_fd_sc_hd__nand2_4
X_84661_ _84660_/CLK _84661_/D _60103_/C sky130_fd_sc_hd__dfxtp_4
X_81873_ _82436_/CLK _78064_/X _81841_/D sky130_fd_sc_hd__dfxtp_4
X_69595_ _88081_/Q _69582_/X _69567_/X _69594_/Y _69595_/X sky130_fd_sc_hd__a211o_4
X_86400_ _86400_/CLK _86400_/D _58576_/B sky130_fd_sc_hd__dfxtp_4
X_83612_ _85555_/CLK _71087_/Y _83612_/Q sky130_fd_sc_hd__dfxtp_4
X_56560_ _56558_/X _72641_/C _56564_/B _56564_/C _56564_/D _56560_/X
+ sky130_fd_sc_hd__a41o_4
X_68546_ _69906_/A _68546_/B _68546_/X sky130_fd_sc_hd__and2_4
X_80824_ _80931_/CLK _83968_/Q _80824_/Q sky130_fd_sc_hd__dfxtp_4
X_87380_ _86914_/CLK _43520_/Y _87380_/Q sky130_fd_sc_hd__dfxtp_4
X_53772_ _53798_/A _53773_/A sky130_fd_sc_hd__buf_2
X_65758_ _65621_/A _65775_/B _84180_/Q _65758_/X sky130_fd_sc_hd__and3_4
X_84592_ _84333_/CLK _84592_/D _79132_/A sky130_fd_sc_hd__dfxtp_4
X_50984_ _50929_/A _50985_/B sky130_fd_sc_hd__buf_2
X_55511_ _55510_/X _55511_/X sky130_fd_sc_hd__buf_2
X_86331_ _86651_/CLK _86331_/D _57820_/B sky130_fd_sc_hd__dfxtp_4
X_52723_ _85766_/Q _52711_/X _52722_/Y _52723_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_512_0_CLK clkbuf_9_256_0_CLK/X _81492_/CLK sky130_fd_sc_hd__clkbuf_1
X_64709_ _64898_/A _64710_/A sky130_fd_sc_hd__buf_2
X_83543_ _83544_/CLK _83543_/D _83543_/Q sky130_fd_sc_hd__dfxtp_4
X_56491_ _56055_/X _56483_/X _56490_/Y _85176_/D sky130_fd_sc_hd__o21ai_4
X_80755_ _80754_/CLK _80755_/D _81131_/D sky130_fd_sc_hd__dfxtp_4
X_68477_ _70001_/A _68477_/X sky130_fd_sc_hd__buf_2
X_65689_ _65704_/A _86480_/Q _65689_/X sky130_fd_sc_hd__and2_4
X_58230_ _58230_/A _58229_/Y _58230_/Y sky130_fd_sc_hd__nand2_4
X_55442_ _55442_/A _55442_/Y sky130_fd_sc_hd__inv_2
X_67428_ _87919_/Q _67355_/X _67405_/X _67427_/X _67428_/X sky130_fd_sc_hd__a211o_4
X_86262_ _85562_/CLK _50111_/Y _86262_/Q sky130_fd_sc_hd__dfxtp_4
X_52654_ _52648_/X _52654_/B _52654_/C _52654_/D _52654_/X sky130_fd_sc_hd__and4_4
X_83474_ _83476_/CLK _71505_/Y _83474_/Q sky130_fd_sc_hd__dfxtp_4
X_80686_ _80719_/CLK _80718_/Q _75239_/A sky130_fd_sc_hd__dfxtp_4
X_88001_ _88001_/CLK _42166_/Y _88001_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_604 sky130_fd_sc_hd__decap_3
X_85213_ _85213_/CLK _56389_/Y _85213_/Q sky130_fd_sc_hd__dfxtp_4
X_51605_ _51617_/A _53131_/B _51605_/Y sky130_fd_sc_hd__nand2_4
X_82425_ _82425_/CLK _82457_/Q _78646_/A sky130_fd_sc_hd__dfxtp_4
X_58161_ _58153_/X _83494_/Q _58160_/Y _58161_/X sky130_fd_sc_hd__o21a_4
XPHY_615 sky130_fd_sc_hd__decap_3
X_55373_ _55288_/Y _55292_/X _55373_/Y sky130_fd_sc_hd__nand2_4
X_67359_ _68347_/A _67359_/X sky130_fd_sc_hd__buf_2
X_86193_ _86193_/CLK _86193_/D _86193_/Q sky130_fd_sc_hd__dfxtp_4
X_52585_ _52583_/Y _52532_/X _52584_/X _85792_/D sky130_fd_sc_hd__a21oi_4
XPHY_626 sky130_fd_sc_hd__decap_3
XPHY_637 sky130_fd_sc_hd__decap_3
XPHY_648 sky130_fd_sc_hd__decap_3
Xclkbuf_10_527_0_CLK clkbuf_9_263_0_CLK/X _81575_/CLK sky130_fd_sc_hd__clkbuf_1
X_57112_ _57086_/X _57112_/X sky130_fd_sc_hd__buf_2
X_54324_ _85463_/Q _54320_/X _54323_/Y _54324_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_6_18_0_CLK clkbuf_5_9_0_CLK/X clkbuf_6_18_0_CLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_659 sky130_fd_sc_hd__decap_3
X_85144_ _85144_/CLK _56620_/X _85144_/Q sky130_fd_sc_hd__dfxtp_4
X_51536_ _85992_/Q _51511_/X _51535_/Y _51536_/Y sky130_fd_sc_hd__o21ai_4
X_70370_ _70370_/A _70375_/C sky130_fd_sc_hd__buf_2
X_58092_ _58087_/Y _58091_/Y _58035_/X _58092_/X sky130_fd_sc_hd__a21o_4
X_82356_ _82349_/CLK _77182_/X _47973_/A sky130_fd_sc_hd__dfxtp_4
X_57043_ _57331_/A _57043_/B _57331_/C _57043_/Y sky130_fd_sc_hd__nand3_4
X_81307_ _81279_/CLK _76995_/X _81275_/D sky130_fd_sc_hd__dfxtp_4
X_69029_ _69026_/X _69029_/B _69029_/Y sky130_fd_sc_hd__nand2_4
X_54255_ _54255_/A _54246_/X _54255_/C _53084_/D _54255_/X sky130_fd_sc_hd__and4_4
X_85075_ _85075_/CLK _85075_/D _45611_/A sky130_fd_sc_hd__dfxtp_4
X_51467_ _51473_/A _51473_/B _51467_/C _52993_/D _51467_/X sky130_fd_sc_hd__and4_4
X_82287_ _82288_/CLK _82287_/D _41034_/A sky130_fd_sc_hd__dfxtp_4
X_41220_ _41219_/X _41220_/X sky130_fd_sc_hd__buf_2
X_72040_ _72040_/A _49055_/A _72040_/Y sky130_fd_sc_hd__nand2_4
X_53206_ _85677_/Q _53198_/X _53205_/Y _53206_/Y sky130_fd_sc_hd__o21ai_4
X_84026_ _86807_/CLK _68151_/X _82066_/D sky130_fd_sc_hd__dfxtp_4
X_50418_ _50415_/Y _50380_/X _50417_/Y _86205_/D sky130_fd_sc_hd__a21boi_4
X_81238_ _85334_/CLK _81046_/Q _81238_/Q sky130_fd_sc_hd__dfxtp_4
X_54186_ _54191_/A _54186_/B _54191_/C _53019_/D _54186_/X sky130_fd_sc_hd__and4_4
X_51398_ _51212_/A _52924_/B _51398_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_2_3_0_CLK clkbuf_2_3_0_CLK/A clkbuf_2_3_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_41151_ _41151_/A _41151_/X sky130_fd_sc_hd__buf_2
X_53137_ _53111_/A _53137_/X sky130_fd_sc_hd__buf_2
X_50349_ _50317_/X _48073_/B _50349_/Y sky130_fd_sc_hd__nand2_4
X_81169_ _81169_/CLK _74956_/B _81169_/Q sky130_fd_sc_hd__dfxtp_4
X_58994_ _58548_/A _83434_/Q _58994_/Y sky130_fd_sc_hd__nor2_4
X_41082_ _41081_/X _41082_/X sky130_fd_sc_hd__buf_2
X_53068_ _85703_/Q _53065_/X _53067_/Y _53068_/Y sky130_fd_sc_hd__o21ai_4
X_57945_ _57884_/X _85489_/Q _57923_/X _57945_/X sky130_fd_sc_hd__o21a_4
X_85977_ _85688_/CLK _85977_/D _85977_/Q sky130_fd_sc_hd__dfxtp_4
X_73991_ _73988_/X _73990_/X _73421_/X _73991_/X sky130_fd_sc_hd__a21o_4
X_44910_ _45612_/A _45824_/B sky130_fd_sc_hd__buf_2
X_52019_ _52027_/A _48016_/B _52019_/Y sky130_fd_sc_hd__nand2_4
X_87716_ _87150_/CLK _87716_/D _67700_/B sky130_fd_sc_hd__dfxtp_4
X_75730_ _75736_/B _75730_/B _75731_/B sky130_fd_sc_hd__xnor2_4
X_72942_ _83171_/Q _72794_/X _72941_/Y _72942_/X sky130_fd_sc_hd__a21o_4
X_84928_ _84926_/CLK _84928_/D _84928_/Q sky130_fd_sc_hd__dfxtp_4
X_45890_ _44120_/Y _45890_/X sky130_fd_sc_hd__buf_2
X_57876_ _57824_/X _85495_/Q _57849_/X _57876_/X sky130_fd_sc_hd__o21a_4
X_59615_ _59615_/A _60403_/C sky130_fd_sc_hd__buf_2
X_44841_ _41720_/Y _44838_/X _86926_/Q _44839_/X _44841_/X sky130_fd_sc_hd__a2bb2o_4
X_56827_ _56820_/Y _56827_/B _56827_/Y sky130_fd_sc_hd__nand2_4
X_75661_ _75650_/Y _75661_/Y sky130_fd_sc_hd__inv_2
X_87647_ _87898_/CLK _87647_/D _87647_/Q sky130_fd_sc_hd__dfxtp_4
X_72873_ _72910_/A _72874_/A sky130_fd_sc_hd__buf_2
X_84859_ _84250_/CLK _58398_/X _84859_/Q sky130_fd_sc_hd__dfxtp_4
X_77400_ _77383_/Y _77382_/X _77386_/A _77400_/Y sky130_fd_sc_hd__a21boi_4
X_74612_ _74549_/Y _74612_/X sky130_fd_sc_hd__buf_2
X_47560_ _47554_/Y _47555_/X _47559_/X _47560_/Y sky130_fd_sc_hd__a21oi_4
X_71824_ _71823_/Y _71824_/Y sky130_fd_sc_hd__inv_2
X_59546_ _59546_/A _59564_/A sky130_fd_sc_hd__buf_2
X_78380_ _78380_/A _78380_/B _78397_/B sky130_fd_sc_hd__nor2_4
X_44772_ _44772_/A _86964_/D sky130_fd_sc_hd__inv_2
X_56758_ _56785_/B _56758_/X sky130_fd_sc_hd__buf_2
X_75592_ _80900_/Q _75594_/B sky130_fd_sc_hd__inv_2
X_87578_ _88060_/CLK _43095_/Y _87578_/Q sky130_fd_sc_hd__dfxtp_4
X_41984_ _42000_/A _41984_/X sky130_fd_sc_hd__buf_2
X_46511_ _54054_/B _49320_/B sky130_fd_sc_hd__buf_2
X_77331_ _77327_/Y _77329_/Y _77332_/C _77334_/A sky130_fd_sc_hd__a21oi_4
X_43723_ _43722_/X _43723_/Y sky130_fd_sc_hd__inv_2
X_55709_ _55706_/X _55708_/X _56127_/B sky130_fd_sc_hd__nand2_4
X_74543_ _74541_/A _46215_/B _44917_/A _74543_/Y sky130_fd_sc_hd__nand3_4
X_86529_ _83589_/CLK _86529_/D _86529_/Q sky130_fd_sc_hd__dfxtp_4
X_40935_ _40935_/A _40935_/X sky130_fd_sc_hd__buf_2
X_47491_ _47517_/A _53076_/B _47491_/Y sky130_fd_sc_hd__nand2_4
X_71755_ _71026_/A _71755_/X sky130_fd_sc_hd__buf_2
X_59477_ _59477_/A _59478_/A sky130_fd_sc_hd__inv_2
X_56689_ _56689_/A _56688_/X _56694_/A sky130_fd_sc_hd__nand2_4
X_49230_ _51256_/A _49113_/B _49091_/C _49230_/X sky130_fd_sc_hd__and3_4
X_46442_ _46441_/Y _51320_/B sky130_fd_sc_hd__buf_2
X_70706_ _74515_/C _70721_/A sky130_fd_sc_hd__buf_2
X_58428_ _58423_/X _83363_/Q _58427_/Y _84851_/D sky130_fd_sc_hd__o21a_4
X_77262_ _77262_/A _82180_/D _77262_/X sky130_fd_sc_hd__xor2_4
X_43654_ _40712_/X _43624_/X _87325_/Q _43625_/X _43654_/X sky130_fd_sc_hd__a2bb2o_4
X_74474_ _46279_/A _74474_/X sky130_fd_sc_hd__buf_2
X_40866_ _40866_/A _40866_/X sky130_fd_sc_hd__buf_2
X_71686_ _71488_/X _71685_/X _71313_/X _71686_/Y sky130_fd_sc_hd__nand3_4
X_79001_ _79001_/A _79001_/B _82711_/D sky130_fd_sc_hd__xor2_4
X_76213_ _81350_/Q _76213_/B _76213_/X sky130_fd_sc_hd__xor2_4
X_42605_ _42568_/X _42569_/X _40890_/X _42604_/Y _42571_/X _87804_/D
+ sky130_fd_sc_hd__o32ai_4
X_73425_ _72721_/X _86183_/Q _73351_/X _73424_/X _73425_/X sky130_fd_sc_hd__a211o_4
X_49161_ _49161_/A _49161_/B _49161_/Y sky130_fd_sc_hd__nor2_4
X_46373_ _51290_/B _53993_/B sky130_fd_sc_hd__buf_2
X_70637_ _70637_/A _70638_/A sky130_fd_sc_hd__buf_2
X_58359_ _63326_/A _58360_/A sky130_fd_sc_hd__buf_2
X_77193_ _77193_/A _77202_/B sky130_fd_sc_hd__buf_2
X_43585_ _51337_/A _43585_/X sky130_fd_sc_hd__buf_2
X_40797_ _40773_/X _82299_/Q _40796_/X _40798_/A sky130_fd_sc_hd__o21ai_4
X_48112_ _48138_/A _48112_/B _48112_/X sky130_fd_sc_hd__and2_4
X_45324_ _55730_/B _45281_/X _45311_/X _45324_/X sky130_fd_sc_hd__o21a_4
X_76144_ _81728_/D _76144_/B _76145_/B sky130_fd_sc_hd__nand2_4
X_42536_ _42554_/A _42536_/X sky130_fd_sc_hd__buf_2
X_49092_ _49085_/Y _49086_/X _49091_/X _86445_/D sky130_fd_sc_hd__a21oi_4
X_61370_ _61364_/Y _61366_/Y _61334_/X _61367_/Y _61369_/Y _61370_/X
+ sky130_fd_sc_hd__a41o_4
X_73356_ _73426_/A _86474_/Q _73356_/X sky130_fd_sc_hd__and2_4
X_70568_ _71865_/A _70549_/X _70568_/C _70568_/D _70568_/Y sky130_fd_sc_hd__nor4_4
X_60321_ _60249_/X _60276_/Y _60165_/A _60367_/B _60320_/Y _84634_/D
+ sky130_fd_sc_hd__a41oi_4
X_72307_ _72305_/X _85362_/Q _72306_/X _72307_/Y sky130_fd_sc_hd__o21ai_4
X_48043_ _48606_/A _48043_/X sky130_fd_sc_hd__buf_2
X_45255_ _45251_/Y _45254_/Y _45212_/X _45255_/X sky130_fd_sc_hd__a21o_4
X_76075_ _81720_/D _76075_/B _76082_/A sky130_fd_sc_hd__xor2_4
X_42467_ _42574_/A _42467_/X sky130_fd_sc_hd__buf_2
X_73287_ _73283_/X _73286_/X _73262_/X _73290_/A sky130_fd_sc_hd__a21o_4
X_70499_ _70502_/A _70500_/D sky130_fd_sc_hd__buf_2
X_44206_ _56670_/A _44207_/A sky130_fd_sc_hd__buf_2
X_79903_ _79903_/A _65888_/C _79903_/Y sky130_fd_sc_hd__nand2_4
X_63040_ _60469_/X _63041_/A sky130_fd_sc_hd__buf_2
X_75026_ _75018_/A _75023_/B _75016_/Y _75026_/Y sky130_fd_sc_hd__o21ai_4
X_41418_ _41486_/A _41418_/X sky130_fd_sc_hd__buf_2
X_60252_ _60263_/A _60367_/C _60285_/A _60252_/X sky130_fd_sc_hd__o21a_4
X_72238_ _72180_/X _85335_/Q _72225_/X _72238_/X sky130_fd_sc_hd__o21a_4
X_45186_ _45179_/X _45183_/Y _45185_/Y _45186_/Y sky130_fd_sc_hd__a21oi_4
X_42398_ _41872_/A _42398_/X sky130_fd_sc_hd__buf_2
X_44137_ _44137_/A _44163_/B sky130_fd_sc_hd__buf_2
X_79834_ _79825_/X _79834_/B _79834_/Y sky130_fd_sc_hd__nand2_4
X_41349_ _41349_/A _88232_/D sky130_fd_sc_hd__inv_2
X_60183_ _60183_/A _59551_/A _60184_/A sky130_fd_sc_hd__and2_4
X_72169_ _72155_/X _85693_/Q _72156_/X _72169_/X sky130_fd_sc_hd__o21a_4
X_49994_ _49915_/A _49994_/X sky130_fd_sc_hd__buf_2
X_48945_ _86459_/Q _48896_/X _48944_/Y _48945_/Y sky130_fd_sc_hd__o21ai_4
X_44068_ _44186_/A _44202_/A _44067_/Y _44068_/Y sky130_fd_sc_hd__nor3_4
X_79765_ _79763_/X _79765_/B _79766_/B sky130_fd_sc_hd__xnor2_4
X_64991_ _64991_/A _64991_/X sky130_fd_sc_hd__buf_2
X_76977_ _76977_/A _84401_/Q _76977_/X sky130_fd_sc_hd__xor2_4
X_43019_ _40361_/A _43013_/X _43019_/B1 _43020_/A sky130_fd_sc_hd__a21o_4
X_66730_ _66727_/X _66729_/X _66706_/X _66730_/Y sky130_fd_sc_hd__a21oi_4
X_78716_ _78715_/X _78716_/Y sky130_fd_sc_hd__inv_2
X_63942_ _63942_/A _59407_/A _63958_/C _63942_/X sky130_fd_sc_hd__and3_4
X_75928_ _75928_/A _75927_/X _75929_/B sky130_fd_sc_hd__xnor2_4
X_48876_ _83625_/Q _48876_/Y sky130_fd_sc_hd__inv_2
X_79696_ _79704_/A _79696_/B _79696_/Y sky130_fd_sc_hd__xnor2_4
X_47827_ _48361_/B _47867_/A _47827_/Y sky130_fd_sc_hd__nand2_4
X_66661_ _84102_/Q _66614_/X _66660_/X _84102_/D sky130_fd_sc_hd__a21bo_4
X_78647_ _78646_/A _82681_/D _78648_/A sky130_fd_sc_hd__nand2_4
X_63873_ _57652_/X _63858_/B _63858_/C _63902_/D _63873_/Y sky130_fd_sc_hd__nand4_4
X_75859_ _75854_/Y _75836_/B _75858_/Y _75860_/B sky130_fd_sc_hd__o21ai_4
X_68400_ _70001_/A _68400_/X sky130_fd_sc_hd__buf_2
X_65612_ _65735_/A _65612_/B _65612_/X sky130_fd_sc_hd__and2_4
X_62824_ _62820_/Y _62772_/X _62821_/Y _62822_/Y _62823_/X _62824_/X
+ sky130_fd_sc_hd__a41o_4
X_69380_ _83928_/Q _69367_/X _69379_/X _69380_/X sky130_fd_sc_hd__a21bo_4
X_47758_ _47758_/A _47777_/B _47777_/C _53230_/D _47758_/X sky130_fd_sc_hd__and4_4
X_66592_ _66589_/X _66591_/X _66547_/X _66597_/A sky130_fd_sc_hd__a21o_4
X_78578_ _78525_/A _78528_/A _78536_/X _78578_/X sky130_fd_sc_hd__a21o_4
X_68331_ _68208_/X _68331_/X sky130_fd_sc_hd__buf_2
X_46709_ _46703_/Y _46704_/X _46708_/X _46709_/Y sky130_fd_sc_hd__a21oi_4
X_65543_ _65543_/A _65543_/B _65543_/Y sky130_fd_sc_hd__nand2_4
X_77529_ _77518_/A _82114_/Q _77529_/Y sky130_fd_sc_hd__nor2_4
X_62755_ _62731_/A _63103_/A _62744_/X _62717_/X _62755_/X sky130_fd_sc_hd__and4_4
X_47689_ _72332_/A _47666_/X _47688_/Y _47689_/Y sky130_fd_sc_hd__o21ai_4
X_61706_ _61755_/A _61706_/X sky130_fd_sc_hd__buf_2
X_49428_ _58720_/B _49415_/X _49427_/Y _49428_/Y sky130_fd_sc_hd__o21ai_4
X_80540_ _80538_/X _80540_/B _80541_/B sky130_fd_sc_hd__xnor2_4
X_68262_ _68246_/X _67602_/Y _68247_/X _68261_/Y _68262_/X sky130_fd_sc_hd__a211o_4
X_65474_ _65673_/A _65474_/X sky130_fd_sc_hd__buf_2
X_62686_ _62677_/Y _62660_/X _62678_/Y _62683_/Y _62685_/X _62686_/X
+ sky130_fd_sc_hd__a41o_4
X_67213_ _67259_/A _87608_/Q _67213_/X sky130_fd_sc_hd__and2_4
X_64425_ _58259_/A _64423_/X _64424_/Y _64425_/Y sky130_fd_sc_hd__o21ai_4
X_49359_ _49357_/Y _49316_/X _49358_/X _86402_/D sky130_fd_sc_hd__a21oi_4
X_61637_ _59430_/A _61637_/X sky130_fd_sc_hd__buf_2
X_80471_ _80471_/A _80471_/B _80471_/X sky130_fd_sc_hd__xor2_4
X_68193_ _67205_/X _67207_/X _68169_/X _68193_/Y sky130_fd_sc_hd__a21oi_4
X_82210_ _81834_/CLK _82242_/Q _77234_/A sky130_fd_sc_hd__dfxtp_4
X_67144_ _67144_/A _67241_/A sky130_fd_sc_hd__buf_2
X_52370_ _52370_/A _52310_/B _52369_/X _52370_/X sky130_fd_sc_hd__and3_4
X_64356_ _58326_/A _64308_/X _64355_/Y _64356_/Y sky130_fd_sc_hd__o21ai_4
X_83190_ _83191_/CLK _72684_/X _83190_/Q sky130_fd_sc_hd__dfxtp_4
X_61568_ _61558_/A _61568_/B _61538_/C _61568_/Y sky130_fd_sc_hd__nand3_4
X_51321_ _65051_/B _51309_/X _51320_/Y _51321_/Y sky130_fd_sc_hd__o21ai_4
X_63307_ _63305_/X _63392_/B _79231_/A _63307_/Y sky130_fd_sc_hd__nor3_4
X_82141_ _82047_/CLK _77984_/Y _77444_/B sky130_fd_sc_hd__dfxtp_4
X_60519_ _60526_/A _60519_/B _79147_/A _60519_/Y sky130_fd_sc_hd__nor3_4
X_67075_ _66717_/A _67075_/X sky130_fd_sc_hd__buf_2
X_64287_ _64287_/A _84851_/Q _64287_/C _64287_/Y sky130_fd_sc_hd__nand3_4
X_61499_ _61499_/A _61499_/B _61459_/X _61499_/Y sky130_fd_sc_hd__nand3_4
X_54040_ _54038_/Y _54015_/X _54039_/X _54040_/Y sky130_fd_sc_hd__a21oi_4
X_66026_ _66023_/X _66025_/X _65880_/X _66030_/A sky130_fd_sc_hd__a21o_4
X_51252_ _51250_/Y _51237_/X _51251_/X _51252_/Y sky130_fd_sc_hd__a21oi_4
X_63238_ _63288_/A _63238_/B _63312_/C _63237_/X _63238_/X sky130_fd_sc_hd__and4_4
X_82072_ _81154_/CLK _82072_/D _82072_/Q sky130_fd_sc_hd__dfxtp_4
X_50203_ _50187_/X _50716_/B _50203_/Y sky130_fd_sc_hd__nand2_4
X_81023_ _84175_/CLK _64663_/C _81023_/Q sky130_fd_sc_hd__dfxtp_4
X_85900_ _86570_/CLK _85900_/D _66209_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_8_1_CLK clkbuf_4_8_1_CLK/A clkbuf_4_8_1_CLK/X sky130_fd_sc_hd__clkbuf_1
X_51183_ _51128_/A _51183_/X sky130_fd_sc_hd__buf_2
X_63169_ _63164_/Y _63166_/X _63167_/X _63168_/X _63125_/X _63169_/Y
+ sky130_fd_sc_hd__o41ai_4
X_86880_ _84418_/CLK _45385_/Y _62629_/A sky130_fd_sc_hd__dfxtp_4
X_50134_ _65037_/B _50113_/X _50133_/Y _50134_/Y sky130_fd_sc_hd__o21ai_4
X_85831_ _86154_/CLK _52396_/Y _65282_/B sky130_fd_sc_hd__dfxtp_4
X_55991_ _55688_/X _55987_/X _55990_/Y _55991_/Y sky130_fd_sc_hd__o21ai_4
X_67977_ _68442_/A _67977_/X sky130_fd_sc_hd__buf_2
X_57730_ _84952_/Q _57691_/X _57723_/X _57729_/X _84952_/D sky130_fd_sc_hd__a2bb2oi_4
X_69716_ _69293_/Y _69644_/X _69672_/X _69715_/Y _69716_/X sky130_fd_sc_hd__a211o_4
X_50065_ _50084_/A _48901_/B _50065_/Y sky130_fd_sc_hd__nand2_4
X_54942_ _54955_/A _54942_/B _46617_/A _53249_/D _54942_/X sky130_fd_sc_hd__and4_4
X_66928_ _87940_/Q _66875_/X _66926_/X _66927_/X _66928_/X sky130_fd_sc_hd__a211o_4
X_85762_ _85764_/CLK _52747_/Y _85762_/Q sky130_fd_sc_hd__dfxtp_4
X_82974_ _82975_/CLK _82782_/Q _82974_/Q sky130_fd_sc_hd__dfxtp_4
X_87501_ _87766_/CLK _43282_/X _87501_/Q sky130_fd_sc_hd__dfxtp_4
X_84713_ _84713_/CLK _59652_/X _80625_/A sky130_fd_sc_hd__dfxtp_4
X_57661_ _57660_/X _57657_/B _57661_/Y sky130_fd_sc_hd__nor2_4
X_69647_ _87565_/Q _69645_/X _68552_/X _69646_/X _69647_/X sky130_fd_sc_hd__a211o_4
X_81925_ _82116_/CLK _78048_/Y _77277_/A sky130_fd_sc_hd__dfxtp_4
X_54873_ _54900_/A _54883_/B sky130_fd_sc_hd__buf_2
X_85693_ _85692_/CLK _53126_/Y _85693_/Q sky130_fd_sc_hd__dfxtp_4
X_66859_ _66859_/A _66858_/X _66859_/Y sky130_fd_sc_hd__nand2_4
X_59400_ _59394_/X _83487_/Q _59399_/Y _59400_/X sky130_fd_sc_hd__o21a_4
X_56612_ _56582_/A _55552_/X _56609_/X _56611_/Y _56613_/A sky130_fd_sc_hd__a211o_4
X_87432_ _87625_/CLK _43416_/Y _87432_/Q sky130_fd_sc_hd__dfxtp_4
X_53824_ _85561_/Q _53816_/X _53823_/Y _53824_/Y sky130_fd_sc_hd__o21ai_4
X_84644_ _84649_/CLK _84644_/D _79826_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_451_0_CLK clkbuf_9_225_0_CLK/X _86301_/CLK sky130_fd_sc_hd__clkbuf_1
X_57592_ _71978_/A _57592_/X sky130_fd_sc_hd__buf_2
X_69578_ _81985_/D _69564_/X _69577_/X _83913_/D sky130_fd_sc_hd__a21bo_4
X_81856_ _82515_/CLK _81888_/Q _77712_/A sky130_fd_sc_hd__dfxtp_4
X_59331_ _57759_/X _59331_/X sky130_fd_sc_hd__buf_2
X_56543_ _56168_/X _56462_/X _56542_/Y _85155_/D sky130_fd_sc_hd__o21ai_4
X_80807_ _83973_/CLK _83951_/Q _80807_/Q sky130_fd_sc_hd__dfxtp_4
X_68529_ _88013_/Q _68527_/X _68501_/X _68528_/X _68529_/X sky130_fd_sc_hd__a211o_4
X_87363_ _86796_/CLK _87363_/D _87363_/Q sky130_fd_sc_hd__dfxtp_4
X_53755_ _53755_/A _53766_/A sky130_fd_sc_hd__buf_2
X_84575_ _84564_/CLK _60753_/Y _84575_/Q sky130_fd_sc_hd__dfxtp_4
X_50967_ _50971_/A _46758_/X _50967_/Y sky130_fd_sc_hd__nand2_4
X_81787_ _80928_/CLK _75925_/X _48426_/A sky130_fd_sc_hd__dfxtp_4
X_86314_ _86312_/CLK _86314_/D _58038_/B sky130_fd_sc_hd__dfxtp_4
X_40720_ _40599_/A _40720_/X sky130_fd_sc_hd__buf_2
X_52706_ _52706_/A _52706_/B _52706_/Y sky130_fd_sc_hd__nand2_4
X_71540_ _71531_/X _83464_/Q _71539_/Y _83464_/D sky130_fd_sc_hd__a21o_4
X_59262_ _59260_/X _85420_/Q _59261_/X _59262_/Y sky130_fd_sc_hd__o21ai_4
X_83526_ _83526_/CLK _71360_/X _83526_/Q sky130_fd_sc_hd__dfxtp_4
X_56474_ _56528_/A _56474_/X sky130_fd_sc_hd__buf_2
X_80738_ _80740_/CLK _75081_/X _81146_/D sky130_fd_sc_hd__dfxtp_4
X_87294_ _87820_/CLK _87294_/D _73299_/A sky130_fd_sc_hd__dfxtp_4
X_53686_ _53684_/Y _53680_/X _53685_/X _85588_/D sky130_fd_sc_hd__a21oi_4
X_50898_ _50908_/A _50045_/X _50897_/X _51761_/D _50898_/X sky130_fd_sc_hd__and4_4
X_58213_ _84906_/Q _63713_/A sky130_fd_sc_hd__inv_2
Xclkbuf_10_466_0_CLK clkbuf_9_233_0_CLK/X _86695_/CLK sky130_fd_sc_hd__clkbuf_1
X_55425_ _55156_/X _55160_/X _57186_/B _55428_/C sky130_fd_sc_hd__a21o_4
X_86245_ _86149_/CLK _50198_/Y _65327_/B sky130_fd_sc_hd__dfxtp_4
X_40651_ _40595_/X _40651_/X sky130_fd_sc_hd__buf_2
XPHY_401 sky130_fd_sc_hd__decap_3
X_52637_ _52637_/A _52637_/B _52637_/Y sky130_fd_sc_hd__nand2_4
X_59193_ _58897_/A _59282_/B sky130_fd_sc_hd__buf_2
X_71471_ _70880_/B _71479_/B _70771_/A _71476_/D _71471_/X sky130_fd_sc_hd__and4_4
X_83457_ _83457_/CLK _83457_/D _83457_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_412 sky130_fd_sc_hd__decap_3
X_80669_ _86841_/CLK _74813_/Y _80669_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_423 sky130_fd_sc_hd__decap_3
X_73210_ _73355_/A _73210_/X sky130_fd_sc_hd__buf_2
XPHY_434 sky130_fd_sc_hd__decap_3
X_58144_ _84922_/Q _58095_/X _58137_/X _58143_/X _84922_/D sky130_fd_sc_hd__a2bb2oi_4
X_70422_ _70421_/Y _70422_/X sky130_fd_sc_hd__buf_2
XPHY_445 sky130_fd_sc_hd__decap_3
X_82408_ _82248_/CLK _82440_/Q _78385_/A sky130_fd_sc_hd__dfxtp_4
X_55356_ _55356_/A _55362_/A _56708_/A sky130_fd_sc_hd__nand2_4
X_43370_ _43178_/X _43396_/A sky130_fd_sc_hd__buf_2
X_74190_ _44738_/Y _73491_/X _74189_/Y _74190_/X sky130_fd_sc_hd__a21o_4
X_86176_ _85566_/CLK _50569_/Y _86176_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_456 sky130_fd_sc_hd__decap_3
X_40582_ _40550_/X _40556_/X _40581_/X _88369_/Q _40568_/X _40583_/A
+ sky130_fd_sc_hd__o32ai_4
X_52568_ _65375_/B _52549_/X _52567_/Y _52568_/Y sky130_fd_sc_hd__o21ai_4
X_83388_ _85404_/CLK _83388_/D _83388_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_467 sky130_fd_sc_hd__decap_3
XPHY_478 sky130_fd_sc_hd__decap_3
X_42321_ _42307_/X _42319_/X _41631_/X _87923_/Q _42320_/X _42321_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54307_ _54312_/A _54325_/B _54312_/C _46688_/Y _54307_/X sky130_fd_sc_hd__and4_4
X_73141_ _48514_/A _73141_/B _73141_/X sky130_fd_sc_hd__xor2_4
XPHY_489 sky130_fd_sc_hd__decap_3
X_85127_ _85128_/CLK _56875_/X _55281_/A sky130_fd_sc_hd__dfxtp_4
X_51519_ _85995_/Q _51511_/X _51518_/Y _51519_/Y sky130_fd_sc_hd__o21ai_4
X_58075_ _58065_/X _85703_/Q _58020_/X _58075_/X sky130_fd_sc_hd__o21a_4
X_70353_ HASH_ADDR[5] _70412_/A sky130_fd_sc_hd__inv_2
X_82339_ _82339_/CLK _77060_/X _48146_/A sky130_fd_sc_hd__dfxtp_4
X_55287_ _55287_/A _55284_/X _55674_/B _55286_/Y _55287_/X sky130_fd_sc_hd__and4_4
X_52499_ _52495_/Y _52496_/X _52498_/X _52499_/Y sky130_fd_sc_hd__a21oi_4
X_45040_ _45720_/A _45040_/X sky130_fd_sc_hd__buf_2
X_57026_ _56551_/X _57026_/X sky130_fd_sc_hd__buf_2
X_42252_ _42204_/X _42252_/X sky130_fd_sc_hd__buf_2
X_54238_ _54235_/Y _54226_/X _54237_/X _54238_/Y sky130_fd_sc_hd__a21oi_4
X_73072_ _73068_/X _73071_/X _73073_/B sky130_fd_sc_hd__nand2_4
X_85058_ _85100_/CLK _85058_/D _55211_/B sky130_fd_sc_hd__dfxtp_4
X_70284_ _70249_/X _70292_/D sky130_fd_sc_hd__buf_2
X_41203_ _41203_/A _41203_/X sky130_fd_sc_hd__buf_2
X_72023_ _83300_/Q _72016_/X _72022_/Y _72023_/Y sky130_fd_sc_hd__o21ai_4
X_76900_ _76901_/A _76893_/Y _76899_/Y _76904_/A sky130_fd_sc_hd__a21o_4
X_84009_ _84074_/CLK _68219_/X _82657_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_510_0_CLK clkbuf_9_510_0_CLK/A clkbuf_9_510_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_42183_ _42137_/A _42183_/X sky130_fd_sc_hd__buf_2
X_54169_ _54184_/A _47352_/A _54169_/Y sky130_fd_sc_hd__nand2_4
X_77880_ _77880_/A _77880_/B _77880_/X sky130_fd_sc_hd__xor2_4
X_41134_ _41133_/Y _41134_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_404_0_CLK clkbuf_9_202_0_CLK/X _85372_/CLK sky130_fd_sc_hd__clkbuf_1
X_76831_ _76831_/A _76831_/Y sky130_fd_sc_hd__inv_2
X_46991_ _46981_/A _47029_/B _46981_/C _52790_/D _46991_/X sky130_fd_sc_hd__and4_4
X_58977_ _58559_/X _83439_/Q _58976_/Y _58977_/X sky130_fd_sc_hd__o21a_4
X_48730_ _48781_/A _48730_/X sky130_fd_sc_hd__buf_2
X_79550_ _84204_/Q _83252_/Q _79550_/Y sky130_fd_sc_hd__nand2_4
X_45942_ _59539_/A _45943_/A sky130_fd_sc_hd__buf_2
X_57928_ _57926_/X _86003_/Q _57927_/X _57928_/Y sky130_fd_sc_hd__o21ai_4
X_41065_ _40941_/A _41065_/X sky130_fd_sc_hd__buf_2
X_76762_ _76758_/Y _76761_/Y _76762_/Y sky130_fd_sc_hd__nand2_4
X_73974_ _73854_/X _85616_/Q _73903_/X _73973_/X _73974_/X sky130_fd_sc_hd__a211o_4
X_78501_ _82800_/Q _78501_/Y sky130_fd_sc_hd__inv_2
X_75713_ _80914_/Q _75715_/A sky130_fd_sc_hd__inv_2
X_48661_ _48661_/A _48851_/B _48661_/Y sky130_fd_sc_hd__nand2_4
X_72925_ _43131_/Y _72830_/X _72799_/X _72924_/Y _72925_/X sky130_fd_sc_hd__a211o_4
X_79481_ _79481_/A _79480_/Y _79481_/Y sky130_fd_sc_hd__nor2_4
X_45873_ _45869_/X _45872_/X _44898_/X _45873_/X sky130_fd_sc_hd__a21o_4
X_57859_ _57801_/X _57857_/Y _57858_/Y _57822_/X _57809_/X _57859_/X
+ sky130_fd_sc_hd__o32a_4
X_76693_ _76688_/A _76687_/Y _76692_/Y _76694_/B sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_419_0_CLK clkbuf_9_209_0_CLK/X _82463_/CLK sky130_fd_sc_hd__clkbuf_1
X_47612_ _86616_/Q _47570_/X _47611_/Y _47612_/Y sky130_fd_sc_hd__o21ai_4
X_78432_ _78432_/A _82667_/D _78434_/A sky130_fd_sc_hd__xor2_4
X_44824_ _44807_/X _44821_/X _41675_/X _67536_/B _44808_/X _44825_/A
+ sky130_fd_sc_hd__o32ai_4
X_75644_ _75642_/X _75631_/X _75643_/X _75644_/X sky130_fd_sc_hd__a21o_4
X_48592_ _83572_/Q _48593_/A sky130_fd_sc_hd__inv_2
X_60870_ _64191_/B _60870_/X sky130_fd_sc_hd__buf_2
X_72856_ _69619_/B _72853_/X _45897_/X _72855_/Y _72856_/X sky130_fd_sc_hd__a211o_4
X_47543_ _83711_/Q _47543_/Y sky130_fd_sc_hd__inv_2
X_71807_ _71805_/X _83369_/Q _71806_/X _83369_/D sky130_fd_sc_hd__a21o_4
X_59529_ _59521_/A _59876_/B _43995_/A _59609_/D _59529_/X sky130_fd_sc_hd__and4_4
X_78363_ _78359_/X _78364_/C _78362_/Y _78363_/Y sky130_fd_sc_hd__a21oi_4
X_44755_ _44650_/A _44755_/X sky130_fd_sc_hd__buf_2
X_75575_ _75575_/A _80818_/Q _75575_/Y sky130_fd_sc_hd__nand2_4
X_41967_ _41967_/A _41967_/X sky130_fd_sc_hd__buf_2
X_72787_ _72755_/X _83080_/Q _72785_/X _72786_/X _72788_/B sky130_fd_sc_hd__a211o_4
X_77314_ _77315_/A _77315_/B _77315_/C _77316_/A sky130_fd_sc_hd__a21o_4
X_43706_ _87301_/Q _69752_/B sky130_fd_sc_hd__inv_2
X_62540_ _62395_/X _62540_/X sky130_fd_sc_hd__buf_2
X_74526_ _52807_/B _74517_/X _74525_/Y _74526_/Y sky130_fd_sc_hd__o21ai_4
X_40918_ _40918_/A _88311_/D sky130_fd_sc_hd__inv_2
X_47474_ _47474_/A _53070_/D sky130_fd_sc_hd__buf_2
X_71738_ _71735_/D _71738_/X sky130_fd_sc_hd__buf_2
X_78294_ _78301_/A _82472_/Q _78298_/A sky130_fd_sc_hd__xor2_4
X_44686_ _44529_/A _44686_/X sky130_fd_sc_hd__buf_2
X_41898_ _41897_/Y _88110_/D sky130_fd_sc_hd__inv_2
X_49213_ _86432_/Q _48548_/X _49212_/Y _49213_/Y sky130_fd_sc_hd__o21ai_4
X_46425_ _47991_/B _46469_/B _46425_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_93_0_CLK clkbuf_8_93_0_CLK/A clkbuf_8_93_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_77245_ _77245_/A _77243_/X _77245_/C _77261_/A sky130_fd_sc_hd__nand3_4
X_43637_ _40667_/A _43634_/X _68732_/B _43636_/X _43637_/X sky130_fd_sc_hd__a2bb2o_4
X_62471_ _62471_/A _62566_/D sky130_fd_sc_hd__buf_2
X_74457_ _83062_/Q _74441_/X _74456_/Y _74457_/Y sky130_fd_sc_hd__o21ai_4
X_40849_ _40848_/X _40849_/X sky130_fd_sc_hd__buf_2
X_71669_ _71669_/A _71669_/X sky130_fd_sc_hd__buf_2
X_64210_ _64210_/A _64457_/C _64208_/Y _64209_/Y _64210_/Y sky130_fd_sc_hd__nand4_4
X_61422_ _64292_/A _61452_/B _61452_/C _61391_/D _61422_/Y sky130_fd_sc_hd__nand4_4
X_49144_ _49144_/A _49144_/X sky130_fd_sc_hd__buf_2
X_73408_ _73359_/X _83056_/Q _73406_/X _73407_/X _73408_/X sky130_fd_sc_hd__a211o_4
X_46356_ _53985_/B _46356_/X sky130_fd_sc_hd__buf_2
X_65190_ _65753_/A _86443_/Q _65190_/X sky130_fd_sc_hd__and2_4
X_77176_ _77159_/Y _77173_/X _77175_/Y _77177_/B sky130_fd_sc_hd__a21oi_4
X_43568_ _43568_/A _43568_/Y sky130_fd_sc_hd__inv_2
X_74388_ _72052_/A _74466_/A sky130_fd_sc_hd__buf_2
X_45307_ _45304_/X _45306_/Y _45275_/X _45307_/Y sky130_fd_sc_hd__a21oi_4
X_64141_ _64137_/Y _64129_/X _64140_/Y _64141_/Y sky130_fd_sc_hd__a21oi_4
X_76127_ _76125_/X _76127_/B _76126_/Y _76127_/X sky130_fd_sc_hd__and3_4
X_42519_ _42556_/A _42519_/X sky130_fd_sc_hd__buf_2
X_49075_ _65100_/B _49052_/X _49074_/Y _49075_/Y sky130_fd_sc_hd__o21ai_4
X_61353_ _61346_/X _61349_/X _61352_/Y _84488_/D sky130_fd_sc_hd__a21oi_4
X_73339_ _73339_/A _73339_/B _73339_/Y sky130_fd_sc_hd__nor2_4
X_46287_ _51251_/B _53959_/B sky130_fd_sc_hd__buf_2
X_43499_ _43466_/X _43499_/X sky130_fd_sc_hd__buf_2
X_48026_ _82351_/Q _47973_/B _48026_/X sky130_fd_sc_hd__or2_4
X_60304_ _60304_/A _60337_/C sky130_fd_sc_hd__buf_2
X_45238_ _55783_/B _45206_/X _45237_/X _45238_/X sky130_fd_sc_hd__o21a_4
X_64072_ _64064_/X _64048_/X _64066_/Y _64069_/Y _64071_/X _64072_/X
+ sky130_fd_sc_hd__a41o_4
X_76058_ _81716_/D _76058_/B _76058_/Y sky130_fd_sc_hd__nand2_4
X_61284_ _61283_/Y _60596_/A _61284_/Y sky130_fd_sc_hd__nor2_4
X_67900_ _81482_/D _67806_/X _67899_/X _84050_/D sky130_fd_sc_hd__a21bo_4
X_63023_ _63021_/Y _63022_/X _61194_/X _63023_/Y sky130_fd_sc_hd__a21oi_4
X_75009_ _75008_/A _75008_/B _75021_/B sky130_fd_sc_hd__nand2_4
X_60235_ _60235_/A _60259_/B sky130_fd_sc_hd__inv_2
X_45169_ _45169_/A _45182_/B _45169_/Y sky130_fd_sc_hd__nand2_4
X_68880_ _68666_/X _68612_/X _68867_/Y _68879_/Y _68880_/X sky130_fd_sc_hd__a211o_4
X_67831_ _67354_/X _67831_/X sky130_fd_sc_hd__buf_2
X_79817_ _79817_/A _79817_/B _79817_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_8_31_0_CLK clkbuf_8_31_0_CLK/A clkbuf_9_63_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_60166_ _60165_/X _60166_/X sky130_fd_sc_hd__buf_2
X_49977_ _40595_/X _49977_/X sky130_fd_sc_hd__buf_2
X_48928_ _48928_/A _48894_/B _48928_/C _48928_/X sky130_fd_sc_hd__and3_4
X_67762_ _67690_/X _87713_/Q _67762_/X sky130_fd_sc_hd__and2_4
X_79748_ _79734_/Y _79731_/Y _79748_/X sky130_fd_sc_hd__and2_4
X_64974_ _65074_/A _64974_/B _64974_/X sky130_fd_sc_hd__and2_4
X_60097_ _60081_/A _60103_/B _60097_/C _60097_/Y sky130_fd_sc_hd__nor3_4
X_69501_ _69013_/X _69016_/X _69500_/X _69501_/Y sky130_fd_sc_hd__a21oi_4
X_66713_ _87437_/Q _66642_/X _66643_/X _66712_/X _66713_/X sky130_fd_sc_hd__a211o_4
X_63925_ _64184_/C _63958_/C sky130_fd_sc_hd__buf_2
X_48859_ _48680_/A _48859_/B _48854_/C _48859_/X sky130_fd_sc_hd__and3_4
X_67693_ _67615_/X _67693_/B _67693_/X sky130_fd_sc_hd__and2_4
X_79679_ _84214_/Q _83262_/Q _79679_/X sky130_fd_sc_hd__xor2_4
X_81710_ _88121_/CLK _81710_/D _41043_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_46_0_CLK clkbuf_8_47_0_CLK/A clkbuf_9_93_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_69432_ _87018_/Q _69414_/X _69430_/X _69431_/X _69432_/X sky130_fd_sc_hd__a211o_4
X_66644_ _68999_/A _66644_/B _66644_/X sky130_fd_sc_hd__and2_4
X_51870_ _51870_/A _51870_/B _51870_/C _52698_/D _51870_/X sky130_fd_sc_hd__and4_4
X_63856_ _64045_/A _63920_/D sky130_fd_sc_hd__buf_2
X_82690_ _81216_/CLK _78805_/X _82678_/D sky130_fd_sc_hd__dfxtp_4
X_50821_ _50728_/A _50822_/A sky130_fd_sc_hd__buf_2
X_62807_ _62805_/X _62779_/X _62806_/Y _84381_/D sky130_fd_sc_hd__a21oi_4
X_81641_ _81671_/CLK _81673_/Q _81641_/Q sky130_fd_sc_hd__dfxtp_4
X_69363_ _87023_/Q _69239_/X _69361_/X _69362_/X _69363_/X sky130_fd_sc_hd__a211o_4
X_66575_ _66553_/X _68742_/A sky130_fd_sc_hd__buf_2
X_63787_ _61367_/A _63772_/B _63721_/C _63787_/D _63787_/Y sky130_fd_sc_hd__nand4_4
X_60999_ _60996_/Y _60998_/X _60895_/X _60901_/X _60999_/X sky130_fd_sc_hd__a211o_4
X_68314_ _82633_/D _68299_/X _68313_/X _68314_/X sky130_fd_sc_hd__a21bo_4
X_53540_ _53448_/X _53540_/X sky130_fd_sc_hd__buf_2
X_65526_ _65524_/X _83075_/Q _65391_/X _65525_/X _65526_/X sky130_fd_sc_hd__a211o_4
X_84360_ _84360_/CLK _84360_/D _79502_/A sky130_fd_sc_hd__dfxtp_4
X_50752_ _50749_/Y _50676_/X _50751_/X _50752_/Y sky130_fd_sc_hd__a21oi_4
X_62738_ _62711_/A _64295_/C _62737_/X _62738_/D _62738_/X sky130_fd_sc_hd__and4_4
X_81572_ _81587_/CLK _84172_/Q _76675_/A sky130_fd_sc_hd__dfxtp_4
X_69294_ _67013_/X _69575_/A sky130_fd_sc_hd__buf_2
X_83311_ _83311_/CLK _71971_/Y _83311_/Q sky130_fd_sc_hd__dfxtp_4
X_80523_ _84767_/Q _84159_/Q _80523_/Y sky130_fd_sc_hd__nand2_4
X_68245_ _84002_/Q _68238_/X _68244_/X _84002_/D sky130_fd_sc_hd__a21bo_4
X_53471_ _53798_/A _53982_/A sky130_fd_sc_hd__buf_2
X_65457_ _64851_/A _65457_/X sky130_fd_sc_hd__buf_2
X_84291_ _84671_/CLK _63851_/Y _84291_/Q sky130_fd_sc_hd__dfxtp_4
X_50683_ _86154_/Q _50680_/X _50682_/Y _50683_/Y sky130_fd_sc_hd__o21ai_4
X_62669_ _62669_/A _63022_/A _62927_/A _62669_/D _62669_/X sky130_fd_sc_hd__and4_4
X_55210_ _72712_/C _55209_/X _83317_/Q _55288_/A sky130_fd_sc_hd__a21o_4
X_86030_ _86030_/CLK _86030_/D _65105_/B sky130_fd_sc_hd__dfxtp_4
X_52422_ _52324_/A _52422_/X sky130_fd_sc_hd__buf_2
X_64408_ _79713_/B _64373_/X _64407_/X _64408_/X sky130_fd_sc_hd__a21o_4
X_83242_ _83242_/CLK _83242_/D _62081_/B sky130_fd_sc_hd__dfxtp_4
X_80454_ _84761_/Q _84153_/Q _80456_/A sky130_fd_sc_hd__xor2_4
X_56190_ _56252_/A _56280_/A sky130_fd_sc_hd__buf_2
X_68176_ _82060_/D _68160_/X _68175_/X _68176_/X sky130_fd_sc_hd__a21bo_4
X_65388_ _65059_/X _85539_/Q _65060_/X _65387_/X _65388_/X sky130_fd_sc_hd__a211o_4
X_55141_ _55125_/A _55142_/A sky130_fd_sc_hd__buf_2
X_67127_ _67126_/X _67149_/A sky130_fd_sc_hd__buf_2
X_52353_ _52349_/A _50144_/B _52353_/Y sky130_fd_sc_hd__nand2_4
X_64339_ _64331_/Y _64338_/X _64328_/X _64339_/X sky130_fd_sc_hd__o21a_4
X_83173_ _84980_/CLK _83173_/D _83173_/Q sky130_fd_sc_hd__dfxtp_4
X_80385_ _80361_/A _80384_/D _80382_/X _80385_/X sky130_fd_sc_hd__a21bo_4
X_51304_ _51296_/A _46412_/B _51304_/Y sky130_fd_sc_hd__nand2_4
X_82124_ _82124_/CLK _82124_/D _82124_/Q sky130_fd_sc_hd__dfxtp_4
X_55072_ _55072_/A _55072_/X sky130_fd_sc_hd__buf_2
X_67058_ _87871_/Q _67056_/X _67032_/X _67057_/X _67058_/X sky130_fd_sc_hd__a211o_4
X_52284_ _64719_/B _52269_/X _52283_/Y _52284_/Y sky130_fd_sc_hd__o21ai_4
X_87981_ _87144_/CLK _42203_/Y _87981_/Q sky130_fd_sc_hd__dfxtp_4
X_58900_ _58810_/A _58900_/X sky130_fd_sc_hd__buf_2
X_54023_ _54021_/Y _54006_/X _54022_/Y _85521_/D sky130_fd_sc_hd__a21boi_4
X_66009_ _64722_/X _85626_/Q _64724_/X _66008_/X _66009_/X sky130_fd_sc_hd__a211o_4
X_51235_ _51240_/A _51235_/B _51235_/Y sky130_fd_sc_hd__nand2_4
X_86932_ _86932_/CLK _86932_/D _67605_/B sky130_fd_sc_hd__dfxtp_4
X_82055_ _83933_/CLK _82055_/D _77780_/B sky130_fd_sc_hd__dfxtp_4
X_59880_ _60418_/D _60174_/D _60407_/A _59552_/C _59880_/X sky130_fd_sc_hd__and4_4
X_81006_ _82515_/CLK _84214_/Q _81006_/Q sky130_fd_sc_hd__dfxtp_4
X_58831_ _86700_/Q _58873_/B _58831_/Y sky130_fd_sc_hd__nor2_4
X_51166_ _51163_/Y _51147_/X _51165_/X _51166_/Y sky130_fd_sc_hd__a21oi_4
X_86863_ _86861_/CLK _45658_/Y _63196_/B sky130_fd_sc_hd__dfxtp_4
X_50117_ _50092_/A _50117_/X sky130_fd_sc_hd__buf_2
X_85814_ _85815_/CLK _52479_/Y _85814_/Q sky130_fd_sc_hd__dfxtp_4
X_58762_ _58758_/Y _58760_/Y _58761_/X _58762_/X sky130_fd_sc_hd__a21o_4
X_51097_ _51097_/A _52787_/B _51097_/Y sky130_fd_sc_hd__nand2_4
X_55974_ _55974_/A _55974_/B _55975_/A sky130_fd_sc_hd__and2_4
X_86794_ _88245_/CLK _46051_/Y _86794_/Q sky130_fd_sc_hd__dfxtp_4
X_57713_ _57712_/X _85729_/Q _44252_/X _57713_/X sky130_fd_sc_hd__o21a_4
X_50048_ _50048_/A _53259_/B _50048_/Y sky130_fd_sc_hd__nand2_4
X_54925_ _85352_/Q _54918_/X _54924_/Y _54925_/Y sky130_fd_sc_hd__o21ai_4
X_85745_ _85745_/CLK _52842_/Y _85745_/Q sky130_fd_sc_hd__dfxtp_4
X_58693_ _58618_/X _86103_/Q _58692_/X _58693_/Y sky130_fd_sc_hd__o21ai_4
X_70971_ _70944_/A _70976_/A sky130_fd_sc_hd__buf_2
X_82957_ _82769_/CLK _82957_/D _82957_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_390_0_CLK clkbuf_9_195_0_CLK/X _83231_/CLK sky130_fd_sc_hd__clkbuf_1
X_72710_ _72710_/A _44907_/A _55285_/A _55274_/X _72710_/X sky130_fd_sc_hd__and4_4
X_57644_ _71970_/A _50385_/B _57644_/Y sky130_fd_sc_hd__nand2_4
X_81908_ _82133_/CLK _81908_/D _82284_/D sky130_fd_sc_hd__dfxtp_4
X_54856_ _54882_/A _54856_/X sky130_fd_sc_hd__buf_2
X_42870_ _42870_/A _42870_/Y sky130_fd_sc_hd__inv_2
X_73690_ _73665_/X _84988_/Q _73614_/X _73689_/X _73690_/X sky130_fd_sc_hd__a211o_4
X_85676_ _84802_/CLK _85676_/D _85676_/Q sky130_fd_sc_hd__dfxtp_4
X_82888_ _82888_/CLK _78123_/B _82888_/Q sky130_fd_sc_hd__dfxtp_4
X_87415_ _87417_/CLK _87415_/D _87415_/Q sky130_fd_sc_hd__dfxtp_4
X_41821_ _41607_/X _41821_/X sky130_fd_sc_hd__buf_2
X_53807_ _53804_/Y _53773_/X _53806_/X _85565_/D sky130_fd_sc_hd__a21oi_4
X_72641_ _72633_/X _72643_/B _72641_/C _72641_/Y sky130_fd_sc_hd__nand3_4
X_84627_ _84624_/CLK _60342_/X _79649_/A sky130_fd_sc_hd__dfxtp_4
X_57575_ _84976_/Q _57550_/X _57574_/Y _57575_/Y sky130_fd_sc_hd__o21ai_4
X_81839_ _81839_/CLK _81839_/D _77409_/A sky130_fd_sc_hd__dfxtp_4
X_88395_ _86824_/CLK _88395_/D _88395_/Q sky130_fd_sc_hd__dfxtp_4
X_54787_ _85378_/Q _54784_/X _54786_/Y _54787_/Y sky130_fd_sc_hd__o21ai_4
X_51999_ _51982_/X _53520_/B _51999_/Y sky130_fd_sc_hd__nand2_4
X_59314_ _59310_/Y _59313_/Y _59278_/X _59314_/X sky130_fd_sc_hd__a21o_4
X_44540_ _44529_/X _44530_/X _40810_/A _44539_/Y _44533_/X _44540_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56526_ _56533_/A _56533_/B _85162_/Q _56526_/Y sky130_fd_sc_hd__nand3_4
X_75360_ _75360_/A _75362_/A sky130_fd_sc_hd__inv_2
X_41752_ _41749_/X _41750_/X _67885_/B _41751_/X _88156_/D sky130_fd_sc_hd__a2bb2o_4
X_87346_ _87345_/CLK _43598_/Y _43596_/A sky130_fd_sc_hd__dfxtp_4
X_53738_ _53763_/A _53748_/C sky130_fd_sc_hd__buf_2
X_72572_ _72572_/A _72572_/B _72572_/X sky130_fd_sc_hd__and2_4
X_84558_ _83216_/CLK _60824_/Y _60822_/C sky130_fd_sc_hd__dfxtp_4
X_74311_ _83103_/Q _74301_/X _74310_/Y _74311_/X sky130_fd_sc_hd__a21bo_4
X_40703_ _40687_/X _40688_/X _40702_/X _88351_/Q _40683_/X _40703_/Y
+ sky130_fd_sc_hd__o32ai_4
X_59245_ _59245_/A _59282_/B _59245_/Y sky130_fd_sc_hd__nor2_4
X_71523_ _71521_/A _70724_/A _71523_/Y sky130_fd_sc_hd__nand2_4
X_83509_ _83508_/CLK _83509_/D _83509_/Q sky130_fd_sc_hd__dfxtp_4
X_44471_ _44447_/X _44448_/X _41173_/X _87091_/Q _44449_/X _44472_/A
+ sky130_fd_sc_hd__o32ai_4
X_56457_ _56279_/A _57364_/D _56174_/X _56459_/A sky130_fd_sc_hd__nand3_4
X_75291_ _75287_/Y _75288_/Y _75291_/C _75291_/X sky130_fd_sc_hd__or3_4
X_87277_ _88087_/CLK _43764_/X _87277_/Q sky130_fd_sc_hd__dfxtp_4
X_41683_ _40565_/Y _41814_/A sky130_fd_sc_hd__buf_2
X_53669_ _53662_/X _74414_/B _53669_/Y sky130_fd_sc_hd__nand2_4
X_84489_ _83218_/CLK _84489_/D _84489_/Q sky130_fd_sc_hd__dfxtp_4
X_46210_ _46210_/A _69611_/A sky130_fd_sc_hd__buf_2
XPHY_220 sky130_fd_sc_hd__decap_3
X_77030_ _77023_/A _77023_/B _77030_/Y sky130_fd_sc_hd__nand2_4
X_43422_ _43518_/A _43422_/X sky130_fd_sc_hd__buf_2
X_55408_ _55403_/A _55408_/B _55403_/B _55415_/B sky130_fd_sc_hd__nand3_4
X_86228_ _86578_/CLK _50301_/Y _86228_/Q sky130_fd_sc_hd__dfxtp_4
X_74242_ _74202_/A _74241_/Y _74242_/Y sky130_fd_sc_hd__nor2_4
XPHY_231 sky130_fd_sc_hd__decap_3
X_40634_ _40633_/X _40596_/X _88363_/Q _40599_/X _88363_/D sky130_fd_sc_hd__a2bb2o_4
X_47190_ _47152_/X _47181_/B _47210_/C _51214_/D _47190_/X sky130_fd_sc_hd__and4_4
X_59176_ _59121_/X _85427_/Q _59175_/X _59176_/Y sky130_fd_sc_hd__o21ai_4
X_71454_ _70682_/A _71626_/C _71450_/C _71454_/Y sky130_fd_sc_hd__nor3_4
X_56388_ _56383_/X _56386_/B _85213_/Q _56388_/Y sky130_fd_sc_hd__nand3_4
XPHY_242 sky130_fd_sc_hd__decap_3
XPHY_253 sky130_fd_sc_hd__decap_3
XPHY_264 sky130_fd_sc_hd__decap_3
X_46141_ _46141_/A _46143_/B sky130_fd_sc_hd__inv_2
X_58127_ _58125_/X _85699_/Q _58126_/X _58127_/X sky130_fd_sc_hd__o21a_4
X_70405_ _71090_/A _70824_/A sky130_fd_sc_hd__buf_2
XPHY_275 sky130_fd_sc_hd__decap_3
X_43353_ _43329_/X _43353_/X sky130_fd_sc_hd__buf_2
X_55339_ _55336_/X _55365_/B _83752_/Q _55445_/B sky130_fd_sc_hd__a21o_4
X_74173_ _74080_/X _86215_/Q _74103_/X _74172_/X _74173_/X sky130_fd_sc_hd__a211o_4
X_86159_ _86256_/CLK _86159_/D _86159_/Q sky130_fd_sc_hd__dfxtp_4
X_40565_ _40344_/A _42446_/A _48162_/A _40565_/Y sky130_fd_sc_hd__a21oi_4
XPHY_286 sky130_fd_sc_hd__decap_3
X_71385_ _71163_/A _71386_/B sky130_fd_sc_hd__buf_2
XPHY_297 sky130_fd_sc_hd__decap_3
X_42304_ _41909_/Y _42304_/X sky130_fd_sc_hd__buf_2
X_73124_ _73124_/A _73124_/B _73124_/Y sky130_fd_sc_hd__nor2_4
X_70336_ _70320_/X _83793_/Q _70335_/X _83793_/D sky130_fd_sc_hd__a21o_4
X_46072_ _41585_/Y _46061_/X _86782_/Q _46062_/X _86782_/D sky130_fd_sc_hd__a2bb2o_4
X_58058_ _58070_/A _58058_/B _58058_/Y sky130_fd_sc_hd__nor2_4
X_43284_ _41157_/X _43277_/X _87499_/Q _43278_/X _87499_/D sky130_fd_sc_hd__a2bb2o_4
X_78981_ _78986_/B _78981_/B _78982_/B sky130_fd_sc_hd__xor2_4
X_40496_ _40325_/X _82316_/Q _40495_/X _40496_/Y sky130_fd_sc_hd__o21ai_4
X_49900_ _49896_/Y _49897_/X _49899_/X _49900_/Y sky130_fd_sc_hd__a21oi_4
X_45023_ _44975_/X _61417_/B _44995_/X _45023_/Y sky130_fd_sc_hd__o21ai_4
X_57009_ _56783_/X _56737_/X _56785_/D _57024_/D _57010_/A _57009_/Y
+ sky130_fd_sc_hd__a41oi_4
X_42235_ _42234_/Y _87968_/D sky130_fd_sc_hd__inv_2
X_77932_ _77916_/B _77929_/X _77931_/Y _77933_/B sky130_fd_sc_hd__a21oi_4
X_73055_ _72798_/X _73055_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_343_0_CLK clkbuf_9_171_0_CLK/X _85741_/CLK sky130_fd_sc_hd__clkbuf_1
X_70267_ _70267_/A _70267_/B _70267_/C _70264_/X _70267_/X sky130_fd_sc_hd__and4_4
X_60020_ _59842_/A _60064_/A sky130_fd_sc_hd__buf_2
X_72006_ _72004_/Y _71978_/X _72005_/X _72006_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_973_0_CLK clkbuf_9_486_0_CLK/X _85547_/CLK sky130_fd_sc_hd__clkbuf_1
X_49831_ _49829_/Y _49815_/X _49830_/X _49831_/Y sky130_fd_sc_hd__a21oi_4
X_42166_ _42166_/A _42166_/Y sky130_fd_sc_hd__inv_2
X_77863_ _82065_/Q _77863_/Y sky130_fd_sc_hd__inv_2
X_70198_ _70200_/A _70200_/B _70198_/C _70200_/D _70198_/X sky130_fd_sc_hd__and4_4
X_79602_ _65294_/C _83255_/Q _79602_/X sky130_fd_sc_hd__or2_4
X_41117_ _41112_/X _41113_/X _41116_/X _88275_/Q _41088_/X _41118_/A
+ sky130_fd_sc_hd__o32ai_4
X_76814_ _76801_/A _76808_/A _76814_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_464_0_CLK clkbuf_8_232_0_CLK/X clkbuf_9_464_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_49762_ _49758_/Y _49759_/X _49761_/X _49762_/Y sky130_fd_sc_hd__a21oi_4
X_46974_ _46970_/Y _46940_/X _46973_/X _86684_/D sky130_fd_sc_hd__a21oi_4
X_42097_ _42083_/X _42094_/X _41016_/X _88037_/Q _42096_/X _42097_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77794_ _82266_/Q _81978_/Q _77819_/A sky130_fd_sc_hd__xnor2_4
X_48713_ _48725_/A _48358_/X _48713_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_358_0_CLK clkbuf_9_179_0_CLK/X _85709_/CLK sky130_fd_sc_hd__clkbuf_1
X_79533_ _79895_/A _79531_/X _79532_/Y _79547_/A sky130_fd_sc_hd__a21boi_4
X_45925_ _65034_/A _64656_/A sky130_fd_sc_hd__buf_2
X_41048_ _41048_/A _41091_/B _41048_/X sky130_fd_sc_hd__or2_4
X_76745_ _76745_/A _76745_/B _76745_/X sky130_fd_sc_hd__xor2_4
X_49693_ _49691_/Y _49677_/X _49692_/X _49693_/Y sky130_fd_sc_hd__a21oi_4
X_61971_ _61969_/X _61924_/B _61971_/C _61971_/D _61971_/Y sky130_fd_sc_hd__nand4_4
X_73957_ _53535_/B _73957_/B _73957_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_10_988_0_CLK clkbuf_9_494_0_CLK/X _86256_/CLK sky130_fd_sc_hd__clkbuf_1
X_63710_ _63701_/A _63701_/B _80279_/B _63710_/Y sky130_fd_sc_hd__nor3_4
X_60922_ _64172_/B _60994_/B sky130_fd_sc_hd__buf_2
X_48644_ _48644_/A _48845_/A sky130_fd_sc_hd__buf_2
X_72908_ _72908_/A _72908_/X sky130_fd_sc_hd__buf_2
X_79464_ _79455_/X _79457_/B _79464_/Y sky130_fd_sc_hd__nand2_4
X_45856_ _85027_/Q _45856_/Y sky130_fd_sc_hd__inv_2
X_64690_ _64687_/Y _64662_/X _64689_/Y _64690_/X sky130_fd_sc_hd__a21o_4
X_76676_ _81477_/Q _76686_/A sky130_fd_sc_hd__inv_2
X_73888_ _73886_/X _73888_/B _73888_/C _73888_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_9_479_0_CLK clkbuf_9_479_0_CLK/A clkbuf_9_479_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_78415_ _78413_/Y _78414_/Y _82761_/D sky130_fd_sc_hd__xnor2_4
X_44807_ _45980_/A _44807_/X sky130_fd_sc_hd__buf_2
X_63641_ _62083_/D _60780_/X _63358_/X _60767_/X _63640_/Y _63641_/X
+ sky130_fd_sc_hd__a2111o_4
X_75627_ _75632_/A _75632_/B _75628_/B sky130_fd_sc_hd__xor2_4
X_48575_ _81774_/Q _48576_/A sky130_fd_sc_hd__inv_2
X_60853_ _60851_/X _60852_/X _63632_/A _60853_/X sky130_fd_sc_hd__and3_4
X_72839_ _73092_/A _72839_/X sky130_fd_sc_hd__buf_2
X_79395_ _79395_/A _79395_/B _79396_/B sky130_fd_sc_hd__xnor2_4
X_45787_ _45787_/A _45746_/B _45787_/Y sky130_fd_sc_hd__nand2_4
X_42999_ _40507_/X _42994_/X _87612_/Q _42995_/X _87612_/D sky130_fd_sc_hd__a2bb2o_4
X_47526_ _47526_/A _47526_/Y sky130_fd_sc_hd__inv_2
X_66360_ _66358_/Y _66343_/X _66359_/X _84138_/D sky130_fd_sc_hd__a21o_4
Xclkbuf_10_911_0_CLK clkbuf_9_455_0_CLK/X _87595_/CLK sky130_fd_sc_hd__clkbuf_1
X_78346_ _78343_/Y _82789_/Q _78344_/Y _78346_/Y sky130_fd_sc_hd__nand3_4
X_44738_ _44738_/A _44738_/Y sky130_fd_sc_hd__inv_2
X_63572_ _60738_/Y _63630_/C sky130_fd_sc_hd__buf_2
X_75558_ _75558_/A _75557_/X _75559_/B sky130_fd_sc_hd__xnor2_4
X_60784_ _60652_/X _63384_/D sky130_fd_sc_hd__buf_2
Xclkbuf_10_0_0_CLK clkbuf_9_0_0_CLK/X _85270_/CLK sky130_fd_sc_hd__clkbuf_1
X_65311_ _65308_/X _86726_/Q _65309_/X _65310_/X _65311_/X sky130_fd_sc_hd__a211o_4
X_62523_ _62463_/A _62623_/D sky130_fd_sc_hd__buf_2
X_74509_ _74509_/A _74509_/B _74509_/C _74509_/X sky130_fd_sc_hd__and3_4
X_47457_ _47453_/Y _47414_/X _47456_/X _47457_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_402_0_CLK clkbuf_9_402_0_CLK/A clkbuf_9_402_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_66291_ _66282_/X _65827_/Y _66290_/Y _66291_/Y sky130_fd_sc_hd__o21ai_4
X_78277_ _78274_/Y _78276_/Y _78278_/B sky130_fd_sc_hd__xor2_4
X_44669_ _44658_/X _44659_/X _40560_/X _87007_/Q _44660_/X _44669_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75489_ _75485_/X _75486_/A _75491_/C sky130_fd_sc_hd__nand2_4
X_68030_ _68451_/A _68405_/A sky130_fd_sc_hd__buf_2
X_46408_ _46408_/A _46407_/X _46408_/Y sky130_fd_sc_hd__nand2_4
X_65242_ _65238_/X _65111_/B _65241_/X _65242_/Y sky130_fd_sc_hd__nand3_4
X_77228_ _77230_/A _77230_/C _77228_/X sky130_fd_sc_hd__and2_4
X_62454_ _62444_/X _62451_/Y _62453_/X _84849_/Q _62440_/X _62454_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47388_ _86640_/Q _47382_/X _47387_/Y _47388_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_926_0_CLK clkbuf_9_463_0_CLK/X _83161_/CLK sky130_fd_sc_hd__clkbuf_1
X_49127_ _86441_/Q _49104_/X _49126_/Y _49127_/Y sky130_fd_sc_hd__o21ai_4
X_61405_ _72529_/C _61406_/C sky130_fd_sc_hd__buf_2
X_46339_ _46339_/A _53978_/B sky130_fd_sc_hd__buf_2
X_65173_ _65155_/A _85803_/Q _65173_/X sky130_fd_sc_hd__and2_4
X_77159_ _77159_/A _77159_/B _77159_/Y sky130_fd_sc_hd__nand2_4
X_62385_ _62344_/X _57670_/A _62565_/C _62355_/X _62385_/X sky130_fd_sc_hd__and4_4
X_64124_ _64118_/Y _64120_/Y _64122_/Y _64123_/Y _64124_/X sky130_fd_sc_hd__and4_4
Xclkbuf_9_417_0_CLK clkbuf_8_208_0_CLK/X clkbuf_9_417_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_49058_ _46447_/B _48699_/B _49058_/Y sky130_fd_sc_hd__nand2_4
X_61336_ _72529_/C _61367_/C sky130_fd_sc_hd__buf_2
X_80170_ _80156_/Y _80162_/B _80169_/X _80171_/B sky130_fd_sc_hd__o21ai_4
X_69981_ _68391_/X _68398_/X _69925_/X _69981_/Y sky130_fd_sc_hd__a21oi_4
X_48009_ _48542_/B _47915_/B _48009_/Y sky130_fd_sc_hd__nand2_4
X_64055_ _64074_/A _64074_/B _80049_/B _64055_/Y sky130_fd_sc_hd__nor3_4
X_68932_ _87580_/Q _68715_/X _66349_/X _68931_/X _68932_/X sky130_fd_sc_hd__a211o_4
X_61267_ _61109_/X _61198_/X _61095_/X _61267_/Y sky130_fd_sc_hd__o21ai_4
X_51020_ _51101_/A _51020_/X sky130_fd_sc_hd__buf_2
Xclkbuf_6_2_0_CLK clkbuf_6_3_0_CLK/A clkbuf_6_2_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_63006_ _63285_/A _63285_/B _79513_/A _63006_/Y sky130_fd_sc_hd__nor3_4
X_60218_ _60218_/A _60344_/B sky130_fd_sc_hd__buf_2
X_68863_ _68860_/X _68862_/X _68748_/X _68863_/X sky130_fd_sc_hd__a21o_4
X_61198_ _64545_/A _61198_/X sky130_fd_sc_hd__buf_2
X_67814_ _86955_/Q _67788_/X _67789_/X _67813_/X _67814_/X sky130_fd_sc_hd__a211o_4
X_60149_ _59875_/X _60118_/X _60073_/Y _59951_/Y _60148_/Y _60149_/X
+ sky130_fd_sc_hd__o41a_4
X_83860_ _82541_/CLK _70062_/X _82540_/D sky130_fd_sc_hd__dfxtp_4
X_68794_ _87490_/Q _68792_/X _68545_/X _68793_/X _68794_/X sky130_fd_sc_hd__a211o_4
X_82811_ _82692_/CLK _82843_/Q _82811_/Q sky130_fd_sc_hd__dfxtp_4
X_67745_ _87150_/Q _67670_/X _67671_/X _67744_/X _67745_/X sky130_fd_sc_hd__a211o_4
X_52971_ _52947_/X _52982_/B _52977_/C _52971_/D _52971_/X sky130_fd_sc_hd__and4_4
X_64957_ _65002_/A _86036_/Q _64957_/X sky130_fd_sc_hd__and2_4
X_83791_ _81631_/CLK _83791_/D _74786_/A sky130_fd_sc_hd__dfxtp_4
X_54710_ _85392_/Q _54703_/X _54709_/Y _54710_/Y sky130_fd_sc_hd__o21ai_4
X_85530_ _85818_/CLK _85530_/D _85530_/Q sky130_fd_sc_hd__dfxtp_4
X_51922_ _52322_/A _51922_/X sky130_fd_sc_hd__buf_2
X_63908_ _61448_/X _63908_/B _63894_/C _63908_/D _63908_/Y sky130_fd_sc_hd__nand4_4
X_82742_ _82147_/CLK _84126_/Q _78994_/A sky130_fd_sc_hd__dfxtp_4
X_55690_ _55690_/A _55690_/X sky130_fd_sc_hd__buf_2
X_67676_ _87909_/Q _67651_/X _67625_/X _67675_/X _67676_/X sky130_fd_sc_hd__a211o_4
X_64888_ _64885_/X _64888_/B _64887_/X _64888_/Y sky130_fd_sc_hd__nand3_4
X_69415_ _69309_/A _69415_/B _69415_/X sky130_fd_sc_hd__and2_4
X_54641_ _54636_/A _54121_/B _54641_/Y sky130_fd_sc_hd__nand2_4
X_66627_ _87953_/Q _66562_/X _66564_/X _66626_/X _66627_/X sky130_fd_sc_hd__a211o_4
X_85461_ _82769_/CLK _54335_/Y _85461_/Q sky130_fd_sc_hd__dfxtp_4
X_51853_ _51853_/A _50987_/B _51853_/Y sky130_fd_sc_hd__nand2_4
X_63839_ _63724_/A _63840_/C sky130_fd_sc_hd__buf_2
X_82673_ _82715_/CLK _82673_/D _82673_/Q sky130_fd_sc_hd__dfxtp_4
X_87200_ _87708_/CLK _87200_/D _87200_/Q sky130_fd_sc_hd__dfxtp_4
X_84412_ _84414_/CLK _84412_/D _84412_/Q sky130_fd_sc_hd__dfxtp_4
X_50804_ _50742_/A _50804_/X sky130_fd_sc_hd__buf_2
X_57360_ _57358_/X _57247_/Y _57359_/Y _85029_/D sky130_fd_sc_hd__a21oi_4
X_81624_ _81696_/CLK _76485_/X _81624_/Q sky130_fd_sc_hd__dfxtp_4
X_69346_ _64806_/A _69346_/X sky130_fd_sc_hd__buf_2
X_88180_ _88180_/CLK _41627_/X _67324_/B sky130_fd_sc_hd__dfxtp_4
X_54572_ _54570_/Y _54558_/X _54571_/X _54572_/Y sky130_fd_sc_hd__a21oi_4
X_66558_ _87135_/Q _66550_/X _66552_/X _66557_/X _66559_/B sky130_fd_sc_hd__a211o_4
X_85392_ _85489_/CLK _85392_/D _85392_/Q sky130_fd_sc_hd__dfxtp_4
X_51784_ _51779_/A _46685_/X _51784_/Y sky130_fd_sc_hd__nand2_4
X_56311_ _45369_/A _56351_/A sky130_fd_sc_hd__buf_2
X_87131_ _87484_/CLK _44393_/X _87131_/Q sky130_fd_sc_hd__dfxtp_4
X_65509_ _65416_/X _86524_/Q _65509_/X sky130_fd_sc_hd__and2_4
X_53523_ _85620_/Q _53506_/X _53522_/Y _53523_/Y sky130_fd_sc_hd__o21ai_4
X_84343_ _84849_/CLK _63222_/X _79321_/A sky130_fd_sc_hd__dfxtp_4
X_50735_ _50768_/A _50735_/X sky130_fd_sc_hd__buf_2
X_57291_ _56726_/X _57268_/X _56739_/X _56740_/X _56852_/A _57291_/Y
+ sky130_fd_sc_hd__a41oi_4
X_81555_ _84087_/CLK _76809_/X _81511_/D sky130_fd_sc_hd__dfxtp_4
X_69277_ _69182_/A _69277_/X sky130_fd_sc_hd__buf_2
X_66489_ _65464_/A _66501_/B sky130_fd_sc_hd__buf_2
X_59030_ _59030_/A _59008_/B _59030_/Y sky130_fd_sc_hd__nor2_4
X_56242_ _56255_/A _56242_/X sky130_fd_sc_hd__buf_2
X_80506_ _80506_/A _80506_/B _80506_/X sky130_fd_sc_hd__xor2_4
X_68228_ _68168_/A _68228_/X sky130_fd_sc_hd__buf_2
X_87062_ _87063_/CLK _44540_/Y _44539_/A sky130_fd_sc_hd__dfxtp_4
X_53454_ _85632_/Q _53449_/X _53453_/Y _53454_/Y sky130_fd_sc_hd__o21ai_4
X_84274_ _84273_/CLK _84274_/D _64108_/C sky130_fd_sc_hd__dfxtp_4
X_50666_ _50657_/A _50153_/B _50666_/Y sky130_fd_sc_hd__nand2_4
X_81486_ _81492_/CLK _81486_/D _81486_/Q sky130_fd_sc_hd__dfxtp_4
X_86013_ _85725_/CLK _51423_/Y _86013_/Q sky130_fd_sc_hd__dfxtp_4
X_52405_ _52400_/X _50708_/B _52405_/Y sky130_fd_sc_hd__nand2_4
X_83225_ _84350_/CLK _72591_/X _79343_/B sky130_fd_sc_hd__dfxtp_4
X_80437_ _80429_/B _80446_/B _80436_/X _80437_/Y sky130_fd_sc_hd__a21boi_4
X_68159_ _68461_/A _68160_/A sky130_fd_sc_hd__buf_2
X_56173_ _56167_/A _56173_/Y sky130_fd_sc_hd__inv_2
X_53385_ _53381_/Y _53382_/X _53384_/X _53385_/Y sky130_fd_sc_hd__a21oi_4
X_50597_ _50597_/A _48955_/X _50597_/Y sky130_fd_sc_hd__nand2_4
X_55124_ _73124_/B _73024_/B sky130_fd_sc_hd__buf_2
X_40350_ _40350_/A _42447_/D _41869_/C sky130_fd_sc_hd__nand2_4
X_52336_ _52320_/A _49031_/A _52336_/X sky130_fd_sc_hd__and2_4
X_71170_ _71170_/A _71181_/C sky130_fd_sc_hd__buf_2
X_83156_ _86213_/CLK _73317_/X _83156_/Q sky130_fd_sc_hd__dfxtp_4
X_80368_ _80358_/A _80357_/X _80367_/Y _80368_/Y sky130_fd_sc_hd__a21boi_4
X_70121_ _70121_/A _70125_/A sky130_fd_sc_hd__inv_2
X_82107_ _82349_/CLK _82107_/D _82107_/Q sky130_fd_sc_hd__dfxtp_4
X_55055_ _85327_/Q _55046_/X _55054_/Y _55055_/Y sky130_fd_sc_hd__o21ai_4
X_59932_ _59929_/C _59935_/A sky130_fd_sc_hd__inv_2
X_52267_ _48894_/A _52267_/B _52267_/C _52267_/X sky130_fd_sc_hd__and3_4
X_87964_ _87446_/CLK _42241_/Y _87964_/Q sky130_fd_sc_hd__dfxtp_4
X_83087_ _83187_/CLK _74352_/X _83087_/Q sky130_fd_sc_hd__dfxtp_4
X_80299_ _80296_/Y _80299_/B _80299_/Y sky130_fd_sc_hd__nand2_4
X_54006_ _53982_/A _54006_/X sky130_fd_sc_hd__buf_2
X_42020_ _88068_/Q _42020_/Y sky130_fd_sc_hd__inv_2
X_51218_ _50946_/A _51218_/X sky130_fd_sc_hd__buf_2
X_70052_ _68843_/X _68845_/X _69992_/X _70054_/A sky130_fd_sc_hd__a21o_4
X_86915_ _86914_/CLK _44861_/X _86915_/Q sky130_fd_sc_hd__dfxtp_4
X_82038_ _82008_/CLK _82038_/D _82038_/Q sky130_fd_sc_hd__dfxtp_4
X_59863_ _59842_/A _59873_/A sky130_fd_sc_hd__buf_2
X_52198_ _52198_/A _52198_/X sky130_fd_sc_hd__buf_2
X_87895_ _87382_/CLK _87895_/D _87895_/Q sky130_fd_sc_hd__dfxtp_4
X_58814_ _58813_/X _85774_/Q _58706_/X _58814_/X sky130_fd_sc_hd__o21a_4
X_51149_ _51149_/A _51160_/B sky130_fd_sc_hd__buf_2
X_74860_ _74850_/Y _74858_/Y _74859_/Y _74860_/Y sky130_fd_sc_hd__o21ai_4
X_86846_ _81117_/CLK _45902_/Y _42447_/C sky130_fd_sc_hd__dfxtp_4
X_59794_ _59794_/A _59794_/X sky130_fd_sc_hd__buf_2
X_73811_ _73786_/X _84983_/Q _73740_/X _73810_/X _73812_/B sky130_fd_sc_hd__a211o_4
X_58745_ _58742_/Y _58744_/Y _58646_/X _58745_/X sky130_fd_sc_hd__a21o_4
X_55957_ _55957_/A _56019_/B sky130_fd_sc_hd__buf_2
X_43971_ _43971_/A _43972_/B sky130_fd_sc_hd__inv_2
X_74791_ _70576_/X _83831_/Q _74764_/A _74791_/X sky130_fd_sc_hd__and3_4
X_86777_ _86814_/CLK _46080_/Y _86777_/Q sky130_fd_sc_hd__dfxtp_4
X_83989_ _81746_/CLK _68298_/X _83989_/Q sky130_fd_sc_hd__dfxtp_4
X_45710_ _85133_/Q _45709_/X _45651_/X _45710_/X sky130_fd_sc_hd__o21a_4
X_76530_ _81371_/Q _81627_/D _81339_/D sky130_fd_sc_hd__xor2_4
X_42922_ _42951_/A _42922_/X sky130_fd_sc_hd__buf_2
X_54908_ _85355_/Q _54892_/X _54907_/Y _54908_/Y sky130_fd_sc_hd__o21ai_4
X_85728_ _85727_/CLK _85728_/D _85728_/Q sky130_fd_sc_hd__dfxtp_4
X_73742_ _73742_/A _86554_/Q _73742_/X sky130_fd_sc_hd__and2_4
X_46690_ _46717_/A _46682_/B _46682_/C _51787_/D _46690_/X sky130_fd_sc_hd__and4_4
X_70954_ _70947_/A _70954_/B _70954_/C _70954_/Y sky130_fd_sc_hd__nand3_4
X_58676_ _58676_/A _58688_/B sky130_fd_sc_hd__buf_2
X_55888_ _55534_/A _55903_/A sky130_fd_sc_hd__buf_2
X_45641_ _45591_/X _61513_/A _45608_/X _45641_/Y sky130_fd_sc_hd__o21ai_4
X_57627_ _72009_/A _57627_/X sky130_fd_sc_hd__buf_2
X_76461_ _76454_/X _76457_/Y _76460_/X _76461_/X sky130_fd_sc_hd__o21a_4
X_42853_ _42832_/A _42853_/X sky130_fd_sc_hd__buf_2
X_54839_ _54892_/A _54839_/X sky130_fd_sc_hd__buf_2
X_73673_ _70125_/C _86754_/D _73672_/X _73673_/Y sky130_fd_sc_hd__o21ai_4
X_85659_ _85433_/CLK _53304_/Y _85659_/Q sky130_fd_sc_hd__dfxtp_4
X_70885_ _70885_/A _70885_/X sky130_fd_sc_hd__buf_2
X_78200_ _78205_/A _78204_/A _78199_/Y _78200_/Y sky130_fd_sc_hd__a21boi_4
X_75412_ _75411_/Y _75413_/C sky130_fd_sc_hd__inv_2
X_41804_ _41802_/X _41803_/X _40371_/X _66621_/B _41792_/X _41805_/A
+ sky130_fd_sc_hd__o32ai_4
X_48360_ _86529_/Q _48350_/X _48359_/Y _48360_/Y sky130_fd_sc_hd__o21ai_4
X_72624_ _79183_/A _61349_/X _72577_/Y _83212_/D sky130_fd_sc_hd__o21ai_4
X_79180_ _79180_/A _66514_/C _79180_/Y sky130_fd_sc_hd__nand2_4
X_45572_ _45572_/A _45617_/B _45572_/Y sky130_fd_sc_hd__nor2_4
X_57558_ _57552_/X _47978_/A _57558_/Y sky130_fd_sc_hd__nand2_4
X_88378_ _87865_/CLK _40521_/X _88378_/Q sky130_fd_sc_hd__dfxtp_4
X_76392_ _76393_/A _81567_/Q _76392_/Y sky130_fd_sc_hd__nor2_4
X_42784_ _42774_/X _42775_/X _41347_/X _87720_/Q _42781_/X _42785_/A
+ sky130_fd_sc_hd__o32ai_4
X_47311_ _47330_/A _47311_/B _47321_/C _52977_/D _47311_/X sky130_fd_sc_hd__and4_4
X_78131_ _78105_/Y _78131_/B _78131_/Y sky130_fd_sc_hd__nand2_4
X_44523_ _44512_/X _44513_/X _40780_/Y _44522_/Y _44516_/X _87068_/D
+ sky130_fd_sc_hd__o32ai_4
X_56509_ _56448_/X _56520_/B sky130_fd_sc_hd__buf_2
X_75343_ _75326_/X _75322_/X _75323_/X _75343_/Y sky130_fd_sc_hd__a21oi_4
X_87329_ _87850_/CLK _87329_/D _87329_/Q sky130_fd_sc_hd__dfxtp_4
X_41735_ _41734_/X _41735_/X sky130_fd_sc_hd__buf_2
X_48291_ _52039_/A _48286_/X _48287_/C _48291_/X sky130_fd_sc_hd__and3_4
X_72555_ _72516_/C _72555_/B _72563_/C _72607_/C _72572_/A sky130_fd_sc_hd__nand4_4
X_57489_ _47819_/A _57489_/B _57489_/Y sky130_fd_sc_hd__nand2_4
X_47242_ _47242_/A _54102_/B sky130_fd_sc_hd__inv_2
X_59228_ _59216_/Y _59145_/X _59223_/X _59227_/X _84759_/D sky130_fd_sc_hd__a22oi_4
X_71506_ _70886_/A _71735_/C _71263_/D _70500_/B _71507_/B sky130_fd_sc_hd__nand4_4
X_78062_ _60789_/C _78062_/B _78062_/X sky130_fd_sc_hd__xor2_4
X_44454_ _44454_/A _44454_/X sky130_fd_sc_hd__buf_2
X_75274_ _75274_/A _75274_/Y sky130_fd_sc_hd__inv_2
X_41666_ _41628_/X _81754_/Q _41665_/X _41666_/X sky130_fd_sc_hd__o21a_4
X_72486_ _63562_/A _72488_/B _72486_/Y sky130_fd_sc_hd__nand2_4
X_77013_ _77013_/A _77013_/B _77013_/Y sky130_fd_sc_hd__nand2_4
X_43405_ _43399_/X _43404_/X _41493_/X _87437_/Q _43378_/X _43405_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74225_ _41973_/Y _73930_/X _73031_/X _74224_/Y _74225_/X sky130_fd_sc_hd__a211o_4
X_40617_ _40616_/Y _40617_/X sky130_fd_sc_hd__buf_2
X_47173_ _83694_/Q _54587_/B sky130_fd_sc_hd__inv_2
X_71437_ _71432_/A _71435_/B _70790_/A _71432_/D _71437_/X sky130_fd_sc_hd__and4_4
X_59159_ _59159_/A _59159_/Y sky130_fd_sc_hd__inv_2
X_44385_ _44385_/A _44385_/Y sky130_fd_sc_hd__inv_2
X_41597_ _41540_/X _41541_/X _41596_/X _88185_/Q _41537_/X _41597_/Y
+ sky130_fd_sc_hd__o32ai_4
X_46124_ _46124_/A _46125_/A sky130_fd_sc_hd__inv_2
X_43336_ _43287_/A _43336_/X sky130_fd_sc_hd__buf_2
X_62170_ _59730_/A _62170_/B _62158_/C _63342_/B _62170_/X sky130_fd_sc_hd__and4_4
X_74156_ _73165_/A _74237_/A sky130_fd_sc_hd__buf_2
X_40548_ _40547_/Y _40548_/X sky130_fd_sc_hd__buf_2
X_71368_ _71090_/A _71439_/C sky130_fd_sc_hd__buf_2
Xclkbuf_10_282_0_CLK clkbuf_9_141_0_CLK/X _83372_/CLK sky130_fd_sc_hd__clkbuf_1
X_61121_ _61120_/Y _64203_/B sky130_fd_sc_hd__buf_2
X_73107_ _69734_/Y _73195_/A _72889_/X _73106_/Y _73107_/X sky130_fd_sc_hd__a211o_4
X_46055_ _46046_/X _46054_/X _41535_/X _86791_/Q _46047_/X _46055_/Y
+ sky130_fd_sc_hd__o32ai_4
X_70319_ _70317_/Y _70157_/A _70318_/Y _70319_/Y sky130_fd_sc_hd__o21ai_4
X_43267_ _41104_/X _43264_/X _87509_/Q _43265_/X _87509_/D sky130_fd_sc_hd__a2bb2o_4
X_74087_ _72880_/A _74087_/X sky130_fd_sc_hd__buf_2
X_78964_ _78970_/B _78964_/B _78965_/B sky130_fd_sc_hd__xnor2_4
X_40479_ _40456_/X _81167_/Q _40478_/X _40479_/X sky130_fd_sc_hd__o21a_4
X_71299_ _48016_/B _71290_/X _71298_/Y _83544_/D sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_64_0_CLK clkbuf_9_32_0_CLK/X _80671_/CLK sky130_fd_sc_hd__clkbuf_1
X_45006_ _83035_/Q _45007_/A sky130_fd_sc_hd__inv_2
X_42218_ _41352_/X _42209_/X _87975_/Q _42210_/X _87975_/D sky130_fd_sc_hd__a2bb2o_4
X_77915_ _77910_/Y _77902_/B _77914_/Y _77916_/B sky130_fd_sc_hd__o21ai_4
X_61052_ _60715_/X _61138_/B sky130_fd_sc_hd__buf_2
X_73038_ _73034_/X _73037_/X _72737_/A _73038_/X sky130_fd_sc_hd__a21o_4
X_43198_ _43197_/Y _43198_/Y sky130_fd_sc_hd__inv_2
X_78895_ _78885_/B _82507_/D sky130_fd_sc_hd__inv_2
Xclkbuf_8_210_0_CLK clkbuf_8_211_0_CLK/A clkbuf_8_210_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_60003_ _59913_/X _60091_/B _60091_/C _60003_/Y sky130_fd_sc_hd__nand3_4
X_49814_ _57991_/B _49798_/X _49813_/Y _49814_/Y sky130_fd_sc_hd__o21ai_4
X_42149_ _41911_/A _42162_/A sky130_fd_sc_hd__buf_2
X_65860_ _65718_/A _65860_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_109_0_CLK clkbuf_6_54_0_CLK/X clkbuf_8_219_0_CLK/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_297_0_CLK clkbuf_9_148_0_CLK/X _84358_/CLK sky130_fd_sc_hd__clkbuf_1
X_77846_ _77844_/Y _77845_/Y _77849_/A sky130_fd_sc_hd__xor2_4
X_64811_ _64809_/X _83306_/Q _64733_/X _64810_/X _64811_/X sky130_fd_sc_hd__a211o_4
X_49745_ _57820_/B _49742_/X _49744_/Y _49745_/Y sky130_fd_sc_hd__o21ai_4
X_46957_ _83717_/Q _54464_/B sky130_fd_sc_hd__inv_2
X_65791_ _65791_/A _65804_/A sky130_fd_sc_hd__buf_2
X_77777_ _77763_/Y _77766_/Y _77777_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_79_0_CLK clkbuf_9_39_0_CLK/X _84420_/CLK sky130_fd_sc_hd__clkbuf_1
X_74989_ _74987_/B _81140_/D _74989_/C _74990_/A sky130_fd_sc_hd__nand3_4
X_79516_ _79503_/A _79503_/B _79515_/Y _79517_/B sky130_fd_sc_hd__a21boi_4
X_67530_ _67575_/A _88235_/Q _67530_/X sky130_fd_sc_hd__and2_4
X_45908_ _44039_/X _45909_/A sky130_fd_sc_hd__buf_2
X_64742_ _64737_/Y _64662_/X _64741_/Y _84229_/D sky130_fd_sc_hd__a21o_4
X_76728_ _76728_/A _76728_/B _76728_/Y sky130_fd_sc_hd__xnor2_4
X_49676_ _86343_/Q _49660_/X _49675_/Y _49676_/Y sky130_fd_sc_hd__o21ai_4
X_61954_ _58335_/A _61954_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_225_0_CLK clkbuf_8_225_0_CLK/A clkbuf_9_451_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_46888_ _46860_/X _51043_/B _46888_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_220_0_CLK clkbuf_9_110_0_CLK/X _84241_/CLK sky130_fd_sc_hd__clkbuf_1
X_48627_ _48627_/A _48628_/B sky130_fd_sc_hd__buf_2
X_60905_ _60997_/A _64081_/C _60889_/X _60864_/X _69814_/A _60905_/Y
+ sky130_fd_sc_hd__a41oi_4
X_67461_ _87918_/Q _67414_/X _67391_/X _67460_/X _67461_/X sky130_fd_sc_hd__a211o_4
X_79447_ _79447_/A _79447_/B _79453_/B sky130_fd_sc_hd__xor2_4
Xclkbuf_10_850_0_CLK clkbuf_9_425_0_CLK/X _85953_/CLK sky130_fd_sc_hd__clkbuf_1
X_45839_ _84996_/Q _55231_/B sky130_fd_sc_hd__inv_2
X_64673_ _64773_/A _86430_/Q _64673_/X sky130_fd_sc_hd__and2_4
X_76659_ _76659_/A _76662_/C sky130_fd_sc_hd__inv_2
X_61885_ _61915_/A _61915_/B _58511_/A _61915_/D _61885_/X sky130_fd_sc_hd__and4_4
X_69200_ _69146_/X _69198_/Y _69095_/X _69199_/Y _69200_/X sky130_fd_sc_hd__a211o_4
X_66412_ _64862_/X _66417_/B _64866_/X _66412_/Y sky130_fd_sc_hd__nand3_4
X_63624_ _63358_/X _63624_/X sky130_fd_sc_hd__buf_2
X_48558_ _48553_/Y _48403_/X _48557_/Y _86512_/D sky130_fd_sc_hd__a21boi_4
X_60836_ _60610_/A _60835_/X _84555_/Q _60836_/X sky130_fd_sc_hd__or3_4
X_67392_ _67342_/A _67392_/B _67392_/X sky130_fd_sc_hd__and2_4
X_79378_ _79364_/Y _79361_/X _79378_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_341_0_CLK clkbuf_9_341_0_CLK/A clkbuf_9_341_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_69131_ _69127_/X _69130_/X _69017_/X _69131_/Y sky130_fd_sc_hd__a21oi_4
X_47509_ _47414_/A _47509_/X sky130_fd_sc_hd__buf_2
X_66343_ _66065_/A _66343_/X sky130_fd_sc_hd__buf_2
X_78329_ _78329_/A _78329_/Y sky130_fd_sc_hd__inv_2
X_63555_ _63553_/Y _63516_/X _63554_/Y _63555_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_235_0_CLK clkbuf_9_117_0_CLK/X _80681_/CLK sky130_fd_sc_hd__clkbuf_1
X_48489_ _52156_/A _48489_/B _48533_/C _48489_/X sky130_fd_sc_hd__and3_4
X_60767_ _60766_/X _60767_/X sky130_fd_sc_hd__buf_2
X_50520_ _50518_/Y _50491_/X _50519_/X _50520_/Y sky130_fd_sc_hd__a21oi_4
X_62506_ _62493_/A _62506_/B _62506_/C _62506_/D _62506_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_10_865_0_CLK clkbuf_9_432_0_CLK/X _83556_/CLK sky130_fd_sc_hd__clkbuf_1
X_81340_ _84049_/CLK _81340_/D _81716_/D sky130_fd_sc_hd__dfxtp_4
X_69062_ _69057_/X _69060_/X _69061_/X _69062_/Y sky130_fd_sc_hd__a21oi_4
X_66274_ _66225_/X _84968_/Q _66186_/X _66273_/X _66274_/X sky130_fd_sc_hd__a211o_4
X_63486_ _58543_/Y _63436_/X _61451_/A _63437_/X _63486_/X sky130_fd_sc_hd__a2bb2o_4
X_60698_ _60697_/Y _60646_/Y _59756_/A _60698_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_10_17_0_CLK clkbuf_9_8_0_CLK/X _85198_/CLK sky130_fd_sc_hd__clkbuf_1
X_68013_ _68371_/A _88151_/Q _68013_/X sky130_fd_sc_hd__and2_4
X_65225_ _65225_/A _65225_/B _65225_/X sky130_fd_sc_hd__and2_4
X_50451_ _52156_/A _50456_/B _50462_/C _50451_/X sky130_fd_sc_hd__and3_4
Xclkbuf_9_356_0_CLK clkbuf_8_178_0_CLK/X clkbuf_9_356_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_62437_ _62276_/X _62479_/C sky130_fd_sc_hd__buf_2
X_81271_ _81257_/CLK _81303_/Q _81271_/Q sky130_fd_sc_hd__dfxtp_4
X_83010_ _82979_/CLK _74626_/Y _45380_/A sky130_fd_sc_hd__dfxtp_4
X_80222_ _80184_/Y _80187_/Y _80199_/X _80197_/Y _80220_/B _80222_/X
+ sky130_fd_sc_hd__a2111o_4
X_53170_ _53181_/A _53159_/B _53169_/X _53170_/D _53170_/X sky130_fd_sc_hd__and4_4
X_65156_ _64999_/X _86156_/Q _65127_/X _65155_/X _65156_/X sky130_fd_sc_hd__a211o_4
X_50382_ _50379_/Y _50380_/X _50381_/Y _50382_/Y sky130_fd_sc_hd__a21boi_4
X_62368_ _62356_/X _62362_/Y _62366_/X _84743_/Q _62367_/X _62368_/Y
+ sky130_fd_sc_hd__o32ai_4
X_52121_ _52121_/A _52121_/B _52121_/Y sky130_fd_sc_hd__nand2_4
X_64107_ _64077_/Y _64102_/Y _64103_/X _64105_/X _64106_/X _64107_/Y
+ sky130_fd_sc_hd__o41ai_4
X_61319_ _61281_/A _61319_/X sky130_fd_sc_hd__buf_2
X_80153_ _80153_/A _63897_/C _80153_/X sky130_fd_sc_hd__xor2_4
X_65087_ _65005_/X _65087_/B _65087_/X sky130_fd_sc_hd__and2_4
X_69964_ _69546_/X _69548_/X _69939_/X _69964_/Y sky130_fd_sc_hd__a21oi_4
X_62299_ _62634_/A _62293_/Y _62299_/C _62298_/Y _62299_/Y sky130_fd_sc_hd__nand4_4
X_52052_ _52070_/A _48073_/B _52052_/Y sky130_fd_sc_hd__nand2_4
X_64038_ _64036_/X _63994_/X _64037_/Y _84279_/D sky130_fd_sc_hd__a21oi_4
X_68915_ _68912_/X _68914_/X _68846_/X _68915_/Y sky130_fd_sc_hd__a21oi_4
X_84961_ _84960_/CLK _84961_/D _84961_/Q sky130_fd_sc_hd__dfxtp_4
X_80084_ _80080_/Y _80083_/Y _80084_/X sky130_fd_sc_hd__xor2_4
X_69895_ _69086_/A _87290_/Q _69895_/X sky130_fd_sc_hd__and2_4
X_51003_ _51003_/A _51003_/B _51003_/Y sky130_fd_sc_hd__nand2_4
X_86700_ _86701_/CLK _86700_/D _86700_/Q sky130_fd_sc_hd__dfxtp_4
X_83912_ _81975_/CLK _69591_/X _83912_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_803_0_CLK clkbuf_9_401_0_CLK/X _82860_/CLK sky130_fd_sc_hd__clkbuf_1
X_56860_ _56859_/X _56860_/X sky130_fd_sc_hd__buf_2
X_68846_ _60109_/A _68846_/X sky130_fd_sc_hd__buf_2
X_87680_ _82888_/CLK _42863_/X _67033_/B sky130_fd_sc_hd__dfxtp_4
X_84892_ _84892_/CLK _84892_/D _84892_/Q sky130_fd_sc_hd__dfxtp_4
X_55811_ _55811_/A _55811_/X sky130_fd_sc_hd__buf_2
X_86631_ _85990_/CLK _86631_/D _86631_/Q sky130_fd_sc_hd__dfxtp_4
X_83843_ _83843_/CLK _70191_/X _83843_/Q sky130_fd_sc_hd__dfxtp_4
X_56791_ _56786_/Y _57673_/A _56790_/X _56791_/Y sky130_fd_sc_hd__nand3_4
X_68777_ _68774_/X _68776_/X _68777_/Y sky130_fd_sc_hd__nand2_4
X_65989_ _65986_/Y _65987_/X _65988_/X _65989_/X sky130_fd_sc_hd__a21o_4
X_58530_ _58530_/A _58530_/Y sky130_fd_sc_hd__inv_2
X_55742_ _45380_/A _55152_/X _55140_/A _55741_/X _55742_/X sky130_fd_sc_hd__a211o_4
X_67728_ _87971_/Q _67651_/X _67625_/X _67727_/X _67728_/X sky130_fd_sc_hd__a211o_4
X_86562_ _86490_/CLK _86562_/D _86562_/Q sky130_fd_sc_hd__dfxtp_4
X_52954_ _52947_/X _52954_/B _52977_/C _52954_/D _52954_/X sky130_fd_sc_hd__and4_4
X_83774_ _86553_/CLK _83774_/D _83774_/Q sky130_fd_sc_hd__dfxtp_4
X_80986_ _80818_/CLK _80986_/D _80986_/Q sky130_fd_sc_hd__dfxtp_4
X_88301_ _88301_/CLK _40969_/X _69224_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_818_0_CLK clkbuf_9_409_0_CLK/X _82924_/CLK sky130_fd_sc_hd__clkbuf_1
X_85513_ _85514_/CLK _54062_/Y _85513_/Q sky130_fd_sc_hd__dfxtp_4
X_51905_ _51887_/A _51898_/B _51893_/C _52730_/D _51905_/X sky130_fd_sc_hd__and4_4
X_58461_ _58461_/A _58498_/B _58461_/Y sky130_fd_sc_hd__nand2_4
X_82725_ _82923_/CLK _66509_/C _78838_/A sky130_fd_sc_hd__dfxtp_4
X_67659_ _67658_/X _67659_/B _67659_/X sky130_fd_sc_hd__and2_4
X_55673_ _55288_/B _55288_/A _55672_/X _55674_/A sky130_fd_sc_hd__nand3_4
X_86493_ _85596_/CLK _86493_/D _65489_/B sky130_fd_sc_hd__dfxtp_4
X_52885_ _52885_/A _52885_/B _52885_/Y sky130_fd_sc_hd__nand2_4
X_57412_ _57408_/X _57410_/Y _57411_/Y _57412_/X sky130_fd_sc_hd__o21a_4
X_88232_ _88232_/CLK _88232_/D _67600_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_309_0_CLK clkbuf_8_154_0_CLK/X clkbuf_9_309_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_54624_ _85408_/Q _54621_/X _54623_/Y _54624_/Y sky130_fd_sc_hd__o21ai_4
X_85444_ _85444_/CLK _85444_/D _85444_/Q sky130_fd_sc_hd__dfxtp_4
X_51836_ _85937_/Q _51817_/X _51835_/Y _51836_/Y sky130_fd_sc_hd__o21ai_4
X_70670_ _70670_/A _70676_/B _70676_/C _70670_/Y sky130_fd_sc_hd__nor3_4
X_58392_ _58388_/X _83349_/Q _58391_/Y _84861_/D sky130_fd_sc_hd__o21a_4
X_82656_ _81783_/CLK _84008_/Q _79086_/A sky130_fd_sc_hd__dfxtp_4
X_57343_ _44287_/X _57339_/X _57340_/Y _57342_/Y _57344_/A sky130_fd_sc_hd__a211o_4
X_81607_ _85003_/CLK _81607_/D _81607_/Q sky130_fd_sc_hd__dfxtp_4
X_69329_ _68300_/X _69329_/X sky130_fd_sc_hd__buf_2
X_88163_ _87150_/CLK _41716_/X _67724_/B sky130_fd_sc_hd__dfxtp_4
X_54555_ _54546_/A _47116_/A _54555_/Y sky130_fd_sc_hd__nand2_4
X_85375_ _85375_/CLK _85375_/D _85375_/Q sky130_fd_sc_hd__dfxtp_4
X_51767_ _51793_/A _51767_/X sky130_fd_sc_hd__buf_2
X_82587_ _82675_/CLK _82619_/Q _78265_/A sky130_fd_sc_hd__dfxtp_4
X_87114_ _87116_/CLK _87114_/D _87114_/Q sky130_fd_sc_hd__dfxtp_4
X_53506_ _53448_/X _53506_/X sky130_fd_sc_hd__buf_2
X_41520_ _41519_/X _41520_/X sky130_fd_sc_hd__buf_2
X_72340_ _72339_/X _85327_/Q _72255_/X _72340_/X sky130_fd_sc_hd__o21a_4
X_84326_ _84355_/CLK _63408_/Y _80588_/B sky130_fd_sc_hd__dfxtp_4
X_50718_ _50718_/A _50740_/A sky130_fd_sc_hd__buf_2
X_81538_ _81346_/CLK _81538_/D _81526_/D sky130_fd_sc_hd__dfxtp_4
X_57274_ _57273_/Y _56672_/Y _57274_/Y sky130_fd_sc_hd__nand2_4
X_88094_ _88108_/CLK _41955_/Y _74051_/A sky130_fd_sc_hd__dfxtp_4
X_54486_ _54486_/A _54486_/X sky130_fd_sc_hd__buf_2
X_51698_ _85962_/Q _51675_/X _51697_/Y _51698_/Y sky130_fd_sc_hd__o21ai_4
X_59013_ _58904_/A _59013_/X sky130_fd_sc_hd__buf_2
X_56225_ _56255_/A _56225_/X sky130_fd_sc_hd__buf_2
X_41451_ _41482_/A _41459_/B sky130_fd_sc_hd__buf_2
X_87045_ _87045_/CLK _87045_/D _44583_/A sky130_fd_sc_hd__dfxtp_4
X_53437_ _53436_/X _53437_/X sky130_fd_sc_hd__buf_2
X_72271_ _59238_/A _72366_/A sky130_fd_sc_hd__buf_2
X_84257_ _84314_/CLK _64313_/X _79797_/B sky130_fd_sc_hd__dfxtp_4
X_50649_ _50607_/A _50649_/B _50649_/Y sky130_fd_sc_hd__nand2_4
X_81469_ _82648_/CLK _76902_/Y _81469_/Q sky130_fd_sc_hd__dfxtp_4
X_74010_ _88352_/Q _73801_/X _73087_/X _74010_/Y sky130_fd_sc_hd__o21ai_4
X_40402_ _40402_/A _40402_/B _40402_/X sky130_fd_sc_hd__or2_4
X_71222_ _71054_/A _71223_/B sky130_fd_sc_hd__buf_2
X_83208_ _83843_/CLK _83208_/D _70176_/C sky130_fd_sc_hd__dfxtp_4
X_44170_ _44170_/A _65768_/A sky130_fd_sc_hd__buf_2
X_56156_ _55745_/D _56167_/A sky130_fd_sc_hd__buf_2
X_53368_ _53365_/Y _53355_/X _53367_/X _53368_/Y sky130_fd_sc_hd__a21oi_4
X_41382_ _41381_/X _41382_/X sky130_fd_sc_hd__buf_2
X_84188_ _83521_/CLK _84188_/D _84188_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_5_9_0_CLK clkbuf_4_4_1_CLK/X clkbuf_5_9_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_55107_ _85317_/Q _55098_/X _55106_/Y _55107_/Y sky130_fd_sc_hd__o21ai_4
X_43121_ _43121_/A _43121_/X sky130_fd_sc_hd__buf_2
X_40333_ _43012_/B _40332_/Y _40343_/A sky130_fd_sc_hd__nor2_4
X_52319_ _52319_/A _52320_/A sky130_fd_sc_hd__buf_2
X_71153_ _48401_/B _71138_/X _71152_/Y _71153_/Y sky130_fd_sc_hd__o21ai_4
X_83139_ _83139_/CLK _73722_/Y _70103_/A sky130_fd_sc_hd__dfxtp_4
X_56087_ _56082_/X _56085_/X _56086_/Y _56087_/Y sky130_fd_sc_hd__o21ai_4
X_53299_ _85659_/Q _53295_/X _53298_/Y _53299_/Y sky130_fd_sc_hd__o21ai_4
X_70104_ _83138_/Q _70107_/B sky130_fd_sc_hd__inv_2
X_43052_ _43052_/A _87594_/D sky130_fd_sc_hd__inv_2
X_55038_ _85330_/Q _55020_/X _55037_/Y _55038_/Y sky130_fd_sc_hd__o21ai_4
X_59915_ _59657_/A _61293_/B _59753_/B _60407_/C _59917_/A sky130_fd_sc_hd__and4_4
X_71084_ _71071_/A _71088_/A sky130_fd_sc_hd__buf_2
X_75961_ _75961_/A _75961_/Y sky130_fd_sc_hd__inv_2
X_87947_ _87950_/CLK _87947_/D _87947_/Q sky130_fd_sc_hd__dfxtp_4
X_42003_ _41998_/X _41993_/X _40806_/X _42002_/Y _42000_/X _42003_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77700_ _77698_/Y _77699_/X _77700_/X sky130_fd_sc_hd__xor2_4
X_74912_ _81132_/D _74912_/B _74912_/X sky130_fd_sc_hd__xor2_4
X_70035_ _69520_/X _69758_/Y _70033_/X _70034_/Y _70035_/X sky130_fd_sc_hd__a211o_4
X_47860_ _46578_/X _46274_/A _47859_/X _47861_/B sky130_fd_sc_hd__o21ai_4
X_59846_ _60781_/A _59846_/X sky130_fd_sc_hd__buf_2
X_78680_ _78680_/A _78680_/B _78680_/Y sky130_fd_sc_hd__nand2_4
X_75892_ _84490_/Q _62995_/C _75892_/X sky130_fd_sc_hd__xor2_4
X_87878_ _88398_/CLK _42407_/Y _87878_/Q sky130_fd_sc_hd__dfxtp_4
X_46811_ _46784_/A _46830_/B _46830_/C _46810_/X _46811_/X sky130_fd_sc_hd__and4_4
X_77631_ _77630_/A _82109_/D _77632_/A sky130_fd_sc_hd__nand2_4
X_86829_ _87990_/CLK _86829_/D _86829_/Q sky130_fd_sc_hd__dfxtp_4
X_74843_ _45909_/X _46167_/B _46167_/A _74843_/Y sky130_fd_sc_hd__nor3_4
X_47791_ _47745_/A _47791_/X sky130_fd_sc_hd__buf_2
X_59777_ _72176_/A _59837_/B sky130_fd_sc_hd__buf_2
X_56989_ _56989_/A _56989_/B _56989_/Y sky130_fd_sc_hd__nand2_4
X_49530_ _49546_/A _46912_/X _49530_/Y sky130_fd_sc_hd__nand2_4
X_46742_ _58727_/A _46719_/X _46741_/Y _46742_/Y sky130_fd_sc_hd__o21ai_4
X_58728_ _58603_/A _58728_/X sky130_fd_sc_hd__buf_2
X_77562_ _77561_/A _77561_/C _77542_/A _77562_/Y sky130_fd_sc_hd__a21oi_4
X_43954_ _43979_/A _43954_/X sky130_fd_sc_hd__buf_2
X_74774_ _70586_/X _83829_/Q _74753_/X _74774_/X sky130_fd_sc_hd__and3_4
X_71986_ _72017_/A _72007_/A sky130_fd_sc_hd__buf_2
X_79301_ _79301_/A _83221_/Q _79301_/X sky130_fd_sc_hd__xor2_4
X_76513_ _76478_/X _76513_/B _76513_/C _76513_/D _76514_/A sky130_fd_sc_hd__and4_4
X_42905_ _42835_/X _42905_/X sky130_fd_sc_hd__buf_2
X_49461_ _49407_/A _49467_/A sky130_fd_sc_hd__buf_2
X_73725_ _87340_/Q _73701_/B _73725_/Y sky130_fd_sc_hd__nor2_4
X_70937_ _70936_/X _70937_/X sky130_fd_sc_hd__buf_2
X_46673_ _46249_/A _46720_/A sky130_fd_sc_hd__buf_2
X_58659_ _58659_/A _86394_/Q _58659_/Y sky130_fd_sc_hd__nor2_4
X_77493_ _77493_/A _77493_/Y sky130_fd_sc_hd__inv_2
X_43885_ _41302_/X _43879_/X _87216_/Q _43880_/X _87216_/D sky130_fd_sc_hd__a2bb2o_4
X_48412_ _48401_/A _52121_/B _48412_/Y sky130_fd_sc_hd__nand2_4
X_79232_ _79230_/Y _79232_/B _79233_/A sky130_fd_sc_hd__or2_4
Xclkbuf_7_71_0_CLK clkbuf_7_70_0_CLK/A clkbuf_7_71_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_45624_ _45591_/X _61502_/A _45608_/X _45624_/Y sky130_fd_sc_hd__o21ai_4
X_76444_ _76432_/X _76444_/Y sky130_fd_sc_hd__inv_2
X_42836_ _42835_/X _42836_/X sky130_fd_sc_hd__buf_2
X_49392_ _49397_/A _49369_/X _49408_/C _51777_/D _49392_/X sky130_fd_sc_hd__and4_4
X_61670_ _61663_/Y _61665_/Y _61594_/X _61666_/Y _61669_/Y _61670_/X
+ sky130_fd_sc_hd__a41o_4
X_73656_ _72861_/X _73656_/X sky130_fd_sc_hd__buf_2
X_70868_ _51800_/B _70855_/X _70867_/Y _70868_/Y sky130_fd_sc_hd__o21ai_4
X_48343_ _48348_/A _50381_/B _48343_/Y sky130_fd_sc_hd__nand2_4
X_60621_ _60620_/Y _60622_/D sky130_fd_sc_hd__inv_2
X_72607_ _72516_/A _72607_/B _72607_/C _72607_/Y sky130_fd_sc_hd__nand3_4
X_79163_ _84786_/Q _66524_/C _79163_/Y sky130_fd_sc_hd__nand2_4
X_45555_ _45550_/X _45554_/X _45523_/X _45555_/X sky130_fd_sc_hd__a21o_4
X_76375_ _81361_/Q _81617_/D _76375_/X sky130_fd_sc_hd__xor2_4
X_42767_ _42745_/A _42767_/X sky130_fd_sc_hd__buf_2
X_73587_ _73584_/X _73586_/X _73383_/X _73590_/A sky130_fd_sc_hd__a21o_4
X_70799_ _70798_/X _71221_/A sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_1_CLK clkbuf_1_1_0_CLK/X clkbuf_1_1_1_CLK/X sky130_fd_sc_hd__clkbuf_1
X_78114_ _82567_/Q _78108_/B _78114_/Y sky130_fd_sc_hd__nand2_4
X_44506_ _41267_/Y _44502_/X _87075_/Q _44503_/X _44506_/X sky130_fd_sc_hd__a2bb2o_4
X_75326_ _75289_/Y _75291_/X _75301_/X _75326_/X sky130_fd_sc_hd__a21o_4
X_63340_ _60454_/A _64545_/B _60441_/B _60473_/B _63340_/X sky130_fd_sc_hd__and4_4
X_41718_ _46317_/A _41718_/X sky130_fd_sc_hd__buf_2
X_48274_ _48903_/A _49215_/A sky130_fd_sc_hd__buf_2
X_72538_ _61278_/B _61281_/C _63733_/X _61260_/A _61319_/X _72539_/B
+ sky130_fd_sc_hd__a32oi_4
X_60552_ _72527_/A _72527_/B _79141_/A _60551_/X _60595_/C _84601_/D
+ sky130_fd_sc_hd__a32o_4
X_79094_ _79095_/A _79095_/B _79094_/X sky130_fd_sc_hd__xor2_4
X_45486_ _85115_/Q _45456_/X _45486_/Y sky130_fd_sc_hd__nor2_4
X_42698_ _41108_/X _42695_/X _69553_/B _42696_/X _42698_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_7_86_0_CLK clkbuf_7_87_0_CLK/A clkbuf_7_86_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_47225_ _47130_/A _47228_/B sky130_fd_sc_hd__buf_2
X_78045_ _78045_/A _78045_/B _81923_/D sky130_fd_sc_hd__nand2_4
X_44437_ _44437_/A _44437_/Y sky130_fd_sc_hd__inv_2
X_63271_ _58498_/A _63250_/X _58400_/A _60493_/X _63271_/X sky130_fd_sc_hd__o22a_4
X_75257_ _75256_/Y _75258_/C sky130_fd_sc_hd__inv_2
X_41649_ _82909_/Q _41624_/B _41649_/X sky130_fd_sc_hd__or2_4
X_60483_ _60482_/Y _60484_/A sky130_fd_sc_hd__buf_2
X_72469_ _57791_/X _85955_/Q _72468_/X _72469_/Y sky130_fd_sc_hd__o21ai_4
X_65010_ _64904_/A _85842_/Q _65010_/X sky130_fd_sc_hd__and2_4
X_62222_ _62336_/A _62236_/A sky130_fd_sc_hd__buf_2
X_74208_ _74205_/X _74207_/X _73602_/X _74208_/X sky130_fd_sc_hd__a21o_4
X_47156_ _47151_/Y _47128_/X _47155_/X _47156_/Y sky130_fd_sc_hd__a21oi_4
X_44368_ _41749_/X _44364_/X _87144_/Q _44365_/X _87144_/D sky130_fd_sc_hd__a2bb2o_4
X_75188_ _75188_/A _75190_/B sky130_fd_sc_hd__inv_2
X_46107_ _46107_/A _46188_/A _46108_/D sky130_fd_sc_hd__nor2_4
X_43319_ _43305_/A _43319_/X sky130_fd_sc_hd__buf_2
X_62153_ _61715_/A _62153_/B _62150_/Y _62152_/Y _62153_/Y sky130_fd_sc_hd__nand4_4
X_74139_ _74139_/A _74139_/X sky130_fd_sc_hd__buf_2
X_47087_ _47087_/A _53364_/B sky130_fd_sc_hd__inv_2
X_44299_ _44299_/A _59238_/A sky130_fd_sc_hd__buf_2
X_79996_ _79995_/Y _80000_/A sky130_fd_sc_hd__inv_2
X_61104_ _61095_/X _61097_/X _61230_/C _61103_/X _60529_/A _61104_/Y
+ sky130_fd_sc_hd__a41oi_4
X_46038_ _46038_/A _46038_/Y sky130_fd_sc_hd__inv_2
X_66961_ _68721_/A _66961_/X sky130_fd_sc_hd__buf_2
X_62084_ _61716_/X _61607_/B _62083_/X _62084_/X sky130_fd_sc_hd__a21o_4
X_78947_ _82737_/Q _78947_/B _82705_/D sky130_fd_sc_hd__xor2_4
X_68700_ _86994_/Q _68570_/X _68571_/X _68699_/X _68700_/X sky130_fd_sc_hd__a211o_4
X_65912_ _65811_/X _84993_/Q _65865_/X _65911_/X _65912_/X sky130_fd_sc_hd__a211o_4
X_61035_ _60998_/X _60996_/Y _60880_/X _61035_/X sky130_fd_sc_hd__a21bo_4
X_69680_ _69680_/A _88331_/Q _69680_/X sky130_fd_sc_hd__and2_4
X_66892_ _66823_/A _66892_/B _66892_/X sky130_fd_sc_hd__and2_4
X_78878_ _78876_/X _78865_/X _78877_/X _78878_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_7_24_0_CLK clkbuf_6_12_0_CLK/X clkbuf_8_49_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_68631_ _68560_/A _68631_/B _68631_/X sky130_fd_sc_hd__and2_4
X_65843_ _65833_/Y _65841_/Y _65842_/X _65843_/Y sky130_fd_sc_hd__a21oi_4
X_77829_ _77822_/Y _77835_/A _77828_/Y _77830_/B sky130_fd_sc_hd__a21oi_4
X_47989_ _73927_/B _47948_/X _47988_/Y _47989_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_8_164_0_CLK clkbuf_7_82_0_CLK/X clkbuf_9_329_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_49728_ _49708_/A _49724_/B _49724_/C _52942_/D _49728_/X sky130_fd_sc_hd__and4_4
X_80840_ _80746_/CLK _80872_/Q _80840_/Q sky130_fd_sc_hd__dfxtp_4
X_68562_ _68559_/X _68561_/X _68327_/X _68562_/Y sky130_fd_sc_hd__a21oi_4
X_65774_ _65969_/A _65855_/A sky130_fd_sc_hd__buf_2
X_62986_ _64328_/A _63516_/A sky130_fd_sc_hd__buf_2
X_67513_ _67513_/A _87212_/Q _67513_/X sky130_fd_sc_hd__and2_4
X_64725_ _64725_/A _64883_/A sky130_fd_sc_hd__buf_2
X_49659_ _49655_/Y _49650_/X _49658_/X _86347_/D sky130_fd_sc_hd__a21oi_4
X_61937_ _59823_/X _61937_/X sky130_fd_sc_hd__buf_2
X_80771_ _80818_/CLK _75888_/Y _80771_/Q sky130_fd_sc_hd__dfxtp_4
X_68493_ _68384_/A _68493_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_280_0_CLK clkbuf_9_281_0_CLK/A clkbuf_9_280_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_7_39_0_CLK clkbuf_7_39_0_CLK/A clkbuf_8_79_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_82510_ _82491_/CLK _82510_/D _82510_/Q sky130_fd_sc_hd__dfxtp_4
X_67444_ _67517_/A _67444_/B _67444_/X sky130_fd_sc_hd__and2_4
X_52670_ _52668_/Y _52647_/X _52669_/X _85776_/D sky130_fd_sc_hd__a21oi_4
X_64656_ _64656_/A _64809_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_179_0_CLK clkbuf_7_89_0_CLK/X clkbuf_8_179_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_83490_ _83491_/CLK _71461_/X _83490_/Q sky130_fd_sc_hd__dfxtp_4
X_61868_ _61787_/X _61915_/D sky130_fd_sc_hd__buf_2
Xclkbuf_10_174_0_CLK clkbuf_9_87_0_CLK/X _83914_/CLK sky130_fd_sc_hd__clkbuf_1
X_51621_ _51621_/A _51621_/X sky130_fd_sc_hd__buf_2
X_63607_ _63655_/A _58487_/A _63581_/X _63595_/D _63607_/X sky130_fd_sc_hd__and4_4
X_82441_ _82820_/CLK _79133_/X _82409_/D sky130_fd_sc_hd__dfxtp_4
X_60819_ _59532_/A _60630_/C _60630_/A _61277_/B sky130_fd_sc_hd__nand3_4
X_67375_ _67372_/X _67374_/X _67255_/X _67375_/Y sky130_fd_sc_hd__a21oi_4
X_64587_ _64676_/A _85857_/Q _64587_/X sky130_fd_sc_hd__and2_4
X_61799_ _61863_/A _61794_/Y _61795_/Y _61798_/Y _61799_/Y sky130_fd_sc_hd__nand4_4
X_69114_ _69958_/A _69114_/B _69114_/Y sky130_fd_sc_hd__nor2_4
X_54340_ _54337_/Y _54338_/X _54339_/X _85460_/D sky130_fd_sc_hd__a21oi_4
X_66326_ _66326_/A _66326_/B _66326_/X sky130_fd_sc_hd__and2_4
X_85160_ _83016_/CLK _56532_/Y _85160_/Q sky130_fd_sc_hd__dfxtp_4
X_51552_ _51552_/A _51553_/C sky130_fd_sc_hd__buf_2
X_63538_ _61499_/B _63487_/X _63535_/X _63537_/X _63538_/X sky130_fd_sc_hd__a211o_4
X_82372_ _84951_/CLK _82180_/Q _82372_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_295_0_CLK clkbuf_9_295_0_CLK/A clkbuf_9_295_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_8_102_0_CLK clkbuf_7_51_0_CLK/X clkbuf_8_102_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_84111_ _84111_/CLK _66502_/X _84111_/Q sky130_fd_sc_hd__dfxtp_4
X_50503_ _50556_/A _50503_/B _50503_/Y sky130_fd_sc_hd__nand2_4
X_81323_ _81344_/CLK _76287_/X _81699_/D sky130_fd_sc_hd__dfxtp_4
X_69045_ _68770_/X _69045_/B _69045_/X sky130_fd_sc_hd__and2_4
X_54271_ _54269_/Y _54051_/X _54270_/X _54271_/Y sky130_fd_sc_hd__a21oi_4
X_66257_ _66225_/X _84969_/Q _66186_/X _66256_/X _66257_/X sky130_fd_sc_hd__a211o_4
X_85091_ _85100_/CLK _85091_/D _85091_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_189_0_CLK clkbuf_9_94_0_CLK/X _81074_/CLK sky130_fd_sc_hd__clkbuf_1
X_51483_ _51473_/A _51494_/B _51494_/C _53008_/D _51483_/X sky130_fd_sc_hd__and4_4
X_63469_ _63517_/A _63517_/B _84321_/Q _63469_/Y sky130_fd_sc_hd__nor3_4
X_56010_ _55997_/X _74312_/C _74310_/C _56010_/X sky130_fd_sc_hd__and3_4
X_53222_ _53302_/A _53222_/X sky130_fd_sc_hd__buf_2
X_65208_ _65208_/A _65207_/X _65208_/Y sky130_fd_sc_hd__nand2_4
X_84042_ _81475_/CLK _84042_/D _81474_/D sky130_fd_sc_hd__dfxtp_4
X_50434_ _53511_/A _50456_/B sky130_fd_sc_hd__buf_2
X_81254_ _81671_/CLK _81286_/Q _76200_/A sky130_fd_sc_hd__dfxtp_4
X_66188_ _66040_/X _84974_/Q _66186_/X _66187_/X _66188_/X sky130_fd_sc_hd__a211o_4
X_80205_ _84949_/Q _84197_/Q _80205_/X sky130_fd_sc_hd__xor2_4
X_53153_ _53147_/X _53153_/B _53153_/Y sky130_fd_sc_hd__nand2_4
X_65139_ _65134_/X _64937_/B _65138_/X _65139_/Y sky130_fd_sc_hd__nand3_4
X_50365_ _50383_/A _50365_/B _50365_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_117_0_CLK clkbuf_7_58_0_CLK/X clkbuf_9_235_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_81185_ _86758_/CLK _75074_/X _81185_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_112_0_CLK clkbuf_9_56_0_CLK/X _84400_/CLK sky130_fd_sc_hd__clkbuf_1
X_52104_ _52101_/Y _52049_/X _52103_/X _52104_/Y sky130_fd_sc_hd__a21oi_4
X_87801_ _87285_/CLK _42613_/Y _73415_/A sky130_fd_sc_hd__dfxtp_4
X_80136_ _80114_/A _80126_/X _80136_/Y sky130_fd_sc_hd__nand2_4
X_57961_ _57868_/X _57958_/Y _57960_/Y _57899_/X _57872_/X _57961_/X
+ sky130_fd_sc_hd__o32a_4
X_53084_ _53107_/A _53069_/X _53074_/C _53084_/D _53084_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_742_0_CLK clkbuf_9_371_0_CLK/X _88002_/CLK sky130_fd_sc_hd__clkbuf_1
X_69947_ _42057_/A _69837_/X _69088_/X _69946_/Y _69947_/X sky130_fd_sc_hd__a211o_4
X_50296_ _50294_/Y _50274_/X _50295_/Y _86229_/D sky130_fd_sc_hd__a21boi_4
X_85993_ _85993_/CLK _85993_/D _85993_/Q sky130_fd_sc_hd__dfxtp_4
X_59700_ _59797_/A _59700_/Y sky130_fd_sc_hd__inv_2
X_52035_ _52032_/Y _51987_/X _52034_/X _85902_/D sky130_fd_sc_hd__a21oi_4
X_56912_ _56912_/A _57272_/D sky130_fd_sc_hd__inv_2
X_87732_ _87990_/CLK _87732_/D _69122_/B sky130_fd_sc_hd__dfxtp_4
X_84944_ _85492_/CLK _57865_/Y _84944_/Q sky130_fd_sc_hd__dfxtp_4
X_80067_ _80059_/X _80060_/X _80066_/Y _80071_/A sky130_fd_sc_hd__a21boi_4
X_57892_ _86646_/Q _57791_/X _57892_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_9_233_0_CLK clkbuf_8_116_0_CLK/X clkbuf_9_233_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_69878_ _87048_/Q _69690_/X _68473_/X _69877_/X _69878_/X sky130_fd_sc_hd__a211o_4
X_59631_ _59689_/B _59631_/B _65680_/A _59631_/Y sky130_fd_sc_hd__nand3_4
X_56843_ _56721_/D _56842_/X _56843_/Y sky130_fd_sc_hd__nand2_4
X_68829_ _69648_/A _43644_/Y _68829_/Y sky130_fd_sc_hd__nor2_4
X_87663_ _82896_/CLK _87663_/D _87663_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_127_0_CLK clkbuf_9_63_0_CLK/X _84518_/CLK sky130_fd_sc_hd__clkbuf_1
X_84875_ _84877_/CLK _84875_/D _58335_/A sky130_fd_sc_hd__dfxtp_4
X_86614_ _85969_/CLK _86614_/D _86614_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_757_0_CLK clkbuf_9_378_0_CLK/X _88084_/CLK sky130_fd_sc_hd__clkbuf_1
X_71840_ _71824_/Y _83356_/Q _71839_/X _83356_/D sky130_fd_sc_hd__a21o_4
X_59562_ _59557_/X _59562_/B _59544_/D _60122_/A sky130_fd_sc_hd__nand3_4
X_83826_ _83187_/CLK _83826_/D _83826_/Q sky130_fd_sc_hd__dfxtp_4
X_56774_ _56774_/A _85133_/Q _56774_/C _56774_/Y sky130_fd_sc_hd__nor3_4
X_87594_ _88111_/CLK _87594_/D _73773_/A sky130_fd_sc_hd__dfxtp_4
X_53986_ _85528_/Q _53955_/X _53985_/Y _53986_/Y sky130_fd_sc_hd__o21ai_4
X_58513_ _58513_/A _58513_/Y sky130_fd_sc_hd__inv_2
X_55725_ _56452_/C _55126_/A _55128_/A _55724_/X _55725_/X sky130_fd_sc_hd__a211o_4
X_86545_ _86222_/CLK _86545_/D _86545_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_248_0_CLK clkbuf_8_124_0_CLK/X clkbuf_9_248_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_40951_ _40944_/X _40946_/X _40950_/X _88305_/Q _40916_/X _40952_/A
+ sky130_fd_sc_hd__o32ai_4
X_52937_ _85727_/Q _52929_/X _52936_/Y _52937_/Y sky130_fd_sc_hd__o21ai_4
X_59493_ _59493_/A _59493_/Y sky130_fd_sc_hd__inv_2
X_71771_ _71762_/X _83382_/Q _71770_/X _71771_/X sky130_fd_sc_hd__a21o_4
X_83757_ _83761_/CLK _70519_/Y _57668_/A sky130_fd_sc_hd__dfxtp_4
X_80969_ _80776_/CLK _75635_/X _75475_/B sky130_fd_sc_hd__dfxtp_4
X_73510_ _43201_/Y _73298_/X _73464_/X _73509_/Y _73510_/X sky130_fd_sc_hd__a211o_4
X_70722_ _70722_/A _70713_/X _70727_/C _70769_/D _70722_/Y sky130_fd_sc_hd__nand4_4
X_58444_ _84846_/Q _63230_/A sky130_fd_sc_hd__inv_2
X_82708_ _82803_/CLK _78975_/X _82664_/D sky130_fd_sc_hd__dfxtp_4
X_43670_ _40749_/X _43656_/X _74226_/A _43657_/X _87318_/D sky130_fd_sc_hd__a2bb2o_4
X_55656_ _55656_/A _55656_/X sky130_fd_sc_hd__buf_2
X_74490_ _74490_/A _48647_/Y _74490_/Y sky130_fd_sc_hd__nand2_4
X_86476_ _86505_/CLK _48824_/Y _86476_/Q sky130_fd_sc_hd__dfxtp_4
X_52868_ _52864_/Y _52865_/X _52867_/X _52868_/Y sky130_fd_sc_hd__a21oi_4
X_40882_ _40881_/X _40821_/X _88318_/Q _40822_/X _40882_/X sky130_fd_sc_hd__a2bb2o_4
X_83688_ _83685_/CLK _70837_/Y _46624_/A sky130_fd_sc_hd__dfxtp_4
X_88215_ _88215_/CLK _88215_/D _88215_/Q sky130_fd_sc_hd__dfxtp_4
X_54607_ _54589_/X _54607_/B _54591_/C _47208_/Y _54607_/X sky130_fd_sc_hd__and4_4
X_42621_ _49210_/B _40921_/A _41888_/X _42620_/Y _42612_/X _42621_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73441_ _43741_/Y _73030_/X _72858_/X _73440_/Y _73441_/X sky130_fd_sc_hd__a211o_4
X_85427_ _85428_/CLK _54523_/Y _85427_/Q sky130_fd_sc_hd__dfxtp_4
X_51819_ _53269_/A _51820_/A sky130_fd_sc_hd__buf_2
X_70653_ _70722_/A _70656_/B _70642_/X _70656_/D _70653_/Y sky130_fd_sc_hd__nand4_4
X_82639_ _84003_/CLK _82639_/D _78921_/A sky130_fd_sc_hd__dfxtp_4
X_58375_ _58341_/X _58372_/Y _58374_/Y _84866_/D sky130_fd_sc_hd__a21oi_4
X_55587_ _55583_/X _55586_/X _44115_/A _55592_/A sky130_fd_sc_hd__a21o_4
X_52799_ _52803_/A _52799_/B _52799_/Y sky130_fd_sc_hd__nand2_4
XPHY_40 sky130_fd_sc_hd__decap_3
X_45340_ _55724_/B _45284_/X _45339_/X _45340_/X sky130_fd_sc_hd__o21a_4
XPHY_51 sky130_fd_sc_hd__decap_3
X_57326_ _57026_/X _57326_/B _57326_/C _57326_/Y sky130_fd_sc_hd__nor3_4
X_76160_ _76158_/X _76159_/Y _81635_/Q _76160_/X sky130_fd_sc_hd__a21o_4
X_88146_ _86834_/CLK _88146_/D _66609_/B sky130_fd_sc_hd__dfxtp_4
X_42552_ _42521_/X _42522_/X _40787_/X _87823_/Q _42540_/X _42553_/A
+ sky130_fd_sc_hd__o32ai_4
X_54538_ _54538_/A _54526_/B _54538_/C _47084_/A _54538_/X sky130_fd_sc_hd__and4_4
X_73372_ _73372_/A _73372_/B _73372_/Y sky130_fd_sc_hd__nor2_4
X_85358_ _86289_/CLK _85358_/D _85358_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_62 sky130_fd_sc_hd__decap_3
X_70584_ _70583_/X _70584_/X sky130_fd_sc_hd__buf_2
XPHY_73 sky130_fd_sc_hd__decap_3
XPHY_84 sky130_fd_sc_hd__decap_3
X_75111_ _75109_/A _75109_/B _75113_/C sky130_fd_sc_hd__nand2_4
X_41503_ _41502_/Y _41503_/X sky130_fd_sc_hd__buf_2
X_72323_ _72323_/A _72323_/Y sky130_fd_sc_hd__inv_2
XPHY_95 sky130_fd_sc_hd__decap_3
X_84309_ _84314_/CLK _63616_/Y _80413_/B sky130_fd_sc_hd__dfxtp_4
X_57257_ _57359_/A _45553_/A _57249_/X _57257_/Y sky130_fd_sc_hd__nor3_4
X_45271_ _83017_/Q _45273_/A sky130_fd_sc_hd__inv_2
X_76091_ _81722_/D _76092_/B _76094_/A sky130_fd_sc_hd__nor2_4
X_88077_ _88081_/CLK _88077_/D _41996_/A sky130_fd_sc_hd__dfxtp_4
X_54469_ _54478_/A _54469_/B _54469_/Y sky130_fd_sc_hd__nand2_4
X_42483_ _73795_/A _68618_/B sky130_fd_sc_hd__inv_2
X_85289_ _83016_/CLK _56141_/Y _85289_/Q sky130_fd_sc_hd__dfxtp_4
X_47010_ _46961_/X _47029_/A sky130_fd_sc_hd__buf_2
X_56208_ _56200_/X _56205_/X _56208_/C _56208_/Y sky130_fd_sc_hd__nand3_4
X_44222_ _68057_/A _69751_/A sky130_fd_sc_hd__buf_2
X_75042_ _75042_/A _75042_/B _75042_/Y sky130_fd_sc_hd__nand2_4
X_87028_ _87032_/CLK _44627_/Y _87028_/Q sky130_fd_sc_hd__dfxtp_4
X_41434_ _41433_/X _41418_/X _88216_/Q _41419_/X _41434_/X sky130_fd_sc_hd__a2bb2o_4
X_72254_ _72137_/X _72251_/Y _72253_/Y _72194_/X _72141_/X _72254_/X
+ sky130_fd_sc_hd__o32a_4
X_57188_ _57188_/A _44239_/A _56818_/X _57188_/Y sky130_fd_sc_hd__nand3_4
X_71205_ _71197_/A _71228_/B _71197_/C _71205_/Y sky130_fd_sc_hd__nand3_4
X_44153_ _44265_/D _44153_/X sky130_fd_sc_hd__buf_2
X_56139_ _56138_/Y _56139_/X sky130_fd_sc_hd__buf_2
X_79850_ _79839_/X _79850_/Y sky130_fd_sc_hd__inv_2
X_41365_ _41358_/X _82898_/Q _41365_/X sky130_fd_sc_hd__or2_4
X_72185_ _59297_/A _72185_/X sky130_fd_sc_hd__buf_2
X_43104_ _43046_/X _43047_/X _40749_/X _43103_/Y _43090_/X _87574_/D
+ sky130_fd_sc_hd__o32ai_4
X_78801_ _78801_/A _78801_/B _78801_/Y sky130_fd_sc_hd__nand2_4
X_71136_ _71136_/A _70758_/C _70827_/C _70627_/A _71137_/B sky130_fd_sc_hd__nand4_4
X_48961_ _48957_/Y _48935_/X _48960_/X _86458_/D sky130_fd_sc_hd__a21oi_4
X_44084_ _43986_/A _87174_/Q _44085_/D sky130_fd_sc_hd__nand2_4
X_79781_ _79774_/X _79781_/B _79781_/Y sky130_fd_sc_hd__nand2_4
X_41296_ _81759_/Q _41292_/B _41296_/X sky130_fd_sc_hd__or2_4
X_76993_ _84545_/Q _76993_/B _76993_/X sky130_fd_sc_hd__xor2_4
X_47912_ _47912_/A _50268_/B _47912_/Y sky130_fd_sc_hd__nand2_4
X_43035_ _42060_/X _43031_/X _40590_/X _43032_/Y _43034_/X _43035_/Y
+ sky130_fd_sc_hd__o32ai_4
X_78732_ _78732_/A _78732_/B _78732_/C _78732_/X sky130_fd_sc_hd__or3_4
Xclkbuf_0_CLK CLK clkbuf_0_CLK/X sky130_fd_sc_hd__clkbuf_16
X_71067_ _48955_/X _71046_/X _71066_/Y _71067_/Y sky130_fd_sc_hd__o21ai_4
X_75944_ _81509_/Q _75944_/B _81790_/D sky130_fd_sc_hd__xor2_4
X_48892_ _48606_/X _81216_/Q _48891_/Y _48893_/A sky130_fd_sc_hd__o21ai_4
X_70018_ _82552_/D _70010_/X _70017_/X _83872_/D sky130_fd_sc_hd__a21bo_4
X_47843_ _73591_/A _50224_/B sky130_fd_sc_hd__buf_2
X_59829_ _59875_/A _59829_/X sky130_fd_sc_hd__buf_2
X_78663_ _78663_/A _78663_/B _78663_/C _78663_/X sky130_fd_sc_hd__or3_4
X_75875_ _75862_/Y _75875_/B _75875_/C _75876_/B sky130_fd_sc_hd__nand3_4
X_77614_ _77614_/A _77614_/B _77614_/C _77614_/X sky130_fd_sc_hd__or3_4
X_74826_ _74826_/A _74826_/Y sky130_fd_sc_hd__inv_2
X_62840_ _62837_/X _62838_/X _62839_/Y _84378_/D sky130_fd_sc_hd__a21oi_4
X_47774_ _72428_/A _47760_/X _47773_/Y _47774_/Y sky130_fd_sc_hd__o21ai_4
X_78594_ _82517_/Q _82773_/D _78594_/X sky130_fd_sc_hd__xor2_4
X_44986_ _45212_/A _44986_/X sky130_fd_sc_hd__buf_2
X_49513_ _58920_/B _49496_/X _49512_/Y _49513_/Y sky130_fd_sc_hd__o21ai_4
X_46725_ _46725_/A _46915_/A sky130_fd_sc_hd__buf_2
X_77545_ _77508_/A _77511_/A _77520_/B _77561_/A sky130_fd_sc_hd__a21o_4
X_43937_ _43937_/A _43937_/Y sky130_fd_sc_hd__inv_2
X_62771_ _57660_/X _62749_/X _62768_/X _62759_/X _62770_/X _62771_/Y
+ sky130_fd_sc_hd__a41oi_4
X_74757_ _83843_/Q _74735_/X _74754_/X _74755_/X _74756_/X _74758_/C
+ sky130_fd_sc_hd__a2111oi_4
X_71969_ _72009_/A _71969_/X sky130_fd_sc_hd__buf_2
X_64510_ _64507_/Y _59655_/X _64509_/Y _64510_/Y sky130_fd_sc_hd__a21oi_4
X_49444_ _49444_/A _49454_/A sky130_fd_sc_hd__buf_2
X_61722_ _61722_/A _61752_/A sky130_fd_sc_hd__buf_2
X_73708_ _73605_/X _86235_/Q _73683_/X _73707_/X _73708_/X sky130_fd_sc_hd__a211o_4
X_46656_ _46845_/A _46682_/B sky130_fd_sc_hd__buf_2
X_65490_ _65453_/X _85597_/Q _65470_/X _65489_/X _65490_/X sky130_fd_sc_hd__a211o_4
X_77476_ _77476_/A _77473_/A _77476_/Y sky130_fd_sc_hd__nand2_4
X_43868_ _43842_/A _43868_/X sky130_fd_sc_hd__buf_2
X_74688_ _74694_/A _45787_/A _74688_/Y sky130_fd_sc_hd__nand2_4
X_79215_ _79215_/A _79215_/X sky130_fd_sc_hd__buf_2
X_45607_ _63158_/B _61492_/A sky130_fd_sc_hd__buf_2
X_76427_ _81269_/Q _81525_/D _76430_/B sky130_fd_sc_hd__nor2_4
X_64441_ _64432_/Y _64434_/X _64435_/X _64439_/Y _64440_/X _64441_/X
+ sky130_fd_sc_hd__o41a_4
X_42819_ _42818_/Y _87702_/D sky130_fd_sc_hd__inv_2
X_49375_ _49373_/Y _49316_/X _49374_/X _49375_/Y sky130_fd_sc_hd__a21oi_4
X_61653_ _72528_/A _61653_/X sky130_fd_sc_hd__buf_2
X_73639_ _73609_/X _85630_/Q _73472_/X _73638_/X _73639_/X sky130_fd_sc_hd__a211o_4
X_46587_ _46547_/A _51389_/B _46587_/Y sky130_fd_sc_hd__nand2_4
X_43799_ _43799_/A _43799_/Y sky130_fd_sc_hd__inv_2
X_48326_ _48320_/Y _48322_/X _48325_/Y _48326_/Y sky130_fd_sc_hd__a21boi_4
X_60604_ _79129_/A _60577_/X _60603_/X _60481_/X _60604_/Y sky130_fd_sc_hd__a2bb2oi_4
X_67160_ _67039_/X _67160_/X sky130_fd_sc_hd__buf_2
X_79146_ _79146_/A _84478_/Q _79146_/X sky130_fd_sc_hd__xor2_4
X_45538_ _85048_/Q _45490_/B _45538_/Y sky130_fd_sc_hd__nor2_4
X_64372_ _79742_/B _64314_/X _64371_/X _64372_/X sky130_fd_sc_hd__a21o_4
X_76358_ _76338_/B _76357_/Y _76358_/Y sky130_fd_sc_hd__nand2_4
X_61584_ _84844_/Q _61323_/B _61584_/X sky130_fd_sc_hd__or2_4
X_66111_ _58124_/A _72155_/A sky130_fd_sc_hd__buf_2
X_63323_ _63289_/X _64525_/C _63341_/C _63332_/D _63323_/X sky130_fd_sc_hd__and4_4
X_75309_ _75309_/A _75308_/Y _81042_/D sky130_fd_sc_hd__xor2_4
X_60535_ _59772_/A _59837_/B _79144_/A _60535_/Y sky130_fd_sc_hd__nor3_4
X_48257_ _48229_/A _48257_/B _48257_/Y sky130_fd_sc_hd__nand2_4
X_67091_ _84084_/Q _66971_/X _67090_/X _84084_/D sky130_fd_sc_hd__a21bo_4
X_79077_ _79076_/Y _79077_/Y sky130_fd_sc_hd__inv_2
X_45469_ _45462_/X _45466_/X _45468_/Y _86875_/D sky130_fd_sc_hd__a21oi_4
X_76289_ _76289_/A _81560_/Q _76290_/B sky130_fd_sc_hd__xor2_4
X_47208_ _82371_/Q _47208_/Y sky130_fd_sc_hd__inv_2
X_66042_ _66040_/X _84984_/Q _66027_/X _66041_/X _66042_/X sky130_fd_sc_hd__a211o_4
X_78028_ _82257_/Q _81969_/Q _78028_/X sky130_fd_sc_hd__xor2_4
X_63254_ _63253_/X _63254_/Y sky130_fd_sc_hd__inv_2
X_48188_ _48478_/A _48188_/X sky130_fd_sc_hd__buf_2
X_60466_ _60420_/A _60466_/X sky130_fd_sc_hd__buf_2
X_62205_ _62620_/A _62249_/A sky130_fd_sc_hd__buf_2
X_47139_ _46902_/A _47140_/A sky130_fd_sc_hd__buf_2
X_63185_ _59419_/A _63170_/X _63161_/C _63149_/X _63185_/X sky130_fd_sc_hd__or4_4
X_60397_ _60459_/B _60473_/B sky130_fd_sc_hd__buf_2
X_69801_ _69374_/X _69377_/X _69728_/X _69801_/Y sky130_fd_sc_hd__a21oi_4
X_50150_ _65096_/B _50137_/X _50149_/Y _50150_/Y sky130_fd_sc_hd__o21ai_4
X_62136_ _61949_/A _62170_/B _62158_/C _63314_/B _62136_/X sky130_fd_sc_hd__and4_4
X_67993_ _87140_/Q _67942_/X _67991_/X _67992_/X _67993_/X sky130_fd_sc_hd__a211o_4
X_79979_ _79978_/Y _79968_/Y _79980_/B sky130_fd_sc_hd__nand2_4
X_69732_ _64732_/A _69732_/X sky130_fd_sc_hd__buf_2
X_50081_ _64755_/B _50061_/X _50080_/Y _50081_/Y sky130_fd_sc_hd__o21ai_4
X_66944_ _66940_/X _66943_/X _66871_/X _66944_/Y sky130_fd_sc_hd__a21oi_4
X_62067_ _62056_/X _62058_/X _62066_/Y _58457_/A _62048_/X _62067_/Y
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_10_1014_0_CLK clkbuf_9_507_0_CLK/X _85581_/CLK sky130_fd_sc_hd__clkbuf_1
X_82990_ _85134_/CLK _74672_/Y _82990_/Q sky130_fd_sc_hd__dfxtp_4
X_61018_ _60866_/A _60962_/A _61018_/Y sky130_fd_sc_hd__nand2_4
X_81941_ _82131_/CLK _81941_/D _81941_/Q sky130_fd_sc_hd__dfxtp_4
X_69663_ _69660_/X _69662_/X _68697_/X _69663_/X sky130_fd_sc_hd__a21o_4
X_66875_ _66758_/X _66875_/X sky130_fd_sc_hd__buf_2
X_68614_ _68614_/A _69685_/A sky130_fd_sc_hd__buf_2
X_53840_ _53837_/Y _53838_/X _53839_/Y _53840_/Y sky130_fd_sc_hd__a21boi_4
X_65826_ _65824_/X _83055_/Q _65707_/X _65825_/X _65827_/B sky130_fd_sc_hd__a211o_4
X_84660_ _84660_/CLK _60108_/Y _60107_/C sky130_fd_sc_hd__dfxtp_4
X_81872_ _81872_/CLK _78063_/X _81840_/D sky130_fd_sc_hd__dfxtp_4
X_69594_ _68360_/X _42548_/Y _69594_/Y sky130_fd_sc_hd__nor2_4
X_83611_ _83613_/CLK _71089_/Y _83611_/Q sky130_fd_sc_hd__dfxtp_4
X_68545_ _68517_/A _68545_/X sky130_fd_sc_hd__buf_2
X_80823_ _80962_/CLK _83967_/Q _75612_/B sky130_fd_sc_hd__dfxtp_4
X_53771_ _85571_/Q _53754_/X _53770_/Y _53771_/Y sky130_fd_sc_hd__o21ai_4
X_65757_ _65757_/A _65757_/X sky130_fd_sc_hd__buf_2
X_84591_ _84458_/CLK _60597_/Y _79131_/A sky130_fd_sc_hd__dfxtp_4
X_50983_ _50957_/A _50983_/X sky130_fd_sc_hd__buf_2
X_62969_ _62988_/A _62988_/B _84365_/Q _62969_/Y sky130_fd_sc_hd__nor3_4
X_55510_ _55470_/A _55510_/X sky130_fd_sc_hd__buf_2
X_86330_ _86647_/CLK _49752_/Y _57832_/B sky130_fd_sc_hd__dfxtp_4
X_52722_ _52718_/A _52722_/B _52722_/Y sky130_fd_sc_hd__nand2_4
X_64708_ _58784_/A _64898_/A sky130_fd_sc_hd__buf_2
X_83542_ _86222_/CLK _83542_/D _83542_/Q sky130_fd_sc_hd__dfxtp_4
X_56490_ _56487_/X _56484_/X _85176_/Q _56490_/Y sky130_fd_sc_hd__nand3_4
X_80754_ _80754_/CLK _80754_/D _81130_/D sky130_fd_sc_hd__dfxtp_4
X_68476_ _87003_/Q _68472_/X _68473_/X _68475_/X _68476_/X sky130_fd_sc_hd__a211o_4
X_65688_ _65685_/X _86192_/Q _65534_/X _65687_/X _65688_/X sky130_fd_sc_hd__a211o_4
X_55441_ _55441_/A _55441_/B _55441_/C _55442_/A sky130_fd_sc_hd__nand3_4
X_67427_ _67333_/A _87663_/Q _67427_/X sky130_fd_sc_hd__and2_4
X_86261_ _85555_/CLK _86261_/D _64931_/B sky130_fd_sc_hd__dfxtp_4
X_52653_ _52626_/A _52654_/C sky130_fd_sc_hd__buf_2
X_64639_ _64634_/Y _60349_/X _64638_/X _84232_/D sky130_fd_sc_hd__a21o_4
X_83473_ _86600_/CLK _83473_/D _47751_/A sky130_fd_sc_hd__dfxtp_4
X_80685_ _81074_/CLK _80685_/D _75226_/A sky130_fd_sc_hd__dfxtp_4
X_88000_ _88001_/CLK _88000_/D _88000_/Q sky130_fd_sc_hd__dfxtp_4
X_85212_ _85244_/CLK _85212_/D _56390_/C sky130_fd_sc_hd__dfxtp_4
X_51604_ _51601_/Y _51585_/X _51603_/X _85980_/D sky130_fd_sc_hd__a21oi_4
X_58160_ _61368_/A _58160_/B _58160_/Y sky130_fd_sc_hd__nand2_4
XPHY_605 sky130_fd_sc_hd__decap_3
X_82424_ _84177_/CLK _82456_/Q _78630_/A sky130_fd_sc_hd__dfxtp_4
X_55372_ _55371_/X _55375_/A sky130_fd_sc_hd__inv_2
X_67358_ _67120_/X _67358_/X sky130_fd_sc_hd__buf_2
X_86192_ _83562_/CLK _50484_/Y _86192_/Q sky130_fd_sc_hd__dfxtp_4
X_52584_ _52588_/A _52594_/B _51919_/C _51756_/D _52584_/X sky130_fd_sc_hd__and4_4
XPHY_616 sky130_fd_sc_hd__decap_3
XPHY_627 sky130_fd_sc_hd__decap_3
XPHY_638 sky130_fd_sc_hd__decap_3
X_57111_ _57109_/X _56607_/X _45500_/A _57110_/X _85082_/D sky130_fd_sc_hd__a2bb2o_4
X_54323_ _54332_/A _52632_/B _54323_/Y sky130_fd_sc_hd__nand2_4
X_66309_ _66266_/X _86213_/Q _66295_/X _66308_/X _66309_/X sky130_fd_sc_hd__a211o_4
XPHY_649 sky130_fd_sc_hd__decap_3
X_85143_ _85057_/CLK _56628_/Y _56627_/B sky130_fd_sc_hd__dfxtp_4
X_51535_ _51514_/A _53060_/B _51535_/Y sky130_fd_sc_hd__nand2_4
X_58091_ _58043_/X _85990_/Q _58090_/X _58091_/Y sky130_fd_sc_hd__o21ai_4
X_82355_ _82343_/CLK _77178_/X _47982_/A sky130_fd_sc_hd__dfxtp_4
X_67289_ _67286_/X _67288_/X _67264_/X _67292_/A sky130_fd_sc_hd__a21o_4
X_81306_ _81304_/CLK _76994_/X _81306_/Q sky130_fd_sc_hd__dfxtp_4
X_57042_ _56837_/X _57331_/C sky130_fd_sc_hd__buf_2
X_69028_ _44738_/A _68818_/X _68819_/X _69027_/X _69029_/B sky130_fd_sc_hd__a211o_4
X_54254_ _54254_/A _54255_/C sky130_fd_sc_hd__buf_2
X_85074_ _85074_/CLK _85074_/D _85074_/Q sky130_fd_sc_hd__dfxtp_4
X_51466_ _51218_/X _51473_/A sky130_fd_sc_hd__buf_2
X_82286_ _82288_/CLK _81910_/Q _82286_/Q sky130_fd_sc_hd__dfxtp_4
X_53205_ _53219_/A _53205_/B _53205_/Y sky130_fd_sc_hd__nand2_4
X_84025_ _81169_/CLK _84025_/D _82065_/D sky130_fd_sc_hd__dfxtp_4
X_50417_ _50556_/A _52119_/B _50417_/Y sky130_fd_sc_hd__nand2_4
X_81237_ _85332_/CLK _81045_/Q _81237_/Q sky130_fd_sc_hd__dfxtp_4
X_54185_ _85488_/Q _54167_/X _54184_/Y _54185_/Y sky130_fd_sc_hd__o21ai_4
X_51397_ _51395_/Y _51391_/X _51396_/X _51397_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_681_0_CLK clkbuf_9_340_0_CLK/X _87646_/CLK sky130_fd_sc_hd__clkbuf_1
X_41150_ _41143_/X _40624_/A _41149_/X _41151_/A sky130_fd_sc_hd__o21ai_4
X_53136_ _85690_/Q _53120_/X _53135_/Y _53136_/Y sky130_fd_sc_hd__o21ai_4
X_50348_ _50346_/Y _50313_/X _50347_/X _86219_/D sky130_fd_sc_hd__a21oi_4
X_81168_ _81179_/CLK _74949_/B _81168_/Q sky130_fd_sc_hd__dfxtp_4
X_58993_ _62186_/A _58993_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_9_172_0_CLK clkbuf_8_86_0_CLK/X clkbuf_9_172_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_80119_ _80098_/B _80115_/X _80118_/Y _80119_/Y sky130_fd_sc_hd__a21oi_4
X_41081_ _41073_/X _81703_/Q _41080_/X _41081_/X sky130_fd_sc_hd__o21a_4
X_53067_ _53080_/A _53067_/B _53067_/Y sky130_fd_sc_hd__nand2_4
X_57944_ _84937_/Q _57944_/Y sky130_fd_sc_hd__inv_2
X_50279_ _50228_/X _50279_/X sky130_fd_sc_hd__buf_2
X_73990_ _43644_/Y _72853_/X _73920_/X _73989_/Y _73990_/X sky130_fd_sc_hd__a211o_4
X_85976_ _85688_/CLK _51626_/Y _85976_/Q sky130_fd_sc_hd__dfxtp_4
X_81099_ _83944_/CLK _79654_/Y _81099_/Q sky130_fd_sc_hd__dfxtp_4
X_52018_ _52016_/Y _51987_/X _52017_/X _52018_/Y sky130_fd_sc_hd__a21oi_4
X_87715_ _87394_/CLK _87715_/D _67727_/B sky130_fd_sc_hd__dfxtp_4
X_72941_ _72939_/X _72940_/Y _72766_/X _72941_/Y sky130_fd_sc_hd__a21oi_4
X_84927_ _86627_/CLK _84927_/D _84927_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_696_0_CLK clkbuf_9_348_0_CLK/X _87189_/CLK sky130_fd_sc_hd__clkbuf_1
X_57875_ _58703_/A _57875_/X sky130_fd_sc_hd__buf_2
X_59614_ _59613_/Y _60162_/A sky130_fd_sc_hd__buf_2
X_44840_ _41715_/A _44838_/X _67719_/B _44839_/X _44840_/X sky130_fd_sc_hd__a2bb2o_4
X_56826_ _56823_/Y _56825_/Y _44137_/A _56827_/B sky130_fd_sc_hd__a21o_4
X_75660_ _75660_/A _75660_/B _75665_/A sky130_fd_sc_hd__nand2_4
X_87646_ _87646_/CLK _87646_/D _67832_/B sky130_fd_sc_hd__dfxtp_4
X_72872_ _72870_/X _86205_/Q _45930_/X _72871_/X _72872_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_9_187_0_CLK clkbuf_8_93_0_CLK/X clkbuf_9_187_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_84858_ _84358_/CLK _58401_/X _58399_/A sky130_fd_sc_hd__dfxtp_4
X_74611_ _45290_/Y _74598_/X _74610_/X _83016_/D sky130_fd_sc_hd__o21ai_4
X_71823_ _71823_/A _70410_/Y _71713_/Y _70854_/A _71823_/Y sky130_fd_sc_hd__nor4_4
X_59545_ _59545_/A _59552_/B sky130_fd_sc_hd__inv_2
X_83809_ _83820_/CLK _83809_/D _74809_/A sky130_fd_sc_hd__dfxtp_4
X_44771_ _44766_/X _44767_/X _41346_/X _86964_/Q _44768_/X _44772_/A
+ sky130_fd_sc_hd__o32ai_4
X_56757_ _57023_/A _56785_/B sky130_fd_sc_hd__buf_2
X_75591_ _75589_/Y _75889_/A _75591_/Y sky130_fd_sc_hd__nand2_4
X_87577_ _87577_/CLK _87577_/D _87577_/Q sky130_fd_sc_hd__dfxtp_4
X_53969_ _53969_/A _53964_/B _53969_/C _53969_/X sky130_fd_sc_hd__and3_4
X_41983_ _88082_/Q _41983_/Y sky130_fd_sc_hd__inv_2
X_84789_ _86695_/CLK _84789_/D _84789_/Q sky130_fd_sc_hd__dfxtp_4
X_46510_ _83634_/Q _54054_/B sky130_fd_sc_hd__inv_2
X_77330_ _77308_/Y _77310_/A _77307_/A _77332_/C sky130_fd_sc_hd__o21ai_4
X_55708_ _83014_/Q _55272_/X _44095_/A _55707_/X _55708_/X sky130_fd_sc_hd__a211o_4
X_43722_ _40866_/A _43716_/X _69823_/B _43718_/X _43722_/X sky130_fd_sc_hd__a2bb2o_4
X_74542_ _55986_/X _74538_/Y _74541_/Y _83041_/D sky130_fd_sc_hd__o21ai_4
X_86528_ _86523_/CLK _48378_/Y _65444_/B sky130_fd_sc_hd__dfxtp_4
X_40934_ _40931_/X _41114_/A _40933_/X _40935_/A sky130_fd_sc_hd__o21ai_4
X_47490_ _47490_/A _53076_/B sky130_fd_sc_hd__buf_2
X_71754_ _52950_/B _71736_/X _71753_/Y _83388_/D sky130_fd_sc_hd__o21ai_4
X_59476_ _84721_/Q _59477_/A sky130_fd_sc_hd__buf_2
X_56688_ _56777_/B _56688_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_110_0_CLK clkbuf_8_55_0_CLK/X clkbuf_9_110_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_46441_ _83640_/Q _46441_/Y sky130_fd_sc_hd__inv_2
X_70705_ _70716_/A _70710_/C sky130_fd_sc_hd__buf_2
X_58427_ _58424_/Y _58426_/X _58427_/Y sky130_fd_sc_hd__nand2_4
X_77261_ _77261_/A _77260_/Y _82180_/D sky130_fd_sc_hd__xnor2_4
X_43653_ _43652_/X _43653_/Y sky130_fd_sc_hd__inv_2
X_55639_ _55636_/X _55638_/X _55615_/A _55643_/A sky130_fd_sc_hd__a21o_4
X_74473_ _74471_/Y _74463_/X _74472_/X _83059_/D sky130_fd_sc_hd__a21oi_4
X_86459_ _85561_/CLK _86459_/D _86459_/Q sky130_fd_sc_hd__dfxtp_4
X_40865_ _40857_/X _82286_/Q _40864_/X _40866_/A sky130_fd_sc_hd__o21a_4
X_71685_ _71641_/A _71685_/X sky130_fd_sc_hd__buf_2
X_79000_ _79000_/A _78999_/Y _79001_/B sky130_fd_sc_hd__xnor2_4
X_76212_ _76209_/Y _76211_/Y _76213_/B sky130_fd_sc_hd__xnor2_4
X_42604_ _73345_/A _42604_/Y sky130_fd_sc_hd__inv_2
X_49160_ _65319_/B _49153_/X _49159_/Y _49160_/Y sky130_fd_sc_hd__o21ai_4
X_73424_ _73353_/A _85863_/Q _73424_/X sky130_fd_sc_hd__and2_4
X_46372_ _46348_/X _48986_/A _46371_/X _51290_/B sky130_fd_sc_hd__o21ai_4
X_70636_ _70625_/Y _70637_/A sky130_fd_sc_hd__buf_2
X_58358_ _84869_/Q _63326_/A sky130_fd_sc_hd__inv_2
X_77192_ _77194_/A _77194_/B _77193_/A sky130_fd_sc_hd__or2_4
Xclkbuf_10_634_0_CLK clkbuf_9_317_0_CLK/X _82327_/CLK sky130_fd_sc_hd__clkbuf_1
X_43584_ _43583_/Y _51337_/A sky130_fd_sc_hd__buf_2
X_40796_ _82875_/Q _40779_/B _40796_/X sky130_fd_sc_hd__or2_4
X_48111_ _48075_/X _82919_/Q _48110_/X _48112_/B sky130_fd_sc_hd__o21ai_4
X_45323_ _45316_/X _45320_/Y _45322_/Y _45323_/Y sky130_fd_sc_hd__a21oi_4
X_76143_ _76143_/A _76143_/B _76145_/A sky130_fd_sc_hd__nand2_4
X_57309_ _57261_/X _57007_/X _57308_/Y _57310_/A sky130_fd_sc_hd__o21ai_4
X_88129_ _88386_/CLK _88129_/D _67003_/B sky130_fd_sc_hd__dfxtp_4
X_42535_ _42517_/X _40748_/Y _42477_/X _42534_/Y _42519_/X _87830_/D
+ sky130_fd_sc_hd__o32ai_4
X_49091_ _52365_/A _48940_/B _49091_/C _49091_/X sky130_fd_sc_hd__and3_4
X_73355_ _73355_/A _73355_/X sky130_fd_sc_hd__buf_2
X_70567_ _71887_/A _71865_/A sky130_fd_sc_hd__buf_2
X_58289_ _58271_/X _83407_/Q _58288_/Y _58289_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_9_125_0_CLK clkbuf_8_62_0_CLK/X clkbuf_9_125_0_CLK/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_9_52_0_CLK clkbuf_9_53_0_CLK/A clkbuf_9_52_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_48042_ _66198_/B _47998_/X _48041_/Y _48042_/Y sky130_fd_sc_hd__o21ai_4
X_60320_ _60317_/A _60319_/X _79722_/A _60320_/Y sky130_fd_sc_hd__nor3_4
X_72306_ _72196_/X _85330_/Q _72255_/X _72306_/X sky130_fd_sc_hd__o21a_4
X_45254_ _85194_/Q _45252_/X _45253_/X _45254_/Y sky130_fd_sc_hd__o21ai_4
X_76074_ _81527_/Q _76074_/B _76074_/X sky130_fd_sc_hd__xor2_4
X_42466_ _42610_/A _42466_/X sky130_fd_sc_hd__buf_2
X_73286_ _73210_/X _85581_/Q _73284_/X _73285_/X _73286_/X sky130_fd_sc_hd__a211o_4
X_70498_ _71115_/C _70700_/A _70700_/B _70609_/A _70502_/A sky130_fd_sc_hd__nand4_4
X_44205_ _44196_/B _56670_/A sky130_fd_sc_hd__buf_2
X_75025_ _81147_/D _75032_/B _75030_/A sky130_fd_sc_hd__xor2_4
X_79902_ _80264_/A _79900_/X _80263_/B _79902_/Y sky130_fd_sc_hd__a21boi_4
X_41417_ _40717_/X _41486_/A sky130_fd_sc_hd__buf_2
X_60251_ _60251_/A _60170_/A _60197_/C _60309_/D _60285_/A sky130_fd_sc_hd__nand4_4
X_72237_ _72358_/A _72237_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_649_0_CLK clkbuf_9_324_0_CLK/X _86965_/CLK sky130_fd_sc_hd__clkbuf_1
X_45185_ _45127_/X _61548_/B _45144_/X _45185_/Y sky130_fd_sc_hd__o21ai_4
X_42397_ _42397_/A _42397_/X sky130_fd_sc_hd__buf_2
X_44136_ _44135_/X _44137_/A sky130_fd_sc_hd__buf_2
X_79833_ _79828_/Y _79832_/Y _79833_/X sky130_fd_sc_hd__xor2_4
X_41348_ _41337_/X _41338_/X _41347_/X _67600_/B _41333_/X _41349_/A
+ sky130_fd_sc_hd__o32ai_4
X_60182_ _60182_/A _60182_/Y sky130_fd_sc_hd__inv_2
X_72168_ _72166_/X _85373_/Q _72167_/X _72168_/Y sky130_fd_sc_hd__o21ai_4
X_49993_ _72366_/B _49986_/X _49992_/Y _49993_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_67_0_CLK clkbuf_9_67_0_CLK/A clkbuf_9_67_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_71119_ _71112_/X _71073_/B _71119_/C _71119_/Y sky130_fd_sc_hd__nand3_4
X_48944_ _48901_/A _48944_/B _48944_/Y sky130_fd_sc_hd__nand2_4
X_44067_ _44054_/Y _44067_/B _44116_/B _44067_/Y sky130_fd_sc_hd__nand3_4
X_79764_ _79764_/A _79764_/B _79765_/B sky130_fd_sc_hd__xor2_4
X_64990_ _64985_/X _64988_/X _64989_/X _64990_/X sky130_fd_sc_hd__a21o_4
X_41279_ _41279_/A _41279_/Y sky130_fd_sc_hd__inv_2
X_72099_ _74391_/A _50710_/B _72099_/Y sky130_fd_sc_hd__nand2_4
X_76976_ _76976_/A _84400_/Q _76976_/X sky130_fd_sc_hd__xor2_4
X_43018_ _41869_/A _42447_/C _41869_/C _43018_/Y sky130_fd_sc_hd__nor3_4
X_78715_ _78689_/Y _78690_/Y _78691_/Y _78715_/X sky130_fd_sc_hd__o21a_4
X_75927_ _81699_/D _75927_/B _75927_/X sky130_fd_sc_hd__xor2_4
X_63941_ _61481_/X _63908_/B _63894_/C _63908_/D _63941_/Y sky130_fd_sc_hd__nand4_4
X_48875_ _48873_/Y _48865_/X _48874_/X _86466_/D sky130_fd_sc_hd__a21oi_4
X_79695_ _79686_/Y _79704_/B _79694_/X _79696_/B sky130_fd_sc_hd__a21boi_4
X_47826_ _82369_/Q _48361_/B sky130_fd_sc_hd__inv_2
X_66660_ _66499_/B _66650_/Y _59782_/X _66659_/Y _66660_/X sky130_fd_sc_hd__a211o_4
X_78646_ _78646_/A _82681_/D _78649_/B sky130_fd_sc_hd__nor2_4
X_63872_ _64012_/A _63902_/D sky130_fd_sc_hd__buf_2
X_75858_ _80927_/Q _75855_/Y _75857_/X _75858_/Y sky130_fd_sc_hd__o21ai_4
X_65611_ _64725_/A _65735_/A sky130_fd_sc_hd__buf_2
X_62823_ _62789_/A _59413_/Y _62848_/C _62789_/D _62823_/X sky130_fd_sc_hd__and4_4
X_74809_ _74809_/A _74796_/B _74796_/C _71016_/A _74810_/D sky130_fd_sc_hd__nand4_4
X_47757_ _47757_/A _53230_/D sky130_fd_sc_hd__buf_2
X_66591_ _87442_/Q _66538_/X _66540_/X _66590_/X _66591_/X sky130_fd_sc_hd__a211o_4
X_78577_ _78561_/B _78560_/B _78560_/A _78577_/X sky130_fd_sc_hd__and3_4
X_44969_ _44968_/X _45033_/B sky130_fd_sc_hd__buf_2
X_75789_ _75779_/Y _75789_/Y sky130_fd_sc_hd__inv_2
X_68330_ _82629_/D _68318_/X _68329_/X _83981_/D sky130_fd_sc_hd__a21bo_4
X_46708_ _46717_/A _46717_/B _46682_/C _46707_/X _46708_/X sky130_fd_sc_hd__and4_4
X_65542_ _65428_/X _83074_/Q _65540_/X _65541_/X _65543_/B sky130_fd_sc_hd__a211o_4
X_77528_ _77528_/A _82198_/D _81910_/D sky130_fd_sc_hd__xor2_4
X_62754_ _61428_/X _62743_/B _62742_/X _62729_/D _62754_/Y sky130_fd_sc_hd__nand4_4
X_47688_ _47696_/A _53187_/B _47688_/Y sky130_fd_sc_hd__nand2_4
X_49427_ _49418_/A _51812_/B _49427_/Y sky130_fd_sc_hd__nand2_4
X_61705_ _61704_/Y _61715_/A sky130_fd_sc_hd__buf_2
X_68261_ _67607_/X _67609_/X _68260_/X _68261_/Y sky130_fd_sc_hd__a21oi_4
X_46639_ _46670_/A _46647_/B _46659_/C _51761_/D _46639_/X sky130_fd_sc_hd__and4_4
X_65473_ _65469_/X _65472_/X _65457_/X _65473_/X sky130_fd_sc_hd__a21o_4
X_77459_ _77452_/A _77433_/A _77459_/X sky130_fd_sc_hd__and2_4
X_62685_ _62669_/A _63033_/A _62704_/C _62669_/D _62685_/X sky130_fd_sc_hd__and4_4
X_67212_ _67093_/X _67259_/A sky130_fd_sc_hd__buf_2
X_64424_ _64380_/X _58382_/A _64381_/X _64424_/Y sky130_fd_sc_hd__nand3_4
X_61636_ _61636_/A _61636_/B _61590_/C _61636_/Y sky130_fd_sc_hd__nand3_4
X_49358_ _51396_/A _49317_/X _49312_/C _49358_/X sky130_fd_sc_hd__and3_4
X_80470_ _80467_/Y _80451_/B _80469_/X _80471_/B sky130_fd_sc_hd__o21ai_4
X_68192_ _84016_/Q _68180_/X _68191_/X _84016_/D sky130_fd_sc_hd__a21bo_4
X_48309_ _48306_/Y _48273_/X _48308_/Y _86538_/D sky130_fd_sc_hd__a21boi_4
X_67143_ _87867_/Q _67117_/X _67046_/X _67142_/X _67143_/X sky130_fd_sc_hd__a211o_4
X_79129_ _79129_/A _79129_/B _82437_/D sky130_fd_sc_hd__xor2_4
X_64355_ _64336_/A _84821_/Q _64323_/X _64355_/Y sky130_fd_sc_hd__nand3_4
X_49289_ _49273_/A _50808_/B _49289_/Y sky130_fd_sc_hd__nand2_4
X_61567_ _61565_/X _61517_/X _61566_/Y _61567_/Y sky130_fd_sc_hd__a21oi_4
X_51320_ _51310_/X _51320_/B _51320_/Y sky130_fd_sc_hd__nand2_4
X_63306_ _63306_/A _63392_/B sky130_fd_sc_hd__buf_2
X_82140_ _82604_/CLK _77970_/X _82096_/D sky130_fd_sc_hd__dfxtp_4
X_60518_ _60488_/B _63004_/C _60556_/B _60518_/X sky130_fd_sc_hd__o21a_4
X_67074_ _66953_/X _67074_/X sky130_fd_sc_hd__buf_2
X_64286_ _64295_/A _64248_/B _64286_/C _64286_/X sky130_fd_sc_hd__and3_4
X_61498_ _61374_/A _61499_/A sky130_fd_sc_hd__buf_2
X_66025_ _65876_/X _85625_/Q _65976_/X _66024_/X _66025_/X sky130_fd_sc_hd__a211o_4
X_51251_ _51278_/A _51251_/B _51251_/X sky130_fd_sc_hd__and2_4
X_63237_ _60459_/B _63237_/X sky130_fd_sc_hd__buf_2
X_82071_ _81154_/CLK _82071_/D _82071_/Q sky130_fd_sc_hd__dfxtp_4
X_60449_ _60438_/A _60420_/A _60440_/X _60439_/X _60473_/C _60572_/B
+ sky130_fd_sc_hd__a41o_4
Xclkbuf_9_8_0_CLK clkbuf_8_4_0_CLK/X clkbuf_9_8_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_50202_ _50200_/Y _50191_/X _50201_/X _86244_/D sky130_fd_sc_hd__a21oi_4
X_81022_ _84210_/CLK _84230_/Q _81022_/Q sky130_fd_sc_hd__dfxtp_4
X_51182_ _51180_/Y _51175_/X _51181_/X _51182_/Y sky130_fd_sc_hd__a21oi_4
X_63168_ _63157_/X _63168_/B _63147_/C _63124_/D _63168_/X sky130_fd_sc_hd__and4_4
X_50133_ _50120_/A _50133_/B _50133_/Y sky130_fd_sc_hd__nand2_4
X_62119_ _61412_/A _62120_/A sky130_fd_sc_hd__buf_2
X_85830_ _85542_/CLK _52404_/Y _65313_/B sky130_fd_sc_hd__dfxtp_4
X_55990_ _56177_/A _45836_/X _55990_/C _55990_/Y sky130_fd_sc_hd__nand3_4
X_67976_ _87448_/Q _67953_/X _67954_/X _67975_/X _67976_/X sky130_fd_sc_hd__a211o_4
X_63099_ _60469_/X _63100_/A sky130_fd_sc_hd__buf_2
X_69715_ _69712_/X _69714_/X _69655_/X _69715_/Y sky130_fd_sc_hd__a21oi_4
X_50064_ _50064_/A _50084_/A sky130_fd_sc_hd__buf_2
X_54941_ _54888_/A _54955_/A sky130_fd_sc_hd__buf_2
X_66927_ _66851_/X _66927_/B _66927_/X sky130_fd_sc_hd__and2_4
X_85761_ _85761_/CLK _52751_/Y _85761_/Q sky130_fd_sc_hd__dfxtp_4
X_82973_ _82973_/CLK _82781_/Q _82973_/Q sky130_fd_sc_hd__dfxtp_4
X_87500_ _88012_/CLK _87500_/D _87500_/Q sky130_fd_sc_hd__dfxtp_4
X_84712_ _84355_/CLK _59677_/Y _80614_/A sky130_fd_sc_hd__dfxtp_4
X_57660_ _84959_/Q _57660_/X sky130_fd_sc_hd__buf_2
X_69646_ _69605_/A _72924_/A _69646_/X sky130_fd_sc_hd__and2_4
X_81924_ _82116_/CLK _78047_/Y _77262_/A sky130_fd_sc_hd__dfxtp_4
X_54872_ _85362_/Q _54865_/X _54871_/Y _54872_/Y sky130_fd_sc_hd__o21ai_4
X_66858_ _87123_/Q _66833_/X _66834_/X _66857_/X _66858_/X sky130_fd_sc_hd__a211o_4
X_85692_ _85692_/CLK _85692_/D _85692_/Q sky130_fd_sc_hd__dfxtp_4
X_56611_ _56629_/B _56580_/B _56616_/A _56616_/B _72654_/C _56611_/Y
+ sky130_fd_sc_hd__a41oi_4
X_87431_ _87436_/CLK _43418_/Y _87431_/Q sky130_fd_sc_hd__dfxtp_4
X_53823_ _53819_/A _71996_/B _53823_/Y sky130_fd_sc_hd__nand2_4
X_65809_ _64729_/A _65809_/X sky130_fd_sc_hd__buf_2
X_84643_ _84333_/CLK _84643_/D _79817_/A sky130_fd_sc_hd__dfxtp_4
X_57591_ _84973_/Q _57562_/X _57590_/Y _57591_/Y sky130_fd_sc_hd__o21ai_4
X_81855_ _81094_/CLK _81887_/Q _77674_/A sky130_fd_sc_hd__dfxtp_4
X_69577_ _69505_/X _69574_/Y _69516_/X _69576_/Y _69577_/X sky130_fd_sc_hd__a211o_4
X_66789_ _66769_/A _88202_/Q _66789_/X sky130_fd_sc_hd__and2_4
X_59330_ _59325_/X _59327_/Y _59328_/Y _59271_/X _59329_/X _59330_/X
+ sky130_fd_sc_hd__o32a_4
X_56542_ _56538_/A _56535_/X _55715_/B _56542_/Y sky130_fd_sc_hd__nand3_4
X_80806_ _83973_/CLK _80806_/D _75750_/B sky130_fd_sc_hd__dfxtp_4
X_68528_ _68553_/A _68528_/B _68528_/X sky130_fd_sc_hd__and2_4
X_87362_ _88245_/CLK _87362_/D _87362_/Q sky130_fd_sc_hd__dfxtp_4
X_53754_ _53729_/A _53754_/X sky130_fd_sc_hd__buf_2
X_84574_ _84454_/CLK _84574_/D _60755_/C sky130_fd_sc_hd__dfxtp_4
X_50966_ _51021_/A _50971_/A sky130_fd_sc_hd__buf_2
X_81786_ _84980_/CLK _76154_/Y _48958_/B sky130_fd_sc_hd__dfxtp_4
X_86313_ _86312_/CLK _86313_/D _86313_/Q sky130_fd_sc_hd__dfxtp_4
X_52705_ _52701_/Y _52702_/X _52704_/X _52705_/Y sky130_fd_sc_hd__a21oi_4
X_59261_ _59135_/X _85644_/Q _59196_/X _59261_/X sky130_fd_sc_hd__o21a_4
X_83525_ _83526_/CLK _71362_/X _83525_/Q sky130_fd_sc_hd__dfxtp_4
X_56473_ _56462_/X _56016_/X _56472_/Y _56473_/Y sky130_fd_sc_hd__o21ai_4
X_68459_ _68301_/X _68446_/Y _68447_/X _68458_/Y _68459_/X sky130_fd_sc_hd__a211o_4
X_80737_ _81121_/CLK _80737_/D _80737_/Q sky130_fd_sc_hd__dfxtp_4
X_87293_ _87813_/CLK _43730_/Y _87293_/Q sky130_fd_sc_hd__dfxtp_4
X_53685_ _52166_/A _53666_/X _53692_/C _53685_/X sky130_fd_sc_hd__and3_4
X_50897_ _50952_/A _50897_/X sky130_fd_sc_hd__buf_2
X_58212_ _58191_/X _58209_/Y _58211_/Y _84907_/D sky130_fd_sc_hd__a21oi_4
X_55424_ _55297_/X _55373_/Y _57186_/B sky130_fd_sc_hd__xnor2_4
X_86244_ _85826_/CLK _86244_/D _86244_/Q sky130_fd_sc_hd__dfxtp_4
X_40650_ _40649_/Y _40650_/X sky130_fd_sc_hd__buf_2
X_52636_ _52633_/Y _52619_/X _52635_/X _85783_/D sky130_fd_sc_hd__a21oi_4
X_59192_ _59117_/A _86353_/Q _59192_/Y sky130_fd_sc_hd__nor2_4
X_71470_ _71418_/B _71479_/B sky130_fd_sc_hd__buf_2
X_83456_ _83457_/CLK _83456_/D _83456_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_402 sky130_fd_sc_hd__decap_3
X_80668_ _84531_/CLK _80668_/D _43945_/A sky130_fd_sc_hd__dfxtp_4
XPHY_413 sky130_fd_sc_hd__decap_3
XPHY_424 sky130_fd_sc_hd__decap_3
X_58143_ _58139_/Y _58142_/Y _58105_/X _58143_/X sky130_fd_sc_hd__a21o_4
X_70421_ _71012_/A _70428_/A _70854_/A _70421_/Y sky130_fd_sc_hd__nor3_4
XPHY_435 sky130_fd_sc_hd__decap_3
X_82407_ _82443_/CLK _82439_/Q _78373_/A sky130_fd_sc_hd__dfxtp_4
X_55355_ _55356_/A _55362_/A _55353_/X _55354_/Y _55369_/A sky130_fd_sc_hd__a211o_4
X_86175_ _85566_/CLK _86175_/D _86175_/Q sky130_fd_sc_hd__dfxtp_4
X_40581_ _40581_/A _40581_/X sky130_fd_sc_hd__buf_2
X_52567_ _52567_/A _46585_/Y _52567_/Y sky130_fd_sc_hd__nand2_4
XPHY_446 sky130_fd_sc_hd__decap_3
X_83387_ _84945_/CLK _83387_/D _83387_/Q sky130_fd_sc_hd__dfxtp_4
X_80599_ _80598_/X _80599_/Y sky130_fd_sc_hd__inv_2
XPHY_457 sky130_fd_sc_hd__decap_3
XPHY_468 sky130_fd_sc_hd__decap_3
X_42320_ _42276_/A _42320_/X sky130_fd_sc_hd__buf_2
X_54306_ _85466_/Q _54294_/X _54305_/Y _54306_/Y sky130_fd_sc_hd__o21ai_4
X_73140_ _73137_/X _73139_/X _73141_/B sky130_fd_sc_hd__nand2_4
XPHY_479 sky130_fd_sc_hd__decap_3
X_85126_ _85134_/CLK _85126_/D _56887_/B sky130_fd_sc_hd__dfxtp_4
X_51518_ _51514_/A _53046_/B _51518_/Y sky130_fd_sc_hd__nand2_4
X_58074_ _58017_/X _85383_/Q _58073_/X _58074_/Y sky130_fd_sc_hd__o21ai_4
X_70352_ HASH_ADDR[3] _70496_/A sky130_fd_sc_hd__inv_2
X_82338_ _82103_/CLK _77049_/X _82338_/Q sky130_fd_sc_hd__dfxtp_4
X_55286_ _56868_/A _55671_/A _56868_/B _55286_/Y sky130_fd_sc_hd__nand3_4
X_52498_ _50802_/A _52446_/B _52498_/C _52498_/X sky130_fd_sc_hd__and3_4
X_57025_ _56800_/X _57024_/Y _57025_/X sky130_fd_sc_hd__xor2_4
X_42251_ _41437_/X _42248_/X _87959_/Q _42249_/X _87959_/D sky130_fd_sc_hd__a2bb2o_4
X_54237_ _54255_/A _54237_/B _54237_/C _53070_/D _54237_/X sky130_fd_sc_hd__and4_4
X_73071_ _72963_/X _83070_/Q _73015_/X _73070_/X _73071_/X sky130_fd_sc_hd__a211o_4
X_85057_ _85057_/CLK _85057_/D _85057_/Q sky130_fd_sc_hd__dfxtp_4
X_51449_ _46612_/A _52688_/A sky130_fd_sc_hd__buf_2
X_70283_ _70247_/X _70292_/B sky130_fd_sc_hd__buf_2
X_82269_ _83514_/CLK _82269_/D _82269_/Q sky130_fd_sc_hd__dfxtp_4
X_41202_ _41184_/X _81136_/Q _41201_/X _41203_/A sky130_fd_sc_hd__o21ai_4
X_72022_ _72017_/X _53848_/B _72022_/Y sky130_fd_sc_hd__nand2_4
X_84008_ _81783_/CLK _68224_/X _84008_/Q sky130_fd_sc_hd__dfxtp_4
X_42182_ _41259_/X _42161_/X _87993_/Q _42162_/X _87993_/D sky130_fd_sc_hd__a2bb2o_4
X_54168_ _54194_/A _54184_/A sky130_fd_sc_hd__buf_2
X_53119_ _53116_/Y _53111_/X _53118_/X _85694_/D sky130_fd_sc_hd__a21oi_4
X_41133_ _41100_/X _81149_/Q _41132_/X _41133_/Y sky130_fd_sc_hd__o21ai_4
X_76830_ _76812_/X _76825_/A _76831_/A sky130_fd_sc_hd__and2_4
X_46990_ _46990_/A _52790_/D sky130_fd_sc_hd__buf_2
X_54099_ _53418_/X _54123_/A sky130_fd_sc_hd__buf_2
X_58976_ _58976_/A _58973_/B _58976_/Y sky130_fd_sc_hd__nand2_4
X_41064_ _41064_/A _41064_/X sky130_fd_sc_hd__buf_2
X_45941_ _45941_/A _59539_/A sky130_fd_sc_hd__buf_2
X_57927_ _57773_/X _85715_/Q _44177_/X _57927_/X sky130_fd_sc_hd__o21a_4
X_76761_ _76746_/A _81357_/D _76760_/X _76761_/Y sky130_fd_sc_hd__o21ai_4
X_73973_ _73972_/X _66155_/B _73973_/X sky130_fd_sc_hd__and2_4
X_85959_ _85959_/CLK _51716_/Y _85959_/Q sky130_fd_sc_hd__dfxtp_4
X_78500_ _82511_/Q _82767_/D _82479_/D sky130_fd_sc_hd__xor2_4
X_75712_ _81009_/Q _75712_/B _75712_/X sky130_fd_sc_hd__xor2_4
X_48660_ _48660_/A _48851_/B sky130_fd_sc_hd__buf_2
X_72924_ _72924_/A _72924_/B _72924_/Y sky130_fd_sc_hd__nor2_4
X_79480_ _79480_/A _79480_/Y sky130_fd_sc_hd__inv_2
X_57858_ _86648_/Q _57845_/X _57858_/Y sky130_fd_sc_hd__nor2_4
X_45872_ _45870_/Y _44968_/X _44875_/X _45871_/Y _45872_/X sky130_fd_sc_hd__a211o_4
X_76692_ _81350_/D _76692_/B _76692_/Y sky130_fd_sc_hd__nand2_4
X_47611_ _47574_/A _53148_/B _47611_/Y sky130_fd_sc_hd__nand2_4
X_78431_ _82506_/Q _82762_/D _82474_/D sky130_fd_sc_hd__xor2_4
X_44823_ _44822_/Y _86936_/D sky130_fd_sc_hd__inv_2
X_56809_ _83322_/Q _56816_/A sky130_fd_sc_hd__buf_2
X_75643_ _75629_/X _75630_/A _75643_/X sky130_fd_sc_hd__and2_4
X_87629_ _88144_/CLK _42961_/X _87629_/Q sky130_fd_sc_hd__dfxtp_4
X_48591_ _48584_/Y _48585_/X _48590_/X _86509_/D sky130_fd_sc_hd__a21oi_4
X_72855_ _72855_/A _73438_/B _72855_/Y sky130_fd_sc_hd__nor2_4
X_57789_ _57788_/X _64621_/A sky130_fd_sc_hd__buf_2
X_47542_ _47538_/Y _47509_/X _47541_/X _86624_/D sky130_fd_sc_hd__a21oi_4
X_71806_ _71779_/A _71422_/C _70852_/C _71806_/X sky130_fd_sc_hd__and3_4
X_59528_ _44216_/X _44217_/X _45941_/A _59609_/D sky130_fd_sc_hd__a21oi_4
X_78362_ _78361_/Y _78362_/Y sky130_fd_sc_hd__inv_2
X_44754_ _44618_/A _44754_/X sky130_fd_sc_hd__buf_2
X_75574_ _75574_/A _75575_/A sky130_fd_sc_hd__inv_2
X_41966_ _88089_/Q _41966_/Y sky130_fd_sc_hd__inv_2
X_72786_ _72758_/X _65444_/B _72786_/X sky130_fd_sc_hd__and2_4
X_77313_ _77312_/Y _77292_/Y _77294_/Y _77315_/C sky130_fd_sc_hd__o21ai_4
X_43705_ _43705_/A _87302_/D sky130_fd_sc_hd__inv_2
X_74525_ _70383_/X _74518_/B _70880_/C _74531_/D _74525_/Y sky130_fd_sc_hd__nand4_4
X_40917_ _40870_/X _40871_/X _40914_/X _69935_/B _40916_/X _40918_/A
+ sky130_fd_sc_hd__o32ai_4
X_47473_ _47473_/A _47474_/A sky130_fd_sc_hd__inv_2
X_71737_ _71736_/X _71737_/X sky130_fd_sc_hd__buf_2
X_59459_ _84726_/Q _59460_/A sky130_fd_sc_hd__inv_2
X_78293_ _82687_/Q _78293_/B _78293_/X sky130_fd_sc_hd__xor2_4
X_44685_ _44593_/X _44594_/X _40616_/Y _44684_/Y _44596_/X _44685_/Y
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_10_573_0_CLK clkbuf_9_286_0_CLK/X _82899_/CLK sky130_fd_sc_hd__clkbuf_1
X_41897_ _41894_/X _41879_/X _40610_/X _73675_/A _41882_/X _41897_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49212_ _49212_/A _49212_/B _49212_/Y sky130_fd_sc_hd__nand2_4
X_46424_ _82930_/Q _47991_/B sky130_fd_sc_hd__inv_2
X_77244_ _77245_/A _77245_/C _77243_/X _77244_/X sky130_fd_sc_hd__a21o_4
X_43636_ _43611_/A _43636_/X sky130_fd_sc_hd__buf_2
X_62470_ _62415_/X _62005_/A _62618_/D _62194_/D _62470_/X sky130_fd_sc_hd__and4_4
X_74456_ _74442_/X _48572_/A _74456_/Y sky130_fd_sc_hd__nand2_4
X_40848_ _40783_/X _41026_/A _40847_/X _40848_/X sky130_fd_sc_hd__o21a_4
X_71668_ _71528_/X _71289_/B _71669_/A sky130_fd_sc_hd__nor2_4
X_49143_ _83599_/Q _49144_/A sky130_fd_sc_hd__inv_2
X_61421_ _61421_/A _61404_/X _61406_/C _61390_/D _61421_/Y sky130_fd_sc_hd__nand4_4
X_73407_ _73407_/A _86504_/Q _73407_/X sky130_fd_sc_hd__and2_4
X_46355_ _83648_/Q _53985_/B sky130_fd_sc_hd__inv_2
X_70619_ _71005_/A _70724_/A sky130_fd_sc_hd__buf_2
X_77175_ _77175_/A _77173_/C _77175_/Y sky130_fd_sc_hd__nand2_4
X_43567_ _43557_/X _43563_/X _40501_/X _87357_/Q _43058_/A _43568_/A
+ sky130_fd_sc_hd__o32ai_4
X_74387_ _46623_/A _74387_/X sky130_fd_sc_hd__buf_2
X_40779_ _82878_/Q _40779_/B _40779_/X sky130_fd_sc_hd__or2_4
X_71599_ _71581_/A _83443_/Q _71598_/Y _83443_/D sky130_fd_sc_hd__a21o_4
X_45306_ _45305_/Y _45272_/X _45306_/Y sky130_fd_sc_hd__nand2_4
X_64140_ _64187_/A _64187_/B _84271_/Q _64140_/Y sky130_fd_sc_hd__nor3_4
X_76126_ _76126_/A _81724_/D _76126_/C _76126_/Y sky130_fd_sc_hd__nand3_4
X_42518_ _42518_/A _42518_/Y sky130_fd_sc_hd__inv_2
X_61352_ _61384_/A _61384_/B _84488_/Q _61352_/Y sky130_fd_sc_hd__nor3_4
X_49074_ _49056_/A _49073_/X _49074_/Y sky130_fd_sc_hd__nand2_4
X_73338_ _73328_/Y _73337_/X _73339_/B sky130_fd_sc_hd__xnor2_4
Xclkbuf_10_588_0_CLK clkbuf_9_294_0_CLK/X _81134_/CLK sky130_fd_sc_hd__clkbuf_1
X_46286_ _46262_/X _48915_/A _46285_/X _51251_/B sky130_fd_sc_hd__o21ai_4
X_43498_ _43513_/A _43498_/X sky130_fd_sc_hd__buf_2
X_48025_ _66168_/B _47998_/X _48024_/Y _48025_/Y sky130_fd_sc_hd__o21ai_4
X_60303_ _60239_/B _60189_/Y _60302_/X _60227_/A _60304_/A sky130_fd_sc_hd__nand4_4
X_45237_ _45237_/A _45237_/X sky130_fd_sc_hd__buf_2
X_64071_ _64162_/A _58452_/A _64071_/C _64071_/X sky130_fd_sc_hd__and3_4
X_76057_ _76063_/B _76063_/C _76057_/Y sky130_fd_sc_hd__nand2_4
X_42449_ _47872_/A _41902_/A _52398_/A _42449_/Y sky130_fd_sc_hd__a21oi_4
X_61283_ _61293_/B _59660_/C _59660_/D _61283_/Y sky130_fd_sc_hd__nand3_4
X_73269_ _73270_/B _73270_/C _73268_/X _73269_/X sky130_fd_sc_hd__a21o_4
X_63022_ _63022_/A _63004_/B _63004_/C _63252_/B _63022_/X sky130_fd_sc_hd__or4_4
X_75008_ _75008_/A _75008_/B _75008_/X sky130_fd_sc_hd__or2_4
X_60234_ _60288_/C _60217_/A _60235_/A sky130_fd_sc_hd__and2_4
X_45168_ _45168_/A _45169_/A sky130_fd_sc_hd__inv_2
Xclkbuf_10_511_0_CLK clkbuf_9_255_0_CLK/X _82769_/CLK sky130_fd_sc_hd__clkbuf_1
X_67830_ _81485_/D _67806_/X _67829_/X _84053_/D sky130_fd_sc_hd__a21bo_4
X_44119_ _44119_/A _86770_/Q _44119_/Y sky130_fd_sc_hd__nand2_4
X_79816_ _84227_/Q _83275_/Q _79816_/X sky130_fd_sc_hd__xor2_4
X_60165_ _60165_/A _59602_/A _60165_/X sky130_fd_sc_hd__and2_4
X_49976_ _86288_/Q _49960_/X _49975_/Y _49976_/Y sky130_fd_sc_hd__o21ai_4
X_45099_ _45092_/X _45096_/Y _45098_/Y _86899_/D sky130_fd_sc_hd__a21oi_4
X_48927_ _48623_/A _48928_/C sky130_fd_sc_hd__buf_2
X_67761_ _67997_/A _67761_/X sky130_fd_sc_hd__buf_2
X_79747_ _79731_/Y _79734_/Y _79747_/X sky130_fd_sc_hd__or2_4
X_64973_ _64601_/A _65074_/A sky130_fd_sc_hd__buf_2
X_60096_ _60058_/B _59995_/X _60095_/X _60096_/Y sky130_fd_sc_hd__a21boi_4
X_76959_ _76792_/Y _81362_/D sky130_fd_sc_hd__inv_2
X_69500_ _69575_/A _69500_/X sky130_fd_sc_hd__buf_2
X_66712_ _66664_/X _86800_/Q _66712_/X sky130_fd_sc_hd__and2_4
X_63924_ _61461_/X _63908_/B _63894_/C _63908_/D _63924_/Y sky130_fd_sc_hd__nand4_4
X_48858_ _48833_/A _48859_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_526_0_CLK clkbuf_9_263_0_CLK/X _81532_/CLK sky130_fd_sc_hd__clkbuf_1
X_79678_ _65142_/C _72357_/Y _79677_/Y _79678_/X sky130_fd_sc_hd__o21a_4
X_67692_ _87908_/Q _67591_/X _67641_/X _67691_/X _67692_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_6_17_0_CLK clkbuf_5_8_0_CLK/X clkbuf_7_35_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_69431_ _69309_/A _69431_/B _69431_/X sky130_fd_sc_hd__and2_4
X_47809_ _47809_/A _53255_/B sky130_fd_sc_hd__buf_2
X_78629_ _78630_/A _82692_/Q _78632_/B sky130_fd_sc_hd__nor2_4
X_66643_ _66540_/A _66643_/X sky130_fd_sc_hd__buf_2
X_63855_ _63448_/B _63900_/B _63900_/C _63820_/D _63859_/B sky130_fd_sc_hd__nand4_4
X_48789_ _86482_/Q _48781_/X _48788_/Y _48789_/Y sky130_fd_sc_hd__o21ai_4
X_50820_ _50819_/X _50820_/X sky130_fd_sc_hd__buf_2
X_62806_ _62792_/X _62839_/B _62806_/C _62806_/Y sky130_fd_sc_hd__nor3_4
X_81640_ _81250_/CLK _76847_/A _81640_/Q sky130_fd_sc_hd__dfxtp_4
X_69362_ _69128_/X _69362_/B _69362_/X sky130_fd_sc_hd__and2_4
X_66574_ _69779_/A _66574_/X sky130_fd_sc_hd__buf_2
X_63786_ _64191_/D _63787_/D sky130_fd_sc_hd__buf_2
X_60998_ _64182_/C _60998_/X sky130_fd_sc_hd__buf_2
X_68313_ _68272_/X _67911_/Y _68308_/X _68312_/Y _68313_/X sky130_fd_sc_hd__a211o_4
X_65525_ _65416_/X _65525_/B _65525_/X sky130_fd_sc_hd__and2_4
X_50751_ _51256_/A _50751_/B _50751_/C _50751_/X sky130_fd_sc_hd__and3_4
X_62737_ _62737_/A _62737_/X sky130_fd_sc_hd__buf_2
X_81571_ _81587_/CLK _84171_/Q _76665_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_2_2_0_CLK clkbuf_2_3_0_CLK/A clkbuf_2_2_1_CLK/A sky130_fd_sc_hd__clkbuf_1
X_69293_ _69290_/X _69292_/X _69293_/Y sky130_fd_sc_hd__nand2_4
X_83310_ _83310_/CLK _71975_/Y _83310_/Q sky130_fd_sc_hd__dfxtp_4
X_80522_ _80530_/A _80522_/B _80522_/Y sky130_fd_sc_hd__xnor2_4
X_68244_ _68221_/X _67506_/Y _68228_/X _68243_/Y _68244_/X sky130_fd_sc_hd__a211o_4
X_53470_ _43177_/Y _53798_/A sky130_fd_sc_hd__buf_2
X_65456_ _65453_/X _85599_/Q _65326_/X _65455_/X _65456_/X sky130_fd_sc_hd__a211o_4
X_84290_ _84287_/CLK _84290_/D _63864_/C sky130_fd_sc_hd__dfxtp_4
X_50682_ _50682_/A _50169_/B _50682_/Y sky130_fd_sc_hd__nand2_4
X_62668_ _62667_/X _62927_/A sky130_fd_sc_hd__buf_2
X_52421_ _52419_/Y _52415_/X _52420_/X _85826_/D sky130_fd_sc_hd__a21oi_4
X_64407_ _64399_/Y _64406_/X _64386_/X _64407_/X sky130_fd_sc_hd__o21a_4
X_83241_ _84333_/CLK _72513_/Y _79513_/B sky130_fd_sc_hd__dfxtp_4
X_61619_ _61608_/X _61618_/X _61619_/C _61619_/Y sky130_fd_sc_hd__nand3_4
X_80453_ _59204_/Y _66164_/C _80452_/Y _80457_/A sky130_fd_sc_hd__o21a_4
X_68175_ _68155_/X _67078_/Y _68168_/X _68174_/Y _68175_/X sky130_fd_sc_hd__a211o_4
X_65387_ _65387_/A _86243_/Q _65387_/X sky130_fd_sc_hd__and2_4
X_62599_ _61665_/B _62504_/X _62534_/X _62621_/D _62600_/D sky130_fd_sc_hd__nand4_4
X_55140_ _55140_/A _55140_/X sky130_fd_sc_hd__buf_2
X_67126_ _68742_/A _67126_/X sky130_fd_sc_hd__buf_2
X_52352_ _52350_/Y _52340_/X _52351_/X _85840_/D sky130_fd_sc_hd__a21oi_4
X_83172_ _84980_/CLK _83172_/D _83172_/Q sky130_fd_sc_hd__dfxtp_4
X_64338_ _64332_/X _64334_/X _64335_/X _64337_/Y _64326_/X _64338_/X
+ sky130_fd_sc_hd__o41a_4
X_80384_ _80361_/A _80382_/X _80361_/B _80384_/D _80384_/Y sky130_fd_sc_hd__nand4_4
X_51303_ _51301_/Y _51289_/X _51302_/X _51303_/Y sky130_fd_sc_hd__a21oi_4
X_82123_ _82532_/CLK _77812_/X _82123_/Q sky130_fd_sc_hd__dfxtp_4
X_55071_ _55068_/Y _55050_/X _55070_/X _85324_/D sky130_fd_sc_hd__a21oi_4
X_67057_ _67057_/A _87615_/Q _67057_/X sky130_fd_sc_hd__and2_4
X_52283_ _52293_/A _48922_/B _52283_/Y sky130_fd_sc_hd__nand2_4
X_64269_ _64328_/A _64269_/X sky130_fd_sc_hd__buf_2
X_87980_ _88158_/CLK _87980_/D _87980_/Q sky130_fd_sc_hd__dfxtp_4
X_54022_ _53998_/A _50808_/B _54022_/Y sky130_fd_sc_hd__nand2_4
X_66008_ _65934_/X _66008_/B _66008_/X sky130_fd_sc_hd__and2_4
X_51234_ _51286_/A _51240_/A sky130_fd_sc_hd__buf_2
X_86931_ _87653_/CLK _86931_/D _67629_/B sky130_fd_sc_hd__dfxtp_4
X_82054_ _84020_/CLK _84014_/Q _77771_/B sky130_fd_sc_hd__dfxtp_4
X_81005_ _84210_/CLK _84213_/Q _81005_/Q sky130_fd_sc_hd__dfxtp_4
X_58830_ _58872_/A _58830_/B _58830_/Y sky130_fd_sc_hd__nor2_4
X_51165_ _51177_/A _51160_/B _51141_/X _52857_/D _51165_/X sky130_fd_sc_hd__and4_4
X_86862_ _80657_/CLK _45671_/Y _63206_/B sky130_fd_sc_hd__dfxtp_4
X_50116_ _64931_/B _50113_/X _50115_/Y _50116_/Y sky130_fd_sc_hd__o21ai_4
X_85813_ _85527_/CLK _52483_/Y _85813_/Q sky130_fd_sc_hd__dfxtp_4
X_58761_ _58939_/A _58761_/X sky130_fd_sc_hd__buf_2
X_51096_ _51092_/Y _51093_/X _51095_/X _86075_/D sky130_fd_sc_hd__a21oi_4
X_55973_ _74545_/C _55690_/X _44102_/X _55972_/X _55974_/B sky130_fd_sc_hd__a211o_4
X_67959_ _68025_/A _88217_/Q _67959_/X sky130_fd_sc_hd__and2_4
X_86793_ _87077_/CLK _46052_/X _86793_/Q sky130_fd_sc_hd__dfxtp_4
X_57712_ _57711_/X _57712_/X sky130_fd_sc_hd__buf_2
X_50047_ _50043_/Y _50029_/X _50046_/X _50047_/Y sky130_fd_sc_hd__a21oi_4
X_54924_ _54919_/X _47762_/Y _54924_/Y sky130_fd_sc_hd__nand2_4
X_85744_ _85748_/CLK _52847_/Y _85744_/Q sky130_fd_sc_hd__dfxtp_4
X_82956_ _82956_/CLK _82956_/D _82956_/Q sky130_fd_sc_hd__dfxtp_4
X_70970_ _50781_/B _70961_/X _70969_/Y _83646_/D sky130_fd_sc_hd__o21ai_4
X_58692_ _58682_/X _85783_/Q _58594_/X _58692_/X sky130_fd_sc_hd__o21a_4
X_57643_ _84963_/Q _57635_/X _57642_/Y _57643_/Y sky130_fd_sc_hd__o21ai_4
X_81907_ _82131_/CLK _81907_/D _82283_/D sky130_fd_sc_hd__dfxtp_4
X_69629_ _69625_/X _69628_/X _69389_/X _69629_/Y sky130_fd_sc_hd__a21oi_4
X_54855_ _85365_/Q _54839_/X _54854_/Y _54855_/Y sky130_fd_sc_hd__o21ai_4
X_85675_ _86400_/CLK _53218_/Y _85675_/Q sky130_fd_sc_hd__dfxtp_4
X_82887_ _82317_/CLK _78112_/B _82887_/Q sky130_fd_sc_hd__dfxtp_4
X_87414_ _87926_/CLK _43454_/Y _87414_/Q sky130_fd_sc_hd__dfxtp_4
X_41820_ _41819_/Y _88136_/D sky130_fd_sc_hd__inv_2
X_53806_ _48928_/A _53806_/B _53806_/C _53806_/X sky130_fd_sc_hd__and3_4
X_72640_ _70178_/C _72631_/X _72639_/Y _83207_/D sky130_fd_sc_hd__a21bo_4
X_84626_ _84623_/CLK _60347_/Y _60346_/C sky130_fd_sc_hd__dfxtp_4
X_57574_ _57552_/X _48014_/Y _57574_/Y sky130_fd_sc_hd__nand2_4
X_81838_ _81883_/CLK _81870_/Q _77406_/A sky130_fd_sc_hd__dfxtp_4
X_88394_ _88394_/CLK _88394_/D _88394_/Q sky130_fd_sc_hd__dfxtp_4
X_54786_ _54790_/A _47516_/A _54786_/Y sky130_fd_sc_hd__nand2_4
X_51998_ _66082_/B _51994_/X _51997_/Y _51998_/Y sky130_fd_sc_hd__o21ai_4
X_59313_ _59286_/X _86056_/Q _59312_/X _59313_/Y sky130_fd_sc_hd__o21ai_4
X_56525_ _56525_/A _56533_/A sky130_fd_sc_hd__buf_2
X_87345_ _87345_/CLK _43601_/Y _87345_/Q sky130_fd_sc_hd__dfxtp_4
X_41751_ _41814_/A _41751_/X sky130_fd_sc_hd__buf_2
X_53737_ _85578_/Q _53729_/X _53736_/Y _53737_/Y sky130_fd_sc_hd__o21ai_4
X_72571_ _79405_/B _61252_/X _72569_/Y _72570_/Y _83231_/D sky130_fd_sc_hd__o22a_4
X_84557_ _84562_/CLK _84557_/D _60826_/C sky130_fd_sc_hd__dfxtp_4
X_50949_ _50944_/Y _50928_/X _50948_/X _50949_/Y sky130_fd_sc_hd__a21oi_4
X_81769_ _82896_/CLK _76025_/X _81769_/Q sky130_fd_sc_hd__dfxtp_4
X_74310_ _74302_/X _74310_/B _74310_/C _74310_/Y sky130_fd_sc_hd__nand3_4
X_40702_ _40702_/A _40702_/X sky130_fd_sc_hd__buf_2
X_59244_ _59117_/A _59244_/B _59244_/Y sky130_fd_sc_hd__nor2_4
X_71522_ _51728_/B _71512_/A _71521_/Y _83468_/D sky130_fd_sc_hd__o21ai_4
X_83508_ _83508_/CLK _71412_/X _83508_/Q sky130_fd_sc_hd__dfxtp_4
X_44470_ _41168_/Y _44464_/X _87092_/Q _44466_/X _44470_/X sky130_fd_sc_hd__a2bb2o_4
X_56456_ _56456_/A _57364_/D sky130_fd_sc_hd__buf_2
X_75290_ _75289_/Y _75291_/C sky130_fd_sc_hd__inv_2
X_41682_ _41799_/A _41682_/X sky130_fd_sc_hd__buf_2
X_87276_ _88056_/CLK _43766_/Y _69236_/B sky130_fd_sc_hd__dfxtp_4
X_53668_ _53664_/Y _53653_/X _53667_/X _53668_/Y sky130_fd_sc_hd__a21oi_4
X_84488_ _84487_/CLK _84488_/D _84488_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_210 sky130_fd_sc_hd__decap_3
X_43421_ _40362_/X _43518_/A sky130_fd_sc_hd__buf_2
X_55407_ _55405_/X _55408_/B sky130_fd_sc_hd__inv_2
X_74241_ _74241_/A _74241_/B _74241_/Y sky130_fd_sc_hd__xnor2_4
X_86227_ _86578_/CLK _86227_/D _86227_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_221 sky130_fd_sc_hd__decap_3
X_52619_ _52619_/A _52619_/X sky130_fd_sc_hd__buf_2
X_40633_ _40632_/Y _40633_/X sky130_fd_sc_hd__buf_2
X_71453_ _71445_/X _83494_/Q _71452_/Y _71453_/X sky130_fd_sc_hd__a21o_4
X_59175_ _59135_/X _85651_/Q _59070_/X _59175_/X sky130_fd_sc_hd__o21a_4
X_83439_ _83402_/CLK _71613_/X _83439_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_232 sky130_fd_sc_hd__decap_3
X_56387_ _56020_/X _56378_/X _56386_/Y _56387_/Y sky130_fd_sc_hd__o21ai_4
X_53599_ _53604_/A _52079_/B _53599_/Y sky130_fd_sc_hd__nand2_4
XPHY_243 sky130_fd_sc_hd__decap_3
XPHY_254 sky130_fd_sc_hd__decap_3
X_70404_ DATA_TO_HASH[0] _71090_/A sky130_fd_sc_hd__buf_2
X_46140_ _46195_/A _46135_/Y _57657_/B _46139_/Y _46140_/X sky130_fd_sc_hd__a211o_4
X_58126_ _58126_/A _58126_/X sky130_fd_sc_hd__buf_2
XPHY_265 sky130_fd_sc_hd__decap_3
X_43352_ _43352_/A _87465_/D sky130_fd_sc_hd__inv_2
X_55338_ _82992_/Q _44061_/X _55312_/X _55337_/X _55365_/B sky130_fd_sc_hd__a211o_4
X_74172_ _74232_/A _66283_/B _74172_/X sky130_fd_sc_hd__and2_4
X_86158_ _85555_/CLK _86158_/D _86158_/Q sky130_fd_sc_hd__dfxtp_4
X_40564_ _40563_/X _48162_/A sky130_fd_sc_hd__buf_2
XPHY_276 sky130_fd_sc_hd__decap_3
X_71384_ _71373_/X _83518_/Q _71383_/Y _71384_/X sky130_fd_sc_hd__a21o_4
XPHY_287 sky130_fd_sc_hd__decap_3
XPHY_298 sky130_fd_sc_hd__decap_3
X_42303_ _42290_/A _42303_/X sky130_fd_sc_hd__buf_2
X_73123_ _83164_/Q _73079_/X _73122_/X _73123_/X sky130_fd_sc_hd__a21o_4
X_85109_ _85074_/CLK _85109_/D _45582_/A sky130_fd_sc_hd__dfxtp_4
X_46071_ _41580_/A _46061_/X _67123_/B _46062_/X _86783_/D sky130_fd_sc_hd__a2bb2o_4
X_58057_ _58048_/Y _57981_/X _58053_/X _58056_/X _84929_/D sky130_fd_sc_hd__a22oi_4
X_70335_ _70338_/A _70333_/B _83089_/Q _70332_/X _70335_/X sky130_fd_sc_hd__and4_4
X_55269_ _55276_/A _57210_/B _55269_/X sky130_fd_sc_hd__and2_4
X_43283_ _41151_/X _43277_/X _87500_/Q _43278_/X _87500_/D sky130_fd_sc_hd__a2bb2o_4
X_78980_ _78968_/A _78967_/Y _78979_/X _78981_/B sky130_fd_sc_hd__o21ai_4
X_86089_ _86089_/CLK _86089_/D _86089_/Q sky130_fd_sc_hd__dfxtp_4
X_40495_ _40416_/A _81164_/Q _40495_/X sky130_fd_sc_hd__or2_4
X_57008_ _56991_/Y _57024_/D sky130_fd_sc_hd__buf_2
X_45022_ _64294_/B _61417_/B sky130_fd_sc_hd__buf_2
X_42234_ _42231_/X _42226_/X _41387_/X _87968_/Q _42228_/X _42234_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77931_ _77920_/A _77919_/Y _77930_/X _77931_/Y sky130_fd_sc_hd__a21oi_4
X_73054_ _42011_/Y _72921_/X _72944_/X _73053_/Y _73054_/X sky130_fd_sc_hd__a211o_4
X_70266_ _70255_/X _74720_/B _70265_/X _70266_/X sky130_fd_sc_hd__a21o_4
X_72005_ _48978_/A _71959_/X _71964_/X _72005_/X sky130_fd_sc_hd__and3_4
X_49830_ _49830_/A _49830_/B _49830_/C _53044_/D _49830_/X sky130_fd_sc_hd__and4_4
X_42165_ _42154_/X _42141_/X _41209_/X _88001_/Q _42142_/X _42166_/A
+ sky130_fd_sc_hd__o32ai_4
X_77862_ _82160_/Q _77862_/B _82128_/D sky130_fd_sc_hd__xor2_4
X_70197_ _70195_/X _83841_/Q _70196_/X _70197_/X sky130_fd_sc_hd__a21o_4
X_79601_ _79605_/A _79605_/B _79601_/X sky130_fd_sc_hd__xor2_4
X_41116_ _41115_/X _41116_/X sky130_fd_sc_hd__buf_2
X_76813_ _76812_/X _76818_/A sky130_fd_sc_hd__inv_2
X_49761_ _49779_/A _49750_/X _49761_/C _52977_/D _49761_/X sky130_fd_sc_hd__and4_4
X_46973_ _46981_/A _46944_/B _46981_/C _52779_/D _46973_/X sky130_fd_sc_hd__and4_4
X_58959_ _58603_/A _58959_/X sky130_fd_sc_hd__buf_2
X_42096_ _42096_/A _42096_/X sky130_fd_sc_hd__buf_2
X_77793_ _82058_/Q _77809_/A sky130_fd_sc_hd__inv_2
X_48712_ _48707_/Y _48403_/X _48711_/Y _48712_/Y sky130_fd_sc_hd__a21boi_4
X_79532_ _65421_/C _83250_/Q _79532_/Y sky130_fd_sc_hd__nand2_4
X_45924_ _45924_/A _65034_/A sky130_fd_sc_hd__buf_2
X_41047_ _41047_/A _88288_/D sky130_fd_sc_hd__inv_2
X_76744_ _76744_/A _76743_/Y _76745_/B sky130_fd_sc_hd__xor2_4
X_49692_ _49685_/A _49669_/B _49685_/C _51214_/D _49692_/X sky130_fd_sc_hd__and4_4
X_61970_ _61747_/X _61971_/D sky130_fd_sc_hd__buf_2
X_73956_ _73956_/A _73955_/X _73957_/B sky130_fd_sc_hd__nand2_4
X_48643_ _48606_/X _49139_/B _48642_/Y _48644_/A sky130_fd_sc_hd__o21ai_4
X_60921_ _63761_/A _60921_/X sky130_fd_sc_hd__buf_2
X_72907_ _72870_/X _86204_/Q _72905_/X _72906_/X _72907_/X sky130_fd_sc_hd__a211o_4
X_79463_ _79481_/A _79462_/Y _82844_/D sky130_fd_sc_hd__xor2_4
X_45855_ _55221_/B _45394_/X _45571_/X _45854_/Y _45855_/X sky130_fd_sc_hd__a211o_4
X_76675_ _76675_/A _76674_/X _81540_/D sky130_fd_sc_hd__xor2_4
X_73887_ _73888_/B _73888_/C _73886_/X _73887_/X sky130_fd_sc_hd__a21o_4
X_78414_ _78400_/B _78426_/C _78426_/B _78414_/Y sky130_fd_sc_hd__a21boi_4
X_44806_ _40554_/X _45980_/A sky130_fd_sc_hd__buf_2
X_63640_ _58277_/A _60748_/X _60724_/A _62544_/Y _60671_/B _63640_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75626_ _75620_/Y _75621_/X _75625_/Y _75632_/B sky130_fd_sc_hd__a21oi_4
X_60852_ _60406_/B _60174_/D _61075_/B _60852_/X sky130_fd_sc_hd__and3_4
X_48574_ _86510_/Q _48536_/X _48573_/Y _48574_/Y sky130_fd_sc_hd__o21ai_4
X_72838_ _72838_/A _73092_/A sky130_fd_sc_hd__buf_2
X_79394_ _79394_/A _79394_/B _79395_/B sky130_fd_sc_hd__xor2_4
X_45786_ _82984_/Q _45787_/A sky130_fd_sc_hd__inv_2
X_42998_ _42998_/A _87613_/D sky130_fd_sc_hd__inv_2
X_47525_ _47525_/A _47553_/A sky130_fd_sc_hd__buf_2
X_78345_ _78343_/Y _78344_/Y _82789_/Q _78345_/X sky130_fd_sc_hd__a21o_4
X_44737_ _49210_/A _50731_/B _40733_/Y _44735_/Y _44736_/X _44737_/Y
+ sky130_fd_sc_hd__o32ai_4
X_63571_ _63523_/A _61997_/X _63571_/X sky130_fd_sc_hd__and2_4
X_75557_ _81089_/Q _75557_/B _75557_/X sky130_fd_sc_hd__xor2_4
X_41949_ _41932_/X _41927_/X _40702_/X _74031_/A _41928_/X _41950_/A
+ sky130_fd_sc_hd__o32ai_4
X_60783_ _63400_/C _63384_/C sky130_fd_sc_hd__buf_2
X_72769_ _72769_/A _72769_/B _72769_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_4_7_1_CLK clkbuf_4_7_0_CLK/X clkbuf_4_7_1_CLK/X sky130_fd_sc_hd__clkbuf_1
X_65310_ _57770_/A _65310_/B _65310_/X sky130_fd_sc_hd__and2_4
X_62522_ _62288_/X _62522_/B _64458_/B _62609_/D _62522_/X sky130_fd_sc_hd__and4_4
X_74508_ _83051_/Q _46250_/X _74507_/Y _74508_/Y sky130_fd_sc_hd__o21ai_4
X_47456_ _47437_/X _47415_/X _47466_/C _53058_/D _47456_/X sky130_fd_sc_hd__and4_4
X_66290_ _66287_/X _66385_/B _66289_/X _66290_/Y sky130_fd_sc_hd__nand3_4
X_78276_ _78268_/Y _78262_/X _78275_/Y _78276_/Y sky130_fd_sc_hd__a21boi_4
X_44668_ _41107_/Y _44665_/X _87008_/Q _44666_/X _44668_/X sky130_fd_sc_hd__a2bb2o_4
X_75488_ _75487_/Y _75506_/D _75488_/Y sky130_fd_sc_hd__nand2_4
X_46407_ _46407_/A _46407_/X sky130_fd_sc_hd__buf_2
X_65241_ _65178_/X _86729_/Q _65239_/X _65240_/X _65241_/X sky130_fd_sc_hd__a211o_4
X_77227_ _77223_/A _77222_/Y _77227_/C _77230_/C sky130_fd_sc_hd__nand3_4
X_43619_ _40633_/X _43604_/X _73752_/A _43607_/X _43619_/X sky130_fd_sc_hd__a2bb2o_4
X_74439_ _48533_/A _46620_/A _46428_/C _74439_/Y sky130_fd_sc_hd__nand3_4
X_62453_ _61521_/B _62390_/X _62436_/X _62407_/X _62452_/X _62453_/X
+ sky130_fd_sc_hd__a41o_4
X_47387_ _47404_/A _53017_/B _47387_/Y sky130_fd_sc_hd__nand2_4
X_44599_ _44593_/X _44594_/X _40924_/Y _44598_/Y _44596_/X _44599_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49126_ _49117_/A _49125_/X _49126_/Y sky130_fd_sc_hd__nand2_4
X_61404_ _72550_/A _61404_/X sky130_fd_sc_hd__buf_2
X_46338_ _46262_/X _48959_/A _46337_/X _46339_/A sky130_fd_sc_hd__o21ai_4
X_65172_ _64817_/A _65172_/X sky130_fd_sc_hd__buf_2
X_77158_ _77149_/Y _77156_/Y _77157_/Y _77159_/B sky130_fd_sc_hd__o21a_4
X_62384_ _62218_/A _62565_/C sky130_fd_sc_hd__buf_2
X_64123_ _58187_/X _64158_/B _64158_/C _64045_/X _64123_/Y sky130_fd_sc_hd__nand4_4
X_76109_ _81723_/D _76109_/B _76109_/Y sky130_fd_sc_hd__nor2_4
X_49057_ _65066_/B _49052_/X _49056_/Y _49057_/Y sky130_fd_sc_hd__o21ai_4
X_61335_ _72550_/A _61367_/B sky130_fd_sc_hd__buf_2
X_46269_ _46257_/Y _46258_/X _46268_/Y _86752_/D sky130_fd_sc_hd__a21boi_4
X_69980_ _83881_/Q _69955_/X _69979_/X _69980_/X sky130_fd_sc_hd__a21bo_4
X_77089_ _82094_/Q _77089_/B _77089_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_10_450_0_CLK clkbuf_9_225_0_CLK/X _83707_/CLK sky130_fd_sc_hd__clkbuf_1
X_48008_ _82353_/Q _48542_/B sky130_fd_sc_hd__inv_2
X_64054_ _64047_/X _64048_/X _64050_/Y _64052_/Y _64053_/X _64054_/X
+ sky130_fd_sc_hd__a41o_4
X_68931_ _69021_/A _74097_/A _68931_/X sky130_fd_sc_hd__and2_4
X_61266_ _61194_/X _61182_/X _61202_/B _61264_/Y _61265_/X _61266_/X
+ sky130_fd_sc_hd__o41a_4
X_63005_ _62997_/X _62998_/Y _63000_/X _63003_/Y _63004_/X _63005_/Y
+ sky130_fd_sc_hd__o41ai_4
X_60217_ _60217_/A _60221_/A sky130_fd_sc_hd__buf_2
X_68862_ _74033_/A _68493_/X _68494_/X _68861_/Y _68862_/X sky130_fd_sc_hd__a211o_4
X_61197_ _64377_/A _64545_/A sky130_fd_sc_hd__buf_2
X_67813_ _67790_/A _67813_/B _67813_/X sky130_fd_sc_hd__and2_4
X_60148_ _72527_/A _72527_/B _60148_/C _60148_/Y sky130_fd_sc_hd__nand3_4
X_49959_ _49956_/Y _49951_/X _49958_/X _49959_/Y sky130_fd_sc_hd__a21oi_4
X_68793_ _68770_/X _68793_/B _68793_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_465_0_CLK clkbuf_9_232_0_CLK/X _83660_/CLK sky130_fd_sc_hd__clkbuf_1
X_82810_ _82743_/CLK _82842_/Q _82810_/Q sky130_fd_sc_hd__dfxtp_4
X_67744_ _67790_/A _88162_/Q _67744_/X sky130_fd_sc_hd__and2_4
X_52970_ _85721_/Q _52957_/X _52969_/Y _52970_/Y sky130_fd_sc_hd__o21ai_4
X_64956_ _64803_/A _65002_/A sky130_fd_sc_hd__buf_2
X_60079_ _59938_/Y _60079_/B _60027_/X _60079_/Y sky130_fd_sc_hd__nand3_4
X_83790_ _81259_/CLK _83790_/D _74780_/A sky130_fd_sc_hd__dfxtp_4
X_51921_ _52398_/A _52322_/A sky130_fd_sc_hd__buf_2
X_63907_ _63761_/A _63908_/D sky130_fd_sc_hd__buf_2
X_82741_ _82152_/CLK _84125_/Q _82741_/Q sky130_fd_sc_hd__dfxtp_4
X_67675_ _67675_/A _67675_/B _67675_/X sky130_fd_sc_hd__and2_4
X_64887_ _64835_/X _83303_/Q _44171_/X _64886_/X _64887_/X sky130_fd_sc_hd__a211o_4
X_69414_ _68394_/A _69414_/X sky130_fd_sc_hd__buf_2
X_54640_ _54637_/Y _54638_/X _54639_/X _85405_/D sky130_fd_sc_hd__a21oi_4
X_66626_ _66651_/A _66626_/B _66626_/X sky130_fd_sc_hd__and2_4
X_85460_ _85459_/CLK _85460_/D _85460_/Q sky130_fd_sc_hd__dfxtp_4
X_51852_ _51849_/Y _51850_/X _51851_/X _51852_/Y sky130_fd_sc_hd__a21oi_4
X_82672_ _82923_/CLK _82672_/D _78182_/A sky130_fd_sc_hd__dfxtp_4
X_63838_ _59501_/X _63820_/B _63900_/C _63820_/D _63838_/Y sky130_fd_sc_hd__nand4_4
X_84411_ _84409_/CLK _84411_/D _62426_/C sky130_fd_sc_hd__dfxtp_4
X_50803_ _50800_/Y _50801_/X _50802_/X _50803_/Y sky130_fd_sc_hd__a21oi_4
X_81623_ _81304_/CLK _76469_/B _81815_/D sky130_fd_sc_hd__dfxtp_4
X_69345_ _87524_/Q _69205_/X _69343_/X _69344_/X _69345_/X sky130_fd_sc_hd__a211o_4
X_54571_ _54565_/A _54559_/B _54565_/C _54571_/D _54571_/X sky130_fd_sc_hd__and4_4
X_66557_ _69853_/A _88211_/Q _66557_/X sky130_fd_sc_hd__and2_4
X_85391_ _85489_/CLK _54717_/Y _85391_/Q sky130_fd_sc_hd__dfxtp_4
X_51783_ _51780_/Y _51767_/X _51782_/X _85947_/D sky130_fd_sc_hd__a21oi_4
X_63769_ _63800_/A _63800_/B _80241_/B _63769_/Y sky130_fd_sc_hd__nor3_4
X_56310_ _56284_/X _56050_/X _56309_/Y _56310_/Y sky130_fd_sc_hd__o21ai_4
X_87130_ _87950_/CLK _87130_/D _87130_/Q sky130_fd_sc_hd__dfxtp_4
X_53522_ _53509_/A _47967_/Y _53522_/Y sky130_fd_sc_hd__nand2_4
X_65508_ _64834_/A _65663_/B sky130_fd_sc_hd__buf_2
X_84342_ _84877_/CLK _84342_/D _79310_/A sky130_fd_sc_hd__dfxtp_4
X_50734_ _86144_/Q _50706_/X _50733_/Y _50734_/Y sky130_fd_sc_hd__o21ai_4
X_81554_ _84087_/CLK _76802_/X _76200_/B sky130_fd_sc_hd__dfxtp_4
X_57290_ _57290_/A _57023_/X _57149_/C _57149_/D _57290_/X sky130_fd_sc_hd__and4_4
X_69276_ _69272_/X _69275_/X _69251_/X _69276_/X sky130_fd_sc_hd__a21o_4
X_66488_ _66475_/X _66258_/Y _66487_/Y _66488_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_403_0_CLK clkbuf_9_201_0_CLK/X _85378_/CLK sky130_fd_sc_hd__clkbuf_1
X_80505_ _84766_/Q _84158_/Q _80505_/X sky130_fd_sc_hd__xor2_4
X_56241_ _56103_/X _56225_/X _56240_/Y _85263_/D sky130_fd_sc_hd__o21ai_4
X_68227_ _84007_/Q _68220_/X _68226_/X _68227_/X sky130_fd_sc_hd__a21bo_4
X_87061_ _88108_/CLK _44542_/Y _73024_/A sky130_fd_sc_hd__dfxtp_4
X_53453_ _53460_/A _73591_/A _53453_/Y sky130_fd_sc_hd__nand2_4
X_65439_ _65184_/A _65439_/B _65439_/X sky130_fd_sc_hd__and2_4
X_84273_ _84273_/CLK _84273_/D _79998_/B sky130_fd_sc_hd__dfxtp_4
X_50665_ _50663_/Y _50644_/X _50664_/Y _86158_/D sky130_fd_sc_hd__a21boi_4
X_81485_ _81428_/CLK _81485_/D _76746_/A sky130_fd_sc_hd__dfxtp_4
X_86012_ _85725_/CLK _86012_/D _86012_/Q sky130_fd_sc_hd__dfxtp_4
X_52404_ _52402_/Y _52390_/X _52403_/X _52404_/Y sky130_fd_sc_hd__a21oi_4
X_83224_ _84487_/CLK _72594_/Y _79330_/B sky130_fd_sc_hd__dfxtp_4
X_56172_ _56172_/A _56175_/A sky130_fd_sc_hd__inv_2
X_80436_ _80436_/A _80436_/B _80436_/X sky130_fd_sc_hd__or2_4
X_68158_ _84024_/Q _68140_/X _68157_/X _84024_/D sky130_fd_sc_hd__a21bo_4
X_53384_ _53371_/A _53388_/B _53388_/C _52867_/D _53384_/X sky130_fd_sc_hd__and4_4
X_50596_ _50596_/A _50597_/A sky130_fd_sc_hd__buf_2
X_55123_ _73195_/A _73124_/B sky130_fd_sc_hd__buf_2
X_67109_ _67105_/X _67108_/X _67085_/X _67109_/X sky130_fd_sc_hd__a21o_4
X_52335_ _85843_/Q _52324_/X _52334_/Y _52335_/Y sky130_fd_sc_hd__o21ai_4
X_83155_ _86535_/CLK _83155_/D _83155_/Q sky130_fd_sc_hd__dfxtp_4
X_80367_ _84752_/Q _84144_/Q _80367_/Y sky130_fd_sc_hd__nand2_4
X_68089_ _68089_/A _68089_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_418_0_CLK clkbuf_9_209_0_CLK/X _82248_/CLK sky130_fd_sc_hd__clkbuf_1
X_70120_ _83514_/Q _83162_/Q _83502_/Q _83150_/Q _70127_/C sky130_fd_sc_hd__a22oi_4
X_82106_ _82343_/CLK _82118_/Q _82106_/Q sky130_fd_sc_hd__dfxtp_4
X_55054_ _55054_/A _54885_/B _55054_/Y sky130_fd_sc_hd__nand2_4
X_59931_ _59931_/A _59931_/X sky130_fd_sc_hd__buf_2
X_52266_ _85856_/Q _52239_/X _52265_/Y _52266_/Y sky130_fd_sc_hd__o21ai_4
X_87963_ _87195_/CLK _87963_/D _87963_/Q sky130_fd_sc_hd__dfxtp_4
X_83086_ _81603_/CLK _83086_/D _83086_/Q sky130_fd_sc_hd__dfxtp_4
X_80298_ _80298_/A _80292_/A _80292_/B _80299_/B sky130_fd_sc_hd__nand3_4
X_54005_ _85524_/Q _53989_/X _54004_/Y _54005_/Y sky130_fd_sc_hd__o21ai_4
X_51217_ _86052_/Q _51209_/X _51216_/Y _51217_/Y sky130_fd_sc_hd__o21ai_4
X_70051_ _82543_/D _70048_/X _70050_/X _70051_/X sky130_fd_sc_hd__a21bo_4
X_86914_ _86914_/CLK _44862_/X _68020_/B sky130_fd_sc_hd__dfxtp_4
X_82037_ _82008_/CLK _82037_/D _82005_/D sky130_fd_sc_hd__dfxtp_4
X_59862_ _59836_/D _59733_/Y _59680_/Y _59862_/X sky130_fd_sc_hd__o21a_4
X_52197_ _85870_/Q _52178_/X _52196_/Y _52197_/Y sky130_fd_sc_hd__o21ai_4
X_87894_ _87382_/CLK _87894_/D _87894_/Q sky130_fd_sc_hd__dfxtp_4
X_58813_ _58813_/A _58813_/X sky130_fd_sc_hd__buf_2
X_51148_ _51012_/A _51149_/A sky130_fd_sc_hd__buf_2
X_86845_ _81117_/CLK _45907_/Y _40350_/A sky130_fd_sc_hd__dfxtp_4
X_59793_ _59680_/A _59731_/Y _59754_/D _59794_/A sky130_fd_sc_hd__nand3_4
Xclkbuf_8_92_0_CLK clkbuf_8_93_0_CLK/A clkbuf_8_92_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_73810_ _73742_/A _86551_/Q _73810_/X sky130_fd_sc_hd__and2_4
X_58744_ _58667_/X _86099_/Q _58743_/X _58744_/Y sky130_fd_sc_hd__o21ai_4
X_43970_ _43970_/A _59571_/C sky130_fd_sc_hd__buf_2
X_51079_ _51077_/Y _51065_/X _51078_/X _86078_/D sky130_fd_sc_hd__a21oi_4
X_55956_ _55956_/A _55956_/B _74297_/C _56003_/B _55957_/A sky130_fd_sc_hd__and4_4
X_74790_ _74764_/A _74790_/B _71010_/X _71735_/D _74790_/X sky130_fd_sc_hd__and4_4
X_86776_ _86784_/CLK _46082_/Y _67296_/B sky130_fd_sc_hd__dfxtp_4
X_83988_ _87671_/CLK _83988_/D _83988_/Q sky130_fd_sc_hd__dfxtp_4
X_42921_ _42680_/A _42951_/A sky130_fd_sc_hd__buf_2
X_54907_ _54893_/X _54907_/B _54907_/Y sky130_fd_sc_hd__nand2_4
X_73741_ _72874_/A _73742_/A sky130_fd_sc_hd__buf_2
X_85727_ _85727_/CLK _52939_/Y _85727_/Q sky130_fd_sc_hd__dfxtp_4
X_70953_ _51261_/B _70936_/X _70952_/Y _83652_/D sky130_fd_sc_hd__o21ai_4
X_58675_ _58687_/A _86392_/Q _58675_/Y sky130_fd_sc_hd__nor2_4
X_82939_ _84981_/CLK _82939_/D _82939_/Q sky130_fd_sc_hd__dfxtp_4
X_55887_ _55884_/X _55886_/X _44115_/A _55891_/A sky130_fd_sc_hd__a21o_4
X_45640_ _63182_/B _61513_/A sky130_fd_sc_hd__buf_2
X_57626_ _84966_/Q _57603_/X _57625_/Y _57626_/Y sky130_fd_sc_hd__o21ai_4
X_76460_ _76458_/Y _76459_/Y _76460_/X sky130_fd_sc_hd__and2_4
X_42852_ _42820_/X _42852_/X sky130_fd_sc_hd__buf_2
X_54838_ _54834_/Y _54830_/X _54837_/X _85369_/D sky130_fd_sc_hd__a21oi_4
X_73672_ _73670_/X _73671_/Y _73546_/X _73672_/X sky130_fd_sc_hd__a21o_4
X_85658_ _85433_/CLK _53308_/Y _85658_/Q sky130_fd_sc_hd__dfxtp_4
X_70884_ _70884_/A _70884_/B _70695_/A _70885_/A sky130_fd_sc_hd__nor3_4
X_75411_ _75411_/A _80965_/Q _75411_/Y sky130_fd_sc_hd__nand2_4
X_41803_ _41825_/A _41803_/X sky130_fd_sc_hd__buf_2
X_72623_ _79184_/B _79183_/A sky130_fd_sc_hd__inv_2
X_84609_ _84606_/CLK _60511_/Y _79149_/A sky130_fd_sc_hd__dfxtp_4
X_45571_ _45720_/A _45571_/X sky130_fd_sc_hd__buf_2
X_57557_ _57554_/Y _57543_/X _57556_/Y _84980_/D sky130_fd_sc_hd__a21boi_4
X_76391_ _76377_/Y _76389_/Y _76390_/Y _76391_/X sky130_fd_sc_hd__o21a_4
X_88377_ _87865_/CLK _88377_/D _88377_/Q sky130_fd_sc_hd__dfxtp_4
X_42783_ _42782_/Y _87721_/D sky130_fd_sc_hd__inv_2
X_54769_ _85381_/Q _54757_/X _54768_/Y _54769_/Y sky130_fd_sc_hd__o21ai_4
X_85589_ _86193_/CLK _85589_/D _85589_/Q sky130_fd_sc_hd__dfxtp_4
X_47310_ _47310_/A _52977_/D sky130_fd_sc_hd__buf_2
X_78130_ _78130_/A _78130_/B _78130_/C _78130_/D _78131_/B sky130_fd_sc_hd__and4_4
X_44522_ _87068_/Q _44522_/Y sky130_fd_sc_hd__inv_2
X_56508_ _56545_/A _56094_/A _56507_/Y _85169_/D sky130_fd_sc_hd__o21ai_4
X_75342_ _75309_/A _75324_/Y _75322_/X _75342_/X sky130_fd_sc_hd__and3_4
X_87328_ _87595_/CLK _87328_/D _87328_/Q sky130_fd_sc_hd__dfxtp_4
X_41734_ _40402_/A _81741_/Q _41733_/X _41734_/X sky130_fd_sc_hd__o21a_4
X_48290_ _86541_/Q _48263_/X _48289_/Y _48290_/Y sky130_fd_sc_hd__o21ai_4
X_72554_ _72539_/B _72579_/A sky130_fd_sc_hd__buf_2
X_57488_ _84994_/Q _57380_/X _57486_/Y _57487_/X _84994_/D sky130_fd_sc_hd__a211o_4
Xclkbuf_8_30_0_CLK clkbuf_8_31_0_CLK/A clkbuf_9_61_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_47241_ _47147_/A _47241_/X sky130_fd_sc_hd__buf_2
X_71505_ _58463_/Y _71486_/A _71504_/Y _71505_/Y sky130_fd_sc_hd__o21ai_4
X_59227_ _59152_/X _59224_/Y _59226_/Y _59169_/X _59156_/X _59227_/X
+ sky130_fd_sc_hd__o32a_4
X_78061_ _84566_/Q _78061_/B _78061_/X sky130_fd_sc_hd__xor2_4
X_44453_ _44602_/A _44453_/X sky130_fd_sc_hd__buf_2
X_56439_ _56439_/A _56439_/X sky130_fd_sc_hd__buf_2
X_75273_ _75254_/Y _75258_/B _75256_/Y _75274_/A sky130_fd_sc_hd__o21a_4
X_41665_ _41319_/B _41653_/X _41665_/X sky130_fd_sc_hd__or2_4
X_87259_ _87273_/CLK _87259_/D _69469_/B sky130_fd_sc_hd__dfxtp_4
X_72485_ _59398_/A _72488_/B sky130_fd_sc_hd__buf_2
X_77012_ _77013_/A _77013_/B _77012_/Y sky130_fd_sc_hd__nor2_4
X_43404_ _43305_/A _43404_/X sky130_fd_sc_hd__buf_2
X_74224_ _74224_/A _73152_/X _74224_/Y sky130_fd_sc_hd__nor2_4
X_40616_ _40585_/X _82875_/Q _40615_/X _40616_/Y sky130_fd_sc_hd__o21ai_4
X_47172_ _47168_/Y _47128_/X _47171_/X _47172_/Y sky130_fd_sc_hd__a21oi_4
X_59158_ _59143_/Y _59145_/X _59151_/X _59157_/X _84765_/D sky130_fd_sc_hd__a22oi_4
X_71436_ _71419_/Y _83500_/Q _71435_/X _83500_/D sky130_fd_sc_hd__a21o_4
X_44384_ _44381_/X _44382_/X _41786_/X _87137_/Q _44383_/X _44385_/A
+ sky130_fd_sc_hd__o32ai_4
X_41596_ _41595_/X _41596_/X sky130_fd_sc_hd__buf_2
X_58109_ _58793_/A _58109_/X sky130_fd_sc_hd__buf_2
X_46123_ _46138_/A _46119_/A _46124_/A sky130_fd_sc_hd__and2_4
X_43335_ _41294_/X _43325_/X _87474_/Q _43326_/X _87474_/D sky130_fd_sc_hd__a2bb2o_4
X_74155_ _73163_/A _74155_/X sky130_fd_sc_hd__buf_2
X_40547_ _40463_/X _41624_/A _40546_/X _40547_/Y sky130_fd_sc_hd__o21ai_4
X_59089_ _58941_/A _86362_/Q _59089_/Y sky130_fd_sc_hd__nor2_4
X_71367_ _71344_/A _83523_/Q _71366_/X _71367_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_8_45_0_CLK clkbuf_8_45_0_CLK/A clkbuf_8_45_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_61120_ _61083_/C _61112_/X _61205_/A _61120_/Y sky130_fd_sc_hd__nand3_4
X_73106_ _73106_/A _44127_/X _73106_/Y sky130_fd_sc_hd__nor2_4
X_46054_ _43030_/A _46054_/X sky130_fd_sc_hd__buf_2
X_70318_ _70318_/A _70183_/A _70183_/B _70183_/D _70318_/Y sky130_fd_sc_hd__nand4_4
X_43266_ _41098_/X _43264_/X _87510_/Q _43265_/X _87510_/D sky130_fd_sc_hd__a2bb2o_4
X_74086_ _74082_/X _74084_/X _74085_/X _74090_/A sky130_fd_sc_hd__a21o_4
X_78963_ _78957_/B _78957_/A _78962_/Y _78964_/B sky130_fd_sc_hd__a21oi_4
X_40478_ _82319_/Q _40471_/X _40478_/X sky130_fd_sc_hd__or2_4
X_71298_ _71303_/A _71303_/B _71297_/X _71298_/Y sky130_fd_sc_hd__nand3_4
X_45005_ _55934_/B _44963_/X _45004_/X _45005_/X sky130_fd_sc_hd__o21a_4
X_42217_ _42217_/A _42217_/Y sky130_fd_sc_hd__inv_2
X_61051_ _60918_/X _60921_/X _60911_/X _61051_/Y sky130_fd_sc_hd__o21ai_4
X_77914_ _82069_/Q _81941_/D _77913_/X _77914_/Y sky130_fd_sc_hd__o21ai_4
X_73037_ _69700_/B _44235_/X _73035_/X _73036_/Y _73037_/X sky130_fd_sc_hd__a211o_4
X_70249_ _70134_/X _70249_/X sky130_fd_sc_hd__buf_2
X_43197_ _43196_/X _43167_/X _40914_/X _73465_/A _43172_/X _43197_/Y
+ sky130_fd_sc_hd__o32ai_4
X_78894_ _78880_/Y _78893_/X _78894_/Y sky130_fd_sc_hd__nand2_4
X_60002_ _59977_/B _60091_/C sky130_fd_sc_hd__buf_2
X_49813_ _49809_/A _53025_/B _49813_/Y sky130_fd_sc_hd__nand2_4
X_42148_ _42137_/A _42148_/X sky130_fd_sc_hd__buf_2
X_77845_ _82271_/Q _81983_/Q _77845_/Y sky130_fd_sc_hd__xnor2_4
X_64810_ _64810_/A _86458_/Q _64810_/X sky130_fd_sc_hd__and2_4
X_49744_ _49757_/A _52959_/B _49744_/Y sky130_fd_sc_hd__nand2_4
X_46956_ _46909_/X _46959_/A sky130_fd_sc_hd__buf_2
X_42079_ _42052_/X _42077_/X _40972_/X _88044_/Q _42078_/X _42080_/A
+ sky130_fd_sc_hd__o32ai_4
X_65790_ _65790_/A _65790_/X sky130_fd_sc_hd__buf_2
X_77776_ _77776_/A _81928_/D _77796_/A sky130_fd_sc_hd__xnor2_4
X_74988_ _74988_/A _74988_/B _74988_/Y sky130_fd_sc_hd__nand2_4
X_79515_ _84816_/Q _84136_/Q _79515_/Y sky130_fd_sc_hd__nand2_4
X_45907_ _45907_/A _45907_/Y sky130_fd_sc_hd__inv_2
X_64741_ _64870_/A _64741_/B _64741_/C _64741_/Y sky130_fd_sc_hd__nor3_4
X_76727_ _81483_/Q _76727_/Y sky130_fd_sc_hd__inv_2
X_49675_ _49661_/X _52889_/B _49675_/Y sky130_fd_sc_hd__nand2_4
X_73939_ _73939_/A _73939_/X sky130_fd_sc_hd__buf_2
X_61953_ _61499_/B _61953_/B _61953_/C _61937_/X _61953_/Y sky130_fd_sc_hd__nand4_4
X_46887_ _52732_/B _51043_/B sky130_fd_sc_hd__buf_2
X_48626_ _83569_/Q _48627_/A sky130_fd_sc_hd__inv_2
X_60904_ _60879_/B _64081_/C sky130_fd_sc_hd__buf_2
X_67460_ _67460_/A _87662_/Q _67460_/X sky130_fd_sc_hd__and2_4
X_79446_ _84811_/Q _84131_/Q _79446_/X sky130_fd_sc_hd__xor2_4
X_45838_ _45829_/X _45833_/Y _45837_/Y _45838_/Y sky130_fd_sc_hd__a21oi_4
X_64672_ _64669_/X _64671_/X _64619_/X _64672_/X sky130_fd_sc_hd__a21o_4
X_76658_ _76657_/Y _81395_/Q _76658_/Y sky130_fd_sc_hd__nand2_4
X_61884_ _59721_/X _61915_/A sky130_fd_sc_hd__buf_2
X_66411_ _66411_/A _66411_/X sky130_fd_sc_hd__buf_2
X_63623_ _63621_/Y _63578_/X _63622_/Y _63623_/Y sky130_fd_sc_hd__a21oi_4
X_75609_ _75602_/Y _75607_/Y _75608_/Y _75609_/Y sky130_fd_sc_hd__a21oi_4
X_48557_ _48557_/A _52188_/B _48557_/Y sky130_fd_sc_hd__nand2_4
X_60835_ _60422_/A _60835_/X sky130_fd_sc_hd__buf_2
X_67391_ _67270_/X _67391_/X sky130_fd_sc_hd__buf_2
X_79377_ _79361_/X _79364_/Y _79377_/X sky130_fd_sc_hd__or2_4
X_45769_ _85065_/Q _45736_/B _45769_/Y sky130_fd_sc_hd__nor2_4
X_76589_ _76588_/X _76589_/Y sky130_fd_sc_hd__inv_2
X_69130_ _87072_/Q _69058_/X _69103_/X _69129_/X _69130_/X sky130_fd_sc_hd__a211o_4
X_47508_ _58132_/A _47478_/X _47507_/Y _47508_/Y sky130_fd_sc_hd__o21ai_4
X_66342_ _66282_/X _65884_/Y _66341_/Y _66342_/Y sky130_fd_sc_hd__o21ai_4
X_78328_ _78330_/A _78330_/B _78329_/A sky130_fd_sc_hd__nor2_4
X_63554_ _63554_/A _63554_/B _63554_/C _63554_/Y sky130_fd_sc_hd__nor3_4
X_48488_ _48545_/A _48533_/C sky130_fd_sc_hd__buf_2
X_60766_ _60652_/X _60724_/B _60624_/X _60659_/A _60766_/X sky130_fd_sc_hd__and4_4
X_62505_ _61570_/B _62504_/X _62449_/X _62475_/X _62506_/D sky130_fd_sc_hd__nand4_4
X_69061_ _68737_/A _69061_/X sky130_fd_sc_hd__buf_2
X_47439_ _54739_/D _53048_/D sky130_fd_sc_hd__buf_2
X_66273_ _66326_/A _86536_/Q _66273_/X sky130_fd_sc_hd__and2_4
X_78259_ _78251_/A _78256_/B _78250_/A _78259_/Y sky130_fd_sc_hd__o21ai_4
X_63485_ _63496_/A _58511_/A _63458_/X _63496_/D _63485_/X sky130_fd_sc_hd__and4_4
X_60697_ _60660_/X _60697_/B _60697_/Y sky130_fd_sc_hd__nand2_4
X_68012_ _67657_/X _68371_/A sky130_fd_sc_hd__buf_2
X_65224_ _65400_/A _65224_/X sky130_fd_sc_hd__buf_2
X_50450_ _86198_/Q _50437_/X _50449_/Y _50450_/Y sky130_fd_sc_hd__o21ai_4
X_62436_ _59950_/C _62436_/X sky130_fd_sc_hd__buf_2
X_81270_ _81697_/CLK _81270_/D _76459_/A sky130_fd_sc_hd__dfxtp_4
X_49109_ _86443_/Q _49104_/X _49108_/Y _49109_/Y sky130_fd_sc_hd__o21ai_4
X_80221_ _80221_/A _80221_/B _80221_/X sky130_fd_sc_hd__and2_4
X_65155_ _65155_/A _65155_/B _65155_/X sky130_fd_sc_hd__and2_4
X_50381_ _50381_/A _50381_/B _50381_/Y sky130_fd_sc_hd__nand2_4
X_62367_ _62214_/A _62367_/X sky130_fd_sc_hd__buf_2
X_52120_ _52116_/Y _52117_/X _52119_/Y _52120_/Y sky130_fd_sc_hd__a21boi_4
X_64106_ _84842_/Q _64136_/B _64106_/X sky130_fd_sc_hd__or2_4
X_61318_ _61313_/A _72575_/A sky130_fd_sc_hd__buf_2
X_80152_ _84944_/Q _84192_/Q _80154_/A sky130_fd_sc_hd__xor2_4
X_65086_ _65083_/X _65085_/X _64989_/X _65086_/X sky130_fd_sc_hd__a21o_4
X_69963_ _69960_/X _69962_/X _60371_/A _69963_/Y sky130_fd_sc_hd__a21oi_4
X_62298_ _61387_/X _62309_/B _62309_/C _62211_/D _62298_/Y sky130_fd_sc_hd__nand4_4
X_52051_ _52048_/Y _52049_/X _52050_/X _52051_/Y sky130_fd_sc_hd__a21oi_4
X_64037_ _64074_/A _64074_/B _64037_/C _64037_/Y sky130_fd_sc_hd__nor3_4
X_68914_ _44725_/A _68472_/X _44246_/A _68913_/X _68914_/X sky130_fd_sc_hd__a211o_4
X_61249_ _60371_/X _59901_/A _63004_/B _44003_/X _59802_/X _61249_/Y
+ sky130_fd_sc_hd__a41oi_4
X_84960_ _84960_/CLK _84960_/D _84960_/Q sky130_fd_sc_hd__dfxtp_4
X_80083_ _80081_/X _80088_/B _80083_/Y sky130_fd_sc_hd__xnor2_4
X_69894_ _69988_/A _69894_/X sky130_fd_sc_hd__buf_2
X_51002_ _50999_/Y _50983_/X _51001_/X _51002_/Y sky130_fd_sc_hd__a21oi_4
X_83911_ _81933_/CLK _83911_/D _81983_/D sky130_fd_sc_hd__dfxtp_4
X_68845_ _44719_/A _68472_/X _44246_/A _68844_/X _68845_/X sky130_fd_sc_hd__a211o_4
X_84891_ _84250_/CLK _84891_/D _84891_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_opt_20_CLK _85555_/CLK _85553_/CLK sky130_fd_sc_hd__clkbuf_16
X_55810_ _55807_/X _55809_/X _55811_/A sky130_fd_sc_hd__and2_4
X_86630_ _85990_/CLK _86630_/D _86630_/Q sky130_fd_sc_hd__dfxtp_4
X_83842_ _83842_/CLK _83842_/D _83842_/Q sky130_fd_sc_hd__dfxtp_4
X_56790_ _56787_/X _56766_/X _57163_/C _56788_/X _57170_/A _56790_/X
+ sky130_fd_sc_hd__a41o_4
X_68776_ _87087_/Q _68353_/X _68354_/X _68775_/X _68776_/X sky130_fd_sc_hd__a211o_4
X_65988_ _65970_/A _65970_/B _84164_/Q _65988_/X sky130_fd_sc_hd__and3_4
X_67727_ _67793_/A _67727_/B _67727_/X sky130_fd_sc_hd__and2_4
X_55741_ _55741_/A _55741_/B _55741_/X sky130_fd_sc_hd__and2_4
X_86561_ _83561_/CLK _86561_/D _73568_/B sky130_fd_sc_hd__dfxtp_4
X_52953_ _53062_/A _52977_/C sky130_fd_sc_hd__buf_2
X_64939_ _64939_/A _64939_/X sky130_fd_sc_hd__buf_2
X_83773_ _84981_/CLK _70443_/Y _47959_/A sky130_fd_sc_hd__dfxtp_4
X_80985_ _80813_/CLK _80985_/D _80985_/Q sky130_fd_sc_hd__dfxtp_4
X_88300_ _88097_/CLK _40974_/Y _88300_/Q sky130_fd_sc_hd__dfxtp_4
X_85512_ _85800_/CLK _85512_/D _85512_/Q sky130_fd_sc_hd__dfxtp_4
X_51904_ _51823_/A _51904_/X sky130_fd_sc_hd__buf_2
X_58460_ _58459_/Y _58461_/A sky130_fd_sc_hd__buf_2
X_82724_ _84115_/CLK _84108_/Q _78831_/A sky130_fd_sc_hd__dfxtp_4
X_55672_ _55287_/A _55674_/B _55672_/X sky130_fd_sc_hd__and2_4
X_67658_ _67657_/X _67658_/X sky130_fd_sc_hd__buf_2
X_86492_ _85596_/CLK _86492_/D _72911_/B sky130_fd_sc_hd__dfxtp_4
X_52884_ _52882_/Y _52865_/X _52883_/X _52884_/Y sky130_fd_sc_hd__a21oi_4
X_57411_ _56694_/Y _57400_/X _57411_/Y sky130_fd_sc_hd__nand2_4
X_88231_ _86930_/CLK _41353_/X _88231_/Q sky130_fd_sc_hd__dfxtp_4
X_54623_ _54636_/A _54097_/B _54623_/Y sky130_fd_sc_hd__nand2_4
X_66609_ _66683_/A _66609_/B _66609_/X sky130_fd_sc_hd__and2_4
X_85443_ _85764_/CLK _85443_/D _85443_/Q sky130_fd_sc_hd__dfxtp_4
X_51835_ _51820_/A _50971_/B _51835_/Y sky130_fd_sc_hd__nand2_4
X_82655_ _81756_/CLK _84007_/Q _82655_/Q sky130_fd_sc_hd__dfxtp_4
X_58391_ _58391_/A _58403_/B _58391_/Y sky130_fd_sc_hd__nand2_4
X_67589_ _67496_/X _67577_/Y _67507_/X _67588_/Y _67589_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_342_0_CLK clkbuf_9_171_0_CLK/X _85645_/CLK sky130_fd_sc_hd__clkbuf_1
X_81606_ _81257_/CLK _76213_/B _81606_/Q sky130_fd_sc_hd__dfxtp_4
X_57342_ _57341_/Y _57342_/Y sky130_fd_sc_hd__inv_2
X_88162_ _87652_/CLK _88162_/D _88162_/Q sky130_fd_sc_hd__dfxtp_4
X_69328_ _81396_/D _69299_/X _69327_/X _83932_/D sky130_fd_sc_hd__a21bo_4
X_54554_ _54552_/Y _54530_/X _54553_/X _54554_/Y sky130_fd_sc_hd__a21oi_4
X_85374_ _83711_/CLK _54811_/Y _85374_/Q sky130_fd_sc_hd__dfxtp_4
X_51766_ _85950_/Q _51763_/X _51765_/Y _51766_/Y sky130_fd_sc_hd__o21ai_4
X_82586_ _82589_/CLK _82586_/D _78248_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_972_0_CLK clkbuf_9_486_0_CLK/X _83282_/CLK sky130_fd_sc_hd__clkbuf_1
X_87113_ _87421_/CLK _87113_/D _87113_/Q sky130_fd_sc_hd__dfxtp_4
X_53505_ _53502_/Y _53498_/X _53504_/Y _85624_/D sky130_fd_sc_hd__a21boi_4
X_84325_ _84321_/CLK _63421_/Y _80579_/B sky130_fd_sc_hd__dfxtp_4
X_50717_ _86147_/Q _50706_/X _50716_/Y _50717_/Y sky130_fd_sc_hd__o21ai_4
X_57273_ _57270_/X _57273_/B _57149_/B _56733_/X _57273_/Y sky130_fd_sc_hd__nand4_4
X_81537_ _83940_/CLK _81537_/D _81537_/Q sky130_fd_sc_hd__dfxtp_4
X_69259_ _69191_/A _87786_/Q _69259_/X sky130_fd_sc_hd__and2_4
X_88093_ _87588_/CLK _88093_/D _41957_/A sky130_fd_sc_hd__dfxtp_4
X_54485_ _54376_/A _54485_/X sky130_fd_sc_hd__buf_2
X_51697_ _51697_/A _53219_/B _51697_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_463_0_CLK clkbuf_8_231_0_CLK/X clkbuf_9_463_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_59012_ _58925_/X _85440_/Q _59011_/X _59012_/Y sky130_fd_sc_hd__o21ai_4
X_56224_ _56070_/X _56210_/X _56223_/Y _56224_/Y sky130_fd_sc_hd__o21ai_4
X_87044_ _88326_/CLK _87044_/D _87044_/Q sky130_fd_sc_hd__dfxtp_4
X_53436_ _51822_/A _53436_/X sky130_fd_sc_hd__buf_2
X_41450_ _40947_/A _41482_/A sky130_fd_sc_hd__buf_2
X_72270_ _44171_/X _72270_/X sky130_fd_sc_hd__buf_2
X_84256_ _83766_/CLK _84256_/D _79784_/B sky130_fd_sc_hd__dfxtp_4
X_50648_ _50643_/Y _50644_/X _50647_/Y _50648_/Y sky130_fd_sc_hd__a21boi_4
X_81468_ _84064_/CLK _81468_/D _81468_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_357_0_CLK clkbuf_9_178_0_CLK/X _84766_/CLK sky130_fd_sc_hd__clkbuf_1
X_40401_ _40400_/X _40342_/X _88397_/Q _40355_/X _88397_/D sky130_fd_sc_hd__a2bb2o_4
X_71221_ _71221_/A _71232_/A sky130_fd_sc_hd__buf_2
X_83207_ _83843_/CLK _83207_/D _70178_/C sky130_fd_sc_hd__dfxtp_4
X_80419_ _84757_/Q _80419_/B _80419_/Y sky130_fd_sc_hd__nand2_4
X_56155_ _56142_/X _56153_/X _56154_/Y _85286_/D sky130_fd_sc_hd__o21ai_4
X_41381_ _41373_/X _41725_/A _41380_/X _41381_/X sky130_fd_sc_hd__o21a_4
X_53367_ _53371_/A _53371_/B _53371_/C _52853_/D _53367_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_987_0_CLK clkbuf_9_493_0_CLK/X _83305_/CLK sky130_fd_sc_hd__clkbuf_1
X_84187_ _84187_/CLK _84187_/D _84187_/Q sky130_fd_sc_hd__dfxtp_4
X_50579_ _50578_/X _71974_/B sky130_fd_sc_hd__buf_2
X_81399_ _81351_/CLK _83935_/Q _76690_/B sky130_fd_sc_hd__dfxtp_4
X_43120_ _43105_/X _43106_/X _40781_/X _43119_/Y _43108_/X _43120_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55106_ _55118_/A _47788_/A _55106_/Y sky130_fd_sc_hd__nand2_4
X_40332_ _41863_/A _40332_/Y sky130_fd_sc_hd__inv_2
X_52318_ _64904_/B _52297_/X _52317_/Y _52318_/Y sky130_fd_sc_hd__o21ai_4
X_71152_ _71178_/A _71155_/B _71152_/C _71160_/D _71152_/Y sky130_fd_sc_hd__nand4_4
X_83138_ _83141_/CLK _73749_/Y _83138_/Q sky130_fd_sc_hd__dfxtp_4
X_56086_ _56100_/A _56086_/B _55851_/B _56086_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_9_478_0_CLK clkbuf_9_479_0_CLK/A clkbuf_9_478_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_53298_ _53298_/A _54473_/B _53298_/Y sky130_fd_sc_hd__nand2_4
X_70103_ _70103_/A _70107_/A sky130_fd_sc_hd__inv_2
X_43051_ _43038_/X _43050_/X _40641_/X _73773_/A _43025_/X _43052_/A
+ sky130_fd_sc_hd__o32ai_4
X_59914_ _59552_/B _61293_/B sky130_fd_sc_hd__buf_2
X_55037_ _55037_/A _54871_/B _55037_/Y sky130_fd_sc_hd__nand2_4
X_52249_ _52246_/Y _52232_/X _52248_/X _85860_/D sky130_fd_sc_hd__a21oi_4
X_71083_ _49006_/X _71070_/X _71082_/Y _71083_/Y sky130_fd_sc_hd__o21ai_4
X_83069_ _83572_/CLK _74427_/Y _83069_/Q sky130_fd_sc_hd__dfxtp_4
X_75960_ _81704_/D _75968_/B _75961_/A sky130_fd_sc_hd__xor2_4
X_87946_ _87950_/CLK _87946_/D _87946_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_910_0_CLK clkbuf_9_455_0_CLK/X _88104_/CLK sky130_fd_sc_hd__clkbuf_1
X_42002_ _42002_/A _42002_/Y sky130_fd_sc_hd__inv_2
X_74911_ _80939_/Q _74911_/B _81188_/D sky130_fd_sc_hd__xor2_4
X_70034_ _68734_/X _68736_/X _70005_/X _70034_/Y sky130_fd_sc_hd__a21oi_4
X_59845_ _59801_/A _60781_/A sky130_fd_sc_hd__buf_2
X_75891_ _75891_/A _80773_/D sky130_fd_sc_hd__inv_2
X_87877_ _87883_/CLK _87877_/D _87877_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_401_0_CLK clkbuf_8_200_0_CLK/X clkbuf_9_401_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_46810_ _46809_/Y _46810_/X sky130_fd_sc_hd__buf_2
Xclkbuf_opt_11_CLK _84914_/CLK _84885_/CLK sky130_fd_sc_hd__clkbuf_16
X_77630_ _77630_/A _82109_/D _77633_/B sky130_fd_sc_hd__nor2_4
X_74842_ _46183_/X _74842_/B _46184_/Y _80672_/D sky130_fd_sc_hd__and3_4
X_86828_ _86824_/CLK _45984_/Y _66810_/B sky130_fd_sc_hd__dfxtp_4
X_47790_ _72447_/A _47760_/X _47789_/Y _47790_/Y sky130_fd_sc_hd__o21ai_4
X_59776_ _59770_/A _72176_/A sky130_fd_sc_hd__buf_2
X_56988_ _56982_/X _56986_/X _56987_/Y _56988_/Y sky130_fd_sc_hd__a21oi_4
X_46741_ _46733_/A _46740_/X _46741_/Y sky130_fd_sc_hd__nand2_4
X_58727_ _58727_/A _58688_/B _58727_/Y sky130_fd_sc_hd__nor2_4
X_77561_ _77561_/A _77561_/B _77561_/C _77561_/D _77561_/X sky130_fd_sc_hd__and4_4
X_43953_ _43949_/X _43952_/X _80669_/Q _43959_/A sky130_fd_sc_hd__a21o_4
X_55939_ _56206_/C _55605_/X _44090_/B _55938_/X _55939_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_925_0_CLK clkbuf_9_462_0_CLK/X _83544_/CLK sky130_fd_sc_hd__clkbuf_1
X_74773_ _74753_/X _70637_/A _74773_/C _74739_/B _74773_/X sky130_fd_sc_hd__and4_4
X_86759_ _80854_/CLK _46220_/Y _44174_/A sky130_fd_sc_hd__dfxtp_4
X_71985_ _71985_/A _71985_/X sky130_fd_sc_hd__buf_2
X_79300_ _84797_/Q _66469_/C _79302_/A sky130_fd_sc_hd__xor2_4
X_76512_ _76511_/X _76517_/A sky130_fd_sc_hd__buf_2
X_42904_ _42903_/Y _87660_/D sky130_fd_sc_hd__inv_2
X_49460_ _49434_/A _49460_/X sky130_fd_sc_hd__buf_2
X_73724_ _42475_/Y _73674_/X _73698_/X _73723_/Y _73724_/X sky130_fd_sc_hd__a211o_4
X_46672_ _46719_/A _46672_/X sky130_fd_sc_hd__buf_2
X_58658_ _58655_/Y _58657_/Y _58646_/X _58658_/X sky130_fd_sc_hd__a21o_4
X_70936_ _70935_/X _70936_/X sky130_fd_sc_hd__buf_2
X_77492_ _77473_/Y _77475_/A _77472_/A _77493_/A sky130_fd_sc_hd__o21a_4
X_43884_ _41298_/X _43879_/X _67395_/B _43880_/X _87217_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_9_416_0_CLK clkbuf_8_208_0_CLK/X clkbuf_9_416_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_48411_ _74389_/B _52121_/B sky130_fd_sc_hd__buf_2
X_79231_ _79231_/A _79231_/B _79232_/B sky130_fd_sc_hd__xnor2_4
X_57609_ _57608_/X _57609_/B _57609_/Y sky130_fd_sc_hd__nand2_4
X_45623_ _63168_/B _61502_/A sky130_fd_sc_hd__buf_2
X_76443_ _76443_/A _76443_/Y sky130_fd_sc_hd__inv_2
X_42835_ _42579_/A _42835_/X sky130_fd_sc_hd__buf_2
X_49391_ _58633_/B _49388_/X _49390_/Y _49391_/Y sky130_fd_sc_hd__o21ai_4
X_73655_ _73651_/X _73654_/X _56549_/X _73655_/X sky130_fd_sc_hd__a21o_4
X_70867_ _70867_/A _70869_/B _70869_/C _70869_/D _70867_/Y sky130_fd_sc_hd__nand4_4
X_58589_ _58701_/A _58589_/X sky130_fd_sc_hd__buf_2
X_48342_ _48342_/A _50381_/B sky130_fd_sc_hd__buf_2
X_60620_ _60353_/B _60620_/B _60620_/C _60620_/Y sky130_fd_sc_hd__nand3_4
X_72606_ _72579_/A _72510_/C _59846_/X _72606_/X sky130_fd_sc_hd__a21o_4
X_79162_ _84786_/Q _66524_/C _79524_/A sky130_fd_sc_hd__or2_4
X_45554_ _45551_/Y _45489_/X _45520_/X _45553_/Y _45554_/X sky130_fd_sc_hd__a211o_4
X_76374_ _76381_/A _76373_/X _81617_/D sky130_fd_sc_hd__xnor2_4
Xclkbuf_6_1_0_CLK clkbuf_6_1_0_CLK/A clkbuf_7_3_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_42766_ _41298_/X _42757_/X _67392_/B _42759_/X _87729_/D sky130_fd_sc_hd__a2bb2o_4
X_73586_ _73449_/X _85632_/Q _73450_/X _73585_/X _73586_/X sky130_fd_sc_hd__a211o_4
X_70798_ _70356_/Y _70423_/X _70907_/B MACRO_WR_SELECT _70798_/X
+ sky130_fd_sc_hd__and4_4
X_78113_ _78105_/Y _78130_/A _78130_/B _78120_/A sky130_fd_sc_hd__nand3_4
X_44505_ _41264_/A _44502_/X _87076_/Q _44503_/X _44505_/X sky130_fd_sc_hd__a2bb2o_4
X_75325_ _75322_/X _75324_/Y _75325_/Y sky130_fd_sc_hd__nand2_4
X_41717_ _40421_/X _41717_/X sky130_fd_sc_hd__buf_2
X_48273_ _48226_/A _48273_/X sky130_fd_sc_hd__buf_2
X_60551_ _60570_/C _60602_/B _60267_/A _60551_/X sky130_fd_sc_hd__o21a_4
X_72537_ _72535_/Y _72537_/B _72537_/Y sky130_fd_sc_hd__nand2_4
X_79093_ _79088_/Y _79070_/B _79092_/Y _79095_/B sky130_fd_sc_hd__o21ai_4
X_45485_ _85083_/Q _45485_/Y sky130_fd_sc_hd__inv_2
X_42697_ _41104_/X _42695_/X _69542_/B _42696_/X _87765_/D sky130_fd_sc_hd__a2bb2o_4
X_47224_ _47128_/A _47224_/X sky130_fd_sc_hd__buf_2
X_78044_ _78044_/A _81922_/D sky130_fd_sc_hd__inv_2
X_44436_ _44425_/X _44427_/X _41596_/X _87109_/Q _44428_/X _44437_/A
+ sky130_fd_sc_hd__o32ai_4
X_75256_ _75255_/A _80943_/D _75256_/Y sky130_fd_sc_hd__nand2_4
X_63270_ _58277_/A _62999_/X _61607_/B _60608_/X _63270_/Y sky130_fd_sc_hd__a2bb2oi_4
X_41648_ _41647_/X _41638_/X _67421_/B _41639_/X _88176_/D sky130_fd_sc_hd__a2bb2o_4
X_60482_ _60482_/A _60482_/Y sky130_fd_sc_hd__inv_2
X_72468_ _72361_/X _85667_/Q _72362_/X _72468_/X sky130_fd_sc_hd__o21a_4
X_62221_ _62572_/A _62362_/A sky130_fd_sc_hd__buf_2
X_74207_ _69055_/B _73030_/X _73035_/X _74206_/Y _74207_/X sky130_fd_sc_hd__a211o_4
X_47155_ _47152_/X _47133_/B _47143_/C _51192_/D _47155_/X sky130_fd_sc_hd__and4_4
X_71419_ _71419_/A _71419_/Y sky130_fd_sc_hd__inv_2
X_44367_ _41745_/X _44364_/X _87145_/Q _44365_/X _44367_/X sky130_fd_sc_hd__a2bb2o_4
X_75187_ _75172_/Y _75169_/Y _75175_/C _75188_/A sky130_fd_sc_hd__o21a_4
X_41579_ _41577_/X _81162_/Q _41578_/X _41580_/A sky130_fd_sc_hd__o21ai_4
X_72399_ _72396_/Y _72398_/Y _57718_/A _72399_/X sky130_fd_sc_hd__a21o_4
X_46106_ _46085_/A _46107_/A sky130_fd_sc_hd__buf_2
X_43318_ _43318_/A _87484_/D sky130_fd_sc_hd__inv_2
X_62152_ _62151_/X _62175_/B _61761_/C _62046_/D _62152_/Y sky130_fd_sc_hd__nand4_4
X_74138_ _70128_/C _73549_/X _74137_/Y _83121_/D sky130_fd_sc_hd__a21o_4
X_47086_ _47080_/Y _47081_/X _47085_/X _86672_/D sky130_fd_sc_hd__a21oi_4
X_44298_ _69442_/A _44299_/A sky130_fd_sc_hd__buf_2
X_79995_ _79985_/A _79985_/B _79994_/Y _79995_/Y sky130_fd_sc_hd__a21boi_4
X_61103_ _61102_/X _61103_/X sky130_fd_sc_hd__buf_2
X_46037_ _46013_/X _46032_/X _41492_/X _86800_/Q _46014_/X _46038_/A
+ sky130_fd_sc_hd__o32ai_4
X_43249_ _41050_/X _43247_/X _87519_/Q _43248_/X _43249_/X sky130_fd_sc_hd__a2bb2o_4
X_66960_ _87939_/Q _66935_/X _66911_/X _66959_/X _66960_/X sky130_fd_sc_hd__a211o_4
X_62083_ _61730_/X _62094_/B _59722_/X _62083_/D _62083_/X sky130_fd_sc_hd__and4_4
X_74069_ _74067_/X _74068_/Y _73982_/X _74069_/X sky130_fd_sc_hd__a21o_4
X_78946_ _78946_/A _78945_/Y _78947_/B sky130_fd_sc_hd__xnor2_4
X_65911_ _65896_/A _73568_/B _65911_/X sky130_fd_sc_hd__and2_4
X_61034_ _60967_/X _60995_/Y _61024_/Y _61032_/X _61033_/X _84534_/D
+ sky130_fd_sc_hd__o41a_4
X_66891_ _66888_/X _66890_/X _66843_/X _66891_/X sky130_fd_sc_hd__a21o_4
X_78877_ _78877_/A _78877_/B _78877_/X sky130_fd_sc_hd__and2_4
X_68630_ _68993_/A _68630_/X sky130_fd_sc_hd__buf_2
X_65842_ _65842_/A _65842_/X sky130_fd_sc_hd__buf_2
X_77828_ _77828_/A _77814_/Y _77828_/Y sky130_fd_sc_hd__nor2_4
X_47988_ _47988_/A _50306_/B _47988_/Y sky130_fd_sc_hd__nand2_4
X_49727_ _86334_/Q _49715_/X _49726_/Y _49727_/Y sky130_fd_sc_hd__o21ai_4
X_68561_ _44688_/A _68455_/X _68509_/X _68560_/X _68561_/X sky130_fd_sc_hd__a211o_4
X_46939_ _59019_/A _46908_/X _46938_/Y _46939_/Y sky130_fd_sc_hd__o21ai_4
X_65773_ _64961_/A _65969_/A sky130_fd_sc_hd__buf_2
X_77759_ _77758_/Y _77745_/Y _77752_/A _77759_/Y sky130_fd_sc_hd__o21ai_4
X_62985_ _59961_/A _64328_/A sky130_fd_sc_hd__buf_2
X_67512_ _67987_/A _67512_/X sky130_fd_sc_hd__buf_2
X_64724_ _65718_/A _64724_/X sky130_fd_sc_hd__buf_2
X_49658_ _49651_/X _49642_/B _49669_/C _52872_/D _49658_/X sky130_fd_sc_hd__and4_4
X_61936_ _61708_/X _61953_/C sky130_fd_sc_hd__buf_2
X_80770_ _80854_/CLK _75887_/Y _80770_/Q sky130_fd_sc_hd__dfxtp_4
X_68492_ _73675_/A _68414_/X _68379_/X _68491_/Y _68492_/X sky130_fd_sc_hd__a211o_4
X_48609_ _48609_/A _50511_/A sky130_fd_sc_hd__buf_2
X_79429_ _79429_/A _79428_/Y _79429_/X sky130_fd_sc_hd__xor2_4
X_67443_ _67438_/X _67441_/X _67442_/X _67443_/X sky130_fd_sc_hd__a21o_4
X_64655_ _64652_/X _64654_/X _64629_/X _64655_/X sky130_fd_sc_hd__a21o_4
X_49589_ _49586_/Y _49570_/X _49588_/X _86360_/D sky130_fd_sc_hd__a21oi_4
X_61867_ _59765_/A _61915_/B sky130_fd_sc_hd__buf_2
X_51620_ _51618_/Y _51613_/X _51619_/X _85977_/D sky130_fd_sc_hd__a21oi_4
X_63606_ _60731_/A _63655_/A sky130_fd_sc_hd__buf_2
X_82440_ _82452_/CLK _79132_/X _82440_/Q sky130_fd_sc_hd__dfxtp_4
X_60818_ _60616_/Y _60704_/Y _60815_/X _60794_/Y _60817_/Y _84559_/D
+ sky130_fd_sc_hd__a41oi_4
X_67374_ _86974_/Q _67348_/X _67278_/X _67373_/X _67374_/X sky130_fd_sc_hd__a211o_4
X_64586_ _64777_/A _64676_/A sky130_fd_sc_hd__buf_2
X_61798_ _61796_/X _61765_/B _61846_/C _61748_/X _61798_/Y sky130_fd_sc_hd__nand4_4
X_69113_ _68385_/A _69113_/X sky130_fd_sc_hd__buf_2
X_66325_ _66322_/X _66324_/X _58882_/A _66325_/X sky130_fd_sc_hd__a21o_4
X_51551_ _85989_/Q _51539_/X _51550_/Y _51551_/Y sky130_fd_sc_hd__o21ai_4
X_63537_ _63512_/A _57680_/A _63537_/C _63537_/X sky130_fd_sc_hd__and3_4
X_82371_ _84951_/CLK _82371_/D _82371_/Q sky130_fd_sc_hd__dfxtp_4
X_60749_ _60646_/Y _63417_/A _60725_/A _60749_/Y sky130_fd_sc_hd__nand3_4
X_84110_ _84111_/CLK _84110_/D _84110_/Q sky130_fd_sc_hd__dfxtp_4
X_50502_ _86188_/Q _50499_/X _50501_/Y _50502_/Y sky130_fd_sc_hd__o21ai_4
X_81322_ _81322_/CLK _76274_/X _81698_/D sky130_fd_sc_hd__dfxtp_4
X_69044_ _69442_/A _69044_/X sky130_fd_sc_hd__buf_2
X_54270_ _54286_/A _54246_/X _54286_/C _46619_/A _54270_/X sky130_fd_sc_hd__and4_4
X_66256_ _66326_/A _66256_/B _66256_/X sky130_fd_sc_hd__and2_4
X_85090_ _85031_/CLK _57085_/X _85090_/Q sky130_fd_sc_hd__dfxtp_4
X_51482_ _86002_/Q _51458_/X _51481_/Y _51482_/Y sky130_fd_sc_hd__o21ai_4
X_63468_ _63468_/A _63517_/B sky130_fd_sc_hd__buf_2
X_53221_ _53221_/A _53302_/A sky130_fd_sc_hd__buf_2
X_65207_ _65099_/X _83290_/Q _65028_/X _65206_/X _65207_/X sky130_fd_sc_hd__a211o_4
X_84041_ _81169_/CLK _68092_/X _82081_/D sky130_fd_sc_hd__dfxtp_4
X_50433_ _86201_/Q _50403_/X _50432_/Y _50433_/Y sky130_fd_sc_hd__o21ai_4
X_62419_ _62448_/A _58528_/A _62375_/C _62421_/C sky130_fd_sc_hd__nand3_4
X_81253_ _81288_/CLK _81285_/Q _76187_/A sky130_fd_sc_hd__dfxtp_4
X_66187_ _66226_/A _86542_/Q _66187_/X sky130_fd_sc_hd__and2_4
X_63399_ _63427_/A _61780_/X _63399_/X sky130_fd_sc_hd__and2_4
X_80204_ _80196_/A _80195_/X _80203_/Y _80204_/Y sky130_fd_sc_hd__a21boi_4
X_53152_ _53149_/Y _53137_/X _53151_/X _53152_/Y sky130_fd_sc_hd__a21oi_4
X_65138_ _65065_/X _83293_/Q _65108_/X _65137_/X _65138_/X sky130_fd_sc_hd__a211o_4
X_50364_ _50500_/A _50383_/A sky130_fd_sc_hd__buf_2
X_81184_ _86758_/CLK _75066_/B _81184_/Q sky130_fd_sc_hd__dfxtp_4
X_52103_ _52103_/A _52135_/B _52097_/X _52103_/X sky130_fd_sc_hd__and3_4
X_87800_ _87544_/CLK _87800_/D _69917_/A sky130_fd_sc_hd__dfxtp_4
X_80135_ _80131_/Y _80134_/Y _80135_/X sky130_fd_sc_hd__xor2_4
X_53083_ _53112_/A _53107_/A sky130_fd_sc_hd__buf_2
X_57960_ _86640_/Q _58039_/B _57960_/Y sky130_fd_sc_hd__nor2_4
X_65069_ _65056_/Y _65068_/Y _65069_/Y sky130_fd_sc_hd__nand2_4
X_69946_ _44149_/A _42620_/Y _69946_/Y sky130_fd_sc_hd__nor2_4
X_50295_ _50279_/X _53520_/B _50295_/Y sky130_fd_sc_hd__nand2_4
X_85992_ _85704_/CLK _85992_/D _85992_/Q sky130_fd_sc_hd__dfxtp_4
X_52034_ _48287_/A _51972_/X _52033_/X _52034_/X sky130_fd_sc_hd__and3_4
X_56911_ _56876_/X _83330_/Q _56985_/D sky130_fd_sc_hd__nor2_4
X_87731_ _88180_/CLK _87731_/D _67333_/B sky130_fd_sc_hd__dfxtp_4
X_84943_ _82386_/CLK _84943_/D _84943_/Q sky130_fd_sc_hd__dfxtp_4
X_80066_ _84935_/Q _65713_/C _80066_/Y sky130_fd_sc_hd__nand2_4
X_57891_ _57952_/A _57891_/B _57891_/Y sky130_fd_sc_hd__nor2_4
X_69877_ _69877_/A _88316_/Q _69877_/X sky130_fd_sc_hd__and2_4
X_59630_ _59961_/A _65680_/A sky130_fd_sc_hd__buf_2
X_56842_ _56842_/A _56842_/X sky130_fd_sc_hd__buf_2
X_68828_ _57803_/A _69648_/A sky130_fd_sc_hd__buf_2
X_87662_ _87915_/CLK _87662_/D _87662_/Q sky130_fd_sc_hd__dfxtp_4
X_84874_ _83451_/CLK _84874_/D _58338_/A sky130_fd_sc_hd__dfxtp_4
X_86613_ _85969_/CLK _86613_/D _86613_/Q sky130_fd_sc_hd__dfxtp_4
X_59561_ _59557_/X _59598_/A _59890_/C _59751_/A sky130_fd_sc_hd__nand3_4
X_83825_ _83187_/CLK _83825_/D _74804_/B sky130_fd_sc_hd__dfxtp_4
X_56773_ _56771_/X _56772_/Y _44292_/A _56773_/Y sky130_fd_sc_hd__a21oi_4
X_68759_ _68759_/A _87236_/Q _68759_/X sky130_fd_sc_hd__and2_4
X_87593_ _87595_/CLK _43056_/Y _87593_/Q sky130_fd_sc_hd__dfxtp_4
X_53985_ _53956_/X _53985_/B _53985_/Y sky130_fd_sc_hd__nand2_4
X_58512_ _58492_/X _58508_/Y _58511_/Y _58512_/Y sky130_fd_sc_hd__a21oi_4
X_55724_ _55245_/A _55724_/B _55724_/X sky130_fd_sc_hd__and2_4
X_86544_ _86549_/CLK _48278_/Y _66159_/B sky130_fd_sc_hd__dfxtp_4
X_52936_ _52944_/A _52936_/B _52936_/Y sky130_fd_sc_hd__nand2_4
X_40950_ _40950_/A _40950_/X sky130_fd_sc_hd__buf_2
X_71770_ _71763_/X _70476_/X _70794_/X _71770_/X sky130_fd_sc_hd__and3_4
X_83756_ _83756_/CLK _83756_/D _57674_/A sky130_fd_sc_hd__dfxtp_4
X_59492_ _84717_/Q _63410_/B sky130_fd_sc_hd__buf_2
X_80968_ _80968_/CLK _80968_/D _80956_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_281_0_CLK clkbuf_9_140_0_CLK/X _83421_/CLK sky130_fd_sc_hd__clkbuf_1
X_70721_ _70721_/A _70769_/D sky130_fd_sc_hd__buf_2
X_58443_ _58423_/X _83479_/Q _58442_/Y _84847_/D sky130_fd_sc_hd__o21a_4
X_82707_ _82665_/CLK _78965_/X _82663_/D sky130_fd_sc_hd__dfxtp_4
X_55655_ _55655_/A _55655_/B _55656_/A sky130_fd_sc_hd__and2_4
X_86475_ _86505_/CLK _86475_/D _86475_/Q sky130_fd_sc_hd__dfxtp_4
X_40881_ _40881_/A _40881_/X sky130_fd_sc_hd__buf_2
X_52867_ _52867_/A _52853_/B _52853_/C _52867_/D _52867_/X sky130_fd_sc_hd__and4_4
X_83687_ _82394_/CLK _70840_/Y _83687_/Q sky130_fd_sc_hd__dfxtp_4
X_80899_ _84074_/CLK _80899_/D _80899_/Q sky130_fd_sc_hd__dfxtp_4
X_88214_ _88208_/CLK _41444_/Y _88214_/Q sky130_fd_sc_hd__dfxtp_4
X_42620_ _73484_/A _42620_/Y sky130_fd_sc_hd__inv_2
X_54606_ _85411_/Q _54593_/X _54605_/Y _54606_/Y sky130_fd_sc_hd__o21ai_4
X_73440_ _73440_/A _73577_/B _73440_/Y sky130_fd_sc_hd__nor2_4
X_85426_ _85651_/CLK _54527_/Y _85426_/Q sky130_fd_sc_hd__dfxtp_4
X_51818_ _50063_/A _53269_/A sky130_fd_sc_hd__buf_2
X_70652_ _70638_/A _70656_/D sky130_fd_sc_hd__buf_2
Xclkbuf_10_63_0_CLK clkbuf_9_31_0_CLK/X _83335_/CLK sky130_fd_sc_hd__clkbuf_1
X_58374_ _58374_/A _58344_/B _58374_/Y sky130_fd_sc_hd__nor2_4
X_82638_ _84003_/CLK _82638_/D _82638_/Q sky130_fd_sc_hd__dfxtp_4
X_55586_ _45460_/A _55571_/X _55610_/A _55585_/Y _55586_/X sky130_fd_sc_hd__a211o_4
X_52798_ _52795_/Y _52783_/X _52797_/X _52798_/Y sky130_fd_sc_hd__a21oi_4
XPHY_30 sky130_fd_sc_hd__decap_3
X_57325_ _57324_/X _57318_/Y _56704_/X _57325_/Y sky130_fd_sc_hd__a21oi_4
XPHY_41 sky130_fd_sc_hd__decap_3
X_88145_ _88398_/CLK _41805_/Y _66621_/B sky130_fd_sc_hd__dfxtp_4
X_42551_ _42536_/X _42547_/X _40781_/X _42550_/Y _42538_/X _42551_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54537_ _54537_/A _54538_/C sky130_fd_sc_hd__buf_2
X_73371_ _69888_/B _73026_/X _73028_/X _73371_/Y sky130_fd_sc_hd__o21ai_4
X_85357_ _86282_/CLK _85357_/D _85357_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_52 sky130_fd_sc_hd__decap_3
X_51749_ _51814_/A _51749_/X sky130_fd_sc_hd__buf_2
X_70583_ _70582_/X _70583_/X sky130_fd_sc_hd__buf_2
X_82569_ _82879_/CLK _82569_/D _82569_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_63 sky130_fd_sc_hd__decap_3
Xclkbuf_7_108_0_CLK clkbuf_6_54_0_CLK/X clkbuf_8_217_0_CLK/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_296_0_CLK clkbuf_9_148_0_CLK/X _84299_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_74 sky130_fd_sc_hd__decap_3
X_75110_ _75110_/A _75113_/A sky130_fd_sc_hd__inv_2
X_41502_ _41481_/X _82329_/Q _41501_/X _41502_/Y sky130_fd_sc_hd__o21ai_4
XPHY_85 sky130_fd_sc_hd__decap_3
X_72322_ _72313_/Y _72237_/X _72318_/X _72321_/X _83265_/D sky130_fd_sc_hd__a22oi_4
X_84308_ _84308_/CLK _63623_/Y _80400_/B sky130_fd_sc_hd__dfxtp_4
X_45270_ _85289_/Q _45269_/X _45229_/X _45270_/X sky130_fd_sc_hd__o21a_4
X_57256_ _57243_/X _56619_/X _85048_/Q _57245_/X _85048_/D sky130_fd_sc_hd__a2bb2o_4
X_76090_ _81529_/Q _76090_/B _76090_/X sky130_fd_sc_hd__xor2_4
XPHY_96 sky130_fd_sc_hd__decap_3
X_42482_ _42482_/A _42482_/Y sky130_fd_sc_hd__inv_2
X_88076_ _87821_/CLK _88076_/D _88076_/Q sky130_fd_sc_hd__dfxtp_4
X_54468_ _54465_/Y _54448_/X _54467_/X _85437_/D sky130_fd_sc_hd__a21oi_4
X_85288_ _83016_/CLK _85288_/D _56145_/C sky130_fd_sc_hd__dfxtp_4
X_44221_ _44146_/A _68057_/A sky130_fd_sc_hd__buf_2
X_56207_ _56031_/X _56195_/X _56206_/Y _56207_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_78_0_CLK clkbuf_9_39_0_CLK/X _86873_/CLK sky130_fd_sc_hd__clkbuf_1
X_75041_ _75039_/X _75051_/B _75041_/Y sky130_fd_sc_hd__nand2_4
X_41433_ _41432_/Y _41433_/X sky130_fd_sc_hd__buf_2
X_87027_ _87032_/CLK _44629_/Y _87027_/Q sky130_fd_sc_hd__dfxtp_4
X_53419_ _53418_/X _53420_/A sky130_fd_sc_hd__buf_2
X_72253_ _86614_/Q _72348_/B _72253_/Y sky130_fd_sc_hd__nor2_4
X_84239_ _84603_/CLK _64510_/Y _79605_/B sky130_fd_sc_hd__dfxtp_4
X_57187_ _57187_/A _57188_/A sky130_fd_sc_hd__buf_2
X_54399_ _54399_/A _54399_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_224_0_CLK clkbuf_8_225_0_CLK/A clkbuf_8_224_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_71204_ _70387_/A _71228_/B sky130_fd_sc_hd__buf_2
X_44152_ _44152_/A _44265_/D sky130_fd_sc_hd__buf_2
X_56138_ _55773_/D _56138_/B _56138_/Y sky130_fd_sc_hd__xnor2_4
X_41364_ _41361_/X _41362_/X _67672_/B _41363_/X _88229_/D sky130_fd_sc_hd__a2bb2o_4
X_72184_ _59368_/X _85980_/Q _72183_/X _72184_/Y sky130_fd_sc_hd__o21ai_4
X_43103_ _43103_/A _43103_/Y sky130_fd_sc_hd__inv_2
X_78800_ _78797_/A _78798_/A _78797_/B _78801_/B sky130_fd_sc_hd__nand3_4
X_71135_ _70428_/A _71137_/A sky130_fd_sc_hd__buf_2
X_48960_ _50599_/A _50599_/B _48917_/X _48960_/X sky130_fd_sc_hd__o21a_4
X_44083_ _55620_/A _44085_/C sky130_fd_sc_hd__buf_2
X_56069_ _74317_/C _56068_/X _56069_/Y sky130_fd_sc_hd__xnor2_4
X_79780_ _79777_/X _79780_/B _79780_/Y sky130_fd_sc_hd__xnor2_4
X_41295_ _41294_/X _41283_/X _67373_/B _41284_/X _88242_/D sky130_fd_sc_hd__a2bb2o_4
X_76992_ _84544_/Q _84416_/Q _76992_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_9_340_0_CLK clkbuf_9_341_0_CLK/A clkbuf_9_340_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_47911_ _57523_/B _50268_/B sky130_fd_sc_hd__buf_2
X_43034_ _43058_/A _43034_/X sky130_fd_sc_hd__buf_2
X_78731_ _78731_/A _78732_/C sky130_fd_sc_hd__inv_2
X_71066_ _71058_/A _71066_/B _71066_/C _71066_/Y sky130_fd_sc_hd__nand3_4
X_75943_ _75940_/Y _75942_/Y _75944_/B sky130_fd_sc_hd__xor2_4
X_87929_ _87417_/CLK _87929_/D _87929_/Q sky130_fd_sc_hd__dfxtp_4
X_48891_ _48642_/A _48891_/B _48891_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_239_0_CLK clkbuf_8_239_0_CLK/A clkbuf_9_479_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_234_0_CLK clkbuf_9_117_0_CLK/X _80817_/CLK sky130_fd_sc_hd__clkbuf_1
X_70017_ _70011_/X _68597_/Y _70012_/X _70016_/Y _70017_/X sky130_fd_sc_hd__a211o_4
X_47842_ _47842_/A _73591_/A sky130_fd_sc_hd__inv_2
X_59828_ _59512_/A _59875_/A sky130_fd_sc_hd__buf_2
X_78662_ _78661_/Y _78663_/C sky130_fd_sc_hd__inv_2
X_75874_ _75870_/Y _75873_/Y _75876_/A sky130_fd_sc_hd__nand2_4
Xclkbuf_10_864_0_CLK clkbuf_9_432_0_CLK/X _86553_/CLK sky130_fd_sc_hd__clkbuf_1
X_77613_ _77612_/Y _77614_/C sky130_fd_sc_hd__inv_2
Xclkbuf_10_16_0_CLK clkbuf_9_8_0_CLK/X _85167_/CLK sky130_fd_sc_hd__clkbuf_1
X_74825_ _74829_/A _46087_/A _74826_/A sky130_fd_sc_hd__nand2_4
X_47773_ _47799_/A _53236_/B _47773_/Y sky130_fd_sc_hd__nand2_4
X_59759_ _59806_/A _59761_/A sky130_fd_sc_hd__buf_2
X_78593_ _78600_/B _78593_/B _82773_/D sky130_fd_sc_hd__xnor2_4
X_44985_ _44887_/X _45212_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_355_0_CLK clkbuf_9_355_0_CLK/A clkbuf_9_355_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_49512_ _49502_/A _51037_/B _49512_/Y sky130_fd_sc_hd__nand2_4
X_46724_ _58700_/A _46719_/X _46723_/Y _46724_/Y sky130_fd_sc_hd__o21ai_4
X_77544_ _77520_/B _77516_/X _77561_/B sky130_fd_sc_hd__nand2_4
X_43936_ _43916_/X _43924_/X _41442_/X _87190_/Q _43917_/X _43937_/A
+ sky130_fd_sc_hd__o32ai_4
X_74756_ _74775_/A _74756_/B _70884_/A _70662_/X _74756_/X sky130_fd_sc_hd__and4_4
X_62770_ _62819_/A _64335_/C _62737_/X _62738_/D _62770_/X sky130_fd_sc_hd__and4_4
X_71968_ _83311_/Q _57635_/X _71967_/Y _71968_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_249_0_CLK clkbuf_9_124_0_CLK/X _81883_/CLK sky130_fd_sc_hd__clkbuf_1
X_49443_ _49415_/A _49443_/X sky130_fd_sc_hd__buf_2
X_61721_ _61412_/A _61722_/A sky130_fd_sc_hd__buf_2
X_73707_ _73607_/A _73707_/B _73707_/X sky130_fd_sc_hd__and2_4
X_46655_ _46892_/A _46845_/A sky130_fd_sc_hd__buf_2
X_70919_ _70867_/A _70914_/B _70914_/C _70919_/D _70919_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_10_879_0_CLK clkbuf_9_439_0_CLK/X _86149_/CLK sky130_fd_sc_hd__clkbuf_1
X_77475_ _77475_/A _77475_/B _77476_/A sky130_fd_sc_hd__nor2_4
X_43867_ _43867_/A _43867_/Y sky130_fd_sc_hd__inv_2
X_74687_ _74687_/A _74687_/Y sky130_fd_sc_hd__inv_2
X_71899_ _56842_/X _71892_/X _71898_/Y _83336_/D sky130_fd_sc_hd__o21ai_4
X_79214_ _84790_/Q _84110_/Q _79215_/A sky130_fd_sc_hd__or2_4
X_45606_ _45604_/Y _45605_/Y _44939_/B _45606_/X sky130_fd_sc_hd__o21a_4
X_64440_ _64440_/A _64440_/X sky130_fd_sc_hd__buf_2
X_76426_ _76426_/A _76430_/A sky130_fd_sc_hd__inv_2
X_42818_ _42816_/X _42817_/X _41442_/X _87702_/Q _42805_/X _42818_/Y
+ sky130_fd_sc_hd__o32ai_4
X_61652_ _61608_/X _61652_/B _61675_/C _61652_/Y sky130_fd_sc_hd__nand3_4
X_49374_ _49374_/A _49369_/X _49380_/C _51761_/D _49374_/X sky130_fd_sc_hd__and4_4
X_73638_ _73638_/A _73638_/B _73638_/X sky130_fd_sc_hd__and2_4
X_46586_ _46585_/Y _51389_/B sky130_fd_sc_hd__buf_2
X_43798_ _43790_/X _43797_/X _41054_/X _69427_/B _43791_/X _43799_/A
+ sky130_fd_sc_hd__o32ai_4
X_60603_ _60435_/C _60341_/A _60603_/C _60578_/Y _60603_/X sky130_fd_sc_hd__and4_4
X_48325_ _48348_/A _50368_/B _48325_/Y sky130_fd_sc_hd__nand2_4
X_79145_ _79145_/A _84477_/Q _79145_/X sky130_fd_sc_hd__xor2_4
X_45537_ _85016_/Q _55539_/B sky130_fd_sc_hd__inv_2
X_64371_ _64360_/Y _64370_/X _64328_/X _64371_/X sky130_fd_sc_hd__o21a_4
X_76357_ _76338_/A _76357_/Y sky130_fd_sc_hd__inv_2
X_42749_ _42749_/A _42749_/Y sky130_fd_sc_hd__inv_2
X_61583_ _61317_/X _72575_/A _61260_/X _61319_/X _61283_/Y _61583_/Y
+ sky130_fd_sc_hd__a41oi_4
X_73569_ _73566_/X _84993_/Q _73385_/X _73568_/X _73569_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_802_0_CLK clkbuf_9_401_0_CLK/X _82015_/CLK sky130_fd_sc_hd__clkbuf_1
X_66110_ _66106_/Y _66065_/X _66109_/Y _84156_/D sky130_fd_sc_hd__a21o_4
X_63322_ _60454_/A _64524_/B _60441_/B _63237_/X _63322_/X sky130_fd_sc_hd__and4_4
X_75308_ _75304_/Y _75283_/Y _75307_/X _75308_/Y sky130_fd_sc_hd__o21ai_4
X_48256_ _47984_/B _48257_/B sky130_fd_sc_hd__buf_2
X_60534_ _60533_/Y _60566_/A _65842_/A _60534_/Y sky130_fd_sc_hd__a21oi_4
X_67090_ _66947_/X _67078_/Y _67031_/X _67089_/Y _67090_/X sky130_fd_sc_hd__a211o_4
X_79076_ _79064_/A _79064_/B _79076_/Y sky130_fd_sc_hd__nor2_4
X_45468_ _45434_/X _61378_/A _45452_/X _45468_/Y sky130_fd_sc_hd__o21ai_4
X_76288_ _81259_/Q _81515_/D _76282_/C _76288_/Y sky130_fd_sc_hd__a21boi_4
X_47207_ _59373_/A _47192_/X _47206_/Y _47207_/Y sky130_fd_sc_hd__o21ai_4
X_66041_ _65980_/X _66041_/B _66041_/X sky130_fd_sc_hd__and2_4
X_78027_ _78021_/C _78027_/B _78031_/A sky130_fd_sc_hd__nand2_4
X_44419_ _41552_/X _44412_/X _87118_/Q _44413_/X _87118_/D sky130_fd_sc_hd__a2bb2o_4
X_63253_ _84844_/Q _63281_/B _63301_/C _63281_/D _63253_/X sky130_fd_sc_hd__or4_4
X_75239_ _75239_/A _80986_/Q _75251_/A sky130_fd_sc_hd__xor2_4
X_48187_ _48535_/A _48478_/A sky130_fd_sc_hd__buf_2
X_60465_ _60421_/B _60488_/A _60488_/B _60476_/C _59980_/X _60465_/Y
+ sky130_fd_sc_hd__a41oi_4
X_45399_ _45393_/Y _45394_/X _45396_/X _45398_/Y _45399_/X sky130_fd_sc_hd__a211o_4
X_62204_ _62203_/Y _62620_/A sky130_fd_sc_hd__buf_2
X_47138_ _86666_/Q _47096_/X _47137_/Y _47138_/Y sky130_fd_sc_hd__o21ai_4
X_63184_ _63177_/Y _63179_/X _63180_/X _63182_/X _63183_/X _63184_/Y
+ sky130_fd_sc_hd__o41ai_4
Xclkbuf_10_817_0_CLK clkbuf_9_408_0_CLK/X _82923_/CLK sky130_fd_sc_hd__clkbuf_1
X_60396_ _60395_/X _60459_/B sky130_fd_sc_hd__buf_2
X_69800_ _69795_/X _69800_/B _69800_/Y sky130_fd_sc_hd__nand2_4
X_62135_ _62037_/X _62021_/B _63672_/B _62020_/X _62135_/X sky130_fd_sc_hd__and4_4
X_47069_ _47069_/A _53353_/B sky130_fd_sc_hd__inv_2
X_67992_ _67992_/A _67992_/B _67992_/X sky130_fd_sc_hd__and2_4
X_79978_ _79973_/Y _79976_/Y _79978_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_308_0_CLK clkbuf_8_154_0_CLK/X clkbuf_9_308_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_69731_ _83901_/Q _69696_/X _69730_/X _83901_/D sky130_fd_sc_hd__a21bo_4
X_50080_ _50084_/A _52287_/B _50080_/Y sky130_fd_sc_hd__nand2_4
X_66943_ _88388_/Q _66868_/X _66919_/X _66942_/X _66943_/X sky130_fd_sc_hd__a211o_4
X_62066_ _59794_/X _62088_/B _62061_/Y _62066_/D _62066_/Y sky130_fd_sc_hd__nand4_4
X_78929_ _82848_/Q _82560_/Q _78930_/B sky130_fd_sc_hd__xnor2_4
X_61017_ _61036_/C _61016_/Y _60952_/X _76987_/A _60898_/X _84539_/D
+ sky130_fd_sc_hd__o32a_4
X_81940_ _82131_/CLK _81940_/D _81940_/Q sky130_fd_sc_hd__dfxtp_4
X_69662_ _88076_/Q _68640_/X _69088_/X _69661_/Y _69662_/X sky130_fd_sc_hd__a211o_4
X_66874_ _80917_/D _66850_/X _66873_/X _84093_/D sky130_fd_sc_hd__a21bo_4
X_68613_ _66540_/A _68613_/X sky130_fd_sc_hd__buf_2
X_65825_ _65825_/A _86503_/Q _65825_/X sky130_fd_sc_hd__and2_4
X_69593_ _87569_/Q _69506_/X _68436_/X _69592_/X _69593_/X sky130_fd_sc_hd__a211o_4
X_81871_ _81872_/CLK _78062_/X _81839_/D sky130_fd_sc_hd__dfxtp_4
X_83610_ _83613_/CLK _71092_/Y _83610_/Q sky130_fd_sc_hd__dfxtp_4
X_80822_ _81994_/CLK _80822_/D _75605_/B sky130_fd_sc_hd__dfxtp_4
X_68544_ _88012_/Q _69796_/A _68540_/X _68543_/X _68544_/X sky130_fd_sc_hd__a211o_4
X_53770_ _53766_/A _48694_/A _53770_/Y sky130_fd_sc_hd__nand2_4
X_65756_ _65747_/Y _65756_/B _65756_/Y sky130_fd_sc_hd__nand2_4
X_84590_ _84590_/CLK _60601_/Y _79130_/A sky130_fd_sc_hd__dfxtp_4
X_50982_ _86095_/Q _50965_/X _50981_/Y _50982_/Y sky130_fd_sc_hd__o21ai_4
X_62968_ _62964_/Y _62886_/X _62965_/Y _62966_/Y _62967_/X _62968_/X
+ sky130_fd_sc_hd__a41o_4
X_52721_ _52719_/Y _52702_/X _52720_/X _52721_/Y sky130_fd_sc_hd__a21oi_4
X_64707_ _64980_/A _64707_/X sky130_fd_sc_hd__buf_2
X_83541_ _86541_/CLK _71307_/Y _48039_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_5_8_0_CLK clkbuf_4_4_1_CLK/X clkbuf_5_8_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_61919_ _61481_/X _61874_/B _61907_/C _61874_/D _61919_/Y sky130_fd_sc_hd__nand4_4
X_80753_ _80746_/CLK _75297_/X _81129_/D sky130_fd_sc_hd__dfxtp_4
X_68475_ _69004_/A _88367_/Q _68475_/X sky130_fd_sc_hd__and2_4
X_65687_ _65702_/A _85872_/Q _65687_/X sky130_fd_sc_hd__and2_4
X_62899_ _84844_/Q _62642_/B _62899_/Y sky130_fd_sc_hd__nor2_4
X_55440_ _55439_/Y _55387_/X _55441_/B sky130_fd_sc_hd__nand2_4
X_67426_ _81502_/D _67331_/X _67425_/X _84070_/D sky130_fd_sc_hd__a21bo_4
X_86260_ _85555_/CLK _86260_/D _64948_/B sky130_fd_sc_hd__dfxtp_4
X_52652_ _85779_/Q _52629_/X _52651_/Y _52652_/Y sky130_fd_sc_hd__o21ai_4
X_64638_ _64637_/X _64638_/B _81024_/D _64638_/X sky130_fd_sc_hd__and3_4
X_83472_ _86600_/CLK _83472_/D _83472_/Q sky130_fd_sc_hd__dfxtp_4
X_80684_ _80681_/CLK _80716_/Q _80684_/Q sky130_fd_sc_hd__dfxtp_4
X_85211_ _85244_/CLK _85211_/D _56392_/C sky130_fd_sc_hd__dfxtp_4
X_51603_ _51619_/A _51603_/B _51603_/C _53129_/D _51603_/X sky130_fd_sc_hd__and4_4
X_82423_ _82463_/CLK _82455_/Q _78611_/A sky130_fd_sc_hd__dfxtp_4
X_55371_ _55325_/X _55384_/A _55371_/X sky130_fd_sc_hd__and2_4
X_67357_ _87922_/Q _67355_/X _67284_/X _67356_/X _67357_/X sky130_fd_sc_hd__a211o_4
X_86191_ _86191_/CLK _50488_/Y _86191_/Q sky130_fd_sc_hd__dfxtp_4
X_52583_ _85792_/Q _52575_/X _52582_/Y _52583_/Y sky130_fd_sc_hd__o21ai_4
XPHY_606 sky130_fd_sc_hd__decap_3
X_64569_ _64611_/A _85825_/Q _64569_/X sky130_fd_sc_hd__and2_4
XPHY_617 sky130_fd_sc_hd__decap_3
XPHY_628 sky130_fd_sc_hd__decap_3
X_57110_ _57221_/A _57110_/X sky130_fd_sc_hd__buf_2
X_54322_ _54322_/A _54332_/A sky130_fd_sc_hd__buf_2
XPHY_639 sky130_fd_sc_hd__decap_3
X_66308_ _66267_/X _85893_/Q _66308_/X sky130_fd_sc_hd__and2_4
X_85142_ _85144_/CLK _85142_/D _55529_/B sky130_fd_sc_hd__dfxtp_4
X_51534_ _51530_/Y _51531_/X _51533_/X _85993_/D sky130_fd_sc_hd__a21oi_4
X_58090_ _58065_/X _85702_/Q _58089_/X _58090_/X sky130_fd_sc_hd__o21a_4
X_82354_ _82558_/CLK _77168_/X _82354_/Q sky130_fd_sc_hd__dfxtp_4
X_67288_ _87349_/Q _67239_/X _67240_/X _67287_/X _67288_/X sky130_fd_sc_hd__a211o_4
X_57041_ _56838_/A _57331_/A sky130_fd_sc_hd__buf_2
X_81305_ _81689_/CLK _76993_/X _81305_/Q sky130_fd_sc_hd__dfxtp_4
X_69027_ _69027_/A _88344_/Q _69027_/X sky130_fd_sc_hd__and2_4
X_54253_ _54253_/A _54253_/X sky130_fd_sc_hd__buf_2
X_66239_ _66236_/X _85610_/Q _66096_/X _66238_/X _66239_/X sky130_fd_sc_hd__a211o_4
X_85073_ _85071_/CLK _85073_/D _57137_/A sky130_fd_sc_hd__dfxtp_4
X_51465_ _86005_/Q _51458_/X _51464_/Y _51465_/Y sky130_fd_sc_hd__o21ai_4
X_82285_ _82301_/CLK _82285_/D _41048_/A sky130_fd_sc_hd__dfxtp_4
X_53204_ _53201_/Y _53189_/X _53203_/X _85678_/D sky130_fd_sc_hd__a21oi_4
X_84024_ _81169_/CLK _84024_/D _84024_/Q sky130_fd_sc_hd__dfxtp_4
X_50416_ _50572_/A _50556_/A sky130_fd_sc_hd__buf_2
X_81236_ _85332_/CLK _81044_/Q _47653_/A sky130_fd_sc_hd__dfxtp_4
X_54184_ _54184_/A _47385_/Y _54184_/Y sky130_fd_sc_hd__nand2_4
X_51396_ _51396_/A _51352_/B _51352_/C _51396_/X sky130_fd_sc_hd__and3_4
X_53135_ _53121_/X _53135_/B _53135_/Y sky130_fd_sc_hd__nand2_4
X_50347_ _52050_/A _50331_/B _50338_/X _50347_/X sky130_fd_sc_hd__and3_4
X_81167_ _81179_/CLK _74940_/B _81167_/Q sky130_fd_sc_hd__dfxtp_4
X_58992_ _58982_/X _83435_/Q _58991_/Y _58992_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_7_70_0_CLK clkbuf_7_70_0_CLK/A clkbuf_7_70_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_80118_ _80105_/X _80116_/X _80117_/X _80118_/Y sky130_fd_sc_hd__a21oi_4
X_41080_ _40901_/B _41079_/X _41080_/X sky130_fd_sc_hd__or2_4
X_53066_ _53147_/A _53080_/A sky130_fd_sc_hd__buf_2
X_57943_ _84938_/Q _57896_/X _57936_/X _57942_/X _57943_/Y sky130_fd_sc_hd__a2bb2oi_4
X_69929_ _69929_/A _69929_/Y sky130_fd_sc_hd__inv_2
X_50278_ _86232_/Q _50250_/X _50277_/Y _50278_/Y sky130_fd_sc_hd__o21ai_4
X_85975_ _85688_/CLK _51631_/Y _85975_/Q sky130_fd_sc_hd__dfxtp_4
X_81098_ _81065_/CLK _79645_/X _81098_/Q sky130_fd_sc_hd__dfxtp_4
X_52017_ _50314_/A _51972_/X _51958_/C _52017_/X sky130_fd_sc_hd__and3_4
X_87714_ _87210_/CLK _87714_/D _87714_/Q sky130_fd_sc_hd__dfxtp_4
X_72940_ _72938_/X _72926_/X _72928_/X _72940_/Y sky130_fd_sc_hd__nand3_4
X_84926_ _84926_/CLK _84926_/D _84926_/Q sky130_fd_sc_hd__dfxtp_4
X_80049_ _60097_/C _80049_/B _80057_/B sky130_fd_sc_hd__xor2_4
X_57874_ _58834_/A _58703_/A sky130_fd_sc_hd__buf_2
Xclkbuf_1_0_1_CLK clkbuf_1_0_0_CLK/X clkbuf_1_0_2_CLK/A sky130_fd_sc_hd__clkbuf_1
X_59613_ _60627_/A _60626_/A _59613_/Y sky130_fd_sc_hd__nor2_4
X_56825_ _56824_/X _85130_/Q _56825_/Y sky130_fd_sc_hd__nand2_4
X_87645_ _87195_/CLK _42932_/X _87645_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_85_0_CLK clkbuf_7_85_0_CLK/A clkbuf_7_85_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_72871_ _73040_/A _85885_/Q _72871_/X sky130_fd_sc_hd__and2_4
X_84857_ _84360_/CLK _84857_/D _84857_/Q sky130_fd_sc_hd__dfxtp_4
X_74610_ _74605_/X _74599_/X _56144_/A _74600_/X _74610_/X sky130_fd_sc_hd__a211o_4
X_71822_ _71804_/Y _83362_/Q _71821_/X _71822_/X sky130_fd_sc_hd__a21o_4
X_83808_ _81807_/CLK _83808_/D _74796_/A sky130_fd_sc_hd__dfxtp_4
X_59544_ _59544_/A _59544_/B _59890_/B _59544_/D _59545_/A sky130_fd_sc_hd__and4_4
X_44770_ _44770_/A _44770_/Y sky130_fd_sc_hd__inv_2
X_56756_ _56755_/X _56756_/X sky130_fd_sc_hd__buf_2
X_75590_ _75889_/A _75589_/Y _75590_/X sky130_fd_sc_hd__or2_4
X_87576_ _87577_/CLK _87576_/D _43098_/A sky130_fd_sc_hd__dfxtp_4
X_41982_ _41998_/A _41982_/X sky130_fd_sc_hd__buf_2
X_53968_ _51814_/A _53969_/C sky130_fd_sc_hd__buf_2
X_84788_ _86695_/CLK _58945_/Y _84788_/Q sky130_fd_sc_hd__dfxtp_4
X_43721_ _87296_/Q _69823_/B sky130_fd_sc_hd__inv_2
X_55707_ _55252_/A _55707_/B _55707_/X sky130_fd_sc_hd__and2_4
X_74541_ _74541_/A _56535_/X _74541_/C _74541_/Y sky130_fd_sc_hd__nand3_4
X_86527_ _86523_/CLK _48389_/Y _72817_/B sky130_fd_sc_hd__dfxtp_4
X_40933_ _82305_/Q _40932_/X _40933_/X sky130_fd_sc_hd__or2_4
X_52919_ _85730_/Q _52902_/X _52918_/Y _52919_/Y sky130_fd_sc_hd__o21ai_4
X_71753_ _71181_/A _71753_/B _71744_/C _71753_/D _71753_/Y sky130_fd_sc_hd__nand4_4
X_59475_ _59462_/X _83458_/Q _59474_/Y _84722_/D sky130_fd_sc_hd__o21a_4
X_83739_ _83736_/CLK _83739_/D _83739_/Q sky130_fd_sc_hd__dfxtp_4
X_56687_ _56671_/X _56685_/X _56686_/X _56687_/X sky130_fd_sc_hd__o21a_4
X_53899_ _85546_/Q _53896_/X _53898_/Y _53899_/Y sky130_fd_sc_hd__o21ai_4
X_46440_ _46435_/Y _46399_/X _46439_/Y _46440_/Y sky130_fd_sc_hd__a21boi_4
X_70704_ _70935_/A _70716_/A sky130_fd_sc_hd__buf_2
X_58426_ _58984_/A _58426_/X sky130_fd_sc_hd__buf_2
X_77260_ _77260_/A _77259_/Y _77260_/Y sky130_fd_sc_hd__nor2_4
X_43652_ _40707_/A _43634_/X _68888_/B _43636_/X _43652_/X sky130_fd_sc_hd__a2bb2o_4
X_55638_ _85057_/Q _55617_/X _55610_/X _55637_/Y _55638_/X sky130_fd_sc_hd__a211o_4
X_86458_ _85555_/CLK _86458_/D _86458_/Q sky130_fd_sc_hd__dfxtp_4
X_74472_ _48609_/A _74478_/B _74478_/C _74472_/X sky130_fd_sc_hd__and3_4
X_40864_ _40864_/A _40883_/B _40864_/X sky130_fd_sc_hd__or2_4
X_71684_ _71682_/Y _83412_/Q _71683_/Y _71684_/X sky130_fd_sc_hd__a21o_4
X_76211_ _76194_/Y _76192_/X _76210_/Y _76211_/Y sky130_fd_sc_hd__a21oi_4
X_42603_ _42603_/A _42603_/Y sky130_fd_sc_hd__inv_2
X_85409_ _85505_/CLK _85409_/D _85409_/Q sky130_fd_sc_hd__dfxtp_4
X_73423_ _44583_/Y _73420_/X _73422_/Y _73434_/C sky130_fd_sc_hd__a21o_4
X_46371_ _46371_/A _46380_/B _46371_/X sky130_fd_sc_hd__or2_4
X_70635_ _70635_/A _70639_/B sky130_fd_sc_hd__buf_2
X_58357_ _58334_/X _61656_/A _58356_/Y _84870_/D sky130_fd_sc_hd__a21oi_4
X_77191_ _82108_/Q _77191_/B _77191_/X sky130_fd_sc_hd__xor2_4
X_43583_ _48144_/A _43583_/Y sky130_fd_sc_hd__inv_2
X_55569_ _56595_/A _55562_/X _56595_/B _55568_/X _55570_/D sky130_fd_sc_hd__and4_4
X_86389_ _83676_/CLK _49430_/Y _58720_/B sky130_fd_sc_hd__dfxtp_4
X_40795_ _40792_/X _40793_/X _88334_/Q _40794_/X _88334_/D sky130_fd_sc_hd__a2bb2o_4
X_48110_ _48110_/A _48086_/B _48110_/X sky130_fd_sc_hd__or2_4
X_45322_ _45277_/X _61649_/B _45294_/X _45322_/Y sky130_fd_sc_hd__o21ai_4
X_57308_ _57306_/Y _57307_/Y _57280_/X _57308_/Y sky130_fd_sc_hd__o21ai_4
X_76142_ _76142_/A _76142_/B _76142_/X sky130_fd_sc_hd__xor2_4
X_88128_ _88128_/CLK _41838_/X _67028_/B sky130_fd_sc_hd__dfxtp_4
X_42534_ _74224_/A _42534_/Y sky130_fd_sc_hd__inv_2
X_73354_ _73257_/X _86186_/Q _73351_/X _73353_/X _73354_/X sky130_fd_sc_hd__a211o_4
X_49090_ _48623_/A _49091_/C sky130_fd_sc_hd__buf_2
X_70566_ DATA_TO_HASH[1] _71887_/A sky130_fd_sc_hd__inv_2
Xclkbuf_7_23_0_CLK clkbuf_7_23_0_CLK/A clkbuf_8_47_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_58288_ _58287_/Y _58280_/B _58288_/Y sky130_fd_sc_hd__nand2_4
X_72305_ _57759_/X _72305_/X sky130_fd_sc_hd__buf_2
X_48041_ _48004_/A _52036_/B _48041_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_163_0_CLK clkbuf_7_81_0_CLK/X clkbuf_9_326_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_45253_ _85162_/Q _45209_/X _45189_/X _45253_/X sky130_fd_sc_hd__o21a_4
X_57239_ _44288_/X _56571_/X _45413_/A _57238_/X _57239_/X sky130_fd_sc_hd__a2bb2o_4
X_76073_ _76073_/A _76073_/B _76074_/B sky130_fd_sc_hd__xnor2_4
X_88059_ _87553_/CLK _42046_/Y _73372_/A sky130_fd_sc_hd__dfxtp_4
X_42465_ _42465_/A _42610_/A sky130_fd_sc_hd__buf_2
X_73285_ _73260_/A _86477_/Q _73285_/X sky130_fd_sc_hd__and2_4
X_70497_ HASH_ADDR[5] _70700_/A sky130_fd_sc_hd__buf_2
X_44204_ _44166_/Y _44204_/Y sky130_fd_sc_hd__inv_2
X_75024_ _80954_/Q _75024_/B _75024_/X sky130_fd_sc_hd__xor2_4
X_79901_ _84922_/Q _65901_/C _80263_/B sky130_fd_sc_hd__nand2_4
X_41416_ _41415_/Y _41416_/X sky130_fd_sc_hd__buf_2
X_60250_ _60170_/A _60218_/A _60324_/B _60367_/C sky130_fd_sc_hd__nand3_4
X_72236_ _72236_/A _72236_/Y sky130_fd_sc_hd__inv_2
X_45184_ _64420_/B _61548_/B sky130_fd_sc_hd__buf_2
X_42396_ _40418_/X _42388_/X _87882_/Q _42389_/X _87882_/D sky130_fd_sc_hd__a2bb2o_4
X_44135_ _44134_/X _44135_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_38_0_CLK clkbuf_7_39_0_CLK/A clkbuf_8_77_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_79832_ _79812_/Y _79852_/B _79831_/X _79832_/Y sky130_fd_sc_hd__a21boi_4
X_41347_ _41346_/X _41347_/X sky130_fd_sc_hd__buf_2
X_72167_ _59292_/X _85341_/Q _59365_/X _72167_/X sky130_fd_sc_hd__o21a_4
X_60181_ _60291_/C _60324_/A sky130_fd_sc_hd__buf_2
X_49992_ _50001_/A _53205_/B _49992_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_178_0_CLK clkbuf_7_89_0_CLK/X clkbuf_8_178_0_CLK/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_173_0_CLK clkbuf_9_86_0_CLK/X _81794_/CLK sky130_fd_sc_hd__clkbuf_1
X_71118_ _70913_/A _71119_/C sky130_fd_sc_hd__buf_2
X_48943_ _71987_/B _48944_/B sky130_fd_sc_hd__buf_2
X_44066_ _44086_/A _44116_/B sky130_fd_sc_hd__buf_2
X_79763_ _84222_/Q _83270_/Q _79763_/X sky130_fd_sc_hd__xor2_4
X_41278_ _41239_/X _41241_/X _41277_/X _69104_/B _41236_/X _41279_/A
+ sky130_fd_sc_hd__o32ai_4
X_72098_ _46259_/A _74391_/A sky130_fd_sc_hd__buf_2
X_76975_ _76975_/A _84399_/Q _76975_/X sky130_fd_sc_hd__xor2_4
X_43017_ _43017_/A _43017_/X sky130_fd_sc_hd__buf_2
X_78714_ _78713_/B _78712_/Y _78709_/Y _78718_/C sky130_fd_sc_hd__o21ai_4
X_63940_ _61922_/X _63876_/B _63905_/C _63892_/D _63940_/Y sky130_fd_sc_hd__nand4_4
X_71049_ _71049_/A _71055_/C sky130_fd_sc_hd__buf_2
X_75926_ _81698_/D _75924_/B _75928_/A sky130_fd_sc_hd__nand2_4
X_48874_ _50069_/A _48874_/B _48874_/X sky130_fd_sc_hd__and2_4
X_79694_ _79678_/X _79682_/B _79694_/X sky130_fd_sc_hd__or2_4
Xclkbuf_9_294_0_CLK clkbuf_9_295_0_CLK/A clkbuf_9_294_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_8_101_0_CLK clkbuf_7_50_0_CLK/X clkbuf_9_203_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_47825_ _47825_/A _48914_/A sky130_fd_sc_hd__buf_2
X_78645_ _82809_/Q _78645_/Y sky130_fd_sc_hd__inv_2
X_63871_ _64305_/B _63920_/B _63840_/C _63920_/D _63871_/Y sky130_fd_sc_hd__nand4_4
X_75857_ _75838_/Y _75840_/B _80926_/Q _80798_/D _75857_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_10_188_0_CLK clkbuf_9_94_0_CLK/X _80719_/CLK sky130_fd_sc_hd__clkbuf_1
X_65610_ _65438_/X _86197_/Q _65576_/X _65609_/X _65610_/X sky130_fd_sc_hd__a211o_4
X_62822_ _61500_/X _62834_/B _62801_/X _62834_/D _62822_/Y sky130_fd_sc_hd__nand4_4
X_74808_ _74723_/X _74808_/B _74745_/D _74810_/C sky130_fd_sc_hd__nand3_4
X_47756_ _81225_/Q _47757_/A sky130_fd_sc_hd__inv_2
X_66590_ _68999_/A _86805_/Q _66590_/X sky130_fd_sc_hd__and2_4
X_78576_ _78575_/X _78600_/A sky130_fd_sc_hd__inv_2
X_44968_ _45734_/A _44968_/X sky130_fd_sc_hd__buf_2
X_75788_ _75771_/A _75784_/A _75788_/Y sky130_fd_sc_hd__nand2_4
X_46707_ _46706_/Y _46707_/X sky130_fd_sc_hd__buf_2
X_65541_ _65474_/X _86522_/Q _65541_/X sky130_fd_sc_hd__and2_4
X_77527_ _77520_/X _77526_/Y _82198_/D sky130_fd_sc_hd__xor2_4
X_43919_ _43918_/Y _87200_/D sky130_fd_sc_hd__inv_2
X_62753_ _62727_/A _62762_/B _61861_/X _62753_/Y sky130_fd_sc_hd__nand3_4
X_74739_ _74716_/A _74739_/B _70732_/X _74739_/Y sky130_fd_sc_hd__nand3_4
X_47687_ _54880_/B _53187_/B sky130_fd_sc_hd__buf_2
X_44899_ _55990_/C _45876_/B _44898_/X _44899_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_8_116_0_CLK clkbuf_7_58_0_CLK/X clkbuf_8_116_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_61704_ _59651_/B _59600_/X _59721_/A _61704_/Y sky130_fd_sc_hd__nand3_4
X_49426_ _49423_/Y _49405_/X _49425_/X _49426_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_111_0_CLK clkbuf_9_55_0_CLK/X _86841_/CLK sky130_fd_sc_hd__clkbuf_1
X_68260_ _68106_/A _68260_/X sky130_fd_sc_hd__buf_2
X_46638_ _46638_/A _51761_/D sky130_fd_sc_hd__buf_2
X_65472_ _65453_/X _85598_/Q _65470_/X _65471_/X _65472_/X sky130_fd_sc_hd__a211o_4
X_77458_ _77454_/X _77458_/B _77458_/X sky130_fd_sc_hd__xor2_4
X_62684_ _62667_/X _62704_/C sky130_fd_sc_hd__buf_2
Xclkbuf_10_741_0_CLK clkbuf_9_370_0_CLK/X _88012_/CLK sky130_fd_sc_hd__clkbuf_1
X_67211_ _66971_/A _67211_/X sky130_fd_sc_hd__buf_2
X_64423_ _64367_/A _64423_/X sky130_fd_sc_hd__buf_2
X_76409_ _76410_/A _81568_/Q _76409_/Y sky130_fd_sc_hd__nor2_4
X_49357_ _86402_/Q _49300_/X _49356_/Y _49357_/Y sky130_fd_sc_hd__o21ai_4
X_61635_ _61633_/X _61576_/X _61634_/Y _61635_/Y sky130_fd_sc_hd__a21oi_4
X_68191_ _68188_/X _67175_/Y _68189_/X _68190_/Y _68191_/X sky130_fd_sc_hd__a211o_4
X_46569_ _51380_/B _54079_/B sky130_fd_sc_hd__buf_2
X_77389_ _77396_/A _77388_/Y _82189_/D sky130_fd_sc_hd__xnor2_4
Xclkbuf_9_232_0_CLK clkbuf_8_116_0_CLK/X clkbuf_9_232_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_48308_ _48275_/X _57609_/B _48308_/Y sky130_fd_sc_hd__nand2_4
X_67142_ _67095_/A _67142_/B _67142_/X sky130_fd_sc_hd__and2_4
X_79128_ _79128_/A _79128_/B _79128_/X sky130_fd_sc_hd__xor2_4
X_64354_ _64344_/X _64307_/B _84829_/Q _64354_/X sky130_fd_sc_hd__and3_4
X_49288_ _65029_/B _49285_/X _49287_/Y _49288_/Y sky130_fd_sc_hd__o21ai_4
X_61566_ _61546_/A _61546_/B _79138_/B _61566_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_10_126_0_CLK clkbuf_9_63_0_CLK/X _84430_/CLK sky130_fd_sc_hd__clkbuf_1
X_63305_ _63528_/A _63305_/X sky130_fd_sc_hd__buf_2
X_48239_ _48229_/A _53516_/B _48239_/Y sky130_fd_sc_hd__nand2_4
X_60517_ _60516_/Y _60517_/Y sky130_fd_sc_hd__inv_2
X_67073_ _67070_/X _67072_/X _67026_/X _67078_/A sky130_fd_sc_hd__a21o_4
X_79059_ _79058_/A _79058_/B _82749_/Q _79059_/X sky130_fd_sc_hd__a21o_4
X_64285_ _64285_/A _64295_/A sky130_fd_sc_hd__buf_2
X_61497_ _61495_/X _61455_/X _61496_/Y _61497_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_756_0_CLK clkbuf_9_378_0_CLK/X _87789_/CLK sky130_fd_sc_hd__clkbuf_1
X_66024_ _65878_/A _66024_/B _66024_/X sky130_fd_sc_hd__and2_4
X_51250_ _64670_/B _51233_/X _51249_/Y _51250_/Y sky130_fd_sc_hd__o21ai_4
X_63236_ _58391_/A _63190_/X _63234_/X _58264_/Y _63235_/X _63236_/Y
+ sky130_fd_sc_hd__o32ai_4
X_82070_ _81154_/CLK _82070_/D _77906_/A sky130_fd_sc_hd__dfxtp_4
X_60448_ _60529_/B _60572_/A sky130_fd_sc_hd__inv_2
Xclkbuf_9_247_0_CLK clkbuf_9_247_0_CLK/A clkbuf_9_247_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_50201_ _51242_/A _50714_/B _50201_/X sky130_fd_sc_hd__and2_4
X_81021_ _85315_/CLK _79836_/A _81021_/Q sky130_fd_sc_hd__dfxtp_4
X_51181_ _51177_/A _51192_/B _51192_/C _52872_/D _51181_/X sky130_fd_sc_hd__and4_4
X_63167_ _63144_/X _64379_/C _63146_/C _63135_/D _63167_/X sky130_fd_sc_hd__and4_4
X_60379_ _60378_/Y _60392_/C sky130_fd_sc_hd__inv_2
X_50132_ _50129_/Y _50117_/X _50131_/X _86258_/D sky130_fd_sc_hd__a21oi_4
X_62118_ _62104_/X _62109_/X _62116_/Y _84872_/Q _62117_/X _62118_/Y
+ sky130_fd_sc_hd__o32ai_4
X_67975_ _68044_/A _67975_/B _67975_/X sky130_fd_sc_hd__and2_4
X_63098_ _63088_/A _64307_/C _63087_/X _63077_/D _63098_/X sky130_fd_sc_hd__and4_4
X_69714_ _44543_/A _69690_/X _69611_/X _69713_/X _69714_/X sky130_fd_sc_hd__a211o_4
X_50063_ _50063_/A _50064_/A sky130_fd_sc_hd__buf_2
X_54940_ _85349_/Q _54918_/X _54939_/Y _54940_/Y sky130_fd_sc_hd__o21ai_4
X_66926_ _67046_/A _66926_/X sky130_fd_sc_hd__buf_2
X_62049_ _62038_/X _62040_/X _62047_/Y _84845_/Q _62048_/X _62049_/Y
+ sky130_fd_sc_hd__o32ai_4
X_85760_ _85761_/CLK _52759_/Y _85760_/Q sky130_fd_sc_hd__dfxtp_4
X_82972_ _83783_/CLK _82780_/Q _82972_/Q sky130_fd_sc_hd__dfxtp_4
X_84711_ _84355_/CLK _59697_/Y _80605_/A sky130_fd_sc_hd__dfxtp_4
X_81923_ _82124_/CLK _81923_/D _81923_/Q sky130_fd_sc_hd__dfxtp_4
X_69645_ _69645_/A _69645_/X sky130_fd_sc_hd__buf_2
X_54871_ _54885_/A _54871_/B _54871_/Y sky130_fd_sc_hd__nand2_4
X_66857_ _66769_/A _66857_/B _66857_/X sky130_fd_sc_hd__and2_4
X_85691_ _85692_/CLK _53134_/Y _85691_/Q sky130_fd_sc_hd__dfxtp_4
X_56610_ _55546_/X _55550_/X _72654_/C sky130_fd_sc_hd__and2_4
X_87430_ _86796_/CLK _43419_/X _87430_/Q sky130_fd_sc_hd__dfxtp_4
X_53822_ _53820_/Y _53799_/X _53821_/Y _53822_/Y sky130_fd_sc_hd__a21boi_4
X_65808_ _65717_/X _85576_/Q _65718_/X _65807_/X _65808_/X sky130_fd_sc_hd__a211o_4
X_84642_ _84645_/CLK _60279_/Y _79806_/A sky130_fd_sc_hd__dfxtp_4
X_57590_ _57564_/X _57590_/B _57590_/Y sky130_fd_sc_hd__nand2_4
X_69576_ _69139_/X _69141_/X _69575_/X _69576_/Y sky130_fd_sc_hd__a21oi_4
X_81854_ _82531_/CLK _81886_/Q _77652_/A sky130_fd_sc_hd__dfxtp_4
X_66788_ _66783_/X _66786_/X _66787_/X _66791_/A sky130_fd_sc_hd__a21o_4
X_56541_ _56164_/X _56462_/X _56540_/Y _56541_/Y sky130_fd_sc_hd__o21ai_4
X_80805_ _80931_/CLK _83949_/Q _75743_/B sky130_fd_sc_hd__dfxtp_4
X_68527_ _69007_/A _68527_/X sky130_fd_sc_hd__buf_2
X_87361_ _86796_/CLK _87361_/D _87361_/Q sky130_fd_sc_hd__dfxtp_4
X_53753_ _53751_/Y _53747_/X _53752_/X _53753_/Y sky130_fd_sc_hd__a21oi_4
X_65739_ _65753_/A _86509_/Q _65739_/X sky130_fd_sc_hd__and2_4
X_84573_ _84583_/CLK _84573_/D _84573_/Q sky130_fd_sc_hd__dfxtp_4
X_50965_ _50819_/X _50965_/X sky130_fd_sc_hd__buf_2
X_81785_ _81475_/CLK _76142_/X _48448_/A sky130_fd_sc_hd__dfxtp_4
X_86312_ _86312_/CLK _86312_/D _58058_/B sky130_fd_sc_hd__dfxtp_4
X_52704_ _52704_/A _52694_/B _52694_/C _52704_/D _52704_/X sky130_fd_sc_hd__and4_4
X_59260_ _59033_/A _59260_/X sky130_fd_sc_hd__buf_2
X_83524_ _83526_/CLK _71364_/X _83524_/Q sky130_fd_sc_hd__dfxtp_4
X_56472_ _56545_/A _56472_/B _85183_/Q _56472_/Y sky130_fd_sc_hd__nand3_4
X_68458_ _68454_/X _68457_/X _68331_/X _68458_/Y sky130_fd_sc_hd__a21oi_4
X_80736_ _81104_/CLK _75922_/X _80704_/D sky130_fd_sc_hd__dfxtp_4
X_87292_ _88062_/CLK _43731_/X _87292_/Q sky130_fd_sc_hd__dfxtp_4
X_53684_ _85588_/Q _53660_/X _53683_/Y _53684_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_709_0_CLK clkbuf_9_354_0_CLK/X _88267_/CLK sky130_fd_sc_hd__clkbuf_1
X_50896_ _51033_/A _50952_/A sky130_fd_sc_hd__buf_2
X_58211_ _58210_/X _58238_/B _58211_/Y sky130_fd_sc_hd__nor2_4
X_55423_ _55422_/Y _55423_/B _55423_/Y sky130_fd_sc_hd__nand2_4
X_67409_ _87472_/Q _67358_/X _67360_/X _67408_/X _67409_/X sky130_fd_sc_hd__a211o_4
X_86243_ _83594_/CLK _50206_/Y _86243_/Q sky130_fd_sc_hd__dfxtp_4
X_52635_ _52643_/A _52654_/B _52643_/C _46716_/X _52635_/X sky130_fd_sc_hd__and4_4
X_59191_ _59182_/Y _59145_/X _59187_/X _59190_/X _84762_/D sky130_fd_sc_hd__a22oi_4
X_83455_ _83457_/CLK _71564_/X _83455_/Q sky130_fd_sc_hd__dfxtp_4
X_80667_ _84531_/CLK _80667_/D _80667_/Q sky130_fd_sc_hd__dfxtp_4
X_68389_ _68389_/A _69678_/A sky130_fd_sc_hd__buf_2
XPHY_403 sky130_fd_sc_hd__decap_3
XPHY_414 sky130_fd_sc_hd__decap_3
X_70420_ _71162_/B _70358_/X _71287_/C _70854_/A sky130_fd_sc_hd__nand3_4
X_58142_ _58140_/X _85986_/Q _58141_/X _58142_/Y sky130_fd_sc_hd__o21ai_4
X_82406_ _82443_/CLK _82438_/Q _78358_/A sky130_fd_sc_hd__dfxtp_4
XPHY_425 sky130_fd_sc_hd__decap_3
X_55354_ _55445_/D _55354_/Y sky130_fd_sc_hd__inv_2
X_86174_ _83307_/CLK _50581_/Y _86174_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_436 sky130_fd_sc_hd__decap_3
X_40580_ _40577_/X _82879_/Q _40579_/X _40581_/A sky130_fd_sc_hd__o21a_4
X_52566_ _52564_/Y _51951_/X _52565_/Y _85796_/D sky130_fd_sc_hd__a21boi_4
X_83386_ _84945_/CLK _83386_/D _83386_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_447 sky130_fd_sc_hd__decap_3
X_80598_ _80598_/A _80598_/B _80598_/C _80598_/X sky130_fd_sc_hd__and3_4
XPHY_458 sky130_fd_sc_hd__decap_3
X_54305_ _54314_/A _46685_/A _54305_/Y sky130_fd_sc_hd__nand2_4
XPHY_469 sky130_fd_sc_hd__decap_3
X_85125_ _85128_/CLK _85125_/D _55207_/A sky130_fd_sc_hd__dfxtp_4
X_51517_ _51515_/Y _51503_/X _51516_/X _85996_/D sky130_fd_sc_hd__a21oi_4
X_58073_ _58030_/X _85479_/Q _58062_/X _58073_/X sky130_fd_sc_hd__o21a_4
X_70351_ _70209_/A _74727_/A _70350_/X _70351_/X sky130_fd_sc_hd__a21o_4
X_82337_ _86758_/CLK _77228_/X _82337_/Q sky130_fd_sc_hd__dfxtp_4
X_55285_ _55285_/A _83318_/Q _55274_/X _55674_/B sky130_fd_sc_hd__nand3_4
X_52497_ _50946_/A _52498_/C sky130_fd_sc_hd__buf_2
X_57024_ _57023_/X _56729_/X _56810_/X _57024_/D _57024_/Y sky130_fd_sc_hd__nand4_4
X_54236_ _54316_/A _54255_/A sky130_fd_sc_hd__buf_2
X_42250_ _41433_/X _42248_/X _87960_/Q _42249_/X _87960_/D sky130_fd_sc_hd__a2bb2o_4
X_73070_ _73239_/A _73070_/B _73070_/X sky130_fd_sc_hd__and2_4
X_85056_ _85152_/CLK _57239_/X _45413_/A sky130_fd_sc_hd__dfxtp_4
X_51448_ _51557_/A _51448_/X sky130_fd_sc_hd__buf_2
X_70282_ _70246_/A _70292_/A sky130_fd_sc_hd__buf_2
X_82268_ _83515_/CLK _82268_/D _82268_/Q sky130_fd_sc_hd__dfxtp_4
X_41201_ _81712_/Q _41197_/B _41201_/X sky130_fd_sc_hd__or2_4
X_72021_ _72019_/Y _72009_/X _72020_/Y _72021_/Y sky130_fd_sc_hd__a21boi_4
X_84007_ _81746_/CLK _68227_/X _84007_/Q sky130_fd_sc_hd__dfxtp_4
X_81219_ _85317_/CLK _81027_/Q _81219_/Q sky130_fd_sc_hd__dfxtp_4
X_42181_ _41250_/X _42161_/X _87994_/Q _42162_/X _42181_/X sky130_fd_sc_hd__a2bb2o_4
X_54167_ _54249_/A _54167_/X sky130_fd_sc_hd__buf_2
X_51379_ _65337_/B _51362_/X _51378_/Y _51379_/Y sky130_fd_sc_hd__o21ai_4
X_82199_ _82390_/CLK _82199_/D _82391_/D sky130_fd_sc_hd__dfxtp_4
X_41132_ _81725_/Q _41102_/B _41132_/X sky130_fd_sc_hd__or2_4
X_53118_ _53133_/A _53113_/B _53133_/C _53118_/D _53118_/X sky130_fd_sc_hd__and4_4
X_54098_ _85504_/Q _53431_/X _54097_/Y _54098_/Y sky130_fd_sc_hd__o21ai_4
X_58975_ _62948_/C _58976_/A sky130_fd_sc_hd__inv_2
X_57926_ _58796_/A _57926_/X sky130_fd_sc_hd__buf_2
X_41063_ _41061_/X _82282_/Q _41062_/X _41064_/A sky130_fd_sc_hd__o21ai_4
X_45940_ _44008_/A _45941_/A sky130_fd_sc_hd__inv_2
X_53049_ _53047_/Y _53028_/X _53048_/X _53049_/Y sky130_fd_sc_hd__a21oi_4
X_76760_ _76746_/Y _76747_/Y _76734_/A _76749_/Y _76760_/X sky130_fd_sc_hd__a2bb2o_4
X_85958_ _85957_/CLK _85958_/D _85958_/Q sky130_fd_sc_hd__dfxtp_4
X_73972_ _72757_/A _73972_/X sky130_fd_sc_hd__buf_2
X_75711_ _75711_/A _75710_/Y _75712_/B sky130_fd_sc_hd__xnor2_4
X_84909_ _84714_/CLK _84909_/D _58201_/A sky130_fd_sc_hd__dfxtp_4
X_72923_ _41996_/Y _72921_/X _72725_/X _72922_/Y _72923_/X sky130_fd_sc_hd__a211o_4
X_45871_ _84994_/Q _45740_/B _45871_/Y sky130_fd_sc_hd__nor2_4
X_57857_ _57806_/X _57857_/B _57857_/Y sky130_fd_sc_hd__nor2_4
X_76691_ _76691_/A _81351_/D _76694_/A sky130_fd_sc_hd__xnor2_4
X_85889_ _85888_/CLK _85889_/D _65423_/B sky130_fd_sc_hd__dfxtp_4
X_47610_ _47610_/A _53148_/B sky130_fd_sc_hd__buf_2
X_78430_ _78450_/C _78429_/Y _82762_/D sky130_fd_sc_hd__xnor2_4
X_44822_ _44807_/X _44821_/X _41666_/X _86936_/Q _44808_/X _44822_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56808_ _56808_/A _56808_/Y sky130_fd_sc_hd__inv_2
X_75642_ _75630_/A _75629_/X _75642_/X sky130_fd_sc_hd__or2_4
X_87628_ _88144_/CLK _42964_/X _87628_/Q sky130_fd_sc_hd__dfxtp_4
X_48590_ _52204_/A _48624_/B _48610_/C _48590_/X sky130_fd_sc_hd__and3_4
X_72854_ _44305_/X _73438_/B sky130_fd_sc_hd__buf_2
X_57788_ _64616_/A _57788_/X sky130_fd_sc_hd__buf_2
X_47541_ _47530_/X _47549_/B _47519_/X _53107_/D _47541_/X sky130_fd_sc_hd__and4_4
X_71805_ _71804_/Y _71805_/X sky130_fd_sc_hd__buf_2
X_59527_ _59602_/C _60175_/A sky130_fd_sc_hd__buf_2
X_78361_ _78343_/Y _82789_/Q _78344_/Y _78361_/Y sky130_fd_sc_hd__a21boi_4
X_44753_ _41298_/A _44665_/X _86973_/Q _44666_/X _86973_/D sky130_fd_sc_hd__a2bb2o_4
X_56739_ _56739_/A _56739_/X sky130_fd_sc_hd__buf_2
X_75573_ _75573_/A _75574_/A _75573_/Y sky130_fd_sc_hd__nand2_4
X_87559_ _87813_/CLK _43145_/Y _73083_/A sky130_fd_sc_hd__dfxtp_4
X_41965_ _41998_/A _41965_/X sky130_fd_sc_hd__buf_2
X_72785_ _73238_/A _72785_/X sky130_fd_sc_hd__buf_2
X_77312_ _77312_/A _77312_/Y sky130_fd_sc_hd__inv_2
X_43704_ _40831_/A _43698_/X _69737_/B _43700_/X _43705_/A sky130_fd_sc_hd__a2bb2o_4
X_74524_ _52803_/B _74517_/X _74523_/Y _74524_/Y sky130_fd_sc_hd__o21ai_4
X_40916_ _40995_/A _40916_/X sky130_fd_sc_hd__buf_2
X_47472_ _47565_/A _47513_/C sky130_fd_sc_hd__buf_2
X_71736_ _71735_/X _71736_/X sky130_fd_sc_hd__buf_2
X_59458_ _59426_/X _59456_/Y _59457_/Y _84727_/D sky130_fd_sc_hd__a21oi_4
X_78292_ _78292_/A _78291_/Y _78293_/B sky130_fd_sc_hd__xor2_4
X_44684_ _87001_/Q _44684_/Y sky130_fd_sc_hd__inv_2
X_41896_ _41895_/Y _41896_/Y sky130_fd_sc_hd__inv_2
X_49211_ _49208_/Y _49189_/X _49210_/Y _49211_/Y sky130_fd_sc_hd__a21oi_4
X_46423_ _47867_/A _46423_/X sky130_fd_sc_hd__buf_2
X_58409_ _58409_/A _58415_/B _58409_/Y sky130_fd_sc_hd__nand2_4
X_77243_ _77241_/Y _77234_/A _77242_/Y _77243_/X sky130_fd_sc_hd__a21bo_4
X_43635_ _87333_/Q _68732_/B sky130_fd_sc_hd__inv_2
X_74455_ _74452_/Y _74430_/X _74454_/X _83063_/D sky130_fd_sc_hd__a21oi_4
X_40847_ _82865_/Q _40847_/B _40847_/X sky130_fd_sc_hd__or2_4
X_71667_ _58530_/Y _71649_/A _71666_/Y _71667_/Y sky130_fd_sc_hd__o21ai_4
X_59389_ _58982_/X _83489_/Q _59388_/Y _59389_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_10_1013_0_CLK clkbuf_9_506_0_CLK/X _83623_/CLK sky130_fd_sc_hd__clkbuf_1
X_73406_ _73238_/A _73406_/X sky130_fd_sc_hd__buf_2
X_49142_ _49137_/Y _49138_/X _49141_/X _86440_/D sky130_fd_sc_hd__a21oi_4
X_61420_ _61429_/A _61419_/X _61429_/C _61420_/Y sky130_fd_sc_hd__nand3_4
X_46354_ _46345_/Y _46346_/X _46353_/Y _86745_/D sky130_fd_sc_hd__a21boi_4
X_70618_ _52995_/B _70583_/X _70617_/Y _83740_/D sky130_fd_sc_hd__o21ai_4
X_77174_ _77173_/B _77174_/B _81920_/Q _77175_/A sky130_fd_sc_hd__nand3_4
X_43566_ _40497_/X _43560_/X _87358_/Q _43561_/X _87358_/D sky130_fd_sc_hd__a2bb2o_4
X_74386_ _74384_/Y _72107_/X _74385_/Y _83077_/D sky130_fd_sc_hd__a21boi_4
X_40778_ _40736_/A _40779_/B sky130_fd_sc_hd__buf_2
X_71598_ _71865_/A _71626_/B _71598_/C _71598_/Y sky130_fd_sc_hd__nor3_4
X_45305_ _83015_/Q _45305_/Y sky130_fd_sc_hd__inv_2
X_76125_ _76110_/X _76124_/Y _76125_/X sky130_fd_sc_hd__or2_4
X_42517_ _42554_/A _42517_/X sky130_fd_sc_hd__buf_2
X_49073_ _53877_/B _49073_/X sky130_fd_sc_hd__buf_2
X_61351_ _61414_/A _61384_/B sky130_fd_sc_hd__buf_2
X_73337_ _48602_/Y _73336_/Y _73337_/X sky130_fd_sc_hd__xor2_4
X_46285_ _46285_/A _46328_/B _46285_/X sky130_fd_sc_hd__or2_4
X_70549_ _71012_/A _70549_/X sky130_fd_sc_hd__buf_2
X_43497_ _43497_/A _43497_/Y sky130_fd_sc_hd__inv_2
X_48024_ _48004_/A _48024_/B _48024_/Y sky130_fd_sc_hd__nand2_4
X_60302_ _60179_/A _60302_/X sky130_fd_sc_hd__buf_2
X_45236_ _45227_/X _45233_/Y _45235_/Y _45236_/Y sky130_fd_sc_hd__a21oi_4
X_76056_ _81717_/D _76056_/B _76063_/C sky130_fd_sc_hd__nand2_4
X_64070_ _63734_/A _64162_/A sky130_fd_sc_hd__buf_2
X_42448_ _42447_/X _52398_/A sky130_fd_sc_hd__buf_2
X_73268_ _48572_/A _73267_/Y _73268_/X sky130_fd_sc_hd__xor2_4
X_61282_ _61281_/X _72507_/A sky130_fd_sc_hd__buf_2
X_75007_ _80952_/Q _75007_/B _75007_/X sky130_fd_sc_hd__xor2_4
X_63021_ _63011_/Y _63012_/X _63014_/X _63017_/X _63020_/X _63021_/Y
+ sky130_fd_sc_hd__o41ai_4
X_60233_ _60189_/A _60239_/A _60233_/Y sky130_fd_sc_hd__nor2_4
X_72219_ _72216_/Y _72218_/Y _72185_/X _72219_/X sky130_fd_sc_hd__a21o_4
X_45167_ _85296_/Q _45120_/X _45153_/X _45167_/X sky130_fd_sc_hd__o21a_4
X_42379_ _42378_/X _42369_/X _41786_/X _87893_/Q _42370_/X _42379_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73199_ _69793_/B _57377_/X _73055_/X _73198_/Y _73199_/X sky130_fd_sc_hd__a211o_4
X_44118_ _44107_/X _44118_/B _44117_/Y _44119_/A sky130_fd_sc_hd__nand3_4
X_79815_ _79807_/A _79807_/B _79814_/Y _79819_/A sky130_fd_sc_hd__a21boi_4
X_60164_ _59830_/Y _60164_/Y sky130_fd_sc_hd__inv_2
X_49975_ _49981_/A _53187_/B _49975_/Y sky130_fd_sc_hd__nand2_4
X_45098_ _45052_/X _61479_/B _45070_/X _45098_/Y sky130_fd_sc_hd__o21ai_4
X_48926_ _48926_/A _48928_/A sky130_fd_sc_hd__buf_2
X_44049_ _44048_/X _44049_/X sky130_fd_sc_hd__buf_2
X_79746_ _79735_/X _79724_/X _79746_/X sky130_fd_sc_hd__and2_4
X_67760_ _84056_/Q _67688_/X _67759_/X _84056_/D sky130_fd_sc_hd__a21bo_4
X_64972_ _64766_/A _64972_/X sky130_fd_sc_hd__buf_2
X_60095_ _60094_/X _60095_/X sky130_fd_sc_hd__buf_2
X_76958_ _76958_/A _76958_/B _76958_/Y sky130_fd_sc_hd__nand2_4
X_66711_ _87949_/Q _66639_/X _66688_/X _66710_/X _66711_/X sky130_fd_sc_hd__a211o_4
X_63923_ _61909_/X _63876_/B _63905_/C _63892_/D _63923_/Y sky130_fd_sc_hd__nand4_4
X_75909_ _75909_/A _62825_/C _80723_/D sky130_fd_sc_hd__xor2_4
X_48857_ _86469_/Q _48836_/X _48856_/Y _48857_/Y sky130_fd_sc_hd__o21ai_4
X_67691_ _67690_/X _67691_/B _67691_/X sky130_fd_sc_hd__and2_4
X_79677_ _79670_/X _79677_/B _79677_/Y sky130_fd_sc_hd__nand2_4
X_76889_ _76901_/A _76889_/B _76889_/X sky130_fd_sc_hd__and2_4
X_69430_ _44245_/A _69430_/X sky130_fd_sc_hd__buf_2
X_47808_ _47808_/A _47809_/A sky130_fd_sc_hd__inv_2
X_66642_ _66642_/A _66642_/X sky130_fd_sc_hd__buf_2
X_78628_ _82808_/Q _78628_/Y sky130_fd_sc_hd__inv_2
X_63854_ _64026_/A _63900_/B sky130_fd_sc_hd__buf_2
X_48788_ _48793_/A _48788_/B _48788_/Y sky130_fd_sc_hd__nand2_4
X_62805_ _62798_/Y _62772_/X _62799_/Y _62802_/Y _62804_/X _62805_/X
+ sky130_fd_sc_hd__a41o_4
X_69361_ _69611_/A _69361_/X sky130_fd_sc_hd__buf_2
X_47739_ _47758_/A _47739_/B _47749_/C _53217_/D _47739_/X sky130_fd_sc_hd__and4_4
X_66573_ _66572_/X _69779_/A sky130_fd_sc_hd__buf_2
X_78559_ _78558_/X _78560_/B sky130_fd_sc_hd__inv_2
X_63785_ _63783_/X _63744_/X _63784_/Y _84295_/D sky130_fd_sc_hd__a21oi_4
X_60997_ _60997_/A _64182_/C sky130_fd_sc_hd__buf_2
X_68312_ _67918_/X _67920_/X _68295_/X _68312_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_680_0_CLK clkbuf_9_340_0_CLK/X _87394_/CLK sky130_fd_sc_hd__clkbuf_1
X_65524_ _65660_/A _65524_/X sky130_fd_sc_hd__buf_2
X_50750_ _50538_/A _50751_/C sky130_fd_sc_hd__buf_2
X_62736_ _62732_/X _62721_/X _62735_/Y _84387_/D sky130_fd_sc_hd__a21oi_4
X_81570_ _81346_/CLK _65901_/C _81570_/Q sky130_fd_sc_hd__dfxtp_4
X_69292_ _87028_/Q _69277_/X _69278_/X _69291_/X _69292_/X sky130_fd_sc_hd__a211o_4
X_49409_ _49404_/Y _49405_/X _49408_/X _86393_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_171_0_CLK clkbuf_8_85_0_CLK/X clkbuf_9_171_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_80521_ _80512_/Y _80513_/A _80520_/X _80522_/B sky130_fd_sc_hd__a21boi_4
X_68243_ _67515_/X _67518_/X _68239_/X _68243_/Y sky130_fd_sc_hd__a21oi_4
X_65455_ _65592_/A _65455_/B _65455_/X sky130_fd_sc_hd__and2_4
X_50681_ _50596_/A _50682_/A sky130_fd_sc_hd__buf_2
X_62667_ _60360_/X _62667_/X sky130_fd_sc_hd__buf_2
X_52420_ _50209_/A _52446_/B _52369_/X _52420_/X sky130_fd_sc_hd__and3_4
X_64406_ _64400_/Y _64401_/X _64403_/X _64405_/Y _64384_/X _64406_/X
+ sky130_fd_sc_hd__o41a_4
X_83240_ _83229_/CLK _72521_/X _79502_/B sky130_fd_sc_hd__dfxtp_4
X_61618_ _59423_/A _61618_/X sky130_fd_sc_hd__buf_2
X_80452_ _80452_/A _80452_/B _80452_/Y sky130_fd_sc_hd__nand2_4
X_68174_ _67086_/X _67088_/X _68173_/X _68174_/Y sky130_fd_sc_hd__a21oi_4
X_65386_ _64725_/A _65387_/A sky130_fd_sc_hd__buf_2
X_62598_ _62620_/A _58296_/A _62532_/X _62600_/C sky130_fd_sc_hd__nand3_4
Xclkbuf_10_695_0_CLK clkbuf_9_347_0_CLK/X _88144_/CLK sky130_fd_sc_hd__clkbuf_1
X_67125_ _67119_/X _67124_/X _67026_/X _67130_/A sky130_fd_sc_hd__a21o_4
X_52351_ _50142_/A _52310_/B _52291_/C _52351_/X sky130_fd_sc_hd__and3_4
X_64337_ _58320_/A _64308_/X _64336_/Y _64337_/Y sky130_fd_sc_hd__o21ai_4
X_83171_ _83161_/CLK _72942_/X _83171_/Q sky130_fd_sc_hd__dfxtp_4
X_61549_ _58382_/A _61549_/X sky130_fd_sc_hd__buf_2
X_80383_ _80372_/X _80383_/B _80384_/D sky130_fd_sc_hd__nand2_4
Xclkbuf_9_186_0_CLK clkbuf_8_93_0_CLK/X clkbuf_9_186_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_51302_ _51298_/A _46407_/A _51302_/X sky130_fd_sc_hd__and2_4
X_82122_ _82485_/CLK _77805_/X _82110_/D sky130_fd_sc_hd__dfxtp_4
X_55070_ _55083_/A _55056_/X _55070_/C _47729_/Y _55070_/X sky130_fd_sc_hd__and4_4
X_67056_ _67055_/X _67056_/X sky130_fd_sc_hd__buf_2
X_52282_ _52278_/Y _52262_/X _52281_/X _52282_/Y sky130_fd_sc_hd__a21oi_4
X_64268_ _64259_/X _64261_/X _64262_/X _64266_/Y _64267_/X _64268_/X
+ sky130_fd_sc_hd__o41a_4
X_54021_ _85521_/Q _54018_/X _54020_/Y _54021_/Y sky130_fd_sc_hd__o21ai_4
X_66007_ _64714_/X _86234_/Q _65904_/X _66006_/X _66007_/X sky130_fd_sc_hd__a211o_4
X_51233_ _50113_/A _51233_/X sky130_fd_sc_hd__buf_2
X_63219_ _60489_/X _63295_/C sky130_fd_sc_hd__buf_2
X_82053_ _82053_/CLK _82053_/D _82053_/Q sky130_fd_sc_hd__dfxtp_4
X_86930_ _86930_/CLK _44831_/X _67654_/B sky130_fd_sc_hd__dfxtp_4
X_64199_ _64508_/A _64490_/B sky130_fd_sc_hd__buf_2
X_81004_ _84210_/CLK _84212_/Q _81004_/Q sky130_fd_sc_hd__dfxtp_4
X_51164_ _51191_/A _51177_/A sky130_fd_sc_hd__buf_2
X_86861_ _86861_/CLK _45687_/Y _63217_/B sky130_fd_sc_hd__dfxtp_4
X_50115_ _50120_/A _49006_/X _50115_/Y sky130_fd_sc_hd__nand2_4
X_85812_ _86422_/CLK _52489_/Y _85812_/Q sky130_fd_sc_hd__dfxtp_4
X_58760_ _58667_/X _86098_/Q _58759_/X _58760_/Y sky130_fd_sc_hd__o21ai_4
X_51095_ _51084_/A _51115_/B _51110_/C _52785_/D _51095_/X sky130_fd_sc_hd__and4_4
X_55972_ _55698_/A _85311_/Q _55972_/X sky130_fd_sc_hd__and2_4
X_67958_ _68644_/A _68025_/A sky130_fd_sc_hd__buf_2
X_86792_ _87086_/CLK _86792_/D _86792_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_633_0_CLK clkbuf_9_316_0_CLK/X _81211_/CLK sky130_fd_sc_hd__clkbuf_1
X_57711_ _57965_/A _57711_/X sky130_fd_sc_hd__buf_2
X_50046_ _50050_/A _50045_/X _51750_/C _53257_/D _50046_/X sky130_fd_sc_hd__and4_4
X_54923_ _54921_/Y _54909_/X _54922_/X _54923_/Y sky130_fd_sc_hd__a21oi_4
X_66909_ _66909_/A _66908_/X _66909_/Y sky130_fd_sc_hd__nand2_4
X_85743_ _85745_/CLK _52854_/Y _85743_/Q sky130_fd_sc_hd__dfxtp_4
X_58691_ _58591_/X _85463_/Q _58690_/X _58691_/Y sky130_fd_sc_hd__o21ai_4
X_82955_ _82769_/CLK _82955_/D _82955_/Q sky130_fd_sc_hd__dfxtp_4
X_67889_ _67817_/X _67889_/B _67889_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_124_0_CLK clkbuf_8_62_0_CLK/X clkbuf_9_124_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_57642_ _71972_/A _48141_/A _57642_/Y sky130_fd_sc_hd__nand2_4
X_81906_ _82131_/CLK _81906_/D _81906_/Q sky130_fd_sc_hd__dfxtp_4
X_69628_ _87067_/Q _44225_/B _57800_/A _69627_/X _69628_/X sky130_fd_sc_hd__a211o_4
X_54854_ _54850_/A _47639_/Y _54854_/Y sky130_fd_sc_hd__nand2_4
X_85674_ _86400_/CLK _53224_/Y _85674_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_51_0_CLK clkbuf_9_51_0_CLK/A clkbuf_9_51_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_82886_ _82886_/CLK _78107_/B _82886_/Q sky130_fd_sc_hd__dfxtp_4
X_87413_ _87926_/CLK _43458_/Y _87413_/Q sky130_fd_sc_hd__dfxtp_4
X_53805_ _53763_/A _53806_/C sky130_fd_sc_hd__buf_2
X_84625_ _81857_/CLK _60352_/X _79629_/A sky130_fd_sc_hd__dfxtp_4
X_57573_ _57570_/Y _57506_/X _57572_/X _84977_/D sky130_fd_sc_hd__a21oi_4
X_69559_ _87008_/Q _44181_/X _69430_/X _69558_/X _69559_/X sky130_fd_sc_hd__a211o_4
X_81837_ _82221_/CLK _81869_/Q _77380_/A sky130_fd_sc_hd__dfxtp_4
X_88393_ _88398_/CLK _40428_/Y _88393_/Q sky130_fd_sc_hd__dfxtp_4
X_54785_ _54758_/A _54790_/A sky130_fd_sc_hd__buf_2
X_51997_ _52027_/A _50293_/B _51997_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_648_0_CLK clkbuf_9_324_0_CLK/X _86930_/CLK sky130_fd_sc_hd__clkbuf_1
X_59312_ _59311_/X _85736_/Q _59263_/X _59312_/X sky130_fd_sc_hd__o21a_4
X_56524_ _56130_/X _56515_/X _56523_/Y _56524_/Y sky130_fd_sc_hd__o21ai_4
X_41750_ _41799_/A _41750_/X sky130_fd_sc_hd__buf_2
X_87344_ _88324_/CLK _87344_/D _87344_/Q sky130_fd_sc_hd__dfxtp_4
X_53736_ _53750_/A _48615_/A _53736_/Y sky130_fd_sc_hd__nand2_4
X_72570_ _72517_/A _72517_/B _72570_/C _72570_/Y sky130_fd_sc_hd__nand3_4
X_84556_ _84590_/CLK _84556_/D _84556_/Q sky130_fd_sc_hd__dfxtp_4
X_50948_ _50963_/A _50941_/B _50948_/C _46728_/X _50948_/X sky130_fd_sc_hd__and4_4
X_81768_ _83133_/CLK _81768_/D _49139_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_139_0_CLK clkbuf_8_69_0_CLK/X clkbuf_9_139_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_40701_ _40698_/X _82861_/Q _40700_/X _40702_/A sky130_fd_sc_hd__o21a_4
X_71521_ _71521_/A _70722_/A _71521_/Y sky130_fd_sc_hd__nand2_4
X_59243_ _59229_/Y _59230_/X _59236_/X _59242_/X _59243_/Y sky130_fd_sc_hd__a22oi_4
X_83507_ _83507_/CLK _71414_/X _83507_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_66_0_CLK clkbuf_9_67_0_CLK/A clkbuf_9_66_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_56455_ _56168_/X _56372_/X _56454_/Y _56455_/Y sky130_fd_sc_hd__o21ai_4
X_80719_ _80719_/CLK _75905_/X _80687_/D sky130_fd_sc_hd__dfxtp_4
X_87275_ _88056_/CLK _43768_/Y _87275_/Q sky130_fd_sc_hd__dfxtp_4
X_41681_ _41680_/Y _41681_/X sky130_fd_sc_hd__buf_2
X_53667_ _50443_/A _53666_/X _53667_/C _53667_/X sky130_fd_sc_hd__and3_4
X_84487_ _84487_/CLK _61363_/Y _84487_/Q sky130_fd_sc_hd__dfxtp_4
X_50879_ _86114_/Q _50820_/X _50878_/Y _50879_/Y sky130_fd_sc_hd__o21ai_4
X_81699_ _84014_/CLK _81699_/D _81699_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_200 sky130_fd_sc_hd__decap_3
X_43420_ _41529_/X _43412_/X _87429_/Q _43413_/X _43420_/X sky130_fd_sc_hd__a2bb2o_4
X_55406_ _56777_/A _55405_/X _55415_/A sky130_fd_sc_hd__nand2_4
X_74240_ _57637_/B _74239_/Y _74241_/B sky130_fd_sc_hd__xor2_4
X_86226_ _85630_/CLK _86226_/D _86226_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_211 sky130_fd_sc_hd__decap_3
X_40632_ _40628_/X _81145_/Q _40631_/X _40632_/Y sky130_fd_sc_hd__o21ai_4
X_52618_ _52618_/A _52619_/A sky130_fd_sc_hd__buf_2
X_59174_ _59115_/X _59172_/Y _59173_/Y _59133_/X _59119_/X _59174_/X
+ sky130_fd_sc_hd__o32a_4
X_71452_ _70679_/A _71626_/C _71450_/C _71452_/Y sky130_fd_sc_hd__nor3_4
X_83438_ _83438_/CLK _83438_/D _83438_/Q sky130_fd_sc_hd__dfxtp_4
X_56386_ _56383_/X _56386_/B _56386_/C _56386_/Y sky130_fd_sc_hd__nand3_4
XPHY_222 sky130_fd_sc_hd__decap_3
X_53598_ _85605_/Q _53586_/X _53597_/Y _53598_/Y sky130_fd_sc_hd__o21ai_4
XPHY_233 sky130_fd_sc_hd__decap_3
XPHY_244 sky130_fd_sc_hd__decap_3
X_58125_ _58846_/A _58125_/X sky130_fd_sc_hd__buf_2
X_70403_ _51389_/B _70364_/A _70402_/Y _70403_/Y sky130_fd_sc_hd__o21ai_4
XPHY_255 sky130_fd_sc_hd__decap_3
X_55337_ _55323_/A _56705_/B _55337_/X sky130_fd_sc_hd__and2_4
X_43351_ _43347_/X _43350_/X _41341_/X _87465_/Q _43330_/X _43352_/A
+ sky130_fd_sc_hd__o32ai_4
X_74171_ _74168_/X _74170_/X _74181_/A sky130_fd_sc_hd__nand2_4
X_86157_ _85837_/CLK _50669_/Y _86157_/Q sky130_fd_sc_hd__dfxtp_4
X_52549_ _51922_/X _52549_/X sky130_fd_sc_hd__buf_2
X_40563_ _41869_/B _42447_/B _41869_/A _42447_/D _40563_/X sky130_fd_sc_hd__and4_4
XPHY_266 sky130_fd_sc_hd__decap_3
X_71383_ _70679_/A _71377_/B _71377_/C _71383_/Y sky130_fd_sc_hd__nor3_4
X_83369_ _83380_/CLK _83369_/D _83369_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_277 sky130_fd_sc_hd__decap_3
XPHY_288 sky130_fd_sc_hd__decap_3
X_42302_ _41586_/X _42290_/X _87931_/Q _42291_/X _87931_/D sky130_fd_sc_hd__a2bb2o_4
X_73122_ _73121_/X _73191_/B _73122_/X sky130_fd_sc_hd__and2_4
X_85108_ _85042_/CLK _85108_/D _45597_/A sky130_fd_sc_hd__dfxtp_4
XPHY_299 sky130_fd_sc_hd__decap_3
X_46070_ _46070_/A _46070_/Y sky130_fd_sc_hd__inv_2
X_58056_ _57989_/X _58054_/Y _58055_/Y _58007_/X _57993_/X _58056_/X
+ sky130_fd_sc_hd__o32a_4
X_70334_ _70320_/X _83794_/Q _70333_/X _83794_/D sky130_fd_sc_hd__a21o_4
X_43282_ _41147_/X _43277_/X _87501_/Q _43278_/X _43282_/X sky130_fd_sc_hd__a2bb2o_4
X_55268_ _45811_/A _55174_/X _55128_/X _55267_/X _55268_/X sky130_fd_sc_hd__a211o_4
X_86088_ _85767_/CLK _51025_/Y _86088_/Q sky130_fd_sc_hd__dfxtp_4
X_40494_ _40494_/A _40494_/Y sky130_fd_sc_hd__inv_2
X_45021_ _45018_/X _45020_/Y _44973_/X _45021_/Y sky130_fd_sc_hd__a21oi_4
X_57007_ _56778_/Y _57007_/X sky130_fd_sc_hd__buf_2
X_42233_ _42232_/Y _87969_/D sky130_fd_sc_hd__inv_2
X_54219_ _54216_/Y _54197_/X _54218_/X _54219_/Y sky130_fd_sc_hd__a21oi_4
X_77930_ _77908_/A _77907_/Y _77920_/A _77919_/Y _77930_/X sky130_fd_sc_hd__o22a_4
X_73053_ _87816_/Q _73053_/B _73053_/Y sky130_fd_sc_hd__nor2_4
X_85039_ _85039_/CLK _57295_/Y _85039_/Q sky130_fd_sc_hd__dfxtp_4
X_70265_ _70267_/A _70267_/B _83178_/Q _70264_/X _70265_/X sky130_fd_sc_hd__and4_4
X_55199_ _55199_/A _55200_/C sky130_fd_sc_hd__buf_2
X_72004_ _83304_/Q _72001_/X _72003_/Y _72004_/Y sky130_fd_sc_hd__o21ai_4
X_42164_ _41203_/X _42161_/X _88002_/Q _42162_/X _88002_/D sky130_fd_sc_hd__a2bb2o_4
X_77861_ _77861_/A _77875_/A _77862_/B sky130_fd_sc_hd__xor2_4
X_70196_ _70200_/A _70200_/B _83201_/Q _70200_/D _70196_/X sky130_fd_sc_hd__and4_4
X_79600_ _79599_/Y _79608_/A sky130_fd_sc_hd__inv_2
X_41115_ _41073_/X _40558_/A _41114_/X _41115_/X sky130_fd_sc_hd__o21a_4
X_76812_ _76812_/A _76811_/Y _76812_/X sky130_fd_sc_hd__xor2_4
X_49760_ _49678_/X _49779_/A sky130_fd_sc_hd__buf_2
X_46972_ _46971_/Y _52779_/D sky130_fd_sc_hd__buf_2
X_42095_ _41881_/A _42096_/A sky130_fd_sc_hd__buf_2
X_58958_ _86690_/Q _58898_/B _58958_/Y sky130_fd_sc_hd__nor2_4
X_77792_ _82153_/Q _77792_/B _77792_/X sky130_fd_sc_hd__xor2_4
X_48711_ _48557_/A _50556_/B _48711_/Y sky130_fd_sc_hd__nand2_4
X_79531_ _65421_/C _83250_/Q _79531_/X sky130_fd_sc_hd__or2_4
X_45923_ _44247_/A _45923_/X sky130_fd_sc_hd__buf_2
X_41046_ _41040_/X _41041_/X _41045_/X _69401_/B _41037_/X _41047_/A
+ sky130_fd_sc_hd__o32ai_4
X_57909_ _58610_/A _57909_/X sky130_fd_sc_hd__buf_2
X_76743_ _76738_/Y _76742_/Y _76743_/Y sky130_fd_sc_hd__nand2_4
X_49691_ _86341_/Q _49687_/X _49690_/Y _49691_/Y sky130_fd_sc_hd__o21ai_4
X_73955_ _73907_/X _84977_/Q _73859_/X _73954_/X _73955_/X sky130_fd_sc_hd__a211o_4
X_58889_ _58877_/X _85928_/Q _58810_/X _58889_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_9_19_0_CLK clkbuf_8_9_0_CLK/X clkbuf_9_19_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_72906_ _73040_/A _65501_/B _72906_/X sky130_fd_sc_hd__and2_4
X_48642_ _48642_/A _48642_/B _48642_/Y sky130_fd_sc_hd__nand2_4
X_60920_ _60920_/A _63761_/A sky130_fd_sc_hd__buf_2
X_79462_ _79442_/Y _79482_/B _79461_/X _79462_/Y sky130_fd_sc_hd__a21boi_4
X_45854_ _85091_/Q _45824_/B _45854_/Y sky130_fd_sc_hd__nor2_4
X_76674_ _76666_/Y _76673_/Y _76674_/X sky130_fd_sc_hd__xor2_4
X_73886_ _47967_/Y _73886_/B _73886_/X sky130_fd_sc_hd__xor2_4
X_78413_ _78413_/A _78412_/Y _78413_/Y sky130_fd_sc_hd__nor2_4
X_44805_ _41453_/Y _46258_/A _86944_/Q _40354_/X _86944_/D sky130_fd_sc_hd__a2bb2o_4
X_75625_ _75625_/A _75625_/Y sky130_fd_sc_hd__inv_2
X_48573_ _48604_/A _48811_/B _48573_/Y sky130_fd_sc_hd__nand2_4
X_60851_ _60162_/A _61287_/A _59716_/B _60851_/X sky130_fd_sc_hd__and3_4
X_72837_ _72806_/X _86206_/Q _72746_/X _72836_/X _72837_/X sky130_fd_sc_hd__a211o_4
X_79393_ _84806_/Q _84126_/Q _79395_/A sky130_fd_sc_hd__xor2_4
X_45785_ _85128_/Q _45709_/X _45743_/X _45785_/X sky130_fd_sc_hd__o21a_4
X_42997_ _42984_/X _42985_/X _40501_/X _67104_/B _42463_/A _42998_/A
+ sky130_fd_sc_hd__o32ai_4
X_47524_ _47619_/A _47524_/X sky130_fd_sc_hd__buf_2
X_78344_ _78344_/A _82661_/D _78344_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_7_0_CLK clkbuf_9_7_0_CLK/A clkbuf_9_7_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_44736_ _44736_/A _44736_/X sky130_fd_sc_hd__buf_2
X_63570_ _58380_/A _63558_/X _61542_/A _63559_/X _63570_/X sky130_fd_sc_hd__a2bb2o_4
X_75556_ _75543_/B _75541_/A _75555_/Y _75557_/B sky130_fd_sc_hd__a21oi_4
X_41948_ _41937_/X _41919_/X _40696_/X _41947_/Y _41939_/X _41948_/Y
+ sky130_fd_sc_hd__o32ai_4
X_72768_ _83177_/Q _72709_/X _72767_/Y _83177_/D sky130_fd_sc_hd__a21o_4
X_60782_ _60686_/X _60689_/Y _60781_/Y _60782_/Y sky130_fd_sc_hd__a21boi_4
X_74507_ _46272_/A _48694_/A _74507_/Y sky130_fd_sc_hd__nand2_4
X_62521_ _64454_/A _60042_/D _62561_/B _62521_/Y sky130_fd_sc_hd__o21ai_4
X_47455_ _54748_/D _53058_/D sky130_fd_sc_hd__buf_2
X_71719_ _70526_/A _71246_/B _70954_/C _71719_/Y sky130_fd_sc_hd__nand3_4
X_78275_ _78262_/A _78262_/B _78275_/Y sky130_fd_sc_hd__nand2_4
X_44667_ _41104_/A _44665_/X _87009_/Q _44666_/X _87009_/D sky130_fd_sc_hd__a2bb2o_4
X_75487_ _75485_/X _75487_/Y sky130_fd_sc_hd__inv_2
X_41879_ _42547_/A _41879_/X sky130_fd_sc_hd__buf_2
X_72699_ _74139_/A _72699_/X sky130_fd_sc_hd__buf_2
X_46406_ _46403_/X _49019_/A _46405_/X _46407_/A sky130_fd_sc_hd__o21ai_4
X_65240_ _65164_/A _86409_/Q _65240_/X sky130_fd_sc_hd__and2_4
X_77226_ _77223_/Y _77225_/Y _77230_/A sky130_fd_sc_hd__nand2_4
X_43618_ _40626_/X _43604_/X _87340_/Q _43607_/X _87340_/D sky130_fd_sc_hd__a2bb2o_4
X_62452_ _62479_/A _63561_/B _62479_/C _62392_/D _62452_/X sky130_fd_sc_hd__and4_4
X_74438_ _83066_/Q _74387_/X _74437_/Y _74438_/Y sky130_fd_sc_hd__o21ai_4
X_47386_ _47385_/Y _53017_/B sky130_fd_sc_hd__buf_2
X_44598_ _87041_/Q _44598_/Y sky130_fd_sc_hd__inv_2
X_49125_ _72077_/B _49125_/X sky130_fd_sc_hd__buf_2
X_61403_ _61334_/A _61403_/X sky130_fd_sc_hd__buf_2
X_46337_ _46337_/A _46328_/B _46337_/X sky130_fd_sc_hd__or2_4
X_65171_ _65167_/Y _65070_/X _65170_/Y _84212_/D sky130_fd_sc_hd__a21o_4
X_77157_ _77157_/A _77157_/B _77157_/Y sky130_fd_sc_hd__nand2_4
X_43549_ _43528_/A _43549_/X sky130_fd_sc_hd__buf_2
X_74369_ _83080_/Q _72066_/X _74368_/Y _74369_/Y sky130_fd_sc_hd__o21ai_4
X_62383_ _62381_/Y _62327_/X _62382_/Y _84414_/D sky130_fd_sc_hd__a21oi_4
X_76108_ _81723_/D _76109_/B _76108_/Y sky130_fd_sc_hd__nand2_4
X_64122_ _64494_/B _64145_/B _64179_/C _64029_/D _64122_/Y sky130_fd_sc_hd__nand4_4
X_49056_ _49056_/A _50649_/B _49056_/Y sky130_fd_sc_hd__nand2_4
X_61334_ _61334_/A _61334_/X sky130_fd_sc_hd__buf_2
X_46268_ _46288_/A _53949_/B _46268_/Y sky130_fd_sc_hd__nand2_4
X_77088_ _77096_/A _77097_/A _77089_/B sky130_fd_sc_hd__xor2_4
X_48007_ _48734_/A _48007_/X sky130_fd_sc_hd__buf_2
X_45219_ _45219_/A _45219_/X sky130_fd_sc_hd__buf_2
X_68930_ _69190_/A _69021_/A sky130_fd_sc_hd__buf_2
X_64053_ _64053_/A _58446_/A _64071_/C _64053_/X sky130_fd_sc_hd__and3_4
X_76039_ _76047_/A _76039_/B _76040_/B sky130_fd_sc_hd__xor2_4
X_61265_ _66518_/B _59771_/X _61265_/C _61265_/X sky130_fd_sc_hd__or3_4
X_46199_ _65464_/A _46199_/X sky130_fd_sc_hd__buf_2
X_63004_ _61323_/A _63004_/B _63004_/C _63252_/B _63004_/X sky130_fd_sc_hd__or4_4
X_60216_ _60193_/A _60217_/A sky130_fd_sc_hd__buf_2
X_68861_ _68746_/A _68861_/B _68861_/Y sky130_fd_sc_hd__nor2_4
X_61196_ _61196_/A _64377_/A sky130_fd_sc_hd__buf_2
X_67812_ _67809_/X _67811_/X _67742_/X _67812_/X sky130_fd_sc_hd__a21o_4
X_60147_ _79907_/B _60148_/C sky130_fd_sc_hd__inv_2
X_49958_ _49973_/A _49943_/B _49973_/C _53170_/D _49958_/X sky130_fd_sc_hd__and4_4
X_68792_ _69442_/A _68792_/X sky130_fd_sc_hd__buf_2
X_48909_ _48902_/Y _48880_/X _48908_/X _86463_/D sky130_fd_sc_hd__a21oi_4
X_67743_ _67738_/X _67741_/X _67742_/X _67743_/X sky130_fd_sc_hd__a21o_4
X_79729_ _79724_/X _79728_/Y _79729_/X sky130_fd_sc_hd__xor2_4
X_64955_ _64817_/X _86132_/Q _64927_/X _64954_/X _64955_/X sky130_fd_sc_hd__a211o_4
X_60078_ _60359_/A _60078_/X sky130_fd_sc_hd__buf_2
X_49889_ _49893_/A _49893_/B _49893_/C _53103_/D _49889_/X sky130_fd_sc_hd__and4_4
X_51920_ _51917_/Y _51904_/X _51919_/X _51920_/Y sky130_fd_sc_hd__a21oi_4
X_63906_ _64067_/A _63908_/B sky130_fd_sc_hd__buf_2
X_82740_ _82740_/CLK _66433_/C _78975_/A sky130_fd_sc_hd__dfxtp_4
X_67674_ _67674_/A _67673_/X _67674_/Y sky130_fd_sc_hd__nand2_4
X_64886_ _64836_/A _86455_/Q _64886_/X sky130_fd_sc_hd__and2_4
X_69413_ _69410_/X _69412_/X _69346_/X _69413_/X sky130_fd_sc_hd__a21o_4
X_66625_ _66625_/A _66651_/A sky130_fd_sc_hd__buf_2
X_51851_ _51851_/A _51851_/B _51851_/C _46791_/X _51851_/X sky130_fd_sc_hd__and4_4
X_63837_ _60996_/B _63900_/C sky130_fd_sc_hd__buf_2
X_82671_ _82671_/CLK _82671_/D _78173_/A sky130_fd_sc_hd__dfxtp_4
X_84410_ _84409_/CLK _84410_/D _62442_/C sky130_fd_sc_hd__dfxtp_4
X_50802_ _50802_/A _50751_/B _50751_/C _50802_/X sky130_fd_sc_hd__and3_4
X_81622_ _81689_/CLK _76449_/B _81622_/Q sky130_fd_sc_hd__dfxtp_4
X_69344_ _69305_/A _87268_/Q _69344_/X sky130_fd_sc_hd__and2_4
X_54570_ _85418_/Q _54567_/X _54569_/Y _54570_/Y sky130_fd_sc_hd__o21ai_4
X_85390_ _85485_/CLK _54722_/Y _85390_/Q sky130_fd_sc_hd__dfxtp_4
X_66556_ _66647_/A _69853_/A sky130_fd_sc_hd__buf_2
X_51782_ _51794_/A _51782_/B _51794_/C _50919_/D _51782_/X sky130_fd_sc_hd__and4_4
X_63768_ _63849_/A _63800_/B sky130_fd_sc_hd__buf_2
X_53521_ _53519_/Y _53498_/X _53520_/Y _85621_/D sky130_fd_sc_hd__a21boi_4
X_65507_ _65502_/X _65506_/X _65389_/X _65507_/X sky130_fd_sc_hd__a21o_4
X_84341_ _84877_/CLK _63246_/X _79301_/A sky130_fd_sc_hd__dfxtp_4
X_50733_ _50738_/A _49212_/B _50733_/Y sky130_fd_sc_hd__nand2_4
X_62719_ _62712_/Y _62713_/X _62715_/Y _62716_/Y _62718_/X _62719_/X
+ sky130_fd_sc_hd__a41o_4
X_81553_ _80912_/CLK _76790_/X _81553_/Q sky130_fd_sc_hd__dfxtp_4
X_69275_ _87529_/Q _69261_/X _69248_/X _69274_/X _69275_/X sky130_fd_sc_hd__a211o_4
X_66487_ _65238_/X _66476_/B _65241_/X _66487_/Y sky130_fd_sc_hd__nand3_4
X_63699_ _58364_/A _63416_/A _63661_/C _63699_/D _63699_/Y sky130_fd_sc_hd__nand4_4
X_56240_ _56250_/A _56243_/B _85263_/Q _56240_/Y sky130_fd_sc_hd__nand3_4
X_80504_ _59143_/Y _66092_/C _80503_/Y _80504_/X sky130_fd_sc_hd__o21a_4
X_68226_ _68221_/X _67387_/Y _68207_/X _68225_/Y _68226_/X sky130_fd_sc_hd__a211o_4
X_87060_ _87063_/CLK _87060_/D _44543_/A sky130_fd_sc_hd__dfxtp_4
X_53452_ _54919_/A _53460_/A sky130_fd_sc_hd__buf_2
X_65438_ _58876_/A _65438_/X sky130_fd_sc_hd__buf_2
X_84272_ _84269_/CLK _84272_/D _64130_/C sky130_fd_sc_hd__dfxtp_4
X_50664_ _50640_/A _53879_/B _50664_/Y sky130_fd_sc_hd__nand2_4
X_81484_ _81431_/CLK _84052_/Q _76734_/A sky130_fd_sc_hd__dfxtp_4
X_86011_ _85725_/CLK _86011_/D _86011_/Q sky130_fd_sc_hd__dfxtp_4
X_52403_ _52385_/A _49163_/A _52403_/X sky130_fd_sc_hd__and2_4
X_83223_ _82272_/CLK _72596_/X _79321_/B sky130_fd_sc_hd__dfxtp_4
X_80435_ _80448_/B _80448_/A _80435_/X sky130_fd_sc_hd__xor2_4
X_56171_ _56171_/A _45904_/X _56171_/C _56172_/A sky130_fd_sc_hd__nand3_4
X_68157_ _68155_/X _66980_/Y _68148_/X _68156_/Y _68157_/X sky130_fd_sc_hd__a211o_4
X_53383_ _53357_/A _53388_/C sky130_fd_sc_hd__buf_2
X_65369_ _65366_/X _65340_/X _65368_/X _65369_/Y sky130_fd_sc_hd__nand3_4
X_50595_ _50595_/A _50596_/A sky130_fd_sc_hd__buf_2
X_55122_ _44305_/X _73195_/A sky130_fd_sc_hd__buf_2
X_67108_ _87357_/Q _67035_/X _67106_/X _67107_/X _67108_/X sky130_fd_sc_hd__a211o_4
X_52334_ _52334_/A _49025_/X _52334_/Y sky130_fd_sc_hd__nand2_4
X_83154_ _86534_/CLK _83154_/D _83154_/Q sky130_fd_sc_hd__dfxtp_4
X_80366_ _80366_/A _80366_/B _80366_/X sky130_fd_sc_hd__xor2_4
X_68088_ _67495_/X _68088_/X sky130_fd_sc_hd__buf_2
X_82105_ _82015_/CLK _82105_/D _82105_/Q sky130_fd_sc_hd__dfxtp_4
X_55053_ _55049_/Y _55050_/X _55052_/X _85328_/D sky130_fd_sc_hd__a21oi_4
X_59930_ _62196_/A _59931_/A sky130_fd_sc_hd__buf_2
X_67039_ _46210_/A _67039_/X sky130_fd_sc_hd__buf_2
X_52265_ _52250_/A _48889_/B _52265_/Y sky130_fd_sc_hd__nand2_4
X_83085_ _83184_/CLK _74356_/X _83085_/Q sky130_fd_sc_hd__dfxtp_4
X_87962_ _87221_/CLK _87962_/D _87962_/Q sky130_fd_sc_hd__dfxtp_4
X_80297_ _80297_/A _80297_/B _80298_/A sky130_fd_sc_hd__nand2_4
X_54004_ _53991_/A _52484_/B _54004_/Y sky130_fd_sc_hd__nand2_4
X_51216_ _51212_/A _47195_/X _51216_/Y sky130_fd_sc_hd__nand2_4
X_86913_ _86914_/CLK _86913_/D _68054_/B sky130_fd_sc_hd__dfxtp_4
X_82036_ _82009_/CLK _82036_/D _82036_/Q sky130_fd_sc_hd__dfxtp_4
X_70050_ _70040_/X _69813_/Y _70033_/X _70049_/Y _70050_/X sky130_fd_sc_hd__a211o_4
X_59861_ _59745_/X _59768_/Y _59858_/Y _59859_/Y _59860_/Y _59861_/Y
+ sky130_fd_sc_hd__a41oi_4
X_52196_ _52210_/A _48811_/B _52196_/Y sky130_fd_sc_hd__nand2_4
X_87893_ _87636_/CLK _87893_/D _87893_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_572_0_CLK clkbuf_9_286_0_CLK/X _87865_/CLK sky130_fd_sc_hd__clkbuf_1
X_58812_ _58703_/X _85454_/Q _58811_/X _58812_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_6_63_0_CLK clkbuf_6_63_0_CLK/A clkbuf_6_63_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_51147_ _51147_/A _51147_/X sky130_fd_sc_hd__buf_2
X_86844_ _81084_/CLK _86844_/D _45889_/A sky130_fd_sc_hd__dfxtp_4
X_59792_ _59791_/X _84700_/D sky130_fd_sc_hd__inv_2
X_58743_ _58714_/X _85779_/Q _58716_/X _58743_/X sky130_fd_sc_hd__o21a_4
X_51078_ _51056_/A _51071_/B _51071_/C _52771_/D _51078_/X sky130_fd_sc_hd__and4_4
X_55955_ _55954_/X _56003_/B sky130_fd_sc_hd__buf_2
X_86775_ _82886_/CLK _86775_/D _86775_/Q sky130_fd_sc_hd__dfxtp_4
X_83987_ _83987_/CLK _68307_/X _82635_/D sky130_fd_sc_hd__dfxtp_4
X_42920_ _42962_/A _42920_/X sky130_fd_sc_hd__buf_2
X_50029_ _40595_/X _50029_/X sky130_fd_sc_hd__buf_2
X_54906_ _54904_/Y _54882_/X _54905_/X _54906_/Y sky130_fd_sc_hd__a21oi_4
X_73740_ _73614_/A _73740_/X sky130_fd_sc_hd__buf_2
X_85726_ _85727_/CLK _85726_/D _85726_/Q sky130_fd_sc_hd__dfxtp_4
X_70952_ _70947_/A _70952_/B _70954_/C _70952_/Y sky130_fd_sc_hd__nand3_4
X_58674_ _58663_/Y _58624_/X _58670_/X _58673_/X _84809_/D sky130_fd_sc_hd__a22oi_4
X_82938_ _81190_/CLK _78311_/Y _46337_/A sky130_fd_sc_hd__dfxtp_4
X_55886_ _85206_/Q _55531_/X _55610_/A _55885_/X _55886_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_587_0_CLK clkbuf_9_293_0_CLK/X _80968_/CLK sky130_fd_sc_hd__clkbuf_1
X_57625_ _57630_/A _53593_/B _57625_/Y sky130_fd_sc_hd__nand2_4
X_54837_ _54857_/A _54843_/B _54857_/C _53144_/D _54837_/X sky130_fd_sc_hd__and4_4
X_42851_ _42850_/Y _42851_/Y sky130_fd_sc_hd__inv_2
X_73671_ _73669_/X _73655_/X _73658_/Y _73671_/Y sky130_fd_sc_hd__nand3_4
X_85657_ _85433_/CLK _85657_/D _85657_/Q sky130_fd_sc_hd__dfxtp_4
X_70883_ _70882_/Y _70884_/B sky130_fd_sc_hd__buf_2
X_82869_ _82349_/CLK _78213_/B _82869_/Q sky130_fd_sc_hd__dfxtp_4
X_75410_ _75411_/A _80965_/Q _75413_/B sky130_fd_sc_hd__nor2_4
X_41802_ _41802_/A _41802_/X sky130_fd_sc_hd__buf_2
X_72622_ _79198_/B _72590_/X _72621_/Y _72612_/X _72622_/X sky130_fd_sc_hd__o22a_4
X_84608_ _83218_/CLK _60514_/X _79148_/A sky130_fd_sc_hd__dfxtp_4
X_45570_ _44891_/X _45570_/X sky130_fd_sc_hd__buf_2
X_57556_ _57597_/A _50300_/B _57556_/Y sky130_fd_sc_hd__nand2_4
X_76390_ _81266_/Q _81522_/D _76390_/Y sky130_fd_sc_hd__nand2_4
X_88376_ _88376_/CLK _88376_/D _88376_/Q sky130_fd_sc_hd__dfxtp_4
X_42782_ _42774_/X _42775_/X _41341_/X _87721_/Q _42781_/X _42782_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54768_ _54758_/X _47490_/A _54768_/Y sky130_fd_sc_hd__nand2_4
X_85588_ _83068_/CLK _85588_/D _85588_/Q sky130_fd_sc_hd__dfxtp_4
X_44521_ _44512_/X _44513_/X _40776_/A _44520_/Y _44516_/X _44521_/Y
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_10_510_0_CLK clkbuf_9_255_0_CLK/X _82768_/CLK sky130_fd_sc_hd__clkbuf_1
X_56507_ _56510_/A _56507_/B _55833_/B _56507_/Y sky130_fd_sc_hd__nand3_4
X_75341_ _75341_/A _75364_/A sky130_fd_sc_hd__inv_2
X_41733_ _82893_/Q _41653_/X _41733_/X sky130_fd_sc_hd__or2_4
X_87327_ _87850_/CLK _87327_/D _87327_/Q sky130_fd_sc_hd__dfxtp_4
X_53719_ _85581_/Q _53687_/X _53718_/Y _53719_/Y sky130_fd_sc_hd__o21ai_4
X_72553_ _72552_/X _83235_/D sky130_fd_sc_hd__inv_2
X_84539_ _84534_/CLK _84539_/D _76987_/A sky130_fd_sc_hd__dfxtp_4
X_57487_ _56927_/A _57440_/A _56927_/C _57487_/X sky130_fd_sc_hd__and3_4
X_54699_ _54616_/X _54699_/X sky130_fd_sc_hd__buf_2
X_47240_ _47382_/A _47240_/X sky130_fd_sc_hd__buf_2
X_59226_ _59226_/A _59226_/B _59226_/Y sky130_fd_sc_hd__nor2_4
X_71504_ _71500_/A _71261_/B _71504_/C _71504_/Y sky130_fd_sc_hd__nand3_4
X_78060_ _84565_/Q _78060_/B _78060_/X sky130_fd_sc_hd__xor2_4
X_56438_ _56134_/X _56426_/X _56437_/Y _85194_/D sky130_fd_sc_hd__o21ai_4
X_44452_ _46298_/A _44602_/A sky130_fd_sc_hd__buf_2
X_75272_ _75268_/Y _75270_/Y _75267_/Y _75272_/Y sky130_fd_sc_hd__o21ai_4
X_87258_ _87776_/CLK _43806_/Y _87258_/Q sky130_fd_sc_hd__dfxtp_4
X_41664_ _41663_/X _41638_/X _67482_/B _41639_/X _88173_/D sky130_fd_sc_hd__a2bb2o_4
X_72484_ _72484_/A _72484_/X sky130_fd_sc_hd__buf_2
X_77011_ _77019_/A _77011_/B _77015_/A sky130_fd_sc_hd__nor2_4
X_43403_ _41485_/X _43396_/X _87438_/Q _43397_/X _43403_/X sky130_fd_sc_hd__a2bb2o_4
X_74223_ _70130_/A _74139_/X _74222_/Y _83117_/D sky130_fd_sc_hd__a21o_4
X_86209_ _85599_/CLK _86209_/D _86209_/Q sky130_fd_sc_hd__dfxtp_4
X_40615_ _40615_/A _40588_/B _40615_/X sky130_fd_sc_hd__or2_4
X_47171_ _47152_/X _47133_/B _47143_/C _52895_/D _47171_/X sky130_fd_sc_hd__and4_4
X_59157_ _59152_/X _59154_/Y _59155_/Y _58943_/X _59156_/X _59157_/X
+ sky130_fd_sc_hd__o32a_4
X_71435_ _71432_/A _71435_/B _71435_/C _71432_/D _71435_/X sky130_fd_sc_hd__and4_4
X_44383_ _44352_/X _44383_/X sky130_fd_sc_hd__buf_2
X_56369_ _56367_/Y _56368_/Y _85218_/D sky130_fd_sc_hd__nand2_4
X_87189_ _87189_/CLK _43938_/X _68044_/B sky130_fd_sc_hd__dfxtp_4
X_41595_ _41344_/X _81159_/Q _41594_/X _41595_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_10_525_0_CLK clkbuf_9_262_0_CLK/X _81344_/CLK sky130_fd_sc_hd__clkbuf_1
X_46122_ _46162_/B _46120_/Y _46121_/Y _46108_/D _45909_/X _46122_/Y
+ sky130_fd_sc_hd__a41oi_4
X_58108_ _58108_/A _58108_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_6_16_0_CLK clkbuf_5_8_0_CLK/X clkbuf_6_16_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_43334_ _41288_/X _43325_/X _87475_/Q _43326_/X _87475_/D sky130_fd_sc_hd__a2bb2o_4
X_74154_ _74151_/X _74153_/X _74085_/X _74154_/X sky130_fd_sc_hd__a21o_4
X_40546_ _40546_/A _40467_/B _40546_/X sky130_fd_sc_hd__or2_4
X_59088_ _59083_/Y _59087_/Y _58939_/X _59088_/X sky130_fd_sc_hd__a21o_4
X_71366_ _71366_/A _70939_/A _70790_/A _71365_/X _71366_/X sky130_fd_sc_hd__and4_4
X_73105_ _69740_/B _72731_/X _56548_/X _73105_/Y sky130_fd_sc_hd__o21ai_4
X_58039_ _86634_/Q _58039_/B _58039_/Y sky130_fd_sc_hd__nor2_4
X_70317_ _70317_/A _70317_/Y sky130_fd_sc_hd__inv_2
X_46053_ _41529_/A _46043_/X _86792_/Q _46044_/X _86792_/D sky130_fd_sc_hd__a2bb2o_4
X_43265_ _43218_/A _43265_/X sky130_fd_sc_hd__buf_2
X_78962_ _78948_/Y _79115_/A _78962_/Y sky130_fd_sc_hd__nor2_4
X_74085_ _72877_/A _74085_/X sky130_fd_sc_hd__buf_2
X_40477_ _44733_/A _40477_/X sky130_fd_sc_hd__buf_2
X_71297_ _70809_/A _71297_/X sky130_fd_sc_hd__buf_2
X_45004_ _45153_/A _45004_/X sky130_fd_sc_hd__buf_2
X_42216_ _42205_/X _42200_/X _41347_/X _87976_/Q _42201_/X _42217_/A
+ sky130_fd_sc_hd__o32ai_4
X_61050_ _60961_/X _60911_/X _60993_/Y _60972_/X _61049_/X _61050_/X
+ sky130_fd_sc_hd__o41a_4
X_77913_ _77899_/Y _77900_/Y _82068_/Q _81940_/D _77913_/X sky130_fd_sc_hd__a2bb2o_4
X_73036_ _73036_/A _73372_/B _73036_/Y sky130_fd_sc_hd__nor2_4
X_70248_ _70247_/X _70260_/B sky130_fd_sc_hd__buf_2
X_43196_ _43162_/A _43196_/X sky130_fd_sc_hd__buf_2
X_78893_ _78881_/A _78888_/A _78893_/X sky130_fd_sc_hd__and2_4
Xclkbuf_2_1_0_CLK clkbuf_2_1_0_CLK/A clkbuf_2_1_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_60001_ _59998_/Y _60000_/Y _59969_/X _80195_/A _59814_/X _84676_/D
+ sky130_fd_sc_hd__o32a_4
X_49812_ _49810_/Y _49787_/X _49811_/X _49812_/Y sky130_fd_sc_hd__a21oi_4
X_42147_ _41157_/X _42137_/X _88011_/Q _42138_/X _88011_/D sky130_fd_sc_hd__a2bb2o_4
X_77844_ _82063_/Q _77844_/Y sky130_fd_sc_hd__inv_2
X_70179_ _70169_/X _83847_/Q _70178_/X _83847_/D sky130_fd_sc_hd__a21o_4
X_49743_ _49688_/X _49757_/A sky130_fd_sc_hd__buf_2
X_46955_ _46767_/A _46955_/X sky130_fd_sc_hd__buf_2
X_42078_ _42025_/A _42078_/X sky130_fd_sc_hd__buf_2
X_77775_ _82264_/Q _77775_/B _81928_/D sky130_fd_sc_hd__xor2_4
X_74987_ _74987_/A _74987_/B _74987_/C _74988_/B sky130_fd_sc_hd__and3_4
X_79514_ _84817_/Q _66364_/C _79517_/A sky130_fd_sc_hd__xor2_4
X_45906_ _42447_/B _45884_/A _46159_/A _45905_/X _45907_/A sky130_fd_sc_hd__a211o_4
X_41029_ _41028_/X _40987_/X _69362_/B _40989_/X _41029_/X sky130_fd_sc_hd__a2bb2o_4
X_64740_ _79836_/A _64741_/C sky130_fd_sc_hd__inv_2
X_76726_ _76726_/A _81450_/D _76726_/X sky130_fd_sc_hd__xor2_4
X_49674_ _49672_/Y _49650_/X _49673_/X _49674_/Y sky130_fd_sc_hd__a21oi_4
X_61952_ _61500_/X _61933_/X _61907_/C _61952_/D _61952_/Y sky130_fd_sc_hd__nand4_4
X_73938_ _70114_/Y _73818_/X _73937_/Y _83130_/D sky130_fd_sc_hd__o21ai_4
X_46886_ _46886_/A _52732_/B sky130_fd_sc_hd__inv_2
X_48625_ _48617_/Y _48585_/X _48624_/X _86506_/D sky130_fd_sc_hd__a21oi_4
X_60903_ _60895_/X _60901_/X _60902_/Y _84552_/Q _60898_/X _84552_/D
+ sky130_fd_sc_hd__o32a_4
X_79445_ _58653_/Y _66402_/C _79444_/Y _79449_/A sky130_fd_sc_hd__o21a_4
X_45837_ _45819_/X _61666_/A _45836_/X _45837_/Y sky130_fd_sc_hd__o21ai_4
X_64671_ _64615_/X _85534_/Q _64642_/X _64670_/X _64671_/X sky130_fd_sc_hd__a211o_4
X_76657_ _76656_/B _76657_/Y sky130_fd_sc_hd__inv_2
X_61883_ _61880_/Y _61881_/X _61882_/Y _61883_/Y sky130_fd_sc_hd__a21oi_4
X_73869_ _72852_/X _73869_/X sky130_fd_sc_hd__buf_2
X_66410_ _66410_/A _66411_/A sky130_fd_sc_hd__buf_2
X_63622_ _63615_/A _63615_/B _80400_/B _63622_/Y sky130_fd_sc_hd__nor3_4
X_75608_ _75607_/B _75891_/A _75608_/Y sky130_fd_sc_hd__nor2_4
X_48556_ _48801_/B _52188_/B sky130_fd_sc_hd__buf_2
X_60834_ _63426_/A _60834_/X sky130_fd_sc_hd__buf_2
X_67390_ _67863_/A _67390_/X sky130_fd_sc_hd__buf_2
X_79376_ _79365_/X _79354_/X _79376_/X sky130_fd_sc_hd__and2_4
X_45768_ _57039_/A _45768_/Y sky130_fd_sc_hd__inv_2
X_76588_ _76586_/X _76560_/Y _76587_/X _76588_/X sky130_fd_sc_hd__and3_4
X_47507_ _47517_/A _53086_/B _47507_/Y sky130_fd_sc_hd__nand2_4
X_66341_ _66338_/X _66385_/B _66340_/X _66341_/Y sky130_fd_sc_hd__nand3_4
X_78327_ _82499_/Q _82755_/D _82467_/D sky130_fd_sc_hd__xor2_4
X_44719_ _44719_/A _44719_/Y sky130_fd_sc_hd__inv_2
X_63553_ _63495_/X _63546_/X _63547_/X _63551_/X _63552_/Y _63553_/Y
+ sky130_fd_sc_hd__o41ai_4
X_75539_ _75503_/Y _75524_/Y _75523_/X _75539_/X sky130_fd_sc_hd__a21bo_4
X_60765_ _60714_/Y _60671_/C _60765_/Y sky130_fd_sc_hd__nand2_4
X_48487_ _48487_/A _52156_/A sky130_fd_sc_hd__buf_2
X_45699_ _63227_/B _61561_/A sky130_fd_sc_hd__buf_2
X_62504_ _62504_/A _62504_/X sky130_fd_sc_hd__buf_2
X_69060_ _86979_/Q _69058_/X _68993_/X _69059_/X _69060_/X sky130_fd_sc_hd__a211o_4
X_47438_ _81803_/Q _54739_/D sky130_fd_sc_hd__inv_2
X_66272_ _66269_/X _66271_/X _66240_/X _66272_/X sky130_fd_sc_hd__a21o_4
X_78258_ _78265_/A _82467_/Q _78263_/A sky130_fd_sc_hd__xor2_4
X_63484_ _63484_/A _63496_/A sky130_fd_sc_hd__buf_2
X_60696_ _60724_/A _60624_/X _60659_/A _60696_/Y sky130_fd_sc_hd__nand3_4
X_68011_ _68008_/X _68010_/X _67917_/X _68011_/X sky130_fd_sc_hd__a21o_4
X_65223_ _64565_/A _65400_/A sky130_fd_sc_hd__buf_2
X_77209_ _77217_/A _77217_/B _77213_/A sky130_fd_sc_hd__xnor2_4
X_62435_ _62406_/A _62435_/B _62432_/Y _62435_/D _62435_/Y sky130_fd_sc_hd__nand4_4
X_47369_ _47369_/A _53008_/D sky130_fd_sc_hd__buf_2
X_78189_ _82673_/Q _78189_/B _78189_/X sky130_fd_sc_hd__xor2_4
X_49108_ _49117_/A _50674_/B _49108_/Y sky130_fd_sc_hd__nand2_4
X_80220_ _80197_/Y _80220_/B _80221_/A sky130_fd_sc_hd__nor2_4
X_65154_ _65154_/A _65153_/X _65154_/Y sky130_fd_sc_hd__nand2_4
X_50380_ _50227_/A _50380_/X sky130_fd_sc_hd__buf_2
X_62366_ _61447_/B _62278_/X _62363_/X _62323_/X _62365_/X _62366_/X
+ sky130_fd_sc_hd__a41o_4
X_64105_ _61611_/A _60967_/X _64104_/Y _64105_/X sky130_fd_sc_hd__a21bo_4
X_49039_ _49039_/A _49029_/B _49039_/Y sky130_fd_sc_hd__nor2_4
X_80151_ _80143_/X _80144_/X _80150_/Y _80151_/Y sky130_fd_sc_hd__a21boi_4
X_61317_ _61317_/A _61317_/X sky130_fd_sc_hd__buf_2
X_65085_ _65059_/X _85551_/Q _65060_/X _65084_/X _65085_/X sky130_fd_sc_hd__a211o_4
X_69962_ _87041_/Q _44181_/X _64600_/A _69961_/X _69962_/X sky130_fd_sc_hd__a211o_4
X_62297_ _62522_/B _62309_/C sky130_fd_sc_hd__buf_2
X_52050_ _52050_/A _52098_/B _52033_/X _52050_/X sky130_fd_sc_hd__and3_4
X_64036_ _64031_/X _63969_/X _64033_/Y _64034_/Y _64035_/X _64036_/X
+ sky130_fd_sc_hd__a41o_4
X_68913_ _69004_/A _88349_/Q _68913_/X sky130_fd_sc_hd__and2_4
X_61248_ _63053_/A _63004_/B sky130_fd_sc_hd__buf_2
X_80082_ _80082_/A _80082_/B _80088_/B sky130_fd_sc_hd__xor2_4
X_69893_ _83889_/Q _69831_/X _69892_/X _83889_/D sky130_fd_sc_hd__a21bo_4
X_51001_ _51018_/A _50985_/B _50985_/C _52694_/D _51001_/X sky130_fd_sc_hd__and4_4
X_83910_ _83906_/CLK _69616_/X _83910_/Q sky130_fd_sc_hd__dfxtp_4
X_68844_ _69004_/A _88352_/Q _68844_/X sky130_fd_sc_hd__and2_4
X_61179_ _61179_/A _61120_/Y _61180_/A sky130_fd_sc_hd__nor2_4
X_84890_ _84921_/CLK _84890_/D _84890_/Q sky130_fd_sc_hd__dfxtp_4
X_83841_ _83835_/CLK _70197_/X _83841_/Q sky130_fd_sc_hd__dfxtp_4
X_68775_ _68938_/A _68775_/B _68775_/X sky130_fd_sc_hd__and2_4
X_65987_ _65757_/A _65987_/X sky130_fd_sc_hd__buf_2
X_55740_ _55737_/X _55739_/X _55740_/Y sky130_fd_sc_hd__nand2_4
X_67726_ _67726_/A _67725_/X _67726_/Y sky130_fd_sc_hd__nand2_4
X_86560_ _86560_/CLK _48180_/Y _73588_/B sky130_fd_sc_hd__dfxtp_4
X_52952_ _53221_/A _53062_/A sky130_fd_sc_hd__buf_2
X_64938_ _64915_/X _64926_/Y _64937_/Y _64938_/Y sky130_fd_sc_hd__o21ai_4
X_83772_ _86578_/CLK _70446_/Y _83772_/Q sky130_fd_sc_hd__dfxtp_4
X_80984_ _80813_/CLK _80984_/D _80984_/Q sky130_fd_sc_hd__dfxtp_4
X_85511_ _85507_/CLK _54072_/Y _85511_/Q sky130_fd_sc_hd__dfxtp_4
X_51903_ _85925_/Q _51900_/X _51902_/Y _51903_/Y sky130_fd_sc_hd__o21ai_4
X_82723_ _84119_/CLK _82723_/D _82723_/Q sky130_fd_sc_hd__dfxtp_4
X_55671_ _55671_/A _55671_/Y sky130_fd_sc_hd__inv_2
X_67657_ _64584_/X _67657_/X sky130_fd_sc_hd__buf_2
X_86491_ _86490_/CLK _86491_/D _65521_/B sky130_fd_sc_hd__dfxtp_4
X_52883_ _52867_/A _52879_/B _52872_/C _51192_/D _52883_/X sky130_fd_sc_hd__and4_4
X_64869_ _84224_/Q _64870_/C sky130_fd_sc_hd__inv_2
X_57410_ _57650_/A _56672_/Y _57409_/Y _57410_/Y sky130_fd_sc_hd__a21oi_4
X_88230_ _86965_/CLK _88230_/D _67647_/B sky130_fd_sc_hd__dfxtp_4
X_54622_ _54594_/X _54636_/A sky130_fd_sc_hd__buf_2
X_66608_ _66608_/A _66608_/X sky130_fd_sc_hd__buf_2
X_85442_ _85764_/CLK _85442_/D _85442_/Q sky130_fd_sc_hd__dfxtp_4
X_51834_ _51831_/Y _51823_/X _51833_/X _51834_/Y sky130_fd_sc_hd__a21oi_4
X_58390_ _58408_/A _58403_/B sky130_fd_sc_hd__buf_2
X_82654_ _81755_/CLK _84006_/Q _82654_/Q sky130_fd_sc_hd__dfxtp_4
X_67588_ _67584_/X _67587_/X _67401_/X _67588_/Y sky130_fd_sc_hd__a21oi_4
X_57341_ _56846_/Y _57340_/C _57341_/Y sky130_fd_sc_hd__nand2_4
X_81605_ _81250_/CLK _76198_/Y _81605_/Q sky130_fd_sc_hd__dfxtp_4
X_69327_ _69300_/X _69324_/Y _69325_/X _69326_/Y _69327_/X sky130_fd_sc_hd__a211o_4
X_88161_ _88158_/CLK _88161_/D _88161_/Q sky130_fd_sc_hd__dfxtp_4
X_54553_ _54538_/A _54559_/B _54538_/C _54553_/D _54553_/X sky130_fd_sc_hd__and4_4
X_66539_ _68347_/A _66540_/A sky130_fd_sc_hd__buf_2
X_85373_ _83707_/CLK _85373_/D _85373_/Q sky130_fd_sc_hd__dfxtp_4
X_51765_ _51779_/A _51765_/B _51765_/Y sky130_fd_sc_hd__nand2_4
X_82585_ _82589_/CLK _82617_/Q _78241_/A sky130_fd_sc_hd__dfxtp_4
X_87112_ _87110_/CLK _44433_/X _87112_/Q sky130_fd_sc_hd__dfxtp_4
X_53504_ _53503_/X _53504_/B _53504_/Y sky130_fd_sc_hd__nand2_4
X_84324_ _84321_/CLK _63433_/Y _80568_/B sky130_fd_sc_hd__dfxtp_4
X_50716_ _50738_/A _50716_/B _50716_/Y sky130_fd_sc_hd__nand2_4
X_81536_ _81475_/CLK _81548_/Q _76142_/A sky130_fd_sc_hd__dfxtp_4
X_57272_ _56729_/X _57023_/A _56674_/X _57272_/D _57273_/B sky130_fd_sc_hd__and4_4
X_69258_ _83937_/Q _69230_/X _69257_/X _69258_/X sky130_fd_sc_hd__a21bo_4
X_88092_ _87834_/CLK _88092_/D _74095_/A sky130_fd_sc_hd__dfxtp_4
X_54484_ _54479_/Y _54475_/X _54483_/X _54484_/Y sky130_fd_sc_hd__a21oi_4
X_51696_ _51692_/Y _51693_/X _51695_/X _85963_/D sky130_fd_sc_hd__a21oi_4
X_59011_ _58961_/X _85664_/Q _59010_/X _59011_/X sky130_fd_sc_hd__o21a_4
X_56223_ _56214_/A _56229_/B _56223_/C _56223_/Y sky130_fd_sc_hd__nand3_4
X_68209_ _68208_/X _68209_/X sky130_fd_sc_hd__buf_2
X_87043_ _88097_/CLK _44592_/Y _87043_/Q sky130_fd_sc_hd__dfxtp_4
X_53435_ _85634_/Q _53431_/X _53434_/Y _53435_/Y sky130_fd_sc_hd__o21ai_4
X_84255_ _83491_/CLK _64340_/X _79775_/B sky130_fd_sc_hd__dfxtp_4
X_50647_ _50640_/A _53863_/A _50647_/Y sky130_fd_sc_hd__nand2_4
X_69189_ _83942_/Q _69161_/X _69188_/X _69189_/X sky130_fd_sc_hd__a21bo_4
X_81467_ _82648_/CLK _76879_/B _81467_/Q sky130_fd_sc_hd__dfxtp_4
X_40400_ _40399_/Y _40400_/X sky130_fd_sc_hd__buf_2
X_71220_ _48843_/B _71216_/X _71219_/Y _71220_/Y sky130_fd_sc_hd__o21ai_4
X_83206_ _83846_/CLK _83206_/D _70181_/A sky130_fd_sc_hd__dfxtp_4
X_80418_ _80425_/B _80418_/B _80418_/X sky130_fd_sc_hd__xor2_4
X_56154_ _56140_/A _56150_/B _55707_/B _56154_/Y sky130_fd_sc_hd__nand3_4
X_41380_ _81743_/Q _41379_/X _41380_/X sky130_fd_sc_hd__or2_4
X_53366_ _53311_/A _53371_/A sky130_fd_sc_hd__buf_2
X_84186_ _84192_/CLK _84186_/D _84186_/Q sky130_fd_sc_hd__dfxtp_4
X_50578_ _50578_/A _50578_/B _50578_/X sky130_fd_sc_hd__or2_4
X_81398_ _81346_/CLK _81398_/D _76683_/B sky130_fd_sc_hd__dfxtp_4
X_55105_ _55101_/Y _55102_/X _55104_/X _85318_/D sky130_fd_sc_hd__a21oi_4
X_40331_ _40330_/Y _40331_/X sky130_fd_sc_hd__buf_2
X_52317_ _52299_/A _48992_/X _52317_/Y sky130_fd_sc_hd__nand2_4
X_71151_ _48391_/X _71138_/X _71150_/Y _83590_/D sky130_fd_sc_hd__o21ai_4
X_83137_ _83141_/CLK _73769_/Y _83137_/Q sky130_fd_sc_hd__dfxtp_4
X_56085_ _56084_/Y _56085_/X sky130_fd_sc_hd__buf_2
X_80349_ _80349_/A _80349_/B _80350_/C sky130_fd_sc_hd__nand2_4
X_53297_ _53352_/A _53298_/A sky130_fd_sc_hd__buf_2
X_70102_ _70102_/A _70099_/Y _70100_/Y _70101_/Y _70102_/Y sky130_fd_sc_hd__nand4_4
X_43050_ _43017_/A _43050_/X sky130_fd_sc_hd__buf_2
X_55036_ _55034_/Y _55024_/X _55035_/X _85331_/D sky130_fd_sc_hd__a21oi_4
X_59913_ _59913_/A _59913_/X sky130_fd_sc_hd__buf_2
X_52248_ _48691_/A _52248_/B _52267_/C _52248_/X sky130_fd_sc_hd__and3_4
X_71082_ _71078_/A _71082_/B _71078_/C _71082_/Y sky130_fd_sc_hd__nand3_4
X_83068_ _83068_/CLK _74432_/Y _83068_/Q sky130_fd_sc_hd__dfxtp_4
X_87945_ _87883_/CLK _42274_/X _87945_/Q sky130_fd_sc_hd__dfxtp_4
X_42001_ _41998_/X _41993_/X _40802_/X _41999_/Y _42000_/X _88076_/D
+ sky130_fd_sc_hd__o32ai_4
X_74910_ _74910_/A _74909_/Y _74911_/B sky130_fd_sc_hd__xnor2_4
X_70033_ _70056_/A _70033_/X sky130_fd_sc_hd__buf_2
X_82019_ _82104_/CLK _77744_/B _81987_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_4_6_1_CLK clkbuf_4_6_1_CLK/A clkbuf_4_6_1_CLK/X sky130_fd_sc_hd__clkbuf_1
X_59844_ _59728_/Y _59744_/Y _59840_/Y _59841_/X _59843_/Y _59844_/Y
+ sky130_fd_sc_hd__a41oi_4
X_52179_ _52215_/A _52210_/A sky130_fd_sc_hd__buf_2
X_87876_ _88394_/CLK _42413_/Y _87876_/Q sky130_fd_sc_hd__dfxtp_4
X_75890_ _75889_/Y _75890_/Y sky130_fd_sc_hd__inv_2
X_74841_ _46186_/X _74842_/B _46189_/Y _80671_/D sky130_fd_sc_hd__and3_4
X_86827_ _86824_/CLK _86827_/D _86827_/Q sky130_fd_sc_hd__dfxtp_4
X_59775_ _59775_/A _59660_/C _59660_/D _59775_/X sky130_fd_sc_hd__and3_4
X_56987_ _57416_/A _57416_/C _44213_/X _56987_/Y sky130_fd_sc_hd__a21oi_4
X_46740_ _52645_/B _46740_/X sky130_fd_sc_hd__buf_2
X_58726_ _58699_/A _86388_/Q _58726_/Y sky130_fd_sc_hd__nor2_4
X_77560_ _77559_/X _77560_/Y sky130_fd_sc_hd__inv_2
X_55938_ _55947_/A _85244_/Q _55938_/X sky130_fd_sc_hd__and2_4
X_43952_ _44293_/B _43979_/A _43945_/A _43951_/Y _43952_/X sky130_fd_sc_hd__a211o_4
X_74772_ _74768_/Y _74772_/B _74772_/C _74771_/Y _74777_/B sky130_fd_sc_hd__and4_4
X_86758_ _86758_/CLK _46227_/Y _44146_/A sky130_fd_sc_hd__dfxtp_4
X_71984_ _71982_/Y _71978_/X _71983_/X _83308_/D sky130_fd_sc_hd__a21oi_4
X_76511_ _76509_/X _76511_/B _76511_/X sky130_fd_sc_hd__and2_4
X_42903_ _42895_/X _42896_/X _41667_/X _87660_/Q _42881_/X _42903_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73723_ _88108_/Q _73649_/X _73723_/Y sky130_fd_sc_hd__nor2_4
X_85709_ _85709_/CLK _85709_/D _85709_/Q sky130_fd_sc_hd__dfxtp_4
X_46671_ _46664_/Y _46654_/X _46670_/X _46671_/Y sky130_fd_sc_hd__a21oi_4
X_58657_ _58112_/X _86106_/Q _58656_/X _58657_/Y sky130_fd_sc_hd__o21ai_4
X_70935_ _70935_/A _70959_/B _71115_/D _71115_/B _70935_/X sky130_fd_sc_hd__and4_4
X_77491_ _77487_/Y _77489_/Y _77486_/Y _77491_/Y sky130_fd_sc_hd__o21ai_4
X_43883_ _41294_/X _43879_/X _87218_/Q _43880_/X _87218_/D sky130_fd_sc_hd__a2bb2o_4
X_55869_ _55866_/X _55868_/X _55517_/X _55872_/A sky130_fd_sc_hd__a21o_4
X_86689_ _86688_/CLK _46927_/Y _58997_/A sky130_fd_sc_hd__dfxtp_4
X_48410_ _83588_/Q _74389_/B sky130_fd_sc_hd__inv_2
X_79230_ _79230_/A _79229_/Y _79230_/Y sky130_fd_sc_hd__nand2_4
X_45622_ _45621_/Y _44975_/A _45622_/X sky130_fd_sc_hd__and2_4
X_57608_ _71993_/A _57608_/X sky130_fd_sc_hd__buf_2
X_76442_ _76419_/Y _76433_/X _76443_/A sky130_fd_sc_hd__nor2_4
X_42834_ _41485_/X _42830_/X _66689_/B _42832_/X _42834_/X sky130_fd_sc_hd__a2bb2o_4
X_49390_ _49410_/A _46662_/X _49390_/Y sky130_fd_sc_hd__nand2_4
X_73654_ _68468_/B _73597_/X _73652_/X _73653_/Y _73654_/X sky130_fd_sc_hd__a211o_4
X_70866_ _70866_/A _70869_/C sky130_fd_sc_hd__buf_2
X_58588_ _86719_/Q _58614_/B _58588_/Y sky130_fd_sc_hd__nor2_4
X_48341_ _66326_/B _48333_/X _48340_/Y _48341_/Y sky130_fd_sc_hd__o21ai_4
X_72605_ _60053_/X _72537_/Y _72569_/C _72569_/A _72604_/Y _72605_/Y
+ sky130_fd_sc_hd__a41oi_4
X_79161_ _79158_/Y _79160_/Y _79161_/Y sky130_fd_sc_hd__nand2_4
X_57539_ _48234_/A _46620_/A _53697_/B _57539_/Y sky130_fd_sc_hd__nand3_4
X_45553_ _45553_/A _45617_/B _45553_/Y sky130_fd_sc_hd__nor2_4
X_76373_ _76355_/Y _76361_/Y _76353_/Y _76373_/X sky130_fd_sc_hd__o21a_4
X_88359_ _86998_/CLK _40658_/Y _88359_/Q sky130_fd_sc_hd__dfxtp_4
X_42765_ _41294_/X _42757_/X _67368_/B _42759_/X _42765_/X sky130_fd_sc_hd__a2bb2o_4
X_73585_ _73497_/A _65921_/B _73585_/X sky130_fd_sc_hd__and2_4
X_70797_ _52876_/B _70761_/A _70796_/Y _70797_/Y sky130_fd_sc_hd__o21ai_4
X_78112_ _78112_/A _78112_/B _78112_/X sky130_fd_sc_hd__xor2_4
X_44504_ _41259_/A _44502_/X _87077_/Q _44503_/X _87077_/D sky130_fd_sc_hd__a2bb2o_4
X_75324_ _75323_/X _75324_/Y sky130_fd_sc_hd__inv_2
X_41716_ _41715_/X _41682_/X _67724_/B _41684_/X _41716_/X sky130_fd_sc_hd__a2bb2o_4
X_48272_ _66159_/B _48241_/X _48271_/Y _48272_/Y sky130_fd_sc_hd__o21ai_4
X_60550_ _60473_/C _60602_/B sky130_fd_sc_hd__buf_2
X_72536_ _72506_/C _72516_/C _72537_/B sky130_fd_sc_hd__nor2_4
X_79092_ _82655_/Q _82527_/D _79091_/X _79092_/Y sky130_fd_sc_hd__o21ai_4
X_45484_ _45478_/X _45481_/X _45483_/Y _45484_/Y sky130_fd_sc_hd__a21oi_4
X_42696_ _42681_/A _42696_/X sky130_fd_sc_hd__buf_2
X_47223_ _57698_/A _47192_/X _47222_/Y _47223_/Y sky130_fd_sc_hd__o21ai_4
X_59209_ _59105_/X _85744_/Q _59106_/X _59209_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_10_464_0_CLK clkbuf_9_232_0_CLK/X _86372_/CLK sky130_fd_sc_hd__clkbuf_1
X_78043_ _78043_/A _78043_/Y sky130_fd_sc_hd__inv_2
X_44435_ _41592_/X _44431_/X _87110_/Q _44432_/X _87110_/D sky130_fd_sc_hd__a2bb2o_4
X_75255_ _75255_/A _80943_/D _75258_/B sky130_fd_sc_hd__nor2_4
X_41647_ _41646_/Y _41647_/X sky130_fd_sc_hd__buf_2
X_60481_ _60481_/A _60481_/X sky130_fd_sc_hd__buf_2
X_72467_ _57709_/X _85347_/Q _72466_/X _72467_/Y sky130_fd_sc_hd__o21ai_4
X_62220_ _62194_/A _58221_/X _62219_/X _62244_/D _62220_/X sky130_fd_sc_hd__and4_4
X_74206_ _74206_/A _73577_/B _74206_/Y sky130_fd_sc_hd__nor2_4
X_47154_ _54576_/D _51192_/D sky130_fd_sc_hd__buf_2
X_71418_ _71221_/A _71418_/B _71419_/A sky130_fd_sc_hd__and2_4
X_44366_ _41741_/X _44364_/X _87146_/Q _44365_/X _44366_/X sky130_fd_sc_hd__a2bb2o_4
X_75186_ _75186_/A _75186_/B _75190_/C sky130_fd_sc_hd__nand2_4
X_41578_ _41358_/X _82314_/Q _41578_/X sky130_fd_sc_hd__or2_4
X_72398_ _72327_/X _85962_/Q _72397_/X _72398_/Y sky130_fd_sc_hd__o21ai_4
X_46105_ _46104_/Y _46214_/C sky130_fd_sc_hd__buf_2
X_43317_ _43316_/X _43305_/X _41234_/X _87484_/Q _43308_/X _43318_/A
+ sky130_fd_sc_hd__o32ai_4
X_62151_ _58983_/A _62151_/X sky130_fd_sc_hd__buf_2
X_74137_ _74117_/A _74136_/Y _74137_/Y sky130_fd_sc_hd__nor2_4
X_40529_ _40528_/X _40508_/X _88376_/Q _40510_/X _88376_/D sky130_fd_sc_hd__a2bb2o_4
X_47085_ _47067_/A _47082_/X _47048_/C _52846_/D _47085_/X sky130_fd_sc_hd__and4_4
X_71349_ _71504_/C _71160_/C _71422_/C _71349_/D _71349_/X sky130_fd_sc_hd__and4_4
X_44297_ _68714_/A _69442_/A sky130_fd_sc_hd__buf_2
X_79994_ _84928_/Q _65817_/C _79994_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_479_0_CLK clkbuf_9_239_0_CLK/X _85773_/CLK sky130_fd_sc_hd__clkbuf_1
X_61102_ _64323_/A _61102_/X sky130_fd_sc_hd__buf_2
X_46036_ _41484_/Y _46029_/X _66691_/B _46030_/X _46036_/X sky130_fd_sc_hd__a2bb2o_4
X_43248_ _43218_/A _43248_/X sky130_fd_sc_hd__buf_2
X_62082_ _59858_/A _61609_/X _62081_/X _62082_/X sky130_fd_sc_hd__a21o_4
X_74068_ _74066_/X _74055_/X _74057_/Y _74068_/Y sky130_fd_sc_hd__nand3_4
X_78945_ _78928_/A _82512_/D _78944_/Y _78945_/Y sky130_fd_sc_hd__a21oi_4
X_65910_ _65907_/X _65909_/X _65809_/X _65910_/X sky130_fd_sc_hd__a21o_4
X_73019_ _53663_/B _73019_/B _73019_/X sky130_fd_sc_hd__xor2_4
X_61033_ _60969_/X _61000_/X _84534_/Q _61033_/X sky130_fd_sc_hd__or3_4
X_43179_ _43178_/X _43180_/A sky130_fd_sc_hd__buf_2
X_66890_ _87366_/Q _66797_/X _66863_/X _66889_/X _66890_/X sky130_fd_sc_hd__a211o_4
X_78876_ _78877_/B _78877_/A _78876_/X sky130_fd_sc_hd__or2_4
Xclkbuf_10_402_0_CLK clkbuf_9_201_0_CLK/X _85342_/CLK sky130_fd_sc_hd__clkbuf_1
X_65841_ _65838_/X _66423_/B _65840_/X _65841_/Y sky130_fd_sc_hd__nand3_4
X_77827_ _77827_/A _77826_/Y _77835_/B sky130_fd_sc_hd__xor2_4
X_47987_ _53531_/B _50306_/B sky130_fd_sc_hd__buf_2
X_49726_ _49716_/X _52940_/B _49726_/Y sky130_fd_sc_hd__nand2_4
X_68560_ _68560_/A _88364_/Q _68560_/X sky130_fd_sc_hd__and2_4
X_46938_ _46948_/A _52760_/B _46938_/Y sky130_fd_sc_hd__nand2_4
X_65772_ _65772_/A _65772_/B _65772_/Y sky130_fd_sc_hd__nand2_4
X_77758_ _77758_/A _77758_/Y sky130_fd_sc_hd__inv_2
X_62984_ _62980_/Y _62642_/B _62981_/Y _62982_/Y _62983_/X _62984_/X
+ sky130_fd_sc_hd__a41o_4
X_67511_ _68392_/A _67987_/A sky130_fd_sc_hd__buf_2
X_64723_ _44175_/A _65718_/A sky130_fd_sc_hd__buf_2
X_76709_ _76696_/X _76709_/B _76709_/X sky130_fd_sc_hd__and2_4
X_49657_ _49657_/A _49669_/C sky130_fd_sc_hd__buf_2
X_61935_ _61490_/X _61933_/X _61907_/C _61952_/D _61935_/Y sky130_fd_sc_hd__nand4_4
X_68491_ _44149_/A _68491_/B _68491_/Y sky130_fd_sc_hd__nor2_4
X_46869_ _46864_/Y _46844_/X _46868_/X _86695_/D sky130_fd_sc_hd__a21oi_4
X_77689_ _77687_/Y _77688_/Y _77690_/B _77689_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_417_0_CLK clkbuf_9_208_0_CLK/X _82820_/CLK sky130_fd_sc_hd__clkbuf_1
X_48608_ _48606_/X _81771_/Q _48607_/Y _48609_/A sky130_fd_sc_hd__o21ai_4
X_67442_ _67203_/X _67442_/X sky130_fd_sc_hd__buf_2
X_79428_ _79433_/A _79433_/B _79428_/Y sky130_fd_sc_hd__xnor2_4
X_64654_ _64589_/X _85567_/Q _64591_/X _64653_/X _64654_/X sky130_fd_sc_hd__a211o_4
X_61866_ _61864_/Y _61801_/X _61865_/Y _61866_/Y sky130_fd_sc_hd__a21oi_4
X_49588_ _49571_/X _49592_/B _49577_/C _52801_/D _49588_/X sky130_fd_sc_hd__and4_4
X_63605_ _63603_/Y _63578_/X _63604_/Y _84310_/D sky130_fd_sc_hd__a21oi_4
X_60817_ _60826_/A _60810_/B _60817_/C _60817_/Y sky130_fd_sc_hd__nor3_4
X_48539_ _48538_/Y _48540_/B sky130_fd_sc_hd__buf_2
X_79359_ _79354_/X _79358_/Y _82834_/D sky130_fd_sc_hd__xor2_4
X_67373_ _67324_/A _67373_/B _67373_/X sky130_fd_sc_hd__and2_4
X_64585_ _64584_/X _64777_/A sky130_fd_sc_hd__buf_2
X_61797_ _61966_/A _61846_/C sky130_fd_sc_hd__buf_2
X_69112_ _88084_/Q _68883_/X _68884_/X _69111_/Y _69112_/X sky130_fd_sc_hd__a211o_4
X_66324_ _58697_/A _85604_/Q _66251_/X _66323_/X _66324_/X sky130_fd_sc_hd__a211o_4
X_51550_ _51545_/A _53076_/B _51550_/Y sky130_fd_sc_hd__nand2_4
X_63536_ _63413_/A _63537_/C sky130_fd_sc_hd__buf_2
X_82370_ _84951_/CLK _82178_/Q _82370_/Q sky130_fd_sc_hd__dfxtp_4
X_60748_ _60667_/A _60748_/X sky130_fd_sc_hd__buf_2
X_50501_ _50575_/A _48820_/B _50501_/Y sky130_fd_sc_hd__nand2_4
X_81321_ _81351_/CLK _81321_/D _81729_/D sky130_fd_sc_hd__dfxtp_4
X_69043_ _87991_/Q _68975_/X _68976_/X _69042_/X _69043_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_8_91_0_CLK clkbuf_8_91_0_CLK/A clkbuf_8_91_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_66255_ _64898_/A _66326_/A sky130_fd_sc_hd__buf_2
X_51481_ _51481_/A _53005_/B _51481_/Y sky130_fd_sc_hd__nand2_4
X_63467_ _63528_/A _63517_/A sky130_fd_sc_hd__buf_2
X_60679_ _60724_/B _63630_/B sky130_fd_sc_hd__buf_2
X_65206_ _65206_/A _86442_/Q _65206_/X sky130_fd_sc_hd__and2_4
X_53220_ _85674_/Q _53198_/X _53219_/Y _53220_/Y sky130_fd_sc_hd__o21ai_4
X_84040_ _81169_/CLK _68095_/X _84040_/Q sky130_fd_sc_hd__dfxtp_4
X_50432_ _50432_/A _52137_/B _50432_/Y sky130_fd_sc_hd__nand2_4
X_62418_ _61502_/A _62472_/B _62386_/C _62431_/D _62421_/B sky130_fd_sc_hd__nand4_4
X_81252_ _81282_/CLK _81284_/Q _76171_/A sky130_fd_sc_hd__dfxtp_4
X_66186_ _65407_/A _66186_/X sky130_fd_sc_hd__buf_2
X_63398_ _63398_/A _63427_/A sky130_fd_sc_hd__buf_2
X_80203_ _84948_/Q _84196_/Q _80203_/Y sky130_fd_sc_hd__nand2_4
X_53151_ _53139_/A _53159_/B _53143_/X _53151_/D _53151_/X sky130_fd_sc_hd__and4_4
X_65137_ _65164_/A _86445_/Q _65137_/X sky130_fd_sc_hd__and2_4
X_50363_ _50594_/A _50363_/X sky130_fd_sc_hd__buf_2
X_62349_ _62632_/A _58506_/A _62632_/C _62351_/C sky130_fd_sc_hd__nand3_4
X_81183_ _86758_/CLK _75059_/X _81183_/Q sky130_fd_sc_hd__dfxtp_4
X_52102_ _51265_/A _52135_/B sky130_fd_sc_hd__buf_2
X_80134_ _80132_/X _80141_/B _80134_/Y sky130_fd_sc_hd__xnor2_4
X_53082_ _53111_/A _53082_/X sky130_fd_sc_hd__buf_2
X_69945_ _43199_/A _69833_/X _68348_/X _69944_/X _69945_/X sky130_fd_sc_hd__a211o_4
X_65068_ _65063_/X _65192_/B _65067_/X _65068_/Y sky130_fd_sc_hd__nand3_4
X_50294_ _86229_/Q _50282_/X _50293_/Y _50294_/Y sky130_fd_sc_hd__o21ai_4
X_85991_ _85700_/CLK _85991_/D _85991_/Q sky130_fd_sc_hd__dfxtp_4
X_52033_ _51956_/X _52033_/X sky130_fd_sc_hd__buf_2
X_56910_ _55218_/Y _56908_/X _56909_/Y _56910_/X sky130_fd_sc_hd__a21o_4
X_87730_ _82906_/CLK _42765_/X _67368_/B sky130_fd_sc_hd__dfxtp_4
X_64019_ _61541_/B _64052_/B _64003_/C _64052_/D _64019_/Y sky130_fd_sc_hd__nand4_4
X_84942_ _85489_/CLK _57895_/Y _84942_/Q sky130_fd_sc_hd__dfxtp_4
X_80065_ _80073_/A _80064_/Y _80065_/Y sky130_fd_sc_hd__xnor2_4
X_57890_ _57886_/Y _57888_/Y _57889_/X _57890_/X sky130_fd_sc_hd__a21o_4
X_69876_ _69872_/X _69875_/X _69678_/X _69876_/X sky130_fd_sc_hd__a21o_4
X_56841_ _56841_/A _85129_/D sky130_fd_sc_hd__inv_2
X_68827_ _73987_/A _68778_/X _68800_/X _68826_/Y _68827_/X sky130_fd_sc_hd__a211o_4
X_87661_ _87471_/CLK _42902_/X _87661_/Q sky130_fd_sc_hd__dfxtp_4
X_84873_ _84299_/CLK _84873_/D _84873_/Q sky130_fd_sc_hd__dfxtp_4
X_86612_ _85969_/CLK _86612_/D _86612_/Q sky130_fd_sc_hd__dfxtp_4
X_83824_ _83187_/CLK _83824_/D _74797_/A sky130_fd_sc_hd__dfxtp_4
X_59560_ _59560_/A _59890_/C sky130_fd_sc_hd__buf_2
X_56772_ _56684_/B _56772_/Y sky130_fd_sc_hd__inv_2
X_68758_ _69357_/A _68759_/A sky130_fd_sc_hd__buf_2
X_87592_ _87045_/CLK _87592_/D _43057_/A sky130_fd_sc_hd__dfxtp_4
X_53984_ _53981_/Y _53982_/X _53983_/Y _53984_/Y sky130_fd_sc_hd__a21boi_4
X_58511_ _58511_/A _58510_/X _58511_/Y sky130_fd_sc_hd__nor2_4
X_55723_ _56267_/C _55126_/A _55133_/X _55722_/X _55723_/X sky130_fd_sc_hd__a211o_4
X_67709_ _67014_/X _67709_/X sky130_fd_sc_hd__buf_2
X_86543_ _86576_/CLK _86543_/D _66171_/B sky130_fd_sc_hd__dfxtp_4
X_52935_ _52932_/Y _52920_/X _52934_/X _85728_/D sky130_fd_sc_hd__a21oi_4
X_59491_ _46159_/X _59488_/Y _59490_/Y _59491_/Y sky130_fd_sc_hd__a21oi_4
X_83755_ _83421_/CLK _83755_/D _83755_/Q sky130_fd_sc_hd__dfxtp_4
X_80967_ _83957_/CLK _80967_/D _80955_/D sky130_fd_sc_hd__dfxtp_4
X_68689_ _68666_/X _68612_/X _68678_/Y _68688_/Y _68689_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_8_44_0_CLK clkbuf_8_45_0_CLK/A clkbuf_9_88_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_70720_ _52773_/B _70699_/X _70719_/Y _70720_/Y sky130_fd_sc_hd__o21ai_4
X_58442_ _58442_/A _58426_/X _58442_/Y sky130_fd_sc_hd__nand2_4
X_82706_ _82665_/CLK _78958_/X _78358_/B sky130_fd_sc_hd__dfxtp_4
X_55654_ _55654_/A _55654_/X sky130_fd_sc_hd__buf_2
X_86474_ _86506_/CLK _86474_/D _86474_/Q sky130_fd_sc_hd__dfxtp_4
X_40880_ _40877_/X _82860_/Q _40879_/X _40881_/A sky130_fd_sc_hd__o21ai_4
X_52866_ _52757_/A _52867_/A sky130_fd_sc_hd__buf_2
X_83686_ _83685_/CLK _70842_/Y _83686_/Q sky130_fd_sc_hd__dfxtp_4
X_80898_ _82067_/CLK _84074_/Q _75568_/A sky130_fd_sc_hd__dfxtp_4
X_88213_ _88215_/CLK _88213_/D _68047_/B sky130_fd_sc_hd__dfxtp_4
X_54605_ _54600_/A _53426_/B _54605_/Y sky130_fd_sc_hd__nand2_4
X_85425_ _85651_/CLK _54532_/Y _85425_/Q sky130_fd_sc_hd__dfxtp_4
X_51817_ _51789_/A _51817_/X sky130_fd_sc_hd__buf_2
X_70651_ _70635_/A _70656_/B sky130_fd_sc_hd__buf_2
X_82637_ _81746_/CLK _83989_/Q _82637_/Q sky130_fd_sc_hd__dfxtp_4
X_58373_ _84866_/Q _58374_/A sky130_fd_sc_hd__buf_2
X_55585_ _44064_/X _55585_/B _55585_/Y sky130_fd_sc_hd__nor2_4
X_52797_ _52784_/X _52818_/B _52789_/X _52797_/D _52797_/X sky130_fd_sc_hd__and4_4
XPHY_20 sky130_fd_sc_hd__decap_3
X_57324_ _56787_/X _56785_/B _57318_/D _56788_/A _56810_/X _57324_/X
+ sky130_fd_sc_hd__a41o_4
XPHY_31 sky130_fd_sc_hd__decap_3
X_88144_ _88144_/CLK _88144_/D _88144_/Q sky130_fd_sc_hd__dfxtp_4
X_42550_ _42550_/A _42550_/Y sky130_fd_sc_hd__inv_2
X_54536_ _54400_/A _54537_/A sky130_fd_sc_hd__buf_2
X_73370_ _73370_/A _73370_/B _73370_/Y sky130_fd_sc_hd__nor2_4
X_85356_ _86282_/CLK _54906_/Y _85356_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_42 sky130_fd_sc_hd__decap_3
X_51748_ _51842_/A _51814_/A sky130_fd_sc_hd__buf_2
X_70582_ _70576_/X _74515_/C _71735_/A _70582_/X sky130_fd_sc_hd__and3_4
X_82568_ _82924_/CLK _82568_/D _82568_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_53 sky130_fd_sc_hd__decap_3
XPHY_64 sky130_fd_sc_hd__decap_3
Xclkbuf_8_59_0_CLK clkbuf_8_59_0_CLK/A clkbuf_8_59_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_41501_ _81177_/Q _41523_/B _41501_/X sky130_fd_sc_hd__or2_4
X_72321_ _72270_/X _72319_/Y _72320_/Y _72296_/X _72274_/X _72321_/X
+ sky130_fd_sc_hd__o32a_4
XPHY_75 sky130_fd_sc_hd__decap_3
X_84307_ _84308_/CLK _63637_/Y _63636_/C sky130_fd_sc_hd__dfxtp_4
X_57255_ _56613_/X _57247_/Y _57254_/Y _57255_/Y sky130_fd_sc_hd__a21oi_4
X_81519_ _82642_/CLK _81563_/Q _81519_/Q sky130_fd_sc_hd__dfxtp_4
X_88075_ _83158_/CLK _42003_/Y _42002_/A sky130_fd_sc_hd__dfxtp_4
XPHY_86 sky130_fd_sc_hd__decap_3
X_42481_ _42466_/X _42467_/X _40641_/X _68588_/A _42480_/X _42482_/A
+ sky130_fd_sc_hd__o32ai_4
X_54467_ _54453_/X _54471_/B _54471_/C _46964_/A _54467_/X sky130_fd_sc_hd__and4_4
X_85287_ _83013_/CLK _56151_/Y _55761_/B sky130_fd_sc_hd__dfxtp_4
X_51679_ _51657_/X _51684_/B _51684_/C _53203_/D _51679_/X sky130_fd_sc_hd__and4_4
XPHY_97 sky130_fd_sc_hd__decap_3
X_82499_ _82924_/CLK _82499_/D _82499_/Q sky130_fd_sc_hd__dfxtp_4
X_44220_ _44220_/A _44220_/B _44220_/Y sky130_fd_sc_hd__nor2_4
X_56206_ _56200_/X _56205_/X _56206_/C _56206_/Y sky130_fd_sc_hd__nand3_4
X_75040_ _81149_/D _75040_/B _75051_/B sky130_fd_sc_hd__nand2_4
X_87026_ _87026_/CLK _44631_/Y _87026_/Q sky130_fd_sc_hd__dfxtp_4
X_41432_ _41412_/X _82886_/Q _41431_/X _41432_/Y sky130_fd_sc_hd__o21ai_4
X_53418_ _53282_/A _53418_/X sky130_fd_sc_hd__buf_2
X_72252_ _57696_/X _72348_/B sky130_fd_sc_hd__buf_2
X_84238_ _84458_/CLK _64519_/X _79581_/B sky130_fd_sc_hd__dfxtp_4
X_57186_ _56691_/A _57186_/B _57187_/A sky130_fd_sc_hd__or2_4
X_54398_ _85449_/Q _54376_/X _54397_/Y _54398_/Y sky130_fd_sc_hd__o21ai_4
X_71203_ _48811_/B _71190_/X _71202_/Y _83574_/D sky130_fd_sc_hd__o21ai_4
X_44151_ _44150_/X _44151_/X sky130_fd_sc_hd__buf_2
X_56137_ _56112_/X _56134_/X _56136_/Y _85290_/D sky130_fd_sc_hd__o21ai_4
X_53349_ _53346_/Y _53328_/X _53348_/X _85650_/D sky130_fd_sc_hd__a21oi_4
X_41363_ _41253_/A _41363_/X sky130_fd_sc_hd__buf_2
X_72183_ _72155_/X _85692_/Q _72156_/X _72183_/X sky130_fd_sc_hd__o21a_4
X_84169_ _82748_/CLK _84169_/D _65916_/C sky130_fd_sc_hd__dfxtp_4
X_43102_ _43101_/Y _87575_/D sky130_fd_sc_hd__inv_2
X_71134_ _50721_/B _71117_/A _71133_/Y _71134_/Y sky130_fd_sc_hd__o21ai_4
X_44082_ _44081_/X _55620_/A sky130_fd_sc_hd__buf_2
X_56068_ _55995_/X _55863_/X _56073_/A _56068_/X sky130_fd_sc_hd__and3_4
X_41294_ _41294_/A _41294_/X sky130_fd_sc_hd__buf_2
X_76991_ _84543_/Q _84415_/Q _76991_/X sky130_fd_sc_hd__xor2_4
X_47910_ _47910_/A _57523_/B sky130_fd_sc_hd__inv_2
X_43033_ _43024_/A _43058_/A sky130_fd_sc_hd__buf_2
X_55019_ _55016_/Y _54998_/X _55018_/X _55019_/Y sky130_fd_sc_hd__a21oi_4
X_78730_ _78729_/A _82686_/D _78731_/A sky130_fd_sc_hd__nand2_4
X_71065_ _48944_/B _71046_/X _71064_/Y _71065_/Y sky130_fd_sc_hd__o21ai_4
X_75942_ _75936_/Y _75941_/Y _75933_/B _75942_/Y sky130_fd_sc_hd__a21oi_4
X_87928_ _88376_/CLK _87928_/D _87928_/Q sky130_fd_sc_hd__dfxtp_4
X_48890_ _86464_/Q _48669_/X _48889_/Y _48890_/Y sky130_fd_sc_hd__o21ai_4
X_70016_ _69689_/X _69692_/X _70001_/X _70016_/Y sky130_fd_sc_hd__a21oi_4
X_47841_ _47841_/A _47855_/A sky130_fd_sc_hd__buf_2
X_59827_ _80413_/A _59822_/X _59826_/Y _59812_/Y _84693_/D sky130_fd_sc_hd__o22a_4
X_78661_ _78661_/A _82694_/Q _78661_/Y sky130_fd_sc_hd__nand2_4
X_75873_ _75875_/C _75873_/Y sky130_fd_sc_hd__inv_2
X_87859_ _87859_/CLK _87859_/D _68361_/A sky130_fd_sc_hd__dfxtp_4
X_77612_ _77612_/A _82108_/D _77612_/Y sky130_fd_sc_hd__nand2_4
X_74824_ _74824_/A _80661_/D sky130_fd_sc_hd__inv_2
X_47772_ _47771_/Y _53236_/B sky130_fd_sc_hd__buf_2
X_59758_ _59687_/Y _59758_/X sky130_fd_sc_hd__buf_2
X_78592_ _78600_/A _78581_/B _78575_/B _78593_/B sky130_fd_sc_hd__o21ai_4
X_44984_ _56390_/C _44945_/X _44983_/X _44984_/Y sky130_fd_sc_hd__o21ai_4
X_49511_ _49509_/Y _49487_/X _49510_/X _86374_/D sky130_fd_sc_hd__a21oi_4
X_46723_ _46733_/A _51807_/B _46723_/Y sky130_fd_sc_hd__nand2_4
X_58709_ _58705_/Y _58708_/Y _58610_/X _58709_/X sky130_fd_sc_hd__a21o_4
X_77543_ _77561_/C _77561_/D _77547_/A sky130_fd_sc_hd__nand2_4
X_43935_ _41437_/X _43928_/X _68000_/B _43929_/X _87191_/D sky130_fd_sc_hd__a2bb2o_4
X_74755_ _70586_/X _74755_/B _74753_/X _74755_/X sky130_fd_sc_hd__and3_4
X_71967_ _71972_/A _48899_/Y _71967_/Y sky130_fd_sc_hd__nand2_4
X_59689_ _59689_/A _59689_/B _59689_/Y sky130_fd_sc_hd__nand2_4
X_61720_ _61703_/X _61715_/Y _61717_/X _58147_/A _61719_/X _61720_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49442_ _49439_/Y _49434_/X _49441_/X _49442_/Y sky130_fd_sc_hd__a21oi_4
X_73706_ _44684_/Y _73420_/X _73705_/Y _73719_/C sky130_fd_sc_hd__a21o_4
X_70918_ _70913_/A _70919_/D sky130_fd_sc_hd__buf_2
X_46654_ _46751_/A _46654_/X sky130_fd_sc_hd__buf_2
X_77474_ _77475_/A _77475_/B _77473_/Y _77478_/B sky130_fd_sc_hd__o21a_4
X_43866_ _43862_/X _43854_/X _41245_/X _87227_/Q _43863_/X _43867_/A
+ sky130_fd_sc_hd__o32ai_4
X_74686_ _82985_/Q _74656_/X _74685_/Y _74687_/A sky130_fd_sc_hd__o21ai_4
X_71898_ _70374_/X _71893_/X _71755_/X _71898_/D _71898_/Y sky130_fd_sc_hd__nand4_4
X_79213_ _79213_/A _79212_/Y _79213_/Y sky130_fd_sc_hd__nand2_4
X_45605_ _85140_/Q _45464_/X _44964_/X _45605_/Y sky130_fd_sc_hd__o21ai_4
X_76425_ _76408_/Y _76409_/Y _76410_/Y _76425_/X sky130_fd_sc_hd__o21a_4
X_42817_ _42723_/A _42817_/X sky130_fd_sc_hd__buf_2
X_49373_ _58587_/B _49360_/X _49372_/Y _49373_/Y sky130_fd_sc_hd__o21ai_4
X_61651_ _61400_/X _61675_/C sky130_fd_sc_hd__buf_2
X_73637_ _73605_/X _86238_/Q _44194_/X _73636_/X _73637_/X sky130_fd_sc_hd__a211o_4
X_46585_ _83779_/Q _46585_/Y sky130_fd_sc_hd__inv_2
X_70849_ _70903_/A _70890_/B _70849_/C _70860_/D _70849_/Y sky130_fd_sc_hd__nand4_4
X_43797_ _43760_/A _43797_/X sky130_fd_sc_hd__buf_2
X_48324_ _48112_/B _50368_/B sky130_fd_sc_hd__buf_2
X_60602_ _60488_/B _60602_/B _60421_/B _60603_/C sky130_fd_sc_hd__nand3_4
X_79144_ _79144_/A _84476_/Q _79144_/X sky130_fd_sc_hd__xor2_4
X_45536_ _45533_/Y _45516_/X _45471_/X _45535_/Y _45536_/X sky130_fd_sc_hd__a211o_4
X_64370_ _64363_/X _64364_/X _64366_/X _64369_/Y _64326_/X _64370_/X
+ sky130_fd_sc_hd__o41a_4
X_76356_ _76356_/A _76325_/A _76356_/Y sky130_fd_sc_hd__nor2_4
X_42748_ _42739_/X _42740_/X _41234_/X _68941_/B _42732_/X _42749_/A
+ sky130_fd_sc_hd__o32ai_4
X_61582_ _61582_/A _72550_/A _72506_/C _61367_/D _61582_/Y sky130_fd_sc_hd__nand4_4
X_73568_ _73588_/A _73568_/B _73568_/X sky130_fd_sc_hd__and2_4
X_63321_ _59436_/Y _63259_/X _63234_/X _58985_/A _63235_/X _63321_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75307_ _75305_/X _75276_/Y _75306_/Y _75307_/X sky130_fd_sc_hd__a21o_4
X_48255_ _66119_/B _48241_/X _48254_/Y _48255_/Y sky130_fd_sc_hd__o21ai_4
X_60533_ _60442_/C _60533_/Y sky130_fd_sc_hd__inv_2
X_72519_ _72555_/B _72597_/C sky130_fd_sc_hd__buf_2
X_79075_ _79087_/B _79075_/Y sky130_fd_sc_hd__inv_2
X_45467_ _63051_/B _61378_/A sky130_fd_sc_hd__buf_2
X_76287_ _81355_/Q _81611_/D _76287_/X sky130_fd_sc_hd__xor2_4
X_42679_ _42651_/X _42679_/X sky130_fd_sc_hd__buf_2
X_73499_ _73496_/X _73498_/X _73383_/X _73502_/A sky130_fd_sc_hd__a21o_4
X_47206_ _47196_/A _51222_/B _47206_/Y sky130_fd_sc_hd__nand2_4
X_66040_ _65595_/X _66040_/X sky130_fd_sc_hd__buf_2
X_78026_ _78025_/X _78027_/B sky130_fd_sc_hd__inv_2
X_44418_ _44418_/A _87119_/D sky130_fd_sc_hd__inv_2
X_63252_ _61580_/X _63252_/B _60602_/B _60570_/C _63252_/Y sky130_fd_sc_hd__nand4_4
X_75238_ _81070_/Q _75240_/A sky130_fd_sc_hd__inv_2
X_48186_ _48186_/A _48535_/A sky130_fd_sc_hd__buf_2
X_60464_ _60515_/C _60476_/C sky130_fd_sc_hd__buf_2
X_45398_ _85057_/Q _45397_/X _45398_/Y sky130_fd_sc_hd__nor2_4
X_62203_ _62203_/A _62203_/Y sky130_fd_sc_hd__inv_2
X_47137_ _47109_/A _52876_/B _47137_/Y sky130_fd_sc_hd__nand2_4
X_44349_ _44348_/Y _87153_/D sky130_fd_sc_hd__inv_2
X_75169_ _80681_/Q _80937_/D _75169_/Y sky130_fd_sc_hd__nor2_4
X_63183_ _63018_/X _63183_/X sky130_fd_sc_hd__buf_2
X_60395_ _60501_/A _60440_/A _60395_/X sky130_fd_sc_hd__and2_4
X_62134_ _62132_/Y _62101_/X _62133_/Y _84431_/D sky130_fd_sc_hd__a21oi_4
X_47068_ _47064_/Y _47035_/X _47067_/X _47068_/Y sky130_fd_sc_hd__a21oi_4
X_67991_ _68370_/A _67991_/X sky130_fd_sc_hd__buf_2
X_79977_ _79977_/A _79973_/Y _79976_/Y _79980_/A sky130_fd_sc_hd__nand3_4
X_46019_ _40527_/Y _46007_/X _67215_/B _46008_/X _46019_/X sky130_fd_sc_hd__a2bb2o_4
X_69730_ _69579_/X _69727_/Y _69672_/X _69729_/Y _69730_/X sky130_fd_sc_hd__a211o_4
X_66942_ _66942_/A _88132_/Q _66942_/X sky130_fd_sc_hd__and2_4
X_62065_ _84836_/Q _62065_/B _62063_/X _62065_/D _62066_/D sky130_fd_sc_hd__nand4_4
Xclkbuf_10_341_0_CLK clkbuf_9_170_0_CLK/X _85738_/CLK sky130_fd_sc_hd__clkbuf_1
X_78928_ _78928_/A _78928_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_971_0_CLK clkbuf_9_485_0_CLK/X _83589_/CLK sky130_fd_sc_hd__clkbuf_1
X_61016_ _60944_/Y _64102_/B _61016_/Y sky130_fd_sc_hd__nand2_4
X_69661_ _69661_/A _69661_/B _69661_/Y sky130_fd_sc_hd__nor2_4
X_66873_ _66757_/X _66859_/Y _66793_/X _66872_/Y _66873_/X sky130_fd_sc_hd__a211o_4
X_78859_ _78858_/Y _78859_/Y sky130_fd_sc_hd__inv_2
X_68612_ _60111_/X _68612_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_462_0_CLK clkbuf_8_231_0_CLK/X clkbuf_9_462_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_65824_ _65595_/X _65824_/X sky130_fd_sc_hd__buf_2
X_69592_ _69580_/A _72800_/A _69592_/X sky130_fd_sc_hd__and2_4
X_81870_ _81883_/CLK _78061_/X _81870_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_356_0_CLK clkbuf_9_178_0_CLK/X _85712_/CLK sky130_fd_sc_hd__clkbuf_1
X_49709_ _49704_/Y _49706_/X _49708_/X _86338_/D sky130_fd_sc_hd__a21oi_4
X_68543_ _68542_/X _68543_/B _68543_/X sky130_fd_sc_hd__and2_4
X_80821_ _80821_/CLK _80821_/D _75599_/B sky130_fd_sc_hd__dfxtp_4
X_65755_ _65752_/X _65741_/B _65754_/X _65756_/B sky130_fd_sc_hd__nand3_4
X_50981_ _50971_/A _50981_/B _50981_/Y sky130_fd_sc_hd__nand2_4
X_62967_ _62967_/A _63326_/A _62939_/X _62967_/D _62967_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_986_0_CLK clkbuf_9_493_0_CLK/X _83306_/CLK sky130_fd_sc_hd__clkbuf_1
X_52720_ _52704_/A _52724_/B _52708_/X _52720_/D _52720_/X sky130_fd_sc_hd__and4_4
X_64706_ _64706_/A _64980_/A sky130_fd_sc_hd__buf_2
X_83540_ _86570_/CLK _83540_/D _83540_/Q sky130_fd_sc_hd__dfxtp_4
X_80752_ _81041_/CLK _75285_/X _81128_/D sky130_fd_sc_hd__dfxtp_4
X_61918_ _57670_/A _61902_/X _61916_/X _61870_/X _61917_/X _61918_/X
+ sky130_fd_sc_hd__a41o_4
X_68474_ _68474_/A _69004_/A sky130_fd_sc_hd__buf_2
X_65686_ _65486_/A _65702_/A sky130_fd_sc_hd__buf_2
X_62898_ _58490_/A _60304_/A _64454_/A _62875_/X _62898_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_9_477_0_CLK clkbuf_8_238_0_CLK/X clkbuf_9_477_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_67425_ _67166_/X _67413_/Y _67390_/X _67424_/Y _67425_/X sky130_fd_sc_hd__a211o_4
X_52651_ _52637_/A _52651_/B _52651_/Y sky130_fd_sc_hd__nand2_4
X_64637_ _66104_/A _64637_/X sky130_fd_sc_hd__buf_2
X_83471_ _85959_/CLK _83471_/D _47771_/A sky130_fd_sc_hd__dfxtp_4
X_61849_ _61865_/A _61865_/B _78073_/B _61849_/Y sky130_fd_sc_hd__nor3_4
X_80683_ _80679_/CLK _80683_/D _80683_/Q sky130_fd_sc_hd__dfxtp_4
X_85210_ _85180_/CLK _85210_/D _56395_/C sky130_fd_sc_hd__dfxtp_4
X_51602_ _51629_/A _51619_/A sky130_fd_sc_hd__buf_2
X_82422_ _82833_/CLK _82454_/Q _78608_/A sky130_fd_sc_hd__dfxtp_4
X_55370_ _55443_/A _55367_/Y _55443_/C _55370_/X sky130_fd_sc_hd__a21bo_4
X_67356_ _67333_/A _67356_/B _67356_/X sky130_fd_sc_hd__and2_4
X_86190_ _86506_/CLK _86190_/D _86190_/Q sky130_fd_sc_hd__dfxtp_4
X_64568_ _64667_/A _64611_/A sky130_fd_sc_hd__buf_2
X_52582_ _52590_/A _46624_/Y _52582_/Y sky130_fd_sc_hd__nand2_4
XPHY_607 sky130_fd_sc_hd__decap_3
XPHY_618 sky130_fd_sc_hd__decap_3
X_54321_ _54321_/A _54322_/A sky130_fd_sc_hd__buf_2
X_66307_ _66305_/Y _66278_/X _66306_/X _84142_/D sky130_fd_sc_hd__a21o_4
XPHY_629 sky130_fd_sc_hd__decap_3
X_85141_ _85057_/CLK _85141_/D _55499_/B sky130_fd_sc_hd__dfxtp_4
X_51533_ _51521_/X _51553_/B _51533_/C _53058_/D _51533_/X sky130_fd_sc_hd__and4_4
Xclkbuf_9_400_0_CLK clkbuf_8_200_0_CLK/X clkbuf_9_400_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_63519_ _63458_/A _63520_/C sky130_fd_sc_hd__buf_2
X_82353_ _87345_/CLK _77161_/X _82353_/Q sky130_fd_sc_hd__dfxtp_4
X_67287_ _67308_/A _67287_/B _67287_/X sky130_fd_sc_hd__and2_4
X_64499_ _64492_/Y _64498_/X _64442_/X _64499_/X sky130_fd_sc_hd__o21a_4
X_57040_ _57038_/X _46178_/X _57039_/Y _57040_/Y sky130_fd_sc_hd__a21oi_4
X_81304_ _81304_/CLK _76992_/X _81304_/Q sky130_fd_sc_hd__dfxtp_4
X_69026_ _69022_/X _69024_/X _69025_/X _69026_/X sky130_fd_sc_hd__a21o_4
X_54252_ _85476_/Q _54249_/X _54251_/Y _54252_/Y sky130_fd_sc_hd__o21ai_4
X_66238_ _66237_/X _66238_/B _66238_/X sky130_fd_sc_hd__and2_4
X_85072_ _85040_/CLK _85072_/D _45659_/A sky130_fd_sc_hd__dfxtp_4
X_51464_ _51481_/A _52991_/B _51464_/Y sky130_fd_sc_hd__nand2_4
X_82284_ _82284_/CLK _82284_/D _40879_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_924_0_CLK clkbuf_9_462_0_CLK/X _83145_/CLK sky130_fd_sc_hd__clkbuf_1
X_53203_ _53211_/A _53211_/B _53195_/X _53203_/D _53203_/X sky130_fd_sc_hd__and4_4
X_84023_ _82067_/CLK _68163_/X _84023_/Q sky130_fd_sc_hd__dfxtp_4
X_50415_ _86205_/Q _50387_/X _50414_/Y _50415_/Y sky130_fd_sc_hd__o21ai_4
X_81235_ _85332_/CLK _81043_/Q _47662_/A sky130_fd_sc_hd__dfxtp_4
X_54183_ _54180_/Y _54171_/X _54182_/X _85489_/D sky130_fd_sc_hd__a21oi_4
X_66169_ _64971_/X _85615_/Q _44261_/X _66168_/X _66169_/X sky130_fd_sc_hd__a211o_4
X_51395_ _65413_/B _51387_/X _51394_/Y _51395_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_415_0_CLK clkbuf_9_415_0_CLK/A clkbuf_9_415_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_53134_ _53132_/Y _53111_/X _53133_/X _53134_/Y sky130_fd_sc_hd__a21oi_4
X_50346_ _86219_/Q _50333_/X _50345_/Y _50346_/Y sky130_fd_sc_hd__o21ai_4
X_81166_ _81125_/CLK _74935_/B _81166_/Q sky130_fd_sc_hd__dfxtp_4
X_58991_ _58990_/Y _58988_/B _58991_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_309_0_CLK clkbuf_9_154_0_CLK/X _85491_/CLK sky130_fd_sc_hd__clkbuf_1
X_80117_ _80103_/Y _80117_/B _80117_/X sky130_fd_sc_hd__and2_4
X_53065_ _53065_/A _53065_/X sky130_fd_sc_hd__buf_2
X_57942_ _57938_/Y _57941_/Y _57909_/X _57942_/X sky130_fd_sc_hd__a21o_4
X_69928_ _83886_/Q _69894_/X _69927_/X _69928_/X sky130_fd_sc_hd__a21bo_4
X_50277_ _50251_/X _47932_/B _50277_/Y sky130_fd_sc_hd__nand2_4
X_85974_ _85974_/CLK _85974_/D _85974_/Q sky130_fd_sc_hd__dfxtp_4
X_81097_ _80679_/CLK _79633_/X _81097_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_939_0_CLK clkbuf_9_469_0_CLK/X _87553_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_0_0_CLK clkbuf_6_1_0_CLK/A clkbuf_6_0_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_52016_ _66141_/B _52013_/X _52015_/Y _52016_/Y sky130_fd_sc_hd__o21ai_4
X_87713_ _87210_/CLK _42798_/Y _87713_/Q sky130_fd_sc_hd__dfxtp_4
X_84925_ _84922_/CLK _84925_/D _84925_/Q sky130_fd_sc_hd__dfxtp_4
X_80048_ _84934_/Q _84182_/Q _80048_/X sky130_fd_sc_hd__xor2_4
X_57873_ _57868_/X _57870_/Y _57871_/Y _57822_/X _57872_/X _57873_/X
+ sky130_fd_sc_hd__o32a_4
X_69859_ _69859_/A _69860_/B sky130_fd_sc_hd__inv_2
X_59612_ _59611_/X _60626_/A sky130_fd_sc_hd__buf_2
X_56824_ _45835_/A _56824_/X sky130_fd_sc_hd__buf_2
X_87644_ _87644_/CLK _42933_/X _87644_/Q sky130_fd_sc_hd__dfxtp_4
X_72870_ _73378_/A _72870_/X sky130_fd_sc_hd__buf_2
X_84856_ _84263_/CLK _84856_/D _84856_/Q sky130_fd_sc_hd__dfxtp_4
X_71821_ _70504_/A _71779_/B _71049_/A _71821_/X sky130_fd_sc_hd__and3_4
X_59543_ _59543_/A _59544_/D sky130_fd_sc_hd__buf_2
X_83807_ _83813_/CLK _83807_/D _83807_/Q sky130_fd_sc_hd__dfxtp_4
X_56755_ _56679_/B _56755_/X sky130_fd_sc_hd__buf_2
X_87575_ _88326_/CLK _87575_/D _74206_/A sky130_fd_sc_hd__dfxtp_4
X_41981_ _41965_/X _41975_/X _40767_/X _41980_/Y _41967_/X _88083_/D
+ sky130_fd_sc_hd__o32ai_4
X_53967_ _85532_/Q _53940_/X _53966_/Y _53967_/Y sky130_fd_sc_hd__o21ai_4
X_84787_ _84787_/CLK _58955_/Y _84787_/Q sky130_fd_sc_hd__dfxtp_4
X_81999_ _82288_/CLK _81999_/D _77098_/A sky130_fd_sc_hd__dfxtp_4
X_43720_ _43719_/X _43720_/Y sky130_fd_sc_hd__inv_2
X_55706_ _55703_/X _55705_/X _55138_/X _55706_/X sky130_fd_sc_hd__a21o_4
X_86526_ _86523_/CLK _86526_/D _72843_/B sky130_fd_sc_hd__dfxtp_4
X_74540_ _74549_/A _74541_/A sky130_fd_sc_hd__buf_2
X_40932_ _40932_/A _40932_/X sky130_fd_sc_hd__buf_2
X_52918_ _52910_/A _52918_/B _52918_/Y sky130_fd_sc_hd__nand2_4
X_71752_ _52944_/B _71737_/X _71751_/Y _71752_/Y sky130_fd_sc_hd__o21ai_4
X_59474_ _59474_/A _59478_/B _59474_/Y sky130_fd_sc_hd__nand2_4
X_83738_ _83736_/CLK _83738_/D _47359_/A sky130_fd_sc_hd__dfxtp_4
X_56686_ _85137_/Q _44253_/X _56686_/X sky130_fd_sc_hd__or2_4
X_53898_ _53898_/A _72072_/B _53898_/Y sky130_fd_sc_hd__nand2_4
X_70703_ _70866_/A _70703_/X sky130_fd_sc_hd__buf_2
X_58425_ _58425_/A _58984_/A sky130_fd_sc_hd__buf_2
X_43651_ _87326_/Q _68888_/B sky130_fd_sc_hd__inv_2
X_55637_ _44087_/B _45393_/Y _55637_/Y sky130_fd_sc_hd__nor2_4
X_74471_ _83059_/Q _74441_/X _74470_/Y _74471_/Y sky130_fd_sc_hd__o21ai_4
X_86457_ _83303_/CLK _86457_/D _86457_/Q sky130_fd_sc_hd__dfxtp_4
X_52849_ _52767_/A _52850_/A sky130_fd_sc_hd__buf_2
X_40863_ _40862_/Y _40863_/Y sky130_fd_sc_hd__inv_2
X_71683_ _71570_/X _71626_/B _71289_/B _71683_/Y sky130_fd_sc_hd__nor3_4
X_83669_ _86091_/CLK _70900_/Y _83669_/Q sky130_fd_sc_hd__dfxtp_4
X_76210_ _76196_/B _76210_/Y sky130_fd_sc_hd__inv_2
X_42602_ _42590_/X _42592_/X _40885_/X _69859_/A _42597_/X _42603_/A
+ sky130_fd_sc_hd__o32ai_4
X_73422_ _88313_/Q _73059_/X _73421_/X _73422_/Y sky130_fd_sc_hd__o21ai_4
X_85408_ _85505_/CLK _85408_/D _85408_/Q sky130_fd_sc_hd__dfxtp_4
X_46370_ _86743_/Q _46364_/X _46369_/Y _46370_/Y sky130_fd_sc_hd__o21ai_4
X_70634_ _70633_/X _70635_/A sky130_fd_sc_hd__buf_2
X_58356_ _58151_/A _58356_/B _58356_/Y sky130_fd_sc_hd__nor2_4
X_77190_ _77202_/A _77189_/Y _77191_/B sky130_fd_sc_hd__xor2_4
X_43582_ _46612_/A _40591_/C _43175_/C _48144_/A sky130_fd_sc_hd__and3_4
X_55568_ _45494_/A _55527_/X _44098_/X _55567_/X _55568_/X sky130_fd_sc_hd__a211o_4
X_86388_ _83676_/CLK _49437_/Y _86388_/Q sky130_fd_sc_hd__dfxtp_4
X_40794_ _40756_/A _40794_/X sky130_fd_sc_hd__buf_2
X_45321_ _63312_/B _61649_/B sky130_fd_sc_hd__buf_2
X_57307_ _85037_/Q _56997_/X _57307_/Y sky130_fd_sc_hd__nor2_4
X_88127_ _87116_/CLK _41843_/Y _88127_/Q sky130_fd_sc_hd__dfxtp_4
X_76141_ _76143_/B _76143_/A _76142_/B sky130_fd_sc_hd__xor2_4
X_42533_ _42532_/Y _87831_/D sky130_fd_sc_hd__inv_2
X_54519_ _85427_/Q _54512_/X _54518_/Y _54519_/Y sky130_fd_sc_hd__o21ai_4
X_73353_ _73353_/A _85866_/Q _73353_/X sky130_fd_sc_hd__and2_4
X_85339_ _85372_/CLK _54993_/Y _85339_/Q sky130_fd_sc_hd__dfxtp_4
X_70565_ _70532_/Y _83748_/Q _70564_/Y _83748_/D sky130_fd_sc_hd__a21o_4
X_58287_ _58287_/A _58287_/Y sky130_fd_sc_hd__inv_2
X_55499_ _55826_/A _55499_/B _55499_/X sky130_fd_sc_hd__and2_4
X_48040_ _57590_/B _52036_/B sky130_fd_sc_hd__buf_2
X_72304_ _72299_/X _72301_/Y _72302_/Y _72194_/X _72303_/X _72304_/X
+ sky130_fd_sc_hd__o32a_4
X_45252_ _45252_/A _45252_/X sky130_fd_sc_hd__buf_2
X_57238_ _57235_/Y _57238_/X sky130_fd_sc_hd__buf_2
X_76072_ _76067_/Y _76068_/A _76071_/Y _76073_/B sky130_fd_sc_hd__a21boi_4
X_88058_ _88062_/CLK _88058_/D _88058_/Q sky130_fd_sc_hd__dfxtp_4
X_42464_ _42460_/X _42049_/X _40590_/X _68440_/B _42463_/X _42464_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73284_ _73284_/A _73284_/X sky130_fd_sc_hd__buf_2
X_70496_ _70496_/A _71115_/C sky130_fd_sc_hd__buf_2
X_44203_ _44201_/Y _44202_/X _44220_/B _87182_/D sky130_fd_sc_hd__a21oi_4
X_75023_ _75023_/A _75023_/B _75024_/B sky130_fd_sc_hd__xnor2_4
X_79900_ _84922_/Q _65901_/C _79900_/X sky130_fd_sc_hd__or2_4
X_87009_ _88283_/CLK _87009_/D _87009_/Q sky130_fd_sc_hd__dfxtp_4
X_41415_ _41412_/X _82889_/Q _41414_/X _41415_/Y sky130_fd_sc_hd__o21ai_4
X_72235_ _72224_/Y _72152_/X _72231_/X _72234_/X _83272_/D sky130_fd_sc_hd__a22oi_4
X_45183_ _45180_/X _45182_/Y _45125_/X _45183_/Y sky130_fd_sc_hd__a21oi_4
X_57169_ _56737_/X _56800_/X _56810_/X _57156_/X _56767_/X _57169_/X
+ sky130_fd_sc_hd__a41o_4
X_42395_ _40408_/X _42388_/X _87883_/Q _42389_/X _87883_/D sky130_fd_sc_hd__a2bb2o_4
X_44134_ _44196_/A _44196_/B _44128_/X _44134_/D _44134_/X sky130_fd_sc_hd__and4_4
X_79831_ _79819_/A _79818_/Y _79830_/X _79831_/X sky130_fd_sc_hd__a21o_4
X_41346_ _41344_/X _81750_/Q _41345_/X _41346_/X sky130_fd_sc_hd__o21a_4
X_60180_ _60179_/Y _60291_/C sky130_fd_sc_hd__buf_2
X_72166_ _57708_/X _72166_/X sky130_fd_sc_hd__buf_2
X_49991_ _49989_/Y _49977_/X _49990_/X _86286_/D sky130_fd_sc_hd__a21oi_4
X_71117_ _71117_/A _71117_/X sky130_fd_sc_hd__buf_2
X_48942_ _83619_/Q _71987_/B sky130_fd_sc_hd__inv_2
X_44065_ _44064_/X _44086_/A sky130_fd_sc_hd__buf_2
X_79762_ _64942_/C _72263_/Y _79761_/Y _79762_/X sky130_fd_sc_hd__o21a_4
X_41277_ _41276_/X _41277_/X sky130_fd_sc_hd__buf_2
X_76974_ _61055_/C _84398_/Q _76974_/X sky130_fd_sc_hd__xor2_4
X_72097_ _83285_/Q _72090_/X _72096_/Y _72097_/Y sky130_fd_sc_hd__o21ai_4
X_43016_ _43030_/A _43017_/A sky130_fd_sc_hd__buf_2
X_78713_ _78709_/Y _78713_/B _78712_/Y _78713_/X sky130_fd_sc_hd__or3_4
X_71048_ _70832_/A _71049_/A sky130_fd_sc_hd__buf_2
X_75925_ _81506_/Q _75925_/B _75925_/X sky130_fd_sc_hd__xor2_4
X_48873_ _86466_/Q _48861_/X _48872_/Y _48873_/Y sky130_fd_sc_hd__o21ai_4
X_79693_ _79689_/Y _79692_/Y _79704_/A sky130_fd_sc_hd__xor2_4
X_47824_ _47820_/Y _47791_/X _47823_/X _86594_/D sky130_fd_sc_hd__a21oi_4
X_78644_ _78644_/A _82776_/D _82488_/D sky130_fd_sc_hd__xor2_4
X_63870_ _60871_/Y _63920_/B sky130_fd_sc_hd__buf_2
X_75856_ _75830_/B _80798_/D sky130_fd_sc_hd__inv_2
X_62821_ _62773_/X _62812_/B _61954_/X _62821_/Y sky130_fd_sc_hd__nand3_4
X_74807_ _74807_/A _74775_/A _70884_/A _70662_/X _74810_/B sky130_fd_sc_hd__nand4_4
X_47755_ _47661_/A _47777_/C sky130_fd_sc_hd__buf_2
X_78575_ _78575_/A _78575_/B _78575_/X sky130_fd_sc_hd__and2_4
X_44967_ _45193_/A _45734_/A sky130_fd_sc_hd__buf_2
X_75787_ _75787_/A _75786_/X _75793_/A sky130_fd_sc_hd__xor2_4
X_72999_ _83169_/Q _72943_/X _72998_/X _72999_/X sky130_fd_sc_hd__a21o_4
X_46706_ _82968_/Q _46706_/Y sky130_fd_sc_hd__inv_2
X_65540_ _65407_/A _65540_/X sky130_fd_sc_hd__buf_2
X_77526_ _77522_/Y _77501_/Y _77525_/X _77526_/Y sky130_fd_sc_hd__o21ai_4
X_43918_ _43916_/X _43902_/X _41387_/X _87200_/Q _43917_/X _43918_/Y
+ sky130_fd_sc_hd__o32ai_4
X_62752_ _60273_/A _62762_/B sky130_fd_sc_hd__buf_2
X_74738_ _74738_/A _74740_/B sky130_fd_sc_hd__inv_2
X_47686_ _83552_/Q _54880_/B sky130_fd_sc_hd__inv_2
X_44898_ _45757_/A _44898_/X sky130_fd_sc_hd__buf_2
X_49425_ _49420_/A _49447_/B _49420_/C _46728_/X _49425_/X sky130_fd_sc_hd__and4_4
X_61703_ _61770_/A _61770_/B _59477_/A _61770_/D _61703_/X sky130_fd_sc_hd__and4_4
X_46637_ _46637_/A _46638_/A sky130_fd_sc_hd__inv_2
X_65471_ _65592_/A _72840_/B _65471_/X sky130_fd_sc_hd__and2_4
X_77457_ _77455_/Y _77456_/X _77458_/B sky130_fd_sc_hd__xor2_4
X_43849_ _43848_/Y _87236_/D sky130_fd_sc_hd__inv_2
X_62683_ _61356_/X _62694_/B _62694_/C _62664_/D _62683_/Y sky130_fd_sc_hd__nand4_4
X_74669_ _74669_/A _82991_/D sky130_fd_sc_hd__inv_2
X_67210_ _80903_/D _67092_/X _67209_/X _67210_/X sky130_fd_sc_hd__a21bo_4
X_64422_ _64402_/X _64421_/X _64422_/C _64422_/X sky130_fd_sc_hd__and3_4
X_76408_ _81652_/Q _76408_/Y sky130_fd_sc_hd__inv_2
X_49356_ _49302_/A _51394_/B _49356_/Y sky130_fd_sc_hd__nand2_4
X_61634_ _61634_/A _61634_/B _79132_/B _61634_/Y sky130_fd_sc_hd__nor3_4
X_68190_ _67181_/X _67184_/X _68169_/X _68190_/Y sky130_fd_sc_hd__a21oi_4
X_46568_ _46525_/X _81189_/Q _46567_/X _51380_/B sky130_fd_sc_hd__o21ai_4
X_77388_ _77396_/B _77374_/B _77387_/X _77388_/Y sky130_fd_sc_hd__o21ai_4
X_48307_ _48079_/B _57609_/B sky130_fd_sc_hd__buf_2
X_67141_ _64608_/A _67141_/X sky130_fd_sc_hd__buf_2
X_79127_ _79127_/A _61690_/C _79127_/X sky130_fd_sc_hd__xor2_4
X_45519_ _57397_/B _45519_/Y sky130_fd_sc_hd__inv_2
X_64353_ _64319_/X _64353_/B _64333_/X _64353_/X sky130_fd_sc_hd__and3_4
X_76339_ _76313_/X _76317_/B _76339_/X sky130_fd_sc_hd__xor2_4
X_49287_ _49287_/A _51316_/B _49287_/Y sky130_fd_sc_hd__nand2_4
X_61565_ _61558_/Y _61560_/Y _61525_/X _61561_/Y _61564_/Y _61565_/X
+ sky130_fd_sc_hd__a41o_4
X_46499_ _46492_/Y _46445_/X _46498_/X _46499_/Y sky130_fd_sc_hd__a21oi_4
X_63304_ _44173_/X _63528_/A sky130_fd_sc_hd__buf_2
X_48238_ _47957_/B _53516_/B sky130_fd_sc_hd__buf_2
X_60516_ _60435_/A _60516_/B _60515_/Y _60516_/Y sky130_fd_sc_hd__nand3_4
X_67072_ _87358_/Q _66997_/X _66998_/X _67071_/X _67072_/X sky130_fd_sc_hd__a211o_4
X_79058_ _79058_/A _79058_/B _82621_/D sky130_fd_sc_hd__nand2_4
X_64284_ _64275_/A _64284_/B _64274_/X _64284_/X sky130_fd_sc_hd__and3_4
X_61496_ _61518_/A _61518_/B _84476_/Q _61496_/Y sky130_fd_sc_hd__nor3_4
X_66023_ _65990_/X _86233_/Q _66021_/X _66022_/X _66023_/X sky130_fd_sc_hd__a211o_4
X_78009_ _78009_/A _78024_/A _78018_/A sky130_fd_sc_hd__xnor2_4
X_63235_ _63118_/A _63235_/X sky130_fd_sc_hd__buf_2
X_48169_ _48897_/A _48169_/X sky130_fd_sc_hd__buf_2
X_60447_ _60447_/A _60447_/B _60515_/A _60529_/B sky130_fd_sc_hd__nor3_4
X_50200_ _86244_/Q _50185_/X _50199_/Y _50200_/Y sky130_fd_sc_hd__o21ai_4
X_81020_ _84150_/CLK _84228_/Q _81020_/Q sky130_fd_sc_hd__dfxtp_4
X_51180_ _86059_/Q _51156_/X _51179_/Y _51180_/Y sky130_fd_sc_hd__o21ai_4
X_63166_ _63154_/X _64378_/B _63165_/X _63121_/D _63166_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_280_0_CLK clkbuf_9_140_0_CLK/X _83482_/CLK sky130_fd_sc_hd__clkbuf_1
X_60378_ _60639_/A _59536_/A _61285_/C _60378_/Y sky130_fd_sc_hd__nand3_4
X_50131_ _50131_/A _53858_/B _50131_/X sky130_fd_sc_hd__and2_4
X_62117_ _62088_/B _62117_/X sky130_fd_sc_hd__buf_2
X_67974_ _66554_/X _68044_/A sky130_fd_sc_hd__buf_2
X_63097_ _63097_/A _64305_/B _63085_/C _63085_/D _63097_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_62_0_CLK clkbuf_9_31_0_CLK/X _85034_/CLK sky130_fd_sc_hd__clkbuf_1
X_69713_ _69680_/A _88328_/Q _69713_/X sky130_fd_sc_hd__and2_4
X_50062_ _47832_/A _50063_/A sky130_fd_sc_hd__buf_2
X_66925_ _66563_/A _67046_/A sky130_fd_sc_hd__buf_2
X_62048_ _61719_/A _62048_/X sky130_fd_sc_hd__buf_2
X_82971_ _82394_/CLK _82779_/Q _46680_/A sky130_fd_sc_hd__dfxtp_4
X_84710_ _84355_/CLK _59703_/Y _80588_/A sky130_fd_sc_hd__dfxtp_4
X_69644_ _64732_/A _69644_/X sky130_fd_sc_hd__buf_2
X_81922_ _82145_/CLK _81922_/D _81922_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_107_0_CLK clkbuf_6_53_0_CLK/X clkbuf_8_215_0_CLK/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_295_0_CLK clkbuf_9_147_0_CLK/X _83402_/CLK sky130_fd_sc_hd__clkbuf_1
X_54870_ _54868_/Y _54856_/X _54869_/X _54870_/Y sky130_fd_sc_hd__a21oi_4
X_66856_ _66853_/X _66855_/X _66787_/X _66859_/A sky130_fd_sc_hd__a21o_4
X_85690_ _85688_/CLK _85690_/D _85690_/Q sky130_fd_sc_hd__dfxtp_4
X_53821_ _71994_/B _53821_/B _53821_/Y sky130_fd_sc_hd__nand2_4
X_65807_ _65807_/A _86472_/Q _65807_/X sky130_fd_sc_hd__and2_4
X_84641_ _84620_/CLK _60287_/X _79797_/A sky130_fd_sc_hd__dfxtp_4
X_69575_ _69575_/A _69575_/X sky130_fd_sc_hd__buf_2
X_81853_ _82515_/CLK _81885_/Q _77630_/A sky130_fd_sc_hd__dfxtp_4
X_66787_ _66547_/A _66787_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_77_0_CLK clkbuf_9_38_0_CLK/X _84418_/CLK sky130_fd_sc_hd__clkbuf_1
X_63999_ _64401_/B _64029_/B _63951_/C _64015_/D _63999_/Y sky130_fd_sc_hd__nand4_4
X_56540_ _56538_/A _56535_/X _55724_/B _56540_/Y sky130_fd_sc_hd__nand3_4
X_80804_ _80804_/CLK _80804_/D _75733_/B sky130_fd_sc_hd__dfxtp_4
X_68526_ _66560_/X _69007_/A sky130_fd_sc_hd__buf_2
X_87360_ _86796_/CLK _87360_/D _87360_/Q sky130_fd_sc_hd__dfxtp_4
X_53752_ _48849_/A _53748_/B _53748_/C _53752_/X sky130_fd_sc_hd__and3_4
Xclkbuf_8_223_0_CLK clkbuf_8_223_0_CLK/A clkbuf_9_446_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_65738_ _64834_/A _65741_/B sky130_fd_sc_hd__buf_2
X_84572_ _84583_/CLK _60764_/Y _84572_/Q sky130_fd_sc_hd__dfxtp_4
X_50964_ _50962_/Y _50957_/X _50963_/X _50964_/Y sky130_fd_sc_hd__a21oi_4
X_81784_ _88121_/CLK _76136_/X _81784_/Q sky130_fd_sc_hd__dfxtp_4
X_86311_ _86627_/CLK _86311_/D _58070_/B sky130_fd_sc_hd__dfxtp_4
X_52703_ _52648_/A _52704_/A sky130_fd_sc_hd__buf_2
X_83523_ _83526_/CLK _71367_/X _83523_/Q sky130_fd_sc_hd__dfxtp_4
X_56471_ _56448_/X _56472_/B sky130_fd_sc_hd__buf_2
X_68457_ _87100_/Q _68455_/X _68370_/X _68456_/X _68457_/X sky130_fd_sc_hd__a211o_4
X_80735_ _82211_/CLK _80735_/D _80703_/D sky130_fd_sc_hd__dfxtp_4
X_87291_ _87553_/CLK _87291_/D _43732_/A sky130_fd_sc_hd__dfxtp_4
X_53683_ _53662_/X _74428_/B _53683_/Y sky130_fd_sc_hd__nand2_4
X_65669_ _65669_/A _65669_/X sky130_fd_sc_hd__buf_2
X_50895_ _46616_/A _51033_/A sky130_fd_sc_hd__buf_2
X_58210_ _64544_/C _58210_/X sky130_fd_sc_hd__buf_2
X_55422_ _56807_/A _56807_/C _55422_/Y sky130_fd_sc_hd__nand2_4
X_86242_ _83594_/CLK _50210_/Y _86242_/Q sky130_fd_sc_hd__dfxtp_4
X_67408_ _67381_/A _87216_/Q _67408_/X sky130_fd_sc_hd__and2_4
X_52634_ _52605_/A _52654_/B sky130_fd_sc_hd__buf_2
X_59190_ _59152_/X _59188_/Y _59189_/Y _59169_/X _59156_/X _59190_/X
+ sky130_fd_sc_hd__o32a_4
X_83454_ _83457_/CLK _71566_/X _83454_/Q sky130_fd_sc_hd__dfxtp_4
X_80666_ _84407_/CLK _74843_/Y _80666_/Q sky130_fd_sc_hd__dfxtp_4
X_68388_ _73577_/A _68384_/X _68385_/X _68387_/Y _68388_/X sky130_fd_sc_hd__a211o_4
XPHY_404 sky130_fd_sc_hd__decap_3
X_58141_ _58065_/X _85698_/Q _58089_/X _58141_/X sky130_fd_sc_hd__o21a_4
X_82405_ _82443_/CLK _82437_/Q _78344_/A sky130_fd_sc_hd__dfxtp_4
XPHY_415 sky130_fd_sc_hd__decap_3
Xclkbuf_8_238_0_CLK clkbuf_8_239_0_CLK/A clkbuf_8_238_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_55353_ _55445_/A _55445_/C _55353_/X sky130_fd_sc_hd__and2_4
X_67339_ _86975_/Q _67311_/X _67313_/X _67338_/X _67339_/X sky130_fd_sc_hd__a211o_4
X_86173_ _83307_/CLK _50585_/Y _86173_/Q sky130_fd_sc_hd__dfxtp_4
X_52565_ _52280_/X _52565_/B _52565_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_233_0_CLK clkbuf_9_116_0_CLK/X _81121_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_426 sky130_fd_sc_hd__decap_3
X_83385_ _83415_/CLK _83385_/D _83385_/Q sky130_fd_sc_hd__dfxtp_4
X_80597_ _80596_/B _80596_/A _80566_/Y _80570_/B _80598_/C sky130_fd_sc_hd__a211o_4
XPHY_437 sky130_fd_sc_hd__decap_3
XPHY_448 sky130_fd_sc_hd__decap_3
X_54304_ _54301_/Y _54285_/X _54303_/X _54304_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_863_0_CLK clkbuf_9_431_0_CLK/X _85527_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_459 sky130_fd_sc_hd__decap_3
X_85124_ _82979_/CLK _85124_/D _56898_/A sky130_fd_sc_hd__dfxtp_4
X_51516_ _51509_/A _51527_/B _51522_/C _53044_/D _51516_/X sky130_fd_sc_hd__and4_4
X_70350_ _70348_/A _70348_/B _83082_/Q _70348_/D _70350_/X sky130_fd_sc_hd__and4_4
X_58072_ _58010_/X _58070_/Y _58071_/Y _58028_/X _58015_/X _58072_/X
+ sky130_fd_sc_hd__o32a_4
X_82336_ _83974_/CLK _77220_/B _82336_/Q sky130_fd_sc_hd__dfxtp_4
X_55284_ _56868_/A _56868_/B _55671_/A _55284_/X sky130_fd_sc_hd__a21o_4
X_52496_ _52496_/A _52496_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_15_0_CLK clkbuf_9_7_0_CLK/X _85311_/CLK sky130_fd_sc_hd__clkbuf_1
X_57023_ _57023_/A _57023_/X sky130_fd_sc_hd__buf_2
X_69009_ _87993_/Q _69007_/X _68916_/X _69008_/X _69009_/X sky130_fd_sc_hd__a211o_4
X_54235_ _85479_/Q _54220_/X _54234_/Y _54235_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_354_0_CLK clkbuf_9_355_0_CLK/A clkbuf_9_354_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_85055_ _85152_/CLK _85055_/D _45426_/A sky130_fd_sc_hd__dfxtp_4
X_51447_ _51010_/A _51557_/A sky130_fd_sc_hd__buf_2
X_70281_ _74762_/A _70157_/A _70280_/Y _83812_/D sky130_fd_sc_hd__o21ai_4
X_82267_ _83515_/CLK _82267_/D _82267_/Q sky130_fd_sc_hd__dfxtp_4
X_41200_ _41199_/X _41181_/X _68775_/B _41182_/X _88259_/D sky130_fd_sc_hd__a2bb2o_4
X_72020_ _71993_/X _53844_/B _72020_/Y sky130_fd_sc_hd__nand2_4
X_84006_ _81746_/CLK _84006_/D _84006_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_248_0_CLK clkbuf_9_124_0_CLK/X _82221_/CLK sky130_fd_sc_hd__clkbuf_1
X_81218_ _85315_/CLK _81026_/Q _81218_/Q sky130_fd_sc_hd__dfxtp_4
X_54166_ _54163_/Y _54144_/X _54165_/X _85492_/D sky130_fd_sc_hd__a21oi_4
X_42180_ _42180_/A _87995_/D sky130_fd_sc_hd__inv_2
X_51378_ _51364_/A _51378_/B _51378_/Y sky130_fd_sc_hd__nand2_4
X_82198_ _82390_/CLK _82198_/D _82390_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_878_0_CLK clkbuf_9_439_0_CLK/X _86592_/CLK sky130_fd_sc_hd__clkbuf_1
X_41131_ _41130_/X _41109_/X _88272_/Q _41110_/X _41131_/X sky130_fd_sc_hd__a2bb2o_4
X_53117_ _53195_/A _53133_/C sky130_fd_sc_hd__buf_2
X_50329_ _86222_/Q _50238_/X _50328_/Y _50329_/Y sky130_fd_sc_hd__o21ai_4
X_81149_ _82284_/CLK _81149_/D _81149_/Q sky130_fd_sc_hd__dfxtp_4
X_54097_ _53434_/A _54097_/B _54097_/Y sky130_fd_sc_hd__nand2_4
X_58974_ _58559_/X _83440_/Q _58973_/Y _84784_/D sky130_fd_sc_hd__o21a_4
Xclkbuf_9_369_0_CLK clkbuf_8_184_0_CLK/X clkbuf_9_369_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_41062_ _40937_/A _41062_/B _41062_/X sky130_fd_sc_hd__or2_4
X_53048_ _53048_/A _53063_/B _53058_/C _53048_/D _53048_/X sky130_fd_sc_hd__and4_4
X_57925_ _57760_/X _85395_/Q _57924_/X _57925_/Y sky130_fd_sc_hd__o21ai_4
X_73971_ _73850_/X _86224_/Q _73948_/X _73970_/X _73971_/X sky130_fd_sc_hd__a211o_4
X_85957_ _85957_/CLK _85957_/D _85957_/Q sky130_fd_sc_hd__dfxtp_4
X_75710_ _75704_/B _75696_/X _75709_/Y _75710_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_801_0_CLK clkbuf_9_400_0_CLK/X _82604_/CLK sky130_fd_sc_hd__clkbuf_1
X_72922_ _87821_/Q _73000_/B _72922_/Y sky130_fd_sc_hd__nor2_4
X_84908_ _84903_/CLK _84908_/D _64534_/C sky130_fd_sc_hd__dfxtp_4
X_45870_ _85026_/Q _45870_/Y sky130_fd_sc_hd__inv_2
X_57856_ _84945_/Q _57819_/X _57847_/X _57855_/X _57856_/Y sky130_fd_sc_hd__a2bb2oi_4
X_76690_ _81687_/Q _76690_/B _81351_/D sky130_fd_sc_hd__xor2_4
X_85888_ _85888_/CLK _52104_/Y _65439_/B sky130_fd_sc_hd__dfxtp_4
X_44821_ _46001_/A _44821_/X sky130_fd_sc_hd__buf_2
X_56807_ _56807_/A _46237_/A _56807_/C _57029_/A sky130_fd_sc_hd__nand3_4
X_87627_ _87883_/CLK _87627_/D _87627_/Q sky130_fd_sc_hd__dfxtp_4
X_75641_ _75641_/A _75641_/B _75641_/Y sky130_fd_sc_hd__nand2_4
X_72853_ _72852_/X _72853_/X sky130_fd_sc_hd__buf_2
X_84839_ _84839_/CLK _84839_/D _64422_/C sky130_fd_sc_hd__dfxtp_4
X_57787_ _64567_/A _64616_/A sky130_fd_sc_hd__buf_2
X_54999_ _54973_/A _55013_/C sky130_fd_sc_hd__buf_2
X_47540_ _47540_/A _53107_/D sky130_fd_sc_hd__buf_2
X_71804_ _71804_/A _71804_/Y sky130_fd_sc_hd__inv_2
X_59526_ _60385_/A _59602_/C sky130_fd_sc_hd__inv_2
X_78360_ _78360_/A _78360_/B _78376_/B _78364_/C sky130_fd_sc_hd__nand3_4
X_44752_ _41294_/A _44665_/X _86974_/Q _44666_/X _44752_/X sky130_fd_sc_hd__a2bb2o_4
X_56738_ _56737_/X _56738_/X sky130_fd_sc_hd__buf_2
X_75572_ _80818_/Q _75573_/A sky130_fd_sc_hd__inv_2
X_87558_ _87553_/CLK _87558_/D _73108_/A sky130_fd_sc_hd__dfxtp_4
X_41964_ _41937_/X _41956_/X _40729_/X _41963_/Y _41939_/X _88090_/D
+ sky130_fd_sc_hd__o32ai_4
X_72784_ _72784_/A _73238_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_816_0_CLK clkbuf_9_408_0_CLK/X _82675_/CLK sky130_fd_sc_hd__clkbuf_1
X_77311_ _77311_/A _77308_/A _77307_/A _77315_/B sky130_fd_sc_hd__nand3_4
X_43703_ _43703_/A _69737_/B sky130_fd_sc_hd__inv_2
X_74523_ _74523_/A _74518_/B _70880_/C _74531_/D _74523_/Y sky130_fd_sc_hd__nand4_4
X_86509_ _85859_/CLK _86509_/D _86509_/Q sky130_fd_sc_hd__dfxtp_4
X_40915_ _40568_/A _40995_/A sky130_fd_sc_hd__buf_2
X_47471_ _86631_/Q _47429_/X _47470_/Y _47471_/Y sky130_fd_sc_hd__o21ai_4
X_71735_ _71735_/A _71115_/D _71735_/C _71735_/D _71735_/X sky130_fd_sc_hd__and4_4
X_59457_ _58548_/A _59457_/B _59457_/Y sky130_fd_sc_hd__nor2_4
X_78291_ _78286_/B _78289_/X _78290_/Y _78291_/Y sky130_fd_sc_hd__a21boi_4
X_44683_ _44682_/Y _87002_/D sky130_fd_sc_hd__inv_2
X_56669_ _56774_/C _56725_/B sky130_fd_sc_hd__buf_2
X_87489_ _87758_/CLK _87489_/D _87489_/Q sky130_fd_sc_hd__dfxtp_4
X_41895_ _41894_/X _41879_/X _40605_/X _73650_/A _41882_/X _41895_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49210_ _49210_/A _49210_/B _53944_/C _49210_/Y sky130_fd_sc_hd__nor3_4
X_46422_ _86738_/Q _46292_/X _46421_/Y _46422_/Y sky130_fd_sc_hd__o21ai_4
X_58408_ _58408_/A _58415_/B sky130_fd_sc_hd__buf_2
Xclkbuf_9_307_0_CLK clkbuf_9_307_0_CLK/A clkbuf_9_307_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_77242_ _77233_/A _82082_/D _77242_/Y sky130_fd_sc_hd__nand2_4
X_43634_ _47834_/A _43634_/X sky130_fd_sc_hd__buf_2
X_74454_ _48567_/A _74478_/B _74425_/X _74454_/X sky130_fd_sc_hd__and3_4
X_40846_ _40845_/X _40821_/X _88324_/Q _40822_/X _88324_/D sky130_fd_sc_hd__a2bb2o_4
X_71666_ _70426_/A _71261_/B _71641_/A _71666_/Y sky130_fd_sc_hd__nand3_4
X_59388_ _59388_/A _58988_/B _59388_/Y sky130_fd_sc_hd__nand2_4
X_49141_ _50693_/A _50693_/B _48908_/A _49141_/X sky130_fd_sc_hd__o21a_4
X_73405_ _73402_/X _73404_/X _73262_/X _73409_/A sky130_fd_sc_hd__a21o_4
X_46353_ _46362_/A _53983_/B _46353_/Y sky130_fd_sc_hd__nand2_4
X_70617_ _70722_/A _70620_/B _70620_/C _70620_/D _70617_/Y sky130_fd_sc_hd__nand4_4
X_58339_ _58338_/Y _58364_/B _58339_/Y sky130_fd_sc_hd__nand2_4
X_77173_ _77173_/A _77173_/B _77173_/C _77173_/X sky130_fd_sc_hd__and3_4
X_43565_ _43564_/Y _43565_/Y sky130_fd_sc_hd__inv_2
X_74385_ _74391_/A _52119_/B _74385_/Y sky130_fd_sc_hd__nand2_4
X_40777_ _40776_/X _40754_/X _69597_/B _40756_/X _88337_/D sky130_fd_sc_hd__a2bb2o_4
X_71597_ _71528_/X _71626_/B sky130_fd_sc_hd__buf_2
X_45304_ _55761_/B _45269_/X _45303_/X _45304_/X sky130_fd_sc_hd__o21a_4
X_76124_ _76112_/A _76126_/A _76127_/B _76124_/Y sky130_fd_sc_hd__nand3_4
X_42516_ _42486_/X _42501_/X _40712_/X _68910_/B _42489_/X _42516_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49072_ _49072_/A _53877_/B sky130_fd_sc_hd__inv_2
X_73336_ _73333_/X _73335_/X _73336_/Y sky130_fd_sc_hd__nand2_4
X_61350_ _72592_/A _61384_/A sky130_fd_sc_hd__buf_2
X_46284_ _86750_/Q _46279_/X _46283_/Y _46284_/Y sky130_fd_sc_hd__o21ai_4
X_70548_ _71857_/A _71698_/A sky130_fd_sc_hd__buf_2
X_43496_ _43495_/X _43475_/X _41735_/X _87391_/Q _43479_/X _43497_/A
+ sky130_fd_sc_hd__o32ai_4
X_48023_ _48022_/Y _48024_/B sky130_fd_sc_hd__buf_2
X_60301_ _79775_/A _59822_/X _60299_/Y _60300_/Y _60301_/X sky130_fd_sc_hd__o22a_4
X_45235_ _45202_/X _61579_/B _45219_/X _45235_/Y sky130_fd_sc_hd__o21ai_4
X_76055_ _81717_/D _76056_/B _76063_/B sky130_fd_sc_hd__or2_4
X_42447_ _42447_/A _42447_/B _42447_/C _42447_/D _42447_/X sky130_fd_sc_hd__and4_4
X_61281_ _61281_/A _72625_/A _61281_/C _61281_/X sky130_fd_sc_hd__and3_4
X_73267_ _73267_/A _73266_/X _73267_/Y sky130_fd_sc_hd__nand2_4
X_70479_ _70387_/A _71815_/B sky130_fd_sc_hd__buf_2
X_63020_ _63020_/A _63020_/X sky130_fd_sc_hd__buf_2
X_75006_ _74999_/X _75005_/Y _75007_/B sky130_fd_sc_hd__xor2_4
X_60232_ _43969_/A _59899_/B _43969_/B _59899_/D _60232_/Y sky130_fd_sc_hd__nand4_4
X_72218_ _59368_/X _85977_/Q _72217_/X _72218_/Y sky130_fd_sc_hd__o21ai_4
X_45166_ _45163_/Y _45165_/Y _45137_/X _45166_/X sky130_fd_sc_hd__a21o_4
X_42378_ _42417_/A _42378_/X sky130_fd_sc_hd__buf_2
X_73198_ _73198_/A _73198_/B _73198_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_5_7_0_CLK clkbuf_5_7_0_CLK/A clkbuf_5_7_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_44117_ _44117_/A _87187_/Q _87186_/Q _44117_/Y sky130_fd_sc_hd__nand3_4
X_79814_ _84226_/Q _83274_/Q _79814_/Y sky130_fd_sc_hd__nand2_4
X_41329_ _41328_/X _41307_/X _88235_/Q _41308_/X _88235_/D sky130_fd_sc_hd__a2bb2o_4
X_60163_ _60162_/X _60387_/A sky130_fd_sc_hd__buf_2
X_72149_ _72145_/Y _72148_/Y _59351_/X _72149_/X sky130_fd_sc_hd__a21o_4
X_49974_ _49972_/Y _49951_/X _49973_/X _86289_/D sky130_fd_sc_hd__a21oi_4
X_45097_ _64353_/B _61479_/B sky130_fd_sc_hd__buf_2
X_48925_ _48881_/X _48405_/A _48924_/Y _48926_/A sky130_fd_sc_hd__o21ai_4
X_44048_ _44047_/X _44048_/X sky130_fd_sc_hd__buf_2
X_79745_ _79745_/A _79745_/Y sky130_fd_sc_hd__inv_2
X_64971_ _58124_/A _64971_/X sky130_fd_sc_hd__buf_2
X_60094_ _60174_/C _61070_/B _60094_/X sky130_fd_sc_hd__and2_4
X_76957_ _76957_/A _81601_/Q _76957_/C _76958_/B sky130_fd_sc_hd__nand3_4
X_66710_ _66689_/A _66710_/B _66710_/X sky130_fd_sc_hd__and2_4
X_63922_ _63916_/Y _63922_/B _63920_/Y _63922_/D _63922_/X sky130_fd_sc_hd__and4_4
X_75908_ _84506_/Q _84378_/Q _75908_/X sky130_fd_sc_hd__xor2_4
X_48856_ _48851_/A _48673_/B _48856_/Y sky130_fd_sc_hd__nand2_4
X_67690_ _68637_/A _67690_/X sky130_fd_sc_hd__buf_2
X_79676_ _79673_/X _79676_/B _79676_/X sky130_fd_sc_hd__xor2_4
X_76888_ _76888_/A _76888_/B _76888_/C _76889_/B sky130_fd_sc_hd__nand3_4
X_47807_ _47620_/X _47819_/A sky130_fd_sc_hd__buf_2
X_66641_ _87888_/Q _66639_/X _66531_/X _66640_/X _66641_/X sky130_fd_sc_hd__a211o_4
X_78627_ _82519_/Q _82775_/D _82487_/D sky130_fd_sc_hd__xor2_4
X_63853_ _61421_/A _63853_/B _63803_/C _63787_/D _63853_/Y sky130_fd_sc_hd__nand4_4
X_75839_ _75839_/A _75839_/B _75840_/B sky130_fd_sc_hd__xnor2_4
X_48787_ _48784_/Y _48785_/X _48786_/X _48787_/Y sky130_fd_sc_hd__a21oi_4
X_45999_ _45994_/X _45987_/X _40473_/X _66975_/B _45995_/X _45999_/Y
+ sky130_fd_sc_hd__o32ai_4
X_62804_ _62789_/A _63150_/A _62848_/C _62789_/D _62804_/X sky130_fd_sc_hd__and4_4
X_69360_ _69355_/X _69359_/X _69138_/X _69360_/X sky130_fd_sc_hd__a21o_4
X_47738_ _55078_/D _53217_/D sky130_fd_sc_hd__buf_2
X_66572_ _44174_/A _66572_/X sky130_fd_sc_hd__buf_2
X_78558_ _78557_/B _78556_/Y _78548_/X _78558_/X sky130_fd_sc_hd__o21a_4
X_63784_ _63800_/A _63800_/B _63784_/C _63784_/Y sky130_fd_sc_hd__nor3_4
X_60996_ _60863_/X _60996_/B _60915_/X _60996_/Y sky130_fd_sc_hd__nor3_4
X_68311_ _83986_/Q _68299_/X _68310_/X _83986_/D sky130_fd_sc_hd__a21bo_4
X_65523_ _65520_/X _65522_/X _65287_/X _65523_/X sky130_fd_sc_hd__a21o_4
X_77509_ _77505_/Y _77509_/B _77508_/Y _77511_/A sky130_fd_sc_hd__or3_4
X_62735_ _62766_/A _62766_/B _84387_/Q _62735_/Y sky130_fd_sc_hd__nor3_4
X_69291_ _69253_/A _88296_/Q _69291_/X sky130_fd_sc_hd__and2_4
X_47669_ _54871_/B _53179_/B sky130_fd_sc_hd__buf_2
X_78489_ _78489_/A _82671_/D _78489_/Y sky130_fd_sc_hd__nand2_4
X_49408_ _49420_/A _49420_/B _49408_/C _52622_/D _49408_/X sky130_fd_sc_hd__and4_4
X_80520_ _80504_/X _80520_/B _80520_/X sky130_fd_sc_hd__or2_4
X_68242_ _84003_/Q _68238_/X _68241_/X _68242_/X sky130_fd_sc_hd__a21bo_4
X_65454_ _65877_/A _65592_/A sky130_fd_sc_hd__buf_2
X_50680_ _50742_/A _50680_/X sky130_fd_sc_hd__buf_2
X_62666_ _62847_/A _62669_/A sky130_fd_sc_hd__buf_2
X_64405_ _58251_/A _64367_/X _64404_/Y _64405_/Y sky130_fd_sc_hd__o21ai_4
X_61617_ _61558_/A _61617_/B _61590_/C _61617_/Y sky130_fd_sc_hd__nand3_4
X_49339_ _49337_/Y _49326_/X _49338_/Y _86407_/D sky130_fd_sc_hd__a21boi_4
X_80451_ _80445_/Y _80451_/B _82256_/D sky130_fd_sc_hd__xor2_4
X_68173_ _68129_/A _68173_/X sky130_fd_sc_hd__buf_2
X_65385_ _65009_/X _86147_/Q _65182_/X _65384_/X _65385_/X sky130_fd_sc_hd__a211o_4
X_62597_ _61666_/A _62597_/B _62501_/X _62597_/D _62600_/B sky130_fd_sc_hd__nand4_4
X_67124_ _87420_/Q _67121_/X _67122_/X _67123_/X _67124_/X sky130_fd_sc_hd__a211o_4
X_52350_ _85840_/Q _52347_/X _52349_/Y _52350_/Y sky130_fd_sc_hd__o21ai_4
X_64336_ _64336_/A _58543_/A _64323_/X _64336_/Y sky130_fd_sc_hd__nand3_4
X_83170_ _83167_/CLK _72972_/X _83170_/Q sky130_fd_sc_hd__dfxtp_4
X_61548_ _61499_/A _61548_/B _61538_/C _61548_/Y sky130_fd_sc_hd__nand3_4
X_80382_ _80383_/B _80372_/X _80382_/X sky130_fd_sc_hd__or2_4
Xclkbuf_7_84_0_CLK clkbuf_7_85_0_CLK/A clkbuf_7_84_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_51301_ _86036_/Q _51285_/X _51300_/Y _51301_/Y sky130_fd_sc_hd__o21ai_4
X_82121_ _82485_/CLK _77792_/X _82109_/D sky130_fd_sc_hd__dfxtp_4
X_67055_ _66560_/X _67055_/X sky130_fd_sc_hd__buf_2
X_52281_ _50578_/A _50578_/B _52280_/X _52281_/X sky130_fd_sc_hd__o21a_4
X_64267_ _64267_/A _64267_/X sky130_fd_sc_hd__buf_2
X_61479_ _61437_/A _61479_/B _61459_/X _61479_/Y sky130_fd_sc_hd__nand3_4
X_54020_ _54020_/A _46433_/A _54020_/Y sky130_fd_sc_hd__nand2_4
X_66006_ _65932_/A _66006_/B _66006_/X sky130_fd_sc_hd__and2_4
X_51232_ _51228_/Y _51229_/X _51231_/X _86050_/D sky130_fd_sc_hd__a21oi_4
X_63218_ _63212_/Y _63214_/X _63215_/X _63217_/X _63183_/X _63218_/Y
+ sky130_fd_sc_hd__o41ai_4
X_82052_ _84074_/CLK _82052_/D _82052_/Q sky130_fd_sc_hd__dfxtp_4
X_64198_ _60034_/X _64490_/A sky130_fd_sc_hd__buf_2
X_81003_ _83238_/CLK _84211_/Q _81003_/Q sky130_fd_sc_hd__dfxtp_4
X_51163_ _86062_/Q _51156_/X _51162_/Y _51163_/Y sky130_fd_sc_hd__o21ai_4
X_63149_ _60508_/A _63149_/X sky130_fd_sc_hd__buf_2
X_86860_ _86861_/CLK _45701_/Y _63227_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_99_0_CLK clkbuf_7_98_0_CLK/A clkbuf_7_99_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_50114_ _50064_/A _50120_/A sky130_fd_sc_hd__buf_2
X_85811_ _86422_/CLK _52493_/Y _64974_/B sky130_fd_sc_hd__dfxtp_4
X_51094_ _51013_/A _51115_/B sky130_fd_sc_hd__buf_2
X_67957_ _67952_/X _67956_/X _67858_/X _67961_/A sky130_fd_sc_hd__a21o_4
X_55971_ _55968_/X _55970_/X _55615_/X _55974_/A sky130_fd_sc_hd__a21o_4
X_86791_ _87077_/CLK _86791_/D _86791_/Q sky130_fd_sc_hd__dfxtp_4
X_57710_ _65034_/A _57965_/A sky130_fd_sc_hd__buf_2
X_50045_ _50929_/A _50045_/X sky130_fd_sc_hd__buf_2
X_54922_ _54932_/A _54910_/B _54932_/C _53230_/D _54922_/X sky130_fd_sc_hd__and4_4
X_85742_ _85745_/CLK _52858_/Y _85742_/Q sky130_fd_sc_hd__dfxtp_4
X_66908_ _87121_/Q _66833_/X _66834_/X _66907_/X _66908_/X sky130_fd_sc_hd__a211o_4
X_58690_ _58605_/X _85943_/Q _58679_/X _58690_/X sky130_fd_sc_hd__o21a_4
X_82954_ _82769_/CLK _82954_/D _82954_/Q sky130_fd_sc_hd__dfxtp_4
X_67888_ _68402_/A _67888_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_22_0_CLK clkbuf_7_23_0_CLK/A clkbuf_8_45_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_57641_ _57638_/Y _57627_/X _57640_/Y _84964_/D sky130_fd_sc_hd__a21boi_4
X_81905_ _81989_/CLK _77453_/X _82281_/D sky130_fd_sc_hd__dfxtp_4
X_69627_ _69865_/A _69627_/B _69627_/X sky130_fd_sc_hd__and2_4
X_54853_ _54851_/Y _54830_/X _54852_/X _54853_/Y sky130_fd_sc_hd__a21oi_4
X_66839_ _87880_/Q _66816_/X _66794_/X _66838_/X _66839_/X sky130_fd_sc_hd__a211o_4
X_85673_ _86400_/CLK _53231_/Y _85673_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_162_0_CLK clkbuf_7_81_0_CLK/X clkbuf_9_325_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_82885_ _82317_/CLK _78101_/B _82885_/Q sky130_fd_sc_hd__dfxtp_4
X_87412_ _88180_/CLK _87412_/D _87412_/Q sky130_fd_sc_hd__dfxtp_4
X_53804_ _85565_/Q _53784_/X _53803_/Y _53804_/Y sky130_fd_sc_hd__o21ai_4
X_84624_ _84624_/CLK _84624_/D _79615_/A sky130_fd_sc_hd__dfxtp_4
X_57572_ _48011_/A _57619_/B _46603_/X _57572_/X sky130_fd_sc_hd__and3_4
X_69558_ _44022_/X _69558_/B _69558_/X sky130_fd_sc_hd__and2_4
X_81836_ _81834_/CLK _81868_/Q _77376_/A sky130_fd_sc_hd__dfxtp_4
X_88392_ _88394_/CLK _40434_/Y _88392_/Q sky130_fd_sc_hd__dfxtp_4
X_54784_ _54892_/A _54784_/X sky130_fd_sc_hd__buf_2
X_51996_ _52185_/A _52027_/A sky130_fd_sc_hd__buf_2
X_59311_ _58904_/A _59311_/X sky130_fd_sc_hd__buf_2
X_56523_ _56523_/A _56533_/B _56523_/C _56523_/Y sky130_fd_sc_hd__nand3_4
X_68509_ _68993_/A _68509_/X sky130_fd_sc_hd__buf_2
X_87343_ _86988_/CLK _43613_/Y _43610_/A sky130_fd_sc_hd__dfxtp_4
X_53735_ _53732_/Y _53715_/X _53734_/X _53735_/Y sky130_fd_sc_hd__a21oi_4
X_84555_ _84555_/CLK _84555_/D _84555_/Q sky130_fd_sc_hd__dfxtp_4
X_50947_ _50973_/A _50963_/A sky130_fd_sc_hd__buf_2
X_81767_ _88175_/CLK _76011_/X _48653_/A sky130_fd_sc_hd__dfxtp_4
X_69489_ _69329_/X _68986_/Y _69405_/X _69488_/Y _69489_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_7_37_0_CLK clkbuf_6_18_0_CLK/X clkbuf_8_75_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_40700_ _40700_/A _40760_/B _40700_/X sky130_fd_sc_hd__or2_4
X_59242_ _59237_/X _59239_/Y _59240_/Y _59169_/X _59241_/X _59242_/X
+ sky130_fd_sc_hd__o32a_4
X_71520_ _53246_/B _71508_/X _71519_/Y _83469_/D sky130_fd_sc_hd__o21ai_4
X_83506_ _83508_/CLK _83506_/D _83506_/Q sky130_fd_sc_hd__dfxtp_4
X_56454_ _56377_/X _56454_/B _56454_/C _56454_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_8_177_0_CLK clkbuf_7_88_0_CLK/X clkbuf_9_355_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_80718_ _81117_/CLK _75904_/X _80718_/Q sky130_fd_sc_hd__dfxtp_4
X_87274_ _87533_/CLK _43769_/X _69262_/B sky130_fd_sc_hd__dfxtp_4
X_53666_ _53733_/A _53666_/X sky130_fd_sc_hd__buf_2
X_41680_ _41659_/X _41330_/A _41679_/X _41680_/Y sky130_fd_sc_hd__o21ai_4
X_84486_ _83231_/CLK _84486_/D _79154_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_172_0_CLK clkbuf_9_86_0_CLK/X _81684_/CLK sky130_fd_sc_hd__clkbuf_1
X_50878_ _50822_/A _51394_/B _50878_/Y sky130_fd_sc_hd__nand2_4
X_81698_ _84020_/CLK _81698_/D _81698_/Q sky130_fd_sc_hd__dfxtp_4
X_55405_ _55405_/A _55405_/X sky130_fd_sc_hd__buf_2
X_86225_ _86222_/CLK _86225_/D _86225_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_201 sky130_fd_sc_hd__decap_3
X_40631_ _40817_/A _82873_/Q _40631_/X sky130_fd_sc_hd__or2_4
X_52617_ _85785_/Q _52601_/X _52616_/Y _52617_/Y sky130_fd_sc_hd__o21ai_4
X_59173_ _86675_/Q _59068_/B _59173_/Y sky130_fd_sc_hd__nor2_4
X_71451_ _71445_/X _83495_/Q _71450_/Y _83495_/D sky130_fd_sc_hd__a21o_4
X_83437_ _83491_/CLK _83437_/D _83437_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_212 sky130_fd_sc_hd__decap_3
X_80649_ _74803_/Y _74713_/Y DATA_FROM_HASH[6] sky130_fd_sc_hd__ebufn_2
X_56385_ _56436_/A _56386_/B sky130_fd_sc_hd__buf_2
X_53597_ _53601_/A _48122_/Y _53597_/Y sky130_fd_sc_hd__nand2_4
XPHY_223 sky130_fd_sc_hd__decap_3
XPHY_234 sky130_fd_sc_hd__decap_3
X_58124_ _58124_/A _58846_/A sky130_fd_sc_hd__buf_2
X_70402_ _70942_/A _74531_/A _70407_/C _70402_/Y sky130_fd_sc_hd__nand3_4
XPHY_245 sky130_fd_sc_hd__decap_3
X_43350_ _43305_/A _43350_/X sky130_fd_sc_hd__buf_2
X_55336_ _55333_/X _55335_/X _55309_/X _55336_/X sky130_fd_sc_hd__a21o_4
X_74170_ _44735_/Y _73491_/X _74169_/Y _74170_/X sky130_fd_sc_hd__a21o_4
X_86156_ _85837_/CLK _50673_/Y _86156_/Q sky130_fd_sc_hd__dfxtp_4
X_40562_ _40350_/A _42447_/B sky130_fd_sc_hd__inv_2
X_52548_ _52546_/Y _52541_/X _52547_/Y _85800_/D sky130_fd_sc_hd__a21boi_4
XPHY_256 sky130_fd_sc_hd__decap_3
X_71382_ _71373_/X _83519_/Q _71381_/Y _71382_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_9_293_0_CLK clkbuf_8_146_0_CLK/X clkbuf_9_293_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_83368_ _83367_/CLK _83368_/D _83368_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_100_0_CLK clkbuf_7_50_0_CLK/X clkbuf_9_201_0_CLK/A sky130_fd_sc_hd__clkbuf_1
XPHY_267 sky130_fd_sc_hd__decap_3
XPHY_278 sky130_fd_sc_hd__decap_3
X_42301_ _41580_/X _42290_/X _87932_/Q _42291_/X _87932_/D sky130_fd_sc_hd__a2bb2o_4
X_73121_ _73121_/A _73120_/X _73121_/X sky130_fd_sc_hd__xor2_4
XPHY_289 sky130_fd_sc_hd__decap_3
X_85107_ _85042_/CLK _85107_/D _85107_/Q sky130_fd_sc_hd__dfxtp_4
X_58055_ _86633_/Q _57954_/X _58055_/Y sky130_fd_sc_hd__nor2_4
X_70333_ _70338_/A _70333_/B _83090_/Q _70332_/X _70333_/X sky130_fd_sc_hd__and4_4
X_82319_ _82327_/CLK _77094_/B _82319_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_187_0_CLK clkbuf_9_93_0_CLK/X _81041_/CLK sky130_fd_sc_hd__clkbuf_1
X_43281_ _43280_/Y _87502_/D sky130_fd_sc_hd__inv_2
X_55267_ _55711_/A _57468_/A _55267_/X sky130_fd_sc_hd__and2_4
X_86087_ _85767_/CLK _51030_/Y _86087_/Q sky130_fd_sc_hd__dfxtp_4
X_40493_ _40477_/X _40488_/X _40491_/X _88383_/Q _40492_/X _40494_/A
+ sky130_fd_sc_hd__o32ai_4
X_52479_ _52477_/Y _52462_/X _52478_/Y _52479_/Y sky130_fd_sc_hd__a21boi_4
X_83299_ _85555_/CLK _83299_/D _83299_/Q sky130_fd_sc_hd__dfxtp_4
X_45020_ _45020_/A _45033_/B _45020_/Y sky130_fd_sc_hd__nand2_4
X_57006_ _85102_/Q _57084_/A _57004_/Y _57005_/Y _85102_/D sky130_fd_sc_hd__a211o_4
X_42232_ _42231_/X _42226_/X _41382_/X _87969_/Q _42228_/X _42232_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54218_ _54208_/X _54237_/B _54209_/C _53052_/D _54218_/X sky130_fd_sc_hd__and4_4
X_85038_ _85037_/CLK _57302_/Y _85038_/Q sky130_fd_sc_hd__dfxtp_4
X_73052_ _72795_/A _73053_/B sky130_fd_sc_hd__buf_2
X_70264_ _70249_/X _70264_/X sky130_fd_sc_hd__buf_2
X_55198_ _55171_/X _55178_/X _55199_/A sky130_fd_sc_hd__and2_4
X_72003_ _72040_/A _48973_/A _72003_/Y sky130_fd_sc_hd__nand2_4
X_42163_ _41199_/X _42161_/X _88003_/Q _42162_/X _88003_/D sky130_fd_sc_hd__a2bb2o_4
X_54149_ _54149_/A _47313_/Y _54149_/Y sky130_fd_sc_hd__nand2_4
X_77860_ _77855_/Y _77860_/B _77875_/A sky130_fd_sc_hd__nand2_4
Xclkbuf_8_115_0_CLK clkbuf_7_57_0_CLK/X clkbuf_9_230_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_70195_ _70209_/A _70195_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_110_0_CLK clkbuf_9_55_0_CLK/X _87183_/CLK sky130_fd_sc_hd__clkbuf_1
X_41114_ _41114_/A _41079_/X _41114_/X sky130_fd_sc_hd__or2_4
X_76811_ _81668_/Q _76811_/B _76811_/Y sky130_fd_sc_hd__xnor2_4
Xclkbuf_10_740_0_CLK clkbuf_9_370_0_CLK/X _87749_/CLK sky130_fd_sc_hd__clkbuf_1
X_46971_ _82396_/Q _46971_/Y sky130_fd_sc_hd__inv_2
X_42094_ _42077_/A _42094_/X sky130_fd_sc_hd__buf_2
X_58957_ _58920_/A _58957_/B _58957_/Y sky130_fd_sc_hd__nor2_4
X_77791_ _77796_/B _77791_/B _77792_/B sky130_fd_sc_hd__xnor2_4
X_86989_ _86989_/CLK _86989_/D _73985_/A sky130_fd_sc_hd__dfxtp_4
X_48710_ _48874_/B _50556_/B sky130_fd_sc_hd__buf_2
X_79530_ _79527_/Y _79529_/Y _79895_/A sky130_fd_sc_hd__nand2_4
X_45922_ _64902_/A _45922_/X sky130_fd_sc_hd__buf_2
X_41045_ _41045_/A _41045_/X sky130_fd_sc_hd__buf_2
X_57908_ _58882_/A _58610_/A sky130_fd_sc_hd__buf_2
X_76742_ _81483_/Q _81355_/D _76741_/X _76742_/Y sky130_fd_sc_hd__o21ai_4
X_49690_ _49699_/A _47184_/X _49690_/Y sky130_fd_sc_hd__nand2_4
X_73954_ _73954_/A _86545_/Q _73954_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_231_0_CLK clkbuf_9_230_0_CLK/A clkbuf_9_231_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_58888_ _58828_/X _58886_/Y _58887_/Y _58874_/X _58832_/X _58888_/X
+ sky130_fd_sc_hd__o32a_4
X_48641_ _86504_/Q _48612_/X _48640_/Y _48641_/Y sky130_fd_sc_hd__o21ai_4
X_72905_ _72905_/A _72905_/X sky130_fd_sc_hd__buf_2
X_79461_ _79449_/A _79448_/Y _79460_/X _79461_/X sky130_fd_sc_hd__a21o_4
X_45853_ _85059_/Q _55221_/B sky130_fd_sc_hd__inv_2
X_57839_ _57739_/X _85722_/Q _57814_/X _57839_/X sky130_fd_sc_hd__o21a_4
X_76673_ _76673_/A _76672_/Y _76673_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_125_0_CLK clkbuf_9_62_0_CLK/X _84393_/CLK sky130_fd_sc_hd__clkbuf_1
X_73885_ _73885_/A _73884_/X _73886_/B sky130_fd_sc_hd__nand2_4
X_78412_ _78412_/A _78412_/Y sky130_fd_sc_hd__inv_2
X_44804_ _41446_/Y _46258_/A _86945_/Q _40354_/X _86945_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_10_755_0_CLK clkbuf_9_377_0_CLK/X _88034_/CLK sky130_fd_sc_hd__clkbuf_1
X_75624_ _75621_/X _75622_/Y _75623_/X _75625_/A sky130_fd_sc_hd__a21oi_4
X_48572_ _48572_/A _48811_/B sky130_fd_sc_hd__buf_2
X_72836_ _72929_/A _72836_/B _72836_/X sky130_fd_sc_hd__and2_4
X_60850_ _60909_/A _60997_/A sky130_fd_sc_hd__buf_2
X_79392_ _58711_/Y _66429_/C _79391_/Y _79392_/X sky130_fd_sc_hd__o21a_4
X_45784_ _45781_/Y _45783_/Y _45757_/X _45784_/X sky130_fd_sc_hd__a21o_4
X_42996_ _40497_/X _42994_/X _87614_/Q _42995_/X _87614_/D sky130_fd_sc_hd__a2bb2o_4
X_47523_ _47518_/Y _47509_/X _47522_/X _86626_/D sky130_fd_sc_hd__a21oi_4
X_59509_ _59508_/X _59509_/X sky130_fd_sc_hd__buf_2
X_78343_ _78342_/Y _78343_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_9_246_0_CLK clkbuf_9_247_0_CLK/A clkbuf_9_246_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_44735_ _86981_/Q _44735_/Y sky130_fd_sc_hd__inv_2
X_75555_ _75555_/A _75555_/Y sky130_fd_sc_hd__inv_2
X_41947_ _88096_/Q _41947_/Y sky130_fd_sc_hd__inv_2
X_60781_ _60781_/A _60780_/X _60781_/Y sky130_fd_sc_hd__nor2_4
X_72767_ _72763_/X _72764_/Y _72766_/X _72767_/Y sky130_fd_sc_hd__a21oi_4
X_62520_ _62520_/A _62561_/B sky130_fd_sc_hd__buf_2
X_74506_ _74504_/Y _74492_/X _74505_/X _74506_/Y sky130_fd_sc_hd__a21oi_4
X_47454_ _81801_/Q _54748_/D sky130_fd_sc_hd__inv_2
X_71718_ _71711_/Y _71718_/X sky130_fd_sc_hd__buf_2
X_78274_ _78274_/A _78284_/B _78274_/Y sky130_fd_sc_hd__nand2_4
X_44666_ _44650_/A _44666_/X sky130_fd_sc_hd__buf_2
X_75486_ _75486_/A _75485_/X _75486_/X sky130_fd_sc_hd__xor2_4
X_41878_ _41878_/A _42547_/A sky130_fd_sc_hd__buf_2
X_72698_ _70241_/C _72686_/X _72697_/Y _83185_/D sky130_fd_sc_hd__a21bo_4
X_46405_ _82932_/Q _46459_/B _46405_/X sky130_fd_sc_hd__or2_4
X_77225_ _77227_/C _77225_/Y sky130_fd_sc_hd__inv_2
X_43617_ _40617_/X _43604_/X _87341_/Q _43607_/X _43617_/X sky130_fd_sc_hd__a2bb2o_4
X_62451_ _62493_/A _62446_/Y _62451_/C _62450_/Y _62451_/Y sky130_fd_sc_hd__nand4_4
X_74437_ _74466_/A _74437_/B _74437_/Y sky130_fd_sc_hd__nand2_4
X_40829_ _40829_/A _40829_/B _40829_/X sky130_fd_sc_hd__or2_4
X_47385_ _47385_/A _47385_/Y sky130_fd_sc_hd__inv_2
X_71649_ _71649_/A _71649_/X sky130_fd_sc_hd__buf_2
X_44597_ _44593_/X _44594_/X _40921_/X _44595_/Y _44596_/X _87042_/D
+ sky130_fd_sc_hd__o32ai_4
X_49124_ _83601_/Q _72077_/B sky130_fd_sc_hd__inv_2
X_61402_ _61377_/A _61399_/X _61429_/C _61402_/Y sky130_fd_sc_hd__nand3_4
X_46336_ _86746_/Q _46279_/X _46335_/Y _46336_/Y sky130_fd_sc_hd__o21ai_4
X_65170_ _65397_/A _65047_/B _65170_/C _65170_/Y sky130_fd_sc_hd__nor3_4
X_77156_ _77157_/A _77157_/B _77156_/Y sky130_fd_sc_hd__nor2_4
X_43548_ _43548_/A _43548_/Y sky130_fd_sc_hd__inv_2
X_62382_ _62342_/A _62341_/X _84414_/Q _62382_/Y sky130_fd_sc_hd__nor3_4
X_74368_ _72068_/A _48367_/Y _74368_/Y sky130_fd_sc_hd__nand2_4
X_64121_ _60879_/B _64179_/C sky130_fd_sc_hd__buf_2
X_76107_ _76107_/A _76107_/Y sky130_fd_sc_hd__inv_2
X_61333_ _61321_/Y _61334_/A sky130_fd_sc_hd__buf_2
X_49055_ _49055_/A _50649_/B sky130_fd_sc_hd__buf_2
X_73319_ _72852_/X _73319_/X sky130_fd_sc_hd__buf_2
X_46267_ _46267_/A _53949_/B sky130_fd_sc_hd__buf_2
X_77087_ _77084_/Y _77087_/B _77097_/A sky130_fd_sc_hd__nand2_4
X_43479_ _43528_/A _43479_/X sky130_fd_sc_hd__buf_2
X_74299_ _74297_/A _74297_/B _55956_/B _74299_/Y sky130_fd_sc_hd__nand3_4
X_48006_ _48759_/A _48734_/A sky130_fd_sc_hd__buf_2
X_45218_ _63238_/B _61568_/B sky130_fd_sc_hd__buf_2
X_64052_ _61560_/B _64052_/B _64150_/C _64052_/D _64052_/Y sky130_fd_sc_hd__nand4_4
X_76038_ _76038_/A _76038_/B _76039_/B sky130_fd_sc_hd__nand2_4
X_61264_ _61264_/A _61264_/B _61264_/Y sky130_fd_sc_hd__nand2_4
X_46198_ _66002_/A _65464_/A sky130_fd_sc_hd__buf_2
X_63003_ _63002_/X _63003_/Y sky130_fd_sc_hd__inv_2
X_60215_ _60192_/Y _60198_/Y _60207_/Y _60300_/B _60214_/Y _84649_/D
+ sky130_fd_sc_hd__a41oi_4
X_45149_ _85265_/Q _45147_/X _45148_/X _45149_/Y sky130_fd_sc_hd__o21ai_4
X_68860_ _74031_/A _68414_/X _68379_/X _68859_/Y _68860_/X sky130_fd_sc_hd__a211o_4
X_61195_ _61195_/A _61196_/A sky130_fd_sc_hd__inv_2
Xclkbuf_10_708_0_CLK clkbuf_9_354_0_CLK/X _87086_/CLK sky130_fd_sc_hd__clkbuf_1
X_67811_ _87455_/Q _67717_/X _67718_/X _67810_/X _67811_/X sky130_fd_sc_hd__a211o_4
X_60146_ _60145_/Y _59230_/X _59968_/B _60005_/Y _60146_/Y sky130_fd_sc_hd__a22oi_4
X_49957_ _49930_/X _49973_/C sky130_fd_sc_hd__buf_2
X_68791_ _88002_/Q _68715_/X _68540_/X _68790_/X _68791_/X sky130_fd_sc_hd__a211o_4
X_77989_ _77950_/A _77965_/A _77957_/A _77980_/C _77989_/X sky130_fd_sc_hd__and4_4
X_48908_ _48908_/A _71970_/B _48908_/X sky130_fd_sc_hd__and2_4
X_67742_ _68442_/A _67742_/X sky130_fd_sc_hd__buf_2
X_79728_ _79725_/Y _79708_/Y _79727_/X _79728_/Y sky130_fd_sc_hd__o21ai_4
X_64954_ _64929_/A _85812_/Q _64954_/X sky130_fd_sc_hd__and2_4
X_60077_ _66064_/A _60359_/A sky130_fd_sc_hd__buf_2
X_49888_ _49861_/A _49893_/B sky130_fd_sc_hd__buf_2
X_63905_ _61891_/X _63876_/B _63905_/C _63892_/D _63905_/Y sky130_fd_sc_hd__nand4_4
X_48839_ _86473_/Q _48836_/X _48838_/Y _48839_/Y sky130_fd_sc_hd__o21ai_4
X_67673_ _86961_/Q _67670_/X _67671_/X _67672_/X _67673_/X sky130_fd_sc_hd__a211o_4
X_79659_ _79657_/X _79668_/B _79659_/Y sky130_fd_sc_hd__xnor2_4
X_64885_ _64882_/X _64884_/X _64729_/X _64885_/X sky130_fd_sc_hd__a21o_4
X_69412_ _87519_/Q _69205_/X _69343_/X _69411_/X _69412_/X sky130_fd_sc_hd__a211o_4
X_66624_ _67816_/A _66625_/A sky130_fd_sc_hd__buf_2
X_51850_ _51823_/A _51850_/X sky130_fd_sc_hd__buf_2
X_63836_ _61406_/A _63772_/B _63803_/C _63787_/D _63836_/Y sky130_fd_sc_hd__nand4_4
X_82670_ _82923_/CLK _82670_/D _82670_/Q sky130_fd_sc_hd__dfxtp_4
X_50801_ _50551_/A _50801_/X sky130_fd_sc_hd__buf_2
X_81621_ _81259_/CLK _76435_/Y _81813_/D sky130_fd_sc_hd__dfxtp_4
X_69343_ _68385_/A _69343_/X sky130_fd_sc_hd__buf_2
X_66555_ _66554_/X _66647_/A sky130_fd_sc_hd__buf_2
X_51781_ _51781_/A _51794_/C sky130_fd_sc_hd__buf_2
X_63767_ _63644_/A _63800_/A sky130_fd_sc_hd__buf_2
X_60979_ _72250_/A _60979_/X sky130_fd_sc_hd__buf_2
X_53520_ _53503_/X _53520_/B _53520_/Y sky130_fd_sc_hd__nand2_4
X_65506_ _65503_/X _85596_/Q _65504_/X _65505_/X _65506_/X sky130_fd_sc_hd__a211o_4
X_84340_ _83216_/CLK _84340_/D _79288_/A sky130_fd_sc_hd__dfxtp_4
X_50732_ _50730_/Y _50676_/X _50731_/Y _86145_/D sky130_fd_sc_hd__a21oi_4
X_62718_ _62669_/A _63069_/A _62704_/C _62717_/X _62718_/X sky130_fd_sc_hd__and4_4
X_81552_ _83918_/CLK _81552_/D _76171_/B sky130_fd_sc_hd__dfxtp_4
X_69274_ _69288_/A _69274_/B _69274_/X sky130_fd_sc_hd__and2_4
X_66486_ _66482_/Y _66483_/X _66485_/Y _84114_/D sky130_fd_sc_hd__a21o_4
X_63698_ _61673_/B _63426_/A _63696_/X _63697_/X _63698_/X sky130_fd_sc_hd__a211o_4
X_80503_ _80496_/X _80498_/B _80503_/Y sky130_fd_sc_hd__nand2_4
X_68225_ _67397_/X _67400_/X _68209_/X _68225_/Y sky130_fd_sc_hd__a21oi_4
X_53451_ _54321_/A _54919_/A sky130_fd_sc_hd__buf_2
X_65437_ _64630_/X _65548_/B _64632_/X _65447_/A sky130_fd_sc_hd__nand3_4
X_84271_ _80728_/CLK _64141_/Y _84271_/Q sky130_fd_sc_hd__dfxtp_4
X_50663_ _86158_/Q _50626_/X _50662_/Y _50663_/Y sky130_fd_sc_hd__o21ai_4
X_62649_ _62886_/A _62949_/B sky130_fd_sc_hd__buf_2
X_81483_ _81482_/CLK _81483_/D _81483_/Q sky130_fd_sc_hd__dfxtp_4
X_86010_ _86008_/CLK _86010_/D _86010_/Q sky130_fd_sc_hd__dfxtp_4
X_52402_ _65313_/B _52397_/X _52401_/Y _52402_/Y sky130_fd_sc_hd__o21ai_4
X_83222_ _83231_/CLK _72599_/Y _79310_/B sky130_fd_sc_hd__dfxtp_4
X_56170_ _56177_/A _56168_/X _56169_/Y _85283_/D sky130_fd_sc_hd__o21ai_4
X_80434_ _80432_/X _80434_/B _80448_/A sky130_fd_sc_hd__xnor2_4
X_68156_ _66987_/X _66990_/X _68129_/X _68156_/Y sky130_fd_sc_hd__a21oi_4
X_53382_ _53355_/A _53382_/X sky130_fd_sc_hd__buf_2
X_65368_ _65342_/X _86724_/Q _65239_/X _65367_/X _65368_/X sky130_fd_sc_hd__a211o_4
X_50594_ _50594_/A _50594_/X sky130_fd_sc_hd__buf_2
X_55121_ _55119_/Y _55102_/X _55120_/X _85314_/D sky130_fd_sc_hd__a21oi_4
X_67107_ _67133_/A _67107_/B _67107_/X sky130_fd_sc_hd__and2_4
X_52333_ _52331_/Y _52314_/X _52332_/X _52333_/Y sky130_fd_sc_hd__a21oi_4
X_64319_ _64377_/A _64319_/X sky130_fd_sc_hd__buf_2
X_83153_ _83153_/CLK _83153_/D _83153_/Q sky130_fd_sc_hd__dfxtp_4
X_80365_ _80338_/Y _80363_/Y _80364_/Y _80366_/B sky130_fd_sc_hd__a21oi_4
X_68087_ _81474_/D _68040_/X _68086_/X _84042_/D sky130_fd_sc_hd__a21bo_4
X_65299_ _72123_/A _86118_/Q _45922_/X _65298_/X _65299_/X sky130_fd_sc_hd__a211o_4
X_82104_ _82104_/CLK _82116_/Q _77161_/A sky130_fd_sc_hd__dfxtp_4
X_55052_ _55043_/X _55030_/X _55070_/C _47691_/A _55052_/X sky130_fd_sc_hd__and4_4
X_67038_ _67034_/X _67037_/X _66964_/X _67038_/X sky130_fd_sc_hd__a21o_4
X_52264_ _52260_/Y _52262_/X _52263_/X _52264_/Y sky130_fd_sc_hd__a21oi_4
X_83084_ _83184_/CLK _83084_/D _70346_/C sky130_fd_sc_hd__dfxtp_4
X_87961_ _87221_/CLK _87961_/D _87961_/Q sky130_fd_sc_hd__dfxtp_4
X_80296_ _80296_/A _80297_/A _80297_/B _80296_/Y sky130_fd_sc_hd__nand3_4
X_54003_ _54001_/Y _53982_/X _54002_/Y _85525_/D sky130_fd_sc_hd__a21boi_4
X_51215_ _51213_/Y _51201_/X _51214_/X _86053_/D sky130_fd_sc_hd__a21oi_4
X_86912_ _87636_/CLK _86912_/D _86912_/Q sky130_fd_sc_hd__dfxtp_4
X_82035_ _82005_/CLK _77888_/B _82035_/Q sky130_fd_sc_hd__dfxtp_4
X_59860_ _59855_/A _59855_/B _80323_/A _59860_/Y sky130_fd_sc_hd__nor3_4
X_52195_ _52191_/Y _52170_/X _52194_/X _85871_/D sky130_fd_sc_hd__a21oi_4
X_87892_ _86914_/CLK _87892_/D _87892_/Q sky130_fd_sc_hd__dfxtp_4
X_58811_ _58730_/X _85934_/Q _58810_/X _58811_/X sky130_fd_sc_hd__o21a_4
X_51146_ _51010_/A _51147_/A sky130_fd_sc_hd__buf_2
X_86843_ _81615_/CLK _86843_/D DATA_AVAILABLE sky130_fd_sc_hd__dfxtp_4
X_59791_ _80484_/A _59787_/X _59789_/Y _59790_/X _59791_/X sky130_fd_sc_hd__a2bb2o_4
X_68989_ _69607_/A _68989_/X sky130_fd_sc_hd__buf_2
X_58742_ _58740_/X _85459_/Q _58741_/X _58742_/Y sky130_fd_sc_hd__o21ai_4
X_51077_ _86078_/Q _51073_/X _51076_/Y _51077_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_1012_0_CLK clkbuf_9_506_0_CLK/X _83564_/CLK sky130_fd_sc_hd__clkbuf_1
X_55954_ _55954_/A _55954_/B _55954_/X sky130_fd_sc_hd__and2_4
X_86774_ _81111_/CLK _46109_/Y _40326_/A sky130_fd_sc_hd__dfxtp_4
X_83986_ _87188_/CLK _83986_/D _83986_/Q sky130_fd_sc_hd__dfxtp_4
X_50028_ _72436_/B _50012_/X _50027_/Y _50028_/Y sky130_fd_sc_hd__o21ai_4
X_54905_ _54910_/A _54910_/B _54910_/C _53211_/D _54905_/X sky130_fd_sc_hd__and4_4
X_85725_ _85725_/CLK _85725_/D _85725_/Q sky130_fd_sc_hd__dfxtp_4
X_70951_ _70939_/A _70954_/C sky130_fd_sc_hd__buf_2
X_58673_ _58631_/X _58671_/Y _58672_/Y _58650_/X _58636_/X _58673_/X
+ sky130_fd_sc_hd__o32a_4
X_82937_ _82933_/CLK _78299_/X _46350_/A sky130_fd_sc_hd__dfxtp_4
X_55885_ _55534_/A _56494_/C _55885_/X sky130_fd_sc_hd__and2_4
X_57624_ _57622_/Y _57581_/X _57623_/Y _57624_/Y sky130_fd_sc_hd__a21boi_4
X_42850_ _42847_/X _42849_/X _41520_/X _66852_/B _42836_/X _42850_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54836_ _54889_/A _54857_/C sky130_fd_sc_hd__buf_2
X_73670_ _73655_/X _73658_/Y _73669_/X _73670_/X sky130_fd_sc_hd__a21o_4
X_85656_ _85431_/CLK _53317_/Y _85656_/Q sky130_fd_sc_hd__dfxtp_4
X_70882_ _70827_/B _71287_/C _70882_/Y sky130_fd_sc_hd__nand2_4
X_82868_ _82343_/CLK _82492_/Q _82868_/Q sky130_fd_sc_hd__dfxtp_4
X_41801_ _40331_/X _41799_/X _66609_/B _41800_/X _88146_/D sky130_fd_sc_hd__a2bb2o_4
X_72621_ _72569_/A _72621_/B _72621_/Y sky130_fd_sc_hd__nand2_4
X_84607_ _84606_/CLK _60520_/Y _79147_/A sky130_fd_sc_hd__dfxtp_4
X_57555_ _46401_/A _57597_/A sky130_fd_sc_hd__buf_2
X_81819_ _83184_/CLK _81819_/D _81819_/Q sky130_fd_sc_hd__dfxtp_4
X_88375_ _87417_/CLK _88375_/D _88375_/Q sky130_fd_sc_hd__dfxtp_4
X_54767_ _54764_/Y _54747_/X _54766_/X _85382_/D sky130_fd_sc_hd__a21oi_4
X_42781_ _42700_/A _42781_/X sky130_fd_sc_hd__buf_2
X_85587_ _86191_/CLK _85587_/D _85587_/Q sky130_fd_sc_hd__dfxtp_4
X_51979_ _51961_/X _47932_/B _51979_/Y sky130_fd_sc_hd__nand2_4
X_82799_ _82425_/CLK _82831_/Q _82799_/Q sky130_fd_sc_hd__dfxtp_4
X_56506_ _56085_/X _56499_/X _56505_/Y _85170_/D sky130_fd_sc_hd__o21ai_4
X_44520_ _87069_/Q _44520_/Y sky130_fd_sc_hd__inv_2
X_75340_ _75340_/A _75339_/Y _75341_/A sky130_fd_sc_hd__and2_4
X_87326_ _87850_/CLK _43653_/Y _87326_/Q sky130_fd_sc_hd__dfxtp_4
X_41732_ _41731_/X _41722_/X _88160_/Q _41723_/X _88160_/D sky130_fd_sc_hd__a2bb2o_4
X_53718_ _53713_/A _48582_/A _53718_/Y sky130_fd_sc_hd__nand2_4
X_84538_ _84538_/CLK _84538_/D _76986_/A sky130_fd_sc_hd__dfxtp_4
X_72552_ _79447_/B _60267_/X _72549_/Y _72551_/X _72552_/X sky130_fd_sc_hd__a2bb2o_4
X_57486_ _72484_/A _72710_/A _46173_/X _57364_/D _56923_/Y _57486_/Y
+ sky130_fd_sc_hd__a41oi_4
X_54698_ _85394_/Q _54676_/X _54697_/Y _54698_/Y sky130_fd_sc_hd__o21ai_4
X_59225_ _57790_/X _59226_/B sky130_fd_sc_hd__buf_2
X_71503_ _71487_/A _83475_/Q _71502_/X _71503_/X sky130_fd_sc_hd__a21o_4
X_44451_ _44451_/A _44451_/Y sky130_fd_sc_hd__inv_2
X_56437_ _56446_/A _56446_/B _85194_/Q _56437_/Y sky130_fd_sc_hd__nand3_4
X_75271_ _75267_/Y _75268_/Y _75270_/Y _75271_/X sky130_fd_sc_hd__or3_4
X_41663_ _41662_/Y _41663_/X sky130_fd_sc_hd__buf_2
X_87257_ _87776_/CLK _87257_/D _69494_/B sky130_fd_sc_hd__dfxtp_4
X_53649_ _48744_/A _53658_/B _53667_/C _53649_/X sky130_fd_sc_hd__and3_4
X_72483_ _83250_/Q _72445_/X _72477_/X _72482_/X _83250_/D sky130_fd_sc_hd__a2bb2oi_4
X_84469_ _84469_/CLK _61578_/Y _61577_/C sky130_fd_sc_hd__dfxtp_4
X_77010_ _77010_/A _77011_/B sky130_fd_sc_hd__inv_2
X_43402_ _41479_/X _43396_/X _87439_/Q _43397_/X _43402_/X sky130_fd_sc_hd__a2bb2o_4
X_74222_ _74202_/A _74221_/Y _74222_/Y sky130_fd_sc_hd__nor2_4
X_86208_ _85599_/CLK _86208_/D _86208_/Q sky130_fd_sc_hd__dfxtp_4
X_40614_ _40614_/A _40614_/Y sky130_fd_sc_hd__inv_2
X_47170_ _47169_/Y _52895_/D sky130_fd_sc_hd__buf_2
X_59156_ _58868_/A _59156_/X sky130_fd_sc_hd__buf_2
X_71434_ _71418_/B _71435_/B sky130_fd_sc_hd__buf_2
X_44382_ _44382_/A _44382_/X sky130_fd_sc_hd__buf_2
X_56368_ _56368_/A _56177_/B _55736_/B _56368_/Y sky130_fd_sc_hd__nand3_4
X_87188_ _87188_/CLK _43942_/X _68071_/B sky130_fd_sc_hd__dfxtp_4
X_41594_ _41604_/A _82311_/Q _41594_/X sky130_fd_sc_hd__or2_4
X_46121_ _46121_/A _46121_/Y sky130_fd_sc_hd__inv_2
X_58107_ _84925_/Q _58095_/X _58099_/X _58106_/X _84925_/D sky130_fd_sc_hd__a2bb2oi_4
X_43333_ _41282_/X _43325_/X _87476_/Q _43326_/X _87476_/D sky130_fd_sc_hd__a2bb2o_4
X_55319_ _85070_/Q _55320_/B sky130_fd_sc_hd__inv_2
X_86139_ _86139_/CLK _86139_/D _86139_/Q sky130_fd_sc_hd__dfxtp_4
X_74153_ _74106_/X _85608_/Q _74107_/X _74152_/X _74153_/X sky130_fd_sc_hd__a211o_4
X_40545_ _40542_/X _40543_/X _88373_/Q _40544_/X _88373_/D sky130_fd_sc_hd__a2bb2o_4
X_59087_ _59085_/X _86074_/Q _59086_/X _59087_/Y sky130_fd_sc_hd__o21ai_4
X_71365_ _71429_/A _71365_/X sky130_fd_sc_hd__buf_2
X_56299_ _56296_/A _56298_/X _85245_/Q _56299_/Y sky130_fd_sc_hd__nand3_4
X_73104_ _73104_/A _73104_/B _73104_/Y sky130_fd_sc_hd__nor2_4
X_46052_ _41524_/Y _46043_/X _86793_/Q _46044_/X _46052_/X sky130_fd_sc_hd__a2bb2o_4
X_58038_ _58070_/A _58038_/B _58038_/Y sky130_fd_sc_hd__nor2_4
X_70316_ _70303_/X _74794_/B _70315_/X _70316_/X sky130_fd_sc_hd__a21o_4
X_43264_ _43180_/A _43264_/X sky130_fd_sc_hd__buf_2
X_74084_ _73449_/X _85611_/Q _73450_/X _74083_/X _74084_/X sky130_fd_sc_hd__a211o_4
X_78961_ _78959_/Y _78960_/Y _78970_/B sky130_fd_sc_hd__xor2_4
X_40476_ _40475_/Y _88386_/D sky130_fd_sc_hd__inv_2
X_71296_ _50310_/B _71290_/X _71295_/Y _83545_/D sky130_fd_sc_hd__o21ai_4
X_45003_ _45000_/Y _45002_/Y _44986_/X _45003_/X sky130_fd_sc_hd__a21o_4
X_42215_ _42215_/A _42215_/Y sky130_fd_sc_hd__inv_2
X_77912_ _77890_/Y _81940_/D sky130_fd_sc_hd__inv_2
X_73035_ _72857_/X _73035_/X sky130_fd_sc_hd__buf_2
X_70247_ _70154_/X _70247_/X sky130_fd_sc_hd__buf_2
X_43195_ _43195_/A _87544_/D sky130_fd_sc_hd__inv_2
X_78892_ _78890_/Y _78892_/B _78900_/A sky130_fd_sc_hd__xor2_4
X_60000_ _60000_/A _59962_/A _60000_/Y sky130_fd_sc_hd__nand2_4
X_49811_ _49807_/A _49830_/B _49795_/X _53023_/D _49811_/X sky130_fd_sc_hd__and4_4
X_42146_ _41151_/X _42137_/X _88012_/Q _42138_/X _42146_/X sky130_fd_sc_hd__a2bb2o_4
X_77843_ _82158_/Q _77843_/B _77843_/X sky130_fd_sc_hd__xor2_4
X_70178_ _70183_/A _70183_/B _70178_/C _70183_/D _70178_/X sky130_fd_sc_hd__and4_4
X_59989_ _80215_/A _59339_/X _59988_/Y _59979_/Y _84678_/D sky130_fd_sc_hd__a2bb2oi_4
Xclkbuf_9_170_0_CLK clkbuf_8_85_0_CLK/X clkbuf_9_170_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_49742_ _49825_/A _49742_/X sky130_fd_sc_hd__buf_2
X_46954_ _46949_/Y _46940_/X _46953_/X _86686_/D sky130_fd_sc_hd__a21oi_4
X_42077_ _42077_/A _42077_/X sky130_fd_sc_hd__buf_2
X_77774_ _82151_/Q _77774_/B _82119_/D sky130_fd_sc_hd__xor2_4
X_74986_ _80766_/Q _74995_/B _74986_/X sky130_fd_sc_hd__xor2_4
X_79513_ _79513_/A _79513_/B _79513_/X sky130_fd_sc_hd__xor2_4
X_45905_ _45893_/B _45883_/B _45904_/X _45905_/X sky130_fd_sc_hd__o21a_4
X_41028_ _41027_/Y _41028_/X sky130_fd_sc_hd__buf_2
X_76725_ _76725_/A _76724_/Y _81450_/D sky130_fd_sc_hd__xor2_4
Xclkbuf_10_694_0_CLK clkbuf_9_347_0_CLK/X _87625_/CLK sky130_fd_sc_hd__clkbuf_1
X_49673_ _49651_/X _49669_/B _49669_/C _52887_/D _49673_/X sky130_fd_sc_hd__and4_4
X_61951_ _61736_/A _61957_/A sky130_fd_sc_hd__buf_2
X_73937_ _73937_/A _74003_/B _73937_/Y sky130_fd_sc_hd__nand2_4
X_46885_ _46881_/Y _46844_/X _46884_/X _86693_/D sky130_fd_sc_hd__a21oi_4
X_48624_ _52218_/A _48624_/B _48657_/C _48624_/X sky130_fd_sc_hd__and3_4
X_60902_ _60881_/B _60543_/B _60902_/Y sky130_fd_sc_hd__nand2_4
X_79444_ _79444_/A _79444_/B _79444_/Y sky130_fd_sc_hd__nand2_4
X_45836_ _46187_/A _45836_/X sky130_fd_sc_hd__buf_2
X_64670_ _64769_/A _64670_/B _64670_/X sky130_fd_sc_hd__and2_4
X_76656_ _76655_/Y _76656_/B _76662_/A sky130_fd_sc_hd__nand2_4
Xclkbuf_9_185_0_CLK clkbuf_8_92_0_CLK/X clkbuf_9_185_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_61882_ _61865_/A _61865_/B _78071_/B _61882_/Y sky130_fd_sc_hd__nor3_4
X_73868_ _70100_/Y _73818_/X _73867_/X _73868_/Y sky130_fd_sc_hd__o21ai_4
X_63621_ _63617_/Y _63618_/Y _63620_/X _58457_/A _63363_/X _63621_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75607_ _75891_/A _75607_/B _75607_/Y sky130_fd_sc_hd__nand2_4
X_60833_ _63487_/A _63426_/A sky130_fd_sc_hd__buf_2
X_72819_ _72813_/X _72819_/B _72820_/B sky130_fd_sc_hd__nand2_4
X_48555_ _48134_/X _48018_/A _48554_/X _48801_/B sky130_fd_sc_hd__o21ai_4
X_79375_ _79374_/X _79375_/Y sky130_fd_sc_hd__inv_2
X_45767_ _45758_/X _45762_/Y _45766_/Y _45767_/Y sky130_fd_sc_hd__a21oi_4
X_76587_ _76541_/B _76559_/A _76587_/X sky130_fd_sc_hd__or2_4
X_42979_ _42970_/X _42971_/X _40452_/X _87621_/Q _42976_/X _42979_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73799_ _72951_/A _73799_/X sky130_fd_sc_hd__buf_2
X_47506_ _47506_/A _53086_/B sky130_fd_sc_hd__buf_2
X_66340_ _64704_/X _84963_/Q _64707_/X _66339_/X _66340_/X sky130_fd_sc_hd__a211o_4
X_78326_ _78325_/X _82755_/D sky130_fd_sc_hd__buf_2
X_44718_ _44718_/A _86989_/D sky130_fd_sc_hd__inv_2
X_63552_ _59421_/A _63541_/B _63514_/C _63541_/D _63552_/Y sky130_fd_sc_hd__nand4_4
X_75538_ _75537_/Y _75538_/B _75546_/A sky130_fd_sc_hd__or2_4
X_48486_ _48471_/X _47955_/A _48485_/Y _48487_/A sky130_fd_sc_hd__o21ai_4
X_60764_ _60707_/X _60692_/X _60820_/B _60714_/Y _60763_/Y _60764_/Y
+ sky130_fd_sc_hd__a41oi_4
X_45698_ _45695_/X _45697_/Y _45561_/X _45698_/Y sky130_fd_sc_hd__a21oi_4
X_62503_ _62533_/A _58487_/A _62491_/C _62506_/C sky130_fd_sc_hd__nand3_4
X_47437_ _47530_/A _47437_/X sky130_fd_sc_hd__buf_2
X_66271_ _66236_/X _85608_/Q _66251_/X _66270_/X _66271_/X sky130_fd_sc_hd__a211o_4
X_78257_ _82682_/Q _78257_/B _78257_/X sky130_fd_sc_hd__xor2_4
X_44649_ _40353_/Y _44650_/A sky130_fd_sc_hd__buf_2
X_63483_ _63481_/Y _63455_/X _63482_/Y _63483_/Y sky130_fd_sc_hd__a21oi_4
X_75469_ _75441_/X _75467_/Y _75468_/Y _75508_/B sky130_fd_sc_hd__a21bo_4
X_60695_ _60652_/X _60724_/A sky130_fd_sc_hd__buf_2
X_68010_ _87383_/Q _67987_/X _67938_/X _68009_/X _68010_/X sky130_fd_sc_hd__a211o_4
X_65222_ _65219_/Y _65195_/X _65221_/Y _84210_/D sky130_fd_sc_hd__a21o_4
X_77208_ _77208_/A _77208_/B _77208_/X sky130_fd_sc_hd__xor2_4
X_62434_ _61510_/X _62492_/B _62420_/C _62404_/X _62435_/D sky130_fd_sc_hd__nand4_4
X_47368_ _81810_/Q _47369_/A sky130_fd_sc_hd__inv_2
Xclkbuf_10_632_0_CLK clkbuf_9_316_0_CLK/X _81197_/CLK sky130_fd_sc_hd__clkbuf_1
X_78188_ _78188_/A _78188_/B _78189_/B sky130_fd_sc_hd__xor2_4
X_49107_ _49106_/Y _50674_/B sky130_fd_sc_hd__buf_2
X_46319_ _46505_/A _48936_/A _46319_/Y sky130_fd_sc_hd__nand2_4
X_65153_ _65099_/X _86732_/Q _65028_/X _65152_/X _65153_/X sky130_fd_sc_hd__a211o_4
X_77139_ _82101_/Q _77139_/B _82350_/D sky130_fd_sc_hd__xor2_4
X_62365_ _62337_/A _61891_/X _62364_/X _62280_/D _62365_/X sky130_fd_sc_hd__and4_4
X_47299_ _47287_/X _52969_/B _47299_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_123_0_CLK clkbuf_8_61_0_CLK/X clkbuf_9_123_0_CLK/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_9_50_0_CLK clkbuf_9_51_0_CLK/A clkbuf_9_50_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_64104_ _62544_/Y _60880_/X _62081_/B _61028_/X _64104_/Y sky130_fd_sc_hd__a2bb2oi_4
X_49038_ _48985_/A _49038_/X sky130_fd_sc_hd__buf_2
X_61316_ _61316_/A _61317_/A sky130_fd_sc_hd__buf_2
X_80150_ _84943_/Q _84191_/Q _80150_/Y sky130_fd_sc_hd__nand2_4
X_65084_ _65012_/A _65084_/B _65084_/X sky130_fd_sc_hd__and2_4
X_69961_ _44022_/X _69961_/B _69961_/X sky130_fd_sc_hd__and2_4
X_62296_ _59896_/X _62309_/B sky130_fd_sc_hd__buf_2
X_68912_ _68909_/X _68911_/X _68470_/X _68912_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_10_647_0_CLK clkbuf_9_323_0_CLK/X _88171_/CLK sky130_fd_sc_hd__clkbuf_1
X_64035_ _64053_/A _58442_/A _64071_/C _64035_/X sky130_fd_sc_hd__and3_4
X_61247_ _63001_/A _63053_/A sky130_fd_sc_hd__buf_2
X_80081_ _84937_/Q _65682_/A _80081_/X sky130_fd_sc_hd__xor2_4
X_69892_ _69832_/X _69890_/Y _69870_/X _69891_/Y _69892_/X sky130_fd_sc_hd__a211o_4
X_51000_ _50973_/A _51018_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_138_0_CLK clkbuf_8_69_0_CLK/X clkbuf_9_138_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_68843_ _68840_/X _68842_/X _68470_/X _68843_/X sky130_fd_sc_hd__a21o_4
X_61178_ _59536_/A _59508_/X _61285_/C _61178_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_9_65_0_CLK clkbuf_9_65_0_CLK/A clkbuf_9_65_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_60129_ _60000_/A _60129_/B _60129_/Y sky130_fd_sc_hd__nand2_4
X_83840_ _83835_/CLK _70199_/X _74799_/C sky130_fd_sc_hd__dfxtp_4
X_68774_ _68769_/X _68772_/X _68773_/X _68774_/X sky130_fd_sc_hd__a21o_4
X_65986_ _65700_/X _65983_/Y _65985_/Y _65986_/Y sky130_fd_sc_hd__o21ai_4
X_67725_ _87151_/Q _67670_/X _67671_/X _67724_/X _67725_/X sky130_fd_sc_hd__a211o_4
X_52951_ _85724_/Q _52929_/X _52950_/Y _52951_/Y sky130_fd_sc_hd__o21ai_4
X_64937_ _64933_/X _64937_/B _64936_/X _64937_/Y sky130_fd_sc_hd__nand3_4
X_83771_ _86578_/CLK _83771_/D _83771_/Q sky130_fd_sc_hd__dfxtp_4
X_80983_ _83944_/CLK _75767_/X _80983_/Q sky130_fd_sc_hd__dfxtp_4
X_85510_ _86118_/CLK _85510_/D _85510_/Q sky130_fd_sc_hd__dfxtp_4
X_51902_ _51902_/A _51037_/B _51902_/Y sky130_fd_sc_hd__nand2_4
X_82722_ _82715_/CLK _66524_/C _82722_/Q sky130_fd_sc_hd__dfxtp_4
X_55670_ _83320_/Q _55670_/B _55676_/C sky130_fd_sc_hd__xor2_4
X_67656_ _67653_/X _67655_/X _67561_/X _67656_/X sky130_fd_sc_hd__a21o_4
X_86490_ _86490_/CLK _48749_/Y _72960_/B sky130_fd_sc_hd__dfxtp_4
X_52882_ _85737_/Q _52874_/X _52881_/Y _52882_/Y sky130_fd_sc_hd__o21ai_4
X_64868_ _60151_/X _64855_/Y _64867_/Y _64868_/Y sky130_fd_sc_hd__o21ai_4
X_54621_ _54540_/A _54621_/X sky130_fd_sc_hd__buf_2
X_66607_ _66599_/X _66603_/X _66606_/X _66607_/X sky130_fd_sc_hd__a21o_4
X_85441_ _85761_/CLK _85441_/D _85441_/Q sky130_fd_sc_hd__dfxtp_4
X_51833_ _51851_/A _51815_/B _51810_/C _52661_/D _51833_/X sky130_fd_sc_hd__and4_4
X_63819_ _61390_/A _63772_/B _63803_/C _63787_/D _63819_/Y sky130_fd_sc_hd__nand4_4
X_82653_ _81746_/CLK _82653_/D _82653_/Q sky130_fd_sc_hd__dfxtp_4
X_67587_ _86965_/Q _67585_/X _67516_/X _67586_/X _67587_/X sky130_fd_sc_hd__a211o_4
X_64799_ _64797_/X _86746_/Q _64772_/X _64798_/X _64800_/B sky130_fd_sc_hd__a211o_4
X_57340_ _57026_/X _57340_/B _57340_/C _57340_/Y sky130_fd_sc_hd__nor3_4
X_81604_ _81668_/CLK _76183_/Y _81796_/D sky130_fd_sc_hd__dfxtp_4
X_69326_ _68706_/X _68709_/X _69295_/X _69326_/Y sky130_fd_sc_hd__a21oi_4
X_88160_ _88158_/CLK _88160_/D _88160_/Q sky130_fd_sc_hd__dfxtp_4
X_54552_ _85421_/Q _54540_/X _54551_/Y _54552_/Y sky130_fd_sc_hd__o21ai_4
X_66538_ _66642_/A _66538_/X sky130_fd_sc_hd__buf_2
X_85372_ _85372_/CLK _85372_/D _85372_/Q sky130_fd_sc_hd__dfxtp_4
X_51764_ _51790_/A _51779_/A sky130_fd_sc_hd__buf_2
X_82584_ _82589_/CLK _82616_/Q _78253_/B sky130_fd_sc_hd__dfxtp_4
X_87111_ _87110_/CLK _87111_/D _87111_/Q sky130_fd_sc_hd__dfxtp_4
X_53503_ _53821_/B _53503_/X sky130_fd_sc_hd__buf_2
X_84323_ _84321_/CLK _84323_/D _80559_/B sky130_fd_sc_hd__dfxtp_4
X_50715_ _50713_/Y _50699_/X _50714_/Y _86148_/D sky130_fd_sc_hd__a21boi_4
X_57271_ _57271_/A _83329_/Q _57270_/X _57271_/Y sky130_fd_sc_hd__nand3_4
X_81535_ _81475_/CLK _76595_/B _76136_/A sky130_fd_sc_hd__dfxtp_4
X_69257_ _69216_/X _69255_/Y _69231_/X _69256_/Y _69257_/X sky130_fd_sc_hd__a211o_4
X_88091_ _88087_/CLK _88091_/D _74121_/A sky130_fd_sc_hd__dfxtp_4
X_54483_ _54483_/A _54471_/B _54483_/C _46990_/A _54483_/X sky130_fd_sc_hd__and4_4
X_66469_ _66501_/A _66419_/X _66469_/C _66469_/X sky130_fd_sc_hd__and3_4
X_51695_ _51695_/A _51715_/B _51695_/C _53217_/D _51695_/X sky130_fd_sc_hd__and4_4
X_59010_ _58810_/A _59010_/X sky130_fd_sc_hd__buf_2
X_56222_ _56064_/X _56210_/X _56221_/Y _85270_/D sky130_fd_sc_hd__o21ai_4
X_68208_ _69654_/A _68208_/X sky130_fd_sc_hd__buf_2
X_87042_ _87851_/CLK _87042_/D _87042_/Q sky130_fd_sc_hd__dfxtp_4
X_53434_ _53434_/A _47212_/Y _53434_/Y sky130_fd_sc_hd__nand2_4
X_84254_ _83766_/CLK _64350_/X _79764_/B sky130_fd_sc_hd__dfxtp_4
X_50646_ _50645_/X _53863_/A sky130_fd_sc_hd__buf_2
X_81466_ _82648_/CLK _81466_/D _81466_/Q sky130_fd_sc_hd__dfxtp_4
X_69188_ _69146_/X _69186_/Y _69095_/X _69187_/Y _69188_/X sky130_fd_sc_hd__a211o_4
X_83205_ _83843_/CLK _83205_/D _70183_/C sky130_fd_sc_hd__dfxtp_4
X_56153_ _56152_/Y _56153_/X sky130_fd_sc_hd__buf_2
X_80417_ _80409_/A _80408_/Y _80416_/X _80418_/B sky130_fd_sc_hd__o21ai_4
X_68139_ _82069_/D _68120_/X _68138_/X _84029_/D sky130_fd_sc_hd__a21bo_4
X_53365_ _85647_/Q _53351_/X _53364_/Y _53365_/Y sky130_fd_sc_hd__o21ai_4
X_84185_ _83508_/CLK _84185_/D _65682_/A sky130_fd_sc_hd__dfxtp_4
X_50577_ _50577_/A _50577_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_18_0_CLK clkbuf_8_9_0_CLK/X clkbuf_9_18_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_81397_ _83933_/CLK _83933_/Q _81397_/Q sky130_fd_sc_hd__dfxtp_4
X_55104_ _55112_/A _55104_/B _55120_/C _47784_/A _55104_/X sky130_fd_sc_hd__and4_4
X_52316_ _52313_/Y _52314_/X _52315_/X _52316_/Y sky130_fd_sc_hd__a21oi_4
X_40330_ _40325_/X _82336_/Q _40329_/X _40330_/Y sky130_fd_sc_hd__o21ai_4
X_71150_ _71175_/A _71155_/B _71152_/C _71160_/D _71150_/Y sky130_fd_sc_hd__nand4_4
X_83136_ _83139_/CLK _73794_/Y _83136_/Q sky130_fd_sc_hd__dfxtp_4
X_80348_ _80344_/X _80360_/B _80349_/B sky130_fd_sc_hd__nand2_4
X_56084_ _55854_/X _56083_/X _56084_/Y sky130_fd_sc_hd__xnor2_4
X_53296_ _50063_/A _53352_/A sky130_fd_sc_hd__buf_2
X_70101_ _83132_/Q _70101_/Y sky130_fd_sc_hd__inv_2
X_55035_ _55017_/X _55030_/X _55026_/C _47663_/A _55035_/X sky130_fd_sc_hd__and4_4
X_59912_ _62501_/A _59913_/A sky130_fd_sc_hd__buf_2
X_52247_ _52247_/A _52267_/C sky130_fd_sc_hd__buf_2
X_71081_ _48992_/X _71070_/X _71080_/Y _71081_/Y sky130_fd_sc_hd__o21ai_4
X_83067_ _86500_/CLK _74436_/Y _83067_/Q sky130_fd_sc_hd__dfxtp_4
X_87944_ _87636_/CLK _87944_/D _87944_/Q sky130_fd_sc_hd__dfxtp_4
X_80279_ _80278_/Y _80279_/B _80280_/C sky130_fd_sc_hd__nand2_4
Xclkbuf_9_6_0_CLK clkbuf_9_7_0_CLK/A clkbuf_9_6_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_42000_ _42000_/A _42000_/X sky130_fd_sc_hd__buf_2
X_70032_ _83868_/Q _70029_/X _70031_/X _70032_/X sky130_fd_sc_hd__a21bo_4
X_82018_ _82104_/CLK _77728_/B _81986_/D sky130_fd_sc_hd__dfxtp_4
X_59843_ _59855_/A _59848_/B _80379_/A _59843_/Y sky130_fd_sc_hd__nor3_4
X_52178_ _52214_/A _52178_/X sky130_fd_sc_hd__buf_2
X_87875_ _88387_/CLK _42416_/X _87875_/Q sky130_fd_sc_hd__dfxtp_4
X_51129_ _51129_/A _51130_/A sky130_fd_sc_hd__buf_2
X_74840_ _74839_/Y _80654_/D sky130_fd_sc_hd__inv_2
X_86826_ _87073_/CLK _45989_/Y _86826_/Q sky130_fd_sc_hd__dfxtp_4
X_59774_ _59773_/X _59774_/Y sky130_fd_sc_hd__inv_2
X_56986_ _56985_/X _56702_/X _56986_/X sky130_fd_sc_hd__xor2_4
X_58725_ _58599_/A _58725_/X sky130_fd_sc_hd__buf_2
X_43951_ _43979_/A _43951_/B _43951_/Y sky130_fd_sc_hd__nor2_4
X_55937_ _55937_/A _55956_/B sky130_fd_sc_hd__buf_2
X_74771_ _74771_/A _74804_/A _74797_/C _71738_/X _74771_/Y sky130_fd_sc_hd__nand4_4
X_86757_ _86757_/CLK _46229_/Y _86757_/Q sky130_fd_sc_hd__dfxtp_4
X_71983_ _48938_/A _71959_/X _71964_/X _71983_/X sky130_fd_sc_hd__and3_4
X_83969_ _80931_/CLK _68585_/X _80825_/D sky130_fd_sc_hd__dfxtp_4
X_76510_ _76510_/A _76510_/B _76510_/C _76511_/B sky130_fd_sc_hd__nand3_4
X_42902_ _41663_/X _42900_/X _87661_/Q _42901_/X _42902_/X sky130_fd_sc_hd__a2bb2o_4
X_73722_ _70107_/A _73697_/X _73721_/X _73722_/Y sky130_fd_sc_hd__o21ai_4
X_85708_ _82390_/CLK _53045_/Y _85708_/Q sky130_fd_sc_hd__dfxtp_4
X_58656_ _58125_/X _85786_/Q _58126_/X _58656_/X sky130_fd_sc_hd__o21a_4
X_46670_ _46670_/A _46682_/B _46682_/C _51777_/D _46670_/X sky130_fd_sc_hd__and4_4
X_70934_ _71093_/C _71115_/B sky130_fd_sc_hd__buf_2
X_77490_ _77486_/Y _77487_/Y _77489_/Y _77495_/A sky130_fd_sc_hd__or3_4
X_43882_ _41288_/X _43879_/X _87219_/Q _43880_/X _87219_/D sky130_fd_sc_hd__a2bb2o_4
X_55868_ _85204_/Q _55511_/X _55513_/X _55867_/X _55868_/X sky130_fd_sc_hd__a211o_4
X_86688_ _86688_/CLK _46935_/Y _86688_/Q sky130_fd_sc_hd__dfxtp_4
X_45621_ _82995_/Q _45401_/X _45620_/X _45621_/Y sky130_fd_sc_hd__o21ai_4
X_57607_ _46259_/A _71993_/A sky130_fd_sc_hd__buf_2
X_76441_ _76437_/X _76440_/X _76441_/X sky130_fd_sc_hd__xor2_4
X_42833_ _41479_/X _42830_/X _87695_/Q _42832_/X _42833_/X sky130_fd_sc_hd__a2bb2o_4
X_54819_ _85372_/Q _54812_/X _54818_/Y _54819_/Y sky130_fd_sc_hd__o21ai_4
X_85639_ _85735_/CLK _53411_/Y _85639_/Q sky130_fd_sc_hd__dfxtp_4
X_73653_ _73653_/A _73599_/B _73653_/Y sky130_fd_sc_hd__nor2_4
X_70865_ _71072_/A _70869_/B sky130_fd_sc_hd__buf_2
X_58587_ _58687_/A _58587_/B _58587_/Y sky130_fd_sc_hd__nor2_4
X_55799_ _55796_/X _55798_/X _55800_/A sky130_fd_sc_hd__and2_4
X_48340_ _48401_/A _50378_/B _48340_/Y sky130_fd_sc_hd__nand2_4
X_72604_ _72581_/A _72604_/B _79279_/B _72604_/Y sky130_fd_sc_hd__nor3_4
X_79160_ _79159_/Y _79160_/B _79160_/Y sky130_fd_sc_hd__nand2_4
X_45552_ _44932_/A _45617_/B sky130_fd_sc_hd__buf_2
X_57538_ _84983_/Q _57527_/X _57537_/Y _57538_/Y sky130_fd_sc_hd__o21ai_4
X_76372_ _76364_/X _76371_/X _76381_/A sky130_fd_sc_hd__xnor2_4
X_42764_ _41288_/X _42757_/X _67333_/B _42759_/X _87731_/D sky130_fd_sc_hd__a2bb2o_4
X_88358_ _87859_/CLK _40663_/Y _68699_/B sky130_fd_sc_hd__dfxtp_4
X_73584_ _73378_/X _86240_/Q _73446_/X _73583_/X _73584_/X sky130_fd_sc_hd__a211o_4
X_70796_ _70905_/A _70791_/B _70794_/X _70841_/D _70796_/Y sky130_fd_sc_hd__nand4_4
X_78111_ _78130_/B _78110_/Y _78112_/B sky130_fd_sc_hd__xnor2_4
X_44503_ _44603_/A _44503_/X sky130_fd_sc_hd__buf_2
X_75323_ _75318_/X _75321_/Y _75322_/A _75323_/X sky130_fd_sc_hd__o21a_4
X_87309_ _83158_/CLK _87309_/D _72924_/A sky130_fd_sc_hd__dfxtp_4
X_41715_ _41715_/A _41715_/X sky130_fd_sc_hd__buf_2
X_48271_ _48244_/A _48016_/B _48271_/Y sky130_fd_sc_hd__nand2_4
X_72535_ _72535_/A _72535_/B _72535_/Y sky130_fd_sc_hd__nand2_4
X_79091_ _79074_/A _79089_/A _82654_/Q _79090_/Y _79091_/X sky130_fd_sc_hd__a2bb2o_4
X_45483_ _45434_/X _61390_/A _45452_/X _45483_/Y sky130_fd_sc_hd__o21ai_4
X_57469_ _44292_/A _57346_/C _57468_/X _57469_/X sky130_fd_sc_hd__o21a_4
X_88289_ _87026_/CLK _41039_/Y _88289_/Q sky130_fd_sc_hd__dfxtp_4
X_42695_ _42651_/X _42695_/X sky130_fd_sc_hd__buf_2
X_47222_ _47196_/A _52924_/B _47222_/Y sky130_fd_sc_hd__nand2_4
X_59208_ _59085_/A _59208_/X sky130_fd_sc_hd__buf_2
X_78042_ _77954_/B _78042_/Y sky130_fd_sc_hd__inv_2
X_44434_ _41586_/X _44431_/X _87111_/Q _44432_/X _87111_/D sky130_fd_sc_hd__a2bb2o_4
X_75254_ _75254_/A _75254_/Y sky130_fd_sc_hd__inv_2
X_41646_ _41588_/X _81758_/Q _41645_/X _41646_/Y sky130_fd_sc_hd__o21ai_4
X_60480_ _60479_/Y _60481_/A sky130_fd_sc_hd__buf_2
X_72466_ _57712_/X _85315_/Q _57736_/A _72466_/X sky130_fd_sc_hd__o21a_4
X_74205_ _69053_/B _44128_/X _73031_/X _74204_/Y _74205_/X sky130_fd_sc_hd__a211o_4
X_47153_ _82377_/Q _54576_/D sky130_fd_sc_hd__inv_2
X_59139_ _59061_/X _86070_/Q _59138_/X _59139_/Y sky130_fd_sc_hd__o21ai_4
X_71417_ _71396_/Y _83506_/Q _71416_/Y _83506_/D sky130_fd_sc_hd__a21o_4
X_44365_ _40509_/X _44365_/X sky130_fd_sc_hd__buf_2
X_75185_ _75186_/B _75186_/A _75190_/A sky130_fd_sc_hd__or2_4
X_41577_ _41061_/A _41577_/X sky130_fd_sc_hd__buf_2
X_72397_ _72361_/X _85674_/Q _72362_/X _72397_/X sky130_fd_sc_hd__o21a_4
X_46104_ _74846_/B _46104_/Y sky130_fd_sc_hd__inv_2
X_43316_ _43296_/A _43316_/X sky130_fd_sc_hd__buf_2
X_74136_ _74126_/Y _74136_/B _74136_/Y sky130_fd_sc_hd__xnor2_4
X_62150_ _61663_/B _62161_/B _62187_/C _61706_/X _62150_/Y sky130_fd_sc_hd__nand4_4
X_40528_ _40527_/Y _40528_/X sky130_fd_sc_hd__buf_2
X_47084_ _47084_/A _52846_/D sky130_fd_sc_hd__buf_2
X_71348_ _70591_/A _71349_/D sky130_fd_sc_hd__buf_2
X_44296_ _44147_/A _68714_/A sky130_fd_sc_hd__buf_2
X_79993_ _79989_/Y _79992_/Y _79993_/X sky130_fd_sc_hd__xor2_4
X_61101_ _61101_/A _64323_/A sky130_fd_sc_hd__buf_2
X_46035_ _41478_/Y _46029_/X _86802_/Q _46030_/X _46035_/X sky130_fd_sc_hd__a2bb2o_4
X_43247_ _43180_/A _43247_/X sky130_fd_sc_hd__buf_2
X_62081_ _62055_/A _62081_/B _61755_/X _61728_/A _62081_/X sky130_fd_sc_hd__and4_4
X_74067_ _74055_/X _74057_/Y _74066_/X _74067_/X sky130_fd_sc_hd__a21o_4
X_78944_ _78937_/A _78937_/B _78938_/A _78944_/Y sky130_fd_sc_hd__a21boi_4
X_40459_ _40458_/X _40459_/X sky130_fd_sc_hd__buf_2
X_71279_ _71178_/A _71276_/B _71279_/C _71276_/D _71279_/Y sky130_fd_sc_hd__nand4_4
X_61032_ _60954_/X _60994_/B _59789_/A _60988_/Y _61032_/X sky130_fd_sc_hd__a211o_4
X_73018_ _73018_/A _73018_/B _73019_/B sky130_fd_sc_hd__nand2_4
X_43178_ _43177_/Y _43178_/X sky130_fd_sc_hd__buf_2
X_78875_ _78873_/Y _78875_/B _78875_/Y sky130_fd_sc_hd__nand2_4
X_42129_ _41104_/X _42125_/X _88021_/Q _42126_/X _42129_/X sky130_fd_sc_hd__a2bb2o_4
X_65840_ _44150_/X _83054_/Q _64980_/X _65839_/X _65840_/X sky130_fd_sc_hd__a211o_4
X_77826_ _82269_/Q _81981_/Q _77826_/Y sky130_fd_sc_hd__xnor2_4
X_47986_ _83770_/Q _53531_/B sky130_fd_sc_hd__inv_2
X_49725_ _49722_/Y _49706_/X _49724_/X _86335_/D sky130_fd_sc_hd__a21oi_4
X_46937_ _54451_/B _52760_/B sky130_fd_sc_hd__buf_2
X_65771_ _65767_/X _65741_/B _65770_/X _65772_/B sky130_fd_sc_hd__nand3_4
X_77757_ _77764_/B _77756_/Y _77757_/X sky130_fd_sc_hd__xor2_4
X_62983_ _62847_/A _63344_/A _62939_/X _62975_/D _62983_/X sky130_fd_sc_hd__and4_4
X_74969_ _74969_/A _74969_/B _74969_/X sky130_fd_sc_hd__xor2_4
X_67510_ _87980_/Q _67414_/X _67508_/X _67509_/X _67510_/X sky130_fd_sc_hd__a211o_4
X_64722_ _64828_/A _64722_/X sky130_fd_sc_hd__buf_2
X_76708_ _76708_/A _76707_/X _76712_/A sky130_fd_sc_hd__xnor2_4
X_61934_ _61856_/A _61952_/D sky130_fd_sc_hd__buf_2
X_49656_ _49520_/A _49657_/A sky130_fd_sc_hd__buf_2
X_68490_ _68490_/A _68491_/B sky130_fd_sc_hd__inv_2
X_46868_ _46868_/A _46845_/X _46868_/C _52720_/D _46868_/X sky130_fd_sc_hd__and4_4
X_77688_ _77688_/A _77688_/B _77688_/Y sky130_fd_sc_hd__nand2_4
X_48607_ _48642_/A _48065_/A _48607_/Y sky130_fd_sc_hd__nand2_4
X_67441_ _87471_/Q _67394_/X _67344_/X _67440_/X _67441_/X sky130_fd_sc_hd__a211o_4
X_79427_ _79427_/A _79427_/B _79433_/B sky130_fd_sc_hd__xor2_4
X_45819_ _45819_/A _45819_/X sky130_fd_sc_hd__buf_2
X_64653_ _64680_/A _86271_/Q _64653_/X sky130_fd_sc_hd__and2_4
X_76639_ _76639_/A _76638_/Y _76639_/Y sky130_fd_sc_hd__nand2_4
X_49587_ _49614_/A _49592_/B sky130_fd_sc_hd__buf_2
X_61865_ _61865_/A _61865_/B _78072_/B _61865_/Y sky130_fd_sc_hd__nor3_4
X_46799_ _46845_/A _46830_/B sky130_fd_sc_hd__buf_2
X_63604_ _63615_/A _63615_/B _80422_/B _63604_/Y sky130_fd_sc_hd__nor3_4
X_48538_ _48538_/A _48538_/Y sky130_fd_sc_hd__inv_2
X_60816_ _60558_/X _60826_/A sky130_fd_sc_hd__buf_2
X_67372_ _67369_/X _67371_/X _67322_/X _67372_/X sky130_fd_sc_hd__a21o_4
X_79358_ _79355_/Y _79339_/B _79357_/X _79358_/Y sky130_fd_sc_hd__o21ai_4
X_64584_ _44020_/A _64584_/X sky130_fd_sc_hd__buf_2
X_61796_ _59463_/A _61796_/X sky130_fd_sc_hd__buf_2
X_69111_ _68669_/A _69110_/Y _69111_/Y sky130_fd_sc_hd__nor2_4
X_66323_ _64923_/A _74234_/B _66323_/X sky130_fd_sc_hd__and2_4
X_78309_ _78309_/A _78309_/B _78309_/C _78309_/Y sky130_fd_sc_hd__nand3_4
X_63535_ _63523_/A _61954_/X _63535_/X sky130_fd_sc_hd__and2_4
X_48469_ _48469_/A _48763_/B _48469_/Y sky130_fd_sc_hd__nand2_4
X_60747_ _61075_/C _60694_/Y _60031_/X _60629_/Y _60746_/Y _60747_/Y
+ sky130_fd_sc_hd__a41oi_4
X_79289_ _79287_/X _79288_/X _79304_/B sky130_fd_sc_hd__xnor2_4
Xclkbuf_10_571_0_CLK clkbuf_9_285_0_CLK/X _87110_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_62_0_CLK clkbuf_6_63_0_CLK/A clkbuf_6_62_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_50500_ _50500_/A _50575_/A sky130_fd_sc_hd__buf_2
X_81320_ _81346_/CLK _81320_/D _81728_/D sky130_fd_sc_hd__dfxtp_4
X_69042_ _69021_/A _69042_/B _69042_/X sky130_fd_sc_hd__and2_4
X_66254_ _66250_/X _66253_/X _66240_/X _66254_/X sky130_fd_sc_hd__a21o_4
X_51480_ _51476_/Y _51477_/X _51479_/X _86003_/D sky130_fd_sc_hd__a21oi_4
X_63466_ _63434_/X _63459_/X _63460_/X _63464_/X _63465_/Y _63466_/Y
+ sky130_fd_sc_hd__o41ai_4
X_60678_ _63478_/A _63416_/A sky130_fd_sc_hd__buf_2
X_65205_ _65202_/X _65204_/X _65122_/X _65208_/A sky130_fd_sc_hd__a21o_4
X_50431_ _50428_/Y _50429_/X _50430_/X _86202_/D sky130_fd_sc_hd__a21oi_4
X_62417_ _62236_/A _62472_/B sky130_fd_sc_hd__buf_2
X_81251_ _81794_/CLK _81283_/Q _76159_/A sky130_fd_sc_hd__dfxtp_4
X_66185_ _66182_/X _66184_/X _66057_/X _66185_/X sky130_fd_sc_hd__a21o_4
X_63397_ _58415_/A _63370_/X _61367_/A _63372_/X _63397_/X sky130_fd_sc_hd__a2bb2o_4
X_80202_ _80197_/Y _80201_/Y _80202_/X sky130_fd_sc_hd__xor2_4
X_53150_ _53097_/X _53159_/B sky130_fd_sc_hd__buf_2
X_65136_ _65782_/A _65164_/A sky130_fd_sc_hd__buf_2
X_50362_ _50655_/A _50594_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_586_0_CLK clkbuf_9_293_0_CLK/X _80746_/CLK sky130_fd_sc_hd__clkbuf_1
X_62348_ _61440_/A _62247_/X _62259_/X _62631_/D _62351_/B sky130_fd_sc_hd__nand4_4
X_81182_ _81182_/CLK _75053_/X _81182_/Q sky130_fd_sc_hd__dfxtp_4
X_52101_ _65439_/B _52089_/X _52100_/Y _52101_/Y sky130_fd_sc_hd__o21ai_4
X_80133_ _60051_/C _80133_/B _80141_/B sky130_fd_sc_hd__xor2_4
X_53081_ _85700_/Q _53065_/X _53080_/Y _53081_/Y sky130_fd_sc_hd__o21ai_4
X_65067_ _65065_/X _83296_/Q _64991_/X _65066_/X _65067_/X sky130_fd_sc_hd__a211o_4
X_69944_ _69906_/A _73487_/A _69944_/X sky130_fd_sc_hd__and2_4
X_50293_ _50285_/A _50293_/B _50293_/Y sky130_fd_sc_hd__nand2_4
X_62279_ _62475_/A _62280_/D sky130_fd_sc_hd__buf_2
X_85990_ _85990_/CLK _85990_/D _85990_/Q sky130_fd_sc_hd__dfxtp_4
X_52032_ _85902_/Q _52013_/X _52031_/Y _52032_/Y sky130_fd_sc_hd__o21ai_4
X_64018_ _61997_/X _63955_/X _64050_/C _64033_/D _64018_/Y sky130_fd_sc_hd__nand4_4
X_84941_ _86322_/CLK _84941_/D _84941_/Q sky130_fd_sc_hd__dfxtp_4
X_80064_ _80056_/B _80073_/B _80063_/X _80064_/Y sky130_fd_sc_hd__a21boi_4
X_69875_ _73341_/A _68467_/X _68385_/X _69874_/Y _69875_/X sky130_fd_sc_hd__a211o_4
X_56840_ _56764_/B _56829_/X _56830_/Y _56839_/Y _56841_/A sky130_fd_sc_hd__a211o_4
X_68826_ _69735_/A _68826_/B _68826_/Y sky130_fd_sc_hd__nor2_4
X_87660_ _86935_/CLK _87660_/D _87660_/Q sky130_fd_sc_hd__dfxtp_4
X_84872_ _84823_/CLK _58349_/X _84872_/Q sky130_fd_sc_hd__dfxtp_4
X_86611_ _86611_/CLK _86611_/D _72295_/A sky130_fd_sc_hd__dfxtp_4
X_83823_ _83787_/CLK _70252_/X _74790_/B sky130_fd_sc_hd__dfxtp_4
X_56771_ _56730_/X _56766_/X _56767_/X _57163_/C _57010_/A _56771_/X
+ sky130_fd_sc_hd__a41o_4
X_68757_ _68757_/A _68757_/X sky130_fd_sc_hd__buf_2
X_87591_ _88111_/CLK _87591_/D _73845_/A sky130_fd_sc_hd__dfxtp_4
X_53983_ _53978_/A _53983_/B _53983_/Y sky130_fd_sc_hd__nand2_4
X_65969_ _65969_/A _65970_/A sky130_fd_sc_hd__buf_2
X_58510_ _58510_/A _58510_/X sky130_fd_sc_hd__buf_2
X_55722_ _55245_/A _55722_/B _55722_/X sky130_fd_sc_hd__and2_4
X_67708_ _86960_/Q _67706_/X _67633_/X _67707_/X _67708_/X sky130_fd_sc_hd__a211o_4
X_86542_ _86222_/CLK _86542_/D _86542_/Q sky130_fd_sc_hd__dfxtp_4
X_52934_ _52922_/A _52954_/B _52926_/X _52934_/D _52934_/X sky130_fd_sc_hd__and4_4
X_83754_ _83421_/CLK _70527_/Y _57682_/A sky130_fd_sc_hd__dfxtp_4
X_59490_ _63396_/B _58532_/X _59490_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_524_0_CLK clkbuf_9_262_0_CLK/X _84049_/CLK sky130_fd_sc_hd__clkbuf_1
X_68688_ _68685_/X _68687_/X _68661_/X _68688_/Y sky130_fd_sc_hd__a21oi_4
X_80966_ _80821_/CLK _80966_/D _75424_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_6_15_0_CLK clkbuf_5_7_0_CLK/X clkbuf_7_31_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_58441_ _58440_/Y _58442_/A sky130_fd_sc_hd__buf_2
X_82705_ _82624_/CLK _82705_/D _82661_/D sky130_fd_sc_hd__dfxtp_4
X_55653_ _55288_/B _55288_/A _55654_/A sky130_fd_sc_hd__and2_4
X_67639_ _67522_/X _67623_/Y _67624_/X _67638_/Y _67639_/X sky130_fd_sc_hd__a211o_4
X_86473_ _86473_/CLK _86473_/D _86473_/Q sky130_fd_sc_hd__dfxtp_4
X_52865_ _52783_/A _52865_/X sky130_fd_sc_hd__buf_2
X_83685_ _83685_/CLK _70845_/Y _83685_/Q sky130_fd_sc_hd__dfxtp_4
X_80897_ _81990_/CLK _80897_/D _80897_/Q sky130_fd_sc_hd__dfxtp_4
X_88212_ _88201_/CLK _88212_/D _88212_/Q sky130_fd_sc_hd__dfxtp_4
X_54604_ _54601_/Y _54584_/X _54603_/X _85412_/D sky130_fd_sc_hd__a21oi_4
X_85424_ _85648_/CLK _85424_/D _85424_/Q sky130_fd_sc_hd__dfxtp_4
X_51816_ _51813_/Y _51793_/X _51815_/X _51816_/Y sky130_fd_sc_hd__a21oi_4
X_70650_ _53033_/B _70632_/X _70649_/Y _83733_/D sky130_fd_sc_hd__o21ai_4
X_58372_ _58372_/A _58372_/Y sky130_fd_sc_hd__inv_2
X_82636_ _88116_/CLK _83988_/Q _82636_/Q sky130_fd_sc_hd__dfxtp_4
X_55584_ _55523_/X _55610_/A sky130_fd_sc_hd__buf_2
X_52796_ _52770_/A _52818_/B sky130_fd_sc_hd__buf_2
XPHY_10 sky130_fd_sc_hd__decap_3
XPHY_21 sky130_fd_sc_hd__decap_3
X_57323_ _44277_/X _57321_/X _57322_/Y _85035_/D sky130_fd_sc_hd__o21ai_4
X_69309_ _69309_/A _88295_/Q _69309_/X sky130_fd_sc_hd__and2_4
X_88143_ _86834_/CLK _88143_/D _66683_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_539_0_CLK clkbuf_9_269_0_CLK/X _84014_/CLK sky130_fd_sc_hd__clkbuf_1
X_54535_ _54481_/A _54538_/A sky130_fd_sc_hd__buf_2
X_85355_ _86282_/CLK _85355_/D _85355_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_32 sky130_fd_sc_hd__decap_3
Xclkbuf_2_0_0_CLK clkbuf_2_1_0_CLK/A clkbuf_2_0_1_CLK/A sky130_fd_sc_hd__clkbuf_1
X_51747_ _51747_/A _51768_/A sky130_fd_sc_hd__buf_2
X_70581_ _74731_/A _71735_/A sky130_fd_sc_hd__buf_2
X_82567_ _82879_/CLK _82567_/D _82567_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_43 sky130_fd_sc_hd__decap_3
XPHY_54 sky130_fd_sc_hd__decap_3
X_41500_ _41500_/A _41500_/Y sky130_fd_sc_hd__inv_2
X_72320_ _86609_/Q _72332_/B _72320_/Y sky130_fd_sc_hd__nor2_4
XPHY_65 sky130_fd_sc_hd__decap_3
X_84306_ _84358_/CLK _63647_/Y _80379_/B sky130_fd_sc_hd__dfxtp_4
X_57254_ _57359_/A _57254_/B _57249_/X _57254_/Y sky130_fd_sc_hd__nor3_4
XPHY_76 sky130_fd_sc_hd__decap_3
X_81518_ _88175_/CLK _81518_/D _81518_/Q sky130_fd_sc_hd__dfxtp_4
X_42480_ _42612_/A _42480_/X sky130_fd_sc_hd__buf_2
X_88074_ _87821_/CLK _88074_/D _88074_/Q sky130_fd_sc_hd__dfxtp_4
X_54466_ _54385_/A _54471_/B sky130_fd_sc_hd__buf_2
X_85286_ _83013_/CLK _85286_/D _55707_/B sky130_fd_sc_hd__dfxtp_4
X_51678_ _85966_/Q _51675_/X _51677_/Y _51678_/Y sky130_fd_sc_hd__o21ai_4
XPHY_87 sky130_fd_sc_hd__decap_3
X_82498_ _82498_/CLK _82498_/D _78314_/A sky130_fd_sc_hd__dfxtp_4
XPHY_98 sky130_fd_sc_hd__decap_3
X_56205_ _56123_/A _56205_/X sky130_fd_sc_hd__buf_2
X_87025_ _87032_/CLK _44633_/Y _87025_/Q sky130_fd_sc_hd__dfxtp_4
X_53417_ _85637_/Q _53404_/X _53416_/Y _53417_/Y sky130_fd_sc_hd__o21ai_4
X_41431_ _81734_/Q _41435_/B _41431_/X sky130_fd_sc_hd__or2_4
X_72251_ _72277_/A _72251_/B _72251_/Y sky130_fd_sc_hd__nor2_4
X_84237_ _84590_/CLK _84237_/D _79568_/B sky130_fd_sc_hd__dfxtp_4
X_50629_ _86164_/Q _50626_/X _50628_/Y _50629_/Y sky130_fd_sc_hd__o21ai_4
X_81449_ _81575_/CLK _76713_/B _81449_/Q sky130_fd_sc_hd__dfxtp_4
X_57185_ _57183_/X _56703_/X _57184_/Y _57185_/Y sky130_fd_sc_hd__a21oi_4
X_54397_ _54378_/A _52706_/B _54397_/Y sky130_fd_sc_hd__nand2_4
X_71202_ _71197_/A _71226_/B _71197_/C _71202_/Y sky130_fd_sc_hd__nand3_4
X_44150_ _44149_/X _44150_/X sky130_fd_sc_hd__buf_2
X_56136_ _56140_/A _56140_/B _85290_/Q _56136_/Y sky130_fd_sc_hd__nand3_4
X_41362_ _41181_/A _41362_/X sky130_fd_sc_hd__buf_2
X_53348_ _53339_/A _53371_/B _53330_/C _52835_/D _53348_/X sky130_fd_sc_hd__and4_4
X_72182_ _72166_/X _85372_/Q _72181_/X _72182_/Y sky130_fd_sc_hd__o21ai_4
X_84168_ _84166_/CLK _84168_/D _84168_/Q sky130_fd_sc_hd__dfxtp_4
X_43101_ _43100_/X _43075_/X _40743_/X _74206_/A _43080_/X _43101_/Y
+ sky130_fd_sc_hd__o32ai_4
X_71133_ _71129_/A _71091_/B _70914_/D _71133_/Y sky130_fd_sc_hd__nand3_4
X_83119_ _86213_/CLK _74183_/X _70129_/A sky130_fd_sc_hd__dfxtp_4
X_44081_ _55549_/A _44081_/X sky130_fd_sc_hd__buf_2
X_56067_ _56058_/X _56064_/X _56066_/Y _85302_/D sky130_fd_sc_hd__o21ai_4
X_53279_ _53277_/Y _53272_/X _53278_/X _53279_/Y sky130_fd_sc_hd__a21oi_4
X_41293_ _41290_/X _82912_/Q _41292_/X _41294_/A sky130_fd_sc_hd__o21ai_4
X_76990_ _76990_/A _84414_/Q _76990_/X sky130_fd_sc_hd__xor2_4
X_84099_ _80928_/CLK _66732_/X _80923_/D sky130_fd_sc_hd__dfxtp_4
X_55018_ _55017_/X _55026_/B _55013_/C _47636_/A _55018_/X sky130_fd_sc_hd__and4_4
X_43032_ _43032_/A _43032_/Y sky130_fd_sc_hd__inv_2
X_75941_ _75933_/A _75941_/Y sky130_fd_sc_hd__inv_2
X_71064_ _71058_/A _71064_/B _71066_/C _71064_/Y sky130_fd_sc_hd__nand3_4
X_87927_ _87417_/CLK _87927_/D _87927_/Q sky130_fd_sc_hd__dfxtp_4
X_70015_ _82553_/D _70010_/X _70014_/X _83873_/D sky130_fd_sc_hd__a21bo_4
X_47840_ _47840_/A _47840_/X sky130_fd_sc_hd__buf_2
X_59826_ _59651_/A _59797_/Y _59825_/X _59680_/Y _59826_/Y sky130_fd_sc_hd__nand4_4
X_78660_ _78661_/A _82694_/Q _78663_/B sky130_fd_sc_hd__nor2_4
X_75872_ _80929_/Q _75872_/B _75875_/C sky130_fd_sc_hd__xor2_4
X_87858_ _86984_/CLK _87858_/D _68380_/A sky130_fd_sc_hd__dfxtp_4
X_77611_ _77612_/A _82108_/D _77614_/B sky130_fd_sc_hd__nor2_4
X_74823_ _74829_/A _46164_/A _74824_/A sky130_fd_sc_hd__nand2_4
X_86809_ _82899_/CLK _86809_/D _86809_/Q sky130_fd_sc_hd__dfxtp_4
X_47771_ _47771_/A _47771_/Y sky130_fd_sc_hd__inv_2
X_59757_ _59683_/A _59753_/Y _59754_/X _80526_/A _59756_/X _84704_/D
+ sky130_fd_sc_hd__o32a_4
X_78591_ _78591_/A _78602_/A _78600_/B sky130_fd_sc_hd__xor2_4
X_44983_ _85180_/Q _44982_/X _44959_/X _44983_/X sky130_fd_sc_hd__o21a_4
X_56969_ _56860_/X _56971_/B sky130_fd_sc_hd__inv_2
X_87789_ _87789_/CLK _87789_/D _69218_/B sky130_fd_sc_hd__dfxtp_4
X_49510_ _49500_/A _49516_/B _49493_/X _52724_/D _49510_/X sky130_fd_sc_hd__and4_4
X_46722_ _52637_/B _51807_/B sky130_fd_sc_hd__buf_2
X_58708_ _58618_/X _86102_/Q _58707_/X _58708_/Y sky130_fd_sc_hd__o21ai_4
X_77542_ _77542_/A _77561_/D sky130_fd_sc_hd__inv_2
X_43934_ _41433_/X _43928_/X _67975_/B _43929_/X _87192_/D sky130_fd_sc_hd__a2bb2o_4
X_74754_ _74753_/X _70637_/A _83835_/Q _74739_/B _74754_/X sky130_fd_sc_hd__and4_4
X_71966_ _71963_/Y _57592_/X _71965_/X _83312_/D sky130_fd_sc_hd__a21oi_4
X_59688_ _59687_/Y _59688_/X sky130_fd_sc_hd__buf_2
X_49441_ _49447_/A _49447_/B _49447_/C _52654_/D _49441_/X sky130_fd_sc_hd__and4_4
X_73705_ _88365_/Q _73633_/X _73704_/X _73705_/Y sky130_fd_sc_hd__o21ai_4
X_46653_ _46653_/A _46751_/A sky130_fd_sc_hd__buf_2
X_70917_ _51022_/B _70909_/X _70916_/Y _83664_/D sky130_fd_sc_hd__o21ai_4
X_58639_ _84811_/Q _58639_/Y sky130_fd_sc_hd__inv_2
X_77473_ _77473_/A _77473_/Y sky130_fd_sc_hd__inv_2
X_43865_ _43865_/A _87228_/D sky130_fd_sc_hd__inv_2
X_74685_ _57331_/A _57331_/C _74685_/C _74685_/Y sky130_fd_sc_hd__nand3_4
X_71897_ _56698_/Y _71892_/X _71896_/Y _83337_/D sky130_fd_sc_hd__o21ai_4
X_79212_ _79212_/A _72617_/A _79212_/Y sky130_fd_sc_hd__nand2_4
X_45604_ _45604_/A _45604_/B _45604_/Y sky130_fd_sc_hd__nor2_4
X_76424_ _76424_/A _76423_/X _76424_/X sky130_fd_sc_hd__xor2_4
X_42816_ _42720_/X _42816_/X sky130_fd_sc_hd__buf_2
X_49372_ _49382_/A _50893_/B _49372_/Y sky130_fd_sc_hd__nand2_4
X_73636_ _73607_/A _73636_/B _73636_/X sky130_fd_sc_hd__and2_4
X_61650_ _59433_/A _61652_/B sky130_fd_sc_hd__buf_2
X_70848_ _70848_/A _70890_/B sky130_fd_sc_hd__buf_2
X_46584_ _46575_/Y _46576_/X _46583_/Y _46584_/Y sky130_fd_sc_hd__a21boi_4
X_43796_ _41050_/X _43770_/X _69411_/B _43772_/X _87263_/D sky130_fd_sc_hd__a2bb2o_4
X_48323_ _49215_/A _48348_/A sky130_fd_sc_hd__buf_2
X_60601_ _60413_/X _60476_/Y _60598_/Y _60599_/X _60600_/Y _60601_/Y
+ sky130_fd_sc_hd__a41oi_4
X_79143_ _79143_/A _84475_/Q _79143_/X sky130_fd_sc_hd__xor2_4
X_45535_ _45535_/A _45597_/B _45535_/Y sky130_fd_sc_hd__nor2_4
X_76355_ _76381_/B _76355_/Y sky130_fd_sc_hd__inv_2
X_42747_ _41230_/X _42745_/X _68918_/B _42746_/X _42747_/X sky130_fd_sc_hd__a2bb2o_4
X_61581_ _61305_/A _61580_/X _72583_/C _61581_/Y sky130_fd_sc_hd__nand3_4
X_73567_ _73165_/A _73588_/A sky130_fd_sc_hd__buf_2
X_70779_ _70869_/A _70779_/B _70791_/C _70791_/D _70779_/Y sky130_fd_sc_hd__nand4_4
X_63320_ _79197_/B _79198_/A sky130_fd_sc_hd__inv_2
X_75306_ _75291_/X _75292_/Y _75294_/A _75306_/Y sky130_fd_sc_hd__a21boi_4
X_48254_ _48244_/A _50302_/B _48254_/Y sky130_fd_sc_hd__nand2_4
X_60532_ _60532_/A _60532_/Y sky130_fd_sc_hd__inv_2
X_72518_ _72502_/A _72597_/B sky130_fd_sc_hd__buf_2
X_79074_ _79074_/A _79089_/A _79087_/B sky130_fd_sc_hd__xor2_4
X_45466_ _45463_/Y _45465_/Y _44901_/X _45466_/X sky130_fd_sc_hd__o21a_4
X_76286_ _76284_/X _76286_/B _81611_/D sky130_fd_sc_hd__xor2_4
X_42678_ _42677_/Y _42678_/Y sky130_fd_sc_hd__inv_2
X_73498_ _73449_/X _85572_/Q _73450_/X _73497_/X _73498_/X sky130_fd_sc_hd__a211o_4
X_47205_ _53426_/B _51222_/B sky130_fd_sc_hd__buf_2
X_78025_ _78024_/Y _78009_/A _78025_/X sky130_fd_sc_hd__and2_4
X_44417_ _44404_/X _44405_/X _41545_/X _87119_/Q _44406_/X _44418_/A
+ sky130_fd_sc_hd__o32ai_4
X_75237_ _75224_/Y _75225_/Y _75226_/Y _75237_/X sky130_fd_sc_hd__o21a_4
X_63251_ _58490_/A _63250_/X _58268_/A _62999_/X _63251_/X sky130_fd_sc_hd__o22a_4
X_41629_ _82913_/Q _41563_/B _41629_/X sky130_fd_sc_hd__or2_4
X_48185_ _48182_/Y _48175_/X _48184_/Y _48185_/Y sky130_fd_sc_hd__a21boi_4
X_60463_ _60570_/A _60488_/B sky130_fd_sc_hd__buf_2
X_72449_ _64758_/X _85317_/Q _57763_/X _72449_/X sky130_fd_sc_hd__o21a_4
X_45397_ _44932_/A _45397_/X sky130_fd_sc_hd__buf_2
X_62202_ _61315_/A _62556_/A _62576_/C _62560_/D _62202_/Y sky130_fd_sc_hd__nand4_4
X_47136_ _53390_/B _52876_/B sky130_fd_sc_hd__buf_2
X_44348_ _44330_/X _44331_/X _41705_/X _87153_/Q _44332_/X _44348_/Y
+ sky130_fd_sc_hd__o32ai_4
X_63182_ _63157_/X _63182_/B _63147_/C _63181_/X _63182_/X sky130_fd_sc_hd__and4_4
X_75168_ _80776_/Q _81032_/D _75168_/X sky130_fd_sc_hd__xor2_4
X_60394_ _60393_/X _60440_/A sky130_fd_sc_hd__buf_2
X_62133_ _62144_/A _62121_/X _78054_/B _62133_/Y sky130_fd_sc_hd__nor3_4
X_74119_ _74119_/A _73370_/B _74119_/Y sky130_fd_sc_hd__nor2_4
X_47067_ _47067_/A _47039_/B _47048_/C _52835_/D _47067_/X sky130_fd_sc_hd__and4_4
X_44279_ _44139_/X _44141_/X _44142_/X _44279_/D _44279_/Y sky130_fd_sc_hd__nand4_4
X_67990_ _67986_/X _67989_/X _67917_/X _67990_/X sky130_fd_sc_hd__a21o_4
X_79976_ _79974_/Y _79975_/Y _79976_/Y sky130_fd_sc_hd__nand2_4
X_75099_ _75099_/A _75099_/Y sky130_fd_sc_hd__inv_2
X_46018_ _40523_/Y _46007_/X _67201_/B _46008_/X _86812_/D sky130_fd_sc_hd__a2bb2o_4
X_66941_ _68474_/A _66942_/A sky130_fd_sc_hd__buf_2
X_62064_ _59766_/X _62065_/D sky130_fd_sc_hd__buf_2
X_78927_ _82735_/Q _78927_/B _82703_/D sky130_fd_sc_hd__xor2_4
X_61015_ _60891_/Y _61012_/Y _60944_/Y _61013_/Y _61014_/Y _61015_/Y
+ sky130_fd_sc_hd__a41oi_4
X_69660_ _43133_/A _68636_/X _68517_/X _69659_/X _69660_/X sky130_fd_sc_hd__a211o_4
X_66872_ _66866_/X _66870_/X _66871_/X _66872_/Y sky130_fd_sc_hd__a21oi_4
X_78858_ _78855_/X _78856_/Y _78857_/X _78858_/Y sky130_fd_sc_hd__a21oi_4
X_68611_ _83968_/Q _68586_/X _68610_/X _68611_/X sky130_fd_sc_hd__a21bo_4
X_65823_ _65820_/X _65822_/X _65642_/X _65827_/A sky130_fd_sc_hd__a21o_4
X_77809_ _77809_/A _77819_/A _77809_/Y sky130_fd_sc_hd__nor2_4
X_69591_ _83912_/Q _69564_/X _69590_/X _69591_/X sky130_fd_sc_hd__a21bo_4
X_47969_ _47988_/A _47969_/B _47969_/Y sky130_fd_sc_hd__nand2_4
X_78789_ _78788_/Y _78789_/Y sky130_fd_sc_hd__inv_2
X_49708_ _49708_/A _49697_/B _49685_/C _47218_/D _49708_/X sky130_fd_sc_hd__and4_4
X_68542_ _69190_/A _68542_/X sky130_fd_sc_hd__buf_2
X_80820_ _81994_/CLK _83964_/Q _80820_/Q sky130_fd_sc_hd__dfxtp_4
X_65754_ _64599_/X _83060_/Q _64600_/X _65753_/X _65754_/X sky130_fd_sc_hd__a211o_4
X_50980_ _50977_/Y _50957_/X _50979_/X _86096_/D sky130_fd_sc_hd__a21oi_4
X_62966_ _61665_/B _62936_/X _62982_/C _62908_/X _62966_/Y sky130_fd_sc_hd__nand4_4
X_64705_ _44244_/A _64706_/A sky130_fd_sc_hd__buf_2
X_49639_ _86350_/Q _49632_/X _49638_/Y _49639_/Y sky130_fd_sc_hd__o21ai_4
X_61917_ _61871_/A _61949_/B _61949_/C _63147_/B _61917_/X sky130_fd_sc_hd__and4_4
X_80751_ _80746_/CLK _80751_/D _81127_/D sky130_fd_sc_hd__dfxtp_4
X_68473_ _69611_/A _68473_/X sky130_fd_sc_hd__buf_2
X_65685_ _65484_/A _65685_/X sky130_fd_sc_hd__buf_2
X_62897_ _62897_/A _62897_/Y sky130_fd_sc_hd__inv_2
X_67424_ _67419_/X _67422_/X _67423_/X _67424_/Y sky130_fd_sc_hd__a21oi_4
X_52650_ _52646_/Y _52647_/X _52649_/X _52650_/Y sky130_fd_sc_hd__a21oi_4
X_83470_ _85957_/CLK _83470_/D _47779_/A sky130_fd_sc_hd__dfxtp_4
X_64636_ _64636_/A _66104_/A sky130_fd_sc_hd__buf_2
X_61848_ _61837_/X _61840_/X _61847_/Y _58177_/A _61815_/X _61848_/Y
+ sky130_fd_sc_hd__o32ai_4
X_80682_ _81065_/CLK _80682_/D _80682_/Q sky130_fd_sc_hd__dfxtp_4
X_51601_ _85980_/Q _51594_/X _51600_/Y _51601_/Y sky130_fd_sc_hd__o21ai_4
X_82421_ _82463_/CLK _82453_/Q _78586_/A sky130_fd_sc_hd__dfxtp_4
X_67355_ _67354_/X _67355_/X sky130_fd_sc_hd__buf_2
X_52581_ _52578_/Y _52532_/X _52580_/X _52581_/Y sky130_fd_sc_hd__a21oi_4
X_64567_ _64567_/A _64667_/A sky130_fd_sc_hd__buf_2
X_61779_ _61364_/B _61795_/B _61795_/C _61778_/X _61779_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_4_5_1_CLK clkbuf_4_5_0_CLK/X clkbuf_4_5_1_CLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_608 sky130_fd_sc_hd__decap_3
X_54320_ _54320_/A _54320_/X sky130_fd_sc_hd__buf_2
XPHY_619 sky130_fd_sc_hd__decap_3
X_66306_ _66231_/X _66319_/B _84142_/Q _66306_/X sky130_fd_sc_hd__and3_4
X_85140_ _85138_/CLK _56641_/X _85140_/Q sky130_fd_sc_hd__dfxtp_4
X_51532_ _51504_/A _51553_/B sky130_fd_sc_hd__buf_2
X_63518_ _63515_/Y _63516_/X _63517_/Y _63518_/Y sky130_fd_sc_hd__a21oi_4
X_82352_ _82299_/CLK _77152_/X _48018_/A sky130_fd_sc_hd__dfxtp_4
X_67286_ _87861_/Q _67236_/X _67284_/X _67285_/X _67286_/X sky130_fd_sc_hd__a211o_4
X_64498_ _64493_/X _64494_/X _64495_/X _64497_/Y _64440_/X _64498_/X
+ sky130_fd_sc_hd__o41a_4
X_81303_ _81801_/CLK _76991_/X _81303_/Q sky130_fd_sc_hd__dfxtp_4
X_69025_ _57716_/A _69025_/X sky130_fd_sc_hd__buf_2
X_54251_ _54961_/A _53080_/B _54251_/Y sky130_fd_sc_hd__nand2_4
X_66237_ _58784_/A _66237_/X sky130_fd_sc_hd__buf_2
X_85071_ _85071_/CLK _85071_/D _85071_/Q sky130_fd_sc_hd__dfxtp_4
X_51463_ _51461_/Y _51448_/X _51462_/X _86006_/D sky130_fd_sc_hd__a21oi_4
X_63449_ _58429_/Y _63436_/X _61421_/A _63437_/X _63449_/X sky130_fd_sc_hd__a2bb2o_4
X_82283_ _82301_/CLK _82283_/D _41057_/A sky130_fd_sc_hd__dfxtp_4
X_53202_ _53097_/X _53211_/B sky130_fd_sc_hd__buf_2
X_84022_ _81169_/CLK _68166_/X _82062_/D sky130_fd_sc_hd__dfxtp_4
X_50414_ _50481_/A _48401_/B _50414_/Y sky130_fd_sc_hd__nand2_4
X_81234_ _81233_/CLK _81042_/Q _47674_/A sky130_fd_sc_hd__dfxtp_4
X_54182_ _54191_/A _54186_/B _54191_/C _53015_/D _54182_/X sky130_fd_sc_hd__and4_4
X_66168_ _65074_/A _66168_/B _66168_/X sky130_fd_sc_hd__and2_4
X_51394_ _51758_/A _51394_/B _51394_/Y sky130_fd_sc_hd__nand2_4
X_53133_ _53133_/A _53133_/B _53133_/C _53133_/D _53133_/X sky130_fd_sc_hd__and4_4
X_65119_ _64616_/A _65227_/A sky130_fd_sc_hd__buf_2
X_50345_ _50398_/A _52047_/B _50345_/Y sky130_fd_sc_hd__nand2_4
X_81165_ _81179_/CLK _74927_/B _41563_/A sky130_fd_sc_hd__dfxtp_4
X_58990_ _58990_/A _58990_/Y sky130_fd_sc_hd__inv_2
X_66099_ _66095_/X _66098_/X _66057_/X _66099_/X sky130_fd_sc_hd__a21o_4
X_80116_ _80117_/B _80103_/Y _80116_/X sky130_fd_sc_hd__or2_4
X_53064_ _53061_/Y _53056_/X _53063_/X _85704_/D sky130_fd_sc_hd__a21oi_4
X_57941_ _57939_/X _86002_/Q _57940_/X _57941_/Y sky130_fd_sc_hd__o21ai_4
X_69927_ _69515_/Y _69916_/X _69870_/X _69926_/Y _69927_/X sky130_fd_sc_hd__a211o_4
X_50276_ _50273_/Y _50274_/X _50275_/Y _50276_/Y sky130_fd_sc_hd__a21boi_4
X_85973_ _84787_/CLK _85973_/D _85973_/Q sky130_fd_sc_hd__dfxtp_4
X_81096_ _82220_/CLK _79624_/X _81096_/Q sky130_fd_sc_hd__dfxtp_4
X_52015_ _52014_/X _50310_/B _52015_/Y sky130_fd_sc_hd__nand2_4
X_87712_ _87210_/CLK _87712_/D _67793_/B sky130_fd_sc_hd__dfxtp_4
X_84924_ _85375_/CLK _84924_/D _58108_/A sky130_fd_sc_hd__dfxtp_4
X_80047_ _57996_/Y _65745_/C _80046_/Y _80047_/X sky130_fd_sc_hd__o21a_4
X_57872_ _57872_/A _57872_/X sky130_fd_sc_hd__buf_2
X_69858_ _81964_/D _69831_/X _69857_/X _83892_/D sky130_fd_sc_hd__a21bo_4
X_59611_ _59557_/A _43995_/A _59609_/D _59611_/X sky130_fd_sc_hd__and3_4
X_56823_ _56821_/X _56738_/X _56822_/Y _56823_/Y sky130_fd_sc_hd__o21ai_4
X_68809_ _86990_/Q _68707_/X _68762_/X _68808_/X _68809_/X sky130_fd_sc_hd__a211o_4
X_87643_ _86920_/CLK _42936_/Y _67912_/B sky130_fd_sc_hd__dfxtp_4
X_84855_ _84263_/CLK _58413_/X _84855_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_463_0_CLK clkbuf_9_231_0_CLK/X _84787_/CLK sky130_fd_sc_hd__clkbuf_1
X_69789_ _64665_/A _69791_/A sky130_fd_sc_hd__buf_2
X_71820_ _71804_/Y _83363_/Q _71819_/X _83363_/D sky130_fd_sc_hd__a21o_4
X_59542_ _44216_/X _44217_/X _44008_/A _59543_/A sky130_fd_sc_hd__a21oi_4
X_83806_ _81807_/CLK _70300_/X _74783_/A sky130_fd_sc_hd__dfxtp_4
X_56754_ _56736_/X _56764_/C sky130_fd_sc_hd__inv_2
X_87574_ _87542_/CLK _87574_/D _43103_/A sky130_fd_sc_hd__dfxtp_4
X_41980_ _41980_/A _41980_/Y sky130_fd_sc_hd__inv_2
X_53966_ _53942_/A _46313_/Y _53966_/Y sky130_fd_sc_hd__nand2_4
X_84786_ _86372_/CLK _84786_/D _84786_/Q sky130_fd_sc_hd__dfxtp_4
X_81998_ _81985_/CLK _81998_/D _81998_/Q sky130_fd_sc_hd__dfxtp_4
X_55705_ _85190_/Q _55272_/A _55128_/X _55704_/X _55705_/X sky130_fd_sc_hd__a211o_4
X_86525_ _86525_/CLK _86525_/D _86525_/Q sky130_fd_sc_hd__dfxtp_4
X_52917_ _52915_/Y _52892_/X _52916_/X _52917_/Y sky130_fd_sc_hd__a21oi_4
X_40931_ _40931_/A _40931_/X sky130_fd_sc_hd__buf_2
X_71751_ _71178_/A _71753_/B _71744_/C _71744_/D _71751_/Y sky130_fd_sc_hd__nand4_4
X_83737_ _83736_/CLK _83737_/D _47372_/A sky130_fd_sc_hd__dfxtp_4
X_59473_ _84722_/Q _59474_/A sky130_fd_sc_hd__inv_2
X_56685_ _56672_/Y _56685_/B _56685_/X sky130_fd_sc_hd__xor2_4
X_80949_ _81211_/CLK _80949_/D _80949_/Q sky130_fd_sc_hd__dfxtp_4
X_53897_ _53956_/A _53898_/A sky130_fd_sc_hd__buf_2
X_70702_ _70712_/A _70866_/A sky130_fd_sc_hd__buf_2
X_58424_ _84851_/Q _58424_/Y sky130_fd_sc_hd__inv_2
X_43650_ _43649_/X _87327_/D sky130_fd_sc_hd__inv_2
X_55636_ _85121_/Q _55617_/X _44052_/A _55635_/Y _55636_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_478_0_CLK clkbuf_9_239_0_CLK/X _86091_/CLK sky130_fd_sc_hd__clkbuf_1
X_74470_ _74442_/X _48602_/Y _74470_/Y sky130_fd_sc_hd__nand2_4
X_86456_ _83303_/CLK _48980_/Y _86456_/Q sky130_fd_sc_hd__dfxtp_4
X_40862_ _40835_/X _40836_/X _40861_/X _88321_/Q _40832_/X _40862_/Y
+ sky130_fd_sc_hd__o32ai_4
X_52848_ _52821_/A _52848_/X sky130_fd_sc_hd__buf_2
X_71682_ _71669_/A _71682_/Y sky130_fd_sc_hd__inv_2
X_83668_ _86091_/CLK _70902_/Y _83668_/Q sky130_fd_sc_hd__dfxtp_4
X_42601_ _42568_/X _40881_/A _42477_/X _42600_/Y _42571_/X _42601_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73421_ _73704_/A _73421_/X sky130_fd_sc_hd__buf_2
X_85407_ _85407_/CLK _54631_/Y _85407_/Q sky130_fd_sc_hd__dfxtp_4
X_70633_ _71115_/C _70412_/X _70933_/B _71287_/C _70633_/X sky130_fd_sc_hd__and4_4
X_58355_ _63316_/A _61656_/A sky130_fd_sc_hd__buf_2
X_82619_ _82589_/CLK _79035_/B _82619_/Q sky130_fd_sc_hd__dfxtp_4
X_43581_ _40591_/B _46612_/A sky130_fd_sc_hd__buf_2
X_55567_ _55534_/A _56604_/B _55567_/X sky130_fd_sc_hd__and2_4
X_86387_ _83673_/CLK _49442_/Y _58750_/B sky130_fd_sc_hd__dfxtp_4
X_52779_ _52775_/A _52775_/B _52775_/C _52779_/D _52779_/X sky130_fd_sc_hd__and4_4
X_40793_ _40793_/A _40793_/X sky130_fd_sc_hd__buf_2
X_83599_ _86145_/CLK _83599_/D _83599_/Q sky130_fd_sc_hd__dfxtp_4
X_57306_ _57304_/Y _57305_/Y _56995_/X _57306_/Y sky130_fd_sc_hd__a21oi_4
X_45320_ _45317_/X _45319_/Y _45275_/X _45320_/Y sky130_fd_sc_hd__a21oi_4
X_76140_ _76138_/Y _76134_/Y _76139_/Y _76143_/A sky130_fd_sc_hd__o21ai_4
X_88126_ _88128_/CLK _88126_/D _88126_/Q sky130_fd_sc_hd__dfxtp_4
X_54518_ _54518_/A _47053_/A _54518_/Y sky130_fd_sc_hd__nand2_4
X_42532_ _42521_/X _42522_/X _40743_/X _69052_/A _42506_/X _42532_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73352_ _73352_/A _73353_/A sky130_fd_sc_hd__buf_2
X_85338_ _85338_/CLK _55001_/Y _85338_/Q sky130_fd_sc_hd__dfxtp_4
X_70564_ _71863_/A _70549_/X _70568_/C _70568_/D _70564_/Y sky130_fd_sc_hd__nor4_4
X_58286_ _58282_/X _58283_/Y _58285_/Y _84888_/D sky130_fd_sc_hd__a21oi_4
X_55498_ _55492_/X _55498_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_401_0_CLK clkbuf_9_200_0_CLK/X _82253_/CLK sky130_fd_sc_hd__clkbuf_1
X_72303_ _72417_/A _72303_/X sky130_fd_sc_hd__buf_2
X_45251_ _56253_/C _45222_/X _45250_/X _45251_/Y sky130_fd_sc_hd__o21ai_4
X_57237_ _56561_/X _57322_/B _56931_/X _85057_/Q _57236_/X _85057_/D
+ sky130_fd_sc_hd__a32o_4
X_76071_ _81718_/D _76062_/B _76071_/Y sky130_fd_sc_hd__nand2_4
X_42463_ _42463_/A _42463_/X sky130_fd_sc_hd__buf_2
X_88057_ _88062_/CLK _42051_/Y _88057_/Q sky130_fd_sc_hd__dfxtp_4
X_54449_ _54435_/A _54440_/B _54429_/C _54449_/D _54449_/X sky130_fd_sc_hd__and4_4
X_73283_ _73257_/X _86189_/Q _73205_/X _73282_/X _73283_/X sky130_fd_sc_hd__a211o_4
X_85269_ _85269_/CLK _56224_/Y _56223_/C sky130_fd_sc_hd__dfxtp_4
X_70495_ _70495_/A _70758_/B sky130_fd_sc_hd__buf_2
X_44202_ _44202_/A _44185_/X _44202_/X sky130_fd_sc_hd__or2_4
X_75022_ _75005_/Y _75019_/X _75021_/Y _75023_/B sky130_fd_sc_hd__a21oi_4
X_41414_ _41414_/A _41435_/B _41414_/X sky130_fd_sc_hd__or2_4
X_87008_ _88283_/CLK _44668_/X _87008_/Q sky130_fd_sc_hd__dfxtp_4
X_72234_ _72172_/X _72232_/Y _72233_/Y _72189_/X _72176_/X _72234_/X
+ sky130_fd_sc_hd__o32a_4
X_45182_ _45182_/A _45182_/B _45182_/Y sky130_fd_sc_hd__nand2_4
X_57168_ _56797_/A _44239_/A _56796_/Y _57175_/A sky130_fd_sc_hd__nand3_4
X_42394_ _40404_/X _42388_/X _87884_/Q _42389_/X _87884_/D sky130_fd_sc_hd__a2bb2o_4
X_44133_ _73614_/A _44130_/X _44133_/Y sky130_fd_sc_hd__nor2_4
X_79830_ _79804_/X _79820_/B _79819_/A _79818_/Y _79830_/X sky130_fd_sc_hd__o22a_4
X_56119_ _56138_/B _55773_/D _55801_/B _55801_/C _56120_/B sky130_fd_sc_hd__nand4_4
X_41345_ _41513_/A _82902_/Q _41345_/X sky130_fd_sc_hd__or2_4
X_72165_ _72165_/A _72165_/Y sky130_fd_sc_hd__inv_2
X_49990_ _49995_/A _49973_/B _50005_/C _53203_/D _49990_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_416_0_CLK clkbuf_9_208_0_CLK/X _82443_/CLK sky130_fd_sc_hd__clkbuf_1
X_57099_ _57221_/A _57099_/X sky130_fd_sc_hd__buf_2
Xclkbuf_opt_0_CLK _84835_/CLK _84839_/CLK sky130_fd_sc_hd__clkbuf_16
X_71116_ _71115_/X _71117_/A sky130_fd_sc_hd__buf_2
X_48941_ _48933_/Y _48935_/X _48940_/X _48941_/Y sky130_fd_sc_hd__a21oi_4
X_44064_ _44063_/X _44064_/X sky130_fd_sc_hd__buf_2
X_79761_ _79761_/A _79761_/B _79761_/Y sky130_fd_sc_hd__nand2_4
X_41276_ _41242_/X _40751_/A _41275_/X _41276_/X sky130_fd_sc_hd__o21a_4
X_72096_ _72091_/X _49166_/Y _72096_/Y sky130_fd_sc_hd__nand2_4
X_76973_ _61057_/C _62606_/C _76973_/X sky130_fd_sc_hd__xor2_4
X_43015_ _43014_/Y _43030_/A sky130_fd_sc_hd__buf_2
X_78712_ _78712_/A _78712_/Y sky130_fd_sc_hd__inv_2
X_71047_ _71046_/X _71047_/X sky130_fd_sc_hd__buf_2
X_75924_ _81698_/D _75924_/B _75925_/B sky130_fd_sc_hd__xor2_4
X_48872_ _50056_/A _48872_/B _48872_/Y sky130_fd_sc_hd__nand2_4
X_79692_ _79692_/A _79692_/B _79692_/Y sky130_fd_sc_hd__xnor2_4
X_47823_ _49374_/A _49364_/B _50886_/C _53261_/D _47823_/X sky130_fd_sc_hd__and4_4
X_59809_ _61966_/A _59810_/A sky130_fd_sc_hd__buf_2
X_78643_ _78639_/Y _78642_/Y _82776_/D sky130_fd_sc_hd__xor2_4
X_75855_ _75840_/B _75855_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_90_0_CLK clkbuf_8_91_0_CLK/A clkbuf_8_90_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_62820_ _57680_/A _62808_/X _62768_/X _62818_/X _62819_/X _62820_/Y
+ sky130_fd_sc_hd__a41oi_4
X_74806_ _83793_/Q _74720_/C _74744_/X _74745_/D _74810_/A sky130_fd_sc_hd__nand4_4
X_47754_ _72405_/A _47714_/X _47753_/Y _47754_/Y sky130_fd_sc_hd__o21ai_4
X_78574_ _78569_/X _78572_/Y _78574_/C _78575_/B sky130_fd_sc_hd__nand3_4
X_44966_ _44966_/A _44966_/Y sky130_fd_sc_hd__inv_2
X_75786_ _81098_/Q _75786_/B _75786_/X sky130_fd_sc_hd__xor2_4
X_72998_ _72997_/X _73191_/B _72998_/X sky130_fd_sc_hd__and2_4
X_46705_ _46845_/A _46717_/B sky130_fd_sc_hd__buf_2
X_77525_ _77512_/A _77523_/Y _77524_/Y _77525_/X sky130_fd_sc_hd__a21bo_4
X_43917_ _43896_/X _43917_/X sky130_fd_sc_hd__buf_2
X_74737_ _70625_/Y _71266_/A _71263_/D _74738_/A sky130_fd_sc_hd__and3_4
X_62751_ _57652_/X _62749_/X _62708_/X _62699_/X _62750_/X _62751_/Y
+ sky130_fd_sc_hd__a41oi_4
X_47685_ _47681_/Y _47651_/X _47684_/X _86609_/D sky130_fd_sc_hd__a21oi_4
X_71949_ _74527_/A _70766_/C _71349_/D _71894_/Y _71949_/Y sky130_fd_sc_hd__nand4_4
X_44897_ _80672_/Q _45757_/A sky130_fd_sc_hd__buf_2
X_49424_ _49451_/A _49447_/B sky130_fd_sc_hd__buf_2
X_61702_ _59721_/X _61770_/A sky130_fd_sc_hd__buf_2
X_46636_ _86719_/Q _46622_/X _46635_/Y _46636_/Y sky130_fd_sc_hd__o21ai_4
X_65470_ _65669_/A _65470_/X sky130_fd_sc_hd__buf_2
X_77456_ _77468_/A _77468_/B _77456_/X sky130_fd_sc_hd__xor2_4
X_43848_ _43846_/X _43824_/X _41193_/X _87236_/Q _43847_/X _43848_/Y
+ sky130_fd_sc_hd__o32ai_4
X_62682_ _62681_/X _62694_/C sky130_fd_sc_hd__buf_2
X_74668_ _74673_/A _57153_/A _74667_/Y _74669_/A sky130_fd_sc_hd__o21ai_4
X_64421_ _64421_/A _64421_/X sky130_fd_sc_hd__buf_2
X_76407_ _81363_/Q _76407_/B _76407_/X sky130_fd_sc_hd__xor2_4
X_49355_ _49353_/Y _48194_/X _49354_/Y _86403_/D sky130_fd_sc_hd__a21boi_4
X_61633_ _61627_/Y _61629_/Y _61594_/X _61630_/Y _61632_/Y _61633_/X
+ sky130_fd_sc_hd__a41o_4
X_73619_ _47853_/Y _73618_/Y _73619_/X sky130_fd_sc_hd__xor2_4
X_46567_ _46567_/A _46527_/X _46567_/X sky130_fd_sc_hd__or2_4
X_77387_ _77387_/A _77387_/B _77387_/X sky130_fd_sc_hd__or2_4
X_43779_ _43774_/X _43760_/X _41004_/X _87271_/Q _43776_/X _43779_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74599_ _74552_/X _74599_/X sky130_fd_sc_hd__buf_2
X_48306_ _66242_/B _48293_/X _48305_/Y _48306_/Y sky130_fd_sc_hd__o21ai_4
X_67140_ _80906_/D _67092_/X _67139_/X _67140_/X sky130_fd_sc_hd__a21bo_4
X_79126_ _60612_/C _84458_/Q _79126_/X sky130_fd_sc_hd__xor2_4
X_45518_ _45515_/Y _45516_/X _45471_/X _45517_/Y _45518_/X sky130_fd_sc_hd__a211o_4
X_76338_ _76338_/A _76338_/B _76356_/A sky130_fd_sc_hd__xor2_4
X_64352_ _64304_/A _64303_/X _84957_/Q _64318_/D _64352_/X sky130_fd_sc_hd__and4_4
X_49286_ _48535_/A _49287_/A sky130_fd_sc_hd__buf_2
X_61564_ _61564_/A _61564_/Y sky130_fd_sc_hd__inv_2
X_46498_ _52528_/A _46487_/B _46472_/C _46498_/X sky130_fd_sc_hd__and3_4
X_63303_ _63248_/X _63298_/Y _63299_/X _63300_/Y _63302_/Y _63303_/X
+ sky130_fd_sc_hd__a41o_4
X_48237_ _73833_/B _48203_/X _48236_/Y _48237_/Y sky130_fd_sc_hd__o21ai_4
X_60515_ _60515_/A _60515_/B _60515_/C _60515_/Y sky130_fd_sc_hd__nand3_4
X_67071_ _67023_/A _67071_/B _67071_/X sky130_fd_sc_hd__and2_4
X_79057_ _79057_/A _79057_/B _79057_/C _79058_/B sky130_fd_sc_hd__nand3_4
X_45449_ _55599_/B _45876_/B _44919_/X _45449_/Y sky130_fd_sc_hd__o21ai_4
X_64283_ _64273_/A _64273_/B _64283_/C _64304_/D _64283_/X sky130_fd_sc_hd__and4_4
X_76269_ _76268_/D _76237_/Y _76236_/X _76269_/Y sky130_fd_sc_hd__nand3_4
X_61495_ _61489_/Y _61491_/Y _61464_/X _61492_/Y _61494_/Y _61495_/X
+ sky130_fd_sc_hd__a41o_4
X_66022_ _65992_/A _66022_/B _66022_/X sky130_fd_sc_hd__and2_4
X_78008_ _82256_/Q _81968_/Q _78024_/A sky130_fd_sc_hd__xnor2_4
X_63234_ _60522_/A _63234_/X sky130_fd_sc_hd__buf_2
X_60446_ _60408_/C _60408_/A _60406_/X _60439_/X _60440_/A _60515_/A
+ sky130_fd_sc_hd__a32oi_4
X_48168_ _48162_/A _48897_/A sky130_fd_sc_hd__buf_2
X_47119_ _82380_/Q _54559_/D sky130_fd_sc_hd__inv_2
X_63165_ _60466_/X _63165_/X sky130_fd_sc_hd__buf_2
X_48099_ _52573_/B _48099_/X sky130_fd_sc_hd__buf_2
X_60377_ _60630_/A _60171_/A _60630_/C _60171_/B _60392_/A sky130_fd_sc_hd__and4_4
Xclkbuf_8_43_0_CLK clkbuf_8_43_0_CLK/A clkbuf_9_87_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_50130_ _50105_/A _50131_/A sky130_fd_sc_hd__buf_2
X_62116_ _62142_/A _62110_/Y _62112_/Y _62115_/Y _62116_/Y sky130_fd_sc_hd__nand4_4
X_67973_ _87960_/Q _67950_/X _67879_/X _67972_/X _67973_/X sky130_fd_sc_hd__a211o_4
X_63096_ _60452_/X _63097_/A sky130_fd_sc_hd__buf_2
X_79959_ _79941_/Y _79959_/Y sky130_fd_sc_hd__inv_2
X_69712_ _69709_/X _69711_/X _69678_/X _69712_/X sky130_fd_sc_hd__a21o_4
X_50061_ _48836_/A _50061_/X sky130_fd_sc_hd__buf_2
X_66924_ _80915_/D _66850_/X _66923_/X _66924_/X sky130_fd_sc_hd__a21bo_4
X_62047_ _62142_/A _62047_/B _62047_/C _62047_/D _62047_/Y sky130_fd_sc_hd__nand4_4
X_82970_ _82206_/CLK _82778_/Q _82970_/Q sky130_fd_sc_hd__dfxtp_4
X_69643_ _81980_/D _69632_/X _69642_/X _83908_/D sky130_fd_sc_hd__a21bo_4
X_81921_ _82124_/CLK _81921_/D _81921_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_58_0_CLK clkbuf_8_59_0_CLK/A clkbuf_8_58_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_66855_ _87431_/Q _66762_/X _66764_/X _66854_/X _66855_/X sky130_fd_sc_hd__a211o_4
X_53820_ _85562_/Q _53816_/X _53819_/Y _53820_/Y sky130_fd_sc_hd__o21ai_4
X_65806_ _65158_/A _65807_/A sky130_fd_sc_hd__buf_2
X_84640_ _84640_/CLK _60295_/Y _79784_/A sky130_fd_sc_hd__dfxtp_4
X_81852_ _82515_/CLK _81852_/D _77612_/A sky130_fd_sc_hd__dfxtp_4
X_69574_ _69571_/X _69574_/B _69574_/Y sky130_fd_sc_hd__nand2_4
X_66786_ _87434_/Q _66762_/X _66764_/X _66785_/X _66786_/X sky130_fd_sc_hd__a211o_4
X_63998_ _84841_/Q _63934_/X _63949_/C _64027_/D _63998_/Y sky130_fd_sc_hd__nand4_4
X_80803_ _83973_/CLK _80803_/D _75726_/B sky130_fd_sc_hd__dfxtp_4
X_68525_ _68525_/A _68525_/B _68525_/Y sky130_fd_sc_hd__nand2_4
X_53751_ _85575_/Q _53729_/X _53750_/Y _53751_/Y sky130_fd_sc_hd__o21ai_4
X_65737_ _65732_/X _65736_/X _65614_/X _65737_/X sky130_fd_sc_hd__a21o_4
X_84571_ _84624_/CLK _60769_/X _78066_/A sky130_fd_sc_hd__dfxtp_4
X_50963_ _50963_/A _50963_/B _50963_/C _52654_/D _50963_/X sky130_fd_sc_hd__and4_4
X_62949_ _60292_/A _62949_/B _62947_/Y _62948_/Y _62949_/Y sky130_fd_sc_hd__nand4_4
X_81783_ _81783_/CLK _76130_/X _48472_/A sky130_fd_sc_hd__dfxtp_4
X_86310_ _86627_/CLK _49863_/Y _58081_/B sky130_fd_sc_hd__dfxtp_4
X_52702_ _52619_/A _52702_/X sky130_fd_sc_hd__buf_2
X_83522_ _83526_/CLK _71370_/X _83522_/Q sky130_fd_sc_hd__dfxtp_4
X_56470_ _56005_/X _56468_/X _56469_/Y _56470_/Y sky130_fd_sc_hd__o21ai_4
X_68456_ _68409_/A _88272_/Q _68456_/X sky130_fd_sc_hd__and2_4
X_80734_ _82211_/CLK _75920_/X _80702_/D sky130_fd_sc_hd__dfxtp_4
X_87290_ _88062_/CLK _43735_/X _87290_/Q sky130_fd_sc_hd__dfxtp_4
X_53682_ _53679_/Y _53680_/X _53681_/X _85589_/D sky130_fd_sc_hd__a21oi_4
X_65668_ _65484_/X _86193_/Q _65534_/X _65667_/X _65668_/X sky130_fd_sc_hd__a211o_4
X_50894_ _86111_/Q _50882_/X _50893_/Y _50894_/Y sky130_fd_sc_hd__o21ai_4
X_55421_ _56807_/A _55421_/B _56807_/C _55421_/Y sky130_fd_sc_hd__nand3_4
X_67407_ _87984_/Q _67355_/X _67405_/X _67406_/X _67407_/X sky130_fd_sc_hd__a211o_4
X_86241_ _83161_/CLK _50217_/Y _86241_/Q sky130_fd_sc_hd__dfxtp_4
X_52633_ _85783_/Q _52629_/X _52632_/Y _52633_/Y sky130_fd_sc_hd__o21ai_4
X_64619_ _64619_/A _64619_/X sky130_fd_sc_hd__buf_2
X_83453_ _83457_/CLK _71569_/X _83453_/Q sky130_fd_sc_hd__dfxtp_4
X_80665_ _86770_/CLK _80665_/D _80665_/Q sky130_fd_sc_hd__dfxtp_4
X_68387_ _69001_/A _68387_/B _68387_/Y sky130_fd_sc_hd__nor2_4
X_65599_ _65599_/A _65599_/B _65599_/Y sky130_fd_sc_hd__nand2_4
X_58140_ _58618_/A _58140_/X sky130_fd_sc_hd__buf_2
X_82404_ _82443_/CLK _82436_/Q _78330_/A sky130_fd_sc_hd__dfxtp_4
XPHY_405 sky130_fd_sc_hd__decap_3
X_55352_ _55352_/A _83753_/Q _55352_/C _55445_/C sky130_fd_sc_hd__nand3_4
X_67338_ _67266_/A _67338_/B _67338_/X sky130_fd_sc_hd__and2_4
X_86172_ _85566_/CLK _86172_/D _86172_/Q sky130_fd_sc_hd__dfxtp_4
X_52564_ _65360_/B _52549_/X _52563_/Y _52564_/Y sky130_fd_sc_hd__o21ai_4
XPHY_416 sky130_fd_sc_hd__decap_3
X_83384_ _83415_/CLK _71767_/X _83384_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_427 sky130_fd_sc_hd__decap_3
X_80596_ _80596_/A _80596_/B _80598_/B sky130_fd_sc_hd__or2_4
XPHY_438 sky130_fd_sc_hd__decap_3
X_54303_ _54312_/A _54325_/B _54312_/C _46680_/Y _54303_/X sky130_fd_sc_hd__and4_4
XPHY_449 sky130_fd_sc_hd__decap_3
X_85123_ _85134_/CLK _85123_/D _56920_/B sky130_fd_sc_hd__dfxtp_4
X_51515_ _85996_/Q _51511_/X _51514_/Y _51515_/Y sky130_fd_sc_hd__o21ai_4
X_58071_ _86631_/Q _58136_/B _58071_/Y sky130_fd_sc_hd__nor2_4
X_82335_ _82335_/CLK _77214_/B _82335_/Q sky130_fd_sc_hd__dfxtp_4
X_55283_ _82983_/Q _55272_/X _55140_/X _55282_/Y _56868_/B sky130_fd_sc_hd__a211o_4
X_67269_ _66910_/A _67269_/X sky130_fd_sc_hd__buf_2
X_52495_ _65000_/B _52422_/X _52494_/Y _52495_/Y sky130_fd_sc_hd__o21ai_4
X_57022_ _45719_/Y _56952_/X _57021_/Y _57022_/Y sky130_fd_sc_hd__o21ai_4
X_69008_ _68987_/A _69008_/B _69008_/X sky130_fd_sc_hd__and2_4
X_54234_ _54230_/A _53067_/B _54234_/Y sky130_fd_sc_hd__nand2_4
X_85054_ _85152_/CLK _85054_/D _45444_/A sky130_fd_sc_hd__dfxtp_4
X_51446_ _86008_/Q _51429_/X _51445_/Y _51446_/Y sky130_fd_sc_hd__o21ai_4
X_82266_ _83514_/CLK _82266_/D _82266_/Q sky130_fd_sc_hd__dfxtp_4
X_70280_ _70280_/A _70160_/X _70162_/X _70164_/X _70280_/Y sky130_fd_sc_hd__nand4_4
X_84005_ _81746_/CLK _84005_/D _82653_/D sky130_fd_sc_hd__dfxtp_4
X_81217_ _82284_/CLK _74890_/X _46239_/A sky130_fd_sc_hd__dfxtp_4
X_54165_ _54160_/A _54186_/B _54146_/X _52997_/D _54165_/X sky130_fd_sc_hd__and4_4
X_51377_ _51375_/Y _51366_/X _51376_/X _86022_/D sky130_fd_sc_hd__a21oi_4
X_82197_ _84766_/CLK _82197_/D _82389_/D sky130_fd_sc_hd__dfxtp_4
X_41130_ _41129_/Y _41130_/X sky130_fd_sc_hd__buf_2
X_53116_ _85694_/Q _53093_/X _53115_/Y _53116_/Y sky130_fd_sc_hd__o21ai_4
X_50328_ _50240_/A _50328_/B _50328_/Y sky130_fd_sc_hd__nand2_4
X_81148_ _82327_/CLK _75042_/A _81148_/Q sky130_fd_sc_hd__dfxtp_4
X_54096_ _54094_/Y _53437_/X _54095_/X _85505_/D sky130_fd_sc_hd__a21oi_4
X_58973_ _58973_/A _58973_/B _58973_/Y sky130_fd_sc_hd__nand2_4
X_41061_ _41061_/A _41061_/X sky130_fd_sc_hd__buf_2
X_53047_ _85707_/Q _53038_/X _53046_/Y _53047_/Y sky130_fd_sc_hd__o21ai_4
X_57924_ _57884_/X _85491_/Q _57923_/X _57924_/X sky130_fd_sc_hd__o21a_4
X_50259_ _50253_/Y _50227_/X _50258_/Y _50259_/Y sky130_fd_sc_hd__a21boi_4
X_73970_ _73949_/A _66153_/B _73970_/X sky130_fd_sc_hd__and2_4
X_85956_ _85471_/CLK _85956_/D _85956_/Q sky130_fd_sc_hd__dfxtp_4
X_81079_ _81121_/CLK _81111_/Q _75381_/B sky130_fd_sc_hd__dfxtp_4
X_72921_ _72722_/X _72921_/X sky130_fd_sc_hd__buf_2
X_84907_ _84903_/CLK _84907_/D _64544_/C sky130_fd_sc_hd__dfxtp_4
X_57855_ _57851_/Y _57854_/Y _57829_/X _57855_/X sky130_fd_sc_hd__a21o_4
X_85887_ _85888_/CLK _85887_/D _65451_/B sky130_fd_sc_hd__dfxtp_4
X_44820_ _43014_/Y _46001_/A sky130_fd_sc_hd__buf_2
X_56806_ _44242_/C _85131_/Q _56805_/X _56806_/Y sky130_fd_sc_hd__a21oi_4
X_75640_ _75640_/A _75616_/A _75641_/B sky130_fd_sc_hd__nor2_4
X_87626_ _87883_/CLK _87626_/D _66795_/B sky130_fd_sc_hd__dfxtp_4
X_72852_ _73186_/A _72852_/X sky130_fd_sc_hd__buf_2
X_84838_ _84838_/CLK _84838_/D _84838_/Q sky130_fd_sc_hd__dfxtp_4
X_57786_ _57952_/A _86333_/Q _57786_/Y sky130_fd_sc_hd__nor2_4
X_54998_ _54253_/A _54998_/X sky130_fd_sc_hd__buf_2
X_71803_ _70500_/D _70830_/B _71804_/A sky130_fd_sc_hd__nor2_4
X_59525_ _59544_/A _59571_/C _59741_/C _59890_/B _60385_/A sky130_fd_sc_hd__and4_4
X_44751_ _41287_/Y _44665_/X _86975_/Q _44666_/X _86975_/D sky130_fd_sc_hd__a2bb2o_4
X_56737_ _56700_/Y _56737_/X sky130_fd_sc_hd__buf_2
X_75571_ _75571_/A _75571_/B _80962_/D sky130_fd_sc_hd__xor2_4
X_87557_ _87814_/CLK _43151_/Y _73126_/A sky130_fd_sc_hd__dfxtp_4
X_41963_ _41963_/A _41963_/Y sky130_fd_sc_hd__inv_2
X_53949_ _53949_/A _53949_/B _53949_/Y sky130_fd_sc_hd__nand2_4
X_72783_ _72780_/X _72782_/X _72735_/X _72783_/X sky130_fd_sc_hd__a21o_4
X_84769_ _86361_/CLK _84769_/D _84769_/Q sky130_fd_sc_hd__dfxtp_4
X_77310_ _77310_/A _77311_/A sky130_fd_sc_hd__inv_2
X_43702_ _43701_/X _87303_/D sky130_fd_sc_hd__inv_2
X_74522_ _70611_/X _74531_/D sky130_fd_sc_hd__buf_2
X_86508_ _86498_/CLK _86508_/D _73310_/B sky130_fd_sc_hd__dfxtp_4
X_40914_ _40913_/X _40914_/X sky130_fd_sc_hd__buf_2
X_47470_ _47444_/A _53067_/B _47470_/Y sky130_fd_sc_hd__nand2_4
X_71734_ _58246_/Y _71711_/Y _71733_/Y _71734_/Y sky130_fd_sc_hd__o21ai_4
X_59456_ _59456_/A _59456_/Y sky130_fd_sc_hd__inv_2
X_78290_ _82590_/Q _78290_/B _78290_/Y sky130_fd_sc_hd__nand2_4
X_56668_ _55489_/B _56553_/Y _56647_/X _56667_/Y _85138_/D sky130_fd_sc_hd__a2bb2o_4
X_44682_ _44679_/X _44680_/X _40610_/X _87002_/Q _44681_/X _44682_/Y
+ sky130_fd_sc_hd__o32ai_4
X_87488_ _87758_/CLK _87488_/D _87488_/Q sky130_fd_sc_hd__dfxtp_4
X_41894_ _43047_/A _41894_/X sky130_fd_sc_hd__buf_2
X_46421_ _46421_/A _50799_/B _46421_/Y sky130_fd_sc_hd__nand2_4
X_58407_ _84856_/Q _58409_/A sky130_fd_sc_hd__inv_2
X_77241_ _77241_/A _77241_/Y sky130_fd_sc_hd__inv_2
X_43633_ _51337_/A _47834_/A sky130_fd_sc_hd__buf_2
X_55619_ _55619_/A _55689_/A sky130_fd_sc_hd__buf_2
X_74453_ _74453_/A _74478_/B sky130_fd_sc_hd__buf_2
X_86439_ _86154_/CLK _86439_/D _65289_/B sky130_fd_sc_hd__dfxtp_4
X_40845_ _40845_/A _40845_/X sky130_fd_sc_hd__buf_2
X_71665_ _58526_/Y _71649_/A _71664_/Y _83419_/D sky130_fd_sc_hd__o21ai_4
X_59387_ _63103_/A _59388_/A sky130_fd_sc_hd__buf_2
X_56599_ _56556_/Y _55570_/D _73078_/A _56598_/Y _56600_/A sky130_fd_sc_hd__a211o_4
Xclkbuf_10_340_0_CLK clkbuf_9_170_0_CLK/X _85643_/CLK sky130_fd_sc_hd__clkbuf_1
X_49140_ _49140_/A _49140_/B _50693_/B sky130_fd_sc_hd__nor2_4
X_73404_ _73355_/X _85576_/Q _73284_/X _73403_/X _73404_/X sky130_fd_sc_hd__a211o_4
X_46352_ _51278_/B _53983_/B sky130_fd_sc_hd__buf_2
X_70616_ _70588_/A _70620_/B sky130_fd_sc_hd__buf_2
X_58338_ _58338_/A _58338_/Y sky130_fd_sc_hd__inv_2
X_77172_ _77172_/A _77172_/B _77177_/A sky130_fd_sc_hd__nor2_4
X_43564_ _43557_/X _43563_/X _40491_/X _87359_/Q _43549_/X _43564_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74384_ _83077_/Q _72090_/X _74383_/Y _74384_/Y sky130_fd_sc_hd__o21ai_4
X_40776_ _40776_/A _40776_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_970_0_CLK clkbuf_9_485_0_CLK/X _86530_/CLK sky130_fd_sc_hd__clkbuf_1
X_71596_ _71581_/A _83444_/Q _71595_/Y _83444_/D sky130_fd_sc_hd__a21o_4
X_45303_ _45651_/A _45303_/X sky130_fd_sc_hd__buf_2
X_76123_ _76112_/A _76107_/A _76126_/A _76127_/B _76123_/Y sky130_fd_sc_hd__nand4_4
X_42515_ _74071_/A _68910_/B sky130_fd_sc_hd__inv_2
X_88109_ _87070_/CLK _41900_/Y _88109_/Q sky130_fd_sc_hd__dfxtp_4
X_49071_ _49066_/Y _49038_/X _49070_/X _86447_/D sky130_fd_sc_hd__a21oi_4
X_73335_ _73163_/X _83059_/Q _72880_/X _73334_/X _73335_/X sky130_fd_sc_hd__a211o_4
X_46283_ _46326_/A _50744_/B _46283_/Y sky130_fd_sc_hd__nand2_4
X_70547_ DATA_TO_HASH[5] _71857_/A sky130_fd_sc_hd__inv_2
X_58269_ _58253_/X _83444_/Q _58268_/Y _84892_/D sky130_fd_sc_hd__o21a_4
X_43495_ _43518_/A _43495_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_461_0_CLK clkbuf_9_461_0_CLK/A clkbuf_9_461_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_60300_ _60367_/B _60300_/B _60300_/C _60300_/Y sky130_fd_sc_hd__nand3_4
X_48022_ _83543_/Q _48022_/Y sky130_fd_sc_hd__inv_2
X_45234_ _64458_/B _61579_/B sky130_fd_sc_hd__buf_2
X_76054_ _76054_/A _81748_/D _76054_/X sky130_fd_sc_hd__xor2_4
X_42446_ _42446_/A _47872_/A sky130_fd_sc_hd__buf_2
X_61280_ _61286_/A _60593_/B _61079_/A _60509_/Y _61281_/A sky130_fd_sc_hd__nor4_4
X_73266_ _73214_/X _83062_/Q _73238_/X _73265_/X _73266_/X sky130_fd_sc_hd__a211o_4
X_70478_ _70466_/Y _58356_/B _70477_/X _83766_/D sky130_fd_sc_hd__a21o_4
Xclkbuf_10_355_0_CLK clkbuf_9_177_0_CLK/X _86637_/CLK sky130_fd_sc_hd__clkbuf_1
X_75005_ _75001_/Y _75004_/X _75005_/Y sky130_fd_sc_hd__nand2_4
X_60231_ _60078_/X _60299_/A _60300_/B _60229_/Y _60230_/Y _60231_/Y
+ sky130_fd_sc_hd__a41oi_4
X_72217_ _72155_/X _85689_/Q _72156_/X _72217_/X sky130_fd_sc_hd__o21a_4
X_45165_ _56420_/C _45102_/X _45164_/X _45165_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_985_0_CLK clkbuf_9_492_0_CLK/X _83562_/CLK sky130_fd_sc_hd__clkbuf_1
X_42377_ _41782_/X _42374_/X _87894_/Q _42375_/X _87894_/D sky130_fd_sc_hd__a2bb2o_4
X_73197_ _69790_/Y _73104_/B _73194_/X _73196_/Y _73197_/X sky130_fd_sc_hd__a211o_4
X_44116_ _43957_/B _44116_/B _43978_/Y _44117_/A sky130_fd_sc_hd__nor3_4
X_79813_ _79829_/A _79812_/Y _79813_/X sky130_fd_sc_hd__xor2_4
X_41328_ _41327_/Y _41328_/X sky130_fd_sc_hd__buf_2
X_60162_ _60162_/A _60636_/B _59615_/A _61287_/A _60162_/X sky130_fd_sc_hd__and4_4
X_72148_ _59381_/X _85983_/Q _72147_/X _72148_/Y sky130_fd_sc_hd__o21ai_4
X_49973_ _49973_/A _49973_/B _49973_/C _53185_/D _49973_/X sky130_fd_sc_hd__and4_4
X_45096_ _45093_/X _45095_/Y _45049_/X _45096_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_476_0_CLK clkbuf_8_238_0_CLK/X clkbuf_9_476_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_48924_ _48924_/A _48699_/B _48924_/Y sky130_fd_sc_hd__nand2_4
X_44047_ _44046_/X _44047_/X sky130_fd_sc_hd__buf_2
X_79744_ _79740_/X _79743_/Y _79745_/A sky130_fd_sc_hd__xor2_4
X_41259_ _41259_/A _41259_/X sky130_fd_sc_hd__buf_2
X_64970_ _64966_/Y _64939_/X _64969_/X _64970_/X sky130_fd_sc_hd__a21o_4
X_60093_ _84663_/Q _59822_/X _59969_/X _60092_/Y _60093_/X sky130_fd_sc_hd__o22a_4
X_72079_ _72075_/A _72079_/B _72079_/Y sky130_fd_sc_hd__nand2_4
X_76956_ _76956_/A _76955_/Y _76958_/A sky130_fd_sc_hd__nand2_4
X_63921_ _57664_/X _63902_/B _63902_/C _63902_/D _63922_/D sky130_fd_sc_hd__nand4_4
X_75907_ _84505_/Q _75907_/B _75907_/X sky130_fd_sc_hd__xor2_4
X_48855_ _48852_/Y _48840_/X _48854_/X _48855_/Y sky130_fd_sc_hd__a21oi_4
X_79675_ _79667_/A _79666_/Y _79674_/X _79676_/B sky130_fd_sc_hd__o21ai_4
X_76887_ _76888_/A _76888_/C _76888_/B _76901_/A sky130_fd_sc_hd__a21o_4
X_47806_ _47714_/A _47806_/X sky130_fd_sc_hd__buf_2
X_66640_ _66689_/A _87632_/Q _66640_/X sky130_fd_sc_hd__and2_4
X_78626_ _78626_/A _78625_/Y _82775_/D sky130_fd_sc_hd__xor2_4
X_75838_ _80927_/Q _75838_/Y sky130_fd_sc_hd__inv_2
X_63852_ _63749_/A _63853_/B sky130_fd_sc_hd__buf_2
X_48786_ _50469_/A _48770_/X _48786_/C _48786_/X sky130_fd_sc_hd__and3_4
X_45998_ _40468_/Y _45974_/X _86822_/Q _45976_/X _45998_/X sky130_fd_sc_hd__a2bb2o_4
X_62803_ _62667_/X _62848_/C sky130_fd_sc_hd__buf_2
X_47737_ _81227_/Q _55078_/D sky130_fd_sc_hd__inv_2
X_66571_ _69162_/A _66571_/X sky130_fd_sc_hd__buf_2
X_78557_ _78548_/X _78557_/B _78556_/Y _78560_/A sky130_fd_sc_hd__or3_4
Xclkbuf_10_923_0_CLK clkbuf_9_461_0_CLK/X _88337_/CLK sky130_fd_sc_hd__clkbuf_1
X_44949_ _55963_/B _44935_/X _45757_/A _44949_/X sky130_fd_sc_hd__o21a_4
X_63783_ _63779_/X _63736_/X _63780_/Y _63781_/Y _63782_/X _63783_/X
+ sky130_fd_sc_hd__a41o_4
X_75769_ _81096_/Q _80808_/Q _75769_/Y sky130_fd_sc_hd__xnor2_4
X_60995_ _60994_/Y _60995_/Y sky130_fd_sc_hd__inv_2
X_68310_ _68301_/X _67887_/Y _68308_/X _68309_/Y _68310_/X sky130_fd_sc_hd__a211o_4
X_65522_ _65362_/X _85595_/Q _65363_/X _65521_/X _65522_/X sky130_fd_sc_hd__a211o_4
X_77508_ _77508_/A _77508_/Y sky130_fd_sc_hd__inv_2
X_62734_ _62672_/A _62766_/B sky130_fd_sc_hd__buf_2
X_69290_ _69287_/X _69289_/X _69251_/X _69290_/X sky130_fd_sc_hd__a21o_4
X_47668_ _47668_/A _54871_/B sky130_fd_sc_hd__inv_2
X_78488_ _78489_/A _82671_/D _78488_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_9_414_0_CLK clkbuf_9_415_0_CLK/A clkbuf_9_414_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_49407_ _49407_/A _49420_/A sky130_fd_sc_hd__buf_2
X_68241_ _68221_/X _67484_/Y _68228_/X _68240_/Y _68241_/X sky130_fd_sc_hd__a211o_4
X_46619_ _46619_/A _52580_/D sky130_fd_sc_hd__buf_2
X_65453_ _65118_/A _65453_/X sky130_fd_sc_hd__buf_2
X_77439_ _77403_/B _77434_/Y _77438_/Y _77439_/Y sky130_fd_sc_hd__a21oi_4
X_62665_ _62910_/A _62847_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_308_0_CLK clkbuf_9_154_0_CLK/X _83431_/CLK sky130_fd_sc_hd__clkbuf_1
X_47599_ _47574_/A _53141_/B _47599_/Y sky130_fd_sc_hd__nand2_4
X_64404_ _64380_/X _84865_/Q _64381_/X _64404_/Y sky130_fd_sc_hd__nand3_4
X_49338_ _49327_/X _54071_/B _49338_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_938_0_CLK clkbuf_9_469_0_CLK/X _87813_/CLK sky130_fd_sc_hd__clkbuf_1
X_61616_ _61614_/X _61576_/X _61615_/Y _61616_/Y sky130_fd_sc_hd__a21oi_4
X_80450_ _80429_/B _80446_/X _80449_/Y _80451_/B sky130_fd_sc_hd__a21oi_4
X_68172_ _82061_/D _68160_/X _68171_/X _68172_/X sky130_fd_sc_hd__a21bo_4
X_65384_ _65184_/A _65384_/B _65384_/X sky130_fd_sc_hd__and2_4
X_62596_ _62269_/X _58201_/X _62618_/C _62608_/D _62596_/X sky130_fd_sc_hd__and4_4
X_67123_ _67023_/A _67123_/B _67123_/X sky130_fd_sc_hd__and2_4
X_79109_ _79109_/A _79109_/B _79107_/A _79110_/B sky130_fd_sc_hd__nand3_4
X_64335_ _64295_/A _64307_/B _64335_/C _64335_/X sky130_fd_sc_hd__and3_4
Xclkbuf_9_429_0_CLK clkbuf_9_429_0_CLK/A clkbuf_9_429_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_61547_ _61545_/X _61517_/X _61546_/Y _61547_/Y sky130_fd_sc_hd__a21oi_4
X_49269_ _49261_/A _46396_/B _49269_/Y sky130_fd_sc_hd__nand2_4
X_80381_ _80394_/A _80394_/B _80404_/B sky130_fd_sc_hd__xor2_4
X_51300_ _51296_/A _46396_/B _51300_/Y sky130_fd_sc_hd__nand2_4
X_82120_ _82485_/CLK _82120_/D _82108_/D sky130_fd_sc_hd__dfxtp_4
X_67054_ _67051_/X _67053_/X _67054_/Y sky130_fd_sc_hd__nand2_4
X_52280_ _52319_/A _52280_/X sky130_fd_sc_hd__buf_2
X_64266_ _59463_/Y _64249_/X _64265_/Y _64266_/Y sky130_fd_sc_hd__o21ai_4
X_61478_ _61473_/X _61455_/X _61477_/Y _84478_/D sky130_fd_sc_hd__a21oi_4
X_66005_ _66001_/Y _65987_/X _66004_/X _66005_/X sky130_fd_sc_hd__a21o_4
X_51231_ _51220_/A _51230_/X _51225_/C _47218_/D _51231_/X sky130_fd_sc_hd__and4_4
X_63217_ _63216_/X _63217_/B _63241_/C _63181_/X _63217_/X sky130_fd_sc_hd__and4_4
X_82051_ _82053_/CLK _84011_/Q _82051_/Q sky130_fd_sc_hd__dfxtp_4
X_60429_ _60472_/A _60433_/A sky130_fd_sc_hd__buf_2
X_64197_ _64193_/X _63741_/X _64194_/Y _64195_/Y _64196_/Y _64197_/X
+ sky130_fd_sc_hd__a41o_4
X_81002_ _84197_/CLK _84210_/Q _81002_/Q sky130_fd_sc_hd__dfxtp_4
X_51162_ _51167_/A _52855_/B _51162_/Y sky130_fd_sc_hd__nand2_4
X_63148_ _63142_/Y _63143_/X _63146_/X _63147_/X _63125_/X _63148_/Y
+ sky130_fd_sc_hd__o41ai_4
X_50113_ _50113_/A _50113_/X sky130_fd_sc_hd__buf_2
X_85810_ _86030_/CLK _52499_/Y _65000_/B sky130_fd_sc_hd__dfxtp_4
X_51093_ _51039_/A _51093_/X sky130_fd_sc_hd__buf_2
X_55970_ _56381_/C _55689_/A _55611_/X _55969_/X _55970_/X sky130_fd_sc_hd__a211o_4
X_67956_ _87449_/Q _67953_/X _67954_/X _67955_/X _67956_/X sky130_fd_sc_hd__a211o_4
X_63079_ _63041_/A _63079_/B _63079_/C _63066_/D _63079_/X sky130_fd_sc_hd__and4_4
X_86790_ _86796_/CLK _86790_/D _66962_/B sky130_fd_sc_hd__dfxtp_4
X_50044_ _51012_/A _50929_/A sky130_fd_sc_hd__buf_2
X_54921_ _85353_/Q _54918_/X _54920_/Y _54921_/Y sky130_fd_sc_hd__o21ai_4
X_66907_ _66956_/A _88197_/Q _66907_/X sky130_fd_sc_hd__and2_4
X_85741_ _85741_/CLK _52862_/Y _85741_/Q sky130_fd_sc_hd__dfxtp_4
X_82953_ _82965_/CLK _82953_/D _82953_/Q sky130_fd_sc_hd__dfxtp_4
X_67887_ _67887_/A _67887_/B _67887_/Y sky130_fd_sc_hd__nand2_4
X_57640_ _71970_/A _50381_/B _57640_/Y sky130_fd_sc_hd__nand2_4
X_81904_ _81990_/CLK _77441_/X _82280_/D sky130_fd_sc_hd__dfxtp_4
X_69626_ _69626_/A _69865_/A sky130_fd_sc_hd__buf_2
X_54852_ _54857_/A _54857_/B _54857_/C _53159_/D _54852_/X sky130_fd_sc_hd__and4_4
X_66838_ _66795_/A _87624_/Q _66838_/X sky130_fd_sc_hd__and2_4
X_85672_ _84815_/CLK _53235_/Y _85672_/Q sky130_fd_sc_hd__dfxtp_4
X_82884_ _88267_/CLK _78095_/Y _82884_/Q sky130_fd_sc_hd__dfxtp_4
X_87411_ _83987_/CLK _87411_/D _87411_/Q sky130_fd_sc_hd__dfxtp_4
X_53803_ _53786_/A _48920_/Y _53803_/Y sky130_fd_sc_hd__nand2_4
X_84623_ _84623_/CLK _60358_/Y _79605_/A sky130_fd_sc_hd__dfxtp_4
X_57571_ _71959_/A _57619_/B sky130_fd_sc_hd__buf_2
X_69557_ _69554_/X _69556_/X _64629_/A _69557_/X sky130_fd_sc_hd__a21o_4
X_81835_ _82220_/CLK _81867_/Q _77353_/A sky130_fd_sc_hd__dfxtp_4
X_88391_ _88394_/CLK _40442_/Y _88391_/Q sky130_fd_sc_hd__dfxtp_4
X_54783_ _54034_/A _54892_/A sky130_fd_sc_hd__buf_2
X_66769_ _66769_/A _88203_/Q _66769_/X sky130_fd_sc_hd__and2_4
X_51995_ _52322_/A _52185_/A sky130_fd_sc_hd__buf_2
X_59310_ _59260_/X _85416_/Q _59309_/X _59310_/Y sky130_fd_sc_hd__o21ai_4
X_56522_ _46187_/A _56533_/B sky130_fd_sc_hd__buf_2
X_68508_ _46210_/A _68993_/A sky130_fd_sc_hd__buf_2
X_87342_ _86988_/CLK _43616_/Y _43614_/A sky130_fd_sc_hd__dfxtp_4
X_53734_ _50511_/A _53748_/B _53734_/C _53734_/X sky130_fd_sc_hd__and3_4
X_84554_ _84375_/CLK _84554_/D _78049_/A sky130_fd_sc_hd__dfxtp_4
X_50946_ _50946_/A _50973_/A sky130_fd_sc_hd__buf_2
X_81766_ _82642_/CLK _76003_/X _81766_/Q sky130_fd_sc_hd__dfxtp_4
X_69488_ _69484_/X _69487_/X _69389_/X _69488_/Y sky130_fd_sc_hd__a21oi_4
X_59241_ _58868_/A _59241_/X sky130_fd_sc_hd__buf_2
X_83505_ _84223_/CLK _83505_/D _83505_/Q sky130_fd_sc_hd__dfxtp_4
X_56453_ _56164_/X _56372_/X _56452_/Y _56453_/Y sky130_fd_sc_hd__o21ai_4
X_80717_ _81084_/CLK _75903_/X _80685_/D sky130_fd_sc_hd__dfxtp_4
X_68439_ _69088_/A _68439_/X sky130_fd_sc_hd__buf_2
X_87273_ _87273_/CLK _43773_/X _69274_/B sky130_fd_sc_hd__dfxtp_4
X_53665_ _50460_/A _53733_/A sky130_fd_sc_hd__buf_2
X_84485_ _82272_/CLK _61385_/Y _79153_/B sky130_fd_sc_hd__dfxtp_4
X_50877_ _50875_/Y _50243_/X _50876_/Y _50877_/Y sky130_fd_sc_hd__a21boi_4
X_81697_ _81697_/CLK _80261_/Y _81697_/Q sky130_fd_sc_hd__dfxtp_4
X_55404_ _55188_/X _55193_/X _55405_/A sky130_fd_sc_hd__and2_4
X_86224_ _83544_/CLK _86224_/D _86224_/Q sky130_fd_sc_hd__dfxtp_4
X_40630_ _48631_/A _40817_/A sky130_fd_sc_hd__buf_2
X_52616_ _52624_/A _54309_/B _52616_/Y sky130_fd_sc_hd__nand2_4
X_59172_ _59117_/A _86355_/Q _59172_/Y sky130_fd_sc_hd__nor2_4
X_71450_ _70676_/A _71626_/C _71450_/C _71450_/Y sky130_fd_sc_hd__nor3_4
X_83436_ _83491_/CLK _83436_/D _83436_/Q sky130_fd_sc_hd__dfxtp_4
X_56384_ _44207_/A _56436_/A sky130_fd_sc_hd__buf_2
XPHY_202 sky130_fd_sc_hd__decap_3
X_80648_ _74793_/X _74712_/Y DATA_FROM_HASH[5] sky130_fd_sc_hd__ebufn_2
X_53596_ _53594_/Y _53574_/X _53595_/Y _85606_/D sky130_fd_sc_hd__a21boi_4
XPHY_213 sky130_fd_sc_hd__decap_3
XPHY_224 sky130_fd_sc_hd__decap_3
X_58123_ _65034_/A _58124_/A sky130_fd_sc_hd__buf_2
X_70401_ _71005_/A _74531_/A sky130_fd_sc_hd__buf_2
XPHY_235 sky130_fd_sc_hd__decap_3
X_55335_ _56989_/B _44060_/X _44046_/X _55334_/Y _55335_/X sky130_fd_sc_hd__a211o_4
X_86155_ _86155_/CLK _86155_/D _86155_/Q sky130_fd_sc_hd__dfxtp_4
X_40561_ _42447_/C _41869_/B sky130_fd_sc_hd__inv_2
XPHY_246 sky130_fd_sc_hd__decap_3
X_52547_ _52542_/X _50854_/B _52547_/Y sky130_fd_sc_hd__nand2_4
X_83367_ _83367_/CLK _83367_/D _83367_/Q sky130_fd_sc_hd__dfxtp_4
X_71381_ _70676_/A _71377_/B _71377_/C _71381_/Y sky130_fd_sc_hd__nor3_4
XPHY_257 sky130_fd_sc_hd__decap_3
X_80579_ _80579_/A _80579_/B _80580_/B sky130_fd_sc_hd__xor2_4
XPHY_268 sky130_fd_sc_hd__decap_3
X_42300_ _42300_/A _42300_/Y sky130_fd_sc_hd__inv_2
X_73120_ _74428_/B _73120_/B _73120_/X sky130_fd_sc_hd__xor2_4
X_85106_ _85074_/CLK _85106_/D _85106_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_279 sky130_fd_sc_hd__decap_3
X_58054_ _57991_/A _86313_/Q _58054_/Y sky130_fd_sc_hd__nor2_4
X_70332_ _70134_/X _70332_/X sky130_fd_sc_hd__buf_2
X_82318_ _82284_/CLK _77089_/B _82318_/Q sky130_fd_sc_hd__dfxtp_4
X_43280_ _43260_/X _43269_/X _41139_/X _87502_/Q _43273_/X _43280_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55266_ _55265_/Y _55288_/C sky130_fd_sc_hd__inv_2
X_86086_ _85767_/CLK _86086_/D _86086_/Q sky130_fd_sc_hd__dfxtp_4
X_40492_ _44736_/A _40492_/X sky130_fd_sc_hd__buf_2
X_52478_ _52468_/A _52478_/B _52478_/Y sky130_fd_sc_hd__nand2_4
X_83298_ _85554_/CLK _72035_/Y _83298_/Q sky130_fd_sc_hd__dfxtp_4
X_57005_ _57427_/A _56750_/Y _56982_/X _57005_/Y sky130_fd_sc_hd__a21oi_4
X_42231_ _42204_/X _42231_/X sky130_fd_sc_hd__buf_2
X_54217_ _54217_/A _54237_/B sky130_fd_sc_hd__buf_2
X_73051_ _83167_/Q _72943_/X _73050_/Y _83167_/D sky130_fd_sc_hd__a21o_4
X_85037_ _85037_/CLK _85037_/D _85037_/Q sky130_fd_sc_hd__dfxtp_4
X_51429_ _51539_/A _51429_/X sky130_fd_sc_hd__buf_2
X_70263_ _70247_/X _70267_/B sky130_fd_sc_hd__buf_2
X_82249_ _82820_/CLK _80375_/X _82249_/Q sky130_fd_sc_hd__dfxtp_4
X_55197_ _55164_/X _55298_/A _55400_/A _55201_/A sky130_fd_sc_hd__nand3_4
X_72002_ _57563_/X _72040_/A sky130_fd_sc_hd__buf_2
X_42162_ _42162_/A _42162_/X sky130_fd_sc_hd__buf_2
X_54148_ _54143_/Y _54144_/X _54147_/X _85496_/D sky130_fd_sc_hd__a21oi_4
X_70194_ _70192_/Y _70157_/X _70193_/Y _83842_/D sky130_fd_sc_hd__o21ai_4
X_41113_ _40946_/A _41113_/X sky130_fd_sc_hd__buf_2
X_76810_ _76810_/A _76812_/A sky130_fd_sc_hd__inv_2
X_46970_ _59057_/A _46955_/X _46969_/Y _46970_/Y sky130_fd_sc_hd__o21ai_4
X_58956_ _58599_/A _58956_/X sky130_fd_sc_hd__buf_2
X_54079_ _53801_/B _54079_/B _54079_/Y sky130_fd_sc_hd__nand2_4
X_42093_ _42093_/A _42093_/Y sky130_fd_sc_hd__inv_2
X_77790_ _77796_/A _77783_/Y _77789_/Y _77791_/B sky130_fd_sc_hd__o21ai_4
X_86988_ _86988_/CLK _86988_/D _44719_/A sky130_fd_sc_hd__dfxtp_4
X_57907_ _57838_/X _86005_/Q _57906_/X _57907_/Y sky130_fd_sc_hd__o21ai_4
X_45921_ _64565_/A _64902_/A sky130_fd_sc_hd__buf_2
X_41044_ _41042_/X _82286_/Q _41043_/X _41045_/A sky130_fd_sc_hd__o21a_4
X_76741_ _76727_/Y _76728_/Y _76714_/A _81354_/D _76741_/X sky130_fd_sc_hd__a2bb2o_4
X_73953_ _73950_/X _73952_/X _73857_/X _73956_/A sky130_fd_sc_hd__a21o_4
X_85939_ _86100_/CLK _85939_/D _85939_/Q sky130_fd_sc_hd__dfxtp_4
X_58887_ _58887_/A _58873_/B _58887_/Y sky130_fd_sc_hd__nor2_4
X_48640_ _48661_/A _48843_/B _48640_/Y sky130_fd_sc_hd__nand2_4
X_72904_ _72898_/X _72904_/B _72904_/Y sky130_fd_sc_hd__nand2_4
X_79460_ _79438_/A _79438_/B _79449_/A _79448_/Y _79460_/X sky130_fd_sc_hd__o22a_4
X_45852_ _45845_/X _45849_/Y _45851_/Y _45852_/Y sky130_fd_sc_hd__a21oi_4
X_57838_ _58618_/A _57838_/X sky130_fd_sc_hd__buf_2
X_76672_ _76668_/X _76672_/B _76669_/Y _76672_/Y sky130_fd_sc_hd__nand3_4
X_73884_ _73786_/X _84980_/Q _73859_/X _73883_/X _73884_/X sky130_fd_sc_hd__a211o_4
X_78411_ _78411_/A _78411_/B _78409_/Y _78412_/A sky130_fd_sc_hd__nand3_4
X_44803_ _44803_/A _46258_/A sky130_fd_sc_hd__buf_2
X_75623_ _80775_/D _75621_/A _75623_/X sky130_fd_sc_hd__and2_4
X_87609_ _82899_/CLK _87609_/D _87609_/Q sky130_fd_sc_hd__dfxtp_4
X_48571_ _48571_/A _48572_/A sky130_fd_sc_hd__inv_2
X_72835_ _44522_/Y _72775_/X _72834_/Y _72835_/X sky130_fd_sc_hd__a21o_4
X_79391_ _79384_/X _79391_/B _79391_/Y sky130_fd_sc_hd__nand2_4
X_57769_ _64923_/A _57770_/A sky130_fd_sc_hd__buf_2
X_45783_ _57340_/B _44933_/X _45782_/X _45783_/Y sky130_fd_sc_hd__o21ai_4
X_42995_ _42951_/A _42995_/X sky130_fd_sc_hd__buf_2
X_47522_ _47513_/A _47549_/B _47519_/X _53099_/D _47522_/X sky130_fd_sc_hd__and4_4
X_59508_ _57689_/A _59508_/X sky130_fd_sc_hd__buf_2
X_78342_ _78344_/A _82661_/D _78342_/Y sky130_fd_sc_hd__nor2_4
X_44734_ _43047_/A _50731_/B sky130_fd_sc_hd__buf_2
X_75554_ _80704_/Q _75554_/B _75555_/A sky130_fd_sc_hd__nand2_4
X_41946_ _41945_/Y _41946_/Y sky130_fd_sc_hd__inv_2
X_60780_ _63371_/A _60780_/X sky130_fd_sc_hd__buf_2
X_72766_ _74140_/A _72766_/X sky130_fd_sc_hd__buf_2
X_74505_ _74505_/A _74509_/B _74501_/C _74505_/X sky130_fd_sc_hd__and3_4
X_47453_ _86633_/Q _47429_/X _47452_/Y _47453_/Y sky130_fd_sc_hd__o21ai_4
X_71717_ _71712_/Y _83401_/Q _71716_/X _83401_/D sky130_fd_sc_hd__a21o_4
X_59439_ _84732_/Q _59439_/Y sky130_fd_sc_hd__inv_2
X_78273_ _78273_/A _78273_/B _78284_/B sky130_fd_sc_hd__nand2_4
X_44665_ _44618_/A _44665_/X sky130_fd_sc_hd__buf_2
X_75485_ _75465_/Y _75470_/Y _75507_/A _75485_/X sky130_fd_sc_hd__o21a_4
X_41877_ _41877_/A _41878_/A sky130_fd_sc_hd__buf_2
X_72697_ _72697_/A _72697_/B _56832_/X _72697_/Y sky130_fd_sc_hd__nand3_4
X_46404_ _46349_/A _46459_/B sky130_fd_sc_hd__buf_2
X_77224_ _82017_/Q _82305_/D _77227_/C sky130_fd_sc_hd__xnor2_4
X_43616_ _43616_/A _43616_/Y sky130_fd_sc_hd__inv_2
X_62450_ _61522_/X _62492_/B _62449_/X _62404_/X _62450_/Y sky130_fd_sc_hd__nand4_4
X_74436_ _74434_/Y _74430_/X _74435_/X _74436_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_61_0_CLK clkbuf_9_30_0_CLK/X _84998_/CLK sky130_fd_sc_hd__clkbuf_1
X_40828_ _40828_/A _40828_/Y sky130_fd_sc_hd__inv_2
X_47384_ _47525_/A _47404_/A sky130_fd_sc_hd__buf_2
X_71648_ _71507_/A _70854_/A _71528_/X _71649_/A sky130_fd_sc_hd__nor3_4
X_44596_ _44533_/A _44596_/X sky130_fd_sc_hd__buf_2
X_61401_ _61400_/X _61429_/C sky130_fd_sc_hd__buf_2
X_49123_ _49118_/Y _49086_/X _49122_/X _86442_/D sky130_fd_sc_hd__a21oi_4
X_46335_ _46326_/A _49241_/B _46335_/Y sky130_fd_sc_hd__nand2_4
X_77155_ _77146_/B _77155_/B _77159_/A sky130_fd_sc_hd__nand2_4
X_43547_ _43542_/X _43546_/X _40446_/X _87366_/Q _43528_/X _43548_/A
+ sky130_fd_sc_hd__o32ai_4
X_62381_ _62371_/X _62378_/Y _62380_/X _84742_/Q _62367_/X _62381_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74367_ _74364_/Y _72059_/X _74366_/X _83081_/D sky130_fd_sc_hd__a21oi_4
X_40759_ _40836_/A _40759_/X sky130_fd_sc_hd__buf_2
X_71579_ _71602_/C _71189_/B _71580_/A sky130_fd_sc_hd__nor2_4
Xclkbuf_7_106_0_CLK clkbuf_6_53_0_CLK/X clkbuf_8_213_0_CLK/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_294_0_CLK clkbuf_9_147_0_CLK/X _84263_/CLK sky130_fd_sc_hd__clkbuf_1
X_64120_ _63655_/B _64091_/B _64178_/C _64091_/D _64120_/Y sky130_fd_sc_hd__nand4_4
X_76106_ _76103_/A _76099_/A _76107_/A sky130_fd_sc_hd__and2_4
X_49054_ _49054_/A _49055_/A sky130_fd_sc_hd__inv_2
X_61332_ _61305_/A _61330_/X _61377_/C _61332_/Y sky130_fd_sc_hd__nand3_4
X_73318_ _73193_/A _73318_/X sky130_fd_sc_hd__buf_2
X_46266_ _46262_/X _81216_/Q _46265_/X _46267_/A sky130_fd_sc_hd__o21ai_4
X_77086_ _77085_/Y _77086_/B _77087_/B sky130_fd_sc_hd__and2_4
X_43478_ _41681_/X _43465_/X _87402_/Q _43467_/X _87402_/D sky130_fd_sc_hd__a2bb2o_4
X_74298_ _70280_/A _74288_/X _74297_/Y _74298_/X sky130_fd_sc_hd__a21bo_4
X_48005_ _66143_/B _47998_/X _48004_/Y _48005_/Y sky130_fd_sc_hd__o21ai_4
X_45217_ _45214_/X _45216_/Y _45200_/X _45217_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_76_0_CLK clkbuf_9_38_0_CLK/X _84407_/CLK sky130_fd_sc_hd__clkbuf_1
X_64051_ _63972_/A _64150_/C sky130_fd_sc_hd__buf_2
X_76037_ _76037_/A _76028_/B _76038_/B sky130_fd_sc_hd__and2_4
X_42429_ _42429_/A _42574_/A sky130_fd_sc_hd__buf_2
X_61263_ _59716_/A _61176_/Y _59710_/Y _61260_/X _61262_/Y _84495_/D
+ sky130_fd_sc_hd__a41oi_4
X_73249_ _72881_/A _73250_/A sky130_fd_sc_hd__buf_2
X_46197_ _57701_/A _66002_/A sky130_fd_sc_hd__inv_2
Xclkbuf_8_222_0_CLK clkbuf_8_223_0_CLK/A clkbuf_9_444_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_63002_ _63281_/B _60438_/A _60417_/A _60508_/A _60392_/C _63002_/X
+ sky130_fd_sc_hd__o41a_4
X_60214_ _60244_/A _60214_/B _60214_/C _60214_/Y sky130_fd_sc_hd__nor3_4
X_45148_ _85233_/Q _45131_/X _45087_/X _45148_/X sky130_fd_sc_hd__o21a_4
X_61194_ _59789_/A _61194_/X sky130_fd_sc_hd__buf_2
X_67810_ _67739_/X _67810_/B _67810_/X sky130_fd_sc_hd__and2_4
X_60145_ _60145_/A _60145_/Y sky130_fd_sc_hd__inv_2
X_49956_ _72277_/B _49934_/X _49955_/Y _49956_/Y sky130_fd_sc_hd__o21ai_4
X_45079_ _45153_/A _45079_/X sky130_fd_sc_hd__buf_2
X_68790_ _68542_/X _68790_/B _68790_/X sky130_fd_sc_hd__and2_4
X_77988_ _78010_/A _77993_/A sky130_fd_sc_hd__inv_2
X_48907_ _52275_/B _71970_/B sky130_fd_sc_hd__buf_2
X_79727_ _79711_/X _79714_/Y _79726_/X _79727_/X sky130_fd_sc_hd__a21o_4
X_67741_ _87394_/Q _67717_/X _67718_/X _67740_/X _67741_/X sky130_fd_sc_hd__a211o_4
X_64953_ _64953_/A _64953_/B _64953_/Y sky130_fd_sc_hd__nand2_4
X_76939_ _76939_/A _76938_/B _76939_/X sky130_fd_sc_hd__or2_4
X_60076_ _60075_/Y _84666_/D sky130_fd_sc_hd__inv_2
X_49887_ _72116_/B _49880_/X _49886_/Y _49887_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_8_237_0_CLK clkbuf_8_237_0_CLK/A clkbuf_9_475_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_232_0_CLK clkbuf_9_116_0_CLK/X _81087_/CLK sky130_fd_sc_hd__clkbuf_1
X_63904_ _60909_/X _63905_/C sky130_fd_sc_hd__buf_2
X_48838_ _48851_/A _48628_/B _48838_/Y sky130_fd_sc_hd__nand2_4
X_67672_ _67696_/A _67672_/B _67672_/X sky130_fd_sc_hd__and2_4
X_79658_ _79658_/A _79658_/B _79668_/B sky130_fd_sc_hd__xor2_4
X_64884_ _64828_/X _85559_/Q _64829_/X _64883_/X _64884_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_862_0_CLK clkbuf_9_431_0_CLK/X _86424_/CLK sky130_fd_sc_hd__clkbuf_1
X_69411_ _69305_/A _69411_/B _69411_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_14_0_CLK clkbuf_9_7_0_CLK/X _83001_/CLK sky130_fd_sc_hd__clkbuf_1
X_66623_ _66620_/X _66622_/X _66623_/Y sky130_fd_sc_hd__nand2_4
X_78609_ _78608_/A _82678_/D _78609_/Y sky130_fd_sc_hd__nand2_4
X_63835_ _63832_/X _63833_/X _63834_/Y _63835_/Y sky130_fd_sc_hd__a21oi_4
X_48769_ _86486_/Q _48754_/X _48768_/Y _48769_/Y sky130_fd_sc_hd__o21ai_4
X_79589_ _79594_/B _79588_/Y _79592_/A sky130_fd_sc_hd__nand2_4
Xclkbuf_9_353_0_CLK clkbuf_8_176_0_CLK/X clkbuf_9_353_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_50800_ _86130_/Q _50727_/X _50799_/Y _50800_/Y sky130_fd_sc_hd__o21ai_4
X_81620_ _81620_/CLK _76423_/X _81620_/Q sky130_fd_sc_hd__dfxtp_4
X_69342_ _88036_/Q _69162_/X _69202_/X _69341_/X _69342_/X sky130_fd_sc_hd__a211o_4
X_66554_ _66553_/X _66554_/X sky130_fd_sc_hd__buf_2
X_51780_ _85947_/Q _51763_/X _51779_/Y _51780_/Y sky130_fd_sc_hd__o21ai_4
X_63766_ _63759_/X _63736_/X _63760_/Y _63762_/Y _63765_/X _63766_/X
+ sky130_fd_sc_hd__a41o_4
X_60978_ _60961_/X _60972_/X _60976_/Y _60958_/X _60977_/X _84546_/D
+ sky130_fd_sc_hd__o41a_4
Xclkbuf_10_247_0_CLK clkbuf_9_123_0_CLK/X _84458_/CLK sky130_fd_sc_hd__clkbuf_1
X_65505_ _65387_/A _72911_/B _65505_/X sky130_fd_sc_hd__and2_4
X_50731_ _50731_/A _50731_/B _53944_/C _50731_/Y sky130_fd_sc_hd__nor3_4
X_62717_ _62717_/A _62717_/X sky130_fd_sc_hd__buf_2
X_81551_ _83918_/CLK _76771_/X _76158_/B sky130_fd_sc_hd__dfxtp_4
X_69273_ _69178_/A _69288_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_877_0_CLK clkbuf_9_438_0_CLK/X _86749_/CLK sky130_fd_sc_hd__clkbuf_1
X_66485_ _66445_/A _66514_/B _66484_/Y _66485_/Y sky130_fd_sc_hd__nor3_4
X_63697_ _63697_/A _64534_/C _63458_/A _63697_/X sky130_fd_sc_hd__and3_4
Xclkbuf_10_29_0_CLK clkbuf_9_14_0_CLK/X _85250_/CLK sky130_fd_sc_hd__clkbuf_1
X_80502_ _80502_/A _80501_/Y _82261_/D sky130_fd_sc_hd__xor2_4
X_68224_ _84008_/Q _68220_/X _68223_/X _68224_/X sky130_fd_sc_hd__a21bo_4
X_53450_ _53450_/A _54321_/A sky130_fd_sc_hd__buf_2
X_65436_ _65433_/Y _65347_/X _65435_/X _84201_/D sky130_fd_sc_hd__a21o_4
X_84270_ _84269_/CLK _84270_/D _79950_/B sky130_fd_sc_hd__dfxtp_4
X_50662_ _50627_/X _49073_/X _50662_/Y sky130_fd_sc_hd__nand2_4
X_81482_ _81482_/CLK _81482_/D _76714_/A sky130_fd_sc_hd__dfxtp_4
X_62648_ _84905_/Q _62924_/C _60220_/A _62644_/X _62647_/Y _62648_/X
+ sky130_fd_sc_hd__a41o_4
Xclkbuf_9_368_0_CLK clkbuf_8_184_0_CLK/X clkbuf_9_368_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_52401_ _52400_/X _50188_/B _52401_/Y sky130_fd_sc_hd__nand2_4
X_83221_ _83227_/CLK _72601_/Y _83221_/Q sky130_fd_sc_hd__dfxtp_4
X_80433_ _80433_/A _84311_/Q _80434_/B sky130_fd_sc_hd__xor2_4
X_68155_ _68097_/A _68155_/X sky130_fd_sc_hd__buf_2
X_53381_ _85644_/Q _53378_/X _53380_/Y _53381_/Y sky130_fd_sc_hd__o21ai_4
X_65367_ _65289_/A _65367_/B _65367_/X sky130_fd_sc_hd__and2_4
X_50593_ _50591_/Y _50577_/X _50592_/Y _86171_/D sky130_fd_sc_hd__a21boi_4
X_62579_ _60055_/A _62129_/X _59936_/X _58194_/A _62579_/Y sky130_fd_sc_hd__a22oi_4
Xclkbuf_10_800_0_CLK clkbuf_9_400_0_CLK/X _82139_/CLK sky130_fd_sc_hd__clkbuf_1
X_55120_ _46647_/B _47877_/A _55120_/C _47822_/A _55120_/X sky130_fd_sc_hd__and4_4
X_67106_ _66628_/X _67106_/X sky130_fd_sc_hd__buf_2
X_52332_ _52320_/A _49021_/A _52332_/X sky130_fd_sc_hd__and2_4
X_64318_ _64304_/A _64303_/X _84960_/Q _64318_/D _64318_/X sky130_fd_sc_hd__and4_4
X_83152_ _86534_/CLK _73414_/X _83152_/Q sky130_fd_sc_hd__dfxtp_4
X_80364_ _80353_/A _80336_/Y _80353_/B _80364_/Y sky130_fd_sc_hd__a21boi_4
X_68086_ _67948_/X _68077_/Y _67983_/X _68085_/Y _68086_/X sky130_fd_sc_hd__a211o_4
X_65298_ _64593_/A _65298_/B _65298_/X sky130_fd_sc_hd__and2_4
X_82103_ _82103_/CLK _82103_/D _77152_/A sky130_fd_sc_hd__dfxtp_4
X_55051_ _54973_/A _55070_/C sky130_fd_sc_hd__buf_2
X_67037_ _87424_/Q _67035_/X _66984_/X _67036_/X _67037_/X sky130_fd_sc_hd__a211o_4
X_52263_ _48885_/A _52267_/B _52267_/C _52263_/X sky130_fd_sc_hd__and3_4
X_64249_ _64249_/A _64249_/X sky130_fd_sc_hd__buf_2
X_87960_ _87952_/CLK _87960_/D _87960_/Q sky130_fd_sc_hd__dfxtp_4
X_83083_ _83184_/CLK _83083_/D _83083_/Q sky130_fd_sc_hd__dfxtp_4
X_80295_ _59866_/Y _80293_/A _80297_/B sky130_fd_sc_hd__nand2_4
X_54002_ _53998_/A _52482_/B _54002_/Y sky130_fd_sc_hd__nand2_4
X_51214_ _51191_/X _51203_/B _51197_/C _51214_/D _51214_/X sky130_fd_sc_hd__and4_4
X_86911_ _86878_/CLK _44909_/Y _62195_/A sky130_fd_sc_hd__dfxtp_4
X_82034_ _82005_/CLK _77880_/X _82034_/Q sky130_fd_sc_hd__dfxtp_4
X_52194_ _52194_/A _52194_/B _52218_/C _52194_/X sky130_fd_sc_hd__and3_4
Xclkbuf_10_815_0_CLK clkbuf_9_407_0_CLK/X _82596_/CLK sky130_fd_sc_hd__clkbuf_1
X_87891_ _87995_/CLK _87891_/D _87891_/Q sky130_fd_sc_hd__dfxtp_4
X_58810_ _58810_/A _58810_/X sky130_fd_sc_hd__buf_2
Xclkbuf_opt_23_CLK _86499_/CLK _86472_/CLK sky130_fd_sc_hd__clkbuf_16
X_51145_ _86065_/Q _51128_/X _51144_/Y _51145_/Y sky130_fd_sc_hd__o21ai_4
X_86842_ _84287_/CLK _86842_/D _86842_/Q sky130_fd_sc_hd__dfxtp_4
X_59790_ _59687_/Y _59790_/B _59790_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_306_0_CLK clkbuf_9_307_0_CLK/A clkbuf_9_306_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_68988_ _87578_/Q _68895_/X _68552_/X _68987_/X _68988_/X sky130_fd_sc_hd__a211o_4
X_58741_ _58641_/X _85939_/Q _58664_/X _58741_/X sky130_fd_sc_hd__o21a_4
X_51076_ _51097_/A _52768_/B _51076_/Y sky130_fd_sc_hd__nand2_4
X_55953_ _44966_/A _55619_/A _44102_/A _55952_/X _55954_/B sky130_fd_sc_hd__a211o_4
X_67939_ _67914_/X _67939_/B _67939_/X sky130_fd_sc_hd__and2_4
X_86773_ _86757_/CLK _46122_/Y _41863_/A sky130_fd_sc_hd__dfxtp_4
X_83985_ _82629_/CLK _68314_/X _82633_/D sky130_fd_sc_hd__dfxtp_4
X_50027_ _50027_/A _53240_/B _50027_/Y sky130_fd_sc_hd__nand2_4
X_54904_ _85356_/Q _54892_/X _54903_/Y _54904_/Y sky130_fd_sc_hd__o21ai_4
X_85724_ _85725_/CLK _85724_/D _85724_/Q sky130_fd_sc_hd__dfxtp_4
X_70950_ _46295_/X _70937_/X _70949_/Y _83653_/D sky130_fd_sc_hd__o21ai_4
X_58672_ _58672_/A _58649_/B _58672_/Y sky130_fd_sc_hd__nor2_4
X_82936_ _82933_/CLK _78293_/X _82936_/Q sky130_fd_sc_hd__dfxtp_4
X_55884_ _56221_/C _55531_/X _44051_/A _55883_/X _55884_/X sky130_fd_sc_hd__a211o_4
X_57623_ _57608_/X _50368_/B _57623_/Y sky130_fd_sc_hd__nand2_4
X_69609_ _88080_/Q _69607_/X _68555_/X _69608_/Y _69609_/X sky130_fd_sc_hd__a211o_4
X_54835_ _54807_/A _54857_/A sky130_fd_sc_hd__buf_2
X_85655_ _85431_/CLK _85655_/D _85655_/Q sky130_fd_sc_hd__dfxtp_4
X_70881_ _46758_/X _70855_/A _70880_/Y _70881_/Y sky130_fd_sc_hd__o21ai_4
X_82867_ _82349_/CLK _82491_/Q _82867_/Q sky130_fd_sc_hd__dfxtp_4
X_41800_ _41814_/A _41800_/X sky130_fd_sc_hd__buf_2
X_84606_ _84606_/CLK _60527_/Y _79146_/A sky130_fd_sc_hd__dfxtp_4
X_72620_ _79211_/A _59868_/X _72618_/X _72619_/Y _72620_/Y sky130_fd_sc_hd__a22oi_4
X_57554_ _84980_/Q _57550_/X _57553_/Y _57554_/Y sky130_fd_sc_hd__o21ai_4
X_81818_ _81304_/CLK _81626_/Q _81818_/Q sky130_fd_sc_hd__dfxtp_4
X_88374_ _88376_/CLK _88374_/D _88374_/Q sky130_fd_sc_hd__dfxtp_4
X_42780_ _42779_/Y _87722_/D sky130_fd_sc_hd__inv_2
X_54766_ _54775_/A _54788_/B _54775_/C _47486_/A _54766_/X sky130_fd_sc_hd__and4_4
X_85586_ _83313_/CLK _53698_/Y _85586_/Q sky130_fd_sc_hd__dfxtp_4
X_51978_ _51976_/Y _51934_/X _51977_/Y _51978_/Y sky130_fd_sc_hd__a21boi_4
X_82798_ _82425_/CLK _82830_/Q _82798_/Q sky130_fd_sc_hd__dfxtp_4
X_56505_ _56510_/A _56507_/B _55848_/B _56505_/Y sky130_fd_sc_hd__nand3_4
X_41731_ _41730_/Y _41731_/X sky130_fd_sc_hd__buf_2
Xclkbuf_5_6_0_CLK clkbuf_5_7_0_CLK/A clkbuf_5_6_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_87325_ _87045_/CLK _43654_/X _87325_/Q sky130_fd_sc_hd__dfxtp_4
X_53717_ _53714_/Y _53715_/X _53716_/X _53717_/Y sky130_fd_sc_hd__a21oi_4
X_72551_ _72572_/B _65680_/A _72551_/X sky130_fd_sc_hd__and2_4
X_84537_ _84280_/CLK _84537_/D _76985_/A sky130_fd_sc_hd__dfxtp_4
X_50929_ _50929_/A _50941_/B sky130_fd_sc_hd__buf_2
X_81749_ _81749_/CLK _76061_/B _41350_/A sky130_fd_sc_hd__dfxtp_4
X_57485_ _57485_/A _57485_/B _57485_/C _57485_/X sky130_fd_sc_hd__and3_4
X_54697_ _54682_/A _47360_/A _54697_/Y sky130_fd_sc_hd__nand2_4
X_59224_ _59154_/A _86351_/Q _59224_/Y sky130_fd_sc_hd__nor2_4
X_71502_ _71308_/A _71777_/B _71496_/C _71502_/X sky130_fd_sc_hd__and3_4
X_44450_ _44447_/X _44448_/X _41115_/X _87103_/Q _44449_/X _44451_/A
+ sky130_fd_sc_hd__o32ai_4
X_56436_ _56436_/A _56446_/B sky130_fd_sc_hd__buf_2
X_75270_ _75269_/Y _75270_/Y sky130_fd_sc_hd__inv_2
X_87256_ _87520_/CLK _43813_/Y _69509_/B sky130_fd_sc_hd__dfxtp_4
X_41662_ _41659_/X _41314_/A _41661_/X _41662_/Y sky130_fd_sc_hd__o21ai_4
X_53648_ _85595_/Q _53626_/X _53647_/Y _53648_/Y sky130_fd_sc_hd__o21ai_4
X_72482_ _72479_/Y _72481_/Y _57779_/X _72482_/X sky130_fd_sc_hd__a21o_4
X_84468_ _83216_/CLK _61588_/X _79136_/B sky130_fd_sc_hd__dfxtp_4
X_43401_ _43400_/Y _87440_/D sky130_fd_sc_hd__inv_2
X_86207_ _86203_/CLK _86207_/D _86207_/Q sky130_fd_sc_hd__dfxtp_4
X_74221_ _74211_/Y _74221_/B _74221_/Y sky130_fd_sc_hd__xnor2_4
X_40613_ _40550_/X _40556_/X _40610_/X _68498_/B _40612_/X _40614_/A
+ sky130_fd_sc_hd__o32ai_4
X_59155_ _86677_/Q _59189_/B _59155_/Y sky130_fd_sc_hd__nor2_4
X_71433_ _71420_/X _83501_/Q _71432_/X _71433_/X sky130_fd_sc_hd__a21o_4
X_83419_ _83761_/CLK _83419_/D _58526_/A sky130_fd_sc_hd__dfxtp_4
X_44381_ _44381_/A _44381_/X sky130_fd_sc_hd__buf_2
X_56367_ _56175_/A _57223_/D _56174_/X _56367_/Y sky130_fd_sc_hd__nand3_4
X_41593_ _41592_/X _41581_/X _88186_/Q _41582_/X _41593_/X sky130_fd_sc_hd__a2bb2o_4
X_87187_ _83753_/CLK _44138_/Y _87187_/Q sky130_fd_sc_hd__dfxtp_4
X_53579_ _53565_/A _50356_/B _53579_/Y sky130_fd_sc_hd__nand2_4
X_84399_ _84424_/CLK _62584_/Y _84399_/Q sky130_fd_sc_hd__dfxtp_4
X_46120_ _46120_/A _46120_/B _41863_/A _46120_/Y sky130_fd_sc_hd__nand3_4
X_58106_ _58102_/Y _58104_/Y _58105_/X _58106_/X sky130_fd_sc_hd__a21o_4
X_43332_ _43332_/A _43332_/Y sky130_fd_sc_hd__inv_2
X_55318_ _85038_/Q _55305_/X _55301_/X _55317_/X _55318_/X sky130_fd_sc_hd__a211o_4
X_74152_ _74152_/A _86568_/Q _74152_/X sky130_fd_sc_hd__and2_4
X_86138_ _85529_/CLK _86138_/D _86138_/Q sky130_fd_sc_hd__dfxtp_4
X_40544_ _40509_/X _40544_/X sky130_fd_sc_hd__buf_2
X_71364_ _71344_/A _83524_/Q _71363_/X _71364_/X sky130_fd_sc_hd__a21o_4
X_59086_ _58846_/X _85754_/Q _58847_/X _59086_/X sky130_fd_sc_hd__o21a_4
X_56298_ _56245_/A _56298_/X sky130_fd_sc_hd__buf_2
X_73103_ _83165_/Q _73079_/X _73102_/Y _73103_/X sky130_fd_sc_hd__a21o_4
X_70315_ _70328_/A _70328_/B _70315_/C _70328_/D _70315_/X sky130_fd_sc_hd__and4_4
X_46051_ _46051_/A _46051_/Y sky130_fd_sc_hd__inv_2
X_58037_ _84931_/Q _58025_/X _58029_/X _58036_/X _84931_/D sky130_fd_sc_hd__a2bb2oi_4
X_43263_ _41093_/X _43247_/X _87511_/Q _43248_/X _87511_/D sky130_fd_sc_hd__a2bb2o_4
X_55249_ _57340_/B _55126_/X _55168_/A _55248_/X _55249_/X sky130_fd_sc_hd__a211o_4
X_74083_ _73497_/A _74083_/B _74083_/X sky130_fd_sc_hd__and2_4
X_78960_ _82787_/D _78960_/B _78960_/Y sky130_fd_sc_hd__xnor2_4
X_86069_ _85751_/CLK _51126_/Y _86069_/Q sky130_fd_sc_hd__dfxtp_4
X_40475_ _40437_/X _40443_/X _40474_/X _88386_/Q _40447_/X _40475_/Y
+ sky130_fd_sc_hd__o32ai_4
X_71295_ _71303_/A _71303_/B _71672_/C _71295_/Y sky130_fd_sc_hd__nand3_4
X_45002_ _56392_/C _44945_/X _45001_/X _45002_/Y sky130_fd_sc_hd__o21ai_4
X_42214_ _42205_/X _42200_/X _41341_/X _87977_/Q _42201_/X _42215_/A
+ sky130_fd_sc_hd__o32ai_4
X_77911_ _77900_/Y _81941_/D sky130_fd_sc_hd__inv_2
X_73034_ _69698_/B _73030_/X _73031_/X _73033_/Y _73034_/X sky130_fd_sc_hd__a211o_4
X_70246_ _70246_/A _70260_/A sky130_fd_sc_hd__buf_2
X_43194_ _43162_/X _43167_/X _40909_/X _73440_/A _43172_/X _43195_/A
+ sky130_fd_sc_hd__o32ai_4
X_78891_ _82844_/Q _82556_/Q _78892_/B sky130_fd_sc_hd__xnor2_4
X_49810_ _57971_/B _49798_/X _49809_/Y _49810_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_opt_14_CLK _84906_/CLK _84778_/CLK sky130_fd_sc_hd__clkbuf_16
X_42145_ _41147_/X _42137_/X _88013_/Q _42138_/X _42145_/X sky130_fd_sc_hd__a2bb2o_4
X_77842_ _77842_/A _77841_/Y _77843_/B sky130_fd_sc_hd__xor2_4
X_70177_ _70169_/X _83848_/Q _70176_/X _83848_/D sky130_fd_sc_hd__a21o_4
X_59988_ _62576_/C _59950_/B _59985_/X _59987_/X _59512_/A _59988_/Y
+ sky130_fd_sc_hd__a41oi_4
X_49741_ _49002_/A _49825_/A sky130_fd_sc_hd__buf_2
X_46953_ _46915_/X _46944_/B _46981_/C _52771_/D _46953_/X sky130_fd_sc_hd__and4_4
X_42076_ _41878_/A _42077_/A sky130_fd_sc_hd__buf_2
X_58939_ _58939_/A _58939_/X sky130_fd_sc_hd__buf_2
X_77773_ _77773_/A _77773_/B _77774_/B sky130_fd_sc_hd__xnor2_4
X_74985_ _80949_/Q _74985_/B _81198_/D sky130_fd_sc_hd__xor2_4
X_79512_ _79510_/Y _79512_/B _79520_/A sky130_fd_sc_hd__nand2_4
X_41027_ _41024_/X _81713_/Q _41026_/X _41027_/Y sky130_fd_sc_hd__o21ai_4
X_45904_ _72973_/B _45904_/X sky130_fd_sc_hd__buf_2
X_76724_ _76719_/Y _76687_/Y _76723_/Y _76724_/Y sky130_fd_sc_hd__o21ai_4
X_61950_ _57680_/A _61902_/X _61916_/X _61948_/X _61949_/X _61950_/X
+ sky130_fd_sc_hd__a41o_4
X_49672_ _86344_/Q _49660_/X _49671_/Y _49672_/Y sky130_fd_sc_hd__o21ai_4
X_73936_ _73191_/B _74003_/B sky130_fd_sc_hd__buf_2
X_46884_ _46868_/A _46845_/X _46868_/C _52730_/D _46884_/X sky130_fd_sc_hd__and4_4
X_60901_ _60901_/A _60901_/B _60882_/X _60910_/B _60901_/X sky130_fd_sc_hd__and4_4
X_48623_ _48623_/A _48657_/C sky130_fd_sc_hd__buf_2
X_79443_ _79459_/A _79442_/Y _79443_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_7_83_0_CLK clkbuf_7_83_0_CLK/A clkbuf_7_83_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_45835_ _45835_/A _46187_/A sky130_fd_sc_hd__buf_2
X_76655_ _81395_/Q _76655_/Y sky130_fd_sc_hd__inv_2
X_61881_ _61645_/A _61881_/X sky130_fd_sc_hd__buf_2
X_73867_ _73865_/X _73866_/Y _73839_/X _73867_/X sky130_fd_sc_hd__a21o_4
X_63620_ _61579_/B _63426_/A _63358_/X _60767_/X _63619_/X _63620_/X
+ sky130_fd_sc_hd__a2111o_4
X_75606_ _75606_/A _80774_/D _75640_/A sky130_fd_sc_hd__xnor2_4
X_48554_ _81776_/Q _48136_/B _48554_/X sky130_fd_sc_hd__or2_4
X_60832_ _60663_/Y _63487_/A sky130_fd_sc_hd__inv_2
X_72818_ _72755_/X _83079_/Q _72785_/X _72817_/X _72819_/B sky130_fd_sc_hd__a211o_4
X_79374_ _79374_/A _79373_/Y _79374_/X sky130_fd_sc_hd__xor2_4
X_45766_ _45748_/X _61611_/A _45765_/X _45766_/Y sky130_fd_sc_hd__o21ai_4
X_76586_ _76585_/Y _76546_/X _76586_/X sky130_fd_sc_hd__or2_4
X_42978_ _42978_/A _42978_/Y sky130_fd_sc_hd__inv_2
X_73798_ _43055_/Y _73627_/X _73772_/X _73797_/Y _73798_/X sky130_fd_sc_hd__a211o_4
X_47505_ _47505_/A _47506_/A sky130_fd_sc_hd__inv_2
X_78325_ _78323_/X _78325_/B _78325_/X sky130_fd_sc_hd__and2_4
X_44717_ _44712_/X _44713_/X _40691_/X _73985_/A _44714_/X _44718_/A
+ sky130_fd_sc_hd__o32ai_4
X_63551_ _61509_/B _63548_/X _63549_/X _63550_/X _63551_/X sky130_fd_sc_hd__a211o_4
X_75537_ _75536_/X _75537_/Y sky130_fd_sc_hd__inv_2
X_41929_ _41894_/X _41927_/X _40661_/X _88102_/Q _41928_/X _41930_/A
+ sky130_fd_sc_hd__o32ai_4
X_72749_ _72744_/X _86209_/Q _72746_/X _72748_/X _72749_/X sky130_fd_sc_hd__a211o_4
X_48485_ _48485_/A _48485_/B _48485_/Y sky130_fd_sc_hd__nand2_4
X_60763_ _60761_/A _60761_/B _84572_/Q _60763_/Y sky130_fd_sc_hd__nor3_4
X_45697_ _45697_/A _45654_/B _45697_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_7_98_0_CLK clkbuf_7_98_0_CLK/A clkbuf_7_98_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_62502_ _61572_/A _62566_/B _62501_/X _62566_/D _62506_/B sky130_fd_sc_hd__nand4_4
X_47436_ _49406_/A _47530_/A sky130_fd_sc_hd__buf_2
X_66270_ _66237_/X _86568_/Q _66270_/X sky130_fd_sc_hd__and2_4
X_78256_ _78263_/B _78256_/B _78257_/B sky130_fd_sc_hd__xnor2_4
X_44648_ _44618_/A _44648_/X sky130_fd_sc_hd__buf_2
X_63482_ _63517_/A _63517_/B _80526_/B _63482_/Y sky130_fd_sc_hd__nor3_4
X_75468_ _75441_/X _75467_/Y _75432_/Y _75468_/Y sky130_fd_sc_hd__o21ai_4
X_60694_ _63389_/B _60694_/B _60694_/C _60694_/Y sky130_fd_sc_hd__nand3_4
X_65221_ _65397_/A _65047_/B _65221_/C _65221_/Y sky130_fd_sc_hd__nor3_4
X_77207_ _77200_/X _77207_/B _77208_/B sky130_fd_sc_hd__xor2_4
X_62433_ _62504_/A _62492_/B sky130_fd_sc_hd__buf_2
X_74419_ _83070_/Q _74412_/X _74418_/Y _74419_/Y sky130_fd_sc_hd__o21ai_4
X_47367_ _47556_/A _47408_/B sky130_fd_sc_hd__buf_2
X_78187_ _78192_/A _78191_/A _78186_/Y _78188_/B sky130_fd_sc_hd__a21boi_4
X_44579_ _44565_/X _44567_/X _40894_/X _73370_/A _44568_/X _44579_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75399_ _75399_/A _75399_/Y sky130_fd_sc_hd__inv_2
X_49106_ _49106_/A _49106_/Y sky130_fd_sc_hd__inv_2
X_65152_ _65206_/A _65152_/B _65152_/X sky130_fd_sc_hd__and2_4
X_46318_ _46318_/A _48936_/A sky130_fd_sc_hd__inv_2
X_77138_ _77135_/Y _77138_/B _77139_/B sky130_fd_sc_hd__xor2_4
X_62364_ _62276_/X _62364_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_21_0_CLK clkbuf_7_21_0_CLK/A clkbuf_8_43_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_47298_ _47297_/Y _52969_/B sky130_fd_sc_hd__buf_2
Xclkbuf_8_161_0_CLK clkbuf_7_80_0_CLK/X clkbuf_9_323_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_64103_ _58400_/A _61003_/Y _84834_/Q _60963_/X _64103_/X sky130_fd_sc_hd__a2bb2o_4
X_49037_ _86450_/Q _49003_/X _49036_/Y _49037_/Y sky130_fd_sc_hd__o21ai_4
X_61315_ _61315_/A _72550_/A _72506_/C _72607_/B _61315_/Y sky130_fd_sc_hd__nand4_4
X_46249_ _46249_/A _46279_/A sky130_fd_sc_hd__buf_2
X_65083_ _65009_/X _86159_/Q _64902_/X _65082_/X _65083_/X sky130_fd_sc_hd__a211o_4
X_69960_ _69957_/X _69959_/X _64629_/A _69960_/X sky130_fd_sc_hd__a21o_4
X_77069_ _77069_/A _82283_/D _77069_/Y sky130_fd_sc_hd__nor2_4
X_62295_ _62249_/A _63424_/B _62632_/C _62299_/C sky130_fd_sc_hd__nand3_4
X_64034_ _61549_/X _64052_/B _64003_/C _64052_/D _64034_/Y sky130_fd_sc_hd__nand4_4
X_68911_ _41957_/A _68384_/X _68745_/X _68910_/Y _68911_/X sky130_fd_sc_hd__a211o_4
X_61246_ _60933_/X _61254_/B _61243_/Y _61264_/B _61245_/Y _84499_/D
+ sky130_fd_sc_hd__a41oi_4
X_80080_ _80068_/X _80069_/X _80079_/Y _80080_/Y sky130_fd_sc_hd__a21boi_4
X_69891_ _69471_/X _69473_/X _69816_/X _69891_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_7_36_0_CLK clkbuf_6_18_0_CLK/X clkbuf_8_73_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_68842_ _88096_/Q _68384_/X _68617_/X _68841_/Y _68842_/X sky130_fd_sc_hd__a211o_4
X_61177_ _61071_/A _61177_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_176_0_CLK clkbuf_7_88_0_CLK/X clkbuf_8_176_0_CLK/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_171_0_CLK clkbuf_9_85_0_CLK/X _80912_/CLK sky130_fd_sc_hd__clkbuf_1
X_60128_ _62269_/A _62194_/A sky130_fd_sc_hd__buf_2
X_49939_ _49937_/Y _49924_/X _49938_/X _49939_/Y sky130_fd_sc_hd__a21oi_4
X_68773_ _57716_/A _68773_/X sky130_fd_sc_hd__buf_2
X_65985_ _65507_/X _66062_/B _65510_/X _65985_/Y sky130_fd_sc_hd__nand3_4
X_67724_ _67790_/A _67724_/B _67724_/X sky130_fd_sc_hd__and2_4
X_64936_ _64934_/X _83301_/Q _64864_/X _64935_/X _64936_/X sky130_fd_sc_hd__a211o_4
X_52950_ _52944_/A _52950_/B _52950_/Y sky130_fd_sc_hd__nand2_4
X_60059_ _60059_/A _60059_/B _60058_/Y _60059_/Y sky130_fd_sc_hd__nand3_4
X_83770_ _86554_/CLK _70451_/Y _83770_/Q sky130_fd_sc_hd__dfxtp_4
X_80982_ _80776_/CLK _80982_/D _80938_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_292_0_CLK clkbuf_8_146_0_CLK/X clkbuf_9_292_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_51901_ _53269_/A _51902_/A sky130_fd_sc_hd__buf_2
X_82721_ _82743_/CLK _79114_/Y _82677_/D sky130_fd_sc_hd__dfxtp_4
X_67655_ _87398_/Q _67628_/X _67581_/X _67654_/X _67655_/X sky130_fd_sc_hd__a211o_4
X_52881_ _52885_/A _52881_/B _52881_/Y sky130_fd_sc_hd__nand2_4
X_64867_ _64862_/X _64867_/B _64866_/X _64867_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_186_0_CLK clkbuf_9_93_0_CLK/X _81040_/CLK sky130_fd_sc_hd__clkbuf_1
X_54620_ _54615_/Y _54611_/X _54619_/X _85409_/D sky130_fd_sc_hd__a21oi_4
X_66606_ _66606_/A _66606_/X sky130_fd_sc_hd__buf_2
X_85440_ _85761_/CLK _85440_/D _85440_/Q sky130_fd_sc_hd__dfxtp_4
X_51832_ _51804_/A _51851_/A sky130_fd_sc_hd__buf_2
X_63818_ _63816_/X _63744_/X _63817_/Y _84293_/D sky130_fd_sc_hd__a21oi_4
X_82652_ _81746_/CLK _82652_/D _79048_/B sky130_fd_sc_hd__dfxtp_4
X_67586_ _67539_/X _88233_/Q _67586_/X sky130_fd_sc_hd__and2_4
X_64798_ _64773_/A _64798_/B _64798_/X sky130_fd_sc_hd__and2_4
X_81603_ _81603_/CLK _81603_/D _81795_/D sky130_fd_sc_hd__dfxtp_4
X_69325_ _68649_/A _69325_/X sky130_fd_sc_hd__buf_2
X_54551_ _54546_/A _53373_/B _54551_/Y sky130_fd_sc_hd__nand2_4
X_66537_ _68057_/A _66642_/A sky130_fd_sc_hd__buf_2
X_85371_ _83707_/CLK _54826_/Y _85371_/Q sky130_fd_sc_hd__dfxtp_4
X_51763_ _51789_/A _51763_/X sky130_fd_sc_hd__buf_2
X_63749_ _63749_/A _64177_/B sky130_fd_sc_hd__buf_2
X_82583_ _82589_/CLK _82615_/Q _82583_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_114_0_CLK clkbuf_7_57_0_CLK/X clkbuf_8_114_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_87110_ _87110_/CLK _87110_/D _87110_/Q sky130_fd_sc_hd__dfxtp_4
X_53502_ _85624_/Q _53476_/X _53501_/Y _53502_/Y sky130_fd_sc_hd__o21ai_4
X_84322_ _84321_/CLK _84322_/D _84322_/Q sky130_fd_sc_hd__dfxtp_4
X_50714_ _50695_/A _50714_/B _50714_/Y sky130_fd_sc_hd__nand2_4
X_57270_ _57270_/A _57270_/X sky130_fd_sc_hd__buf_2
X_81534_ _81703_/CLK _81546_/Q _76130_/A sky130_fd_sc_hd__dfxtp_4
X_69256_ _68579_/X _68582_/X _69212_/X _69256_/Y sky130_fd_sc_hd__a21oi_4
X_88090_ _88086_/CLK _88090_/D _41963_/A sky130_fd_sc_hd__dfxtp_4
X_54482_ _54401_/A _54483_/C sky130_fd_sc_hd__buf_2
X_66468_ _65307_/A _66501_/A sky130_fd_sc_hd__buf_2
X_51694_ _51694_/A _51715_/B sky130_fd_sc_hd__buf_2
X_56221_ _56214_/A _56229_/B _56221_/C _56221_/Y sky130_fd_sc_hd__nand3_4
X_68207_ _68168_/A _68207_/X sky130_fd_sc_hd__buf_2
X_87041_ _83139_/CLK _44599_/Y _87041_/Q sky130_fd_sc_hd__dfxtp_4
X_53433_ _54194_/A _53434_/A sky130_fd_sc_hd__buf_2
X_65419_ _65415_/X _65340_/X _65418_/X _65419_/Y sky130_fd_sc_hd__nand3_4
X_84253_ _83766_/CLK _64359_/X _79755_/B sky130_fd_sc_hd__dfxtp_4
X_50645_ _50645_/A _50645_/B _50645_/X sky130_fd_sc_hd__or2_4
X_81465_ _81433_/CLK _81465_/D _81465_/Q sky130_fd_sc_hd__dfxtp_4
X_69187_ _68454_/X _68457_/X _69061_/X _69187_/Y sky130_fd_sc_hd__a21oi_4
X_66399_ _66366_/X _64800_/Y _66398_/Y _66399_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_230_0_CLK clkbuf_9_230_0_CLK/A clkbuf_9_230_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_83204_ _83843_/CLK _72649_/X _70188_/C sky130_fd_sc_hd__dfxtp_4
X_80416_ _80416_/A _80416_/B _80416_/X sky130_fd_sc_hd__or2_4
X_56152_ _56127_/B _56127_/C _56152_/Y sky130_fd_sc_hd__xnor2_4
X_68138_ _68121_/X _66859_/Y _68128_/X _68137_/Y _68138_/X sky130_fd_sc_hd__a211o_4
X_53364_ _53353_/A _53364_/B _53364_/Y sky130_fd_sc_hd__nand2_4
X_84184_ _84194_/CLK _84184_/D _65698_/C sky130_fd_sc_hd__dfxtp_4
X_50576_ _86174_/Q _50499_/X _50575_/Y _50576_/Y sky130_fd_sc_hd__o21ai_4
X_81396_ _83933_/CLK _81396_/D _76967_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_129_0_CLK clkbuf_7_64_0_CLK/X clkbuf_9_259_0_CLK/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_124_0_CLK clkbuf_9_62_0_CLK/X _84396_/CLK sky130_fd_sc_hd__clkbuf_1
X_55103_ _49520_/A _55120_/C sky130_fd_sc_hd__buf_2
X_52315_ _52295_/A _48988_/A _52315_/X sky130_fd_sc_hd__and2_4
X_83135_ _83141_/CLK _83135_/D _83135_/Q sky130_fd_sc_hd__dfxtp_4
X_56083_ _55993_/Y _55994_/X _56083_/C _56083_/X sky130_fd_sc_hd__and3_4
X_80347_ _80347_/A _80347_/B _80349_/A sky130_fd_sc_hd__xnor2_4
X_68069_ _68640_/A _68069_/X sky130_fd_sc_hd__buf_2
X_53295_ _51900_/A _53295_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_754_0_CLK clkbuf_9_377_0_CLK/X _87767_/CLK sky130_fd_sc_hd__clkbuf_1
X_70100_ _83133_/Q _70100_/Y sky130_fd_sc_hd__inv_2
X_55034_ _85331_/Q _55020_/X _55033_/Y _55034_/Y sky130_fd_sc_hd__o21ai_4
X_59911_ _59910_/X _62501_/A sky130_fd_sc_hd__buf_2
X_52246_ _85860_/Q _52239_/X _52245_/Y _52246_/Y sky130_fd_sc_hd__o21ai_4
X_71080_ _71078_/A _71080_/B _71078_/C _71080_/Y sky130_fd_sc_hd__nand3_4
X_83066_ _83313_/CLK _83066_/D _83066_/Q sky130_fd_sc_hd__dfxtp_4
X_87943_ _88133_/CLK _42281_/Y _87943_/Q sky130_fd_sc_hd__dfxtp_4
X_80278_ _80277_/B _80278_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_9_245_0_CLK clkbuf_9_245_0_CLK/A clkbuf_9_245_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_82017_ _82047_/CLK _82017_/D _82017_/Q sky130_fd_sc_hd__dfxtp_4
X_70031_ _70011_/X _68701_/Y _70012_/X _70030_/Y _70031_/X sky130_fd_sc_hd__a211o_4
X_59842_ _59842_/A _59855_/A sky130_fd_sc_hd__buf_2
X_52177_ _52177_/A _52214_/A sky130_fd_sc_hd__buf_2
X_87874_ _88387_/CLK _42419_/Y _87874_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_139_0_CLK clkbuf_9_69_0_CLK/X _81265_/CLK sky130_fd_sc_hd__clkbuf_1
X_51128_ _51128_/A _51128_/X sky130_fd_sc_hd__buf_2
X_86825_ _87073_/CLK _45991_/Y _86825_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_769_0_CLK clkbuf_9_384_0_CLK/X _82515_/CLK sky130_fd_sc_hd__clkbuf_1
X_59773_ _59758_/X _59762_/Y _59763_/X _59768_/Y _59772_/Y _59773_/X
+ sky130_fd_sc_hd__a41o_4
X_56985_ _56684_/B _57149_/B _57149_/C _56985_/D _56985_/X sky130_fd_sc_hd__and4_4
X_58724_ _58711_/Y _58624_/X _58719_/X _58723_/X _84805_/D sky130_fd_sc_hd__a22oi_4
X_43950_ _43950_/A _43951_/B sky130_fd_sc_hd__inv_2
X_51059_ _86081_/Q _51047_/X _51058_/Y _51059_/Y sky130_fd_sc_hd__o21ai_4
X_55936_ _55936_/A _55936_/B _55937_/A sky130_fd_sc_hd__and2_4
X_74770_ _74770_/A _74796_/B _74797_/C _74769_/D _74772_/C sky130_fd_sc_hd__nand4_4
X_86756_ _81084_/CLK _86756_/D _42447_/D sky130_fd_sc_hd__dfxtp_4
X_71982_ _83308_/Q _57615_/X _71981_/Y _71982_/Y sky130_fd_sc_hd__o21ai_4
X_83968_ _81990_/CLK _68611_/X _83968_/Q sky130_fd_sc_hd__dfxtp_4
X_42901_ _42832_/A _42901_/X sky130_fd_sc_hd__buf_2
X_85707_ _85704_/CLK _53049_/Y _85707_/Q sky130_fd_sc_hd__dfxtp_4
X_73721_ _73718_/X _73719_/Y _73720_/X _73721_/X sky130_fd_sc_hd__a21o_4
X_58655_ _58625_/X _85466_/Q _58654_/X _58655_/Y sky130_fd_sc_hd__o21ai_4
X_70933_ HASH_ADDR[5] _70933_/B _71093_/C sky130_fd_sc_hd__nor2_4
X_82919_ _82923_/CLK _78168_/X _82919_/Q sky130_fd_sc_hd__dfxtp_4
X_43881_ _41282_/X _43879_/X _69125_/B _43880_/X _43881_/X sky130_fd_sc_hd__a2bb2o_4
X_55867_ _55549_/A _56501_/C _55867_/X sky130_fd_sc_hd__and2_4
X_86687_ _86688_/CLK _46945_/Y _59019_/A sky130_fd_sc_hd__dfxtp_4
X_83899_ _82116_/CLK _83899_/D _81971_/D sky130_fd_sc_hd__dfxtp_4
X_45620_ _85139_/Q _45507_/X _45429_/X _45620_/X sky130_fd_sc_hd__o21a_4
X_57606_ _84970_/Q _57603_/X _57605_/Y _57606_/Y sky130_fd_sc_hd__o21ai_4
X_76440_ _76440_/A _76439_/X _76440_/X sky130_fd_sc_hd__xor2_4
X_42832_ _42832_/A _42832_/X sky130_fd_sc_hd__buf_2
X_54818_ _54823_/A _47572_/Y _54818_/Y sky130_fd_sc_hd__nand2_4
X_73652_ _56934_/X _73652_/X sky130_fd_sc_hd__buf_2
X_85638_ _86054_/CLK _53415_/Y _85638_/Q sky130_fd_sc_hd__dfxtp_4
X_70864_ _46701_/X _70855_/X _70863_/Y _70864_/Y sky130_fd_sc_hd__o21ai_4
X_58586_ _58080_/A _58687_/A sky130_fd_sc_hd__buf_2
X_55798_ _83020_/Q _55306_/X _44095_/X _55797_/X _55798_/X sky130_fd_sc_hd__a211o_4
X_72603_ _72602_/X _72562_/A _72520_/X _83220_/Q _59509_/X _72603_/X
+ sky130_fd_sc_hd__o32a_4
X_45551_ _57401_/B _45551_/Y sky130_fd_sc_hd__inv_2
X_57537_ _57528_/X _57537_/B _57537_/Y sky130_fd_sc_hd__nand2_4
X_76371_ _76369_/X _76370_/Y _76371_/X sky130_fd_sc_hd__and2_4
X_88357_ _86998_/CLK _88357_/D _68735_/B sky130_fd_sc_hd__dfxtp_4
X_42763_ _41282_/X _42757_/X _69122_/B _42759_/X _87732_/D sky130_fd_sc_hd__a2bb2o_4
X_54749_ _54746_/Y _54747_/X _54748_/X _54749_/Y sky130_fd_sc_hd__a21oi_4
X_73583_ _73583_/A _73583_/B _73583_/X sky130_fd_sc_hd__and2_4
X_85569_ _83564_/CLK _53783_/Y _85569_/Q sky130_fd_sc_hd__dfxtp_4
X_70795_ _70862_/A _70841_/D sky130_fd_sc_hd__buf_2
X_78110_ _78105_/Y _78130_/A _78109_/Y _78110_/Y sky130_fd_sc_hd__a21boi_4
X_44502_ _44602_/A _44502_/X sky130_fd_sc_hd__buf_2
X_75322_ _75322_/A _75318_/X _75321_/Y _75322_/X sky130_fd_sc_hd__or3_4
X_87308_ _83158_/CLK _43689_/X _72947_/A sky130_fd_sc_hd__dfxtp_4
X_41714_ _41659_/X _41369_/A _41713_/X _41715_/A sky130_fd_sc_hd__o21ai_4
X_48270_ _48266_/Y _48233_/X _48269_/X _86545_/D sky130_fd_sc_hd__a21oi_4
X_72534_ _79476_/B _70085_/X _72533_/A _83238_/D sky130_fd_sc_hd__a21bo_4
X_79090_ _79064_/B _79090_/Y sky130_fd_sc_hd__inv_2
X_45482_ _63066_/B _61390_/A sky130_fd_sc_hd__buf_2
X_57468_ _57468_/A _56551_/X _57468_/X sky130_fd_sc_hd__or2_4
Xclkbuf_10_707_0_CLK clkbuf_9_353_0_CLK/X _87077_/CLK sky130_fd_sc_hd__clkbuf_1
X_88288_ _88288_/CLK _88288_/D _69401_/B sky130_fd_sc_hd__dfxtp_4
X_42694_ _41098_/X _42679_/X _69531_/B _42681_/X _87766_/D sky130_fd_sc_hd__a2bb2o_4
X_47221_ _47221_/A _52924_/B sky130_fd_sc_hd__buf_2
X_59207_ _59146_/X _85424_/Q _59206_/X _59207_/Y sky130_fd_sc_hd__o21ai_4
X_78041_ _77919_/Y _81943_/D sky130_fd_sc_hd__inv_2
X_44433_ _41580_/X _44431_/X _87112_/Q _44432_/X _44433_/X sky130_fd_sc_hd__a2bb2o_4
X_56419_ _56458_/A _56094_/X _56418_/Y _85201_/D sky130_fd_sc_hd__o21ai_4
X_75253_ _75251_/Y _75252_/Y _75261_/A sky130_fd_sc_hd__and2_4
X_87239_ _87758_/CLK _87239_/D _68681_/B sky130_fd_sc_hd__dfxtp_4
X_41645_ _82910_/Q _41624_/B _41645_/X sky130_fd_sc_hd__or2_4
X_72465_ _72465_/A _72465_/Y sky130_fd_sc_hd__inv_2
X_57399_ _57394_/X _56619_/X _85016_/Q _57395_/X _85016_/D sky130_fd_sc_hd__a2bb2o_4
X_74204_ _74204_/A _74095_/B _74204_/Y sky130_fd_sc_hd__nor2_4
X_47152_ _46961_/X _47152_/X sky130_fd_sc_hd__buf_2
X_59138_ _59073_/X _85750_/Q _59124_/X _59138_/X sky130_fd_sc_hd__o21a_4
X_71416_ _70692_/A _71411_/B _71450_/C _71416_/Y sky130_fd_sc_hd__nor3_4
X_44364_ _44363_/X _44364_/X sky130_fd_sc_hd__buf_2
X_75184_ _80682_/Q _80938_/D _75186_/A sky130_fd_sc_hd__xor2_4
X_41576_ _41576_/A _41576_/Y sky130_fd_sc_hd__inv_2
X_72396_ _57709_/X _85354_/Q _72395_/X _72396_/Y sky130_fd_sc_hd__o21ai_4
X_46103_ _58981_/A _72484_/A sky130_fd_sc_hd__buf_2
X_43315_ _41230_/X _43300_/X _87485_/Q _43302_/X _43315_/X sky130_fd_sc_hd__a2bb2o_4
X_74135_ _48081_/Y _74135_/B _74136_/B sky130_fd_sc_hd__xor2_4
X_40527_ _40463_/X _81158_/Q _40526_/X _40527_/Y sky130_fd_sc_hd__o21ai_4
X_47083_ _47083_/A _47084_/A sky130_fd_sc_hd__inv_2
X_59069_ _59027_/X _59066_/Y _59068_/Y _59046_/X _59031_/X _59069_/X
+ sky130_fd_sc_hd__o32a_4
X_71347_ DATA_TO_HASH[7] _71422_/C sky130_fd_sc_hd__buf_2
X_44295_ _44293_/Y _44294_/X _44277_/X _44295_/Y sky130_fd_sc_hd__a21oi_4
X_79992_ _79965_/Y _79990_/Y _79991_/Y _79992_/Y sky130_fd_sc_hd__a21oi_4
X_61100_ _61122_/A _61101_/A sky130_fd_sc_hd__inv_2
X_46034_ _46034_/A _46034_/Y sky130_fd_sc_hd__inv_2
X_43246_ _43246_/A _43246_/Y sky130_fd_sc_hd__inv_2
X_74066_ _48051_/Y _74066_/B _74066_/X sky130_fd_sc_hd__xor2_4
X_62080_ _62078_/Y _62033_/X _62079_/Y _62080_/Y sky130_fd_sc_hd__a21oi_4
X_78943_ _78930_/B _82512_/D sky130_fd_sc_hd__inv_2
X_40458_ _40456_/X _81170_/Q _40457_/X _40458_/X sky130_fd_sc_hd__o21a_4
X_71278_ _71026_/A _71279_/C sky130_fd_sc_hd__buf_2
X_61031_ _60953_/X _61030_/Y _61010_/Y _76983_/A _61020_/X _84535_/D
+ sky130_fd_sc_hd__o32a_4
X_73017_ _72963_/X _83072_/Q _73015_/X _73016_/X _73018_/B sky130_fd_sc_hd__a211o_4
X_70229_ _70229_/A _70229_/B _70229_/C _70229_/D _70229_/X sky130_fd_sc_hd__and4_4
X_43177_ _53900_/A _43177_/Y sky130_fd_sc_hd__inv_2
X_78874_ _78874_/A _78874_/B _78875_/B sky130_fd_sc_hd__nor2_4
X_40389_ _82333_/Q _40385_/B _40389_/X sky130_fd_sc_hd__or2_4
X_42128_ _41098_/X _42125_/X _88022_/Q _42126_/X _88022_/D sky130_fd_sc_hd__a2bb2o_4
X_77825_ _77825_/A _77827_/A sky130_fd_sc_hd__inv_2
X_47985_ _47980_/Y _47954_/X _47984_/X _47985_/Y sky130_fd_sc_hd__a21oi_4
X_49724_ _49708_/A _49724_/B _49724_/C _52938_/D _49724_/X sky130_fd_sc_hd__and4_4
X_46936_ _46936_/A _54451_/B sky130_fd_sc_hd__inv_2
X_42059_ _42059_/A _43129_/A sky130_fd_sc_hd__buf_2
X_65770_ _65660_/X _83059_/Q _65768_/X _65769_/X _65770_/X sky130_fd_sc_hd__a211o_4
X_77756_ _82261_/Q _81973_/Q _77756_/Y sky130_fd_sc_hd__xnor2_4
X_62982_ _61683_/X _62936_/X _62982_/C _60228_/A _62982_/Y sky130_fd_sc_hd__nand4_4
X_74968_ _74971_/B _74968_/B _74969_/B sky130_fd_sc_hd__xnor2_4
X_64721_ _65034_/A _64828_/A sky130_fd_sc_hd__buf_2
X_76707_ _76707_/A _76707_/B _76707_/X sky130_fd_sc_hd__xor2_4
X_49655_ _86347_/Q _49632_/X _49654_/Y _49655_/Y sky130_fd_sc_hd__o21ai_4
X_61933_ _62185_/B _61933_/X sky130_fd_sc_hd__buf_2
X_73919_ _41938_/Y _72899_/A _45897_/X _73918_/Y _73919_/X sky130_fd_sc_hd__a211o_4
X_46867_ _46866_/Y _52720_/D sky130_fd_sc_hd__buf_2
X_77687_ _77686_/Y _77687_/B _77687_/Y sky130_fd_sc_hd__nand2_4
X_74899_ _74899_/A _74894_/A _74899_/Y sky130_fd_sc_hd__nand2_4
X_48606_ _48606_/A _48606_/X sky130_fd_sc_hd__buf_2
X_67440_ _67513_/A _67440_/B _67440_/X sky130_fd_sc_hd__and2_4
X_79426_ _84809_/Q _84129_/Q _79433_/A sky130_fd_sc_hd__xor2_4
X_45818_ _45815_/X _45817_/Y _45803_/X _45818_/Y sky130_fd_sc_hd__a21oi_4
X_64652_ _64650_/X _86175_/Q _64583_/X _64651_/X _64652_/X sky130_fd_sc_hd__a211o_4
X_76638_ _76637_/X _76638_/Y sky130_fd_sc_hd__inv_2
X_49586_ _86360_/Q _49579_/X _49585_/Y _49586_/Y sky130_fd_sc_hd__o21ai_4
X_61864_ _61851_/X _61854_/X _61863_/Y _84745_/Q _61815_/X _61864_/Y
+ sky130_fd_sc_hd__o32ai_4
X_46798_ _46751_/A _46798_/X sky130_fd_sc_hd__buf_2
X_63603_ _63556_/X _63595_/X _63596_/X _63599_/X _63602_/Y _63603_/Y
+ sky130_fd_sc_hd__o41ai_4
X_48537_ _48613_/A _48604_/A sky130_fd_sc_hd__buf_2
X_60815_ _60622_/C _60599_/A _60182_/Y _60815_/X sky130_fd_sc_hd__and3_4
X_67371_ _87474_/Q _67274_/X _67344_/X _67370_/X _67371_/X sky130_fd_sc_hd__a211o_4
X_79357_ _79341_/Y _79344_/Y _79356_/X _79357_/X sky130_fd_sc_hd__a21o_4
X_45749_ _63265_/B _61597_/A sky130_fd_sc_hd__buf_2
X_64583_ _64776_/A _64583_/X sky130_fd_sc_hd__buf_2
X_76569_ _76566_/Y _81373_/Q _76567_/Y _76569_/Y sky130_fd_sc_hd__nand3_4
X_61795_ _61375_/B _61795_/B _61795_/C _61778_/X _61795_/Y sky130_fd_sc_hd__nand4_4
X_69110_ _69110_/A _69110_/Y sky130_fd_sc_hd__inv_2
X_66322_ _66266_/X _86212_/Q _66295_/X _66321_/X _66322_/X sky130_fd_sc_hd__a211o_4
X_78308_ _78309_/A _78309_/C _78309_/B _78308_/Y sky130_fd_sc_hd__a21oi_4
X_63534_ _58557_/A _63497_/X _61502_/A _63498_/X _63534_/X sky130_fd_sc_hd__a2bb2o_4
X_48468_ _74414_/B _48763_/B sky130_fd_sc_hd__buf_2
X_60746_ _60700_/A _60752_/B _60746_/C _60746_/Y sky130_fd_sc_hd__nor3_4
X_79288_ _79288_/A _83220_/Q _79288_/X sky130_fd_sc_hd__xor2_4
X_69041_ _80806_/D _68954_/X _69040_/X _83950_/D sky130_fd_sc_hd__a21bo_4
X_47419_ _47413_/Y _47414_/X _47418_/X _86637_/D sky130_fd_sc_hd__a21oi_4
X_66253_ _66236_/X _85609_/Q _66251_/X _66252_/X _66253_/X sky130_fd_sc_hd__a211o_4
X_78239_ _78252_/A _78239_/B _78240_/B sky130_fd_sc_hd__xor2_4
X_63465_ _59388_/A _63465_/B _63465_/C _63465_/D _63465_/Y sky130_fd_sc_hd__nand4_4
X_48399_ _83589_/Q _74383_/B sky130_fd_sc_hd__inv_2
X_60677_ _60677_/A _63478_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_1011_0_CLK clkbuf_9_505_0_CLK/X _85566_/CLK sky130_fd_sc_hd__clkbuf_1
X_65204_ _65118_/X _85546_/Q _65146_/X _65203_/X _65204_/X sky130_fd_sc_hd__a211o_4
X_50430_ _52135_/A _50430_/B _50435_/C _50430_/X sky130_fd_sc_hd__and3_4
X_62416_ _62415_/X _57680_/A _62565_/C _62355_/X _62416_/X sky130_fd_sc_hd__and4_4
X_81250_ _81250_/CLK _81250_/D _76155_/A sky130_fd_sc_hd__dfxtp_4
X_66184_ _66053_/X _85614_/Q _66096_/X _66183_/X _66184_/X sky130_fd_sc_hd__a211o_4
X_63396_ _63410_/A _63396_/B _63410_/C _63384_/D _63396_/X sky130_fd_sc_hd__and4_4
X_80201_ _80189_/A _80221_/B _80200_/X _80201_/Y sky130_fd_sc_hd__a21boi_4
X_65135_ _64601_/A _65782_/A sky130_fd_sc_hd__buf_2
X_50361_ _50359_/Y _50313_/X _50360_/X _50361_/Y sky130_fd_sc_hd__a21oi_4
X_62347_ _62196_/X _61876_/X _62346_/X _62347_/X sky130_fd_sc_hd__a21o_4
X_81181_ _81197_/CLK _75045_/B _81181_/Q sky130_fd_sc_hd__dfxtp_4
X_52100_ _52100_/A _48368_/X _52100_/Y sky130_fd_sc_hd__nand2_4
X_80132_ _84942_/Q _84190_/Q _80132_/X sky130_fd_sc_hd__xor2_4
X_53080_ _53080_/A _53080_/B _53080_/Y sky130_fd_sc_hd__nand2_4
X_65066_ _65005_/X _65066_/B _65066_/X sky130_fd_sc_hd__and2_4
X_69943_ _68823_/A _69943_/X sky130_fd_sc_hd__buf_2
X_50292_ _50290_/Y _50274_/X _50291_/Y _50292_/Y sky130_fd_sc_hd__a21boi_4
X_62278_ _62623_/C _62278_/X sky130_fd_sc_hd__buf_2
X_52031_ _52014_/X _50328_/B _52031_/Y sky130_fd_sc_hd__nand2_4
X_64017_ _64011_/Y _64013_/Y _64017_/C _64017_/D _64017_/X sky130_fd_sc_hd__and4_4
X_61229_ _61254_/C _61190_/X _61167_/Y _64454_/B _61228_/Y _84503_/D
+ sky130_fd_sc_hd__a41oi_4
X_84940_ _85489_/CLK _84940_/D _84940_/Q sky130_fd_sc_hd__dfxtp_4
X_80063_ _80047_/X _80050_/Y _80063_/X sky130_fd_sc_hd__or2_4
X_69874_ _69687_/A _69873_/Y _69874_/Y sky130_fd_sc_hd__nor2_4
X_68825_ _87841_/Q _68826_/B sky130_fd_sc_hd__inv_2
X_84871_ _84299_/CLK _58353_/Y _84871_/Q sky130_fd_sc_hd__dfxtp_4
X_86610_ _86610_/CLK _47677_/Y _72302_/A sky130_fd_sc_hd__dfxtp_4
X_83822_ _83787_/CLK _83822_/D _74778_/B sky130_fd_sc_hd__dfxtp_4
X_56770_ _83325_/Q _57010_/A sky130_fd_sc_hd__buf_2
X_68756_ _88004_/Q _68650_/X _68651_/X _68755_/X _68756_/X sky130_fd_sc_hd__a211o_4
X_87590_ _88108_/CLK _43065_/Y _73873_/A sky130_fd_sc_hd__dfxtp_4
X_53982_ _53982_/A _53982_/X sky130_fd_sc_hd__buf_2
X_65968_ _65903_/X _65494_/Y _65967_/Y _65968_/Y sky130_fd_sc_hd__o21ai_4
X_55721_ _55794_/A _56165_/C _55140_/A _55721_/Y sky130_fd_sc_hd__a21oi_4
X_67707_ _67658_/X _67707_/B _67707_/X sky130_fd_sc_hd__and2_4
X_86541_ _86541_/CLK _86541_/D _86541_/Q sky130_fd_sc_hd__dfxtp_4
X_52933_ _52852_/A _52954_/B sky130_fd_sc_hd__buf_2
X_64919_ _65669_/A _64919_/X sky130_fd_sc_hd__buf_2
X_83753_ _83753_/CLK _70542_/X _83753_/Q sky130_fd_sc_hd__dfxtp_4
X_68687_ _87091_/Q _68580_/X _68630_/X _68686_/X _68687_/X sky130_fd_sc_hd__a211o_4
X_80965_ _80962_/CLK _75604_/X _80965_/Q sky130_fd_sc_hd__dfxtp_4
X_65899_ _65789_/X _65410_/Y _65898_/Y _65899_/Y sky130_fd_sc_hd__o21ai_4
X_58440_ _84847_/Q _58440_/Y sky130_fd_sc_hd__inv_2
X_82704_ _82491_/CLK _82704_/D _78330_/B sky130_fd_sc_hd__dfxtp_4
X_67638_ _67631_/X _67635_/X _67637_/X _67638_/Y sky130_fd_sc_hd__a21oi_4
X_55652_ _83318_/Q _55652_/Y sky130_fd_sc_hd__inv_2
X_86472_ _86472_/CLK _86472_/D _86472_/Q sky130_fd_sc_hd__dfxtp_4
X_52864_ _85740_/Q _52848_/X _52863_/Y _52864_/Y sky130_fd_sc_hd__o21ai_4
X_83684_ _84807_/CLK _70847_/Y _83684_/Q sky130_fd_sc_hd__dfxtp_4
X_80896_ _81994_/CLK _75860_/X _80896_/Q sky130_fd_sc_hd__dfxtp_4
X_88211_ _87484_/CLK _41462_/X _88211_/Q sky130_fd_sc_hd__dfxtp_4
X_54603_ _54589_/X _54607_/B _54591_/C _47201_/A _54603_/X sky130_fd_sc_hd__and4_4
X_85423_ _85648_/CLK _54545_/Y _85423_/Q sky130_fd_sc_hd__dfxtp_4
X_51815_ _51805_/A _51815_/B _51810_/C _46736_/X _51815_/X sky130_fd_sc_hd__and4_4
X_58371_ _58366_/X _83763_/Q _58370_/Y _84867_/D sky130_fd_sc_hd__o21a_4
X_82635_ _87416_/CLK _82635_/D _82635_/Q sky130_fd_sc_hd__dfxtp_4
X_55583_ _85117_/Q _55527_/X _44049_/X _55582_/Y _55583_/X sky130_fd_sc_hd__a211o_4
X_67569_ _67093_/X _67569_/X sky130_fd_sc_hd__buf_2
X_52795_ _85753_/Q _52792_/X _52794_/Y _52795_/Y sky130_fd_sc_hd__o21ai_4
X_57322_ _56814_/A _57322_/B _57322_/Y sky130_fd_sc_hd__nand2_4
XPHY_11 sky130_fd_sc_hd__decap_3
X_69308_ _64777_/A _69309_/A sky130_fd_sc_hd__buf_2
X_88142_ _88398_/CLK _88142_/D _66704_/B sky130_fd_sc_hd__dfxtp_4
X_54534_ _85424_/Q _54512_/X _54533_/Y _54534_/Y sky130_fd_sc_hd__o21ai_4
X_85354_ _85354_/CLK _85354_/D _85354_/Q sky130_fd_sc_hd__dfxtp_4
X_51746_ _46892_/A _51747_/A sky130_fd_sc_hd__buf_2
XPHY_22 sky130_fd_sc_hd__decap_3
X_70580_ _70579_/Y _74731_/A sky130_fd_sc_hd__buf_2
X_82566_ _82879_/CLK _82598_/Q _82566_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_33 sky130_fd_sc_hd__decap_3
XPHY_44 sky130_fd_sc_hd__decap_3
XPHY_55 sky130_fd_sc_hd__decap_3
X_84305_ _84308_/CLK _84305_/D _80371_/B sky130_fd_sc_hd__dfxtp_4
X_57253_ _56774_/A _57359_/A sky130_fd_sc_hd__buf_2
X_81517_ _81749_/CLK _81561_/Q _81517_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_66 sky130_fd_sc_hd__decap_3
X_69239_ _69485_/A _69239_/X sky130_fd_sc_hd__buf_2
X_88073_ _88326_/CLK _42009_/Y _73033_/A sky130_fd_sc_hd__dfxtp_4
X_54465_ _85437_/Q _54457_/X _54464_/Y _54465_/Y sky130_fd_sc_hd__o21ai_4
X_85285_ _83013_/CLK _56161_/Y _85285_/Q sky130_fd_sc_hd__dfxtp_4
X_51677_ _51697_/A _53200_/B _51677_/Y sky130_fd_sc_hd__nand2_4
XPHY_77 sky130_fd_sc_hd__decap_3
X_82497_ _82589_/CLK _78801_/Y _78241_/B sky130_fd_sc_hd__dfxtp_4
XPHY_88 sky130_fd_sc_hd__decap_3
XPHY_99 sky130_fd_sc_hd__decap_3
X_56204_ _56026_/X _56195_/X _56203_/Y _85277_/D sky130_fd_sc_hd__o21ai_4
X_41430_ _41429_/X _41418_/X _88217_/Q _41419_/X _41430_/X sky130_fd_sc_hd__a2bb2o_4
X_87024_ _87032_/CLK _87024_/D _87024_/Q sky130_fd_sc_hd__dfxtp_4
X_53416_ _53405_/X _47184_/A _53416_/Y sky130_fd_sc_hd__nand2_4
X_72250_ _72250_/A _72250_/X sky130_fd_sc_hd__buf_2
X_84236_ _82797_/CLK _84236_/D _79554_/B sky130_fd_sc_hd__dfxtp_4
X_50628_ _50627_/X _49015_/X _50628_/Y sky130_fd_sc_hd__nand2_4
X_57184_ _85066_/Q _57026_/X _57184_/Y sky130_fd_sc_hd__nor2_4
X_81448_ _81575_/CLK _81448_/D _81448_/Q sky130_fd_sc_hd__dfxtp_4
X_54396_ _54393_/Y _54394_/X _54395_/X _85450_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_693_0_CLK clkbuf_9_346_0_CLK/X _87883_/CLK sky130_fd_sc_hd__clkbuf_1
X_71201_ _70382_/A _71226_/B sky130_fd_sc_hd__buf_2
X_56135_ _56104_/A _56140_/A sky130_fd_sc_hd__buf_2
X_41361_ _41360_/Y _41361_/X sky130_fd_sc_hd__buf_2
X_53347_ _53347_/A _53371_/B sky130_fd_sc_hd__buf_2
X_72181_ _72180_/X _85340_/Q _59365_/X _72181_/X sky130_fd_sc_hd__o21a_4
X_84167_ _84166_/CLK _65944_/X _84167_/Q sky130_fd_sc_hd__dfxtp_4
X_50559_ _86177_/Q _50533_/X _50558_/Y _50559_/Y sky130_fd_sc_hd__o21ai_4
X_81379_ _80784_/CLK _83915_/Q _76804_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_184_0_CLK clkbuf_8_92_0_CLK/X clkbuf_9_184_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_43100_ _43146_/A _43100_/X sky130_fd_sc_hd__buf_2
X_71132_ _50716_/B _71117_/A _71131_/Y _71132_/Y sky130_fd_sc_hd__o21ai_4
X_83118_ _86213_/CLK _74203_/X _70129_/B sky130_fd_sc_hd__dfxtp_4
X_44080_ _44079_/X _55549_/A sky130_fd_sc_hd__buf_2
X_56066_ _56052_/A _56086_/B _55889_/B _56066_/Y sky130_fd_sc_hd__nand3_4
X_41292_ _41634_/B _41292_/B _41292_/X sky130_fd_sc_hd__or2_4
X_53278_ _51914_/A _53274_/B _53293_/C _52763_/D _53278_/X sky130_fd_sc_hd__and4_4
X_84098_ _80928_/CLK _84098_/D _84098_/Q sky130_fd_sc_hd__dfxtp_4
X_43031_ _43189_/A _43031_/X sky130_fd_sc_hd__buf_2
X_55017_ _46614_/X _55017_/X sky130_fd_sc_hd__buf_2
X_52229_ _52226_/Y _52203_/X _52228_/X _85864_/D sky130_fd_sc_hd__a21oi_4
X_71063_ _52287_/B _71046_/X _71062_/Y _83620_/D sky130_fd_sc_hd__o21ai_4
X_75940_ _81701_/D _75940_/B _75940_/Y sky130_fd_sc_hd__xnor2_4
X_83049_ _83049_/CLK _74519_/Y _83049_/Q sky130_fd_sc_hd__dfxtp_4
X_87926_ _87926_/CLK _42314_/Y _87926_/Q sky130_fd_sc_hd__dfxtp_4
X_70014_ _70011_/X _68574_/Y _70012_/X _70013_/Y _70014_/X sky130_fd_sc_hd__a211o_4
X_59825_ _59794_/A _59825_/B _59825_/X sky130_fd_sc_hd__and2_4
X_75871_ _81105_/Q _80817_/Q _75872_/B sky130_fd_sc_hd__xor2_4
X_87857_ _86984_/CLK _87857_/D _87857_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_199_0_CLK clkbuf_8_99_0_CLK/X clkbuf_9_199_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_77610_ _82236_/Q _77614_/A sky130_fd_sc_hd__inv_2
X_74822_ _74822_/A _74822_/Y sky130_fd_sc_hd__inv_2
X_86808_ _86807_/CLK _86808_/D _67287_/B sky130_fd_sc_hd__dfxtp_4
X_47770_ _47765_/Y _47745_/X _47769_/X _86600_/D sky130_fd_sc_hd__a21oi_4
X_59756_ _59756_/A _59756_/X sky130_fd_sc_hd__buf_2
X_78590_ _78588_/X _78589_/Y _78602_/A sky130_fd_sc_hd__and2_4
X_44982_ _45281_/A _44982_/X sky130_fd_sc_hd__buf_2
X_56968_ _56966_/X _56643_/X _85107_/Q _56989_/A _85107_/D sky130_fd_sc_hd__a2bb2o_4
X_87788_ _87544_/CLK _42646_/Y _87788_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_631_0_CLK clkbuf_9_315_0_CLK/X _82009_/CLK sky130_fd_sc_hd__clkbuf_1
X_46721_ _46721_/A _52637_/B sky130_fd_sc_hd__inv_2
X_58707_ _58682_/X _85782_/Q _58706_/X _58707_/X sky130_fd_sc_hd__o21a_4
X_77541_ _77540_/B _77540_/C _77540_/A _77542_/A sky130_fd_sc_hd__o21a_4
X_43933_ _41429_/X _43928_/X _67955_/B _43929_/X _87193_/D sky130_fd_sc_hd__a2bb2o_4
X_55919_ _55620_/A _56306_/C _55919_/X sky130_fd_sc_hd__and2_4
X_74753_ _74731_/A _74753_/X sky130_fd_sc_hd__buf_2
X_86739_ _85815_/CLK _46418_/Y _86739_/Q sky130_fd_sc_hd__dfxtp_4
X_71965_ _48893_/A _71959_/X _71964_/X _71965_/X sky130_fd_sc_hd__and3_4
X_59687_ _59687_/A _59687_/B _59687_/C _59686_/Y _59687_/Y sky130_fd_sc_hd__nand4_4
X_56899_ _56675_/X _56876_/X _83330_/Q _56899_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_9_122_0_CLK clkbuf_8_61_0_CLK/X clkbuf_9_122_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_49440_ _49493_/A _49447_/C sky130_fd_sc_hd__buf_2
X_73704_ _73704_/A _73704_/X sky130_fd_sc_hd__buf_2
X_70916_ _70863_/A _70914_/B _70914_/C _70914_/D _70916_/Y sky130_fd_sc_hd__nand4_4
X_46652_ _86717_/Q _46622_/X _46651_/Y _46652_/Y sky130_fd_sc_hd__o21ai_4
X_58638_ _58623_/Y _58624_/X _58630_/X _58637_/X _84812_/D sky130_fd_sc_hd__a22oi_4
X_77472_ _77472_/A _77475_/B sky130_fd_sc_hd__inv_2
X_43864_ _43862_/X _43854_/X _41234_/X _68944_/B _43863_/X _43865_/A
+ sky130_fd_sc_hd__o32ai_4
X_74684_ _74684_/A _74684_/Y sky130_fd_sc_hd__inv_2
X_71896_ _70368_/X _71893_/X _71755_/X _71898_/D _71896_/Y sky130_fd_sc_hd__nand4_4
X_79211_ _79211_/A _79211_/B _79213_/A sky130_fd_sc_hd__nand2_4
X_45603_ _45598_/X _45601_/X _45602_/X _45603_/X sky130_fd_sc_hd__a21o_4
X_76423_ _76419_/Y _76422_/Y _76423_/X sky130_fd_sc_hd__xor2_4
X_42815_ _41437_/X _42802_/X _87703_/Q _42803_/X _87703_/D sky130_fd_sc_hd__a2bb2o_4
X_49371_ _49367_/Y _49316_/X _49370_/X _86400_/D sky130_fd_sc_hd__a21oi_4
X_73635_ _44675_/Y _73420_/X _73634_/Y _73635_/X sky130_fd_sc_hd__a21o_4
X_46583_ _57497_/A _52565_/B _46583_/Y sky130_fd_sc_hd__nand2_4
X_70847_ _46662_/X _70830_/Y _70846_/Y _70847_/Y sky130_fd_sc_hd__o21ai_4
X_58569_ _58100_/X _85953_/Q _58568_/X _58569_/X sky130_fd_sc_hd__o21a_4
X_43795_ _43795_/A _43795_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_646_0_CLK clkbuf_9_323_0_CLK/X _87915_/CLK sky130_fd_sc_hd__clkbuf_1
X_48322_ _49247_/A _48322_/X sky130_fd_sc_hd__buf_2
X_60600_ _60612_/A _60612_/B _79130_/A _60600_/Y sky130_fd_sc_hd__nor3_4
X_79142_ _79142_/A _79142_/B _79142_/X sky130_fd_sc_hd__xor2_4
X_45534_ _45612_/A _45597_/B sky130_fd_sc_hd__buf_2
X_76354_ _76352_/X _76353_/Y _76381_/B sky130_fd_sc_hd__and2_4
X_42746_ _42681_/A _42746_/X sky130_fd_sc_hd__buf_2
X_73566_ _73163_/A _73566_/X sky130_fd_sc_hd__buf_2
X_61580_ _84860_/Q _61580_/X sky130_fd_sc_hd__buf_2
X_70778_ _70778_/A _70869_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_137_0_CLK clkbuf_8_68_0_CLK/X clkbuf_9_137_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_75305_ _75269_/Y _75271_/X _75293_/X _75305_/X sky130_fd_sc_hd__a21bo_4
X_48253_ _48250_/Y _48226_/X _48252_/Y _86548_/D sky130_fd_sc_hd__a21boi_4
Xclkbuf_9_64_0_CLK clkbuf_9_65_0_CLK/A clkbuf_9_64_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_60531_ _60481_/X _60517_/Y _60571_/B _60529_/Y _60530_/Y _60531_/Y
+ sky130_fd_sc_hd__a41oi_4
X_72517_ _72517_/A _72517_/B _72517_/Y sky130_fd_sc_hd__nand2_4
X_79073_ _82831_/Q _82543_/Q _79089_/A sky130_fd_sc_hd__xnor2_4
X_45465_ _55590_/B _45464_/X _44919_/X _45465_/Y sky130_fd_sc_hd__o21ai_4
X_76285_ _76272_/Y _76267_/A _76267_/B _76286_/B sky130_fd_sc_hd__a21boi_4
X_42677_ _42665_/X _42666_/X _41054_/X _87774_/Q _42673_/X _42677_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73497_ _73497_/A _86468_/Q _73497_/X sky130_fd_sc_hd__and2_4
X_47204_ _47204_/A _53426_/B sky130_fd_sc_hd__inv_2
X_78024_ _78024_/A _78024_/Y sky130_fd_sc_hd__inv_2
X_44416_ _44415_/Y _87120_/D sky130_fd_sc_hd__inv_2
X_63250_ _60460_/A _63250_/X sky130_fd_sc_hd__buf_2
X_75236_ _80781_/Q _81037_/D _80749_/D sky130_fd_sc_hd__xor2_4
X_41628_ _40380_/A _41628_/X sky130_fd_sc_hd__buf_2
X_60462_ _60515_/B _60488_/A sky130_fd_sc_hd__buf_2
X_72448_ _72413_/X _72446_/Y _72447_/Y _57793_/X _72417_/X _72448_/X
+ sky130_fd_sc_hd__o32a_4
X_48184_ _48184_/A _50234_/B _48184_/Y sky130_fd_sc_hd__nand2_4
X_45396_ _45395_/X _45396_/X sky130_fd_sc_hd__buf_2
X_62201_ _60084_/A _62560_/D sky130_fd_sc_hd__buf_2
X_47135_ _47135_/A _53390_/B sky130_fd_sc_hd__inv_2
X_44347_ _41701_/X _44345_/X _87154_/Q _44346_/X _87154_/D sky130_fd_sc_hd__a2bb2o_4
X_63181_ _60482_/Y _63181_/X sky130_fd_sc_hd__buf_2
X_75167_ _75163_/X _75167_/B _81032_/D sky130_fd_sc_hd__xor2_4
X_41559_ _41548_/X _82318_/Q _41558_/X _41559_/Y sky130_fd_sc_hd__o21ai_4
X_60393_ _59613_/Y _59639_/A _60222_/C _59532_/A _60393_/X sky130_fd_sc_hd__and4_4
X_72379_ _57800_/X _72377_/Y _72378_/Y _72296_/X _59833_/X _72379_/X
+ sky130_fd_sc_hd__o32a_4
Xclkbuf_9_79_0_CLK clkbuf_9_79_0_CLK/A clkbuf_9_79_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_62132_ _62125_/X _62127_/X _62131_/Y _58352_/A _62117_/X _62132_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74118_ _83122_/Q _73549_/X _74117_/Y _83122_/D sky130_fd_sc_hd__a21o_4
X_47066_ _54526_/D _52835_/D sky130_fd_sc_hd__buf_2
X_44278_ _44266_/Y _44268_/Y _44277_/X _44278_/Y sky130_fd_sc_hd__a21oi_4
X_79975_ _79971_/X _79972_/Y _79975_/Y sky130_fd_sc_hd__nand2_4
X_75098_ _75098_/A _75100_/A _75099_/A _75104_/C sky130_fd_sc_hd__nand3_4
X_46017_ _40519_/Y _46007_/X _67179_/B _46008_/X _46017_/X sky130_fd_sc_hd__a2bb2o_4
X_43229_ _43167_/A _43229_/X sky130_fd_sc_hd__buf_2
X_66940_ _66937_/X _66939_/X _66843_/X _66940_/X sky130_fd_sc_hd__a21o_4
X_62063_ _59637_/A _62063_/X sky130_fd_sc_hd__buf_2
X_74049_ _74047_/X _74048_/Y _73982_/X _74049_/X sky130_fd_sc_hd__a21o_4
X_78926_ _78931_/B _78925_/Y _78927_/B sky130_fd_sc_hd__xnor2_4
X_61014_ _60946_/X _60838_/X _84540_/Q _61014_/Y sky130_fd_sc_hd__nor3_4
X_66871_ _66410_/A _66871_/X sky130_fd_sc_hd__buf_2
X_78857_ _78857_/A _78857_/B _78857_/X sky130_fd_sc_hd__and2_4
X_68610_ _68516_/X _68597_/Y _68447_/X _68609_/Y _68610_/X sky130_fd_sc_hd__a211o_4
X_65822_ _65638_/X _85575_/Q _65669_/X _65821_/X _65822_/X sky130_fd_sc_hd__a211o_4
X_77808_ _77806_/Y _77807_/Y _77808_/X sky130_fd_sc_hd__xor2_4
X_69590_ _69579_/X _69588_/Y _69516_/X _69589_/Y _69590_/X sky130_fd_sc_hd__a211o_4
X_47968_ _47967_/Y _47969_/B sky130_fd_sc_hd__buf_2
X_78788_ _78788_/A _82700_/Q _78788_/Y sky130_fd_sc_hd__nand2_4
X_49707_ _49678_/X _49708_/A sky130_fd_sc_hd__buf_2
X_68541_ _66565_/A _69190_/A sky130_fd_sc_hd__buf_2
X_46919_ _46914_/Y _46891_/X _46918_/X _86690_/D sky130_fd_sc_hd__a21oi_4
X_65753_ _65753_/A _73310_/B _65753_/X sky130_fd_sc_hd__and2_4
X_77739_ _78045_/A _78045_/B _77738_/Y _77739_/Y sky130_fd_sc_hd__a21oi_4
X_62965_ _62965_/A _62664_/B _62151_/X _62965_/Y sky130_fd_sc_hd__nand3_4
X_47899_ _47899_/A _73717_/A sky130_fd_sc_hd__inv_2
Xclkbuf_9_17_0_CLK clkbuf_8_8_0_CLK/X clkbuf_9_17_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_64704_ _64564_/X _64704_/X sky130_fd_sc_hd__buf_2
X_49638_ _49638_/A _52855_/B _49638_/Y sky130_fd_sc_hd__nand2_4
X_61916_ _61787_/X _61916_/X sky130_fd_sc_hd__buf_2
X_80750_ _80849_/CLK _75250_/X _81126_/D sky130_fd_sc_hd__dfxtp_4
X_68472_ _68472_/A _68472_/X sky130_fd_sc_hd__buf_2
X_65684_ _65679_/Y _65681_/X _65683_/Y _84185_/D sky130_fd_sc_hd__a21o_4
X_62896_ _60257_/X _61580_/X _62679_/X _60281_/A _84892_/Q _62897_/A
+ sky130_fd_sc_hd__a32o_4
X_67423_ _66410_/A _67423_/X sky130_fd_sc_hd__buf_2
X_79409_ _79401_/B _79418_/B _79408_/X _79410_/B sky130_fd_sc_hd__a21boi_4
X_64635_ _45943_/A _64636_/A sky130_fd_sc_hd__buf_2
X_49569_ _49569_/A _49570_/A sky130_fd_sc_hd__buf_2
X_61847_ _61863_/A _61847_/B _61843_/Y _61846_/Y _61847_/Y sky130_fd_sc_hd__nand4_4
X_80681_ _80681_/CLK _80681_/D _80681_/Q sky130_fd_sc_hd__dfxtp_4
X_51600_ _51617_/A _53127_/B _51600_/Y sky130_fd_sc_hd__nand2_4
X_82420_ _82820_/CLK _82452_/Q _78566_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_5_0_CLK clkbuf_9_5_0_CLK/A clkbuf_9_5_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_67354_ _68714_/A _67354_/X sky130_fd_sc_hd__buf_2
X_52580_ _52588_/A _52594_/B _51919_/C _52580_/D _52580_/X sky130_fd_sc_hd__and4_4
X_64566_ _64766_/A _64566_/X sky130_fd_sc_hd__buf_2
X_61778_ _59766_/X _61778_/X sky130_fd_sc_hd__buf_2
XPHY_609 sky130_fd_sc_hd__decap_3
X_66305_ _66294_/X _66303_/Y _66304_/Y _66305_/Y sky130_fd_sc_hd__o21ai_4
X_51531_ _51557_/A _51531_/X sky130_fd_sc_hd__buf_2
X_63517_ _63517_/A _63517_/B _63517_/C _63517_/Y sky130_fd_sc_hd__nor3_4
X_82351_ _82343_/CLK _77147_/X _82351_/Q sky130_fd_sc_hd__dfxtp_4
X_60729_ _78074_/A _60673_/X _60069_/Y _60702_/Y _84579_/D sky130_fd_sc_hd__a2bb2oi_4
X_67285_ _67259_/A _67285_/B _67285_/X sky130_fd_sc_hd__and2_4
X_64497_ _58973_/A _64423_/X _64496_/Y _64497_/Y sky130_fd_sc_hd__o21ai_4
X_81302_ _81257_/CLK _76990_/X _81270_/D sky130_fd_sc_hd__dfxtp_4
X_69024_ _88088_/Q _68792_/X _68933_/X _69023_/Y _69024_/X sky130_fd_sc_hd__a211o_4
X_54250_ _54250_/A _54961_/A sky130_fd_sc_hd__buf_2
X_66236_ _66053_/A _66236_/X sky130_fd_sc_hd__buf_2
X_85070_ _85039_/CLK _57161_/Y _85070_/Q sky130_fd_sc_hd__dfxtp_4
X_51462_ _51456_/A _51473_/B _51467_/C _52989_/D _51462_/X sky130_fd_sc_hd__and4_4
X_63448_ _63448_/A _63448_/B _63410_/C _63410_/D _63448_/X sky130_fd_sc_hd__and4_4
X_82282_ _82288_/CLK _81906_/Q _82282_/Q sky130_fd_sc_hd__dfxtp_4
X_53201_ _85678_/Q _53198_/X _53200_/Y _53201_/Y sky130_fd_sc_hd__o21ai_4
X_84021_ _82067_/CLK _68172_/X _82061_/D sky130_fd_sc_hd__dfxtp_4
X_50413_ _50411_/Y _50395_/X _50412_/X _50413_/Y sky130_fd_sc_hd__a21oi_4
X_81233_ _81233_/CLK _81041_/Q _81233_/Q sky130_fd_sc_hd__dfxtp_4
X_54181_ _53418_/X _54191_/A sky130_fd_sc_hd__buf_2
X_66167_ _72155_/A _86223_/Q _64692_/X _66166_/X _66167_/X sky130_fd_sc_hd__a211o_4
X_51393_ _51390_/Y _51391_/X _51392_/X _51393_/Y sky130_fd_sc_hd__a21oi_4
X_63379_ _63443_/A _63418_/C sky130_fd_sc_hd__buf_2
X_53132_ _85691_/Q _53120_/X _53131_/Y _53132_/Y sky130_fd_sc_hd__o21ai_4
X_65118_ _65118_/A _65118_/X sky130_fd_sc_hd__buf_2
X_50344_ _50342_/Y _50299_/X _50343_/Y _86220_/D sky130_fd_sc_hd__a21boi_4
X_81164_ _80792_/CLK _74920_/B _81164_/Q sky130_fd_sc_hd__dfxtp_4
X_66098_ _66053_/X _85620_/Q _66096_/X _66097_/X _66098_/X sky130_fd_sc_hd__a211o_4
X_80115_ _80107_/A _80098_/A _80115_/X sky130_fd_sc_hd__and2_4
X_65049_ _57788_/X _65049_/B _65049_/X sky130_fd_sc_hd__and2_4
X_53063_ _53074_/A _53063_/B _53074_/C _53063_/D _53063_/X sky130_fd_sc_hd__and4_4
X_57940_ _57852_/X _85714_/Q _57878_/X _57940_/X sky130_fd_sc_hd__o21a_4
X_69926_ _69922_/X _69924_/X _69925_/X _69926_/Y sky130_fd_sc_hd__a21oi_4
X_50275_ _50230_/A _50275_/B _50275_/Y sky130_fd_sc_hd__nand2_4
X_85972_ _85969_/CLK _85972_/D _85972_/Q sky130_fd_sc_hd__dfxtp_4
X_81095_ _82084_/CLK _79613_/X _81095_/Q sky130_fd_sc_hd__dfxtp_4
X_52014_ _51922_/X _52014_/X sky130_fd_sc_hd__buf_2
X_87711_ _87394_/CLK _42801_/X _67808_/B sky130_fd_sc_hd__dfxtp_4
X_84923_ _85372_/CLK _84923_/D _84923_/Q sky130_fd_sc_hd__dfxtp_4
X_80046_ _80039_/X _80046_/B _80046_/Y sky130_fd_sc_hd__nand2_4
X_57871_ _86647_/Q _57845_/X _57871_/Y sky130_fd_sc_hd__nor2_4
X_69857_ _69832_/X _69855_/Y _69815_/X _69856_/Y _69857_/X sky130_fd_sc_hd__a211o_4
X_59610_ _59609_/X _60627_/A sky130_fd_sc_hd__buf_2
X_56822_ _56758_/X _56756_/X _56761_/X _56821_/X _45957_/A _56822_/Y
+ sky130_fd_sc_hd__a41oi_4
X_68808_ _68785_/A _88354_/Q _68808_/X sky130_fd_sc_hd__and2_4
X_87642_ _86920_/CLK _87642_/D _67927_/B sky130_fd_sc_hd__dfxtp_4
X_84854_ _84732_/CLK _84854_/D _84854_/Q sky130_fd_sc_hd__dfxtp_4
X_69788_ _81969_/D _69763_/X _69787_/X _83897_/D sky130_fd_sc_hd__a21bo_4
X_83805_ _81807_/CLK _83805_/D _74770_/A sky130_fd_sc_hd__dfxtp_4
X_59541_ _59540_/Y _60407_/A sky130_fd_sc_hd__buf_2
X_56753_ _56753_/A _85134_/Q _56753_/Y sky130_fd_sc_hd__nand2_4
X_68739_ _68725_/Y _68358_/X _68649_/X _68738_/Y _68739_/X sky130_fd_sc_hd__a211o_4
X_87573_ _87826_/CLK _43109_/Y _87573_/Q sky130_fd_sc_hd__dfxtp_4
X_53965_ _53962_/Y _53892_/X _53964_/X _85533_/D sky130_fd_sc_hd__a21oi_4
X_84785_ _84906_/CLK _58971_/X _84785_/Q sky130_fd_sc_hd__dfxtp_4
X_81997_ _82133_/CLK _82029_/Q _81997_/Q sky130_fd_sc_hd__dfxtp_4
X_55704_ _55276_/A _56536_/C _55704_/X sky130_fd_sc_hd__and2_4
X_86524_ _83282_/CLK _86524_/D _86524_/Q sky130_fd_sc_hd__dfxtp_4
X_40930_ _40929_/X _40904_/X _69972_/B _40905_/X _88308_/D sky130_fd_sc_hd__a2bb2o_4
X_52916_ _52895_/A _52916_/B _52900_/C _51225_/D _52916_/X sky130_fd_sc_hd__and4_4
X_71750_ _52940_/B _71737_/X _71749_/Y _83390_/D sky130_fd_sc_hd__o21ai_4
X_59472_ _59462_/X _83459_/Q _59471_/Y _84723_/D sky130_fd_sc_hd__o21a_4
X_83736_ _83736_/CLK _83736_/D _47385_/A sky130_fd_sc_hd__dfxtp_4
X_56684_ _57270_/A _56684_/B _56684_/C _56739_/A _56685_/B sky130_fd_sc_hd__nand4_4
X_80948_ _81197_/CLK _80948_/D _80948_/Q sky130_fd_sc_hd__dfxtp_4
X_53896_ _53921_/A _53896_/X sky130_fd_sc_hd__buf_2
X_70701_ _70701_/A _70712_/A sky130_fd_sc_hd__buf_2
X_58423_ _58423_/A _58423_/X sky130_fd_sc_hd__buf_2
X_55635_ _44087_/B _55635_/B _55635_/Y sky130_fd_sc_hd__nor2_4
X_86455_ _83303_/CLK _48990_/Y _86455_/Q sky130_fd_sc_hd__dfxtp_4
X_40861_ _40861_/A _40861_/X sky130_fd_sc_hd__buf_2
X_52847_ _52844_/Y _52839_/X _52846_/X _52847_/Y sky130_fd_sc_hd__a21oi_4
X_71681_ _58485_/Y _71669_/X _71680_/Y _71681_/Y sky130_fd_sc_hd__o21ai_4
X_83667_ _86091_/CLK _70904_/Y _46824_/A sky130_fd_sc_hd__dfxtp_4
X_80879_ _80804_/CLK _75693_/B _80847_/D sky130_fd_sc_hd__dfxtp_4
X_42600_ _42600_/A _42600_/Y sky130_fd_sc_hd__inv_2
X_73420_ _56274_/X _73420_/X sky130_fd_sc_hd__buf_2
X_85406_ _85407_/CLK _85406_/D _85406_/Q sky130_fd_sc_hd__dfxtp_4
X_70632_ _70631_/X _70632_/X sky130_fd_sc_hd__buf_2
X_58354_ _84870_/Q _63316_/A sky130_fd_sc_hd__inv_2
X_82618_ _82503_/CLK _79028_/B _82586_/D sky130_fd_sc_hd__dfxtp_4
X_43580_ _40548_/X _53455_/A _87348_/Q _43185_/A _87348_/D sky130_fd_sc_hd__a2bb2o_4
X_55566_ _83002_/Q _55527_/X _44098_/X _55565_/X _56595_/B sky130_fd_sc_hd__a211o_4
X_86386_ _86384_/CLK _86386_/D _58763_/B sky130_fd_sc_hd__dfxtp_4
X_40792_ _40792_/A _40792_/X sky130_fd_sc_hd__buf_2
X_52778_ _85756_/Q _52765_/X _52777_/Y _52778_/Y sky130_fd_sc_hd__o21ai_4
X_83598_ _85542_/CLK _71126_/Y _49157_/A sky130_fd_sc_hd__dfxtp_4
X_57305_ _57010_/A _57268_/X _56767_/X _57163_/C _57305_/Y sky130_fd_sc_hd__nand4_4
X_88125_ _87116_/CLK _88125_/D _88125_/Q sky130_fd_sc_hd__dfxtp_4
X_42531_ _42517_/X _42527_/X _40739_/X _69023_/B _42519_/X _42531_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54517_ _54515_/Y _54502_/X _54516_/X _54517_/Y sky130_fd_sc_hd__a21oi_4
X_73351_ _73351_/A _73351_/X sky130_fd_sc_hd__buf_2
X_85337_ _85338_/CLK _85337_/D _85337_/Q sky130_fd_sc_hd__dfxtp_4
X_51729_ _85956_/Q _50220_/X _51728_/Y _51729_/Y sky130_fd_sc_hd__o21ai_4
X_70563_ _71215_/C _70568_/D sky130_fd_sc_hd__buf_2
X_58285_ _63655_/B _58248_/B _58285_/Y sky130_fd_sc_hd__nor2_4
X_82549_ _82369_/CLK _82549_/D _78833_/B sky130_fd_sc_hd__dfxtp_4
X_55497_ _55494_/X _55496_/X _44111_/X _55501_/A sky130_fd_sc_hd__a21o_4
X_72302_ _72302_/A _72348_/B _72302_/Y sky130_fd_sc_hd__nor2_4
X_57236_ _57235_/Y _57236_/X sky130_fd_sc_hd__buf_2
X_45250_ _55774_/B _45206_/X _45237_/X _45250_/X sky130_fd_sc_hd__o21a_4
X_76070_ _81719_/D _76070_/B _76073_/A sky130_fd_sc_hd__xor2_4
X_88056_ _88056_/CLK _42054_/Y _73438_/A sky130_fd_sc_hd__dfxtp_4
X_42462_ _42488_/A _42463_/A sky130_fd_sc_hd__buf_2
X_54448_ _54475_/A _54448_/X sky130_fd_sc_hd__buf_2
X_73282_ _73206_/X _85869_/Q _73282_/X sky130_fd_sc_hd__and2_4
X_85268_ _86900_/CLK _85268_/D _85268_/Q sky130_fd_sc_hd__dfxtp_4
X_70494_ _70696_/B _70500_/B sky130_fd_sc_hd__buf_2
X_44201_ _44139_/X _44141_/X _44142_/X _44166_/Y _44201_/Y sky130_fd_sc_hd__nand4_4
X_75021_ _75020_/Y _75021_/B _75021_/Y sky130_fd_sc_hd__nand2_4
X_87007_ _87859_/CLK _87007_/D _87007_/Q sky130_fd_sc_hd__dfxtp_4
X_41413_ _41186_/A _41435_/B sky130_fd_sc_hd__buf_2
X_72233_ _86616_/Q _72162_/B _72233_/Y sky130_fd_sc_hd__nor2_4
X_84219_ _81227_/CLK _84219_/D _84219_/Q sky130_fd_sc_hd__dfxtp_4
X_45181_ _45181_/A _45182_/A sky130_fd_sc_hd__inv_2
X_57167_ _55186_/B _57106_/X _57166_/X _85069_/D sky130_fd_sc_hd__o21ai_4
X_42393_ _40400_/X _42388_/X _87885_/Q _42389_/X _42393_/X sky130_fd_sc_hd__a2bb2o_4
X_54379_ _85453_/Q _54376_/X _54378_/Y _54379_/Y sky130_fd_sc_hd__o21ai_4
X_85199_ _85198_/CLK _85199_/D _56424_/C sky130_fd_sc_hd__dfxtp_4
X_44132_ _72784_/A _73614_/A sky130_fd_sc_hd__buf_2
X_56118_ _56118_/A _56138_/B sky130_fd_sc_hd__buf_2
X_41344_ _40365_/X _41344_/X sky130_fd_sc_hd__buf_2
X_72164_ _72151_/Y _72152_/X _72159_/X _72163_/X _83278_/D sky130_fd_sc_hd__a22oi_4
X_57098_ _57093_/Y _57221_/A sky130_fd_sc_hd__buf_2
X_71115_ _70913_/A _71115_/B _71115_/C _71115_/D _71115_/X sky130_fd_sc_hd__and4_4
X_48940_ _52291_/A _48940_/B _48928_/C _48940_/X sky130_fd_sc_hd__and3_4
X_44063_ _55470_/A _44063_/X sky130_fd_sc_hd__buf_2
X_56049_ _56171_/A _56171_/C _56048_/Y _56049_/Y sky130_fd_sc_hd__nand3_4
X_79760_ _79767_/B _79760_/B _79760_/X sky130_fd_sc_hd__xor2_4
X_41275_ _81699_/Q _41275_/B _41275_/X sky130_fd_sc_hd__or2_4
X_72095_ _72093_/Y _72083_/X _72094_/Y _83286_/D sky130_fd_sc_hd__a21boi_4
X_76972_ _84524_/Q _62616_/C _76972_/X sky130_fd_sc_hd__xor2_4
X_43014_ _43013_/X _43014_/Y sky130_fd_sc_hd__inv_2
X_78711_ _78710_/A _82685_/D _78712_/A sky130_fd_sc_hd__nand2_4
X_71046_ _71046_/A _71046_/X sky130_fd_sc_hd__buf_2
X_75923_ _61089_/C _75923_/B _80737_/D sky130_fd_sc_hd__xor2_4
X_87909_ _88220_/CLK _87909_/D _87909_/Q sky130_fd_sc_hd__dfxtp_4
X_48871_ _48869_/Y _48865_/X _48870_/X _86467_/D sky130_fd_sc_hd__a21oi_4
X_79691_ _79691_/A _79691_/B _79692_/B sky130_fd_sc_hd__xor2_4
Xclkbuf_10_570_0_CLK clkbuf_9_285_0_CLK/X _88180_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_61_0_CLK clkbuf_6_61_0_CLK/A clkbuf_6_61_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_47822_ _47822_/A _53261_/D sky130_fd_sc_hd__buf_2
X_59808_ _59824_/B _61966_/A sky130_fd_sc_hd__buf_2
X_78642_ _78605_/Y _78640_/X _78641_/Y _78642_/Y sky130_fd_sc_hd__a21oi_4
X_75854_ _75853_/X _75854_/Y sky130_fd_sc_hd__inv_2
X_74805_ _70158_/Y _70669_/A _83833_/Q _74716_/X _74805_/X sky130_fd_sc_hd__a2bb2o_4
X_47753_ _47715_/X _53227_/B _47753_/Y sky130_fd_sc_hd__nand2_4
X_59739_ _62640_/C _62717_/A sky130_fd_sc_hd__buf_2
X_78573_ _78569_/X _78574_/C _78572_/Y _78575_/A sky130_fd_sc_hd__a21o_4
X_44965_ _56027_/C _44963_/X _44964_/X _44965_/X sky130_fd_sc_hd__o21a_4
X_75785_ _81017_/Q _80889_/D _80985_/D sky130_fd_sc_hd__xor2_4
X_72997_ _72984_/Y _72996_/X _72997_/X sky130_fd_sc_hd__xor2_4
X_46704_ _46751_/A _46704_/X sky130_fd_sc_hd__buf_2
X_77524_ _77512_/A _77523_/Y _77495_/Y _77524_/Y sky130_fd_sc_hd__o21ai_4
X_43916_ _43810_/A _43916_/X sky130_fd_sc_hd__buf_2
X_62750_ _62711_/A _64307_/C _62737_/X _62738_/D _62750_/X sky130_fd_sc_hd__and4_4
X_74736_ _74716_/A _70586_/X _74731_/X _74736_/X sky130_fd_sc_hd__a21o_4
X_47684_ _47692_/A _47692_/B _47692_/C _53185_/D _47684_/X sky130_fd_sc_hd__and4_4
X_71948_ _55652_/Y _71939_/X _71947_/Y _83318_/D sky130_fd_sc_hd__o21ai_4
X_44896_ _44895_/X _45876_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_585_0_CLK clkbuf_9_292_0_CLK/X _81130_/CLK sky130_fd_sc_hd__clkbuf_1
X_49423_ _58699_/B _49415_/X _49422_/Y _49423_/Y sky130_fd_sc_hd__o21ai_4
X_61701_ _61698_/X _61699_/X _61700_/Y _61701_/Y sky130_fd_sc_hd__a21oi_4
X_46635_ _46651_/A _50893_/B _46635_/Y sky130_fd_sc_hd__nand2_4
X_77455_ _77455_/A _77455_/Y sky130_fd_sc_hd__inv_2
X_43847_ _43776_/A _43847_/X sky130_fd_sc_hd__buf_2
X_74667_ _74679_/A _74667_/B _74667_/Y sky130_fd_sc_hd__nand2_4
X_62681_ _60179_/Y _62681_/X sky130_fd_sc_hd__buf_2
X_71879_ _71857_/A _71883_/B _71873_/X _71883_/D _71879_/Y sky130_fd_sc_hd__nor4_4
X_76406_ _76406_/A _76405_/Y _76407_/B sky130_fd_sc_hd__xor2_4
X_64420_ _64377_/X _64420_/B _64391_/X _64420_/X sky130_fd_sc_hd__and3_4
X_49354_ _48917_/X _54087_/B _49354_/Y sky130_fd_sc_hd__nand2_4
X_61632_ _61632_/A _61632_/Y sky130_fd_sc_hd__inv_2
X_73618_ _73618_/A _73617_/X _73618_/Y sky130_fd_sc_hd__nand2_4
X_46566_ _86725_/Q _46543_/X _46565_/Y _46566_/Y sky130_fd_sc_hd__o21ai_4
X_77386_ _77386_/A _77386_/B _77396_/A sky130_fd_sc_hd__xor2_4
X_43778_ _43777_/Y _87272_/D sky130_fd_sc_hd__inv_2
X_74598_ _74549_/Y _74598_/X sky130_fd_sc_hd__buf_2
X_48305_ _48319_/A _48073_/B _48305_/Y sky130_fd_sc_hd__nand2_4
X_79125_ _78833_/Y _82501_/D sky130_fd_sc_hd__inv_2
X_45517_ _85113_/Q _45456_/X _45517_/Y sky130_fd_sc_hd__nor2_4
X_64351_ _59407_/A _64316_/B _64351_/Y sky130_fd_sc_hd__nor2_4
X_76337_ _76337_/A _76338_/B sky130_fd_sc_hd__buf_2
X_42729_ _42728_/Y _87748_/D sky130_fd_sc_hd__inv_2
X_61563_ _58446_/A _61563_/B _61563_/C _61563_/D _61564_/A sky130_fd_sc_hd__nand4_4
X_49285_ _48548_/A _49285_/X sky130_fd_sc_hd__buf_2
X_73549_ _73193_/A _73549_/X sky130_fd_sc_hd__buf_2
X_46497_ _54047_/A _52528_/A sky130_fd_sc_hd__buf_2
X_63302_ _63301_/X _63302_/Y sky130_fd_sc_hd__inv_2
X_60514_ _60376_/X _60512_/Y _60399_/Y _60445_/A _60513_/X _60514_/X
+ sky130_fd_sc_hd__o41a_4
X_48236_ _48204_/X _48236_/B _48236_/Y sky130_fd_sc_hd__nand2_4
X_67070_ _87870_/Q _66994_/X _67046_/X _67069_/X _67070_/X sky130_fd_sc_hd__a211o_4
X_79056_ _79057_/A _79057_/B _79057_/C _79058_/A sky130_fd_sc_hd__a21o_4
X_45448_ _45448_/A _44894_/B _45448_/Y sky130_fd_sc_hd__nor2_4
X_64282_ _64282_/A _64301_/B _64282_/Y sky130_fd_sc_hd__nor2_4
X_76268_ _76209_/Y _76223_/Y _76239_/X _76268_/D _76268_/Y sky130_fd_sc_hd__nand4_4
X_61494_ _61494_/A _61494_/Y sky130_fd_sc_hd__inv_2
X_66021_ _65400_/A _66021_/X sky130_fd_sc_hd__buf_2
X_78007_ _78007_/A _78006_/Y _78007_/Y sky130_fd_sc_hd__nand2_4
X_63233_ _79310_/A _63189_/X _63232_/Y _84342_/D sky130_fd_sc_hd__a21o_4
X_75219_ _75196_/Y _75217_/Y _75218_/Y _75219_/Y sky130_fd_sc_hd__a21oi_4
X_48167_ _48166_/Y _86561_/D sky130_fd_sc_hd__inv_2
X_60445_ _60445_/A _60444_/Y _60445_/Y sky130_fd_sc_hd__nor2_4
X_45379_ _55741_/B _45343_/X _45378_/X _45379_/X sky130_fd_sc_hd__o21a_4
X_76199_ _81349_/Q _76199_/B _76199_/Y sky130_fd_sc_hd__xnor2_4
Xclkbuf_10_523_0_CLK clkbuf_9_261_0_CLK/X _82648_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_14_0_CLK clkbuf_5_7_0_CLK/X clkbuf_7_28_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_47118_ _86668_/Q _47096_/X _47117_/Y _47118_/Y sky130_fd_sc_hd__o21ai_4
X_63164_ _58557_/A _63131_/X _63117_/X _58335_/Y _63118_/X _63164_/Y
+ sky130_fd_sc_hd__o32ai_4
X_48098_ _57619_/A _50360_/A sky130_fd_sc_hd__buf_2
X_60376_ _59875_/A _60376_/X sky130_fd_sc_hd__buf_2
X_62115_ _62113_/X _62175_/B _62046_/C _62046_/D _62115_/Y sky130_fd_sc_hd__nand4_4
X_47049_ _47044_/Y _47035_/X _47048_/X _86676_/D sky130_fd_sc_hd__a21oi_4
X_63095_ _58535_/Y _63073_/X _63059_/X _58314_/A _63060_/X _63095_/Y
+ sky130_fd_sc_hd__o32ai_4
X_67972_ _67972_/A _67972_/B _67972_/X sky130_fd_sc_hd__and2_4
X_79958_ _79958_/A _79957_/Y _79961_/A sky130_fd_sc_hd__nand2_4
X_69711_ _88072_/Q _69607_/X _68617_/X _69710_/Y _69711_/X sky130_fd_sc_hd__a211o_4
X_50060_ _50057_/Y _48865_/X _50059_/X _50060_/Y sky130_fd_sc_hd__a21oi_4
X_66923_ _66899_/X _66909_/Y _66910_/X _66922_/Y _66923_/X sky130_fd_sc_hd__a211o_4
X_62046_ _63610_/B _61999_/B _62046_/C _62046_/D _62047_/D sky130_fd_sc_hd__nand4_4
X_78909_ _82733_/Q _78909_/B _78909_/X sky130_fd_sc_hd__xor2_4
X_79889_ _79889_/A _79890_/B sky130_fd_sc_hd__inv_2
Xclkbuf_10_538_0_CLK clkbuf_9_269_0_CLK/X _82053_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_29_0_CLK clkbuf_6_29_0_CLK/A clkbuf_7_58_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_69642_ _69579_/X _69640_/Y _69604_/X _69641_/Y _69642_/X sky130_fd_sc_hd__a211o_4
X_81920_ _82015_/CLK _77708_/Y _81920_/Q sky130_fd_sc_hd__dfxtp_4
X_66854_ _66785_/A _86794_/Q _66854_/X sky130_fd_sc_hd__and2_4
X_65805_ _65623_/X _86184_/Q _65790_/X _65804_/X _65805_/X sky130_fd_sc_hd__a211o_4
X_81851_ _81872_/CLK _81883_/Q _77601_/A sky130_fd_sc_hd__dfxtp_4
X_69573_ _44514_/A _69457_/X _69458_/X _69572_/X _69574_/B sky130_fd_sc_hd__a211o_4
X_66785_ _66785_/A _66785_/B _66785_/X sky130_fd_sc_hd__and2_4
X_63997_ _63196_/B _63947_/B _64040_/C _64025_/D _63997_/Y sky130_fd_sc_hd__nand4_4
X_80802_ _83973_/CLK _80802_/D _75714_/B sky130_fd_sc_hd__dfxtp_4
X_68524_ _87001_/Q _68023_/X _68024_/X _68523_/X _68525_/B sky130_fd_sc_hd__a211o_4
X_53750_ _53750_/A _48647_/Y _53750_/Y sky130_fd_sc_hd__nand2_4
X_65736_ _65733_/X _85581_/Q _65734_/X _65735_/X _65736_/X sky130_fd_sc_hd__a211o_4
X_84570_ _84603_/CLK _60774_/X _84570_/Q sky130_fd_sc_hd__dfxtp_4
X_50962_ _86099_/Q _50936_/X _50961_/Y _50962_/Y sky130_fd_sc_hd__o21ai_4
X_62948_ _62927_/A _62926_/B _62948_/C _62948_/Y sky130_fd_sc_hd__nand3_4
X_81782_ _81703_/CLK _76121_/X _48484_/A sky130_fd_sc_hd__dfxtp_4
X_52701_ _85770_/Q _52684_/X _52700_/Y _52701_/Y sky130_fd_sc_hd__o21ai_4
X_83521_ _83521_/CLK _83521_/D _83521_/Q sky130_fd_sc_hd__dfxtp_4
X_80733_ _84280_/CLK _80733_/D _80733_/Q sky130_fd_sc_hd__dfxtp_4
X_68455_ _68059_/A _68455_/X sky130_fd_sc_hd__buf_2
X_53681_ _52161_/A _53666_/X _53692_/C _53681_/X sky130_fd_sc_hd__and3_4
X_65667_ _65667_/A _85873_/Q _65667_/X sky130_fd_sc_hd__and2_4
X_50893_ _50906_/A _50893_/B _50893_/Y sky130_fd_sc_hd__nand2_4
X_62879_ _61560_/B _62858_/X _62859_/X _62889_/D _62879_/Y sky130_fd_sc_hd__nand4_4
X_55420_ _55416_/Y _55296_/B _55417_/Y _56807_/C sky130_fd_sc_hd__nand3_4
X_67406_ _67333_/A _67406_/B _67406_/X sky130_fd_sc_hd__and2_4
X_86240_ _86436_/CLK _50231_/Y _86240_/Q sky130_fd_sc_hd__dfxtp_4
X_52632_ _52637_/A _52632_/B _52632_/Y sky130_fd_sc_hd__nand2_4
X_64618_ _64615_/X _85536_/Q _64571_/X _64617_/X _64618_/X sky130_fd_sc_hd__a211o_4
X_83452_ _83451_/CLK _71573_/X _83452_/Q sky130_fd_sc_hd__dfxtp_4
X_80664_ _80664_/CLK _80664_/D _46085_/A sky130_fd_sc_hd__dfxtp_4
X_68386_ _68386_/A _69001_/A sky130_fd_sc_hd__buf_2
X_65598_ _65596_/X _83070_/Q _65540_/X _65597_/X _65599_/B sky130_fd_sc_hd__a211o_4
X_82403_ _82797_/CLK _82435_/Q _78316_/A sky130_fd_sc_hd__dfxtp_4
X_55351_ _55352_/A _55352_/C _83753_/Q _55445_/A sky130_fd_sc_hd__a21o_4
X_67337_ _67334_/X _67336_/X _67264_/X _67340_/A sky130_fd_sc_hd__a21o_4
X_86171_ _85566_/CLK _86171_/D _86171_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_406 sky130_fd_sc_hd__decap_3
X_52563_ _52567_/A _52563_/B _52563_/Y sky130_fd_sc_hd__nand2_4
X_64549_ _64544_/X _64545_/X _64546_/X _64548_/Y _64219_/B _64549_/X
+ sky130_fd_sc_hd__o41a_4
X_83383_ _83415_/CLK _83383_/D _83383_/Q sky130_fd_sc_hd__dfxtp_4
X_80595_ _80557_/X _80561_/B _80572_/X _80570_/Y _80592_/Y _80598_/A
+ sky130_fd_sc_hd__a2111o_4
XPHY_417 sky130_fd_sc_hd__decap_3
XPHY_428 sky130_fd_sc_hd__decap_3
X_54302_ _54329_/A _54325_/B sky130_fd_sc_hd__buf_2
XPHY_439 sky130_fd_sc_hd__decap_3
X_85122_ _82980_/CLK _56929_/X _85122_/Q sky130_fd_sc_hd__dfxtp_4
X_51514_ _51514_/A _53041_/B _51514_/Y sky130_fd_sc_hd__nand2_4
X_58070_ _58070_/A _58070_/B _58070_/Y sky130_fd_sc_hd__nor2_4
X_82334_ _88268_/CLK _77208_/B _82334_/Q sky130_fd_sc_hd__dfxtp_4
X_55282_ _55145_/A _55282_/B _55282_/Y sky130_fd_sc_hd__nor2_4
X_67268_ _67268_/A _67267_/X _67268_/Y sky130_fd_sc_hd__nand2_4
X_52494_ _52448_/A _52494_/B _52494_/Y sky130_fd_sc_hd__nand2_4
X_57021_ _57019_/X _57020_/Y _56952_/A _57021_/Y sky130_fd_sc_hd__o21ai_4
X_69007_ _69007_/A _69007_/X sky130_fd_sc_hd__buf_2
X_54233_ _54231_/Y _54226_/X _54232_/X _54233_/Y sky130_fd_sc_hd__a21oi_4
X_66219_ _66217_/Y _66205_/X _66218_/X _66219_/X sky130_fd_sc_hd__a21o_4
X_85053_ _85114_/CLK _85053_/D _45460_/A sky130_fd_sc_hd__dfxtp_4
X_51445_ _51430_/X _52973_/B _51445_/Y sky130_fd_sc_hd__nand2_4
X_82265_ _83520_/CLK _80544_/X _82265_/Q sky130_fd_sc_hd__dfxtp_4
X_67199_ _87865_/Q _67176_/X _67153_/X _67198_/X _67199_/X sky130_fd_sc_hd__a211o_4
X_84004_ _81746_/CLK _68237_/X _82652_/D sky130_fd_sc_hd__dfxtp_4
X_81216_ _81216_/CLK _81216_/D _81216_/Q sky130_fd_sc_hd__dfxtp_4
X_54164_ _54217_/A _54186_/B sky130_fd_sc_hd__buf_2
X_51376_ _51367_/X _51376_/B _51376_/X sky130_fd_sc_hd__and2_4
X_82196_ _85491_/CLK _82196_/D _82196_/Q sky130_fd_sc_hd__dfxtp_4
X_53115_ _53115_/A _53115_/B _53115_/Y sky130_fd_sc_hd__nand2_4
X_50327_ _50325_/Y _50299_/X _50326_/Y _50327_/Y sky130_fd_sc_hd__a21boi_4
X_81147_ _81197_/CLK _81147_/D _40615_/A sky130_fd_sc_hd__dfxtp_4
X_54095_ _53420_/A _53428_/X _54111_/C _52927_/D _54095_/X sky130_fd_sc_hd__and4_4
X_58972_ _84784_/Q _58973_/A sky130_fd_sc_hd__inv_2
X_53046_ _53040_/X _53046_/B _53046_/Y sky130_fd_sc_hd__nand2_4
X_57923_ _58793_/A _57923_/X sky130_fd_sc_hd__buf_2
X_41060_ _41059_/X _40987_/X _88285_/Q _40989_/X _41060_/X sky130_fd_sc_hd__a2bb2o_4
X_69909_ _88057_/Q _68377_/X _69465_/X _69908_/Y _69909_/X sky130_fd_sc_hd__a211o_4
X_50258_ _47886_/X _50475_/B _50257_/X _50258_/Y sky130_fd_sc_hd__nand3_4
X_85955_ _85955_/CLK _85955_/D _85955_/Q sky130_fd_sc_hd__dfxtp_4
X_81078_ _81121_/CLK _81110_/Q _75360_/A sky130_fd_sc_hd__dfxtp_4
X_72920_ _83172_/Q _72794_/X _72919_/Y _83172_/D sky130_fd_sc_hd__a21o_4
X_80029_ _80025_/Y _80043_/B _80030_/A sky130_fd_sc_hd__xor2_4
X_84906_ _84906_/CLK _84906_/D _84906_/Q sky130_fd_sc_hd__dfxtp_4
X_57854_ _57838_/X _86009_/Q _57853_/X _57854_/Y sky130_fd_sc_hd__o21ai_4
X_50189_ _65315_/B _50185_/X _50188_/Y _50189_/Y sky130_fd_sc_hd__o21ai_4
X_85886_ _85888_/CLK _85886_/D _72836_/B sky130_fd_sc_hd__dfxtp_4
X_56805_ _56801_/X _57170_/B _56804_/Y _56805_/X sky130_fd_sc_hd__o21a_4
X_87625_ _87625_/CLK _42968_/Y _66808_/B sky130_fd_sc_hd__dfxtp_4
X_72851_ _74139_/A _73050_/A sky130_fd_sc_hd__buf_2
X_84837_ _84837_/CLK _84837_/D _84837_/Q sky130_fd_sc_hd__dfxtp_4
X_57785_ _58749_/A _57952_/A sky130_fd_sc_hd__buf_2
X_54997_ _85338_/Q _54994_/X _54996_/Y _54997_/Y sky130_fd_sc_hd__o21ai_4
X_71802_ _71800_/Y _83370_/Q _71801_/X _83370_/D sky130_fd_sc_hd__a21o_4
X_59524_ _59563_/A _59890_/B sky130_fd_sc_hd__buf_2
X_56736_ _56730_/X _56732_/X _56733_/X _56735_/X _56736_/X sky130_fd_sc_hd__and4_4
X_44750_ _44749_/Y _86976_/D sky130_fd_sc_hd__inv_2
X_75570_ _75570_/A _75887_/A _75571_/B sky130_fd_sc_hd__xor2_4
X_87556_ _87821_/CLK _43153_/Y _87556_/Q sky130_fd_sc_hd__dfxtp_4
X_41962_ _41961_/Y _88091_/D sky130_fd_sc_hd__inv_2
X_53948_ _53838_/A _53948_/X sky130_fd_sc_hd__buf_2
X_72782_ _72750_/X _85600_/Q _44130_/X _72781_/X _72782_/X sky130_fd_sc_hd__a211o_4
X_84768_ _85342_/CLK _59114_/Y _84768_/Q sky130_fd_sc_hd__dfxtp_4
X_43701_ _40826_/A _43698_/X _69722_/B _43700_/X _43701_/X sky130_fd_sc_hd__a2bb2o_4
X_74521_ _52799_/B _74517_/X _74520_/Y _74521_/Y sky130_fd_sc_hd__o21ai_4
X_86507_ _85859_/CLK _48611_/Y _86507_/Q sky130_fd_sc_hd__dfxtp_4
X_40913_ _40324_/X _82853_/Q _40912_/X _40913_/X sky130_fd_sc_hd__o21a_4
X_83719_ _83721_/CLK _83719_/D _46936_/A sky130_fd_sc_hd__dfxtp_4
X_71733_ _71729_/A _71261_/B _71724_/X _71733_/Y sky130_fd_sc_hd__nand3_4
X_59455_ _59442_/X _83464_/Q _59454_/Y _59455_/X sky130_fd_sc_hd__o21a_4
X_44681_ _44714_/A _44681_/X sky130_fd_sc_hd__buf_2
X_56667_ _56666_/Y _56667_/Y sky130_fd_sc_hd__inv_2
X_87487_ _87487_/CLK _87487_/D _87487_/Q sky130_fd_sc_hd__dfxtp_4
X_41893_ _42059_/A _43047_/A sky130_fd_sc_hd__buf_2
X_53879_ _53844_/A _53879_/B _53879_/Y sky130_fd_sc_hd__nand2_4
X_84699_ _84329_/CLK _84699_/D _80475_/A sky130_fd_sc_hd__dfxtp_4
X_46420_ _52494_/B _50799_/B sky130_fd_sc_hd__buf_2
X_58406_ _58423_/A _58406_/X sky130_fd_sc_hd__buf_2
X_77240_ _77233_/A _82082_/D _77241_/A sky130_fd_sc_hd__nor2_4
X_43632_ _43632_/A _43632_/Y sky130_fd_sc_hd__inv_2
X_55618_ _55617_/X _55619_/A sky130_fd_sc_hd__buf_2
X_74452_ _83063_/Q _74441_/X _74451_/Y _74452_/Y sky130_fd_sc_hd__o21ai_4
X_86438_ _85542_/CLK _86438_/D _65319_/B sky130_fd_sc_hd__dfxtp_4
X_40844_ _40817_/X _82290_/Q _40843_/X _40845_/A sky130_fd_sc_hd__o21ai_4
X_71664_ _71660_/A _71232_/B _71660_/C _71664_/Y sky130_fd_sc_hd__nand3_4
X_59386_ _84745_/Q _63103_/A sky130_fd_sc_hd__inv_2
X_56598_ _56629_/B _56580_/B _55552_/X _72652_/C _56597_/X _56598_/Y
+ sky130_fd_sc_hd__a41oi_4
X_73403_ _73426_/A _86472_/Q _73403_/X sky130_fd_sc_hd__and2_4
X_70615_ _70786_/A _70722_/A sky130_fd_sc_hd__buf_2
X_46351_ _46348_/X _48967_/A _46350_/X _51278_/B sky130_fd_sc_hd__o21ai_4
X_58337_ _58334_/X _58335_/Y _58336_/Y _84875_/D sky130_fd_sc_hd__a21oi_4
X_77171_ _77171_/A _77172_/B sky130_fd_sc_hd__inv_2
X_43563_ _43760_/A _43563_/X sky130_fd_sc_hd__buf_2
X_55549_ _55549_/A _56614_/B _55549_/X sky130_fd_sc_hd__and2_4
X_86369_ _83721_/CLK _49538_/Y _86369_/Q sky130_fd_sc_hd__dfxtp_4
X_74383_ _72091_/X _74383_/B _74383_/Y sky130_fd_sc_hd__nand2_4
X_40775_ _40773_/X _82303_/Q _40774_/X _40776_/A sky130_fd_sc_hd__o21ai_4
X_71595_ _71570_/X _71590_/B _71598_/C _71595_/Y sky130_fd_sc_hd__nor3_4
X_45302_ _45299_/Y _45301_/Y _45287_/X _45302_/X sky130_fd_sc_hd__a21o_4
X_76122_ _81726_/D _76133_/B _76122_/X sky130_fd_sc_hd__xor2_4
X_88108_ _88108_/CLK _41913_/X _88108_/Q sky130_fd_sc_hd__dfxtp_4
X_42514_ _42514_/A _42514_/Y sky130_fd_sc_hd__inv_2
X_49070_ _52355_/A _48940_/B _48928_/C _49070_/X sky130_fd_sc_hd__and3_4
X_73334_ _73386_/A _86507_/Q _73334_/X sky130_fd_sc_hd__and2_4
X_46282_ _52440_/B _50744_/B sky130_fd_sc_hd__buf_2
X_70546_ _70533_/X _83752_/Q _70545_/Y _70546_/X sky130_fd_sc_hd__a21o_4
X_58268_ _58268_/A _58268_/B _58268_/Y sky130_fd_sc_hd__nand2_4
X_43494_ _41731_/X _43484_/X _87392_/Q _43485_/X _87392_/D sky130_fd_sc_hd__a2bb2o_4
X_48021_ _48017_/Y _48007_/X _48020_/X _86576_/D sky130_fd_sc_hd__a21oi_4
X_45233_ _45230_/X _45232_/Y _45200_/X _45233_/Y sky130_fd_sc_hd__a21oi_4
X_57219_ _57068_/X _57153_/B _57218_/Y _85061_/D sky130_fd_sc_hd__a21o_4
X_76053_ _76063_/A _76052_/Y _81748_/D sky130_fd_sc_hd__xor2_4
X_88039_ _88044_/CLK _88039_/D _88039_/Q sky130_fd_sc_hd__dfxtp_4
X_42445_ _40556_/A _51238_/B sky130_fd_sc_hd__buf_2
X_73265_ _73407_/A _86510_/Q _73265_/X sky130_fd_sc_hd__and2_4
X_70477_ _71706_/A _70483_/B _70476_/X _70477_/X sky130_fd_sc_hd__and3_4
X_58199_ _58191_/X _58196_/Y _58198_/Y _58199_/Y sky130_fd_sc_hd__a21oi_4
X_75004_ _74995_/Y _75002_/Y _75003_/Y _75004_/X sky130_fd_sc_hd__o21a_4
X_72216_ _72166_/X _85369_/Q _72215_/X _72216_/Y sky130_fd_sc_hd__o21ai_4
X_60230_ _60244_/A _60214_/B _79872_/A _60230_/Y sky130_fd_sc_hd__nor3_4
X_45164_ _56510_/C _45134_/X _45116_/X _45164_/X sky130_fd_sc_hd__o21a_4
X_42376_ _41778_/X _42374_/X _87895_/Q _42375_/X _87895_/D sky130_fd_sc_hd__a2bb2o_4
X_73196_ _73196_/A _73196_/B _73196_/Y sky130_fd_sc_hd__nor2_4
X_44115_ _44115_/A _44118_/B sky130_fd_sc_hd__buf_2
X_79812_ _79809_/Y _79793_/B _79811_/X _79812_/Y sky130_fd_sc_hd__o21ai_4
X_41327_ _41324_/X _41674_/A _41326_/X _41327_/Y sky130_fd_sc_hd__o21ai_4
X_60161_ _60222_/C _61287_/A sky130_fd_sc_hd__buf_2
X_72147_ _72123_/X _85695_/Q _72146_/X _72147_/X sky130_fd_sc_hd__o21a_4
X_49972_ _86289_/Q _49960_/X _49971_/Y _49972_/Y sky130_fd_sc_hd__o21ai_4
X_45095_ _45095_/A _45067_/B _45095_/Y sky130_fd_sc_hd__nand2_4
X_48923_ _86461_/Q _48896_/X _48922_/Y _48923_/Y sky130_fd_sc_hd__o21ai_4
X_44046_ _44045_/X _44046_/X sky130_fd_sc_hd__buf_2
X_79743_ _79741_/X _79742_/X _79743_/Y sky130_fd_sc_hd__xnor2_4
X_41258_ _41255_/X _40732_/A _41257_/X _41259_/A sky130_fd_sc_hd__o21ai_4
X_72078_ _83289_/Q _72051_/X _72077_/Y _72078_/Y sky130_fd_sc_hd__o21ai_4
X_76955_ _81601_/Q _76955_/Y sky130_fd_sc_hd__inv_2
X_60092_ _60042_/D _60092_/B _60091_/Y _60058_/Y _60092_/Y sky130_fd_sc_hd__nand4_4
X_63920_ _64343_/B _63920_/B _63951_/C _63920_/D _63920_/Y sky130_fd_sc_hd__nand4_4
X_75906_ _61223_/C _62864_/C _75906_/X sky130_fd_sc_hd__xor2_4
X_71029_ _70994_/A _71175_/A sky130_fd_sc_hd__buf_2
Xclkbuf_4_4_1_CLK clkbuf_4_4_1_CLK/A clkbuf_4_4_1_CLK/X sky130_fd_sc_hd__clkbuf_1
X_48854_ _48667_/A _48849_/B _48854_/C _48854_/X sky130_fd_sc_hd__and3_4
X_79674_ _79660_/A _79659_/Y _79674_/X sky130_fd_sc_hd__or2_4
X_41189_ _41189_/A _41189_/X sky130_fd_sc_hd__buf_2
X_76886_ _76885_/X _76888_/B sky130_fd_sc_hd__inv_2
X_47805_ _47800_/Y _47791_/X _47804_/X _86596_/D sky130_fd_sc_hd__a21oi_4
X_78625_ _78605_/Y _78640_/B _78640_/A _78625_/Y sky130_fd_sc_hd__a21boi_4
X_63851_ _63847_/X _63833_/X _63850_/Y _63851_/Y sky130_fd_sc_hd__a21oi_4
X_75837_ _81022_/Q _80894_/D _80990_/D sky130_fd_sc_hd__xor2_4
X_48785_ _48840_/A _48785_/X sky130_fd_sc_hd__buf_2
X_45997_ _45996_/Y _86823_/D sky130_fd_sc_hd__inv_2
X_62802_ _61481_/X _62834_/B _62801_/X _62834_/D _62802_/Y sky130_fd_sc_hd__nand4_4
X_47736_ _72384_/A _47714_/X _47735_/Y _47736_/Y sky130_fd_sc_hd__o21ai_4
X_66570_ _68392_/A _69162_/A sky130_fd_sc_hd__buf_2
X_78556_ _78555_/Y _78556_/Y sky130_fd_sc_hd__inv_2
X_44948_ _44944_/Y _44947_/Y _44889_/X _44948_/X sky130_fd_sc_hd__a21o_4
X_63782_ _63765_/A _63389_/A _63765_/C _63782_/X sky130_fd_sc_hd__and3_4
X_75768_ _80920_/Q _75768_/Y sky130_fd_sc_hd__inv_2
X_60994_ _60994_/A _60994_/B _60993_/B _60994_/Y sky130_fd_sc_hd__nand3_4
X_65521_ _65285_/A _65521_/B _65521_/X sky130_fd_sc_hd__and2_4
X_77507_ _77507_/A _82101_/D _77508_/A sky130_fd_sc_hd__nand2_4
X_62733_ _62671_/A _62766_/A sky130_fd_sc_hd__buf_2
X_74719_ _70732_/X _74804_/D sky130_fd_sc_hd__buf_2
X_47667_ _47620_/X _47696_/A sky130_fd_sc_hd__buf_2
X_78487_ _82799_/Q _78487_/Y sky130_fd_sc_hd__inv_2
X_44879_ _44932_/A _45827_/B sky130_fd_sc_hd__buf_2
X_75699_ _75688_/Y _80783_/D sky130_fd_sc_hd__inv_2
X_49406_ _49406_/A _49407_/A sky130_fd_sc_hd__buf_2
X_68240_ _67489_/X _67491_/X _68239_/X _68240_/Y sky130_fd_sc_hd__a21oi_4
X_46618_ _82977_/Q _46619_/A sky130_fd_sc_hd__inv_2
X_65452_ _65350_/X _86207_/Q _65400_/X _65451_/X _65452_/X sky130_fd_sc_hd__a211o_4
X_77438_ _77418_/X _77436_/Y _77437_/Y _77438_/Y sky130_fd_sc_hd__a21oi_4
X_62664_ _61330_/X _62664_/B _60324_/A _62664_/D _62664_/Y sky130_fd_sc_hd__nand4_4
X_47598_ _47598_/A _53141_/B sky130_fd_sc_hd__buf_2
X_64403_ _64402_/X _64379_/B _84841_/Q _64403_/X sky130_fd_sc_hd__and3_4
X_49337_ _65279_/B _49334_/X _49336_/Y _49337_/Y sky130_fd_sc_hd__o21ai_4
X_61615_ _61634_/A _61634_/B _79134_/B _61615_/Y sky130_fd_sc_hd__nor3_4
X_68171_ _68144_/X _67054_/Y _68168_/X _68170_/Y _68171_/X sky130_fd_sc_hd__a211o_4
X_46549_ _82919_/Q _46527_/X _46549_/X sky130_fd_sc_hd__or2_4
X_65383_ _65379_/X _65548_/B _65383_/C _65395_/A sky130_fd_sc_hd__nand3_4
X_77369_ _77387_/A _77387_/B _77369_/X sky130_fd_sc_hd__xor2_4
X_62595_ _62592_/Y _62593_/X _62594_/Y _84398_/D sky130_fd_sc_hd__a21oi_4
X_67122_ _66879_/A _67122_/X sky130_fd_sc_hd__buf_2
X_79108_ _79104_/Y _79108_/B _79110_/A sky130_fd_sc_hd__nand2_4
X_64334_ _64319_/X _64334_/B _64333_/X _64334_/X sky130_fd_sc_hd__and3_4
X_49268_ _49266_/Y _49247_/X _49267_/Y _49268_/Y sky130_fd_sc_hd__a21boi_4
X_61546_ _61546_/A _61546_/B _61546_/C _61546_/Y sky130_fd_sc_hd__nor3_4
X_80380_ _80378_/X _80380_/B _80394_/B sky130_fd_sc_hd__xnor2_4
Xclkbuf_10_462_0_CLK clkbuf_9_231_0_CLK/X _85969_/CLK sky130_fd_sc_hd__clkbuf_1
X_48219_ _48204_/X _47924_/B _48219_/Y sky130_fd_sc_hd__nand2_4
X_67053_ _87115_/Q _66954_/X _66955_/X _67052_/X _67053_/X sky130_fd_sc_hd__a211o_4
X_79039_ _79029_/Y _79031_/B _79038_/Y _79044_/C sky130_fd_sc_hd__o21a_4
X_64265_ _64287_/A _84853_/Q _64287_/C _64265_/Y sky130_fd_sc_hd__nand3_4
X_49199_ _46600_/B _46348_/A _49199_/Y sky130_fd_sc_hd__nand2_4
X_61477_ _61518_/A _61518_/B _84478_/Q _61477_/Y sky130_fd_sc_hd__nor3_4
X_66004_ _65970_/A _66004_/B _84163_/Q _66004_/X sky130_fd_sc_hd__and3_4
X_51230_ _51149_/A _51230_/X sky130_fd_sc_hd__buf_2
X_63216_ _60469_/X _63216_/X sky130_fd_sc_hd__buf_2
X_82050_ _84074_/CLK _82050_/D _82050_/Q sky130_fd_sc_hd__dfxtp_4
X_60428_ _64386_/A _72577_/B sky130_fd_sc_hd__buf_2
X_64196_ _84866_/Q _64136_/B _64196_/Y sky130_fd_sc_hd__nor2_4
X_81001_ _80776_/CLK _84209_/Q _75635_/A sky130_fd_sc_hd__dfxtp_4
X_51161_ _51159_/Y _51147_/X _51160_/X _51161_/Y sky130_fd_sc_hd__a21oi_4
X_63147_ _63100_/A _63147_/B _63147_/C _63124_/D _63147_/X sky130_fd_sc_hd__and4_4
X_60359_ _60359_/A _60359_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_477_0_CLK clkbuf_9_238_0_CLK/X _85770_/CLK sky130_fd_sc_hd__clkbuf_1
X_50112_ _48808_/A _50113_/A sky130_fd_sc_hd__buf_2
X_51092_ _86075_/Q _51073_/X _51091_/Y _51092_/Y sky130_fd_sc_hd__o21ai_4
X_67955_ _67955_/A _67955_/B _67955_/X sky130_fd_sc_hd__and2_4
X_63078_ _63342_/C _63079_/C sky130_fd_sc_hd__buf_2
X_50043_ _72471_/B _48170_/X _50042_/Y _50043_/Y sky130_fd_sc_hd__o21ai_4
X_54920_ _54919_/X _47752_/A _54920_/Y sky130_fd_sc_hd__nand2_4
X_66906_ _66901_/X _66904_/X _66905_/X _66909_/A sky130_fd_sc_hd__a21o_4
X_62029_ _62027_/X _61999_/B _62046_/C _61971_/D _62030_/D sky130_fd_sc_hd__nand4_4
X_85740_ _85741_/CLK _52868_/Y _85740_/Q sky130_fd_sc_hd__dfxtp_4
X_82952_ _82965_/CLK _82760_/Q _82952_/Q sky130_fd_sc_hd__dfxtp_4
X_67886_ _87144_/Q _67788_/X _67789_/X _67885_/X _67887_/B sky130_fd_sc_hd__a211o_4
Xclkbuf_10_400_0_CLK clkbuf_9_200_0_CLK/X _82263_/CLK sky130_fd_sc_hd__clkbuf_1
X_81903_ _81985_/CLK _81903_/D _77036_/B sky130_fd_sc_hd__dfxtp_4
X_69625_ _69620_/X _69623_/X _69624_/X _69625_/X sky130_fd_sc_hd__a21o_4
X_54851_ _85366_/Q _54839_/X _54850_/Y _54851_/Y sky130_fd_sc_hd__o21ai_4
X_66837_ _66832_/X _66836_/X _66837_/Y sky130_fd_sc_hd__nand2_4
X_85671_ _84815_/CLK _85671_/D _85671_/Q sky130_fd_sc_hd__dfxtp_4
X_82883_ _82886_/CLK _78085_/Y _82883_/Q sky130_fd_sc_hd__dfxtp_4
X_87410_ _87922_/CLK _43462_/X _87410_/Q sky130_fd_sc_hd__dfxtp_4
X_53802_ _53797_/Y _53799_/X _53801_/Y _53802_/Y sky130_fd_sc_hd__a21boi_4
X_84622_ _84620_/CLK _60366_/Y _79581_/A sky130_fd_sc_hd__dfxtp_4
X_57570_ _84977_/Q _57562_/X _57569_/Y _57570_/Y sky130_fd_sc_hd__o21ai_4
X_81834_ _81834_/CLK _81866_/Q _77338_/A sky130_fd_sc_hd__dfxtp_4
X_69556_ _87508_/Q _69468_/X _59036_/A _69555_/X _69556_/X sky130_fd_sc_hd__a211o_4
X_88390_ _88394_/CLK _88390_/D _88390_/Q sky130_fd_sc_hd__dfxtp_4
X_54782_ _54778_/Y _54774_/X _54781_/X _85379_/D sky130_fd_sc_hd__a21oi_4
X_66768_ _66647_/A _66769_/A sky130_fd_sc_hd__buf_2
X_51994_ _51928_/X _51994_/X sky130_fd_sc_hd__buf_2
X_56521_ _56121_/X _56515_/X _56520_/Y _85164_/D sky130_fd_sc_hd__o21ai_4
X_68507_ _68503_/X _68506_/X _68429_/X _68507_/X sky130_fd_sc_hd__a21o_4
X_87341_ _87070_/CLK _43617_/X _87341_/Q sky130_fd_sc_hd__dfxtp_4
X_53733_ _53733_/A _53748_/B sky130_fd_sc_hd__buf_2
X_65719_ _65779_/A _86478_/Q _65719_/X sky130_fd_sc_hd__and2_4
X_84553_ _84529_/CLK _60899_/X _84553_/Q sky130_fd_sc_hd__dfxtp_4
X_50945_ _50256_/A _50946_/A sky130_fd_sc_hd__buf_2
X_81765_ _84003_/CLK _75996_/X _48675_/A sky130_fd_sc_hd__dfxtp_4
X_69487_ _87014_/Q _69485_/X _69361_/X _69486_/X _69487_/X sky130_fd_sc_hd__a211o_4
X_66699_ _87886_/Q _66697_/X _66675_/X _66698_/X _66699_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_415_0_CLK clkbuf_9_207_0_CLK/X _85332_/CLK sky130_fd_sc_hd__clkbuf_1
X_59240_ _59240_/A _59226_/B _59240_/Y sky130_fd_sc_hd__nor2_4
X_83504_ _84223_/CLK _71425_/X _83504_/Q sky130_fd_sc_hd__dfxtp_4
X_56452_ _56377_/X _56454_/B _56452_/C _56452_/Y sky130_fd_sc_hd__nand3_4
X_80716_ _80681_/CLK _75902_/X _80716_/Q sky130_fd_sc_hd__dfxtp_4
X_68438_ _43032_/A _68066_/X _68436_/X _68437_/X _68438_/X sky130_fd_sc_hd__a211o_4
X_87272_ _88044_/CLK _87272_/D _69288_/B sky130_fd_sc_hd__dfxtp_4
X_53664_ _85592_/Q _53660_/X _53663_/Y _53664_/Y sky130_fd_sc_hd__o21ai_4
X_84484_ _84481_/CLK _84484_/D _79152_/B sky130_fd_sc_hd__dfxtp_4
X_50876_ _50228_/X _54087_/B _50876_/Y sky130_fd_sc_hd__nand2_4
X_81696_ _81696_/CLK _80248_/X _76773_/A sky130_fd_sc_hd__dfxtp_4
X_55403_ _55403_/A _55403_/B _56777_/A sky130_fd_sc_hd__nand2_4
X_86223_ _83544_/CLK _50327_/Y _86223_/Q sky130_fd_sc_hd__dfxtp_4
X_52615_ _52613_/Y _52592_/X _52614_/X _52615_/Y sky130_fd_sc_hd__a21oi_4
X_59171_ _59159_/Y _59145_/X _59166_/X _59170_/X _59171_/Y sky130_fd_sc_hd__a22oi_4
X_83435_ _83491_/CLK _83435_/D _83435_/Q sky130_fd_sc_hd__dfxtp_4
X_56383_ _56439_/A _56383_/X sky130_fd_sc_hd__buf_2
X_80647_ _74785_/X _74711_/Y DATA_FROM_HASH[4] sky130_fd_sc_hd__ebufn_2
X_68369_ _68363_/X _68368_/X _68033_/X _68369_/X sky130_fd_sc_hd__a21o_4
X_53595_ _53604_/A _50372_/B _53595_/Y sky130_fd_sc_hd__nand2_4
XPHY_203 sky130_fd_sc_hd__decap_3
XPHY_214 sky130_fd_sc_hd__decap_3
X_58122_ _57983_/X _85379_/Q _58121_/X _58122_/Y sky130_fd_sc_hd__o21ai_4
X_70400_ _70400_/A _71005_/A sky130_fd_sc_hd__buf_2
XPHY_225 sky130_fd_sc_hd__decap_3
X_55334_ _55306_/X _45659_/Y _55334_/Y sky130_fd_sc_hd__nor2_4
X_86154_ _86154_/CLK _50685_/Y _86154_/Q sky130_fd_sc_hd__dfxtp_4
X_40560_ _40559_/X _40560_/X sky130_fd_sc_hd__buf_2
X_52546_ _85800_/Q _52500_/X _52545_/Y _52546_/Y sky130_fd_sc_hd__o21ai_4
XPHY_236 sky130_fd_sc_hd__decap_3
X_71380_ _71373_/X _83520_/Q _71379_/Y _83520_/D sky130_fd_sc_hd__a21o_4
X_83366_ _83367_/CLK _83366_/D _83366_/Q sky130_fd_sc_hd__dfxtp_4
X_80578_ _84773_/Q _65970_/C _80580_/A sky130_fd_sc_hd__xor2_4
XPHY_247 sky130_fd_sc_hd__decap_3
XPHY_258 sky130_fd_sc_hd__decap_3
XPHY_269 sky130_fd_sc_hd__decap_3
X_85105_ _85041_/CLK _85105_/D _85105_/Q sky130_fd_sc_hd__dfxtp_4
X_70331_ _70154_/X _70333_/B sky130_fd_sc_hd__buf_2
X_58053_ _58050_/Y _58052_/Y _58003_/X _58053_/X sky130_fd_sc_hd__a21o_4
X_82317_ _82317_/CLK _77081_/B _40489_/A sky130_fd_sc_hd__dfxtp_4
X_55265_ _55290_/A _55678_/A _55263_/X _55264_/Y _55265_/Y sky130_fd_sc_hd__nand4_4
X_86085_ _85764_/CLK _86085_/D _86085_/Q sky130_fd_sc_hd__dfxtp_4
X_40491_ _40490_/X _40491_/X sky130_fd_sc_hd__buf_2
X_52477_ _85814_/Q _52470_/X _52476_/Y _52477_/Y sky130_fd_sc_hd__o21ai_4
X_83297_ _83297_/CLK _72039_/Y _83297_/Q sky130_fd_sc_hd__dfxtp_4
X_57004_ _46155_/X _57004_/B _57004_/C _57004_/Y sky130_fd_sc_hd__nor3_4
X_42230_ _42230_/A _87970_/D sky130_fd_sc_hd__inv_2
X_54216_ _85482_/Q _54193_/X _54215_/Y _54216_/Y sky130_fd_sc_hd__o21ai_4
X_73050_ _73050_/A _73049_/Y _73050_/Y sky130_fd_sc_hd__nor2_4
X_85036_ _84998_/CLK _57317_/Y _85036_/Q sky130_fd_sc_hd__dfxtp_4
X_51428_ _50991_/A _51539_/A sky130_fd_sc_hd__buf_2
X_70262_ _70246_/A _70267_/A sky130_fd_sc_hd__buf_2
X_82248_ _82248_/CLK _80366_/X _82248_/Q sky130_fd_sc_hd__dfxtp_4
X_55196_ _55196_/A _55196_/B _55400_/A sky130_fd_sc_hd__and2_4
X_72001_ _72001_/A _72001_/X sky130_fd_sc_hd__buf_2
X_54147_ _54127_/X _54160_/B _54146_/X _52977_/D _54147_/X sky130_fd_sc_hd__and4_4
X_42161_ _42137_/A _42161_/X sky130_fd_sc_hd__buf_2
X_51359_ _86025_/Q _51332_/X _51358_/Y _51359_/Y sky130_fd_sc_hd__o21ai_4
X_70193_ _70193_/A _70160_/X _70162_/X _70164_/X _70193_/Y sky130_fd_sc_hd__nand4_4
X_82179_ _84951_/CLK _82179_/D _82371_/D sky130_fd_sc_hd__dfxtp_4
X_41112_ _40999_/A _41112_/X sky130_fd_sc_hd__buf_2
X_42092_ _42083_/X _42077_/X _41009_/X _88038_/Q _42078_/X _42093_/A
+ sky130_fd_sc_hd__o32ai_4
X_58955_ _58946_/Y _58857_/X _58951_/X _58954_/X _58955_/Y sky130_fd_sc_hd__a22oi_4
X_54078_ _85509_/Q _54067_/X _54077_/Y _54078_/Y sky130_fd_sc_hd__o21ai_4
X_86987_ _86998_/CLK _44722_/Y _86987_/Q sky130_fd_sc_hd__dfxtp_4
X_45920_ _45920_/A _64565_/A sky130_fd_sc_hd__buf_2
X_41043_ _41007_/A _41043_/B _41043_/X sky130_fd_sc_hd__or2_4
X_53029_ _52620_/A _53112_/A sky130_fd_sc_hd__buf_2
X_57906_ _57852_/X _85717_/Q _57878_/X _57906_/X sky130_fd_sc_hd__o21a_4
X_76740_ _76715_/Y _81354_/D sky130_fd_sc_hd__inv_2
X_73952_ _73854_/X _85617_/Q _73903_/X _73951_/X _73952_/X sky130_fd_sc_hd__a211o_4
X_85938_ _86096_/CLK _51834_/Y _85938_/Q sky130_fd_sc_hd__dfxtp_4
X_58886_ _58872_/A _86376_/Q _58886_/Y sky130_fd_sc_hd__nor2_4
X_72903_ _44526_/Y _72899_/X _72902_/Y _72904_/B sky130_fd_sc_hd__a21o_4
X_57837_ _57837_/A _58618_/A sky130_fd_sc_hd__buf_2
X_45851_ _45819_/X _61676_/A _45836_/X _45851_/Y sky130_fd_sc_hd__o21ai_4
X_76671_ _76668_/X _76669_/Y _76672_/B _76673_/A sky130_fd_sc_hd__a21o_4
X_85869_ _85859_/CLK _85869_/D _85869_/Q sky130_fd_sc_hd__dfxtp_4
X_73883_ _73954_/A _66101_/B _73883_/X sky130_fd_sc_hd__and2_4
X_78410_ _78411_/A _78411_/B _78409_/Y _78413_/A sky130_fd_sc_hd__a21oi_4
X_44802_ _44802_/A _44802_/Y sky130_fd_sc_hd__inv_2
X_87608_ _82899_/CLK _43004_/X _87608_/Q sky130_fd_sc_hd__dfxtp_4
X_75622_ _75622_/A _75622_/Y sky130_fd_sc_hd__inv_2
X_48570_ _48562_/Y _48517_/X _48569_/X _86511_/D sky130_fd_sc_hd__a21oi_4
X_72834_ _69612_/B _72803_/X _72776_/X _72834_/Y sky130_fd_sc_hd__o21ai_4
X_79390_ _79387_/X _79390_/B _82837_/D sky130_fd_sc_hd__xor2_4
X_45782_ _55248_/B _45705_/X _45389_/X _45782_/X sky130_fd_sc_hd__o21a_4
X_57768_ _58784_/A _64923_/A sky130_fd_sc_hd__buf_2
X_42994_ _52021_/A _42994_/X sky130_fd_sc_hd__buf_2
X_47521_ _47521_/A _53099_/D sky130_fd_sc_hd__buf_2
X_59507_ _46159_/X _59504_/Y _59506_/Y _59507_/Y sky130_fd_sc_hd__a21oi_4
X_78341_ _78341_/A _82756_/D _78341_/X sky130_fd_sc_hd__xor2_4
X_44733_ _44733_/A _49210_/A sky130_fd_sc_hd__buf_2
X_56719_ _56719_/A _56719_/B _46237_/A _56724_/A sky130_fd_sc_hd__nand3_4
X_75553_ _75562_/A _75552_/X _75553_/Y sky130_fd_sc_hd__nand2_4
X_87539_ _88087_/CLK _43205_/X _87539_/Q sky130_fd_sc_hd__dfxtp_4
X_41945_ _41932_/X _41927_/X _40691_/X _73987_/A _41928_/X _41945_/Y
+ sky130_fd_sc_hd__o32ai_4
X_72765_ _72765_/A _74140_/A sky130_fd_sc_hd__buf_2
X_57699_ _58602_/A _58098_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_42_0_CLK clkbuf_8_43_0_CLK/A clkbuf_8_42_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_74504_ _83052_/Q _46250_/X _74503_/Y _74504_/Y sky130_fd_sc_hd__o21ai_4
X_47452_ _47444_/A _53054_/B _47452_/Y sky130_fd_sc_hd__nand2_4
X_71716_ _71160_/C _71716_/B _70763_/A _71716_/D _71716_/X sky130_fd_sc_hd__and4_4
X_59438_ _59426_/X _59436_/Y _59437_/Y _59438_/Y sky130_fd_sc_hd__a21oi_4
X_78272_ _78271_/X _78274_/A sky130_fd_sc_hd__buf_2
X_44664_ _41098_/A _44648_/X _87010_/Q _44650_/X _44664_/X sky130_fd_sc_hd__a2bb2o_4
X_75484_ _75506_/D _75486_/A sky130_fd_sc_hd__inv_2
X_41876_ _41875_/Y _88114_/D sky130_fd_sc_hd__inv_2
X_72696_ _70239_/C _72686_/X _72695_/Y _83186_/D sky130_fd_sc_hd__a21bo_4
X_46403_ _47904_/A _46403_/X sky130_fd_sc_hd__buf_2
X_77223_ _77223_/A _77222_/Y _77223_/Y sky130_fd_sc_hd__nand2_4
X_43615_ _40610_/A _43609_/X _68495_/B _43611_/X _43616_/A sky130_fd_sc_hd__a2bb2o_4
X_74435_ _48522_/A _74420_/X _74425_/X _74435_/X sky130_fd_sc_hd__and3_4
X_40827_ _40758_/X _40759_/X _40826_/X _69725_/B _40744_/X _40828_/A
+ sky130_fd_sc_hd__o32ai_4
X_47383_ _57563_/A _47525_/A sky130_fd_sc_hd__buf_2
X_59369_ _59219_/X _85731_/Q _59220_/X _59369_/X sky130_fd_sc_hd__o21a_4
X_71647_ _59504_/Y _71628_/A _71646_/Y _71647_/Y sky130_fd_sc_hd__o21ai_4
X_44595_ _87042_/Q _44595_/Y sky130_fd_sc_hd__inv_2
X_49122_ _49080_/A _53902_/B _49122_/X sky130_fd_sc_hd__and2_4
X_61400_ _61302_/Y _61400_/X sky130_fd_sc_hd__buf_2
X_46334_ _53976_/B _49241_/B sky130_fd_sc_hd__buf_2
X_77154_ _77154_/A _77151_/A _77155_/B sky130_fd_sc_hd__and2_4
X_43546_ _43760_/A _43546_/X sky130_fd_sc_hd__buf_2
X_62380_ _61460_/B _62278_/X _62363_/X _62323_/X _62379_/X _62380_/X
+ sky130_fd_sc_hd__a41o_4
X_74366_ _74366_/A _72113_/B _74366_/C _74366_/X sky130_fd_sc_hd__and3_4
X_40758_ _40835_/A _40758_/X sky130_fd_sc_hd__buf_2
X_71578_ _71556_/Y _83450_/Q _71577_/Y _71578_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_8_57_0_CLK clkbuf_8_57_0_CLK/A clkbuf_8_57_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_76105_ _81724_/D _76126_/C _76112_/A sky130_fd_sc_hd__xor2_4
X_49053_ _48898_/A _49056_/A sky130_fd_sc_hd__buf_2
X_73317_ _83156_/Q _73193_/X _73316_/Y _73317_/X sky130_fd_sc_hd__a21o_4
X_61331_ _72563_/C _61377_/C sky130_fd_sc_hd__buf_2
X_46265_ _46265_/A _46328_/B _46265_/X sky130_fd_sc_hd__or2_4
X_70529_ _70694_/A _71823_/A sky130_fd_sc_hd__buf_2
X_77085_ _77077_/A _77066_/A _82284_/D _77085_/Y sky130_fd_sc_hd__nand3_4
X_43477_ _43477_/A _43477_/Y sky130_fd_sc_hd__inv_2
X_74297_ _74297_/A _74297_/B _74297_/C _74297_/Y sky130_fd_sc_hd__nand3_4
X_40689_ _40689_/A _40654_/B _40689_/X sky130_fd_sc_hd__or2_4
X_48004_ _48004_/A _50310_/B _48004_/Y sky130_fd_sc_hd__nand2_4
X_45216_ _45216_/A _45199_/B _45216_/Y sky130_fd_sc_hd__nand2_4
X_64050_ _62027_/X _64095_/B _64050_/C _64095_/D _64050_/Y sky130_fd_sc_hd__nand4_4
X_76036_ _76028_/A _81712_/D _76036_/C _76037_/A sky130_fd_sc_hd__nand3_4
X_42428_ _40507_/X _42414_/X _87868_/Q _42415_/X _42428_/X sky130_fd_sc_hd__a2bb2o_4
X_61262_ _61262_/A _72544_/B _61262_/C _61262_/Y sky130_fd_sc_hd__nor3_4
X_73248_ _69820_/Y _73224_/X _73194_/X _73247_/Y _73248_/X sky130_fd_sc_hd__a211o_4
X_46196_ _46196_/A _74842_/B _46195_/Y _86762_/D sky130_fd_sc_hd__and3_4
X_63001_ _63001_/A _63281_/B sky130_fd_sc_hd__buf_2
X_60213_ _60105_/X _60244_/A sky130_fd_sc_hd__buf_2
X_45147_ _45297_/A _45147_/X sky130_fd_sc_hd__buf_2
X_42359_ _42350_/X _42346_/X _41735_/X _87903_/Q _42347_/X _42360_/A
+ sky130_fd_sc_hd__o32ai_4
X_61193_ _61190_/X _61154_/X _61170_/Y _61173_/Y _61192_/Y _84510_/D
+ sky130_fd_sc_hd__a41oi_4
X_73179_ _73176_/X _73178_/X _72866_/X _73179_/X sky130_fd_sc_hd__a21o_4
X_60144_ _60143_/X _60144_/Y sky130_fd_sc_hd__inv_2
X_49955_ _49955_/A _53167_/B _49955_/Y sky130_fd_sc_hd__nand2_4
X_45078_ _45075_/Y _45077_/Y _45063_/X _45078_/X sky130_fd_sc_hd__a21o_4
X_77987_ _77999_/A _77999_/B _78010_/A sky130_fd_sc_hd__xor2_4
X_48906_ _46240_/A _48384_/Y _48905_/Y _52275_/B sky130_fd_sc_hd__a21o_4
X_44029_ _64731_/A _60371_/A sky130_fd_sc_hd__buf_2
X_67740_ _67739_/X _86926_/Q _67740_/X sky130_fd_sc_hd__and2_4
X_79726_ _79702_/A _79701_/Y _79711_/X _79714_/Y _79726_/X sky130_fd_sc_hd__o22a_4
X_64952_ _64797_/X _83300_/Q _64772_/X _64951_/X _64953_/B sky130_fd_sc_hd__a211o_4
X_60075_ _60071_/X _60073_/Y _59969_/X _80091_/A _60074_/X _60075_/Y
+ sky130_fd_sc_hd__o32ai_4
X_76938_ _76939_/A _76938_/B _76938_/X sky130_fd_sc_hd__xor2_4
X_49886_ _49901_/A _53101_/B _49886_/Y sky130_fd_sc_hd__nand2_4
X_63903_ _63899_/Y _63903_/B _63901_/Y _63903_/D _63903_/X sky130_fd_sc_hd__and4_4
X_48837_ _48837_/A _48851_/A sky130_fd_sc_hd__buf_2
X_79657_ _84212_/Q _83260_/Q _79657_/X sky130_fd_sc_hd__xor2_4
X_67671_ _67312_/X _67671_/X sky130_fd_sc_hd__buf_2
X_64883_ _64883_/A _86263_/Q _64883_/X sky130_fd_sc_hd__and2_4
X_76869_ _81497_/Q _76867_/Y _76868_/X _76869_/Y sky130_fd_sc_hd__o21ai_4
X_69410_ _88031_/Q _69162_/X _69202_/X _69409_/X _69410_/X sky130_fd_sc_hd__a211o_4
X_66622_ _88401_/Q _66593_/X _66594_/X _66621_/X _66622_/X sky130_fd_sc_hd__a211o_4
X_78608_ _78608_/A _82678_/D _78608_/Y sky130_fd_sc_hd__nor2_4
X_63834_ _63800_/A _63800_/B _84292_/Q _63834_/Y sky130_fd_sc_hd__nor3_4
X_48768_ _48777_/A _48482_/B _48768_/Y sky130_fd_sc_hd__nand2_4
X_79588_ _79588_/A _79586_/A _79585_/Y _79588_/Y sky130_fd_sc_hd__nand3_4
X_69341_ _69302_/A _87780_/Q _69341_/X sky130_fd_sc_hd__and2_4
X_47719_ _72368_/A _47714_/X _47718_/Y _47719_/Y sky130_fd_sc_hd__o21ai_4
X_66553_ _44019_/A _66553_/X sky130_fd_sc_hd__buf_2
X_78539_ _78538_/X _78539_/Y sky130_fd_sc_hd__inv_2
X_63765_ _63765_/A _63380_/A _63765_/C _63765_/X sky130_fd_sc_hd__and3_4
X_48699_ _48697_/Y _48699_/B _48699_/Y sky130_fd_sc_hd__nand2_4
X_60977_ _60969_/X _60835_/X _84546_/Q _60977_/X sky130_fd_sc_hd__or3_4
X_65504_ _64829_/A _65504_/X sky130_fd_sc_hd__buf_2
X_50730_ _86145_/Q _50727_/X _50729_/Y _50730_/Y sky130_fd_sc_hd__o21ai_4
X_62716_ _61387_/X _62694_/B _62694_/C _62664_/D _62716_/Y sky130_fd_sc_hd__nand4_4
X_81550_ _80912_/CLK _81550_/D _76155_/B sky130_fd_sc_hd__dfxtp_4
X_69272_ _88041_/Q _69217_/X _69245_/X _69271_/X _69272_/X sky130_fd_sc_hd__a211o_4
X_66484_ _84114_/Q _66484_/Y sky130_fd_sc_hd__inv_2
X_63696_ _63696_/A _62162_/X _63696_/X sky130_fd_sc_hd__and2_4
X_80501_ _80487_/Y _80492_/Y _80500_/X _80501_/Y sky130_fd_sc_hd__o21ai_4
X_68223_ _68221_/X _67367_/Y _68207_/X _68222_/Y _68223_/X sky130_fd_sc_hd__a211o_4
X_65435_ _65449_/A _65294_/B _84201_/Q _65435_/X sky130_fd_sc_hd__and3_4
X_50661_ _50658_/Y _50609_/X _50660_/X _86159_/D sky130_fd_sc_hd__a21oi_4
X_62647_ _59450_/Y _60284_/A _62646_/Y _62647_/Y sky130_fd_sc_hd__o21ai_4
X_81481_ _81344_/CLK _81481_/D _76708_/A sky130_fd_sc_hd__dfxtp_4
X_52400_ _52602_/A _52400_/X sky130_fd_sc_hd__buf_2
X_83220_ _84487_/CLK _72603_/X _83220_/Q sky130_fd_sc_hd__dfxtp_4
X_80432_ _84759_/Q _84151_/Q _80432_/X sky130_fd_sc_hd__xor2_4
X_68154_ _82065_/D _68140_/X _68153_/X _84025_/D sky130_fd_sc_hd__a21bo_4
X_53380_ _53386_/A _47116_/A _53380_/Y sky130_fd_sc_hd__nand2_4
X_65366_ _65361_/X _65365_/X _65287_/X _65366_/X sky130_fd_sc_hd__a21o_4
X_50592_ _50580_/A _71989_/B _50592_/Y sky130_fd_sc_hd__nand2_4
X_62578_ _62577_/Y _59945_/Y _62948_/C _59931_/A _62578_/X sky130_fd_sc_hd__a2bb2o_4
X_67105_ _87869_/Q _67056_/X _67032_/X _67104_/X _67105_/X sky130_fd_sc_hd__a211o_4
X_52331_ _85844_/Q _52324_/X _52330_/Y _52331_/Y sky130_fd_sc_hd__o21ai_4
X_64317_ _64221_/A _64318_/D sky130_fd_sc_hd__buf_2
X_83151_ _86535_/CLK _83151_/D _83151_/Q sky130_fd_sc_hd__dfxtp_4
X_61529_ _61686_/A _61563_/B sky130_fd_sc_hd__buf_2
X_80363_ _80337_/Y _80353_/Y _80363_/Y sky130_fd_sc_hd__nor2_4
X_68085_ _68082_/X _68084_/X _68062_/X _68085_/Y sky130_fd_sc_hd__a21oi_4
X_65297_ _64656_/A _72123_/A sky130_fd_sc_hd__buf_2
X_82102_ _82343_/CLK _82114_/Q _82102_/Q sky130_fd_sc_hd__dfxtp_4
X_55050_ _55102_/A _55050_/X sky130_fd_sc_hd__buf_2
X_67036_ _66961_/X _86787_/Q _67036_/X sky130_fd_sc_hd__and2_4
X_52262_ _52262_/A _52262_/X sky130_fd_sc_hd__buf_2
X_64248_ _64248_/A _64248_/B _64248_/C _64248_/X sky130_fd_sc_hd__and3_4
X_83082_ _83184_/CLK _74362_/X _83082_/Q sky130_fd_sc_hd__dfxtp_4
X_80294_ _80293_/Y _80294_/B _80297_/A sky130_fd_sc_hd__nand2_4
X_54001_ _85525_/Q _53989_/X _54000_/Y _54001_/Y sky130_fd_sc_hd__o21ai_4
X_51213_ _86053_/Q _51209_/X _51212_/Y _51213_/Y sky130_fd_sc_hd__o21ai_4
X_86910_ _84538_/CLK _44924_/Y _64223_/B sky130_fd_sc_hd__dfxtp_4
X_82033_ _82005_/CLK _82033_/D _82001_/D sky130_fd_sc_hd__dfxtp_4
X_52193_ _52247_/A _52218_/C sky130_fd_sc_hd__buf_2
X_64179_ _64545_/B _64179_/B _64179_/C _64179_/D _64181_/C sky130_fd_sc_hd__nand4_4
X_87890_ _87995_/CLK _42384_/X _87890_/Q sky130_fd_sc_hd__dfxtp_4
X_51144_ _51130_/A _52837_/B _51144_/Y sky130_fd_sc_hd__nand2_4
X_86841_ _86841_/CLK _45939_/Y _86841_/Q sky130_fd_sc_hd__dfxtp_4
X_68987_ _68987_/A _74145_/A _68987_/X sky130_fd_sc_hd__and2_4
X_58740_ _58858_/A _58740_/X sky130_fd_sc_hd__buf_2
X_55952_ _44085_/C _56027_/C _55952_/X sky130_fd_sc_hd__and2_4
X_51075_ _51129_/A _51097_/A sky130_fd_sc_hd__buf_2
X_67938_ _68450_/A _67938_/X sky130_fd_sc_hd__buf_2
X_86772_ _86772_/CLK _46140_/X _43012_/B sky130_fd_sc_hd__dfxtp_4
X_83984_ _87671_/CLK _83984_/D _82632_/D sky130_fd_sc_hd__dfxtp_4
X_50026_ _50024_/Y _50003_/X _50025_/X _50026_/Y sky130_fd_sc_hd__a21oi_4
X_54903_ _54893_/X _54903_/B _54903_/Y sky130_fd_sc_hd__nand2_4
X_85723_ _84746_/CLK _85723_/D _85723_/Q sky130_fd_sc_hd__dfxtp_4
X_58671_ _58659_/A _86393_/Q _58671_/Y sky130_fd_sc_hd__nor2_4
X_82935_ _82933_/CLK _78287_/X _46371_/A sky130_fd_sc_hd__dfxtp_4
X_55883_ _44081_/X _56317_/C _55883_/X sky130_fd_sc_hd__and2_4
X_67869_ _67891_/A _86921_/Q _67869_/X sky130_fd_sc_hd__and2_4
X_57622_ _84967_/Q _57603_/X _57621_/Y _57622_/Y sky130_fd_sc_hd__o21ai_4
X_69608_ _69648_/A _42550_/Y _69608_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_9_460_0_CLK clkbuf_9_461_0_CLK/A clkbuf_9_460_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_54834_ _85369_/Q _54812_/X _54833_/Y _54834_/Y sky130_fd_sc_hd__o21ai_4
X_85654_ _85751_/CLK _85654_/D _85654_/Q sky130_fd_sc_hd__dfxtp_4
X_70880_ _70905_/A _70880_/B _70880_/C _70875_/X _70880_/Y sky130_fd_sc_hd__nand4_4
X_82866_ _82855_/CLK _78199_/B _82866_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_354_0_CLK clkbuf_9_177_0_CLK/X _86317_/CLK sky130_fd_sc_hd__clkbuf_1
X_84605_ _84606_/CLK _60531_/Y _79145_/A sky130_fd_sc_hd__dfxtp_4
X_57553_ _57552_/X _47967_/Y _57553_/Y sky130_fd_sc_hd__nand2_4
X_81817_ _81689_/CLK _81625_/Q _81817_/Q sky130_fd_sc_hd__dfxtp_4
X_69539_ _69080_/X _69082_/X _69500_/X _69539_/Y sky130_fd_sc_hd__a21oi_4
X_88373_ _87416_/CLK _88373_/D _88373_/Q sky130_fd_sc_hd__dfxtp_4
X_54765_ _54656_/X _54788_/B sky130_fd_sc_hd__buf_2
X_85585_ _86193_/CLK _85585_/D _85585_/Q sky130_fd_sc_hd__dfxtp_4
X_51977_ _51941_/A _50275_/B _51977_/Y sky130_fd_sc_hd__nand2_4
X_82797_ _82797_/CLK _82829_/Q _82797_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_984_0_CLK clkbuf_9_492_0_CLK/X _86498_/CLK sky130_fd_sc_hd__clkbuf_1
X_56504_ _56079_/X _56499_/X _56503_/Y _85171_/D sky130_fd_sc_hd__o21ai_4
X_87324_ _87577_/CLK _87324_/D _74097_/A sky130_fd_sc_hd__dfxtp_4
X_41730_ _41717_/X _81742_/Q _41729_/X _41730_/Y sky130_fd_sc_hd__o21ai_4
X_53716_ _52199_/A _53720_/B _53734_/C _53716_/X sky130_fd_sc_hd__and3_4
X_72550_ _72550_/A _72555_/B _72550_/C _72572_/B sky130_fd_sc_hd__nand3_4
X_84536_ _84531_/CLK _84536_/D _84536_/Q sky130_fd_sc_hd__dfxtp_4
X_50928_ _50957_/A _50928_/X sky130_fd_sc_hd__buf_2
X_57484_ _57484_/A _57225_/Y _57485_/C sky130_fd_sc_hd__nand2_4
X_81748_ _81514_/CLK _81748_/D _41699_/B sky130_fd_sc_hd__dfxtp_4
X_54696_ _54692_/Y _54694_/X _54695_/X _54696_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_475_0_CLK clkbuf_9_475_0_CLK/A clkbuf_9_475_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_59223_ _59218_/Y _59222_/Y _59165_/X _59223_/X sky130_fd_sc_hd__a21o_4
X_71501_ _58454_/Y _71486_/A _71500_/Y _83476_/D sky130_fd_sc_hd__o21ai_4
X_56435_ _56435_/A _56446_/A sky130_fd_sc_hd__buf_2
X_87255_ _87260_/CLK _87255_/D _69523_/B sky130_fd_sc_hd__dfxtp_4
X_53647_ _53656_/A _53647_/B _53647_/Y sky130_fd_sc_hd__nand2_4
X_41661_ _41661_/A _41660_/X _41661_/X sky130_fd_sc_hd__or2_4
X_72481_ _57697_/X _85954_/Q _72480_/X _72481_/Y sky130_fd_sc_hd__o21ai_4
X_84467_ _82452_/CLK _84467_/D _79135_/B sky130_fd_sc_hd__dfxtp_4
X_50859_ _86119_/Q _50856_/X _50858_/Y _50859_/Y sky130_fd_sc_hd__o21ai_4
X_81679_ _81259_/CLK _80065_/Y _76917_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_369_0_CLK clkbuf_9_184_0_CLK/X _83046_/CLK sky130_fd_sc_hd__clkbuf_1
X_43400_ _43399_/X _43375_/X _41473_/X _87440_/Q _43378_/X _43400_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74220_ _48122_/Y _74220_/B _74221_/B sky130_fd_sc_hd__xor2_4
X_86206_ _86490_/CLK _50413_/Y _86206_/Q sky130_fd_sc_hd__dfxtp_4
X_40612_ _40832_/A _40612_/X sky130_fd_sc_hd__buf_2
X_71432_ _71432_/A _71432_/B _70782_/A _71432_/D _71432_/X sky130_fd_sc_hd__and4_4
X_59154_ _59154_/A _86357_/Q _59154_/Y sky130_fd_sc_hd__nor2_4
X_83418_ _83414_/CLK _71667_/Y _58530_/A sky130_fd_sc_hd__dfxtp_4
X_44380_ _41782_/X _44377_/X _87138_/Q _44379_/X _87138_/D sky130_fd_sc_hd__a2bb2o_4
X_56366_ _56168_/X _56284_/X _56365_/Y _85219_/D sky130_fd_sc_hd__o21ai_4
X_41592_ _41591_/Y _41592_/X sky130_fd_sc_hd__buf_2
X_87186_ _83753_/CLK _87186_/D _87186_/Q sky130_fd_sc_hd__dfxtp_4
X_53578_ _85609_/Q _53540_/X _53577_/Y _53578_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_999_0_CLK clkbuf_9_499_0_CLK/X _86516_/CLK sky130_fd_sc_hd__clkbuf_1
X_84398_ _83242_/CLK _84398_/D _84398_/Q sky130_fd_sc_hd__dfxtp_4
X_58105_ _58610_/A _58105_/X sky130_fd_sc_hd__buf_2
X_43331_ _43316_/X _43319_/X _41277_/X _87477_/Q _43330_/X _43332_/A
+ sky130_fd_sc_hd__o32ai_4
X_55317_ _55317_/A _55317_/B _55317_/X sky130_fd_sc_hd__and2_4
X_74151_ _74080_/X _86216_/Q _74103_/X _74150_/X _74151_/X sky130_fd_sc_hd__a211o_4
X_86137_ _85529_/CLK _50770_/Y _86137_/Q sky130_fd_sc_hd__dfxtp_4
X_40543_ _40409_/X _40543_/X sky130_fd_sc_hd__buf_2
X_52529_ _52527_/Y _52496_/X _52528_/X _52529_/Y sky130_fd_sc_hd__a21oi_4
X_59085_ _59085_/A _59085_/X sky130_fd_sc_hd__buf_2
X_71363_ _71366_/A _71351_/X _71435_/C _71363_/D _71363_/X sky130_fd_sc_hd__and4_4
X_83349_ _83763_/CLK _83349_/D _83349_/Q sky130_fd_sc_hd__dfxtp_4
X_56297_ _56020_/X _56290_/X _56296_/Y _56297_/Y sky130_fd_sc_hd__o21ai_4
X_73102_ _73100_/X _73101_/Y _72970_/X _73102_/Y sky130_fd_sc_hd__a21oi_4
X_46050_ _46046_/X _46032_/X _41519_/X _86794_/Q _46047_/X _46051_/A
+ sky130_fd_sc_hd__o32ai_4
X_58036_ _58032_/Y _58034_/Y _58035_/X _58036_/X sky130_fd_sc_hd__a21o_4
X_70314_ _70303_/X _74808_/B _70313_/X _70314_/X sky130_fd_sc_hd__a21o_4
X_55248_ _55135_/A _55248_/B _55248_/X sky130_fd_sc_hd__and2_4
X_43262_ _43261_/Y _43262_/Y sky130_fd_sc_hd__inv_2
X_74082_ _74080_/X _86219_/Q _73446_/X _74081_/X _74082_/X sky130_fd_sc_hd__a211o_4
X_86068_ _85748_/CLK _86068_/D _86068_/Q sky130_fd_sc_hd__dfxtp_4
X_40474_ _40473_/X _40474_/X sky130_fd_sc_hd__buf_2
X_71294_ _71185_/B _71303_/B sky130_fd_sc_hd__buf_2
X_45001_ _55931_/B _44982_/X _44959_/X _45001_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_10_922_0_CLK clkbuf_9_461_0_CLK/X _87070_/CLK sky130_fd_sc_hd__clkbuf_1
X_42213_ _42212_/Y _87978_/D sky130_fd_sc_hd__inv_2
X_77910_ _77909_/X _77910_/Y sky130_fd_sc_hd__inv_2
X_73033_ _73033_/A _73372_/B _73033_/Y sky130_fd_sc_hd__nor2_4
X_85019_ _85013_/CLK _57393_/Y _57392_/B sky130_fd_sc_hd__dfxtp_4
X_70245_ _70127_/X _70246_/A sky130_fd_sc_hd__buf_2
X_43193_ _43031_/X _43125_/X _40903_/X _43192_/Y _43142_/X _43193_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55179_ _55171_/X _55178_/X _83748_/Q _55179_/X sky130_fd_sc_hd__a21o_4
X_78890_ _82636_/Q _78890_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_9_413_0_CLK clkbuf_9_413_0_CLK/A clkbuf_9_413_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_42144_ _42143_/Y _88014_/D sky130_fd_sc_hd__inv_2
X_77841_ _77841_/A _77840_/Y _77841_/Y sky130_fd_sc_hd__nand2_4
X_70176_ _70183_/A _70183_/B _70176_/C _70183_/D _70176_/X sky130_fd_sc_hd__and4_4
X_59987_ _62609_/D _59987_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_307_0_CLK clkbuf_9_153_0_CLK/X _83367_/CLK sky130_fd_sc_hd__clkbuf_1
X_49740_ _49737_/Y _49732_/X _49739_/X _86332_/D sky130_fd_sc_hd__a21oi_4
X_46952_ _46952_/A _52771_/D sky130_fd_sc_hd__buf_2
X_42075_ _40968_/X _42072_/X _88045_/Q _42073_/X _42075_/X sky130_fd_sc_hd__a2bb2o_4
X_58938_ _58796_/X _86084_/Q _58937_/X _58938_/Y sky130_fd_sc_hd__o21ai_4
X_77772_ _77763_/Y _77766_/Y _77771_/Y _77773_/B sky130_fd_sc_hd__o21ai_4
X_74984_ _74981_/Y _74983_/Y _74985_/B sky130_fd_sc_hd__xor2_4
Xclkbuf_10_937_0_CLK clkbuf_9_468_0_CLK/X _88326_/CLK sky130_fd_sc_hd__clkbuf_1
X_79511_ _79500_/Y _79504_/B _79512_/B sky130_fd_sc_hd__or2_4
X_41026_ _41026_/A _41091_/B _41026_/X sky130_fd_sc_hd__or2_4
X_45903_ _44128_/X _72973_/B sky130_fd_sc_hd__buf_2
X_76723_ _76703_/Y _76719_/A _76722_/X _76723_/Y sky130_fd_sc_hd__a21oi_4
X_49671_ _49661_/X _52885_/B _49671_/Y sky130_fd_sc_hd__nand2_4
X_73935_ _73924_/Y _73935_/B _73937_/A sky130_fd_sc_hd__xor2_4
X_46883_ _54423_/D _52730_/D sky130_fd_sc_hd__buf_2
X_58869_ _58864_/X _58866_/Y _58867_/Y _58766_/X _58868_/X _58869_/X
+ sky130_fd_sc_hd__o32a_4
Xclkbuf_9_428_0_CLK clkbuf_9_429_0_CLK/A clkbuf_9_428_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_48622_ _47872_/A _48623_/A sky130_fd_sc_hd__buf_2
X_60900_ _60888_/Y _60910_/B sky130_fd_sc_hd__buf_2
X_79442_ _79439_/Y _79422_/Y _79441_/X _79442_/Y sky130_fd_sc_hd__o21ai_4
X_45834_ _63324_/B _61666_/A sky130_fd_sc_hd__buf_2
X_76654_ _76651_/Y _76653_/Y _76648_/A _76664_/A sky130_fd_sc_hd__a21oi_4
X_61880_ _61869_/X _61872_/X _61879_/Y _84744_/Q _61815_/X _61880_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73866_ _73864_/X _73866_/B _73866_/C _73866_/Y sky130_fd_sc_hd__nand3_4
X_75605_ _81110_/Q _75605_/B _80774_/D sky130_fd_sc_hd__xor2_4
X_48553_ _86512_/Q _48548_/X _48552_/Y _48553_/Y sky130_fd_sc_hd__o21ai_4
X_72817_ _72816_/X _72817_/B _72817_/X sky130_fd_sc_hd__and2_4
X_60831_ _60830_/X _84556_/D sky130_fd_sc_hd__inv_2
X_79373_ _79373_/A _79373_/B _79373_/Y sky130_fd_sc_hd__xnor2_4
X_45765_ _45765_/A _45765_/X sky130_fd_sc_hd__buf_2
X_76585_ _76541_/B _76559_/Y _76541_/A _76560_/Y _76585_/Y sky130_fd_sc_hd__nand4_4
X_42977_ _42970_/X _42971_/X _40446_/X _87622_/Q _42976_/X _42978_/A
+ sky130_fd_sc_hd__o32ai_4
X_73797_ _73797_/A _73701_/B _73797_/Y sky130_fd_sc_hd__nor2_4
X_47504_ _47500_/Y _47462_/X _47503_/X _47504_/Y sky130_fd_sc_hd__a21oi_4
X_78324_ _78317_/X _78324_/B _78335_/A _78325_/B sky130_fd_sc_hd__nand3_4
X_44716_ _44716_/A _86990_/D sky130_fd_sc_hd__inv_2
X_63550_ _63512_/A _84954_/Q _63537_/C _63550_/X sky130_fd_sc_hd__and3_4
X_75536_ _75536_/A _75523_/X _75503_/Y _75524_/Y _75536_/X sky130_fd_sc_hd__and4_4
X_41928_ _42000_/A _41928_/X sky130_fd_sc_hd__buf_2
X_48484_ _48484_/A _48485_/A sky130_fd_sc_hd__inv_2
X_60762_ _60739_/X _60759_/Y _60722_/Y _60726_/Y _60761_/Y _84573_/D
+ sky130_fd_sc_hd__a41oi_4
X_72748_ _72929_/A _65423_/B _72748_/X sky130_fd_sc_hd__and2_4
X_45696_ _82990_/Q _45697_/A sky130_fd_sc_hd__inv_2
X_62501_ _62501_/A _62501_/X sky130_fd_sc_hd__buf_2
X_47435_ _46610_/A _49406_/A sky130_fd_sc_hd__buf_2
X_78255_ _78239_/B _78252_/X _78254_/Y _78256_/B sky130_fd_sc_hd__a21oi_4
X_44647_ _44647_/A _44647_/Y sky130_fd_sc_hd__inv_2
X_75467_ _75467_/A _75467_/Y sky130_fd_sc_hd__inv_2
X_63481_ _63434_/X _63472_/X _63473_/X _63477_/X _63480_/Y _63481_/Y
+ sky130_fd_sc_hd__o41ai_4
X_41859_ _40542_/X _48226_/A _67290_/B _40599_/A _88117_/D sky130_fd_sc_hd__a2bb2o_4
X_72679_ _72683_/A _72683_/B _55392_/A _72679_/Y sky130_fd_sc_hd__nand3_4
X_60693_ _63478_/A _63389_/B sky130_fd_sc_hd__buf_2
X_65220_ _84210_/Q _65221_/C sky130_fd_sc_hd__inv_2
X_77206_ _77201_/Y _77177_/B _77205_/X _77207_/B sky130_fd_sc_hd__o21ai_4
X_74418_ _74413_/X _73073_/A _74418_/Y sky130_fd_sc_hd__nand2_4
X_62432_ _62448_/A _58533_/A _62375_/C _62432_/Y sky130_fd_sc_hd__nand3_4
X_47366_ _49504_/A _47556_/A sky130_fd_sc_hd__buf_2
X_78186_ _78193_/B _78174_/B _78186_/Y sky130_fd_sc_hd__nand2_4
X_44578_ _44554_/X _44555_/X _40889_/Y _44577_/Y _44557_/X _87048_/D
+ sky130_fd_sc_hd__o32ai_4
X_75398_ _75378_/Y _75375_/Y _75376_/Y _75399_/A sky130_fd_sc_hd__o21a_4
X_49105_ _48898_/A _49117_/A sky130_fd_sc_hd__buf_2
X_46317_ _46317_/A _46505_/A sky130_fd_sc_hd__buf_2
X_65151_ _65673_/A _65206_/A sky130_fd_sc_hd__buf_2
X_77137_ _77143_/B _81916_/Q _77136_/Y _77138_/B sky130_fd_sc_hd__a21oi_4
X_43529_ _43518_/X _43523_/X _40395_/X _87374_/Q _43528_/X _43529_/Y
+ sky130_fd_sc_hd__o32ai_4
X_62363_ _59950_/C _62363_/X sky130_fd_sc_hd__buf_2
X_74349_ _74351_/A _74342_/X _56117_/B _74349_/Y sky130_fd_sc_hd__nand3_4
X_47297_ _47297_/A _47297_/Y sky130_fd_sc_hd__inv_2
X_64102_ _58277_/A _64102_/B _64102_/Y sky130_fd_sc_hd__nor2_4
X_61314_ _72550_/C _72607_/B sky130_fd_sc_hd__buf_2
X_49036_ _49007_/A _52338_/B _49036_/Y sky130_fd_sc_hd__nand2_4
X_46248_ _47002_/A _46249_/A sky130_fd_sc_hd__buf_2
X_65082_ _64904_/A _85839_/Q _65082_/X sky130_fd_sc_hd__and2_4
X_77068_ _77068_/A _77068_/B _77068_/Y sky130_fd_sc_hd__nand2_4
X_62294_ _62609_/D _62632_/C sky130_fd_sc_hd__buf_2
X_64033_ _63585_/B _64095_/B _64050_/C _64033_/D _64033_/Y sky130_fd_sc_hd__nand4_4
X_68910_ _69001_/A _68910_/B _68910_/Y sky130_fd_sc_hd__nor2_4
X_76019_ _76009_/Y _76019_/B _76023_/A sky130_fd_sc_hd__nand2_4
X_61245_ _61262_/A _61250_/B _75901_/A _61245_/Y sky130_fd_sc_hd__nor3_4
X_46179_ _46178_/X _46179_/X sky130_fd_sc_hd__buf_2
X_69890_ _69887_/X _69889_/X _69890_/Y sky130_fd_sc_hd__nand2_4
X_68841_ _57804_/A _42509_/Y _68841_/Y sky130_fd_sc_hd__nor2_4
X_61176_ _61202_/B _61176_/B _61176_/Y sky130_fd_sc_hd__nand2_4
X_60127_ _59943_/A _59973_/A _62269_/A sky130_fd_sc_hd__and2_4
X_49938_ _49925_/X _49915_/X _49953_/C _53151_/D _49938_/X sky130_fd_sc_hd__and4_4
X_68772_ _87491_/Q _68472_/A _68545_/X _68771_/X _68772_/X sky130_fd_sc_hd__a211o_4
X_65984_ _65984_/A _66062_/B sky130_fd_sc_hd__buf_2
X_67723_ _68644_/A _67790_/A sky130_fd_sc_hd__buf_2
X_79709_ _79703_/Y _79708_/Y _79709_/X sky130_fd_sc_hd__xor2_4
X_64935_ _64877_/X _86453_/Q _64935_/X sky130_fd_sc_hd__and2_4
X_60058_ _60528_/A _60058_/B _60058_/Y sky130_fd_sc_hd__nor2_4
X_49869_ _58116_/B _49853_/X _49868_/Y _49869_/Y sky130_fd_sc_hd__o21ai_4
X_80981_ _80931_/CLK _75748_/X _80937_/D sky130_fd_sc_hd__dfxtp_4
X_51900_ _51900_/A _51900_/X sky130_fd_sc_hd__buf_2
X_82720_ _82624_/CLK _82720_/D _82720_/Q sky130_fd_sc_hd__dfxtp_4
X_67654_ _67582_/A _67654_/B _67654_/X sky130_fd_sc_hd__and2_4
X_52880_ _52877_/Y _52865_/X _52879_/X _52880_/Y sky130_fd_sc_hd__a21oi_4
X_64866_ _64809_/X _86744_/Q _64864_/X _64865_/X _64866_/X sky130_fd_sc_hd__a211o_4
X_66605_ _68389_/A _66606_/A sky130_fd_sc_hd__buf_2
X_51831_ _85938_/Q _51817_/X _51830_/Y _51831_/Y sky130_fd_sc_hd__o21ai_4
X_63817_ _63800_/A _63800_/B _80206_/B _63817_/Y sky130_fd_sc_hd__nor3_4
X_82651_ _84003_/CLK _84003_/Q _82651_/Q sky130_fd_sc_hd__dfxtp_4
X_67585_ _67466_/X _67585_/X sky130_fd_sc_hd__buf_2
X_64797_ _64797_/A _64797_/X sky130_fd_sc_hd__buf_2
X_81602_ _81794_/CLK _81602_/D _81602_/Q sky130_fd_sc_hd__dfxtp_4
X_69324_ _69320_/X _69323_/X _69324_/Y sky130_fd_sc_hd__nand2_4
X_54550_ _54547_/Y _54530_/X _54549_/X _85422_/D sky130_fd_sc_hd__a21oi_4
X_66536_ _87955_/Q _66529_/X _66531_/X _66535_/X _66536_/X sky130_fd_sc_hd__a211o_4
X_85370_ _83275_/CLK _85370_/D _85370_/Q sky130_fd_sc_hd__dfxtp_4
X_51762_ _51759_/Y _51391_/X _51761_/X _51762_/Y sky130_fd_sc_hd__a21oi_4
X_63748_ _60930_/A _63749_/A sky130_fd_sc_hd__buf_2
X_82582_ _82711_/CLK _82614_/Q _78228_/A sky130_fd_sc_hd__dfxtp_4
X_53501_ _53478_/A _53501_/B _53501_/Y sky130_fd_sc_hd__nand2_4
X_84321_ _84321_/CLK _63470_/Y _84321_/Q sky130_fd_sc_hd__dfxtp_4
X_50713_ _86148_/Q _50706_/X _50712_/Y _50713_/Y sky130_fd_sc_hd__o21ai_4
X_81533_ _81703_/CLK _81545_/Q _81533_/Q sky130_fd_sc_hd__dfxtp_4
X_69255_ _69255_/A _69254_/X _69255_/Y sky130_fd_sc_hd__nand2_4
X_54481_ _54481_/A _54483_/A sky130_fd_sc_hd__buf_2
X_66467_ _60110_/X _65126_/Y _66466_/Y _66467_/Y sky130_fd_sc_hd__o21ai_4
X_51693_ _51639_/A _51693_/X sky130_fd_sc_hd__buf_2
X_63679_ _63578_/A _63679_/X sky130_fd_sc_hd__buf_2
X_56220_ _56060_/X _56210_/X _56219_/Y _85271_/D sky130_fd_sc_hd__o21ai_4
X_68206_ _82052_/D _68200_/X _68205_/X _68206_/X sky130_fd_sc_hd__a21bo_4
X_87040_ _87068_/CLK _44601_/Y _87040_/Q sky130_fd_sc_hd__dfxtp_4
X_53432_ _47832_/X _54194_/A sky130_fd_sc_hd__buf_2
X_65418_ _65342_/X _86722_/Q _65391_/X _65417_/X _65418_/X sky130_fd_sc_hd__a211o_4
X_84252_ _83766_/CLK _64372_/X _79742_/B sky130_fd_sc_hd__dfxtp_4
X_50644_ _50577_/A _50644_/X sky130_fd_sc_hd__buf_2
X_81464_ _81431_/CLK _81464_/D _81464_/Q sky130_fd_sc_hd__dfxtp_4
X_69186_ _69181_/X _69186_/B _69186_/Y sky130_fd_sc_hd__nand2_4
X_66398_ _66010_/X _66397_/X _66013_/X _66398_/Y sky130_fd_sc_hd__nand3_4
X_83203_ _83843_/CLK _83203_/D _83203_/Q sky130_fd_sc_hd__dfxtp_4
X_56151_ _56142_/X _56148_/X _56150_/Y _56151_/Y sky130_fd_sc_hd__o21ai_4
X_80415_ _80411_/Y _80414_/Y _80425_/B sky130_fd_sc_hd__xor2_4
X_68137_ _66866_/X _66870_/X _68133_/X _68137_/Y sky130_fd_sc_hd__a21oi_4
X_53363_ _53361_/Y _53355_/X _53362_/X _85648_/D sky130_fd_sc_hd__a21oi_4
X_65349_ _65346_/Y _65347_/X _65348_/X _84205_/D sky130_fd_sc_hd__a21o_4
X_84183_ _84194_/CLK _84183_/D _65713_/C sky130_fd_sc_hd__dfxtp_4
X_50575_ _50575_/A _48912_/B _50575_/Y sky130_fd_sc_hd__nand2_4
X_81395_ _83932_/CLK _83931_/Q _81395_/Q sky130_fd_sc_hd__dfxtp_4
X_55102_ _55102_/A _55102_/X sky130_fd_sc_hd__buf_2
X_52314_ _52262_/A _52314_/X sky130_fd_sc_hd__buf_2
X_83134_ _84980_/CLK _73841_/Y _83134_/Q sky130_fd_sc_hd__dfxtp_4
X_80346_ _80343_/X _80344_/X _80360_/B _80350_/B sky130_fd_sc_hd__nand3_4
X_56082_ _56142_/A _56082_/X sky130_fd_sc_hd__buf_2
X_68068_ _87956_/Q _68066_/X _67997_/X _68067_/X _68068_/X sky130_fd_sc_hd__a211o_4
X_53294_ _53291_/Y _53272_/X _53293_/X _53294_/Y sky130_fd_sc_hd__a21oi_4
X_55033_ _55037_/A _54867_/B _55033_/Y sky130_fd_sc_hd__nand2_4
X_59910_ _59909_/Y _59910_/X sky130_fd_sc_hd__buf_2
X_67019_ _66972_/X _87616_/Q _67019_/X sky130_fd_sc_hd__and2_4
X_52245_ _52250_/A _48684_/B _52245_/Y sky130_fd_sc_hd__nand2_4
X_83065_ _85581_/CLK _74446_/Y _83065_/Q sky130_fd_sc_hd__dfxtp_4
X_87942_ _88387_/CLK _87942_/D _87942_/Q sky130_fd_sc_hd__dfxtp_4
X_80277_ _80276_/Y _80277_/B _80280_/B sky130_fd_sc_hd__nand2_4
X_70030_ _69739_/X _69741_/X _70001_/X _70030_/Y sky130_fd_sc_hd__a21oi_4
X_82016_ _82604_/CLK _82016_/D _77222_/A sky130_fd_sc_hd__dfxtp_4
X_59841_ _59825_/B _59841_/X sky130_fd_sc_hd__buf_2
X_52176_ _52174_/Y _52170_/X _52175_/X _85874_/D sky130_fd_sc_hd__a21oi_4
X_87873_ _88387_/CLK _42421_/Y _87873_/Q sky130_fd_sc_hd__dfxtp_4
X_51127_ _50991_/A _51128_/A sky130_fd_sc_hd__buf_2
X_86824_ _86824_/CLK _86824_/D _86824_/Q sky130_fd_sc_hd__dfxtp_4
X_59772_ _59772_/A _59771_/X _80517_/A _59772_/Y sky130_fd_sc_hd__nor3_4
X_56984_ _56682_/X _57149_/C sky130_fd_sc_hd__buf_2
Xclkbuf_10_60_0_CLK clkbuf_9_30_0_CLK/X _85005_/CLK sky130_fd_sc_hd__clkbuf_1
X_58723_ _58631_/X _58720_/Y _58722_/Y _58650_/X _58636_/X _58723_/X
+ sky130_fd_sc_hd__o32a_4
X_51058_ _51058_/A _52748_/B _51058_/Y sky130_fd_sc_hd__nand2_4
X_55935_ _83035_/Q _55619_/A _44102_/A _55934_/X _55936_/B sky130_fd_sc_hd__a211o_4
X_86755_ _84407_/CLK _46232_/Y _86755_/Q sky130_fd_sc_hd__dfxtp_4
X_71981_ _71957_/A _48931_/A _71981_/Y sky130_fd_sc_hd__nand2_4
X_83967_ _83967_/CLK _83967_/D _83967_/Q sky130_fd_sc_hd__dfxtp_4
X_50009_ _49930_/X _50025_/C sky130_fd_sc_hd__buf_2
X_42900_ _42962_/A _42900_/X sky130_fd_sc_hd__buf_2
X_73720_ _73367_/A _73720_/X sky130_fd_sc_hd__buf_2
X_85706_ _85704_/CLK _53053_/Y _85706_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_105_0_CLK clkbuf_6_52_0_CLK/X clkbuf_8_211_0_CLK/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_293_0_CLK clkbuf_9_146_0_CLK/X _83464_/CLK sky130_fd_sc_hd__clkbuf_1
X_70932_ _71115_/C _70959_/B sky130_fd_sc_hd__buf_2
X_58654_ _58641_/X _85946_/Q _58109_/X _58654_/X sky130_fd_sc_hd__o21a_4
X_82918_ _81198_/CLK _78160_/X _82918_/Q sky130_fd_sc_hd__dfxtp_4
X_43880_ _43869_/X _43880_/X sky130_fd_sc_hd__buf_2
X_55866_ _85268_/Q _55505_/X _55506_/X _55865_/X _55866_/X sky130_fd_sc_hd__a211o_4
X_86686_ _86686_/CLK _86686_/D _59030_/A sky130_fd_sc_hd__dfxtp_4
X_83898_ _82299_/CLK _69775_/X _83898_/Q sky130_fd_sc_hd__dfxtp_4
X_57605_ _57630_/A _57605_/B _57605_/Y sky130_fd_sc_hd__nand2_4
X_42831_ _42680_/A _42832_/A sky130_fd_sc_hd__buf_2
X_54817_ _54815_/Y _54802_/X _54816_/X _85373_/D sky130_fd_sc_hd__a21oi_4
X_73651_ _68465_/B _73250_/X _73344_/X _73650_/Y _73651_/X sky130_fd_sc_hd__a211o_4
X_85637_ _85635_/CLK _85637_/D _85637_/Q sky130_fd_sc_hd__dfxtp_4
X_70863_ _70863_/A _71088_/C _70863_/C _70869_/D _70863_/Y sky130_fd_sc_hd__nand4_4
X_58585_ _58696_/A _58585_/X sky130_fd_sc_hd__buf_2
X_82849_ _82740_/CLK _82849_/D _82849_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_75_0_CLK clkbuf_9_37_0_CLK/X _86882_/CLK sky130_fd_sc_hd__clkbuf_1
X_55797_ _55761_/A _56124_/C _55797_/X sky130_fd_sc_hd__and2_4
X_72602_ _72602_/A _72575_/A _72602_/X sky130_fd_sc_hd__and2_4
X_45550_ _55520_/B _45516_/X _45548_/X _45549_/Y _45550_/X sky130_fd_sc_hd__a211o_4
X_57536_ _57534_/Y _57515_/X _57535_/Y _84984_/D sky130_fd_sc_hd__a21boi_4
X_76370_ _76369_/B _76368_/Y _76369_/A _76370_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_8_221_0_CLK clkbuf_8_221_0_CLK/A clkbuf_9_443_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_88356_ _82538_/CLK _88356_/D _68750_/B sky130_fd_sc_hd__dfxtp_4
X_54748_ _54748_/A _54755_/B _54748_/C _54748_/D _54748_/X sky130_fd_sc_hd__and4_4
X_42762_ _42762_/A _42762_/Y sky130_fd_sc_hd__inv_2
X_73582_ _73582_/A _73581_/Y _73582_/Y sky130_fd_sc_hd__nand2_4
X_85568_ _83307_/CLK _53790_/Y _85568_/Q sky130_fd_sc_hd__dfxtp_4
X_70794_ _70772_/A _70794_/X sky130_fd_sc_hd__buf_2
X_44501_ _41249_/Y _44474_/X _87078_/Q _44475_/X _87078_/D sky130_fd_sc_hd__a2bb2o_4
X_75321_ _75320_/Y _75321_/Y sky130_fd_sc_hd__inv_2
X_87307_ _83158_/CLK _87307_/D _87307_/Q sky130_fd_sc_hd__dfxtp_4
X_41713_ _82897_/Q _41660_/X _41713_/X sky130_fd_sc_hd__or2_4
X_72533_ _72533_/A _72527_/Y _72532_/X _83239_/D sky130_fd_sc_hd__nand3_4
X_84519_ _84508_/CLK _84519_/D _61132_/C sky130_fd_sc_hd__dfxtp_4
X_45481_ _45479_/Y _45480_/Y _44939_/B _45481_/X sky130_fd_sc_hd__o21a_4
X_57467_ _57466_/Y _84999_/D sky130_fd_sc_hd__inv_2
X_42693_ _41093_/X _42679_/X _69521_/B _42681_/X _42693_/X sky130_fd_sc_hd__a2bb2o_4
X_88287_ _87022_/CLK _88287_/D _69415_/B sky130_fd_sc_hd__dfxtp_4
X_54679_ _85398_/Q _54676_/X _54678_/Y _54679_/Y sky130_fd_sc_hd__o21ai_4
X_85499_ _85499_/CLK _85499_/D _85499_/Q sky130_fd_sc_hd__dfxtp_4
X_47220_ _83393_/Q _47221_/A sky130_fd_sc_hd__inv_2
X_59206_ _59160_/X _85648_/Q _59205_/X _59206_/X sky130_fd_sc_hd__o21a_4
X_78040_ _77907_/Y _81942_/D sky130_fd_sc_hd__inv_2
X_44432_ _44454_/A _44432_/X sky130_fd_sc_hd__buf_2
X_56418_ _56418_/A _56418_/B _85201_/Q _56418_/Y sky130_fd_sc_hd__nand3_4
X_75252_ _75239_/A _80986_/Q _75252_/Y sky130_fd_sc_hd__nand2_4
X_41644_ _41643_/X _41638_/X _67385_/B _41639_/X _41644_/X sky130_fd_sc_hd__a2bb2o_4
X_87238_ _88012_/CLK _43844_/X _87238_/Q sky130_fd_sc_hd__dfxtp_4
X_72464_ _79549_/B _72358_/X _72460_/X _72463_/X _83252_/D sky130_fd_sc_hd__a22oi_4
X_57398_ _56613_/X _57391_/Y _57397_/Y _85017_/D sky130_fd_sc_hd__a21oi_4
X_74203_ _70129_/B _74139_/X _74202_/Y _74203_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_8_236_0_CLK clkbuf_8_237_0_CLK/A clkbuf_8_236_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_59137_ _59121_/X _85430_/Q _59136_/X _59137_/Y sky130_fd_sc_hd__o21ai_4
X_47151_ _86665_/Q _47145_/X _47150_/Y _47151_/Y sky130_fd_sc_hd__o21ai_4
X_71415_ _71342_/B _71450_/C sky130_fd_sc_hd__buf_2
X_44363_ _46298_/A _44363_/X sky130_fd_sc_hd__buf_2
X_56349_ _56134_/X _56337_/X _56348_/Y _85226_/D sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_231_0_CLK clkbuf_9_115_0_CLK/X _84441_/CLK sky130_fd_sc_hd__clkbuf_1
X_75183_ _80777_/Q _81033_/D _75183_/X sky130_fd_sc_hd__xor2_4
X_87169_ _87169_/CLK _87169_/D _87169_/Q sky130_fd_sc_hd__dfxtp_4
X_41575_ _41540_/X _41541_/X _41574_/X _67100_/B _41537_/X _41576_/A
+ sky130_fd_sc_hd__o32ai_4
X_72395_ _57712_/X _85322_/Q _72324_/X _72395_/X sky130_fd_sc_hd__o21a_4
X_46102_ _45955_/X _58981_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_861_0_CLK clkbuf_9_430_0_CLK/X _85815_/CLK sky130_fd_sc_hd__clkbuf_1
X_43314_ _43314_/A _87486_/D sky130_fd_sc_hd__inv_2
X_74134_ _74134_/A _74133_/X _74135_/B sky130_fd_sc_hd__nand2_4
X_40526_ _82310_/Q _40467_/B _40526_/X sky130_fd_sc_hd__or2_4
X_47082_ _46941_/A _47082_/X sky130_fd_sc_hd__buf_2
X_59068_ _59068_/A _59068_/B _59068_/Y sky130_fd_sc_hd__nor2_4
X_71346_ _71418_/B _71504_/C sky130_fd_sc_hd__buf_2
X_44294_ _44216_/X _44217_/X _45950_/A _44268_/A _44294_/X sky130_fd_sc_hd__a211o_4
X_79991_ _79980_/A _79963_/Y _79980_/B _79991_/Y sky130_fd_sc_hd__a21boi_4
Xclkbuf_10_13_0_CLK clkbuf_9_6_0_CLK/X _85184_/CLK sky130_fd_sc_hd__clkbuf_1
X_46033_ _46013_/X _46032_/X _41472_/X _86803_/Q _46014_/X _46034_/A
+ sky130_fd_sc_hd__o32ai_4
X_58019_ _58017_/X _85388_/Q _58018_/X _58019_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_352_0_CLK clkbuf_8_176_0_CLK/X clkbuf_9_352_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_43245_ _43241_/X _43244_/X _41045_/X _87520_/Q _43232_/X _43246_/A
+ sky130_fd_sc_hd__o32ai_4
X_74065_ _74065_/A _74065_/B _74066_/B sky130_fd_sc_hd__nand2_4
X_78942_ _78942_/A _78953_/A _78946_/A sky130_fd_sc_hd__xor2_4
X_40457_ _82322_/Q _40907_/B _40457_/X sky130_fd_sc_hd__or2_4
X_71277_ _53200_/B _71265_/X _71276_/Y _83550_/D sky130_fd_sc_hd__o21ai_4
X_61030_ _61030_/A _60966_/A _61030_/Y sky130_fd_sc_hd__nand2_4
X_73016_ _72816_/X _73016_/B _73016_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_246_0_CLK clkbuf_9_123_0_CLK/X _84564_/CLK sky130_fd_sc_hd__clkbuf_1
X_70228_ _70224_/X _83830_/Q _70227_/X _83830_/D sky130_fd_sc_hd__a21o_4
X_43176_ _43175_/X _53900_/A sky130_fd_sc_hd__buf_2
X_78873_ _78866_/A _78868_/A _78873_/Y sky130_fd_sc_hd__nor2_4
X_40388_ _40387_/X _40342_/X _88400_/Q _40355_/X _40388_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_10_876_0_CLK clkbuf_9_438_0_CLK/X _86436_/CLK sky130_fd_sc_hd__clkbuf_1
X_42127_ _41093_/X _42125_/X _88023_/Q _42126_/X _42127_/X sky130_fd_sc_hd__a2bb2o_4
X_77824_ _82156_/Q _77824_/B _82124_/D sky130_fd_sc_hd__xor2_4
Xclkbuf_10_28_0_CLK clkbuf_9_14_0_CLK/X _85156_/CLK sky130_fd_sc_hd__clkbuf_1
X_70159_ _70127_/X _70348_/A sky130_fd_sc_hd__buf_2
X_47984_ _47981_/X _47984_/B _47984_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_367_0_CLK clkbuf_9_367_0_CLK/A clkbuf_9_367_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_49723_ _49641_/A _49724_/B sky130_fd_sc_hd__buf_2
X_46935_ _46931_/Y _46891_/X _46934_/X _46935_/Y sky130_fd_sc_hd__a21oi_4
X_42058_ _42035_/X _42049_/X _40921_/X _42057_/Y _42037_/X _88054_/D
+ sky130_fd_sc_hd__o32ai_4
X_77755_ _82053_/Q _77764_/B sky130_fd_sc_hd__inv_2
X_74967_ _74963_/B _74971_/A _74966_/Y _74968_/B sky130_fd_sc_hd__a21boi_4
X_62981_ _62927_/A _62664_/B _62174_/X _62981_/Y sky130_fd_sc_hd__nand3_4
X_64720_ _64714_/X _86173_/Q _64716_/X _64719_/X _64720_/X sky130_fd_sc_hd__a211o_4
X_41009_ _41009_/A _41009_/X sky130_fd_sc_hd__buf_2
X_76706_ _76706_/A _81448_/D _81544_/D sky130_fd_sc_hd__xor2_4
X_49654_ _49638_/A _52869_/B _49654_/Y sky130_fd_sc_hd__nand2_4
X_61932_ _57672_/X _61902_/X _61916_/X _61870_/X _61931_/X _61932_/X
+ sky130_fd_sc_hd__a41o_4
X_73918_ _42499_/A _72829_/X _73918_/Y sky130_fd_sc_hd__nor2_4
X_46866_ _82951_/Q _46866_/Y sky130_fd_sc_hd__inv_2
X_77686_ _77688_/A _77686_/Y sky130_fd_sc_hd__inv_2
X_74898_ _74872_/Y _74897_/X _74904_/A sky130_fd_sc_hd__nand2_4
X_48605_ _86507_/Q _48536_/X _48604_/Y _48605_/Y sky130_fd_sc_hd__o21ai_4
X_79425_ _79415_/A _79414_/X _79424_/Y _79429_/A sky130_fd_sc_hd__a21boi_4
X_45817_ _74694_/B _45832_/B _45817_/Y sky130_fd_sc_hd__nand2_4
X_64651_ _64676_/A _85855_/Q _64651_/X sky130_fd_sc_hd__and2_4
X_76637_ _81537_/D _76637_/B _76637_/X sky130_fd_sc_hd__xor2_4
X_49585_ _49580_/X _52799_/B _49585_/Y sky130_fd_sc_hd__nand2_4
X_61863_ _61863_/A _61857_/Y _61860_/Y _61862_/Y _61863_/Y sky130_fd_sc_hd__nand4_4
X_73849_ _86995_/Q _73776_/X _73848_/X _73866_/C sky130_fd_sc_hd__o21ai_4
X_46797_ _58807_/A _46767_/X _46796_/Y _46797_/Y sky130_fd_sc_hd__o21ai_4
X_63602_ _58446_/A _63600_/X _63575_/C _63661_/D _63602_/Y sky130_fd_sc_hd__nand4_4
X_60814_ _60707_/X _60812_/Y _60748_/X _60732_/Y _60813_/Y _84560_/D
+ sky130_fd_sc_hd__a41oi_4
X_48536_ _48612_/A _48536_/X sky130_fd_sc_hd__buf_2
X_67370_ _67320_/A _87218_/Q _67370_/X sky130_fd_sc_hd__and2_4
X_79356_ _79346_/A _79346_/B _79341_/Y _79344_/Y _79356_/X sky130_fd_sc_hd__o22a_4
X_45748_ _45668_/A _45748_/X sky130_fd_sc_hd__buf_2
X_64582_ _64582_/A _64582_/B _64582_/Y sky130_fd_sc_hd__nand2_4
X_76568_ _76566_/Y _76567_/Y _81373_/Q _76568_/Y sky130_fd_sc_hd__a21oi_4
X_61794_ _61376_/X _61794_/B _59810_/A _61776_/D _61794_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_10_814_0_CLK clkbuf_9_407_0_CLK/X _82557_/CLK sky130_fd_sc_hd__clkbuf_1
X_66321_ _66267_/X _74232_/B _66321_/X sky130_fd_sc_hd__and2_4
X_78307_ _78309_/A _78309_/C _78307_/X sky130_fd_sc_hd__and2_4
X_63533_ _63496_/A _58528_/A _63520_/C _63546_/D _63533_/X sky130_fd_sc_hd__and4_4
X_75519_ _75519_/A _75516_/Y _75519_/C _75519_/X sky130_fd_sc_hd__or3_4
X_48467_ _83583_/Q _74414_/B sky130_fd_sc_hd__inv_2
X_60745_ _60671_/C _60737_/Y _60743_/X _60694_/Y _60744_/Y _84577_/D
+ sky130_fd_sc_hd__a41oi_4
X_79287_ _84796_/Q _84116_/Q _79287_/X sky130_fd_sc_hd__xor2_4
X_45679_ _45674_/X _45677_/Y _45678_/X _45679_/X sky130_fd_sc_hd__a21o_4
X_76499_ _76497_/X _76498_/Y _76499_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_9_305_0_CLK clkbuf_8_152_0_CLK/X clkbuf_9_305_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_69040_ _68929_/X _69029_/Y _68824_/X _69039_/Y _69040_/X sky130_fd_sc_hd__a211o_4
X_47418_ _47418_/A _47415_/X _47377_/X _53036_/D _47418_/X sky130_fd_sc_hd__and4_4
X_66252_ _66237_/X _74129_/B _66252_/X sky130_fd_sc_hd__and2_4
X_78238_ _78234_/Y _78237_/X _78239_/B sky130_fd_sc_hd__nand2_4
X_63464_ _61427_/B _63426_/X _63462_/X _63463_/X _63464_/X sky130_fd_sc_hd__a211o_4
X_60676_ _60632_/A _60677_/A sky130_fd_sc_hd__inv_2
X_48398_ _48393_/Y _48383_/X _48397_/X _86526_/D sky130_fd_sc_hd__a21oi_4
X_65203_ _65227_/A _86250_/Q _65203_/X sky130_fd_sc_hd__and2_4
X_62415_ _62269_/A _62415_/X sky130_fd_sc_hd__buf_2
X_47349_ _47380_/A _47349_/B _47370_/C _52997_/D _47349_/X sky130_fd_sc_hd__and4_4
X_66183_ _66054_/X _66183_/B _66183_/X sky130_fd_sc_hd__and2_4
X_78169_ _78177_/A _78177_/B _78172_/A sky130_fd_sc_hd__xor2_4
X_63395_ _63458_/A _63410_/C sky130_fd_sc_hd__buf_2
Xclkbuf_10_829_0_CLK clkbuf_9_414_0_CLK/X _86582_/CLK sky130_fd_sc_hd__clkbuf_1
X_80200_ _80184_/Y _80187_/Y _80199_/X _80200_/X sky130_fd_sc_hd__a21o_4
X_65134_ _65131_/X _65133_/X _64959_/X _65134_/X sky130_fd_sc_hd__a21o_4
X_50360_ _50360_/A _50331_/B _50338_/X _50360_/X sky130_fd_sc_hd__and3_4
X_62346_ _62288_/X _62285_/X _64320_/B _62609_/D _62346_/X sky130_fd_sc_hd__and4_4
X_81180_ _81197_/CLK _75036_/X _81180_/Q sky130_fd_sc_hd__dfxtp_4
X_49019_ _49019_/A _49009_/B _49019_/Y sky130_fd_sc_hd__nor2_4
X_80131_ _80125_/A _80124_/X _80130_/Y _80131_/Y sky130_fd_sc_hd__a21boi_4
X_65065_ _64809_/A _65065_/X sky130_fd_sc_hd__buf_2
X_69942_ _81957_/D _69894_/X _69941_/X _83885_/D sky130_fd_sc_hd__a21bo_4
X_50291_ _50279_/X _53516_/B _50291_/Y sky130_fd_sc_hd__nand2_4
X_62277_ _62276_/X _62623_/C sky130_fd_sc_hd__buf_2
X_52030_ _52028_/Y _52022_/X _52029_/Y _52030_/Y sky130_fd_sc_hd__a21boi_4
X_64016_ _83248_/Q _64046_/B _64046_/C _64016_/D _64017_/D sky130_fd_sc_hd__nand4_4
X_80062_ _80058_/X _80074_/B _80073_/A sky130_fd_sc_hd__xor2_4
X_61228_ _61234_/A _61250_/B _84503_/Q _61228_/Y sky130_fd_sc_hd__nor3_4
X_69873_ _87292_/Q _69873_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_5_5_0_CLK clkbuf_4_2_1_CLK/X clkbuf_5_5_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_68824_ _68649_/A _68824_/X sky130_fd_sc_hd__buf_2
X_61159_ _61082_/X _64456_/C sky130_fd_sc_hd__buf_2
X_84870_ _84892_/CLK _84870_/D _84870_/Q sky130_fd_sc_hd__dfxtp_4
X_83821_ _83819_/CLK _70257_/X _74771_/A sky130_fd_sc_hd__dfxtp_4
X_68755_ _68779_/A _68755_/B _68755_/X sky130_fd_sc_hd__and2_4
X_53981_ _85529_/Q _53955_/X _53980_/Y _53981_/Y sky130_fd_sc_hd__o21ai_4
X_65967_ _65962_/X _65967_/B _65966_/X _65967_/Y sky130_fd_sc_hd__nand3_4
X_55720_ _55276_/A _55794_/A sky130_fd_sc_hd__buf_2
X_86540_ _86570_/CLK _86540_/D _66214_/B sky130_fd_sc_hd__dfxtp_4
X_67706_ _67466_/X _67706_/X sky130_fd_sc_hd__buf_2
X_52932_ _85728_/Q _52929_/X _52931_/Y _52932_/Y sky130_fd_sc_hd__o21ai_4
X_64918_ _44175_/A _65669_/A sky130_fd_sc_hd__buf_2
X_83752_ _84280_/CLK _70546_/X _83752_/Q sky130_fd_sc_hd__dfxtp_4
X_68686_ _68735_/A _68686_/B _68686_/X sky130_fd_sc_hd__and2_4
X_80964_ _81990_/CLK _75597_/X _75393_/B sky130_fd_sc_hd__dfxtp_4
X_65898_ _65894_/X _65868_/B _65897_/X _65898_/Y sky130_fd_sc_hd__nand3_4
X_82703_ _82610_/CLK _82703_/D _82659_/D sky130_fd_sc_hd__dfxtp_4
X_55651_ _74539_/A _56171_/A sky130_fd_sc_hd__buf_2
X_67637_ _68129_/A _67637_/X sky130_fd_sc_hd__buf_2
X_86471_ _86471_/CLK _48850_/Y _86471_/Q sky130_fd_sc_hd__dfxtp_4
X_52863_ _52850_/A _52863_/B _52863_/Y sky130_fd_sc_hd__nand2_4
X_64849_ _64846_/X _85560_/Q _64642_/X _64848_/X _64849_/X sky130_fd_sc_hd__a211o_4
X_83683_ _85786_/CLK _70850_/Y _83683_/Q sky130_fd_sc_hd__dfxtp_4
X_80895_ _83967_/CLK _80895_/D _80895_/Q sky130_fd_sc_hd__dfxtp_4
X_88210_ _87888_/CLK _41466_/X _88210_/Q sky130_fd_sc_hd__dfxtp_4
X_54602_ _54521_/A _54607_/B sky130_fd_sc_hd__buf_2
X_85422_ _85648_/CLK _85422_/D _85422_/Q sky130_fd_sc_hd__dfxtp_4
X_51814_ _51814_/A _51815_/B sky130_fd_sc_hd__buf_2
X_82634_ _87926_/CLK _83986_/Q _78870_/A sky130_fd_sc_hd__dfxtp_4
X_58370_ _58370_/A _58369_/X _58370_/Y sky130_fd_sc_hd__nand2_4
X_55582_ _55572_/X _45455_/Y _55582_/Y sky130_fd_sc_hd__nor2_4
X_67568_ _67806_/A _67568_/X sky130_fd_sc_hd__buf_2
X_52794_ _52803_/A _52794_/B _52794_/Y sky130_fd_sc_hd__nand2_4
X_57321_ _45909_/A _45738_/Y _57320_/X _57321_/X sky130_fd_sc_hd__o21a_4
X_69307_ _69303_/X _69306_/X _69116_/X _69307_/X sky130_fd_sc_hd__a21o_4
X_88141_ _87373_/CLK _41810_/X _88141_/Q sky130_fd_sc_hd__dfxtp_4
X_54533_ _54518_/A _53360_/B _54533_/Y sky130_fd_sc_hd__nand2_4
X_66519_ _66517_/Y _66518_/Y _60529_/A _66519_/X sky130_fd_sc_hd__a21o_4
X_85353_ _86600_/CLK _54923_/Y _85353_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_12 sky130_fd_sc_hd__decap_3
X_51745_ _85953_/Q _51387_/X _51744_/Y _51745_/Y sky130_fd_sc_hd__o21ai_4
X_82565_ _82942_/CLK _82565_/D _82565_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_23 sky130_fd_sc_hd__decap_3
X_67499_ _67144_/A _67572_/A sky130_fd_sc_hd__buf_2
XPHY_34 sky130_fd_sc_hd__decap_3
XPHY_45 sky130_fd_sc_hd__decap_3
X_84304_ _84358_/CLK _63664_/Y _80357_/B sky130_fd_sc_hd__dfxtp_4
X_57252_ _57243_/X _56607_/X _45504_/A _57245_/X _85050_/D sky130_fd_sc_hd__a2bb2o_4
X_81516_ _81755_/CLK _81560_/Q _81516_/Q sky130_fd_sc_hd__dfxtp_4
X_69238_ _69235_/X _69237_/X _69138_/X _69238_/X sky130_fd_sc_hd__a21o_4
XPHY_56 sky130_fd_sc_hd__decap_3
X_88072_ _87821_/CLK _42012_/Y _88072_/Q sky130_fd_sc_hd__dfxtp_4
X_54464_ _54478_/A _54464_/B _54464_/Y sky130_fd_sc_hd__nand2_4
X_85284_ _83013_/CLK _85284_/D _56165_/C sky130_fd_sc_hd__dfxtp_4
XPHY_67 sky130_fd_sc_hd__decap_3
X_51676_ _50222_/X _51697_/A sky130_fd_sc_hd__buf_2
X_82496_ _82671_/CLK _82496_/D _82496_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_78 sky130_fd_sc_hd__decap_3
XPHY_89 sky130_fd_sc_hd__decap_3
X_56203_ _56200_/X _56192_/B _56203_/C _56203_/Y sky130_fd_sc_hd__nand3_4
X_87023_ _88301_/CLK _87023_/D _87023_/Q sky130_fd_sc_hd__dfxtp_4
X_53415_ _53413_/Y _53408_/X _53414_/X _53415_/Y sky130_fd_sc_hd__a21oi_4
X_84235_ _82786_/CLK _84235_/D _64542_/A sky130_fd_sc_hd__dfxtp_4
X_50627_ _50596_/A _50627_/X sky130_fd_sc_hd__buf_2
X_81447_ _81575_/CLK _81447_/D _81447_/Q sky130_fd_sc_hd__dfxtp_4
X_57183_ _56816_/Y _57182_/X _57183_/X sky130_fd_sc_hd__xor2_4
X_69169_ _69073_/A _88305_/Q _69169_/X sky130_fd_sc_hd__and2_4
X_54395_ _54395_/A _54395_/B _54395_/C _54395_/D _54395_/X sky130_fd_sc_hd__and4_4
X_71200_ _48561_/B _71190_/X _71199_/Y _71200_/Y sky130_fd_sc_hd__o21ai_4
X_56134_ _56134_/A _56134_/X sky130_fd_sc_hd__buf_2
X_41360_ _41261_/X _41703_/B _41359_/X _41360_/Y sky130_fd_sc_hd__o21ai_4
X_53346_ _85650_/Q _53324_/X _53345_/Y _53346_/Y sky130_fd_sc_hd__o21ai_4
X_72180_ _57711_/X _72180_/X sky130_fd_sc_hd__buf_2
X_84166_ _84166_/CLK _84166_/D _84166_/Q sky130_fd_sc_hd__dfxtp_4
X_50558_ _50541_/A _48878_/B _50558_/Y sky130_fd_sc_hd__nand2_4
X_81378_ _83914_/CLK _83914_/Q _76792_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_82_0_CLK clkbuf_7_83_0_CLK/A clkbuf_7_82_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_71131_ _71129_/A _71064_/B _70914_/D _71131_/Y sky130_fd_sc_hd__nand3_4
X_83117_ _86213_/CLK _83117_/D _70130_/A sky130_fd_sc_hd__dfxtp_4
X_80329_ _80324_/Y _80328_/Y _80329_/Y sky130_fd_sc_hd__nand2_4
X_56065_ _45765_/A _56086_/B sky130_fd_sc_hd__buf_2
X_41291_ _41186_/A _41292_/B sky130_fd_sc_hd__buf_2
X_53277_ _85663_/Q _53268_/X _53276_/Y _53277_/Y sky130_fd_sc_hd__o21ai_4
X_84097_ _80928_/CLK _84097_/D _80921_/D sky130_fd_sc_hd__dfxtp_4
X_50489_ _50465_/X _48811_/B _50489_/Y sky130_fd_sc_hd__nand2_4
X_43030_ _43030_/A _43189_/A sky130_fd_sc_hd__buf_2
X_55016_ _85334_/Q _54994_/X _55015_/Y _55016_/Y sky130_fd_sc_hd__o21ai_4
X_52228_ _48845_/A _52248_/B _52223_/C _52228_/X sky130_fd_sc_hd__and3_4
X_71062_ _71058_/A _70952_/B _71066_/C _71062_/Y sky130_fd_sc_hd__nand3_4
X_87925_ _87926_/CLK _87925_/D _87925_/Q sky130_fd_sc_hd__dfxtp_4
X_83048_ _83049_/CLK _74521_/Y _83048_/Q sky130_fd_sc_hd__dfxtp_4
X_70013_ _69679_/X _69681_/X _70001_/X _70013_/Y sky130_fd_sc_hd__a21oi_4
X_59824_ _59588_/Y _59824_/B _59823_/X _59825_/B sky130_fd_sc_hd__nand3_4
X_52159_ _85877_/Q _52152_/X _52158_/Y _52159_/Y sky130_fd_sc_hd__o21ai_4
X_75870_ _75862_/Y _75875_/B _75870_/Y sky130_fd_sc_hd__nand2_4
X_87856_ _87068_/CLK _42464_/Y _87856_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_97_0_CLK clkbuf_7_96_0_CLK/A clkbuf_7_97_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_74821_ _74829_/A _46111_/B _74822_/A sky130_fd_sc_hd__nand2_4
X_86807_ _86807_/CLK _46026_/X _86807_/Q sky130_fd_sc_hd__dfxtp_4
X_59755_ _59755_/A _59756_/A sky130_fd_sc_hd__buf_2
X_44981_ _56206_/C _44911_/X _44980_/X _44981_/Y sky130_fd_sc_hd__o21ai_4
X_56967_ _56966_/X _56639_/X _45597_/A _56989_/A _85108_/D sky130_fd_sc_hd__a2bb2o_4
X_87787_ _87544_/CLK _42650_/Y _87787_/Q sky130_fd_sc_hd__dfxtp_4
X_84999_ _83335_/CLK _84999_/D _84999_/Q sky130_fd_sc_hd__dfxtp_4
X_46720_ _46720_/A _46733_/A sky130_fd_sc_hd__buf_2
X_58706_ _58928_/A _58706_/X sky130_fd_sc_hd__buf_2
X_77540_ _77540_/A _77540_/B _77540_/C _77561_/C sky130_fd_sc_hd__or3_4
X_43932_ _43932_/A _43932_/Y sky130_fd_sc_hd__inv_2
X_55918_ _55918_/A _55928_/C sky130_fd_sc_hd__buf_2
X_74752_ _74752_/A _74745_/Y _74748_/Y _74751_/Y _74758_/B sky130_fd_sc_hd__and4_4
X_86738_ _86246_/CLK _46429_/Y _86738_/Q sky130_fd_sc_hd__dfxtp_4
X_71964_ _71964_/A _71964_/X sky130_fd_sc_hd__buf_2
X_59686_ _59637_/A _59806_/A _59699_/A _59686_/Y sky130_fd_sc_hd__o21ai_4
X_56898_ _56898_/A _59498_/A _56898_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_7_20_0_CLK clkbuf_7_21_0_CLK/A clkbuf_8_41_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_73703_ _73700_/X _73702_/X _73679_/X _73719_/B sky130_fd_sc_hd__a21o_4
X_70915_ _51016_/B _70909_/X _70914_/Y _70915_/Y sky130_fd_sc_hd__o21ai_4
X_46651_ _46651_/A _51770_/B _46651_/Y sky130_fd_sc_hd__nand2_4
X_58637_ _58631_/X _58633_/Y _58634_/Y _58007_/X _58636_/X _58637_/X
+ sky130_fd_sc_hd__o32a_4
X_77471_ _77471_/A _77471_/B _77472_/A sky130_fd_sc_hd__nand2_4
X_55849_ _85202_/Q _55462_/X _55512_/X _55848_/X _55849_/X sky130_fd_sc_hd__a211o_4
X_43863_ _43776_/A _43863_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_160_0_CLK clkbuf_7_80_0_CLK/X clkbuf_8_160_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_74683_ _74675_/X _56820_/A _74682_/Y _74684_/A sky130_fd_sc_hd__o21ai_4
X_86669_ _86351_/CLK _86669_/D _59245_/A sky130_fd_sc_hd__dfxtp_4
X_71895_ _71894_/Y _71898_/D sky130_fd_sc_hd__buf_2
X_79210_ _79208_/Y _79209_/Y _82821_/D sky130_fd_sc_hd__xor2_4
X_45602_ _45678_/A _45602_/X sky130_fd_sc_hd__buf_2
X_76422_ _76387_/B _76420_/X _76421_/Y _76422_/Y sky130_fd_sc_hd__a21oi_4
X_42814_ _41433_/X _42802_/X _67972_/B _42803_/X _42814_/X sky130_fd_sc_hd__a2bb2o_4
X_49370_ _49374_/A _49369_/X _49380_/C _51756_/D _49370_/X sky130_fd_sc_hd__and4_4
X_73634_ _88368_/Q _73633_/X _73028_/X _73634_/Y sky130_fd_sc_hd__o21ai_4
X_46582_ _51384_/B _52565_/B sky130_fd_sc_hd__buf_2
X_70846_ _70873_/A _70846_/B _70849_/C _70860_/D _70846_/Y sky130_fd_sc_hd__nand4_4
X_58568_ _58679_/A _58568_/X sky130_fd_sc_hd__buf_2
X_43794_ _43790_/X _43781_/X _41045_/X _69397_/B _43791_/X _43795_/A
+ sky130_fd_sc_hd__o32ai_4
X_48321_ _48934_/A _49247_/A sky130_fd_sc_hd__buf_2
X_79141_ _79141_/A _79141_/B _79141_/X sky130_fd_sc_hd__xor2_4
X_45533_ _85080_/Q _45533_/Y sky130_fd_sc_hd__inv_2
X_57519_ _84987_/Q _57493_/X _57518_/Y _57519_/Y sky130_fd_sc_hd__o21ai_4
X_76353_ _76348_/X _76353_/B _76349_/Y _76353_/Y sky130_fd_sc_hd__nand3_4
X_88339_ _88337_/CLK _88339_/D _88339_/Q sky130_fd_sc_hd__dfxtp_4
X_42745_ _42745_/A _42745_/X sky130_fd_sc_hd__buf_2
X_73565_ _73562_/X _73564_/X _73383_/X _73570_/A sky130_fd_sc_hd__a21o_4
X_70777_ _70382_/A _70778_/A sky130_fd_sc_hd__buf_2
X_58499_ _58448_/X _83410_/Q _58498_/Y _84834_/D sky130_fd_sc_hd__o21a_4
Xclkbuf_7_35_0_CLK clkbuf_7_35_0_CLK/A clkbuf_8_71_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_75304_ _75304_/A _75304_/Y sky130_fd_sc_hd__inv_2
X_60530_ _60526_/A _60526_/B _79145_/A _60530_/Y sky130_fd_sc_hd__nor3_4
X_48252_ _48229_/A _50300_/B _48252_/Y sky130_fd_sc_hd__nand2_4
X_72516_ _72516_/A _72516_/B _72516_/C _72517_/B sky130_fd_sc_hd__nand3_4
Xclkbuf_8_175_0_CLK clkbuf_7_87_0_CLK/X clkbuf_9_351_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_79072_ _82655_/Q _79074_/A sky130_fd_sc_hd__inv_2
X_45464_ _44895_/X _45464_/X sky130_fd_sc_hd__buf_2
X_76284_ _76293_/A _76283_/Y _76284_/X sky130_fd_sc_hd__or2_4
Xclkbuf_10_170_0_CLK clkbuf_9_85_0_CLK/X _81587_/CLK sky130_fd_sc_hd__clkbuf_1
X_42676_ _41050_/X _42652_/X _69409_/B _42653_/X _87775_/D sky130_fd_sc_hd__a2bb2o_4
X_73496_ _73378_/X _86180_/Q _73446_/X _73495_/X _73496_/X sky130_fd_sc_hd__a211o_4
X_47203_ _47197_/Y _47177_/X _47202_/X _47203_/Y sky130_fd_sc_hd__a21oi_4
X_78023_ _78020_/Y _78022_/Y _82144_/D sky130_fd_sc_hd__nor2_4
X_44415_ _44404_/X _44405_/X _41536_/X _87120_/Q _44406_/X _44415_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75235_ _75242_/A _75234_/Y _81037_/D sky130_fd_sc_hd__xnor2_4
X_41627_ _41626_/X _41581_/X _67324_/B _41582_/X _41627_/X sky130_fd_sc_hd__a2bb2o_4
X_48183_ _47861_/B _50234_/B sky130_fd_sc_hd__buf_2
X_60461_ _79154_/A _60246_/X _60571_/B _60445_/Y _84614_/D sky130_fd_sc_hd__a2bb2oi_4
X_72447_ _72447_/A _72476_/B _72447_/Y sky130_fd_sc_hd__nor2_4
X_45395_ _80671_/Q _45395_/X sky130_fd_sc_hd__buf_2
X_62200_ _62572_/A _62212_/A sky130_fd_sc_hd__buf_2
X_47134_ _47126_/Y _47128_/X _47133_/X _47134_/Y sky130_fd_sc_hd__a21oi_4
X_44346_ _40509_/X _44346_/X sky130_fd_sc_hd__buf_2
X_63180_ _63144_/X _84826_/Q _63146_/C _63135_/D _63180_/X sky130_fd_sc_hd__and4_4
Xclkbuf_9_291_0_CLK clkbuf_9_291_0_CLK/A clkbuf_9_291_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_75166_ _75164_/Y _75135_/Y _75165_/X _75167_/B sky130_fd_sc_hd__o21ai_4
X_41558_ _81166_/Q _41584_/B _41558_/X sky130_fd_sc_hd__or2_4
X_60392_ _60392_/A _60392_/B _60392_/C _60512_/A _60501_/A sky130_fd_sc_hd__and4_4
X_72378_ _72378_/A _72401_/B _72378_/Y sky130_fd_sc_hd__nor2_4
X_62131_ _59794_/X _62088_/B _62131_/C _62131_/D _62131_/Y sky130_fd_sc_hd__nand4_4
X_74117_ _74117_/A _74116_/Y _74117_/Y sky130_fd_sc_hd__nor2_4
X_40509_ _40353_/Y _40509_/X sky130_fd_sc_hd__buf_2
X_47065_ _82386_/Q _54526_/D sky130_fd_sc_hd__inv_2
X_71329_ _71335_/A _71335_/B _71302_/X _71329_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_185_0_CLK clkbuf_9_92_0_CLK/X _80720_/CLK sky130_fd_sc_hd__clkbuf_1
X_44277_ _57331_/B _44277_/X sky130_fd_sc_hd__buf_2
X_79974_ _60136_/C _84271_/Q _79974_/Y sky130_fd_sc_hd__xnor2_4
X_75097_ _80676_/Q _80932_/D _75099_/A sky130_fd_sc_hd__nand2_4
X_41489_ _41336_/X _41489_/X sky130_fd_sc_hd__buf_2
X_46016_ _46016_/A _46016_/Y sky130_fd_sc_hd__inv_2
X_43228_ _43227_/Y _87528_/D sky130_fd_sc_hd__inv_2
X_62062_ _61747_/X _62065_/B sky130_fd_sc_hd__buf_2
X_74048_ _74046_/X _74048_/B _74048_/C _74048_/Y sky130_fd_sc_hd__nand3_4
X_78925_ _78918_/Y _78919_/A _78924_/Y _78925_/Y sky130_fd_sc_hd__a21oi_4
X_61013_ _61202_/A _60908_/X _61013_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_8_113_0_CLK clkbuf_7_56_0_CLK/X clkbuf_8_113_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_66870_ _88391_/Q _66868_/X _66801_/X _66869_/X _66870_/X sky130_fd_sc_hd__a211o_4
X_43159_ _43146_/X _43149_/X _40861_/X _73228_/A _43154_/X _43160_/A
+ sky130_fd_sc_hd__o32ai_4
X_78856_ _78856_/A _78856_/Y sky130_fd_sc_hd__inv_2
X_65821_ _65704_/A _86471_/Q _65821_/X sky130_fd_sc_hd__and2_4
X_77807_ _82267_/Q _81979_/Q _77807_/Y sky130_fd_sc_hd__xnor2_4
X_47967_ _83772_/Q _47967_/Y sky130_fd_sc_hd__inv_2
X_78787_ _78782_/Y _78786_/X _78795_/A sky130_fd_sc_hd__nand2_4
X_75999_ _76005_/B _76005_/C _75999_/Y sky130_fd_sc_hd__nand2_4
X_49706_ _49787_/A _49706_/X sky130_fd_sc_hd__buf_2
X_68540_ _66180_/A _68540_/X sky130_fd_sc_hd__buf_2
X_46918_ _46915_/X _46896_/B _46926_/C _52746_/D _46918_/X sky130_fd_sc_hd__and4_4
X_65752_ _65749_/X _65751_/X _65614_/X _65752_/X sky130_fd_sc_hd__a21o_4
X_77738_ _82051_/Q _77738_/Y sky130_fd_sc_hd__inv_2
X_62964_ _58201_/X _62924_/C _62827_/X _62818_/X _62963_/X _62964_/Y
+ sky130_fd_sc_hd__a41oi_4
X_47898_ _47841_/A _47912_/A sky130_fd_sc_hd__buf_2
X_64703_ _65607_/A _64712_/B sky130_fd_sc_hd__buf_2
Xclkbuf_8_128_0_CLK clkbuf_7_64_0_CLK/X clkbuf_8_128_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_61915_ _61915_/A _61915_/B _58520_/A _61915_/D _61915_/X sky130_fd_sc_hd__and4_4
X_49637_ _49635_/Y _49623_/X _49636_/X _49637_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_123_0_CLK clkbuf_9_61_0_CLK/X _84671_/CLK sky130_fd_sc_hd__clkbuf_1
X_68471_ _68466_/X _68469_/X _68470_/X _68471_/X sky130_fd_sc_hd__a21o_4
X_46849_ _46843_/Y _46844_/X _46848_/X _86697_/D sky130_fd_sc_hd__a21oi_4
X_65683_ _65634_/A _65802_/B _65683_/C _65683_/Y sky130_fd_sc_hd__nor3_4
X_77669_ _77596_/B _77663_/X _77668_/Y _77695_/B sky130_fd_sc_hd__a21oi_4
X_62895_ _62892_/X _62893_/X _62894_/Y _62895_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_753_0_CLK clkbuf_9_376_0_CLK/X _87273_/CLK sky130_fd_sc_hd__clkbuf_1
X_79408_ _79392_/X _79396_/B _79408_/X sky130_fd_sc_hd__or2_4
X_67422_ _87164_/Q _67348_/X _67398_/X _67421_/X _67422_/X sky130_fd_sc_hd__a211o_4
X_64634_ _64561_/X _64623_/Y _64633_/Y _64634_/Y sky130_fd_sc_hd__o21ai_4
X_49568_ _86363_/Q _49551_/X _49567_/Y _49568_/Y sky130_fd_sc_hd__o21ai_4
X_61846_ _61844_/X _61846_/B _61846_/C _61846_/D _61846_/Y sky130_fd_sc_hd__nand4_4
X_80680_ _80681_/CLK _80680_/D _80680_/Q sky130_fd_sc_hd__dfxtp_4
X_48519_ _48461_/A _48565_/B sky130_fd_sc_hd__buf_2
Xclkbuf_9_244_0_CLK clkbuf_9_245_0_CLK/A clkbuf_9_244_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_67353_ _81505_/D _67331_/X _67352_/X _67353_/X sky130_fd_sc_hd__a21bo_4
X_79339_ _79333_/Y _79339_/B _82832_/D sky130_fd_sc_hd__xor2_4
X_64565_ _64565_/A _64766_/A sky130_fd_sc_hd__buf_2
X_61777_ _61777_/A _61795_/C sky130_fd_sc_hd__buf_2
X_49499_ _86376_/Q _49496_/X _49498_/Y _49499_/Y sky130_fd_sc_hd__o21ai_4
X_66304_ _65838_/X _66276_/B _65840_/X _66304_/Y sky130_fd_sc_hd__nand3_4
X_51530_ _85993_/Q _51511_/X _51529_/Y _51530_/Y sky130_fd_sc_hd__o21ai_4
X_63516_ _63516_/A _63516_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_138_0_CLK clkbuf_9_69_0_CLK/X _81361_/CLK sky130_fd_sc_hd__clkbuf_1
X_82350_ _82369_/CLK _82350_/D _82350_/Q sky130_fd_sc_hd__dfxtp_4
X_60728_ _84580_/Q _60719_/X _60671_/Y _60727_/Y _60728_/X sky130_fd_sc_hd__o22a_4
X_67284_ _67046_/A _67284_/X sky130_fd_sc_hd__buf_2
X_64496_ _64515_/A _59427_/A _64515_/C _64496_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_768_0_CLK clkbuf_9_384_0_CLK/X _82531_/CLK sky130_fd_sc_hd__clkbuf_1
X_81301_ _81689_/CLK _76989_/X _81301_/Q sky130_fd_sc_hd__dfxtp_4
X_69023_ _68934_/X _69023_/B _69023_/Y sky130_fd_sc_hd__nor2_4
X_66235_ _66125_/X _86218_/Q _66180_/X _66234_/X _66235_/X sky130_fd_sc_hd__a211o_4
X_51461_ _86006_/Q _51458_/X _51460_/Y _51461_/Y sky130_fd_sc_hd__o21ai_4
X_63447_ _63445_/Y _63391_/X _63446_/Y _84323_/D sky130_fd_sc_hd__a21oi_4
X_82281_ _82288_/CLK _82281_/D _82281_/Q sky130_fd_sc_hd__dfxtp_4
X_60659_ _60659_/A _60660_/A sky130_fd_sc_hd__buf_2
X_53200_ _53219_/A _53200_/B _53200_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_259_0_CLK clkbuf_9_259_0_CLK/A clkbuf_9_259_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_84020_ _84020_/CLK _68176_/X _82060_/D sky130_fd_sc_hd__dfxtp_4
X_50412_ _53636_/A _50430_/B _50435_/C _50412_/X sky130_fd_sc_hd__and3_4
X_81232_ _81233_/CLK _81040_/Q _81232_/Q sky130_fd_sc_hd__dfxtp_4
X_54180_ _85489_/Q _54167_/X _54179_/Y _54180_/Y sky130_fd_sc_hd__o21ai_4
X_66166_ _57694_/X _66166_/B _66166_/X sky130_fd_sc_hd__and2_4
X_51392_ _47857_/X _46591_/A _51392_/X sky130_fd_sc_hd__and2_4
X_63378_ _63632_/A _63443_/A sky130_fd_sc_hd__buf_2
X_53131_ _53121_/X _53131_/B _53131_/Y sky130_fd_sc_hd__nand2_4
X_65117_ _65117_/A _65118_/A sky130_fd_sc_hd__buf_2
X_50343_ _50356_/A _48297_/X _50343_/Y sky130_fd_sc_hd__nand2_4
X_62329_ _62326_/Y _62327_/X _62328_/Y _84418_/D sky130_fd_sc_hd__a21oi_4
X_81163_ _81125_/CLK _74911_/B _41572_/A sky130_fd_sc_hd__dfxtp_4
X_66097_ _66054_/X _66097_/B _66097_/X sky130_fd_sc_hd__and2_4
X_80114_ _80114_/A _80114_/Y sky130_fd_sc_hd__inv_2
X_53062_ _53062_/A _53074_/C sky130_fd_sc_hd__buf_2
X_65048_ _65043_/Y _64939_/X _65047_/Y _65048_/X sky130_fd_sc_hd__a21o_4
X_69925_ _69655_/A _69925_/X sky130_fd_sc_hd__buf_2
X_50274_ _50227_/A _50274_/X sky130_fd_sc_hd__buf_2
X_85971_ _84787_/CLK _51652_/Y _85971_/Q sky130_fd_sc_hd__dfxtp_4
X_81094_ _81094_/CLK _81094_/D _81094_/Q sky130_fd_sc_hd__dfxtp_4
X_52013_ _52152_/A _52013_/X sky130_fd_sc_hd__buf_2
X_87710_ _87644_/CLK _42804_/X _87710_/Q sky130_fd_sc_hd__dfxtp_4
X_84922_ _84922_/CLK _84922_/D _84922_/Q sky130_fd_sc_hd__dfxtp_4
X_80045_ _80052_/B _80045_/B _80045_/X sky130_fd_sc_hd__xor2_4
X_57870_ _57971_/A _57870_/B _57870_/Y sky130_fd_sc_hd__nor2_4
X_69856_ _69429_/X _69432_/X _69816_/X _69856_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_706_0_CLK clkbuf_9_353_0_CLK/X _86796_/CLK sky130_fd_sc_hd__clkbuf_1
X_56821_ _56816_/A _56821_/X sky130_fd_sc_hd__buf_2
X_68807_ _68803_/X _68805_/X _68806_/X _68807_/X sky130_fd_sc_hd__a21o_4
X_87641_ _87195_/CLK _87641_/D _87641_/Q sky130_fd_sc_hd__dfxtp_4
X_84853_ _84732_/CLK _58419_/X _84853_/Q sky130_fd_sc_hd__dfxtp_4
X_69787_ _69746_/X _69785_/Y _69733_/X _69786_/Y _69787_/X sky130_fd_sc_hd__a211o_4
X_66999_ _66902_/X _86820_/Q _66999_/X sky130_fd_sc_hd__and2_4
X_59540_ _60593_/A _59540_/Y sky130_fd_sc_hd__inv_2
X_83804_ _83813_/CLK _83804_/D _83804_/Q sky130_fd_sc_hd__dfxtp_4
X_56752_ _56752_/A _56798_/B _56765_/A sky130_fd_sc_hd__nand2_4
X_68738_ _68734_/X _68736_/X _68737_/X _68738_/Y sky130_fd_sc_hd__a21oi_4
X_87572_ _88326_/CLK _87572_/D _74266_/A sky130_fd_sc_hd__dfxtp_4
X_53964_ _53964_/A _53964_/B _53888_/C _53964_/X sky130_fd_sc_hd__and3_4
X_84784_ _84823_/CLK _84784_/D _84784_/Q sky130_fd_sc_hd__dfxtp_4
X_81996_ _81996_/CLK _81996_/D _77066_/A sky130_fd_sc_hd__dfxtp_4
X_55703_ _85254_/Q _55174_/X _44044_/X _55702_/X _55703_/X sky130_fd_sc_hd__a211o_4
X_86523_ _86523_/CLK _48432_/Y _65525_/B sky130_fd_sc_hd__dfxtp_4
X_52915_ _85731_/Q _52902_/X _52914_/Y _52915_/Y sky130_fd_sc_hd__o21ai_4
X_83735_ _83736_/CLK _83735_/D _83735_/Q sky130_fd_sc_hd__dfxtp_4
X_59471_ _59471_/A _59478_/B _59471_/Y sky130_fd_sc_hd__nand2_4
X_56683_ _56682_/X _56739_/A sky130_fd_sc_hd__buf_2
X_80947_ _80740_/CLK _80991_/Q _74969_/A sky130_fd_sc_hd__dfxtp_4
X_68669_ _68669_/A _68669_/B _68669_/Y sky130_fd_sc_hd__nor2_4
X_53895_ _53661_/A _53921_/A sky130_fd_sc_hd__buf_2
X_70700_ _70700_/A _70700_/B _71115_/C _70701_/A sky130_fd_sc_hd__nor3_4
X_58422_ _58406_/X _83364_/Q _58421_/Y _84852_/D sky130_fd_sc_hd__o21a_4
X_55634_ _55634_/A _56564_/C sky130_fd_sc_hd__buf_2
X_86454_ _85555_/CLK _49000_/Y _86454_/Q sky130_fd_sc_hd__dfxtp_4
X_40860_ _40857_/X _41034_/A _40859_/X _40861_/A sky130_fd_sc_hd__o21a_4
X_52846_ _52853_/A _52831_/B _52853_/C _52846_/D _52846_/X sky130_fd_sc_hd__and4_4
X_71680_ _71680_/A _71671_/X _71680_/C _71680_/Y sky130_fd_sc_hd__nand3_4
X_83666_ _83666_/CLK _83666_/D _83666_/Q sky130_fd_sc_hd__dfxtp_4
X_80878_ _80754_/CLK _75686_/B _80878_/Q sky130_fd_sc_hd__dfxtp_4
X_85405_ _85499_/CLK _85405_/D _85405_/Q sky130_fd_sc_hd__dfxtp_4
X_70631_ _70630_/X _70631_/X sky130_fd_sc_hd__buf_2
X_58353_ _58341_/X _58350_/Y _58352_/Y _58353_/Y sky130_fd_sc_hd__a21oi_4
X_82617_ _82617_/CLK _79019_/B _82617_/Q sky130_fd_sc_hd__dfxtp_4
X_55565_ _55843_/A _85146_/Q _55565_/X sky130_fd_sc_hd__and2_4
X_86385_ _83673_/CLK _86385_/D _86385_/Q sky130_fd_sc_hd__dfxtp_4
X_40791_ _40628_/X _82876_/Q _40790_/X _40792_/A sky130_fd_sc_hd__o21ai_4
X_52777_ _52773_/A _52777_/B _52777_/Y sky130_fd_sc_hd__nand2_4
X_83597_ _86149_/CLK _83597_/D _83597_/Q sky130_fd_sc_hd__dfxtp_4
X_57304_ _57303_/Y _57010_/Y _57304_/Y sky130_fd_sc_hd__nand2_4
X_88124_ _87675_/CLK _41849_/X _67136_/B sky130_fd_sc_hd__dfxtp_4
X_42530_ _74184_/A _69023_/B sky130_fd_sc_hd__inv_2
X_54516_ _54509_/A _54503_/B _54509_/C _47047_/A _54516_/X sky130_fd_sc_hd__and4_4
X_85336_ _85334_/CLK _55010_/Y _85336_/Q sky130_fd_sc_hd__dfxtp_4
X_73350_ _44577_/Y _73006_/X _73349_/Y _73365_/C sky130_fd_sc_hd__a21o_4
X_51728_ _51737_/A _51728_/B _51728_/Y sky130_fd_sc_hd__nand2_4
X_70562_ _71570_/A _71863_/A sky130_fd_sc_hd__buf_2
X_58284_ _84888_/Q _63655_/B sky130_fd_sc_hd__buf_2
X_82548_ _82541_/CLK _83868_/Q _79123_/B sky130_fd_sc_hd__dfxtp_4
X_55496_ _45585_/A _55454_/X _55457_/X _55495_/Y _55496_/X sky130_fd_sc_hd__a211o_4
X_72301_ _72347_/A _72301_/B _72301_/Y sky130_fd_sc_hd__nor2_4
X_57235_ _45886_/X _45882_/A _45898_/X _56183_/X _44038_/X _57235_/Y
+ sky130_fd_sc_hd__a41oi_4
X_88055_ _88056_/CLK _42056_/Y _73462_/A sky130_fd_sc_hd__dfxtp_4
X_42461_ _87856_/Q _68440_/B sky130_fd_sc_hd__inv_2
X_54447_ _85440_/Q _54431_/X _54446_/Y _54447_/Y sky130_fd_sc_hd__o21ai_4
X_73281_ _87051_/Q _73129_/X _73280_/X _73281_/Y sky130_fd_sc_hd__o21ai_4
X_85267_ _85168_/CLK _56230_/Y _85267_/Q sky130_fd_sc_hd__dfxtp_4
X_51659_ _51654_/Y _51639_/X _51658_/X _51659_/Y sky130_fd_sc_hd__a21oi_4
X_70493_ _70907_/B _70696_/B sky130_fd_sc_hd__buf_2
X_82479_ _82855_/CLK _82479_/D _78108_/B sky130_fd_sc_hd__dfxtp_4
X_44200_ _44167_/Y _44186_/X _44220_/B _44200_/Y sky130_fd_sc_hd__a21oi_4
X_75020_ _75008_/X _80768_/Q _75020_/C _75020_/Y sky130_fd_sc_hd__nand3_4
X_41412_ _41411_/X _41412_/X sky130_fd_sc_hd__buf_2
X_87006_ _86984_/CLK _44672_/Y _87006_/Q sky130_fd_sc_hd__dfxtp_4
X_72232_ _72220_/A _72232_/B _72232_/Y sky130_fd_sc_hd__nor2_4
X_84218_ _84220_/CLK _84218_/D _84218_/Q sky130_fd_sc_hd__dfxtp_4
X_45180_ _55826_/B _45120_/X _45153_/X _45180_/X sky130_fd_sc_hd__o21a_4
X_57166_ _57162_/Y _57165_/X _57192_/A _57166_/X sky130_fd_sc_hd__a21o_4
X_42392_ _42392_/A _87886_/D sky130_fd_sc_hd__inv_2
X_54378_ _54378_/A _52686_/B _54378_/Y sky130_fd_sc_hd__nand2_4
X_85198_ _85198_/CLK _85198_/D _85198_/Q sky130_fd_sc_hd__dfxtp_4
X_44131_ _44131_/A _72784_/A sky130_fd_sc_hd__inv_2
X_56117_ _56117_/A _56117_/B _56117_/C _56118_/A sky130_fd_sc_hd__and3_4
X_41343_ _41343_/A _41343_/Y sky130_fd_sc_hd__inv_2
X_53329_ _53302_/A _53330_/C sky130_fd_sc_hd__buf_2
X_72163_ _59237_/X _72160_/Y _72162_/Y _59301_/X _59241_/X _72163_/X
+ sky130_fd_sc_hd__o32a_4
X_84149_ _82746_/CLK _84149_/D _80419_/B sky130_fd_sc_hd__dfxtp_4
X_57097_ _57096_/Y _57097_/X sky130_fd_sc_hd__buf_2
X_71114_ _50169_/B _71095_/A _71113_/Y _71114_/Y sky130_fd_sc_hd__o21ai_4
X_44062_ _44061_/X _55470_/A sky130_fd_sc_hd__buf_2
X_56048_ _55928_/A _74310_/C _55928_/C _56045_/Y _56047_/Y _56048_/Y
+ sky130_fd_sc_hd__a32oi_4
X_41274_ _41013_/A _41275_/B sky130_fd_sc_hd__buf_2
X_72094_ _72075_/A _53919_/B _72094_/Y sky130_fd_sc_hd__nand2_4
X_76971_ _76971_/A _84395_/Q _76971_/X sky130_fd_sc_hd__xor2_4
X_43013_ _43175_/C _43013_/X sky130_fd_sc_hd__buf_2
X_78710_ _78710_/A _82685_/D _78713_/B sky130_fd_sc_hd__nor2_4
X_71045_ _70828_/A _70959_/B _70959_/C _71115_/B _71046_/A sky130_fd_sc_hd__and4_4
X_75922_ _84520_/Q _84392_/Q _75922_/X sky130_fd_sc_hd__xor2_4
X_87908_ _87898_/CLK _87908_/D _87908_/Q sky130_fd_sc_hd__dfxtp_4
X_48870_ _48702_/A _48859_/B _48854_/C _48870_/X sky130_fd_sc_hd__and3_4
X_79690_ _84215_/Q _83263_/Q _79692_/A sky130_fd_sc_hd__xor2_4
X_47821_ _81218_/Q _47822_/A sky130_fd_sc_hd__inv_2
X_59807_ _59807_/A _59840_/A sky130_fd_sc_hd__buf_2
X_78641_ _78640_/A _78640_/C _78621_/A _78641_/Y sky130_fd_sc_hd__a21oi_4
X_75853_ _75831_/A _75841_/A _75853_/X sky130_fd_sc_hd__and2_4
X_87839_ _87850_/CLK _42512_/Y _87839_/Q sky130_fd_sc_hd__dfxtp_4
X_57999_ _57983_/X _85389_/Q _57998_/X _57999_/Y sky130_fd_sc_hd__o21ai_4
X_74804_ _74804_/A _74804_/B _74804_/C _74804_/D _74804_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_1010_0_CLK clkbuf_9_505_0_CLK/X _83310_/CLK sky130_fd_sc_hd__clkbuf_1
X_47752_ _47752_/A _53227_/B sky130_fd_sc_hd__buf_2
X_59738_ _59727_/X _59728_/Y _59686_/Y _59733_/Y _59737_/Y _59738_/Y
+ sky130_fd_sc_hd__a41oi_4
X_78572_ _78572_/A _78572_/Y sky130_fd_sc_hd__inv_2
X_44964_ _44887_/X _44964_/X sky130_fd_sc_hd__buf_2
X_75784_ _75784_/A _75783_/Y _80889_/D sky130_fd_sc_hd__xnor2_4
X_72996_ _74403_/B _72996_/B _72996_/X sky130_fd_sc_hd__xor2_4
X_46703_ _58677_/A _46672_/X _46702_/Y _46703_/Y sky130_fd_sc_hd__o21ai_4
X_77523_ _77512_/B _77523_/Y sky130_fd_sc_hd__inv_2
X_43915_ _43914_/Y _43915_/Y sky130_fd_sc_hd__inv_2
X_74735_ _74734_/Y _74735_/X sky130_fd_sc_hd__buf_2
X_47683_ _47682_/Y _53185_/D sky130_fd_sc_hd__buf_2
X_71947_ _70383_/X _70766_/C _71349_/D _71945_/D _71947_/Y sky130_fd_sc_hd__nand4_4
X_59669_ _45923_/X _64738_/A sky130_fd_sc_hd__buf_2
X_44895_ _45193_/A _44895_/X sky130_fd_sc_hd__buf_2
X_49422_ _49418_/A _51807_/B _49422_/Y sky130_fd_sc_hd__nand2_4
X_61700_ _61690_/A _61690_/B _84458_/Q _61700_/Y sky130_fd_sc_hd__nor3_4
X_46634_ _54277_/B _50893_/B sky130_fd_sc_hd__buf_2
X_77454_ _77447_/A _77444_/Y _77446_/A _77454_/X sky130_fd_sc_hd__o21a_4
X_43846_ _43810_/A _43846_/X sky130_fd_sc_hd__buf_2
X_62680_ _62679_/X _62694_/B sky130_fd_sc_hd__buf_2
X_74666_ _74675_/A _74679_/A sky130_fd_sc_hd__buf_2
X_71878_ _71319_/B _71883_/D sky130_fd_sc_hd__buf_2
X_76405_ _76387_/B _76387_/A _76404_/X _76405_/Y sky130_fd_sc_hd__a21boi_4
X_61631_ _58348_/A _61598_/X _61677_/C _61563_/D _61632_/A sky130_fd_sc_hd__nand4_4
X_49353_ _65381_/B _49334_/X _49352_/Y _49353_/Y sky130_fd_sc_hd__o21ai_4
X_73617_ _72829_/X _84991_/Q _73614_/X _73616_/X _73617_/X sky130_fd_sc_hd__a211o_4
X_46565_ _46547_/A _51378_/B _46565_/Y sky130_fd_sc_hd__nand2_4
X_70829_ _70832_/A _70830_/B sky130_fd_sc_hd__inv_2
X_77385_ _77385_/A _77386_/B sky130_fd_sc_hd__buf_2
X_43777_ _43774_/X _43760_/X _40994_/X _69288_/B _43776_/X _43777_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74597_ _45216_/A _74582_/X _74596_/X _83021_/D sky130_fd_sc_hd__o21ai_4
X_40989_ _40989_/A _40989_/X sky130_fd_sc_hd__buf_2
X_48304_ _48301_/Y _48302_/X _48303_/X _86539_/D sky130_fd_sc_hd__a21oi_4
X_79124_ _79123_/Y _79124_/Y sky130_fd_sc_hd__inv_2
X_45516_ _45596_/A _45516_/X sky130_fd_sc_hd__buf_2
X_64350_ _79764_/B _64314_/X _64349_/X _64350_/X sky130_fd_sc_hd__a21o_4
X_76336_ _76336_/A _76336_/B _76337_/A sky130_fd_sc_hd__and2_4
X_42728_ _42721_/X _42723_/X _41193_/X _68755_/B _42700_/X _42728_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49284_ _49280_/Y _49281_/X _49283_/X _49284_/Y sky130_fd_sc_hd__a21oi_4
X_61562_ _61380_/A _61563_/D sky130_fd_sc_hd__buf_2
X_73548_ _83146_/Q _73437_/X _73547_/Y _73548_/X sky130_fd_sc_hd__a21o_4
X_46496_ _46493_/X _82924_/Q _46495_/Y _54047_/A sky130_fd_sc_hd__o21ai_4
X_63301_ _84871_/Q _63281_/B _63301_/C _63281_/D _63301_/X sky130_fd_sc_hd__or4_4
X_48235_ _48232_/Y _48233_/X _48234_/X _48235_/Y sky130_fd_sc_hd__a21oi_4
X_60513_ _60513_/A _60513_/B _79148_/A _60513_/X sky130_fd_sc_hd__or3_4
X_79055_ _79055_/A _79055_/B _79057_/C sky130_fd_sc_hd__nor2_4
X_45447_ _45441_/X _45445_/X _45446_/X _45447_/X sky130_fd_sc_hd__a21o_4
X_64281_ _84260_/Q _64255_/X _64280_/X _84260_/D sky130_fd_sc_hd__a21o_4
X_76267_ _76267_/A _76267_/B _76273_/A sky130_fd_sc_hd__nand2_4
X_42659_ _42647_/X _42648_/X _41004_/X _87783_/Q _42658_/X _42659_/Y
+ sky130_fd_sc_hd__o32ai_4
X_61493_ _59411_/A _61484_/B _61484_/C _61452_/D _61494_/A sky130_fd_sc_hd__nand4_4
X_73479_ _48672_/A _73478_/Y _73479_/X sky130_fd_sc_hd__xor2_4
X_66020_ _66366_/A _66020_/X sky130_fd_sc_hd__buf_2
X_78006_ _78003_/A _78006_/B _78006_/Y sky130_fd_sc_hd__nand2_4
X_63232_ _63228_/Y _63230_/X _63231_/X _63232_/Y sky130_fd_sc_hd__a21oi_4
X_75218_ _75207_/Y _75190_/Y _75205_/A _75218_/Y sky130_fd_sc_hd__a21oi_4
X_48166_ _73568_/B _40568_/X _48165_/X _48166_/Y sky130_fd_sc_hd__o21ai_4
X_60444_ _60515_/C _60476_/D _60399_/B _72296_/A _72176_/A _60444_/Y
+ sky130_fd_sc_hd__o32ai_4
X_45378_ _45651_/A _45378_/X sky130_fd_sc_hd__buf_2
X_76198_ _76199_/B _76198_/Y sky130_fd_sc_hd__inv_2
X_47117_ _47109_/A _52863_/B _47117_/Y sky130_fd_sc_hd__nand2_4
X_44329_ _44587_/A _44381_/A sky130_fd_sc_hd__buf_2
X_63163_ _79372_/A _63130_/X _63162_/Y _63163_/X sky130_fd_sc_hd__a21o_4
X_75149_ _75147_/Y _75148_/Y _81031_/D sky130_fd_sc_hd__xor2_4
X_48097_ _47867_/X _82920_/Q _48096_/Y _57619_/A sky130_fd_sc_hd__o21ai_4
X_60375_ _60359_/X _60252_/X _60229_/Y _60363_/Y _60374_/Y _84618_/D
+ sky130_fd_sc_hd__a41oi_4
X_62114_ _61712_/X _62175_/B sky130_fd_sc_hd__buf_2
X_47048_ _47029_/A _47039_/B _47048_/C _52827_/D _47048_/X sky130_fd_sc_hd__and4_4
X_67971_ _81479_/D _67925_/X _67970_/X _84047_/D sky130_fd_sc_hd__a21bo_4
X_63094_ _79436_/A _63072_/X _63093_/Y _84354_/D sky130_fd_sc_hd__a21o_4
X_79957_ _79957_/A _79957_/B _79957_/C _79957_/Y sky130_fd_sc_hd__nand3_4
X_69710_ _69687_/A _69710_/B _69710_/Y sky130_fd_sc_hd__nor2_4
X_66922_ _66918_/X _66921_/X _66871_/X _66922_/Y sky130_fd_sc_hd__a21oi_4
X_62045_ _59699_/A _62046_/D sky130_fd_sc_hd__buf_2
X_78908_ _78908_/A _78907_/Y _78909_/B sky130_fd_sc_hd__xnor2_4
X_79888_ _79883_/X _79888_/B _79889_/A sky130_fd_sc_hd__xnor2_4
X_69641_ _69208_/X _69210_/X _69575_/X _69641_/Y sky130_fd_sc_hd__a21oi_4
X_66853_ _87943_/Q _66759_/X _66807_/X _66852_/X _66853_/X sky130_fd_sc_hd__a211o_4
X_78839_ _82838_/Q _78839_/B _78839_/X sky130_fd_sc_hd__xor2_4
X_48999_ _49022_/A _72014_/B _48999_/X sky130_fd_sc_hd__and2_4
X_65804_ _65804_/A _85864_/Q _65804_/X sky130_fd_sc_hd__and2_4
X_81850_ _82221_/CLK _81882_/Q _77582_/A sky130_fd_sc_hd__dfxtp_4
X_69572_ _69586_/A _88339_/Q _69572_/X sky130_fd_sc_hd__and2_4
X_66784_ _68614_/A _66785_/A sky130_fd_sc_hd__buf_2
X_63996_ _63993_/X _63994_/X _63995_/Y _84282_/D sky130_fd_sc_hd__a21oi_4
X_80801_ _81065_/CLK _75872_/B _80801_/Q sky130_fd_sc_hd__dfxtp_4
X_68523_ _68444_/A _88365_/Q _68523_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_692_0_CLK clkbuf_9_346_0_CLK/X _88398_/CLK sky130_fd_sc_hd__clkbuf_1
X_65735_ _65735_/A _86477_/Q _65735_/X sky130_fd_sc_hd__and2_4
X_50961_ _50938_/X _50961_/B _50961_/Y sky130_fd_sc_hd__nand2_4
X_62947_ _61637_/X _62926_/B _62681_/X _60228_/A _62947_/Y sky130_fd_sc_hd__nand4_4
X_81781_ _81703_/CLK _76113_/X _81781_/Q sky130_fd_sc_hd__dfxtp_4
X_52700_ _52706_/A _52700_/B _52700_/Y sky130_fd_sc_hd__nand2_4
X_83520_ _83520_/CLK _83520_/D _83520_/Q sky130_fd_sc_hd__dfxtp_4
X_80732_ _83749_/CLK _75918_/X _80732_/Q sky130_fd_sc_hd__dfxtp_4
X_68454_ _68449_/X _68453_/X _68429_/X _68454_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_9_183_0_CLK clkbuf_8_91_0_CLK/X clkbuf_9_183_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_53680_ _53747_/A _53680_/X sky130_fd_sc_hd__buf_2
X_65666_ _65664_/Y _65602_/X _65665_/X _84186_/D sky130_fd_sc_hd__a21o_4
X_50892_ _50889_/Y _50839_/X _50891_/X _50892_/Y sky130_fd_sc_hd__a21oi_4
X_62878_ _62869_/A _62935_/B _62027_/X _62878_/Y sky130_fd_sc_hd__nand3_4
X_67405_ _67046_/A _67405_/X sky130_fd_sc_hd__buf_2
X_52631_ _52657_/A _52637_/A sky130_fd_sc_hd__buf_2
X_64617_ _64769_/A _64617_/B _64617_/X sky130_fd_sc_hd__and2_4
X_83451_ _83451_/CLK _83451_/D _58336_/B sky130_fd_sc_hd__dfxtp_4
X_61829_ _61399_/X _61794_/B _61809_/C _61776_/D _61829_/Y sky130_fd_sc_hd__nand4_4
X_80663_ _80657_/CLK _74817_/Y _46188_/A sky130_fd_sc_hd__dfxtp_4
X_68385_ _68385_/A _68385_/X sky130_fd_sc_hd__buf_2
X_65597_ _65474_/X _73070_/B _65597_/X sky130_fd_sc_hd__and2_4
X_82402_ _82786_/CLK _82434_/Q _78312_/A sky130_fd_sc_hd__dfxtp_4
X_55350_ _82993_/Q _44061_/X _55312_/X _55349_/X _55352_/C sky130_fd_sc_hd__a211o_4
X_67336_ _87475_/Q _67239_/X _67240_/X _67335_/X _67336_/X sky130_fd_sc_hd__a211o_4
X_86170_ _83306_/CLK _86170_/D _86170_/Q sky130_fd_sc_hd__dfxtp_4
X_52562_ _52560_/Y _52541_/X _52561_/Y _85797_/D sky130_fd_sc_hd__a21boi_4
X_64548_ _58990_/Y _64226_/X _64547_/Y _64548_/Y sky130_fd_sc_hd__o21ai_4
X_83382_ _83415_/CLK _71771_/X _83382_/Q sky130_fd_sc_hd__dfxtp_4
X_80594_ _80593_/Y _80571_/X _80594_/X sky130_fd_sc_hd__and2_4
XPHY_407 sky130_fd_sc_hd__decap_3
XPHY_418 sky130_fd_sc_hd__decap_3
X_54301_ _85467_/Q _54294_/X _54300_/Y _54301_/Y sky130_fd_sc_hd__o21ai_4
XPHY_429 sky130_fd_sc_hd__decap_3
X_85121_ _85074_/CLK _56942_/X _85121_/Q sky130_fd_sc_hd__dfxtp_4
X_51513_ _51622_/A _51514_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_198_0_CLK clkbuf_8_99_0_CLK/X clkbuf_9_198_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_82333_ _82284_/CLK _77199_/B _82333_/Q sky130_fd_sc_hd__dfxtp_4
X_67267_ _88374_/Q _67193_/X _67194_/X _67266_/X _67267_/X sky130_fd_sc_hd__a211o_4
X_55281_ _55281_/A _55282_/B sky130_fd_sc_hd__inv_2
X_52493_ _52491_/Y _52486_/X _52492_/Y _52493_/Y sky130_fd_sc_hd__a21boi_4
X_64479_ _58277_/A _61085_/X _64478_/Y _64479_/Y sky130_fd_sc_hd__o21ai_4
X_57020_ _56797_/A _56796_/Y _44213_/X _57020_/Y sky130_fd_sc_hd__a21oi_4
X_69006_ _69003_/X _69005_/X _60014_/X _69006_/Y sky130_fd_sc_hd__a21oi_4
X_54232_ _54208_/X _54237_/B _54237_/C _53063_/D _54232_/X sky130_fd_sc_hd__and4_4
X_66218_ _66123_/A _66151_/B _84148_/Q _66218_/X sky130_fd_sc_hd__and3_4
X_85052_ _85050_/CLK _85052_/D _85052_/Q sky130_fd_sc_hd__dfxtp_4
X_51444_ _51441_/Y _51420_/X _51443_/X _86009_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_630_0_CLK clkbuf_9_315_0_CLK/X _82133_/CLK sky130_fd_sc_hd__clkbuf_1
X_82264_ _83515_/CLK _82264_/D _82264_/Q sky130_fd_sc_hd__dfxtp_4
X_67198_ _67131_/A _87609_/Q _67198_/X sky130_fd_sc_hd__and2_4
X_84003_ _84003_/CLK _68242_/X _84003_/Q sky130_fd_sc_hd__dfxtp_4
X_81215_ _82284_/CLK _74874_/X _81215_/Q sky130_fd_sc_hd__dfxtp_4
X_54163_ _85492_/Q _54140_/X _54162_/Y _54163_/Y sky130_fd_sc_hd__o21ai_4
X_66149_ _66068_/X _65676_/Y _66148_/Y _66149_/Y sky130_fd_sc_hd__o21ai_4
X_51375_ _86022_/Q _51362_/X _51374_/Y _51375_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_121_0_CLK clkbuf_8_60_0_CLK/X clkbuf_9_121_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_82195_ _85491_/CLK _82195_/D _82387_/D sky130_fd_sc_hd__dfxtp_4
X_53114_ _53110_/Y _53111_/X _53113_/X _85695_/D sky130_fd_sc_hd__a21oi_4
X_50326_ _50356_/A _50326_/B _50326_/Y sky130_fd_sc_hd__nand2_4
X_81146_ _82327_/CLK _81146_/D _40624_/A sky130_fd_sc_hd__dfxtp_4
X_54094_ _85505_/Q _53431_/X _54093_/Y _54094_/Y sky130_fd_sc_hd__o21ai_4
X_58971_ _58559_/X _83441_/Q _58970_/Y _58971_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_10_645_0_CLK clkbuf_9_322_0_CLK/X _83987_/CLK sky130_fd_sc_hd__clkbuf_1
X_53045_ _53042_/Y _53028_/X _53044_/X _53045_/Y sky130_fd_sc_hd__a21oi_4
X_57922_ _84939_/Q _57922_/Y sky130_fd_sc_hd__inv_2
X_69908_ _69908_/A _42611_/Y _69908_/Y sky130_fd_sc_hd__nor2_4
X_50257_ _50918_/A _50257_/X sky130_fd_sc_hd__buf_2
X_85954_ _85471_/CLK _51743_/Y _85954_/Q sky130_fd_sc_hd__dfxtp_4
X_81077_ _81121_/CLK _81109_/Q _75348_/A sky130_fd_sc_hd__dfxtp_4
X_80028_ _80026_/X _80027_/X _80043_/B sky130_fd_sc_hd__xnor2_4
X_84905_ _84905_/CLK _84905_/D _84905_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_136_0_CLK clkbuf_8_68_0_CLK/X clkbuf_9_136_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_57853_ _57852_/X _85721_/Q _57814_/X _57853_/X sky130_fd_sc_hd__o21a_4
X_69839_ _73275_/A _69837_/X _69779_/X _69838_/Y _69839_/X sky130_fd_sc_hd__a211o_4
X_50188_ _50187_/X _50188_/B _50188_/Y sky130_fd_sc_hd__nand2_4
X_85885_ _83572_/CLK _52120_/Y _85885_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_63_0_CLK clkbuf_9_63_0_CLK/A clkbuf_9_63_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_56804_ _56758_/X _56756_/X _56788_/X _57163_/C _45835_/A _56804_/Y
+ sky130_fd_sc_hd__a41oi_4
X_87624_ _87883_/CLK _87624_/D _87624_/Q sky130_fd_sc_hd__dfxtp_4
X_72850_ _83174_/Q _72794_/X _72849_/Y _83174_/D sky130_fd_sc_hd__a21o_4
X_84836_ _84308_/CLK _84836_/D _84836_/Q sky130_fd_sc_hd__dfxtp_4
X_57784_ _69182_/A _58749_/A sky130_fd_sc_hd__buf_2
X_54996_ _55011_/A _47589_/Y _54996_/Y sky130_fd_sc_hd__nand2_4
X_71801_ _70370_/A _71716_/B _71439_/C _71716_/D _71801_/X sky130_fd_sc_hd__and4_4
X_59523_ _59519_/C _59741_/C sky130_fd_sc_hd__buf_2
X_56735_ _57149_/D _56735_/X sky130_fd_sc_hd__buf_2
X_41961_ _41960_/X _41951_/X _40724_/X _74121_/A _41953_/X _41961_/Y
+ sky130_fd_sc_hd__o32ai_4
X_87555_ _88060_/CLK _43156_/Y _87555_/Q sky130_fd_sc_hd__dfxtp_4
X_53947_ _85536_/Q _53921_/X _53946_/Y _53947_/Y sky130_fd_sc_hd__o21ai_4
X_72781_ _73535_/A _65441_/B _72781_/X sky130_fd_sc_hd__and2_4
X_84767_ _86361_/CLK _59128_/Y _84767_/Q sky130_fd_sc_hd__dfxtp_4
X_81979_ _82234_/CLK _83907_/Q _81979_/Q sky130_fd_sc_hd__dfxtp_4
X_43700_ _43606_/A _43700_/X sky130_fd_sc_hd__buf_2
X_74520_ _70374_/X _74518_/B _70880_/C _74518_/D _74520_/Y sky130_fd_sc_hd__nand4_4
X_86506_ _86506_/CLK _86506_/D _86506_/Q sky130_fd_sc_hd__dfxtp_4
X_40912_ _40829_/A _40912_/B _40912_/X sky130_fd_sc_hd__or2_4
X_71732_ _58240_/Y _71711_/Y _71731_/Y _71732_/Y sky130_fd_sc_hd__o21ai_4
X_59454_ _59454_/A _59444_/X _59454_/Y sky130_fd_sc_hd__nand2_4
X_83718_ _83721_/CLK _70718_/Y _83718_/Q sky130_fd_sc_hd__dfxtp_4
X_44680_ _41936_/A _44680_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_78_0_CLK clkbuf_9_79_0_CLK/A clkbuf_9_78_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_56666_ _56972_/A _56650_/Y _56665_/Y _56666_/Y sky130_fd_sc_hd__a21oi_4
X_87486_ _87487_/CLK _87486_/D _87486_/Q sky130_fd_sc_hd__dfxtp_4
X_41892_ _41887_/X _41888_/X _40590_/X _41889_/Y _41891_/X _41892_/Y
+ sky130_fd_sc_hd__o32ai_4
X_53878_ _85550_/Q _53846_/X _53877_/Y _53878_/Y sky130_fd_sc_hd__o21ai_4
X_84698_ _84713_/CLK _59800_/Y _80464_/A sky130_fd_sc_hd__dfxtp_4
X_58405_ _58981_/A _58423_/A sky130_fd_sc_hd__buf_2
X_43631_ _40660_/X _43609_/X _68695_/B _43611_/X _43632_/A sky130_fd_sc_hd__a2bb2o_4
X_55617_ _55617_/A _55617_/X sky130_fd_sc_hd__buf_2
X_74451_ _74442_/X _48559_/Y _74451_/Y sky130_fd_sc_hd__nand2_4
X_86437_ _86436_/CLK _86437_/D _86437_/Q sky130_fd_sc_hd__dfxtp_4
X_40843_ _82866_/Q _40842_/X _40843_/X sky130_fd_sc_hd__or2_4
X_52829_ _52843_/A _52829_/B _52829_/Y sky130_fd_sc_hd__nand2_4
X_59385_ _84746_/Q _59339_/X _59378_/X _59384_/X _59385_/Y sky130_fd_sc_hd__a2bb2oi_4
X_71663_ _58522_/Y _71649_/A _71662_/Y _83420_/D sky130_fd_sc_hd__o21ai_4
X_83649_ _82774_/CLK _70963_/Y _83649_/Q sky130_fd_sc_hd__dfxtp_4
X_56597_ _55562_/X _55568_/X _56597_/X sky130_fd_sc_hd__and2_4
X_73402_ _73257_/X _86184_/Q _73351_/X _73401_/X _73402_/X sky130_fd_sc_hd__a211o_4
X_46350_ _46350_/A _46380_/B _46350_/X sky130_fd_sc_hd__or2_4
X_70614_ _52991_/B _70584_/X _70613_/Y _83741_/D sky130_fd_sc_hd__o21ai_4
X_58336_ _58151_/A _58336_/B _58336_/Y sky130_fd_sc_hd__nor2_4
X_77170_ _77170_/A _77170_/B _77171_/A sky130_fd_sc_hd__nand2_4
X_43562_ _40485_/X _43560_/X _87360_/Q _43561_/X _87360_/D sky130_fd_sc_hd__a2bb2o_4
X_55548_ _83000_/Q _55511_/X _55532_/X _55547_/X _56616_/B sky130_fd_sc_hd__a211o_4
X_74382_ _74380_/Y _74370_/X _74381_/X _74382_/Y sky130_fd_sc_hd__a21oi_4
X_86368_ _83721_/CLK _49545_/Y _86368_/Q sky130_fd_sc_hd__dfxtp_4
X_40774_ _82879_/Q _40765_/B _40774_/X sky130_fd_sc_hd__or2_4
X_71594_ _71189_/B _71598_/C sky130_fd_sc_hd__buf_2
X_45301_ _56444_/C _45252_/X _45300_/X _45301_/Y sky130_fd_sc_hd__o21ai_4
X_76121_ _81533_/Q _76121_/B _76121_/X sky130_fd_sc_hd__xor2_4
X_88107_ _87595_/CLK _88107_/D _41914_/A sky130_fd_sc_hd__dfxtp_4
X_42513_ _42495_/X _42496_/X _40707_/X _87838_/Q _42506_/X _42514_/A
+ sky130_fd_sc_hd__o32ai_4
X_73333_ _73330_/X _73332_/X _72877_/X _73333_/X sky130_fd_sc_hd__a21o_4
X_85319_ _85351_/CLK _55097_/Y _85319_/Q sky130_fd_sc_hd__dfxtp_4
X_46281_ _83654_/Q _52440_/B sky130_fd_sc_hd__inv_2
X_70545_ _71586_/A _70692_/B _70538_/X _70550_/D _70545_/Y sky130_fd_sc_hd__nor4_4
X_58267_ _84892_/Q _58268_/A sky130_fd_sc_hd__inv_2
X_43493_ _41727_/X _43484_/X _87393_/Q _43485_/X _43493_/X sky130_fd_sc_hd__a2bb2o_4
X_55479_ _55474_/X _55478_/X _55646_/A sky130_fd_sc_hd__and2_4
X_86299_ _86301_/CLK _49921_/Y _72192_/B sky130_fd_sc_hd__dfxtp_4
X_48020_ _47981_/X _48020_/B _48020_/X sky130_fd_sc_hd__and2_4
X_45232_ _45232_/A _45199_/B _45232_/Y sky130_fd_sc_hd__nand2_4
X_57218_ _57216_/Y _57217_/Y _57112_/X _57218_/Y sky130_fd_sc_hd__a21oi_4
X_76052_ _76048_/Y _76051_/X _76052_/Y sky130_fd_sc_hd__nand2_4
X_42444_ _40548_/X _42434_/X _87860_/Q _42435_/X _42444_/X sky130_fd_sc_hd__a2bb2o_4
X_88038_ _88044_/CLK _42093_/Y _88038_/Q sky130_fd_sc_hd__dfxtp_4
X_73264_ _73516_/A _73407_/A sky130_fd_sc_hd__buf_2
X_70476_ _70382_/A _70476_/X sky130_fd_sc_hd__buf_2
X_58198_ _58198_/A _58184_/B _58198_/Y sky130_fd_sc_hd__nor2_4
X_75003_ _81143_/D _75003_/B _75003_/Y sky130_fd_sc_hd__nand2_4
X_72215_ _72180_/X _85337_/Q _59365_/X _72215_/X sky130_fd_sc_hd__o21a_4
X_45163_ _85264_/Q _45147_/X _45162_/X _45163_/Y sky130_fd_sc_hd__o21ai_4
X_57149_ _56700_/Y _57149_/B _57149_/C _57149_/D _57149_/X sky130_fd_sc_hd__and4_4
X_42375_ _42304_/X _42375_/X sky130_fd_sc_hd__buf_2
X_73195_ _73195_/A _73196_/B sky130_fd_sc_hd__buf_2
Xclkbuf_9_16_0_CLK clkbuf_8_8_0_CLK/X clkbuf_9_16_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_44114_ _44113_/X _44115_/A sky130_fd_sc_hd__buf_2
X_79811_ _79795_/X _79798_/Y _79810_/X _79811_/X sky130_fd_sc_hd__a21o_4
X_41326_ _41326_/A _41325_/X _41326_/X sky130_fd_sc_hd__or2_4
X_72146_ _59037_/A _72146_/X sky130_fd_sc_hd__buf_2
X_60160_ _59574_/A _60160_/B _60222_/C sky130_fd_sc_hd__and2_4
X_49971_ _49981_/A _53183_/B _49971_/Y sky130_fd_sc_hd__nand2_4
X_45094_ _45094_/A _45095_/A sky130_fd_sc_hd__inv_2
X_48922_ _48901_/A _48922_/B _48922_/Y sky130_fd_sc_hd__nand2_4
X_44045_ _44044_/X _44045_/X sky130_fd_sc_hd__buf_2
X_79742_ _79742_/A _79742_/B _79742_/X sky130_fd_sc_hd__xor2_4
X_41257_ _81703_/Q _41280_/B _41257_/X sky130_fd_sc_hd__or2_4
X_60091_ _60091_/A _60091_/B _60091_/C _60091_/Y sky130_fd_sc_hd__nand3_4
X_72077_ _72053_/A _72077_/B _72077_/Y sky130_fd_sc_hd__nand2_4
X_76954_ _76957_/A _76957_/C _76956_/A sky130_fd_sc_hd__nand2_4
Xclkbuf_9_4_0_CLK clkbuf_9_5_0_CLK/A clkbuf_9_4_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_71028_ _53153_/B _71013_/X _71027_/Y _83631_/D sky130_fd_sc_hd__o21ai_4
X_75905_ _84503_/Q _62873_/C _75905_/X sky130_fd_sc_hd__xor2_4
X_48853_ _48853_/A _48854_/C sky130_fd_sc_hd__buf_2
X_79673_ _79669_/X _79672_/Y _79673_/X sky130_fd_sc_hd__xor2_4
X_41188_ _41184_/X _81139_/Q _41187_/X _41189_/A sky130_fd_sc_hd__o21ai_4
X_76885_ _81500_/Q _76884_/X _76885_/X sky130_fd_sc_hd__xor2_4
X_47804_ _47804_/A _49364_/B _50886_/C _53253_/D _47804_/X sky130_fd_sc_hd__and4_4
X_78624_ _78586_/Y _78588_/X _78623_/A _78640_/A sky130_fd_sc_hd__a21o_4
X_63850_ _63848_/X _63849_/X _84291_/Q _63850_/Y sky130_fd_sc_hd__nor3_4
X_75836_ _75836_/A _75836_/B _80894_/D sky130_fd_sc_hd__xor2_4
X_48784_ _86483_/Q _48781_/X _48783_/Y _48784_/Y sky130_fd_sc_hd__o21ai_4
X_45996_ _45994_/X _45987_/X _40458_/X _66938_/B _45995_/X _45996_/Y
+ sky130_fd_sc_hd__o32ai_4
X_62801_ _62681_/X _62801_/X sky130_fd_sc_hd__buf_2
X_47735_ _47715_/X _53213_/B _47735_/Y sky130_fd_sc_hd__nand2_4
X_78555_ _78555_/A _78552_/A _78555_/Y sky130_fd_sc_hd__nand2_4
X_44947_ _56386_/C _44945_/X _44946_/X _44947_/Y sky130_fd_sc_hd__o21ai_4
X_63781_ _61356_/X _63781_/B _63781_/C _63761_/X _63781_/Y sky130_fd_sc_hd__nand4_4
X_75767_ _81015_/Q _80887_/D _75767_/X sky130_fd_sc_hd__xor2_4
X_60993_ _60992_/X _60993_/B _60934_/X _60993_/Y sky130_fd_sc_hd__nor3_4
X_72979_ _44272_/X _72979_/X sky130_fd_sc_hd__buf_2
X_65520_ _65334_/X _86203_/Q _65517_/X _65519_/X _65520_/X sky130_fd_sc_hd__a211o_4
X_77506_ _77507_/A _82101_/D _77509_/B sky130_fd_sc_hd__nor2_4
X_62732_ _62726_/Y _62713_/X _62727_/Y _62729_/Y _62731_/X _62732_/X
+ sky130_fd_sc_hd__a41o_4
X_74718_ _74739_/B _74720_/C sky130_fd_sc_hd__buf_2
X_47666_ _47619_/A _47666_/X sky130_fd_sc_hd__buf_2
X_78486_ _78472_/X _82798_/Q _78485_/Y _78486_/Y sky130_fd_sc_hd__a21oi_4
X_44878_ _45387_/A _44932_/A sky130_fd_sc_hd__buf_2
X_75698_ _75684_/Y _75697_/X _75703_/A sky130_fd_sc_hd__nand2_4
X_49405_ _49405_/A _49405_/X sky130_fd_sc_hd__buf_2
X_46617_ _46617_/A _46659_/C sky130_fd_sc_hd__buf_2
X_65451_ _65401_/A _65451_/B _65451_/X sky130_fd_sc_hd__and2_4
X_77437_ _77412_/X _77413_/Y _77416_/A _77437_/Y sky130_fd_sc_hd__a21boi_4
X_43829_ _43810_/X _43824_/X _41139_/X _87246_/Q _43811_/X _43830_/A
+ sky130_fd_sc_hd__o32ai_4
X_62663_ _60202_/A _62664_/D sky130_fd_sc_hd__buf_2
X_74649_ _74638_/X _56619_/A _83000_/Q _74645_/X _74649_/X sky130_fd_sc_hd__a2bb2o_4
X_47597_ _47597_/A _47598_/A sky130_fd_sc_hd__inv_2
X_64402_ _64285_/A _64402_/X sky130_fd_sc_hd__buf_2
X_49336_ _49352_/A _50858_/B _49336_/Y sky130_fd_sc_hd__nand2_4
X_61614_ _61607_/Y _61610_/Y _61583_/Y _61611_/Y _61613_/Y _61614_/X
+ sky130_fd_sc_hd__a41o_4
X_68170_ _67061_/X _67065_/X _68169_/X _68170_/Y sky130_fd_sc_hd__a21oi_4
X_46548_ _86727_/Q _46543_/X _46547_/Y _46548_/Y sky130_fd_sc_hd__o21ai_4
X_65382_ _44150_/X _86723_/Q _64980_/X _65381_/X _65383_/C sky130_fd_sc_hd__a211o_4
X_77368_ _82220_/Q _77367_/X _77387_/B sky130_fd_sc_hd__xnor2_4
X_62594_ _62551_/X _62553_/X _84398_/Q _62594_/Y sky130_fd_sc_hd__nor3_4
X_67121_ _67120_/X _67121_/X sky130_fd_sc_hd__buf_2
X_79107_ _79107_/A _79108_/B sky130_fd_sc_hd__inv_2
X_76319_ _76319_/A _76319_/Y sky130_fd_sc_hd__inv_2
X_64333_ _64274_/A _64333_/X sky130_fd_sc_hd__buf_2
X_49267_ _49263_/A _52482_/B _49267_/Y sky130_fd_sc_hd__nand2_4
X_61545_ _61538_/Y _61541_/Y _61525_/X _61542_/Y _61544_/Y _61545_/X
+ sky130_fd_sc_hd__a41o_4
X_46479_ _86733_/Q _46474_/X _46478_/Y _46479_/Y sky130_fd_sc_hd__o21ai_4
X_77299_ _77297_/Y _77295_/X _77296_/Y _77300_/A sky130_fd_sc_hd__nand3_4
X_48218_ _48216_/Y _48194_/X _48217_/X _48218_/Y sky130_fd_sc_hd__a21oi_4
X_67052_ _67028_/A _67052_/B _67052_/X sky130_fd_sc_hd__and2_4
X_79038_ _79037_/C _79021_/A _79021_/B _79038_/Y sky130_fd_sc_hd__nand3_4
X_64264_ _64323_/A _64287_/C sky130_fd_sc_hd__buf_2
X_49198_ _86434_/Q _49153_/X _49197_/Y _49198_/Y sky130_fd_sc_hd__o21ai_4
X_61476_ _61476_/A _61518_/B sky130_fd_sc_hd__buf_2
X_66003_ _66003_/A _66004_/B sky130_fd_sc_hd__buf_2
X_63215_ _63203_/X _64422_/C _63204_/X _63239_/D _63215_/X sky130_fd_sc_hd__and4_4
X_60427_ _60427_/A _60435_/A sky130_fd_sc_hd__inv_2
X_48149_ _48143_/Y _48109_/X _48148_/X _86563_/D sky130_fd_sc_hd__a21oi_4
X_64195_ _84906_/Q _63761_/X _60895_/X _64195_/Y sky130_fd_sc_hd__o21ai_4
X_81000_ _81134_/CLK _65268_/C _75628_/A sky130_fd_sc_hd__dfxtp_4
X_51160_ _51160_/A _51160_/B _51141_/X _52853_/D _51160_/X sky130_fd_sc_hd__and4_4
X_63146_ _63144_/X _84829_/Q _63146_/C _63135_/D _63146_/X sky130_fd_sc_hd__and4_4
X_60358_ _60344_/Y _60300_/C _60284_/B _60356_/Y _60357_/Y _60358_/Y
+ sky130_fd_sc_hd__a41oi_4
X_50111_ _50109_/Y _50092_/X _50110_/X _50111_/Y sky130_fd_sc_hd__a21oi_4
X_51091_ _51097_/A _52781_/B _51091_/Y sky130_fd_sc_hd__nand2_4
X_67954_ _69779_/A _67954_/X sky130_fd_sc_hd__buf_2
X_63077_ _63039_/A _64286_/C _63028_/X _63077_/D _63077_/X sky130_fd_sc_hd__and4_4
X_60289_ _60288_/X _60325_/B sky130_fd_sc_hd__inv_2
X_50042_ _50048_/A _53255_/B _50042_/Y sky130_fd_sc_hd__nand2_4
X_66905_ _66547_/A _66905_/X sky130_fd_sc_hd__buf_2
X_62028_ _61777_/A _62046_/C sky130_fd_sc_hd__buf_2
X_82951_ _82961_/CLK _82759_/Q _82951_/Q sky130_fd_sc_hd__dfxtp_4
X_67885_ _67909_/A _67885_/B _67885_/X sky130_fd_sc_hd__and2_4
X_81902_ _81985_/CLK _81902_/D _77023_/B sky130_fd_sc_hd__dfxtp_4
X_69624_ _69768_/A _69624_/X sky130_fd_sc_hd__buf_2
X_54850_ _54850_/A _47632_/A _54850_/Y sky130_fd_sc_hd__nand2_4
X_66836_ _87124_/Q _66833_/X _66834_/X _66835_/X _66836_/X sky130_fd_sc_hd__a211o_4
X_85670_ _84815_/CLK _53245_/Y _85670_/Q sky130_fd_sc_hd__dfxtp_4
X_82882_ _82327_/CLK _78082_/B _82882_/Q sky130_fd_sc_hd__dfxtp_4
X_53801_ _71974_/B _53801_/B _53801_/Y sky130_fd_sc_hd__nand2_4
X_84621_ _84620_/CLK _60368_/X _79566_/B sky130_fd_sc_hd__dfxtp_4
X_69555_ _69626_/A _69555_/B _69555_/X sky130_fd_sc_hd__and2_4
X_81833_ _84441_/CLK _81865_/Q _77324_/A sky130_fd_sc_hd__dfxtp_4
X_54781_ _54798_/A _54788_/B _54798_/C _47511_/Y _54781_/X sky130_fd_sc_hd__and4_4
X_66767_ _66761_/X _66766_/X _66667_/X _66771_/A sky130_fd_sc_hd__a21o_4
X_51993_ _51991_/Y _51981_/X _51992_/Y _85910_/D sky130_fd_sc_hd__a21boi_4
X_63979_ _61513_/A _63947_/B _64040_/C _64025_/D _63979_/Y sky130_fd_sc_hd__nand4_4
X_56520_ _56523_/A _56520_/B _85164_/Q _56520_/Y sky130_fd_sc_hd__nand3_4
X_68506_ _87502_/Q _68504_/X _68450_/X _68505_/X _68506_/X sky130_fd_sc_hd__a211o_4
X_87340_ _87045_/CLK _87340_/D _87340_/Q sky130_fd_sc_hd__dfxtp_4
X_53732_ _85579_/Q _53729_/X _53731_/Y _53732_/Y sky130_fd_sc_hd__o21ai_4
X_65718_ _65718_/A _65718_/X sky130_fd_sc_hd__buf_2
X_84552_ _84529_/CLK _84552_/D _84552_/Q sky130_fd_sc_hd__dfxtp_4
X_50944_ _86102_/Q _50936_/X _50943_/Y _50944_/Y sky130_fd_sc_hd__o21ai_4
X_81764_ _81783_/CLK _75987_/X _81764_/Q sky130_fd_sc_hd__dfxtp_4
X_69486_ _69612_/A _69486_/B _69486_/X sky130_fd_sc_hd__and2_4
X_66698_ _66651_/A _66698_/B _66698_/X sky130_fd_sc_hd__and2_4
X_83503_ _83498_/CLK _83503_/D _83503_/Q sky130_fd_sc_hd__dfxtp_4
X_56451_ _56159_/X _56439_/X _56450_/Y _85189_/D sky130_fd_sc_hd__o21ai_4
X_80715_ _80679_/CLK _75901_/X _80683_/D sky130_fd_sc_hd__dfxtp_4
X_68437_ _68437_/A _87344_/Q _68437_/X sky130_fd_sc_hd__and2_4
X_87271_ _87782_/CLK _43780_/Y _87271_/Q sky130_fd_sc_hd__dfxtp_4
X_53663_ _53662_/X _53663_/B _53663_/Y sky130_fd_sc_hd__nand2_4
X_65649_ _65045_/A _65802_/B sky130_fd_sc_hd__buf_2
X_84483_ _84187_/CLK _61416_/Y _79151_/B sky130_fd_sc_hd__dfxtp_4
X_50875_ _86115_/Q _50856_/X _50874_/Y _50875_/Y sky130_fd_sc_hd__o21ai_4
X_81695_ _81695_/CLK _80237_/X _81695_/Q sky130_fd_sc_hd__dfxtp_4
X_55402_ _55399_/X _55400_/Y _55181_/B _55403_/B sky130_fd_sc_hd__nand3_4
X_86222_ _86222_/CLK _50332_/Y _86222_/Q sky130_fd_sc_hd__dfxtp_4
X_52614_ _52614_/A _52605_/X _52622_/C _51787_/D _52614_/X sky130_fd_sc_hd__and4_4
X_59170_ _59152_/X _59167_/Y _59168_/Y _59169_/X _59156_/X _59170_/X
+ sky130_fd_sc_hd__o32a_4
X_83434_ _83338_/CLK _71623_/X _83434_/Q sky130_fd_sc_hd__dfxtp_4
X_56382_ _56372_/X _56016_/X _56381_/Y _85215_/D sky130_fd_sc_hd__o21ai_4
X_80646_ _74777_/Y _74710_/Y DATA_FROM_HASH[3] sky130_fd_sc_hd__ebufn_2
X_68368_ _73554_/A _68365_/X _68053_/X _68367_/Y _68368_/X sky130_fd_sc_hd__a211o_4
X_53594_ _85606_/Q _53586_/X _53593_/Y _53594_/Y sky130_fd_sc_hd__o21ai_4
XPHY_204 sky130_fd_sc_hd__decap_3
X_58121_ _57997_/X _85475_/Q _58109_/X _58121_/X sky130_fd_sc_hd__o21a_4
XPHY_215 sky130_fd_sc_hd__decap_3
X_55333_ _57283_/B _44060_/X _55301_/X _55332_/X _55333_/X sky130_fd_sc_hd__a211o_4
X_67319_ _67082_/A _67320_/A sky130_fd_sc_hd__buf_2
X_86153_ _86154_/CLK _86153_/D _86153_/Q sky130_fd_sc_hd__dfxtp_4
X_52545_ _52501_/X _52545_/B _52545_/Y sky130_fd_sc_hd__nand2_4
XPHY_226 sky130_fd_sc_hd__decap_3
X_83365_ _83362_/CLK _71816_/X _83365_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_237 sky130_fd_sc_hd__decap_3
X_80577_ _80567_/X _80569_/B _80576_/Y _80596_/A sky130_fd_sc_hd__a21boi_4
X_68299_ _68338_/A _68299_/X sky130_fd_sc_hd__buf_2
Xclkbuf_6_60_0_CLK clkbuf_6_61_0_CLK/A clkbuf_6_60_0_CLK/X sky130_fd_sc_hd__clkbuf_1
XPHY_248 sky130_fd_sc_hd__decap_3
XPHY_259 sky130_fd_sc_hd__decap_3
X_85104_ _85041_/CLK _85104_/D _56989_/B sky130_fd_sc_hd__dfxtp_4
X_58052_ _57926_/X _85993_/Q _58051_/X _58052_/Y sky130_fd_sc_hd__o21ai_4
X_70330_ _70127_/X _70338_/A sky130_fd_sc_hd__buf_2
X_82316_ _86758_/CLK _77074_/B _82316_/Q sky130_fd_sc_hd__dfxtp_4
X_55264_ _55264_/A _83321_/Q _55264_/C _55264_/Y sky130_fd_sc_hd__nand3_4
X_86084_ _85764_/CLK _51046_/Y _86084_/Q sky130_fd_sc_hd__dfxtp_4
X_52476_ _52476_/A _46376_/Y _52476_/Y sky130_fd_sc_hd__nand2_4
X_40490_ _40456_/X _41563_/A _40489_/X _40490_/X sky130_fd_sc_hd__o21a_4
X_83296_ _83304_/CLK _72045_/Y _83296_/Q sky130_fd_sc_hd__dfxtp_4
X_57003_ _56738_/X _57003_/B _56740_/X _56994_/D _57004_/C sky130_fd_sc_hd__and4_4
X_54215_ _54215_/A _47442_/Y _54215_/Y sky130_fd_sc_hd__nand2_4
X_85035_ _85031_/CLK _85035_/D _85035_/Q sky130_fd_sc_hd__dfxtp_4
X_51427_ _51425_/Y _51420_/X _51426_/X _86012_/D sky130_fd_sc_hd__a21oi_4
X_70261_ _70255_/X _74751_/A _70260_/X _70261_/X sky130_fd_sc_hd__a21o_4
X_82247_ _83521_/CLK _80355_/X _82247_/Q sky130_fd_sc_hd__dfxtp_4
X_55195_ _55188_/X _83749_/Q _55193_/X _55196_/B sky130_fd_sc_hd__nand3_4
X_72000_ _47003_/A _72001_/A sky130_fd_sc_hd__buf_2
X_42160_ _42159_/Y _88004_/D sky130_fd_sc_hd__inv_2
X_54146_ _54254_/A _54146_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_584_0_CLK clkbuf_9_292_0_CLK/X _80792_/CLK sky130_fd_sc_hd__clkbuf_1
X_51358_ _51350_/A _51358_/B _51358_/Y sky130_fd_sc_hd__nand2_4
X_70192_ _83842_/Q _70192_/Y sky130_fd_sc_hd__inv_2
X_82178_ _84951_/CLK _82178_/D _82178_/Q sky130_fd_sc_hd__dfxtp_4
X_41111_ _41108_/X _41109_/X _69558_/B _41110_/X _41111_/X sky130_fd_sc_hd__a2bb2o_4
X_50309_ _50307_/Y _50243_/X _50308_/X _86226_/D sky130_fd_sc_hd__a21oi_4
X_81129_ _81125_/CLK _81129_/D _40722_/A sky130_fd_sc_hd__dfxtp_4
X_58954_ _58864_/X _58952_/Y _58953_/Y _58943_/X _58868_/X _58954_/X
+ sky130_fd_sc_hd__o32a_4
X_42091_ _42090_/Y _88039_/D sky130_fd_sc_hd__inv_2
X_54077_ _54068_/X _54077_/B _54077_/Y sky130_fd_sc_hd__nand2_4
X_51289_ _51263_/A _51289_/X sky130_fd_sc_hd__buf_2
X_86986_ _86998_/CLK _44724_/Y _86986_/Q sky130_fd_sc_hd__dfxtp_4
X_41042_ _49140_/B _41042_/X sky130_fd_sc_hd__buf_2
X_53028_ _53111_/A _53028_/X sky130_fd_sc_hd__buf_2
X_57905_ _57875_/X _85397_/Q _57904_/X _57905_/Y sky130_fd_sc_hd__o21ai_4
X_85937_ _86096_/CLK _51839_/Y _85937_/Q sky130_fd_sc_hd__dfxtp_4
X_73951_ _73829_/X _66143_/B _73951_/X sky130_fd_sc_hd__and2_4
X_58885_ _84793_/Q _58871_/X _58875_/X _58884_/X _58885_/Y sky130_fd_sc_hd__a2bb2oi_4
Xclkbuf_10_599_0_CLK clkbuf_9_299_0_CLK/X _82234_/CLK sky130_fd_sc_hd__clkbuf_1
X_72902_ _88334_/Q _72900_/X _72901_/X _72902_/Y sky130_fd_sc_hd__o21ai_4
X_45850_ _63333_/B _61676_/A sky130_fd_sc_hd__buf_2
X_57836_ _57811_/X _85402_/Q _57835_/X _57836_/Y sky130_fd_sc_hd__o21ai_4
X_76670_ _81476_/Q _76672_/B sky130_fd_sc_hd__inv_2
X_73882_ _73879_/X _73881_/X _73857_/X _73885_/A sky130_fd_sc_hd__a21o_4
X_85868_ _83562_/CLK _85868_/D _85868_/Q sky130_fd_sc_hd__dfxtp_4
X_44801_ _44512_/A _41887_/A _41441_/X _86946_/Q _44516_/A _44802_/A
+ sky130_fd_sc_hd__o32ai_4
X_75621_ _75621_/A _80775_/D _75621_/X sky130_fd_sc_hd__or2_4
X_87607_ _87073_/CLK _87607_/D _87607_/Q sky130_fd_sc_hd__dfxtp_4
X_72833_ _72826_/X _72832_/X _72737_/X _72848_/B sky130_fd_sc_hd__a21o_4
X_84819_ _83451_/CLK _84819_/D _84819_/Q sky130_fd_sc_hd__dfxtp_4
X_45781_ _85096_/Q _44880_/X _45780_/X _45781_/Y sky130_fd_sc_hd__o21ai_4
X_57767_ _64567_/A _58784_/A sky130_fd_sc_hd__buf_2
X_42993_ _51949_/A _52021_/A sky130_fd_sc_hd__buf_2
X_54979_ _54964_/A _54978_/X _54974_/C _47558_/A _54979_/X sky130_fd_sc_hd__and4_4
X_85799_ _86119_/CLK _52554_/Y _65270_/B sky130_fd_sc_hd__dfxtp_4
X_47520_ _81794_/Q _47521_/A sky130_fd_sc_hd__inv_2
X_59506_ _63448_/B _58230_/A _59506_/Y sky130_fd_sc_hd__nor2_4
X_78340_ _78325_/B _78340_/B _82756_/D sky130_fd_sc_hd__xnor2_4
X_44732_ _44707_/X _44708_/X _40729_/A _44731_/Y _44710_/X _86982_/D
+ sky130_fd_sc_hd__o32ai_4
X_56718_ _56636_/X _56706_/X _56717_/Y _85136_/D sky130_fd_sc_hd__a21o_4
X_75552_ _75517_/Y _75519_/X _75543_/X _75552_/X sky130_fd_sc_hd__a21o_4
X_87538_ _88084_/CLK _43206_/X _87538_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_522_0_CLK clkbuf_9_261_0_CLK/X _84064_/CLK sky130_fd_sc_hd__clkbuf_1
X_41944_ _41944_/A _41944_/Y sky130_fd_sc_hd__inv_2
X_72764_ _72762_/X _72738_/X _72764_/C _72764_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_6_13_0_CLK clkbuf_5_6_0_CLK/X clkbuf_7_26_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_57698_ _57698_/A _57697_/X _57698_/Y sky130_fd_sc_hd__nor2_4
X_74503_ _46272_/A _48683_/A _74503_/Y sky130_fd_sc_hd__nand2_4
X_47451_ _47451_/A _53054_/B sky130_fd_sc_hd__buf_2
X_71715_ _71714_/Y _71716_/B sky130_fd_sc_hd__buf_2
X_59437_ _58548_/A _59437_/B _59437_/Y sky130_fd_sc_hd__nor2_4
X_78271_ _78273_/A _78273_/B _78271_/X sky130_fd_sc_hd__or2_4
X_44663_ _41092_/Y _44648_/X _87011_/Q _44650_/X _87011_/D sky130_fd_sc_hd__a2bb2o_4
X_56649_ _56593_/A _56649_/X sky130_fd_sc_hd__buf_2
X_75483_ _75481_/X _75482_/Y _75506_/D sky130_fd_sc_hd__and2_4
X_87469_ _87708_/CLK _87469_/D _87469_/Q sky130_fd_sc_hd__dfxtp_4
X_41875_ _57491_/B _50731_/A _40573_/X _88114_/Q _41872_/X _41875_/Y
+ sky130_fd_sc_hd__o32ai_4
X_72695_ _72697_/A _72697_/B _55426_/X _72695_/Y sky130_fd_sc_hd__nand3_4
X_46402_ _48631_/A _47904_/A sky130_fd_sc_hd__buf_2
X_77222_ _77222_/A _77222_/B _77222_/Y sky130_fd_sc_hd__nand2_4
X_43614_ _43614_/A _68495_/B sky130_fd_sc_hd__inv_2
X_74434_ _83067_/Q _74412_/X _74433_/Y _74434_/Y sky130_fd_sc_hd__o21ai_4
X_40826_ _40826_/A _40826_/X sky130_fd_sc_hd__buf_2
X_47382_ _47382_/A _47382_/X sky130_fd_sc_hd__buf_2
X_71646_ _71241_/A _71261_/B _71644_/C _71646_/Y sky130_fd_sc_hd__nand3_4
X_59368_ _59085_/A _59368_/X sky130_fd_sc_hd__buf_2
X_44594_ _44530_/A _44594_/X sky130_fd_sc_hd__buf_2
X_49121_ _49121_/A _53902_/B sky130_fd_sc_hd__buf_2
X_46333_ _83650_/Q _53976_/B sky130_fd_sc_hd__inv_2
Xclkbuf_10_537_0_CLK clkbuf_9_268_0_CLK/X _84079_/CLK sky130_fd_sc_hd__clkbuf_1
X_58319_ _58319_/A _58320_/A sky130_fd_sc_hd__inv_2
X_77153_ _77174_/B _81920_/Q _77173_/A sky130_fd_sc_hd__xor2_4
Xclkbuf_6_28_0_CLK clkbuf_6_29_0_CLK/A clkbuf_7_57_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_43545_ _43166_/A _43760_/A sky130_fd_sc_hd__buf_2
X_74365_ _71964_/A _74366_/C sky130_fd_sc_hd__buf_2
X_40757_ _40753_/X _40754_/X _88341_/Q _40756_/X _88341_/D sky130_fd_sc_hd__a2bb2o_4
X_59299_ _59238_/X _86345_/Q _59299_/Y sky130_fd_sc_hd__nor2_4
X_71577_ _71576_/X _71583_/B _71574_/C _71577_/Y sky130_fd_sc_hd__nor3_4
X_76104_ _81531_/Q _76104_/B _76104_/X sky130_fd_sc_hd__xor2_4
X_49052_ _49052_/A _49052_/X sky130_fd_sc_hd__buf_2
X_61330_ _84856_/Q _61330_/X sky130_fd_sc_hd__buf_2
X_73316_ _73314_/X _73315_/Y _73221_/X _73316_/Y sky130_fd_sc_hd__a21oi_4
X_70528_ _70410_/Y _71507_/A sky130_fd_sc_hd__buf_2
X_46264_ _46349_/A _46328_/B sky130_fd_sc_hd__buf_2
X_77084_ _77084_/A _77083_/X _77084_/Y sky130_fd_sc_hd__nand2_4
X_43476_ _43472_/X _43475_/X _41676_/X _87403_/Q _43456_/X _43477_/A
+ sky130_fd_sc_hd__o32ai_4
X_74296_ _70277_/C _74288_/X _74295_/Y _74296_/X sky130_fd_sc_hd__a21bo_4
X_40688_ _40836_/A _40688_/X sky130_fd_sc_hd__buf_2
X_48003_ _53535_/B _50310_/B sky130_fd_sc_hd__buf_2
X_45215_ _45215_/A _45216_/A sky130_fd_sc_hd__inv_2
X_76035_ _76023_/Y _76034_/X _76038_/A sky130_fd_sc_hd__nand2_4
X_42427_ _42427_/A _42427_/Y sky130_fd_sc_hd__inv_2
X_61261_ _72564_/A _72544_/B sky130_fd_sc_hd__buf_2
X_73247_ _73247_/A _73196_/B _73247_/Y sky130_fd_sc_hd__nor2_4
X_46195_ _46195_/A _46162_/C _46217_/B _46195_/D _46195_/Y sky130_fd_sc_hd__nand4_4
X_70459_ _70455_/Y _71337_/A sky130_fd_sc_hd__buf_2
X_63000_ _59450_/Y _62999_/X _61315_/A _60555_/A _63000_/X sky130_fd_sc_hd__a2bb2o_4
X_60212_ _60212_/A _60300_/B sky130_fd_sc_hd__buf_2
X_45146_ _45138_/X _45142_/Y _45145_/Y _45146_/Y sky130_fd_sc_hd__a21oi_4
X_42358_ _41731_/X _42356_/X _87904_/Q _42357_/X _87904_/D sky130_fd_sc_hd__a2bb2o_4
X_61192_ _61234_/A _61165_/B _61192_/C _61192_/Y sky130_fd_sc_hd__nor3_4
X_73178_ _69780_/B _73227_/A _72979_/X _73177_/Y _73178_/X sky130_fd_sc_hd__a211o_4
X_41309_ _41306_/X _41307_/X _67444_/B _41308_/X _41309_/X sky130_fd_sc_hd__a2bb2o_4
X_60143_ _60042_/A _59988_/Y _60141_/Y _79937_/A _59802_/X _60143_/X
+ sky130_fd_sc_hd__a32o_4
X_72129_ _72129_/A _72193_/B _72129_/Y sky130_fd_sc_hd__nor2_4
X_49954_ _49950_/Y _49951_/X _49953_/X _86293_/D sky130_fd_sc_hd__a21oi_4
X_45077_ _85206_/Q _45027_/X _45076_/X _45077_/Y sky130_fd_sc_hd__o21ai_4
X_42289_ _51584_/A _42290_/A sky130_fd_sc_hd__buf_2
X_77986_ _82254_/Q _81966_/Q _77999_/B sky130_fd_sc_hd__xnor2_4
X_48905_ _81215_/Q _48976_/A _48905_/Y sky130_fd_sc_hd__nor2_4
X_44028_ _69654_/A _64731_/A sky130_fd_sc_hd__buf_2
X_79725_ _79702_/X _79715_/X _79725_/Y sky130_fd_sc_hd__nand2_4
X_64951_ _64924_/A _64951_/B _64951_/X sky130_fd_sc_hd__and2_4
X_60074_ _59508_/X _60074_/X sky130_fd_sc_hd__buf_2
X_76937_ _76932_/Y _76914_/B _76936_/Y _76938_/B sky130_fd_sc_hd__o21ai_4
X_49885_ _49883_/Y _49870_/X _49884_/X _49885_/Y sky130_fd_sc_hd__a21oi_4
X_63902_ _57660_/X _63902_/B _63902_/C _63902_/D _63903_/D sky130_fd_sc_hd__nand4_4
X_48836_ _48836_/A _48836_/X sky130_fd_sc_hd__buf_2
X_67670_ _67550_/X _67670_/X sky130_fd_sc_hd__buf_2
X_79656_ _79648_/X _79650_/B _79655_/Y _79660_/A sky130_fd_sc_hd__a21boi_4
X_64882_ _64752_/X _86167_/Q _64716_/X _64881_/X _64882_/X sky130_fd_sc_hd__a211o_4
X_76868_ _76858_/A _76857_/Y _81496_/Q _81368_/D _76868_/X sky130_fd_sc_hd__a2bb2o_4
X_66621_ _69853_/A _66621_/B _66621_/X sky130_fd_sc_hd__and2_4
X_78607_ _82518_/Q _82774_/D _82486_/D sky130_fd_sc_hd__xor2_4
X_75819_ _75817_/Y _75818_/A _75820_/A sky130_fd_sc_hd__nand2_4
X_63833_ _63578_/A _63833_/X sky130_fd_sc_hd__buf_2
X_48767_ _48764_/Y _48760_/X _48766_/X _86487_/D sky130_fd_sc_hd__a21oi_4
X_79587_ _79587_/A _79587_/B _79594_/B sky130_fd_sc_hd__nand2_4
X_45979_ _40417_/Y _45974_/X _86829_/Q _45976_/X _86829_/D sky130_fd_sc_hd__a2bb2o_4
X_76799_ _81489_/Q _81361_/D _76798_/X _76800_/B sky130_fd_sc_hd__o21ai_4
X_69340_ _64789_/A _69340_/X sky130_fd_sc_hd__buf_2
X_47718_ _47715_/X _53205_/B _47718_/Y sky130_fd_sc_hd__nand2_4
X_66552_ _69183_/A _66552_/X sky130_fd_sc_hd__buf_2
X_78538_ _78529_/Y _78511_/X _78538_/X sky130_fd_sc_hd__and2_4
X_63764_ _64184_/C _63765_/C sky130_fd_sc_hd__buf_2
X_60976_ _60954_/X _61012_/C _61012_/A _60976_/Y sky130_fd_sc_hd__a21boi_4
X_48698_ _48631_/A _48699_/B sky130_fd_sc_hd__buf_2
X_65503_ _64828_/A _65503_/X sky130_fd_sc_hd__buf_2
X_62715_ _62727_/A _62727_/B _61811_/X _62715_/Y sky130_fd_sc_hd__nand3_4
X_69271_ _69191_/A _87785_/Q _69271_/X sky130_fd_sc_hd__and2_4
X_47649_ _47649_/A _53167_/B _47649_/Y sky130_fd_sc_hd__nand2_4
X_66483_ _66377_/A _66483_/X sky130_fd_sc_hd__buf_2
X_78469_ _78469_/A _82765_/D _78469_/X sky130_fd_sc_hd__xor2_4
X_63695_ _59439_/Y _63626_/X _61676_/A _63627_/X _63695_/X sky130_fd_sc_hd__a2bb2o_4
X_80500_ _80482_/Y _80485_/Y _80500_/X sky130_fd_sc_hd__or2_4
X_68222_ _67372_/X _67374_/X _68209_/X _68222_/Y sky130_fd_sc_hd__a21oi_4
X_65434_ _64967_/X _65449_/A sky130_fd_sc_hd__buf_2
X_50660_ _52355_/A _50651_/X _50668_/C _50660_/X sky130_fd_sc_hd__and3_4
X_62646_ _61301_/X _62646_/B _60291_/C _60227_/A _62646_/Y sky130_fd_sc_hd__nand4_4
X_81480_ _81344_/CLK _84048_/Q _76709_/B sky130_fd_sc_hd__dfxtp_4
X_49319_ _49315_/Y _49316_/X _49318_/X _86411_/D sky130_fd_sc_hd__a21oi_4
X_80431_ _59229_/Y _66193_/C _80430_/Y _80448_/B sky130_fd_sc_hd__o21a_4
X_68153_ _68097_/X _66958_/Y _68148_/X _68152_/Y _68153_/X sky130_fd_sc_hd__a211o_4
X_65365_ _65362_/X _85508_/Q _65363_/X _65364_/X _65365_/X sky130_fd_sc_hd__a211o_4
X_50591_ _86171_/Q _50499_/X _50590_/Y _50591_/Y sky130_fd_sc_hd__o21ai_4
X_62577_ _45308_/A _62577_/Y sky130_fd_sc_hd__inv_2
X_67104_ _67131_/A _67104_/B _67104_/X sky130_fd_sc_hd__and2_4
X_52330_ _52334_/A _49015_/X _52330_/Y sky130_fd_sc_hd__nand2_4
X_64316_ _59392_/A _64316_/B _64316_/Y sky130_fd_sc_hd__nor2_4
X_83150_ _86218_/CLK _83150_/D _83150_/Q sky130_fd_sc_hd__dfxtp_4
X_61528_ _61528_/A _61542_/B _61542_/C _61512_/X _61528_/Y sky130_fd_sc_hd__nand4_4
X_80362_ _80362_/A _80366_/A sky130_fd_sc_hd__inv_2
X_68084_ _87136_/Q _68059_/X _67991_/X _68083_/X _68084_/X sky130_fd_sc_hd__a211o_4
X_65296_ _65296_/A _65296_/X sky130_fd_sc_hd__buf_2
X_82101_ _82047_/CLK _82101_/D _82101_/Q sky130_fd_sc_hd__dfxtp_4
X_67035_ _66915_/A _67035_/X sky130_fd_sc_hd__buf_2
X_52261_ _52618_/A _52262_/A sky130_fd_sc_hd__buf_2
X_64247_ _64306_/A _64248_/B sky130_fd_sc_hd__buf_2
X_83081_ _86525_/CLK _83081_/D _83081_/Q sky130_fd_sc_hd__dfxtp_4
X_61459_ _72561_/C _61459_/X sky130_fd_sc_hd__buf_2
X_80293_ _80293_/A _80293_/Y sky130_fd_sc_hd__inv_2
X_54000_ _53991_/A _52480_/B _54000_/Y sky130_fd_sc_hd__nand2_4
X_51212_ _51212_/A _47184_/X _51212_/Y sky130_fd_sc_hd__nand2_4
X_82032_ _82005_/CLK _77862_/B _82032_/Q sky130_fd_sc_hd__dfxtp_4
X_52192_ _50537_/A _52247_/A sky130_fd_sc_hd__buf_2
X_64178_ _63703_/B _64190_/B _64178_/C _64190_/D _64181_/B sky130_fd_sc_hd__nand4_4
X_51143_ _51140_/Y _51119_/X _51142_/X _86066_/D sky130_fd_sc_hd__a21oi_4
X_63129_ _84351_/Q _63072_/X _63128_/Y _84351_/D sky130_fd_sc_hd__a21o_4
X_86840_ _86841_/CLK _86840_/D _86840_/Q sky130_fd_sc_hd__dfxtp_4
X_68986_ _68982_/X _68985_/X _68986_/Y sky130_fd_sc_hd__nand2_4
X_51074_ _51074_/A _51129_/A sky130_fd_sc_hd__buf_2
X_55951_ _55948_/X _55950_/X _55615_/A _55954_/A sky130_fd_sc_hd__a21o_4
X_67937_ _87962_/Q _67888_/X _67865_/X _67936_/X _67937_/X sky130_fd_sc_hd__a211o_4
X_86771_ _84276_/CLK _86771_/D _43175_/B sky130_fd_sc_hd__dfxtp_4
X_83983_ _87671_/CLK _83983_/D _83983_/Q sky130_fd_sc_hd__dfxtp_4
X_50025_ _50025_/A _50040_/B _50025_/C _53238_/D _50025_/X sky130_fd_sc_hd__and4_4
X_54902_ _54899_/Y _54882_/X _54901_/X _85357_/D sky130_fd_sc_hd__a21oi_4
X_85722_ _84746_/CLK _85722_/D _85722_/Q sky130_fd_sc_hd__dfxtp_4
X_58670_ _58666_/Y _58669_/Y _58646_/X _58670_/X sky130_fd_sc_hd__a21o_4
X_82934_ _82933_/CLK _78278_/X _46380_/A sky130_fd_sc_hd__dfxtp_4
X_67868_ _67987_/A _67868_/X sky130_fd_sc_hd__buf_2
X_55882_ _55882_/A _74317_/C sky130_fd_sc_hd__buf_2
X_57621_ _57630_/A _53588_/B _57621_/Y sky130_fd_sc_hd__nand2_4
X_69607_ _69607_/A _69607_/X sky130_fd_sc_hd__buf_2
X_54833_ _54823_/A _47598_/A _54833_/Y sky130_fd_sc_hd__nand2_4
X_85653_ _85431_/CLK _53335_/Y _85653_/Q sky130_fd_sc_hd__dfxtp_4
X_66819_ _66819_/A _66819_/B _66819_/X sky130_fd_sc_hd__and2_4
X_82865_ _82859_/CLK _82489_/Q _82865_/Q sky130_fd_sc_hd__dfxtp_4
X_67799_ _68429_/A _67799_/X sky130_fd_sc_hd__buf_2
X_84604_ _84333_/CLK _60537_/Y _79144_/A sky130_fd_sc_hd__dfxtp_4
X_57552_ _72017_/A _57552_/X sky130_fd_sc_hd__buf_2
X_81816_ _81696_/CLK _81624_/Q _81816_/Q sky130_fd_sc_hd__dfxtp_4
X_69538_ _69535_/X _69537_/X _69433_/X _69538_/Y sky130_fd_sc_hd__a21oi_4
X_88372_ _87416_/CLK _40549_/X _88372_/Q sky130_fd_sc_hd__dfxtp_4
X_54764_ _85382_/Q _54757_/X _54763_/Y _54764_/Y sky130_fd_sc_hd__o21ai_4
X_85584_ _83562_/CLK _85584_/D _85584_/Q sky130_fd_sc_hd__dfxtp_4
X_51976_ _66022_/B _51960_/X _51975_/Y _51976_/Y sky130_fd_sc_hd__o21ai_4
X_82796_ _82463_/CLK _82828_/Q _82796_/Q sky130_fd_sc_hd__dfxtp_4
X_56503_ _56510_/A _56507_/B _55857_/B _56503_/Y sky130_fd_sc_hd__nand3_4
X_87323_ _88327_/CLK _43663_/Y _43660_/A sky130_fd_sc_hd__dfxtp_4
X_53715_ _53747_/A _53715_/X sky130_fd_sc_hd__buf_2
X_84535_ _84534_/CLK _84535_/D _76983_/A sky130_fd_sc_hd__dfxtp_4
X_50927_ _86105_/Q _50910_/X _50926_/Y _50927_/Y sky130_fd_sc_hd__o21ai_4
X_81747_ _81756_/CLK _81747_/D _41703_/B sky130_fd_sc_hd__dfxtp_4
X_57483_ _44282_/X _55219_/B _57440_/A _57485_/B sky130_fd_sc_hd__or3_4
X_69469_ _69305_/A _69469_/B _69469_/X sky130_fd_sc_hd__and2_4
X_54695_ _54674_/A _54707_/B _54674_/C _47355_/Y _54695_/X sky130_fd_sc_hd__and4_4
X_71500_ _71500_/A _71256_/B _71500_/C _71500_/Y sky130_fd_sc_hd__nand3_4
X_59222_ _59208_/X _86063_/Q _59221_/X _59222_/Y sky130_fd_sc_hd__o21ai_4
X_56434_ _56130_/X _56426_/X _56433_/Y _85195_/D sky130_fd_sc_hd__o21ai_4
X_41660_ _41482_/A _41660_/X sky130_fd_sc_hd__buf_2
X_87254_ _87790_/CLK _43815_/X _87254_/Q sky130_fd_sc_hd__dfxtp_4
X_53646_ _53644_/Y _53603_/X _53645_/Y _85596_/D sky130_fd_sc_hd__a21boi_4
X_72480_ _65308_/X _85666_/Q _72422_/X _72480_/X sky130_fd_sc_hd__o21a_4
X_84466_ _84469_/CLK _61616_/Y _79134_/B sky130_fd_sc_hd__dfxtp_4
X_50858_ _50857_/X _50858_/B _50858_/Y sky130_fd_sc_hd__nand2_4
X_81678_ _81259_/CLK _80056_/X _76907_/A sky130_fd_sc_hd__dfxtp_4
X_86205_ _85884_/CLK _86205_/D _86205_/Q sky130_fd_sc_hd__dfxtp_4
X_40611_ _40568_/A _40832_/A sky130_fd_sc_hd__buf_2
X_59153_ _59238_/A _59154_/A sky130_fd_sc_hd__buf_2
X_71431_ _71420_/X _83502_/Q _71430_/X _83502_/D sky130_fd_sc_hd__a21o_4
X_83417_ _83415_/CLK _71673_/Y _83417_/Q sky130_fd_sc_hd__dfxtp_4
X_56365_ _56360_/A _56363_/B _55713_/B _56365_/Y sky130_fd_sc_hd__nand3_4
X_80629_ _80629_/A _80629_/B _80630_/B sky130_fd_sc_hd__xor2_4
X_87185_ _83753_/CLK _87185_/D _44160_/B sky130_fd_sc_hd__dfxtp_4
X_53577_ _53548_/A _48081_/Y _53577_/Y sky130_fd_sc_hd__nand2_4
X_41591_ _41588_/X _82312_/Q _41590_/X _41591_/Y sky130_fd_sc_hd__o21ai_4
X_84397_ _84393_/CLK _84397_/D _62606_/C sky130_fd_sc_hd__dfxtp_4
X_50789_ _50786_/Y _50768_/X _50788_/Y _86133_/D sky130_fd_sc_hd__a21boi_4
Xclkbuf_4_3_1_CLK clkbuf_4_3_0_CLK/X clkbuf_5_7_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_58104_ _58043_/X _85989_/Q _58103_/X _58104_/Y sky130_fd_sc_hd__o21ai_4
X_55316_ _55310_/X _55315_/X _83751_/Q _55316_/X sky130_fd_sc_hd__a21o_4
X_43330_ _43329_/X _43330_/X sky130_fd_sc_hd__buf_2
X_74150_ _74232_/A _85896_/Q _74150_/X sky130_fd_sc_hd__and2_4
X_86136_ _85529_/CLK _86136_/D _86136_/Q sky130_fd_sc_hd__dfxtp_4
X_40542_ _40541_/Y _40542_/X sky130_fd_sc_hd__buf_2
X_52528_ _52528_/A _52509_/B _52498_/C _52528_/X sky130_fd_sc_hd__and3_4
X_59084_ _64621_/A _59085_/A sky130_fd_sc_hd__buf_2
X_71362_ _71344_/X _83525_/Q _71361_/X _71362_/X sky130_fd_sc_hd__a21o_4
X_83348_ _82251_/CLK _83348_/D _83348_/Q sky130_fd_sc_hd__dfxtp_4
X_56296_ _56296_/A _56270_/B _55958_/B _56296_/Y sky130_fd_sc_hd__nand3_4
X_73101_ _73099_/X _73101_/B _73101_/C _73101_/Y sky130_fd_sc_hd__nand3_4
X_58035_ _58610_/A _58035_/X sky130_fd_sc_hd__buf_2
X_70313_ _70328_/A _70328_/B _70313_/C _70328_/D _70313_/X sky130_fd_sc_hd__and4_4
X_43261_ _43260_/X _43244_/X _41087_/X _87512_/Q _43250_/X _43261_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55247_ _85096_/Q _55272_/A _44044_/X _55246_/X _55247_/X sky130_fd_sc_hd__a211o_4
X_74081_ _73583_/A _85899_/Q _74081_/X sky130_fd_sc_hd__and2_4
X_86067_ _85748_/CLK _51138_/Y _86067_/Q sky130_fd_sc_hd__dfxtp_4
X_40473_ _40456_/X _81168_/Q _40472_/X _40473_/X sky130_fd_sc_hd__o21a_4
X_52459_ _52457_/Y _52430_/X _52458_/Y _85818_/D sky130_fd_sc_hd__a21boi_4
X_71293_ _71308_/A _71303_/A sky130_fd_sc_hd__buf_2
X_83279_ _86301_/CLK _83279_/D _83279_/Q sky130_fd_sc_hd__dfxtp_4
X_45000_ _56208_/C _44998_/X _44999_/X _45000_/Y sky130_fd_sc_hd__o21ai_4
X_42212_ _42205_/X _42200_/X _41332_/X _87978_/Q _42201_/X _42212_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73032_ _44305_/X _73372_/B sky130_fd_sc_hd__buf_2
X_85018_ _85049_/CLK _85018_/D _85018_/Q sky130_fd_sc_hd__dfxtp_4
X_70244_ _70238_/X _74797_/A _70243_/X _83824_/D sky130_fd_sc_hd__a21o_4
X_43192_ _87545_/Q _43192_/Y sky130_fd_sc_hd__inv_2
X_55178_ _45727_/A _44059_/X _55172_/X _55177_/Y _55178_/X sky130_fd_sc_hd__a211o_4
X_42143_ _42120_/X _42141_/X _41139_/X _88014_/Q _42142_/X _42143_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54129_ _54126_/Y _54117_/X _54128_/X _85499_/D sky130_fd_sc_hd__a21oi_4
X_77840_ _77825_/A _81933_/D _77839_/X _77840_/Y sky130_fd_sc_hd__o21ai_4
X_70175_ _70233_/A _70183_/D sky130_fd_sc_hd__buf_2
X_59986_ _59943_/X _62609_/D sky130_fd_sc_hd__buf_2
X_46951_ _82398_/Q _46952_/A sky130_fd_sc_hd__inv_2
X_42074_ _40964_/X _42072_/X _88046_/Q _42073_/X _42074_/X sky130_fd_sc_hd__a2bb2o_4
X_58937_ _58846_/X _85764_/Q _58847_/X _58937_/X sky130_fd_sc_hd__o21a_4
X_77771_ _81926_/D _77771_/B _77771_/Y sky130_fd_sc_hd__nand2_4
X_74983_ _74988_/A _74987_/A _74982_/Y _74983_/Y sky130_fd_sc_hd__a21boi_4
X_86969_ _87397_/CLK _86969_/D _86969_/Q sky130_fd_sc_hd__dfxtp_4
X_79510_ _79510_/A _79510_/B _79510_/Y sky130_fd_sc_hd__nand2_4
X_45902_ _45901_/X _45902_/Y sky130_fd_sc_hd__inv_2
X_41025_ _40932_/A _41091_/B sky130_fd_sc_hd__buf_2
X_76722_ _76720_/X _76709_/X _76721_/X _76722_/X sky130_fd_sc_hd__a21o_4
X_49670_ _49667_/Y _49650_/X _49669_/X _86345_/D sky130_fd_sc_hd__a21oi_4
X_73934_ _53531_/B _73933_/Y _73935_/B sky130_fd_sc_hd__xor2_4
X_46882_ _82949_/Q _54423_/D sky130_fd_sc_hd__inv_2
X_58868_ _58868_/A _58868_/X sky130_fd_sc_hd__buf_2
X_48621_ _48621_/A _52218_/A sky130_fd_sc_hd__buf_2
X_79441_ _79429_/A _79428_/Y _79440_/X _79441_/X sky130_fd_sc_hd__a21o_4
X_45833_ _45830_/X _45832_/Y _45803_/X _45833_/Y sky130_fd_sc_hd__a21oi_4
X_57819_ _57896_/A _57819_/X sky130_fd_sc_hd__buf_2
X_76653_ _76652_/Y _81394_/Q _76653_/Y sky130_fd_sc_hd__nand2_4
X_73865_ _73866_/B _73866_/C _73864_/X _73865_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_10_461_0_CLK clkbuf_9_230_0_CLK/X _85688_/CLK sky130_fd_sc_hd__clkbuf_1
X_58799_ _58795_/Y _58798_/Y _58761_/X _58799_/X sky130_fd_sc_hd__a21o_4
X_75604_ _80997_/Q _75604_/B _75604_/X sky130_fd_sc_hd__xor2_4
X_48552_ _49212_/A _48551_/X _48552_/Y sky130_fd_sc_hd__nand2_4
X_60830_ _60812_/Y _60702_/Y _59654_/X _60820_/B _60829_/Y _60830_/X
+ sky130_fd_sc_hd__a41o_4
X_72816_ _73516_/A _72816_/X sky130_fd_sc_hd__buf_2
X_79372_ _79372_/A _79372_/B _79373_/B sky130_fd_sc_hd__xor2_4
X_45764_ _45369_/A _45765_/A sky130_fd_sc_hd__buf_2
X_76584_ _76584_/A _76517_/A _76584_/C _76584_/D _76584_/X sky130_fd_sc_hd__and4_4
X_42976_ _42488_/A _42976_/X sky130_fd_sc_hd__buf_2
X_73796_ _41920_/Y _73529_/X _73698_/X _73795_/Y _73796_/X sky130_fd_sc_hd__a211o_4
X_47503_ _47513_/A _47463_/X _47513_/C _53084_/D _47503_/X sky130_fd_sc_hd__and4_4
X_78323_ _78317_/X _78335_/A _78324_/B _78323_/X sky130_fd_sc_hd__a21o_4
X_44715_ _44712_/X _44713_/X _40682_/X _86990_/Q _44714_/X _44716_/A
+ sky130_fd_sc_hd__o32ai_4
X_75535_ _75535_/A _75535_/B _75535_/Y sky130_fd_sc_hd__nor2_4
X_41927_ _42024_/A _41927_/X sky130_fd_sc_hd__buf_2
X_48483_ _73070_/B _48478_/X _48482_/Y _48483_/Y sky130_fd_sc_hd__o21ai_4
X_60761_ _60761_/A _60761_/B _84573_/Q _60761_/Y sky130_fd_sc_hd__nor3_4
X_72747_ _73183_/A _72929_/A sky130_fd_sc_hd__buf_2
X_45695_ _85134_/Q _45556_/X _45651_/X _45695_/X sky130_fd_sc_hd__o21a_4
X_62500_ _62487_/X _83245_/Q _62628_/C _62219_/X _62500_/X sky130_fd_sc_hd__and4_4
X_47434_ _86635_/Q _47429_/X _47433_/Y _47434_/Y sky130_fd_sc_hd__o21ai_4
X_78254_ _78254_/A _78252_/C _78254_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_476_0_CLK clkbuf_9_238_0_CLK/X _86089_/CLK sky130_fd_sc_hd__clkbuf_1
X_44646_ _44638_/X _44639_/X _41053_/X _87018_/Q _44640_/X _44647_/A
+ sky130_fd_sc_hd__o32ai_4
X_63480_ _59392_/A _63491_/B _63465_/C _63491_/D _63480_/Y sky130_fd_sc_hd__nand4_4
X_75466_ _75466_/A _75466_/B _75466_/X sky130_fd_sc_hd__and2_4
X_41858_ _48164_/A _48226_/A sky130_fd_sc_hd__buf_2
X_60692_ _60727_/A _60692_/X sky130_fd_sc_hd__buf_2
X_72678_ _70219_/C _72672_/X _72677_/Y _83193_/D sky130_fd_sc_hd__a21bo_4
X_77205_ _77205_/A _77202_/C _77204_/Y _77205_/X sky130_fd_sc_hd__and3_4
X_62431_ _61513_/A _62472_/B _62490_/C _62431_/D _62435_/B sky130_fd_sc_hd__nand4_4
X_74417_ _74415_/Y _74405_/X _74416_/X _83071_/D sky130_fd_sc_hd__a21oi_4
X_40809_ _40773_/X _82296_/Q _40808_/X _40810_/A sky130_fd_sc_hd__o21ai_4
X_47365_ _46612_/A _49504_/A sky130_fd_sc_hd__buf_2
X_71629_ _71527_/Y _71655_/A sky130_fd_sc_hd__inv_2
X_78185_ _78191_/B _78191_/C _78188_/A sky130_fd_sc_hd__nand2_4
X_44577_ _87048_/Q _44577_/Y sky130_fd_sc_hd__inv_2
X_75397_ _75393_/Y _75396_/C _75396_/A _75397_/Y sky130_fd_sc_hd__o21ai_4
X_41789_ _82882_/Q _48946_/A _41789_/X sky130_fd_sc_hd__or2_4
X_49104_ _49052_/A _49104_/X sky130_fd_sc_hd__buf_2
X_46316_ _86748_/Q _46292_/X _46315_/Y _46316_/Y sky130_fd_sc_hd__o21ai_4
X_65150_ _58784_/A _65673_/A sky130_fd_sc_hd__buf_2
X_77136_ _77130_/A _77129_/X _77141_/A _77136_/Y sky130_fd_sc_hd__a21boi_4
X_43528_ _43528_/A _43528_/X sky130_fd_sc_hd__buf_2
X_62362_ _62362_/A _62358_/Y _62359_/Y _62361_/Y _62362_/Y sky130_fd_sc_hd__nand4_4
X_74348_ _83089_/Q _74340_/X _74347_/Y _83089_/D sky130_fd_sc_hd__a21bo_4
X_47296_ _47291_/Y _47271_/X _47295_/X _86650_/D sky130_fd_sc_hd__a21oi_4
X_64101_ _64099_/X _64073_/X _64100_/Y _64101_/Y sky130_fd_sc_hd__a21oi_4
X_49035_ _53856_/B _52338_/B sky130_fd_sc_hd__buf_2
X_61313_ _61313_/A _72550_/C sky130_fd_sc_hd__buf_2
X_46247_ _46247_/A _46247_/Y sky130_fd_sc_hd__inv_2
XPHY_590 sky130_fd_sc_hd__decap_3
X_65081_ _65078_/X _65056_/B _65080_/X _65090_/A sky130_fd_sc_hd__nand3_4
X_77067_ _77067_/A _77067_/B _77068_/B sky130_fd_sc_hd__and2_4
X_43459_ _41626_/X _43446_/X _87412_/Q _43447_/X _87412_/D sky130_fd_sc_hd__a2bb2o_4
X_62293_ _61390_/A _62247_/X _62259_/X _62631_/D _62293_/Y sky130_fd_sc_hd__nand4_4
X_74279_ _48153_/A _74278_/Y _74279_/X sky130_fd_sc_hd__xor2_4
X_64032_ _64032_/A _64095_/B sky130_fd_sc_hd__buf_2
X_76018_ _76010_/A _76015_/A _76019_/B sky130_fd_sc_hd__and2_4
X_61244_ _72543_/A _61262_/A sky130_fd_sc_hd__buf_2
X_46178_ _44253_/X _46178_/X sky130_fd_sc_hd__buf_2
X_45129_ _45127_/X _61499_/B _45070_/X _45129_/Y sky130_fd_sc_hd__o21ai_4
X_68840_ _87584_/Q _68463_/X _68613_/X _68839_/X _68840_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_414_0_CLK clkbuf_9_207_0_CLK/X _83627_/CLK sky130_fd_sc_hd__clkbuf_1
X_61175_ _61086_/X _61162_/X _61170_/Y _61173_/Y _61174_/Y _84514_/D
+ sky130_fd_sc_hd__a41oi_4
X_60126_ _60119_/Y _60095_/X _60155_/D _60123_/Y _60125_/Y _60126_/Y
+ sky130_fd_sc_hd__a41oi_4
X_49937_ _72232_/B _49934_/X _49936_/Y _49937_/Y sky130_fd_sc_hd__o21ai_4
X_68771_ _68770_/X _87235_/Q _68771_/X sky130_fd_sc_hd__and2_4
X_65983_ _65983_/A _65982_/X _65983_/Y sky130_fd_sc_hd__nand2_4
X_77969_ _77968_/X _77970_/B sky130_fd_sc_hd__buf_2
X_67722_ _68742_/A _68644_/A sky130_fd_sc_hd__buf_2
X_79708_ _79686_/Y _79704_/X _79707_/Y _79708_/Y sky130_fd_sc_hd__a21oi_4
X_64934_ _64809_/A _64934_/X sky130_fd_sc_hd__buf_2
X_60057_ _63055_/A _60528_/A sky130_fd_sc_hd__buf_2
X_49868_ _49864_/A _53080_/B _49868_/Y sky130_fd_sc_hd__nand2_4
X_80980_ _80962_/CLK _80980_/D _75151_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_429_0_CLK clkbuf_9_214_0_CLK/X _83167_/CLK sky130_fd_sc_hd__clkbuf_1
X_48819_ _48817_/Y _48813_/X _48818_/X _86477_/D sky130_fd_sc_hd__a21oi_4
X_67653_ _87910_/Q _67651_/X _67625_/X _67652_/X _67653_/X sky130_fd_sc_hd__a211o_4
X_79639_ _79652_/A _79638_/Y _79639_/X sky130_fd_sc_hd__xor2_4
X_64865_ _64810_/A _86424_/Q _64865_/X sky130_fd_sc_hd__and2_4
X_49799_ _49688_/X _49809_/A sky130_fd_sc_hd__buf_2
X_66604_ _44012_/A _68389_/A sky130_fd_sc_hd__buf_2
X_51830_ _51820_/A _46758_/X _51830_/Y sky130_fd_sc_hd__nand2_4
X_63816_ _63809_/X _63810_/X _63812_/Y _63814_/Y _63815_/X _63816_/X
+ sky130_fd_sc_hd__a41o_4
X_82650_ _81755_/CLK _84002_/Q _79021_/A sky130_fd_sc_hd__dfxtp_4
X_67584_ _67580_/X _67583_/X _67561_/X _67584_/X sky130_fd_sc_hd__a21o_4
X_64796_ _64793_/X _64795_/X _64619_/X _64800_/A sky130_fd_sc_hd__a21o_4
X_81601_ _83940_/CLK _84201_/Q _81601_/Q sky130_fd_sc_hd__dfxtp_4
X_69323_ _87026_/Q _69277_/X _69278_/X _69322_/X _69323_/X sky130_fd_sc_hd__a211o_4
X_66535_ _69633_/A _66535_/B _66535_/X sky130_fd_sc_hd__and2_4
X_51761_ _51768_/A _51782_/B _51755_/X _51761_/D _51761_/X sky130_fd_sc_hd__and4_4
X_63747_ _61338_/A _60870_/X _63721_/C _61012_/A _63747_/Y sky130_fd_sc_hd__nand4_4
X_82581_ _82491_/CLK _82613_/Q _78213_/A sky130_fd_sc_hd__dfxtp_4
X_60959_ _60610_/A _60835_/X _60959_/C _60959_/X sky130_fd_sc_hd__or3_4
X_53500_ _53496_/Y _53498_/X _53499_/Y _53500_/Y sky130_fd_sc_hd__a21boi_4
X_84320_ _84321_/CLK _63483_/Y _80526_/B sky130_fd_sc_hd__dfxtp_4
X_50712_ _50738_/A _50712_/B _50712_/Y sky130_fd_sc_hd__nand2_4
X_81532_ _81532_/CLK _76533_/B _76113_/A sky130_fd_sc_hd__dfxtp_4
X_69254_ _87031_/Q _69182_/X _69183_/X _69253_/X _69254_/X sky130_fd_sc_hd__a211o_4
X_54480_ _54344_/A _54481_/A sky130_fd_sc_hd__buf_2
X_66466_ _66200_/X _66397_/X _66203_/C _66466_/Y sky130_fd_sc_hd__nand3_4
X_51692_ _85963_/Q _51675_/X _51691_/Y _51692_/Y sky130_fd_sc_hd__o21ai_4
X_63678_ _63624_/X _63672_/X _63673_/X _63676_/X _63677_/Y _63678_/Y
+ sky130_fd_sc_hd__o41ai_4
X_68205_ _68196_/X _67268_/Y _68189_/X _68204_/Y _68205_/X sky130_fd_sc_hd__a211o_4
X_53431_ _53351_/A _53431_/X sky130_fd_sc_hd__buf_2
X_65417_ _65416_/X _86402_/Q _65417_/X sky130_fd_sc_hd__and2_4
X_84251_ _84877_/CLK _64388_/X _79733_/B sky130_fd_sc_hd__dfxtp_4
X_50643_ _86161_/Q _50626_/X _50642_/Y _50643_/Y sky130_fd_sc_hd__o21ai_4
X_62629_ _62629_/A _62629_/Y sky130_fd_sc_hd__inv_2
X_81463_ _81431_/CLK _76845_/B _81463_/Q sky130_fd_sc_hd__dfxtp_4
X_69185_ _87036_/Q _69182_/X _69183_/X _69184_/X _69186_/B sky130_fd_sc_hd__a211o_4
X_66397_ _66104_/A _66397_/X sky130_fd_sc_hd__buf_2
X_83202_ _83843_/CLK _83202_/D _70193_/A sky130_fd_sc_hd__dfxtp_4
X_80414_ _80412_/X _80413_/X _80414_/Y sky130_fd_sc_hd__xnor2_4
X_56150_ _56140_/A _56150_/B _55761_/B _56150_/Y sky130_fd_sc_hd__nand3_4
X_68136_ _82070_/D _68120_/X _68135_/X _68136_/X sky130_fd_sc_hd__a21bo_4
X_53362_ _53339_/A _53371_/B _53371_/C _52846_/D _53362_/X sky130_fd_sc_hd__and4_4
X_65348_ _65268_/A _65294_/B _65348_/C _65348_/X sky130_fd_sc_hd__and3_4
X_84182_ _83507_/CLK _84182_/D _84182_/Q sky130_fd_sc_hd__dfxtp_4
X_50574_ _50571_/Y _50474_/X _50573_/Y _86175_/D sky130_fd_sc_hd__a21boi_4
X_81394_ _83932_/CLK _83930_/Q _81394_/Q sky130_fd_sc_hd__dfxtp_4
X_55101_ _85318_/Q _55098_/X _55100_/Y _55101_/Y sky130_fd_sc_hd__o21ai_4
X_52313_ _85847_/Q _52297_/X _52312_/Y _52313_/Y sky130_fd_sc_hd__o21ai_4
X_83133_ _83133_/CLK _73868_/Y _83133_/Q sky130_fd_sc_hd__dfxtp_4
X_56081_ _56058_/X _56079_/X _56080_/Y _85299_/D sky130_fd_sc_hd__o21ai_4
X_80345_ _84751_/Q _84143_/Q _80360_/B sky130_fd_sc_hd__nand2_4
X_68067_ _68437_/A _68067_/B _68067_/X sky130_fd_sc_hd__and2_4
X_53293_ _53293_/A _53293_/B _53293_/C _52779_/D _53293_/X sky130_fd_sc_hd__and4_4
X_65279_ _65206_/A _65279_/B _65279_/X sky130_fd_sc_hd__and2_4
X_55032_ _55029_/Y _55024_/X _55031_/X _85332_/D sky130_fd_sc_hd__a21oi_4
X_67018_ _80911_/D _66971_/X _67017_/X _84087_/D sky130_fd_sc_hd__a21bo_4
X_52244_ _52242_/Y _52232_/X _52243_/X _85861_/D sky130_fd_sc_hd__a21oi_4
X_83064_ _86498_/CLK _83064_/D _83064_/Q sky130_fd_sc_hd__dfxtp_4
X_87941_ _88387_/CLK _87941_/D _87941_/Q sky130_fd_sc_hd__dfxtp_4
X_80276_ _80279_/B _80276_/Y sky130_fd_sc_hd__inv_2
X_82015_ _82015_/CLK _82015_/D _77217_/A sky130_fd_sc_hd__dfxtp_4
X_59840_ _59840_/A _59840_/Y sky130_fd_sc_hd__inv_2
X_52175_ _52175_/A _52194_/B _52182_/C _52175_/X sky130_fd_sc_hd__and3_4
X_87872_ _88128_/CLK _87872_/D _87872_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_41_0_CLK clkbuf_8_41_0_CLK/A clkbuf_9_83_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_51126_ _51124_/Y _51119_/X _51125_/X _51126_/Y sky130_fd_sc_hd__a21oi_4
X_86823_ _88245_/CLK _86823_/D _66938_/B sky130_fd_sc_hd__dfxtp_4
X_59771_ _65044_/A _59771_/X sky130_fd_sc_hd__buf_2
X_56983_ _56684_/C _57149_/B sky130_fd_sc_hd__buf_2
X_68969_ _68966_/X _68968_/X _68922_/X _68969_/X sky130_fd_sc_hd__a21o_4
X_58722_ _58722_/A _58764_/B _58722_/Y sky130_fd_sc_hd__nor2_4
X_51057_ _51054_/Y _51039_/X _51056_/X _51057_/Y sky130_fd_sc_hd__a21oi_4
X_55934_ _44085_/C _55934_/B _55934_/X sky130_fd_sc_hd__and2_4
X_86754_ _83115_/CLK _86754_/D _86754_/Q sky130_fd_sc_hd__dfxtp_4
X_71980_ _71977_/Y _71978_/X _71979_/X _71980_/Y sky130_fd_sc_hd__a21oi_4
X_83966_ _81994_/CLK _83966_/D _80822_/D sky130_fd_sc_hd__dfxtp_4
X_50008_ _72400_/B _49986_/X _50007_/Y _50008_/Y sky130_fd_sc_hd__o21ai_4
X_85705_ _86686_/CLK _53059_/Y _85705_/Q sky130_fd_sc_hd__dfxtp_4
X_70931_ _46912_/X _70909_/A _70930_/Y _70931_/Y sky130_fd_sc_hd__o21ai_4
X_58653_ _58653_/A _58653_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_56_0_CLK clkbuf_8_57_0_CLK/A clkbuf_8_56_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_82917_ _82931_/CLK _78153_/X _46567_/A sky130_fd_sc_hd__dfxtp_4
X_55865_ _55549_/A _55865_/B _55865_/X sky130_fd_sc_hd__and2_4
X_86685_ _86686_/CLK _86685_/D _86685_/Q sky130_fd_sc_hd__dfxtp_4
X_83897_ _82299_/CLK _83897_/D _81969_/D sky130_fd_sc_hd__dfxtp_4
X_57604_ _72017_/A _57630_/A sky130_fd_sc_hd__buf_2
X_54816_ _54825_/A _54816_/B _54831_/C _53125_/D _54816_/X sky130_fd_sc_hd__and4_4
X_42830_ _42820_/X _42830_/X sky130_fd_sc_hd__buf_2
X_73650_ _73650_/A _73649_/X _73650_/Y sky130_fd_sc_hd__nor2_4
X_85636_ _86054_/CLK _53425_/Y _85636_/Q sky130_fd_sc_hd__dfxtp_4
X_70862_ _70862_/A _70869_/D sky130_fd_sc_hd__buf_2
X_58584_ _84816_/Q _58095_/X _58578_/X _58583_/X _58584_/Y sky130_fd_sc_hd__a2bb2oi_4
X_82848_ _82152_/CLK _82848_/D _82848_/Q sky130_fd_sc_hd__dfxtp_4
X_55796_ _55793_/X _55795_/X _44110_/X _55796_/X sky130_fd_sc_hd__a21o_4
X_72601_ _83221_/Q _72445_/X _72588_/Y _72600_/Y _72601_/Y sky130_fd_sc_hd__a2bb2oi_4
X_57535_ _57531_/A _53504_/B _57535_/Y sky130_fd_sc_hd__nand2_4
X_42761_ _42739_/X _42740_/X _41277_/X _87733_/Q _42750_/X _42762_/A
+ sky130_fd_sc_hd__o32ai_4
X_88355_ _88363_/CLK _88355_/D _88355_/Q sky130_fd_sc_hd__dfxtp_4
X_54747_ _54693_/X _54747_/X sky130_fd_sc_hd__buf_2
X_73581_ _87006_/Q _57092_/X _73580_/X _73581_/Y sky130_fd_sc_hd__o21ai_4
X_85567_ _83307_/CLK _85567_/D _85567_/Q sky130_fd_sc_hd__dfxtp_4
X_51959_ _51955_/Y _51951_/X _51958_/X _51959_/Y sky130_fd_sc_hd__a21oi_4
X_70793_ _70824_/A _70905_/A sky130_fd_sc_hd__buf_2
X_82779_ _82206_/CLK _82779_/D _82779_/Q sky130_fd_sc_hd__dfxtp_4
X_44500_ _44500_/A _44500_/Y sky130_fd_sc_hd__inv_2
X_75320_ _75320_/A _81075_/Q _75320_/Y sky130_fd_sc_hd__nand2_4
X_87306_ _83158_/CLK _87306_/D _87306_/Q sky130_fd_sc_hd__dfxtp_4
X_41712_ _41712_/A _41712_/Y sky130_fd_sc_hd__inv_2
X_72532_ _72569_/A _72531_/Y _61202_/A _72532_/X sky130_fd_sc_hd__a21o_4
X_84518_ _84518_/CLK _61139_/Y _84518_/Q sky130_fd_sc_hd__dfxtp_4
X_45480_ _85148_/Q _45464_/X _44919_/X _45480_/Y sky130_fd_sc_hd__o21ai_4
X_57466_ _57440_/X _57464_/X _57465_/X _57466_/Y sky130_fd_sc_hd__o21ai_4
X_88286_ _87253_/CLK _41056_/Y _69431_/B sky130_fd_sc_hd__dfxtp_4
X_42692_ _42692_/A _42692_/Y sky130_fd_sc_hd__inv_2
X_54678_ _54682_/A _47324_/A _54678_/Y sky130_fd_sc_hd__nand2_4
X_85498_ _83745_/CLK _85498_/D _85498_/Q sky130_fd_sc_hd__dfxtp_4
X_59205_ _59081_/A _59205_/X sky130_fd_sc_hd__buf_2
X_44431_ _44363_/X _44431_/X sky130_fd_sc_hd__buf_2
X_56417_ _56085_/X _56409_/X _56416_/Y _56417_/Y sky130_fd_sc_hd__o21ai_4
X_75251_ _75251_/A _81070_/Q _75251_/Y sky130_fd_sc_hd__nand2_4
X_87237_ _88012_/CLK _87237_/D _68718_/B sky130_fd_sc_hd__dfxtp_4
X_41643_ _41642_/Y _41643_/X sky130_fd_sc_hd__buf_2
X_53629_ _85599_/Q _53626_/X _53628_/Y _53629_/Y sky130_fd_sc_hd__o21ai_4
X_72463_ _57800_/X _72461_/Y _72462_/Y _64761_/B _59833_/X _72463_/X
+ sky130_fd_sc_hd__o32a_4
X_84449_ _84449_/CLK _61866_/Y _78072_/B sky130_fd_sc_hd__dfxtp_4
X_57397_ _57359_/A _57397_/B _57372_/X _57397_/Y sky130_fd_sc_hd__nor3_4
X_74202_ _74202_/A _74201_/Y _74202_/Y sky130_fd_sc_hd__nor2_4
X_47150_ _47150_/A _52881_/B _47150_/Y sky130_fd_sc_hd__nand2_4
X_59136_ _59135_/X _85654_/Q _59070_/X _59136_/X sky130_fd_sc_hd__o21a_4
X_71414_ _71396_/Y _83507_/Q _71413_/Y _71414_/X sky130_fd_sc_hd__a21o_4
X_44362_ _44362_/A _46298_/A sky130_fd_sc_hd__buf_2
X_56348_ _56358_/A _56345_/B _55774_/B _56348_/Y sky130_fd_sc_hd__nand3_4
X_75182_ _75182_/A _75181_/Y _81033_/D sky130_fd_sc_hd__xnor2_4
X_41574_ _41573_/X _41574_/X sky130_fd_sc_hd__buf_2
X_87168_ _87169_/CLK _44320_/Y _43950_/A sky130_fd_sc_hd__dfxtp_4
X_72394_ _72394_/A _72394_/Y sky130_fd_sc_hd__inv_2
X_46101_ _46101_/A _46214_/D sky130_fd_sc_hd__buf_2
X_43313_ _43296_/X _43305_/X _41225_/X _87486_/Q _43308_/X _43314_/A
+ sky130_fd_sc_hd__o32ai_4
X_74133_ _73566_/X _84969_/Q _74087_/X _74132_/X _74133_/X sky130_fd_sc_hd__a211o_4
X_86119_ _86119_/CLK _86119_/D _86119_/Q sky130_fd_sc_hd__dfxtp_4
X_40525_ _40524_/X _40508_/X _88377_/Q _40510_/X _88377_/D sky130_fd_sc_hd__a2bb2o_4
X_47081_ _47081_/A _47081_/X sky130_fd_sc_hd__buf_2
X_59067_ _58897_/A _59068_/B sky130_fd_sc_hd__buf_2
X_71345_ _71462_/B _71418_/B sky130_fd_sc_hd__buf_2
X_44293_ _44268_/A _44293_/B _72498_/B _44293_/Y sky130_fd_sc_hd__nand3_4
X_56279_ _56279_/A _57223_/D _56174_/X _56281_/A sky130_fd_sc_hd__nand3_4
X_79990_ _79964_/Y _79982_/A _79990_/Y sky130_fd_sc_hd__nor2_4
X_87099_ _88272_/CLK _44459_/X _87099_/Q sky130_fd_sc_hd__dfxtp_4
X_46032_ _43030_/A _46032_/X sky130_fd_sc_hd__buf_2
X_58018_ _57903_/X _85484_/Q _57962_/X _58018_/X sky130_fd_sc_hd__o21a_4
X_43244_ _43167_/A _43244_/X sky130_fd_sc_hd__buf_2
X_74064_ _72730_/X _84972_/Q _74021_/X _74063_/X _74065_/B sky130_fd_sc_hd__a211o_4
X_78941_ _82849_/Q _82561_/Q _78953_/A sky130_fd_sc_hd__xnor2_4
X_40456_ _40783_/A _40456_/X sky130_fd_sc_hd__buf_2
X_71276_ _71175_/A _71276_/B _71276_/C _71276_/D _71276_/Y sky130_fd_sc_hd__nand4_4
X_73015_ _73238_/A _73015_/X sky130_fd_sc_hd__buf_2
X_70227_ _70229_/A _70229_/B _83190_/Q _70229_/D _70227_/X sky130_fd_sc_hd__and4_4
X_43175_ _43175_/A _43175_/B _43175_/C _43175_/X sky130_fd_sc_hd__and3_4
X_78872_ _78886_/A _78896_/A _78881_/A sky130_fd_sc_hd__xor2_4
X_40387_ _40386_/Y _40387_/X sky130_fd_sc_hd__buf_2
X_42126_ _41912_/A _42126_/X sky130_fd_sc_hd__buf_2
X_77823_ _77835_/A _77822_/Y _77824_/B sky130_fd_sc_hd__xor2_4
X_70158_ _83849_/Q _70158_/Y sky130_fd_sc_hd__inv_2
X_47983_ _47971_/X _82931_/Q _47982_/X _47984_/B sky130_fd_sc_hd__o21ai_4
X_59969_ _59968_/X _59969_/X sky130_fd_sc_hd__buf_2
X_49722_ _57731_/B _49715_/X _49721_/Y _49722_/Y sky130_fd_sc_hd__o21ai_4
X_46934_ _46915_/X _46896_/B _46926_/C _52758_/D _46934_/X sky130_fd_sc_hd__and4_4
X_42057_ _42057_/A _42057_/Y sky130_fd_sc_hd__inv_2
X_77754_ _82148_/Q _77754_/B _82116_/D sky130_fd_sc_hd__xor2_4
X_62980_ _58210_/X _62924_/C _60220_/A _62644_/X _62979_/X _62980_/Y
+ sky130_fd_sc_hd__a41oi_4
X_74966_ _80762_/Q _74957_/B _74966_/Y sky130_fd_sc_hd__nand2_4
X_70089_ _69071_/X _69074_/X _69156_/X _70089_/Y sky130_fd_sc_hd__a21oi_4
X_41008_ _40429_/X _40829_/B _41007_/X _41009_/A sky130_fd_sc_hd__o21a_4
X_76705_ _76697_/Y _76704_/Y _81448_/D sky130_fd_sc_hd__xor2_4
X_49653_ _49649_/Y _49650_/X _49652_/X _86348_/D sky130_fd_sc_hd__a21oi_4
X_61931_ _61949_/A _61949_/B _61949_/C _63158_/B _61931_/X sky130_fd_sc_hd__and4_4
X_73917_ _68750_/B _56939_/X _72741_/X _73917_/Y sky130_fd_sc_hd__o21ai_4
X_46865_ _46915_/A _46868_/A sky130_fd_sc_hd__buf_2
X_77685_ _77688_/B _77688_/A _77685_/X sky130_fd_sc_hd__xor2_4
X_74897_ _74897_/A _74897_/B _74899_/A _74894_/A _74897_/X sky130_fd_sc_hd__and4_4
X_48604_ _48604_/A _50508_/B _48604_/Y sky130_fd_sc_hd__nand2_4
X_79424_ _84808_/Q _66415_/C _79424_/Y sky130_fd_sc_hd__nand2_4
X_45816_ _82982_/Q _74694_/B sky130_fd_sc_hd__inv_2
X_64650_ _64817_/A _64650_/X sky130_fd_sc_hd__buf_2
X_76636_ _76636_/A _76635_/X _76637_/B sky130_fd_sc_hd__xnor2_4
X_49584_ _49582_/Y _49570_/X _49583_/X _86361_/D sky130_fd_sc_hd__a21oi_4
X_61862_ _61861_/X _61846_/B _61846_/C _61846_/D _61862_/Y sky130_fd_sc_hd__nand4_4
X_73848_ _88359_/Q _73777_/X _73656_/X _73848_/X sky130_fd_sc_hd__o21a_4
X_46796_ _46806_/A _50987_/B _46796_/Y sky130_fd_sc_hd__nand2_4
X_63601_ _63540_/A _63661_/D sky130_fd_sc_hd__buf_2
X_48535_ _48535_/A _48612_/A sky130_fd_sc_hd__buf_2
X_60813_ _60792_/A _60810_/B _84560_/Q _60813_/Y sky130_fd_sc_hd__nor3_4
X_79355_ _79332_/X _79355_/B _79355_/Y sky130_fd_sc_hd__nand2_4
X_45747_ _45744_/X _45746_/Y _45714_/X _45747_/Y sky130_fd_sc_hd__a21oi_4
X_64581_ _64577_/X _86753_/Q _64579_/X _64580_/X _64582_/B sky130_fd_sc_hd__a211o_4
X_76567_ _76563_/X _76562_/Y _76567_/Y sky130_fd_sc_hd__nand2_4
X_42959_ _42944_/X _42945_/X _40395_/X _66698_/B _42954_/X _42960_/A
+ sky130_fd_sc_hd__o32ai_4
X_61793_ _61736_/A _61863_/A sky130_fd_sc_hd__buf_2
X_73779_ _86998_/Q _73776_/X _73778_/X _73779_/Y sky130_fd_sc_hd__o21ai_4
X_66320_ _66317_/Y _66278_/X _66319_/X _84141_/D sky130_fd_sc_hd__a21o_4
X_78306_ _78302_/A _78302_/B _78306_/C _78309_/C sky130_fd_sc_hd__nand3_4
X_63532_ _63471_/A _63546_/D sky130_fd_sc_hd__buf_2
X_75518_ _75517_/Y _75519_/C sky130_fd_sc_hd__inv_2
X_60744_ _60700_/A _60752_/B _60744_/C _60744_/Y sky130_fd_sc_hd__nor3_4
X_48466_ _48457_/Y _48459_/X _48465_/X _86520_/D sky130_fd_sc_hd__a21oi_4
X_79286_ _58843_/Y _66478_/Y _79285_/Y _79286_/X sky130_fd_sc_hd__o21a_4
X_45678_ _45678_/A _45678_/X sky130_fd_sc_hd__buf_2
X_76498_ _76485_/A _76484_/Y _76513_/C _76498_/Y sky130_fd_sc_hd__o21ai_4
X_47417_ _47417_/A _53036_/D sky130_fd_sc_hd__buf_2
X_66251_ _65976_/A _66251_/X sky130_fd_sc_hd__buf_2
X_78237_ _78228_/Y _78235_/Y _78236_/Y _78237_/X sky130_fd_sc_hd__o21a_4
X_44629_ _44628_/Y _44629_/Y sky130_fd_sc_hd__inv_2
X_63463_ _63463_/A _84961_/Q _63463_/C _63463_/X sky130_fd_sc_hd__and3_4
X_75449_ _75441_/X _75467_/A _75466_/A sky130_fd_sc_hd__xnor2_4
X_48397_ _53636_/A _48364_/X _48354_/X _48397_/X sky130_fd_sc_hd__and3_4
X_60675_ _60694_/B _60654_/X _60697_/B _60804_/B _59512_/X _60675_/Y
+ sky130_fd_sc_hd__a41oi_4
X_65202_ _65199_/X _86154_/Q _65022_/X _65201_/X _65202_/X sky130_fd_sc_hd__a211o_4
X_62414_ _62410_/Y _62396_/X _62413_/Y _84412_/D sky130_fd_sc_hd__a21oi_4
X_47348_ _47348_/A _52997_/D sky130_fd_sc_hd__buf_2
X_66182_ _66125_/X _86222_/Q _66180_/X _66181_/X _66182_/X sky130_fd_sc_hd__a211o_4
X_78168_ _82670_/Q _78168_/B _78168_/X sky130_fd_sc_hd__xor2_4
X_63394_ _60720_/A _63458_/A sky130_fd_sc_hd__buf_2
X_65133_ _65035_/X _85549_/Q _65036_/X _65132_/X _65133_/X sky130_fd_sc_hd__a211o_4
X_77119_ _77127_/A _77127_/B _77122_/A sky130_fd_sc_hd__xor2_4
X_62345_ _62344_/X _57656_/X _62315_/C _62286_/X _62345_/X sky130_fd_sc_hd__and4_4
X_47279_ _47241_/X _52959_/B _47279_/Y sky130_fd_sc_hd__nand2_4
X_78099_ _78093_/Y _78098_/Y _78090_/B _78099_/Y sky130_fd_sc_hd__a21oi_4
X_49018_ _48946_/A _49018_/X sky130_fd_sc_hd__buf_2
X_80130_ _84941_/Q _84189_/Q _80130_/Y sky130_fd_sc_hd__nand2_4
X_65064_ _64834_/A _65192_/B sky130_fd_sc_hd__buf_2
X_69941_ _69832_/X _69937_/Y _69938_/X _69940_/Y _69941_/X sky130_fd_sc_hd__a211o_4
X_50290_ _86230_/Q _50282_/X _50289_/Y _50290_/Y sky130_fd_sc_hd__o21ai_4
X_62276_ _59923_/Y _62276_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_353_0_CLK clkbuf_9_176_0_CLK/X _86640_/CLK sky130_fd_sc_hd__clkbuf_1
X_64015_ _64411_/B _64029_/B _64029_/C _64015_/D _64017_/C sky130_fd_sc_hd__nand4_4
X_61227_ _61226_/X _64454_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_983_0_CLK clkbuf_9_491_0_CLK/X _83303_/CLK sky130_fd_sc_hd__clkbuf_1
X_80061_ _80059_/X _80060_/X _80074_/B sky130_fd_sc_hd__xnor2_4
X_69872_ _42041_/A _68463_/X _69478_/X _69871_/Y _69872_/X sky130_fd_sc_hd__a211o_4
X_68823_ _68823_/A _68823_/X sky130_fd_sc_hd__buf_2
X_61158_ _60933_/X _61149_/X _61154_/X _61156_/X _61157_/Y _84517_/D
+ sky130_fd_sc_hd__a41oi_4
Xclkbuf_9_474_0_CLK clkbuf_9_475_0_CLK/A clkbuf_9_474_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_60109_ _60109_/A _65607_/A sky130_fd_sc_hd__buf_2
X_83820_ _83820_/CLK _83820_/D _74764_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_368_0_CLK clkbuf_9_184_0_CLK/X _86359_/CLK sky130_fd_sc_hd__clkbuf_1
X_68754_ _69233_/A _68779_/A sky130_fd_sc_hd__buf_2
X_53980_ _53956_/X _53980_/B _53980_/Y sky130_fd_sc_hd__nand2_4
X_65966_ _65308_/X _84989_/Q _65309_/X _65965_/X _65966_/X sky130_fd_sc_hd__a211o_4
X_61089_ _72592_/A _61414_/A _61089_/C _61089_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_10_998_0_CLK clkbuf_9_499_0_CLK/X _83584_/CLK sky130_fd_sc_hd__clkbuf_1
X_67705_ _67701_/X _67704_/X _67681_/X _67705_/X sky130_fd_sc_hd__a21o_4
X_52931_ _52944_/A _52931_/B _52931_/Y sky130_fd_sc_hd__nand2_4
X_64917_ _64666_/X _86133_/Q _64766_/X _64916_/X _64917_/X sky130_fd_sc_hd__a211o_4
X_83751_ _83753_/CLK _83751_/D _83751_/Q sky130_fd_sc_hd__dfxtp_4
X_80963_ _81985_/CLK _75587_/X _75376_/B sky130_fd_sc_hd__dfxtp_4
X_68685_ _68680_/X _68682_/X _68684_/X _68685_/X sky130_fd_sc_hd__a21o_4
X_65897_ _65811_/X _83050_/Q _65865_/X _65896_/X _65897_/X sky130_fd_sc_hd__a211o_4
X_82702_ _82702_/CLK _78920_/X _82658_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_489_0_CLK clkbuf_9_489_0_CLK/A clkbuf_9_489_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_55650_ _55650_/A _55649_/Y _74539_/A sky130_fd_sc_hd__nand2_4
X_67636_ _45923_/X _68129_/A sky130_fd_sc_hd__buf_2
X_86470_ _86470_/CLK _48855_/Y _86470_/Q sky130_fd_sc_hd__dfxtp_4
X_52862_ _52860_/Y _52839_/X _52861_/X _52862_/Y sky130_fd_sc_hd__a21oi_4
X_64848_ _64948_/A _86264_/Q _64848_/X sky130_fd_sc_hd__and2_4
X_83682_ _83681_/CLK _70853_/Y _83682_/Q sky130_fd_sc_hd__dfxtp_4
X_80894_ _80961_/CLK _80894_/D _80894_/Q sky130_fd_sc_hd__dfxtp_4
X_54601_ _85412_/Q _54593_/X _54600_/Y _54601_/Y sky130_fd_sc_hd__o21ai_4
X_85421_ _85645_/CLK _54554_/Y _85421_/Q sky130_fd_sc_hd__dfxtp_4
X_51813_ _85941_/Q _51789_/X _51812_/Y _51813_/Y sky130_fd_sc_hd__o21ai_4
X_82633_ _82301_/CLK _82633_/D _78877_/B sky130_fd_sc_hd__dfxtp_4
X_55581_ _55580_/X _72648_/C sky130_fd_sc_hd__buf_2
Xclkbuf_10_921_0_CLK clkbuf_9_460_0_CLK/X _83115_/CLK sky130_fd_sc_hd__clkbuf_1
X_67567_ _84064_/Q _67449_/X _67566_/X _67567_/X sky130_fd_sc_hd__a21bo_4
X_52793_ _52767_/A _52803_/A sky130_fd_sc_hd__buf_2
X_64779_ _64650_/X _86139_/Q _64776_/X _64778_/X _64779_/X sky130_fd_sc_hd__a211o_4
X_57320_ _57318_/Y _56808_/Y _58981_/A _57319_/X _57320_/X sky130_fd_sc_hd__a211o_4
X_69306_ _87527_/Q _69205_/X _69113_/X _69305_/X _69306_/X sky130_fd_sc_hd__a211o_4
X_88140_ _88144_/CLK _88140_/D _88140_/Q sky130_fd_sc_hd__dfxtp_4
X_54532_ _54529_/Y _54530_/X _54531_/X _54532_/Y sky130_fd_sc_hd__a21oi_4
X_66518_ _65379_/X _66518_/B _65383_/C _66518_/Y sky130_fd_sc_hd__nand3_4
X_85352_ _85351_/CLK _85352_/D _85352_/Q sky130_fd_sc_hd__dfxtp_4
X_51744_ _51758_/A _51744_/B _51744_/Y sky130_fd_sc_hd__nand2_4
X_82564_ _82596_/CLK _82564_/D _78088_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_412_0_CLK clkbuf_9_413_0_CLK/A clkbuf_9_412_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_13 sky130_fd_sc_hd__decap_3
X_67498_ _87916_/Q _67473_/X _67405_/X _67497_/X _67498_/X sky130_fd_sc_hd__a211o_4
XPHY_24 sky130_fd_sc_hd__decap_3
XPHY_35 sky130_fd_sc_hd__decap_3
X_84303_ _84308_/CLK _84303_/D _80347_/B sky130_fd_sc_hd__dfxtp_4
X_57251_ _56600_/X _57247_/Y _57250_/Y _85051_/D sky130_fd_sc_hd__a21oi_4
X_81515_ _81514_/CLK _81515_/D _81515_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_46 sky130_fd_sc_hd__decap_3
X_69237_ _87532_/Q _69098_/X _69124_/X _69236_/X _69237_/X sky130_fd_sc_hd__a211o_4
X_88071_ _87553_/CLK _88071_/D _73081_/A sky130_fd_sc_hd__dfxtp_4
X_54463_ _54461_/Y _54448_/X _54462_/X _85438_/D sky130_fd_sc_hd__a21oi_4
X_66449_ _66377_/A _66449_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_306_0_CLK clkbuf_9_153_0_CLK/X _83338_/CLK sky130_fd_sc_hd__clkbuf_1
X_85283_ _83012_/CLK _85283_/D _85283_/Q sky130_fd_sc_hd__dfxtp_4
X_51675_ _51621_/A _51675_/X sky130_fd_sc_hd__buf_2
XPHY_57 sky130_fd_sc_hd__decap_3
X_82495_ _82692_/CLK _78769_/Y _82495_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_68 sky130_fd_sc_hd__decap_3
XPHY_79 sky130_fd_sc_hd__decap_3
X_56202_ _56020_/X _56195_/X _56201_/Y _85278_/D sky130_fd_sc_hd__o21ai_4
X_87022_ _87022_/CLK _87022_/D _87022_/Q sky130_fd_sc_hd__dfxtp_4
X_53414_ _53397_/A _53402_/B _53410_/C _52900_/D _53414_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_936_0_CLK clkbuf_9_468_0_CLK/X _87814_/CLK sky130_fd_sc_hd__clkbuf_1
X_84234_ _84624_/CLK _64560_/Y _79529_/B sky130_fd_sc_hd__dfxtp_4
X_50626_ _50594_/A _50626_/X sky130_fd_sc_hd__buf_2
X_57182_ _56755_/X _57023_/X _56759_/X _56877_/X _57182_/X sky130_fd_sc_hd__and4_4
X_81446_ _82053_/CLK _81446_/D _81446_/Q sky130_fd_sc_hd__dfxtp_4
X_69168_ _44245_/A _69168_/X sky130_fd_sc_hd__buf_2
X_54394_ _54366_/A _54394_/X sky130_fd_sc_hd__buf_2
X_68119_ _82074_/D _68101_/X _68118_/X _68119_/X sky130_fd_sc_hd__a21bo_4
X_56133_ _55801_/B _55801_/A _56134_/A sky130_fd_sc_hd__xnor2_4
X_53345_ _53332_/A _53345_/B _53345_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_427_0_CLK clkbuf_9_427_0_CLK/A clkbuf_9_427_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_84165_ _84166_/CLK _84165_/D _65970_/C sky130_fd_sc_hd__dfxtp_4
X_50557_ _50555_/Y _50474_/X _50556_/Y _50557_/Y sky130_fd_sc_hd__a21boi_4
X_81377_ _83940_/CLK _76949_/X _81377_/Q sky130_fd_sc_hd__dfxtp_4
X_69099_ _69357_/A _69236_/A sky130_fd_sc_hd__buf_2
X_71130_ _50712_/B _71117_/A _71129_/Y _83596_/D sky130_fd_sc_hd__o21ai_4
X_83116_ _85895_/CLK _74243_/X _70130_/B sky130_fd_sc_hd__dfxtp_4
X_56064_ _56063_/Y _56064_/X sky130_fd_sc_hd__buf_2
X_80328_ _80326_/X _80327_/Y _80328_/Y sky130_fd_sc_hd__nand2_4
X_41290_ _41143_/A _41290_/X sky130_fd_sc_hd__buf_2
X_53276_ _53276_/A _54451_/B _53276_/Y sky130_fd_sc_hd__nand2_4
X_84096_ _81169_/CLK _66806_/X _84096_/Q sky130_fd_sc_hd__dfxtp_4
X_50488_ _50486_/Y _50455_/X _50487_/X _50488_/Y sky130_fd_sc_hd__a21oi_4
X_55015_ _55011_/A _47632_/A _55015_/Y sky130_fd_sc_hd__nand2_4
X_52227_ _52198_/A _52248_/B sky130_fd_sc_hd__buf_2
X_71061_ _48922_/B _71047_/X _71060_/Y _83621_/D sky130_fd_sc_hd__o21ai_4
X_83047_ _83049_/CLK _74524_/Y _83047_/Q sky130_fd_sc_hd__dfxtp_4
X_87924_ _88180_/CLK _42317_/X _87924_/Q sky130_fd_sc_hd__dfxtp_4
X_80259_ _80259_/A _80259_/B _80261_/A sky130_fd_sc_hd__nand2_4
X_70012_ _70012_/A _70012_/X sky130_fd_sc_hd__buf_2
X_59823_ _59664_/A _59823_/X sky130_fd_sc_hd__buf_2
X_52158_ _52168_/A _52158_/B _52158_/Y sky130_fd_sc_hd__nand2_4
X_87855_ _88345_/CLK _87855_/D _87855_/Q sky130_fd_sc_hd__dfxtp_4
X_51109_ _51191_/A _51115_/A sky130_fd_sc_hd__buf_2
X_74820_ _74831_/A _74829_/A sky130_fd_sc_hd__buf_2
X_86806_ _87888_/CLK _46027_/X _66544_/B sky130_fd_sc_hd__dfxtp_4
X_59754_ _59754_/A _59731_/Y _59754_/C _59754_/D _59754_/X sky130_fd_sc_hd__and4_4
X_52089_ _52152_/A _52089_/X sky130_fd_sc_hd__buf_2
X_44980_ _85244_/Q _44979_/X _44926_/X _44980_/X sky130_fd_sc_hd__o21a_4
X_56966_ _57019_/A _56966_/X sky130_fd_sc_hd__buf_2
X_87786_ _87789_/CLK _42654_/X _87786_/Q sky130_fd_sc_hd__dfxtp_4
X_84998_ _84998_/CLK _84998_/D _57468_/A sky130_fd_sc_hd__dfxtp_4
X_58705_ _58703_/X _85462_/Q _58704_/X _58705_/Y sky130_fd_sc_hd__o21ai_4
X_43931_ _43916_/X _43924_/X _41424_/X _67939_/B _43917_/X _43932_/A
+ sky130_fd_sc_hd__o32ai_4
X_74751_ _74751_/A _74804_/A _74797_/C _71738_/X _74751_/Y sky130_fd_sc_hd__nand4_4
X_55917_ _55907_/X _55912_/X _55914_/X _55916_/X _55918_/A sky130_fd_sc_hd__and4_4
X_86737_ _85815_/CLK _46440_/Y _86737_/Q sky130_fd_sc_hd__dfxtp_4
X_71963_ _83312_/Q _57615_/X _71962_/Y _71963_/Y sky130_fd_sc_hd__o21ai_4
X_83949_ _80776_/CLK _83949_/D _83949_/Q sky130_fd_sc_hd__dfxtp_4
X_59685_ _59684_/X _59699_/A sky130_fd_sc_hd__buf_2
X_56897_ _56892_/Y _56897_/B _85125_/D sky130_fd_sc_hd__nand2_4
X_73702_ _43041_/Y _73627_/X _73652_/X _73701_/Y _73702_/X sky130_fd_sc_hd__a211o_4
X_46650_ _46650_/A _51770_/B sky130_fd_sc_hd__buf_2
X_70914_ _70860_/A _70914_/B _70914_/C _70914_/D _70914_/Y sky130_fd_sc_hd__nand4_4
X_58636_ _58868_/A _58636_/X sky130_fd_sc_hd__buf_2
X_77470_ _77471_/A _77471_/B _77475_/A sky130_fd_sc_hd__nor2_4
X_43862_ _43810_/A _43862_/X sky130_fd_sc_hd__buf_2
X_55848_ _44079_/X _55848_/B _55848_/X sky130_fd_sc_hd__and2_4
X_74682_ _74679_/A _45761_/A _74682_/Y sky130_fd_sc_hd__nand2_4
X_86668_ _86351_/CLK _47122_/Y _86668_/Q sky130_fd_sc_hd__dfxtp_4
X_71894_ _70530_/Y _71894_/Y sky130_fd_sc_hd__inv_2
X_45601_ _45599_/Y _45570_/X _45520_/X _45600_/Y _45601_/X sky130_fd_sc_hd__a211o_4
X_76421_ _76404_/X _76400_/X _76401_/X _76421_/Y sky130_fd_sc_hd__a21oi_4
X_42813_ _41429_/X _42802_/X _87705_/Q _42803_/X _87705_/D sky130_fd_sc_hd__a2bb2o_4
X_73633_ _74244_/B _73633_/X sky130_fd_sc_hd__buf_2
X_85619_ _86549_/CLK _53530_/Y _85619_/Q sky130_fd_sc_hd__dfxtp_4
X_70845_ _51770_/B _70831_/X _70844_/Y _70845_/Y sky130_fd_sc_hd__o21ai_4
X_58567_ _58079_/X _58564_/Y _58566_/Y _58098_/X _58083_/X _58567_/X
+ sky130_fd_sc_hd__o32a_4
X_46581_ _46578_/X _49179_/A _46580_/X _51384_/B sky130_fd_sc_hd__o21ai_4
X_43793_ _43792_/Y _87265_/D sky130_fd_sc_hd__inv_2
X_55779_ _55761_/A _85290_/Q _55779_/X sky130_fd_sc_hd__and2_4
X_86599_ _85961_/CLK _86599_/D _72428_/A sky130_fd_sc_hd__dfxtp_4
X_48320_ _74177_/B _48293_/X _48319_/Y _48320_/Y sky130_fd_sc_hd__o21ai_4
X_79140_ _79140_/A _61546_/C _79140_/X sky130_fd_sc_hd__xor2_4
X_45532_ _45524_/X _45528_/Y _45531_/Y _45532_/Y sky130_fd_sc_hd__a21oi_4
X_57518_ _57499_/A _73717_/A _57518_/Y sky130_fd_sc_hd__nand2_4
X_88338_ _88337_/CLK _40772_/X _88338_/Q sky130_fd_sc_hd__dfxtp_4
X_76352_ _76348_/X _76349_/Y _76353_/B _76352_/X sky130_fd_sc_hd__a21o_4
X_42744_ _51949_/A _42745_/A sky130_fd_sc_hd__buf_2
X_73564_ _73449_/X _85633_/Q _73450_/X _73563_/X _73564_/X sky130_fd_sc_hd__a211o_4
X_70776_ _52850_/B _70761_/X _70775_/Y _70776_/Y sky130_fd_sc_hd__o21ai_4
X_58498_ _58498_/A _58498_/B _58498_/Y sky130_fd_sc_hd__nand2_4
X_75303_ _75294_/Y _75303_/B _75304_/A sky130_fd_sc_hd__and2_4
X_48251_ _47975_/B _50300_/B sky130_fd_sc_hd__buf_2
X_72515_ _72563_/B _72508_/A _72607_/C _72515_/D _72517_/A sky130_fd_sc_hd__nand4_4
X_79071_ _79071_/A _79071_/B _79071_/X sky130_fd_sc_hd__xor2_4
X_45463_ _83005_/Q _44894_/B _45463_/Y sky130_fd_sc_hd__nor2_4
X_57449_ _57441_/X _56821_/X _57448_/X _57449_/X sky130_fd_sc_hd__o21a_4
X_76283_ _76283_/A _76283_/Y sky130_fd_sc_hd__inv_2
X_88269_ _88272_/CLK _88269_/D _88269_/Q sky130_fd_sc_hd__dfxtp_4
X_42675_ _42674_/Y _87776_/D sky130_fd_sc_hd__inv_2
X_73495_ _73495_/A _85860_/Q _73495_/X sky130_fd_sc_hd__and2_4
X_47202_ _47210_/A _47181_/B _47210_/C _51220_/D _47202_/X sky130_fd_sc_hd__and4_4
X_78022_ _78022_/A _78022_/Y sky130_fd_sc_hd__inv_2
X_44414_ _41529_/X _44412_/X _87121_/Q _44413_/X _44414_/X sky130_fd_sc_hd__a2bb2o_4
X_75234_ _75216_/Y _75219_/Y _75233_/X _75234_/Y sky130_fd_sc_hd__o21ai_4
X_41626_ _41625_/Y _41626_/X sky130_fd_sc_hd__buf_2
X_60460_ _60460_/A _60571_/B sky130_fd_sc_hd__buf_2
X_72446_ _72414_/X _86277_/Q _72446_/Y sky130_fd_sc_hd__nor2_4
X_48182_ _65939_/B _48170_/X _48181_/Y _48182_/Y sky130_fd_sc_hd__o21ai_4
X_45394_ _44891_/X _45394_/X sky130_fd_sc_hd__buf_2
X_47133_ _47113_/A _47133_/B _47091_/X _52872_/D _47133_/X sky130_fd_sc_hd__and4_4
X_59119_ _58923_/A _59119_/X sky130_fd_sc_hd__buf_2
X_44345_ _40409_/X _44345_/X sky130_fd_sc_hd__buf_2
X_75165_ _75131_/Y _75145_/Y _75144_/Y _75165_/X sky130_fd_sc_hd__a21o_4
X_41557_ _41556_/X _41530_/X _67011_/B _41531_/X _88193_/D sky130_fd_sc_hd__a2bb2o_4
X_60391_ _61183_/A _59905_/B _60512_/A sky130_fd_sc_hd__nor2_4
X_72377_ _72461_/A _72377_/B _72377_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_opt_3_CLK _83246_/CLK _84840_/CLK sky130_fd_sc_hd__clkbuf_16
X_62130_ _62129_/X _61748_/X _59608_/A _62130_/D _62131_/D sky130_fd_sc_hd__nand4_4
X_74116_ _74102_/Y _74116_/B _74116_/Y sky130_fd_sc_hd__xnor2_4
X_40508_ _40409_/X _40508_/X sky130_fd_sc_hd__buf_2
X_47064_ _59189_/A _47050_/X _47063_/Y _47064_/Y sky130_fd_sc_hd__o21ai_4
X_71328_ _50365_/B _71320_/X _71327_/Y _83535_/D sky130_fd_sc_hd__o21ai_4
X_44276_ _57327_/B _57331_/B sky130_fd_sc_hd__buf_2
X_79973_ _79973_/A _79971_/X _79972_/Y _79973_/Y sky130_fd_sc_hd__nand3_4
X_75096_ _75096_/A _75098_/A sky130_fd_sc_hd__inv_2
X_41488_ _41485_/X _41486_/X _66694_/B _41487_/X _88206_/D sky130_fd_sc_hd__a2bb2o_4
X_46015_ _46013_/X _46001_/X _40514_/X _86814_/Q _46014_/X _46016_/A
+ sky130_fd_sc_hd__o32ai_4
X_43227_ _43226_/X _43207_/X _40994_/X _87528_/Q _43212_/X _43227_/Y
+ sky130_fd_sc_hd__o32ai_4
X_62061_ _84892_/Q _62128_/B _62010_/X _62060_/X _62061_/Y sky130_fd_sc_hd__nand4_4
X_78924_ _78912_/A _78912_/B _78924_/Y sky130_fd_sc_hd__nor2_4
X_74047_ _74048_/B _74048_/C _74046_/X _74047_/X sky130_fd_sc_hd__a21o_4
X_40439_ _40421_/X _81173_/Q _40438_/X _40439_/X sky130_fd_sc_hd__o21a_4
X_71259_ _50264_/B _71239_/A _71258_/Y _83555_/D sky130_fd_sc_hd__o21ai_4
X_61012_ _61012_/A _60918_/X _61012_/C _61012_/Y sky130_fd_sc_hd__nand3_4
X_43158_ _43158_/A _43158_/Y sky130_fd_sc_hd__inv_2
X_78855_ _78857_/B _78857_/A _78855_/X sky130_fd_sc_hd__or2_4
X_42109_ _42109_/A _42109_/Y sky130_fd_sc_hd__inv_2
X_65820_ _65685_/X _86183_/Q _65701_/X _65819_/X _65820_/X sky130_fd_sc_hd__a211o_4
X_77806_ _82059_/Q _77806_/Y sky130_fd_sc_hd__inv_2
X_47966_ _47962_/Y _47954_/X _47965_/X _47966_/Y sky130_fd_sc_hd__a21oi_4
X_43089_ _87580_/Q _43089_/Y sky130_fd_sc_hd__inv_2
X_78786_ _78752_/A _78758_/A _78778_/B _78786_/X sky130_fd_sc_hd__a21o_4
X_75998_ _81333_/Q _81421_/Q _76005_/C sky130_fd_sc_hd__nand2_4
X_49705_ _49569_/A _49787_/A sky130_fd_sc_hd__buf_2
X_46917_ _46916_/Y _52746_/D sky130_fd_sc_hd__buf_2
X_65751_ _65733_/X _85580_/Q _65734_/X _65750_/X _65751_/X sky130_fd_sc_hd__a211o_4
X_77737_ _77736_/Y _77737_/B _78045_/B sky130_fd_sc_hd__nand2_4
X_62963_ _62971_/A _64525_/C _60302_/X _62979_/D _62963_/X sky130_fd_sc_hd__and4_4
X_74949_ _80944_/Q _74949_/B _74949_/X sky130_fd_sc_hd__xor2_4
X_47897_ _47840_/A _47897_/X sky130_fd_sc_hd__buf_2
X_64702_ _64695_/X _64700_/X _64701_/X _64702_/X sky130_fd_sc_hd__a21o_4
X_49636_ _49625_/A _49614_/X _49629_/X _52853_/D _49636_/X sky130_fd_sc_hd__and4_4
X_61914_ _61912_/Y _61881_/X _61913_/Y _61914_/Y sky130_fd_sc_hd__a21oi_4
X_68470_ _69678_/A _68470_/X sky130_fd_sc_hd__buf_2
X_46848_ _46830_/A _46845_/X _46830_/C _52709_/D _46848_/X sky130_fd_sc_hd__and4_4
X_65682_ _65682_/A _65683_/C sky130_fd_sc_hd__inv_2
X_77668_ _77667_/X _77668_/Y sky130_fd_sc_hd__inv_2
X_62894_ _62894_/A _62852_/X _84373_/Q _62894_/Y sky130_fd_sc_hd__nor3_4
X_67421_ _67517_/A _67421_/B _67421_/X sky130_fd_sc_hd__and2_4
X_79407_ _79419_/A _79419_/B _79418_/A sky130_fd_sc_hd__xor2_4
X_64633_ _64630_/X _64633_/B _64632_/X _64633_/Y sky130_fd_sc_hd__nand3_4
X_76619_ _81664_/Q _76619_/Y sky130_fd_sc_hd__inv_2
X_61845_ _61856_/A _61846_/B sky130_fd_sc_hd__buf_2
X_49567_ _49558_/A _52781_/B _49567_/Y sky130_fd_sc_hd__nand2_4
X_46779_ _52667_/B _50976_/B sky130_fd_sc_hd__buf_2
X_77599_ _77599_/A _77603_/A sky130_fd_sc_hd__inv_2
X_48518_ _81779_/Q _48520_/A sky130_fd_sc_hd__inv_2
X_67352_ _67166_/X _67340_/Y _67269_/X _67351_/Y _67352_/X sky130_fd_sc_hd__a211o_4
X_79338_ _79316_/Y _79334_/X _79337_/Y _79339_/B sky130_fd_sc_hd__a21oi_4
X_64564_ _64696_/A _64564_/X sky130_fd_sc_hd__buf_2
X_49498_ _49502_/A _51022_/B _49498_/Y sky130_fd_sc_hd__nand2_4
X_61776_ _61365_/X _61794_/B _59810_/A _61776_/D _61776_/Y sky130_fd_sc_hd__nand4_4
X_66303_ _66300_/X _66303_/B _66303_/Y sky130_fd_sc_hd__nand2_4
X_63515_ _63495_/X _63509_/X _63510_/X _63513_/X _63514_/Y _63515_/Y
+ sky130_fd_sc_hd__o41ai_4
X_48449_ _48449_/A _48449_/B _48449_/Y sky130_fd_sc_hd__nand2_4
X_60727_ _60727_/A _60723_/X _60726_/Y _60727_/Y sky130_fd_sc_hd__nand3_4
X_67283_ _80900_/D _67211_/X _67282_/X _84076_/D sky130_fd_sc_hd__a21bo_4
X_79269_ _79282_/A _79268_/Y _79292_/B sky130_fd_sc_hd__xor2_4
X_64495_ _64474_/A _64421_/X _84888_/Q _64495_/X sky130_fd_sc_hd__and3_4
X_81300_ _81259_/CLK _76988_/X _81300_/Q sky130_fd_sc_hd__dfxtp_4
X_69022_ _43098_/A _68975_/X _66349_/X _69021_/X _69022_/X sky130_fd_sc_hd__a211o_4
X_66234_ _66181_/A _74104_/B _66234_/X sky130_fd_sc_hd__and2_4
X_51460_ _51481_/A _52986_/B _51460_/Y sky130_fd_sc_hd__nand2_4
X_63446_ _63456_/A _63456_/B _80559_/B _63446_/Y sky130_fd_sc_hd__nor3_4
X_82280_ _82288_/CLK _82280_/D _82280_/Q sky130_fd_sc_hd__dfxtp_4
X_60658_ _63540_/A _60697_/B sky130_fd_sc_hd__buf_2
X_50411_ _86206_/Q _50403_/X _50410_/Y _50411_/Y sky130_fd_sc_hd__o21ai_4
X_81231_ _81233_/CLK _81039_/Q _81231_/Q sky130_fd_sc_hd__dfxtp_4
X_66165_ _66162_/Y _66137_/X _66164_/Y _66165_/X sky130_fd_sc_hd__a21o_4
X_51391_ _51793_/A _51391_/X sky130_fd_sc_hd__buf_2
X_63377_ _61329_/B _60834_/X _63374_/X _63376_/X _63377_/X sky130_fd_sc_hd__a211o_4
X_60589_ _60440_/X _60439_/X _60588_/X _63272_/A sky130_fd_sc_hd__a21oi_4
Xclkbuf_7_104_0_CLK clkbuf_6_52_0_CLK/X clkbuf_8_209_0_CLK/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_292_0_CLK clkbuf_9_146_0_CLK/X _84732_/CLK sky130_fd_sc_hd__clkbuf_1
X_53130_ _53128_/Y _53111_/X _53129_/X _85692_/D sky130_fd_sc_hd__a21oi_4
X_65116_ _64944_/X _86125_/Q _65022_/X _65115_/X _65116_/X sky130_fd_sc_hd__a211o_4
X_50342_ _86220_/Q _50316_/X _50341_/Y _50342_/Y sky130_fd_sc_hd__o21ai_4
X_62328_ _62267_/A _62267_/B _62328_/C _62328_/Y sky130_fd_sc_hd__nor3_4
X_81162_ _80835_/CLK _74906_/B _81162_/Q sky130_fd_sc_hd__dfxtp_4
X_66096_ _65976_/A _66096_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_74_0_CLK clkbuf_9_37_0_CLK/X _83012_/CLK sky130_fd_sc_hd__clkbuf_1
X_80113_ _80109_/X _80112_/Y _80114_/A sky130_fd_sc_hd__xor2_4
X_53061_ _85704_/Q _53038_/X _53060_/Y _53061_/Y sky130_fd_sc_hd__o21ai_4
X_65047_ _65047_/A _65047_/B _65047_/C _65047_/Y sky130_fd_sc_hd__nor3_4
X_69924_ _87044_/Q _69690_/X _68473_/X _69923_/X _69924_/X sky130_fd_sc_hd__a211o_4
X_50273_ _86233_/Q _50250_/X _50272_/Y _50273_/Y sky130_fd_sc_hd__o21ai_4
X_62259_ _59976_/A _62259_/X sky130_fd_sc_hd__buf_2
X_85970_ _85679_/CLK _51659_/Y _85970_/Q sky130_fd_sc_hd__dfxtp_4
X_81093_ _81928_/CLK _81093_/D _81093_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_220_0_CLK clkbuf_8_221_0_CLK/A clkbuf_9_441_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_52012_ _52010_/Y _51987_/X _52011_/X _52012_/Y sky130_fd_sc_hd__a21oi_4
X_80044_ _80030_/Y _80035_/Y _80043_/X _80045_/B sky130_fd_sc_hd__o21ai_4
X_84921_ _84921_/CLK _58148_/Y _61323_/A sky130_fd_sc_hd__dfxtp_4
X_69855_ _69852_/X _69855_/B _69855_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_7_119_0_CLK clkbuf_6_59_0_CLK/X clkbuf_8_239_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_56820_ _56820_/A _56725_/B _56820_/Y sky130_fd_sc_hd__nand2_4
X_68806_ _69035_/A _68806_/X sky130_fd_sc_hd__buf_2
X_87640_ _86920_/CLK _42941_/Y _67985_/B sky130_fd_sc_hd__dfxtp_4
X_84852_ _84732_/CLK _84852_/D _84852_/Q sky130_fd_sc_hd__dfxtp_4
X_69786_ _69360_/X _69363_/X _69728_/X _69786_/Y sky130_fd_sc_hd__a21oi_4
X_66998_ _66879_/A _66998_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_89_0_CLK clkbuf_9_44_0_CLK/X _84409_/CLK sky130_fd_sc_hd__clkbuf_1
X_83803_ _81807_/CLK _70307_/X _74748_/A sky130_fd_sc_hd__dfxtp_4
X_56751_ _57427_/A _56750_/Y _56752_/A sky130_fd_sc_hd__nand2_4
X_68737_ _68737_/A _68737_/X sky130_fd_sc_hd__buf_2
X_87571_ _83153_/CLK _43114_/Y _87571_/Q sky130_fd_sc_hd__dfxtp_4
X_53963_ _53874_/A _53964_/B sky130_fd_sc_hd__buf_2
X_65949_ _65946_/X _65948_/X _65937_/X _65949_/X sky130_fd_sc_hd__a21o_4
X_84783_ _84906_/CLK _58977_/X _62948_/C sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_235_0_CLK clkbuf_8_235_0_CLK/A clkbuf_9_471_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_81995_ _82131_/CLK _82027_/Q _77069_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_230_0_CLK clkbuf_9_115_0_CLK/X _82211_/CLK sky130_fd_sc_hd__clkbuf_1
X_55702_ _55711_/A _55702_/B _55702_/X sky130_fd_sc_hd__and2_4
X_86522_ _85593_/CLK _48443_/Y _86522_/Q sky130_fd_sc_hd__dfxtp_4
X_52914_ _52910_/A _51222_/B _52914_/Y sky130_fd_sc_hd__nand2_4
X_59470_ _84723_/Q _59471_/A sky130_fd_sc_hd__inv_2
X_83734_ _86317_/CLK _83734_/D _83734_/Q sky130_fd_sc_hd__dfxtp_4
X_56682_ _56682_/A _56682_/X sky130_fd_sc_hd__buf_2
X_80946_ _80813_/CLK _80990_/Q _80946_/Q sky130_fd_sc_hd__dfxtp_4
X_68668_ _68668_/A _68669_/B sky130_fd_sc_hd__inv_2
Xclkbuf_10_860_0_CLK clkbuf_9_430_0_CLK/X _86127_/CLK sky130_fd_sc_hd__clkbuf_1
X_53894_ _53891_/Y _53892_/X _53893_/X _53894_/Y sky130_fd_sc_hd__a21oi_4
X_58421_ _58421_/A _58415_/B _58421_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_12_0_CLK clkbuf_9_6_0_CLK/X _85248_/CLK sky130_fd_sc_hd__clkbuf_1
X_67619_ _68442_/A _67619_/X sky130_fd_sc_hd__buf_2
X_55633_ _55630_/X _55632_/X _55634_/A sky130_fd_sc_hd__and2_4
X_86453_ _86453_/CLK _86453_/D _86453_/Q sky130_fd_sc_hd__dfxtp_4
X_52845_ _52845_/A _52853_/C sky130_fd_sc_hd__buf_2
X_83665_ _83666_/CLK _70915_/Y _46840_/A sky130_fd_sc_hd__dfxtp_4
X_80877_ _80849_/CLK _75675_/B _80877_/Q sky130_fd_sc_hd__dfxtp_4
X_68599_ _68599_/A _87754_/Q _68599_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_351_0_CLK clkbuf_9_351_0_CLK/A clkbuf_9_351_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_85404_ _85404_/CLK _54646_/Y _85404_/Q sky130_fd_sc_hd__dfxtp_4
X_70630_ _71735_/A _70630_/B _71115_/D _71735_/C _70630_/X sky130_fd_sc_hd__and4_4
X_58352_ _58352_/A _58344_/B _58352_/Y sky130_fd_sc_hd__nor2_4
X_82616_ _82503_/CLK _79011_/B _82616_/Q sky130_fd_sc_hd__dfxtp_4
X_55564_ _55836_/A _55843_/A sky130_fd_sc_hd__buf_2
X_86384_ _86384_/CLK _86384_/D _86384_/Q sky130_fd_sc_hd__dfxtp_4
X_40790_ _40817_/A _40790_/B _40790_/X sky130_fd_sc_hd__or2_4
X_52776_ _52774_/Y _52755_/X _52775_/X _52776_/Y sky130_fd_sc_hd__a21oi_4
X_83596_ _86149_/CLK _83596_/D _49175_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_245_0_CLK clkbuf_9_122_0_CLK/X _84590_/CLK sky130_fd_sc_hd__clkbuf_1
X_57303_ _57268_/X _56783_/X _56785_/D _57303_/Y sky130_fd_sc_hd__nand3_4
X_88123_ _87417_/CLK _41851_/Y _88123_/Q sky130_fd_sc_hd__dfxtp_4
X_54515_ _85428_/Q _54512_/X _54514_/Y _54515_/Y sky130_fd_sc_hd__o21ai_4
X_85335_ _85335_/CLK _55014_/Y _85335_/Q sky130_fd_sc_hd__dfxtp_4
X_51727_ _51725_/Y _51719_/X _51726_/X _85957_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_875_0_CLK clkbuf_9_437_0_CLK/X _86237_/CLK sky130_fd_sc_hd__clkbuf_1
X_70561_ DATA_TO_HASH[2] _71570_/A sky130_fd_sc_hd__inv_2
X_58283_ _58283_/A _58283_/Y sky130_fd_sc_hd__inv_2
X_82547_ _82541_/CLK _82547_/D _82547_/Q sky130_fd_sc_hd__dfxtp_4
X_55495_ _44061_/X _45584_/Y _55495_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_27_0_CLK clkbuf_9_13_0_CLK/X _82993_/CLK sky130_fd_sc_hd__clkbuf_1
X_72300_ _59255_/A _72347_/A sky130_fd_sc_hd__buf_2
X_57234_ _57326_/C _57322_/B sky130_fd_sc_hd__buf_2
X_88054_ _87542_/CLK _88054_/D _42057_/A sky130_fd_sc_hd__dfxtp_4
X_42460_ _41841_/X _42460_/X sky130_fd_sc_hd__buf_2
X_54446_ _54446_/A _54446_/B _54446_/Y sky130_fd_sc_hd__nand2_4
X_73280_ _69842_/B _73279_/X _73202_/X _73280_/X sky130_fd_sc_hd__o21a_4
X_85266_ _85167_/CLK _56234_/Y _56233_/C sky130_fd_sc_hd__dfxtp_4
X_51658_ _51657_/X _51651_/B _51651_/C _53181_/D _51658_/X sky130_fd_sc_hd__and4_4
Xclkbuf_9_366_0_CLK clkbuf_9_367_0_CLK/A clkbuf_9_366_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_70492_ _70491_/Y _71136_/A sky130_fd_sc_hd__buf_2
X_82478_ _82563_/CLK _78483_/X _78102_/B sky130_fd_sc_hd__dfxtp_4
X_41411_ _47867_/A _41411_/X sky130_fd_sc_hd__buf_2
X_87005_ _86984_/CLK _44674_/Y _87005_/Q sky130_fd_sc_hd__dfxtp_4
X_72231_ _72227_/Y _72230_/Y _72185_/X _72231_/X sky130_fd_sc_hd__a21o_4
X_84217_ _81227_/CLK _65048_/X _84217_/Q sky130_fd_sc_hd__dfxtp_4
X_50609_ _50551_/A _50609_/X sky130_fd_sc_hd__buf_2
X_57165_ _57010_/Y _57163_/Y _57164_/X _57126_/A _57165_/X sky130_fd_sc_hd__a211o_4
X_81429_ _84049_/CLK _81461_/Q _76056_/B sky130_fd_sc_hd__dfxtp_4
X_54377_ _54322_/A _54378_/A sky130_fd_sc_hd__buf_2
X_42391_ _42378_/X _42369_/X _40395_/X _87886_/Q _42370_/X _42392_/A
+ sky130_fd_sc_hd__o32ai_4
X_85197_ _85257_/CLK _56430_/Y _85197_/Q sky130_fd_sc_hd__dfxtp_4
X_51589_ _51583_/Y _51585_/X _51588_/X _85983_/D sky130_fd_sc_hd__a21oi_4
X_44130_ _73284_/A _44130_/X sky130_fd_sc_hd__buf_2
X_56116_ _56112_/X _56114_/X _56115_/Y _85293_/D sky130_fd_sc_hd__o21ai_4
X_53328_ _53355_/A _53328_/X sky130_fd_sc_hd__buf_2
X_41342_ _41337_/X _41338_/X _41341_/X _88233_/Q _41333_/X _41343_/A
+ sky130_fd_sc_hd__o32ai_4
X_72162_ _72162_/A _72162_/B _72162_/Y sky130_fd_sc_hd__nor2_4
X_84148_ _82746_/CLK _66219_/X _84148_/Q sky130_fd_sc_hd__dfxtp_4
X_57096_ _44236_/X _57096_/Y sky130_fd_sc_hd__inv_2
X_71113_ _71112_/X _71091_/B _70890_/D _71113_/Y sky130_fd_sc_hd__nand3_4
X_44061_ _44060_/X _44061_/X sky130_fd_sc_hd__buf_2
X_56047_ _74306_/C _56047_/Y sky130_fd_sc_hd__inv_2
X_41273_ _41272_/X _41251_/X _88246_/Q _41253_/X _41273_/X sky130_fd_sc_hd__a2bb2o_4
X_53259_ _53259_/A _53259_/B _53259_/Y sky130_fd_sc_hd__nand2_4
X_72093_ _83286_/Q _72090_/X _72092_/Y _72093_/Y sky130_fd_sc_hd__o21ai_4
X_76970_ _84522_/Q _62636_/C _76970_/X sky130_fd_sc_hd__xor2_4
X_84079_ _84079_/CLK _67210_/X _80903_/D sky130_fd_sc_hd__dfxtp_4
X_43012_ _41863_/A _43012_/B _43175_/C sky130_fd_sc_hd__nor2_4
X_71044_ _53179_/B _71013_/A _71043_/Y _71044_/Y sky130_fd_sc_hd__o21ai_4
X_75921_ _61132_/C _84391_/Q _80735_/D sky130_fd_sc_hd__xor2_4
X_87907_ _87394_/CLK _87907_/D _87907_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_813_0_CLK clkbuf_9_406_0_CLK/X _82855_/CLK sky130_fd_sc_hd__clkbuf_1
X_47820_ _72476_/A _47806_/X _47819_/Y _47820_/Y sky130_fd_sc_hd__o21ai_4
X_59806_ _59806_/A _59721_/A _59722_/A _59807_/A sky130_fd_sc_hd__and3_4
X_78640_ _78640_/A _78640_/B _78640_/C _78621_/Y _78640_/X sky130_fd_sc_hd__and4_4
X_75852_ _75852_/A _75867_/A _75860_/A sky130_fd_sc_hd__xnor2_4
X_87838_ _87850_/CLK _42514_/Y _87838_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_304_0_CLK clkbuf_8_152_0_CLK/X clkbuf_9_304_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_57998_ _57997_/X _85485_/Q _57923_/X _57998_/X sky130_fd_sc_hd__o21a_4
X_74803_ _74741_/X _74798_/X _74802_/Y _74803_/Y sky130_fd_sc_hd__nand3_4
X_47751_ _47751_/A _47752_/A sky130_fd_sc_hd__inv_2
X_59737_ _59737_/A _59711_/B _80548_/A _59737_/Y sky130_fd_sc_hd__nor3_4
X_78571_ _78552_/Y _78554_/A _78551_/A _78572_/A sky130_fd_sc_hd__o21a_4
X_44963_ _44895_/X _44963_/X sky130_fd_sc_hd__buf_2
X_56949_ _44213_/X _56949_/X sky130_fd_sc_hd__buf_2
X_75783_ _80920_/Q _75781_/Y _75782_/Y _75783_/Y sky130_fd_sc_hd__a21oi_4
X_87769_ _87520_/CLK _87769_/D _87769_/Q sky130_fd_sc_hd__dfxtp_4
X_72995_ _72995_/A _72994_/X _72996_/B sky130_fd_sc_hd__nand2_4
X_46702_ _46712_/A _46701_/X _46702_/Y sky130_fd_sc_hd__nand2_4
X_77522_ _77521_/Y _77522_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_828_0_CLK clkbuf_9_414_0_CLK/X _82925_/CLK sky130_fd_sc_hd__clkbuf_1
X_43914_ _43895_/X _43902_/X _41382_/X _87201_/Q _43897_/X _43914_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74734_ _70669_/A _74734_/Y sky130_fd_sc_hd__inv_2
X_47682_ _81233_/Q _47682_/Y sky130_fd_sc_hd__inv_2
X_71946_ _55671_/Y _71939_/X _71945_/Y _83319_/D sky130_fd_sc_hd__o21ai_4
X_59668_ _59588_/Y _59668_/B _59763_/A sky130_fd_sc_hd__nand2_4
X_44894_ _74541_/C _44894_/B _44894_/Y sky130_fd_sc_hd__nor2_4
X_49421_ _49419_/Y _49405_/X _49420_/X _86391_/D sky130_fd_sc_hd__a21oi_4
X_46633_ _83687_/Q _54277_/B sky130_fd_sc_hd__inv_2
X_58619_ _58571_/X _85789_/Q _58594_/X _58619_/X sky130_fd_sc_hd__o21a_4
X_77453_ _77453_/A _82193_/D _77453_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_9_319_0_CLK clkbuf_9_318_0_CLK/A clkbuf_9_319_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_43845_ _41189_/X _43842_/X _68718_/B _43843_/X _87237_/D sky130_fd_sc_hd__a2bb2o_4
X_74665_ _74694_/A _74673_/A sky130_fd_sc_hd__buf_2
X_71877_ _71871_/X _83344_/Q _71876_/Y _71877_/X sky130_fd_sc_hd__a21o_4
X_59599_ _60630_/A _60630_/C _60636_/B sky130_fd_sc_hd__and2_4
X_76404_ _76368_/A _76369_/X _76379_/X _76404_/X sky130_fd_sc_hd__a21o_4
X_49352_ _49352_/A _51389_/B _49352_/Y sky130_fd_sc_hd__nand2_4
X_61630_ _61630_/A _61611_/B _61611_/C _61572_/D _61630_/Y sky130_fd_sc_hd__nand4_4
X_73616_ _73641_/A _65939_/B _73616_/X sky130_fd_sc_hd__and2_4
X_46564_ _54077_/B _51378_/B sky130_fd_sc_hd__buf_2
X_70828_ _70828_/A _70832_/A sky130_fd_sc_hd__buf_2
X_77384_ _77382_/X _77383_/Y _77385_/A sky130_fd_sc_hd__and2_4
X_43776_ _43776_/A _43776_/X sky130_fd_sc_hd__buf_2
X_74596_ _74591_/X _74583_/X _56114_/A _74584_/X _74596_/X sky130_fd_sc_hd__a211o_4
X_40988_ _40755_/A _40989_/A sky130_fd_sc_hd__buf_2
X_48303_ _52050_/A _48286_/X _48287_/C _48303_/X sky130_fd_sc_hd__and3_4
X_79123_ _82836_/Q _79123_/B _79123_/Y sky130_fd_sc_hd__xnor2_4
X_45515_ _57113_/B _45515_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_5_4_0_CLK clkbuf_4_2_1_CLK/X clkbuf_6_9_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_76335_ _76331_/Y _76333_/Y _76330_/Y _76336_/B sky130_fd_sc_hd__o21ai_4
X_42727_ _41189_/X _42717_/X _87749_/Q _42718_/X _87749_/D sky130_fd_sc_hd__a2bb2o_4
X_49283_ _50802_/A _49283_/B _49234_/X _49283_/X sky130_fd_sc_hd__and3_4
X_73547_ _73544_/X _73545_/Y _73546_/X _73547_/Y sky130_fd_sc_hd__a21oi_4
X_61561_ _61561_/A _61542_/B _61542_/C _61512_/X _61561_/Y sky130_fd_sc_hd__nand4_4
X_70759_ _70764_/A _70760_/B sky130_fd_sc_hd__inv_2
X_46495_ _46505_/A _46495_/B _46495_/Y sky130_fd_sc_hd__nand2_4
X_63300_ _63272_/A _61640_/A _63280_/C _63300_/Y sky130_fd_sc_hd__nand3_4
X_48234_ _48234_/A _48201_/B _48195_/X _48234_/X sky130_fd_sc_hd__and3_4
X_60512_ _60512_/A _60512_/Y sky130_fd_sc_hd__inv_2
X_79054_ _79054_/A _79055_/B sky130_fd_sc_hd__inv_2
X_45446_ _45678_/A _45446_/X sky130_fd_sc_hd__buf_2
X_64280_ _64272_/Y _64279_/X _64269_/X _64280_/X sky130_fd_sc_hd__o21a_4
X_76266_ _76261_/X _76264_/Y _76262_/Y _76267_/B sky130_fd_sc_hd__nand3_4
X_42658_ _42580_/A _42658_/X sky130_fd_sc_hd__buf_2
X_61492_ _61492_/A _61468_/B _61467_/X _61451_/D _61492_/Y sky130_fd_sc_hd__nand4_4
X_73478_ _73478_/A _73477_/X _73478_/Y sky130_fd_sc_hd__nand2_4
X_78005_ _78003_/Y _78004_/Y _78007_/A sky130_fd_sc_hd__nand2_4
X_63231_ _63231_/A _63231_/X sky130_fd_sc_hd__buf_2
X_75217_ _75217_/A _75217_/B _75217_/Y sky130_fd_sc_hd__nor2_4
X_41609_ _41540_/X _41541_/X _41606_/X _88183_/Q _41608_/X _41610_/A
+ sky130_fd_sc_hd__o32ai_4
X_48165_ _48164_/A _57491_/C _48164_/Y _48165_/X sky130_fd_sc_hd__o21a_4
X_60443_ _60443_/A _60476_/D sky130_fd_sc_hd__buf_2
X_72429_ _72413_/X _72427_/Y _72428_/Y _57793_/X _72417_/X _72429_/X
+ sky130_fd_sc_hd__o32a_4
X_45377_ _45374_/Y _45376_/Y _45361_/X _45377_/X sky130_fd_sc_hd__a21o_4
X_76197_ _76195_/X _76196_/Y _76199_/B sky130_fd_sc_hd__nand2_4
X_42589_ _42465_/A _42590_/A sky130_fd_sc_hd__buf_2
X_47116_ _47116_/A _52863_/B sky130_fd_sc_hd__buf_2
X_44328_ _41651_/X _44326_/X _87163_/Q _44327_/X _87163_/D sky130_fd_sc_hd__a2bb2o_4
X_75148_ _75130_/Y _75135_/Y _75131_/Y _75148_/Y sky130_fd_sc_hd__o21ai_4
X_63162_ _63159_/Y _63161_/X _63114_/X _63162_/Y sky130_fd_sc_hd__a21oi_4
X_48096_ _48642_/B _48449_/B _48096_/Y sky130_fd_sc_hd__nand2_4
X_60374_ _60477_/A _60519_/B _60374_/C _60374_/Y sky130_fd_sc_hd__nor3_4
X_62113_ _84784_/Q _62113_/X sky130_fd_sc_hd__buf_2
X_47047_ _47047_/A _52827_/D sky130_fd_sc_hd__buf_2
X_44259_ _64850_/A _65880_/A sky130_fd_sc_hd__buf_2
X_67970_ _67948_/X _67961_/Y _67863_/X _67969_/Y _67970_/X sky130_fd_sc_hd__a211o_4
X_63093_ _63090_/Y _63092_/X _63056_/X _63093_/Y sky130_fd_sc_hd__a21oi_4
X_79956_ _79956_/A _79955_/Y _79958_/A sky130_fd_sc_hd__nand2_4
X_75079_ _75086_/A _75079_/B _75080_/B sky130_fd_sc_hd__xor2_4
X_66921_ _88389_/Q _66868_/X _66919_/X _66920_/X _66921_/X sky130_fd_sc_hd__a211o_4
X_62044_ _58264_/A _63610_/B sky130_fd_sc_hd__buf_2
X_78907_ _82636_/Q _82508_/D _78906_/Y _78907_/Y sky130_fd_sc_hd__a21oi_4
X_79887_ _79887_/A _79886_/Y _79888_/B sky130_fd_sc_hd__xor2_4
X_69640_ _69637_/X _69639_/X _69640_/Y sky130_fd_sc_hd__nand2_4
X_66852_ _66851_/X _66852_/B _66852_/X sky130_fd_sc_hd__and2_4
X_78838_ _78838_/A _78838_/B _78838_/X sky130_fd_sc_hd__xor2_4
X_48998_ _48998_/A _72014_/B sky130_fd_sc_hd__buf_2
X_65803_ _65800_/Y _65757_/X _65802_/Y _84177_/D sky130_fd_sc_hd__a21o_4
X_69571_ _69566_/X _69569_/X _69570_/X _69571_/X sky130_fd_sc_hd__a21o_4
X_47949_ _47841_/A _47988_/A sky130_fd_sc_hd__buf_2
X_66783_ _87946_/Q _66759_/X _66688_/X _66782_/X _66783_/X sky130_fd_sc_hd__a211o_4
X_78769_ _78769_/A _78769_/B _78769_/Y sky130_fd_sc_hd__nor2_4
X_63995_ _63960_/A _63960_/B _63995_/C _63995_/Y sky130_fd_sc_hd__nor3_4
X_80800_ _80821_/CLK _75867_/Y _80800_/Q sky130_fd_sc_hd__dfxtp_4
X_68522_ _68519_/X _68521_/X _68442_/X _68525_/A sky130_fd_sc_hd__a21o_4
X_65734_ _64829_/A _65734_/X sky130_fd_sc_hd__buf_2
X_50960_ _50956_/Y _50957_/X _50959_/X _86100_/D sky130_fd_sc_hd__a21oi_4
X_81780_ _81703_/CLK _76104_/X _81780_/Q sky130_fd_sc_hd__dfxtp_4
X_62946_ _62644_/X _58194_/A _60253_/A _60220_/A _62946_/X sky130_fd_sc_hd__and4_4
X_49619_ _49610_/A _49614_/X _49615_/C _52835_/D _49619_/X sky130_fd_sc_hd__and4_4
Xclkbuf_7_81_0_CLK clkbuf_7_81_0_CLK/A clkbuf_7_81_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_68453_ _87504_/Q _68365_/X _68450_/X _68452_/X _68453_/X sky130_fd_sc_hd__a211o_4
X_80731_ _81048_/CLK _75917_/X _80699_/D sky130_fd_sc_hd__dfxtp_4
X_65665_ _65621_/A _65559_/B _84186_/Q _65665_/X sky130_fd_sc_hd__and3_4
X_50891_ _50908_/A _50045_/X _50886_/C _51756_/D _50891_/X sky130_fd_sc_hd__and4_4
X_62877_ _63598_/A _62875_/X _62876_/Y _62877_/X sky130_fd_sc_hd__o21a_4
X_67404_ _84071_/Q _67331_/X _67403_/X _67404_/X sky130_fd_sc_hd__a21bo_4
X_52630_ _52630_/A _52657_/A sky130_fd_sc_hd__buf_2
X_64616_ _64616_/A _64769_/A sky130_fd_sc_hd__buf_2
X_83450_ _83451_/CLK _71578_/X _83450_/Q sky130_fd_sc_hd__dfxtp_4
X_61828_ _58241_/X _61824_/X _61756_/X _61790_/X _61827_/X _61828_/X
+ sky130_fd_sc_hd__a41o_4
X_80662_ _80657_/CLK _74828_/Y _46129_/A sky130_fd_sc_hd__dfxtp_4
X_68384_ _68384_/A _68384_/X sky130_fd_sc_hd__buf_2
X_65596_ _65595_/X _65596_/X sky130_fd_sc_hd__buf_2
X_82401_ _82965_/CLK _82209_/Q _82401_/Q sky130_fd_sc_hd__dfxtp_4
X_67335_ _67308_/A _87219_/Q _67335_/X sky130_fd_sc_hd__and2_4
X_52561_ _52542_/X _54079_/B _52561_/Y sky130_fd_sc_hd__nand2_4
X_64547_ _64250_/A _59443_/A _61102_/X _64547_/Y sky130_fd_sc_hd__nand3_4
X_83381_ _83414_/CLK _71773_/X _83381_/Q sky130_fd_sc_hd__dfxtp_4
X_61759_ _61356_/X _62183_/A _59810_/A _59754_/A _61766_/B sky130_fd_sc_hd__nand4_4
X_80593_ _80570_/Y _80592_/Y _80593_/Y sky130_fd_sc_hd__nor2_4
XPHY_408 sky130_fd_sc_hd__decap_3
X_54300_ _54314_/A _46676_/A _54300_/Y sky130_fd_sc_hd__nand2_4
XPHY_419 sky130_fd_sc_hd__decap_3
X_85120_ _85152_/CLK _85120_/D _45409_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_96_0_CLK clkbuf_7_96_0_CLK/A clkbuf_7_96_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_51512_ _51074_/A _51622_/A sky130_fd_sc_hd__buf_2
X_82332_ _82288_/CLK _77191_/B _82332_/Q sky130_fd_sc_hd__dfxtp_4
X_55280_ _55277_/X _55279_/X _55138_/X _56868_/A sky130_fd_sc_hd__a21o_4
X_67266_ _67266_/A _88118_/Q _67266_/X sky130_fd_sc_hd__and2_4
X_52492_ _52487_/X _46417_/B _52492_/Y sky130_fd_sc_hd__nand2_4
X_64478_ _61182_/X _61609_/X _64211_/C _64478_/Y sky130_fd_sc_hd__nand3_4
X_69005_ _86981_/Q _68472_/X _44246_/A _69004_/X _69005_/X sky130_fd_sc_hd__a211o_4
X_54231_ _85480_/Q _54220_/X _54230_/Y _54231_/Y sky130_fd_sc_hd__o21ai_4
X_66217_ _66217_/A _66216_/Y _66217_/Y sky130_fd_sc_hd__nand2_4
X_85051_ _85089_/CLK _85051_/D _85051_/Q sky130_fd_sc_hd__dfxtp_4
X_51443_ _51456_/A _51421_/X _51467_/C _52971_/D _51443_/X sky130_fd_sc_hd__and4_4
X_63429_ _61386_/B _63426_/X _63427_/X _63428_/X _63429_/X sky130_fd_sc_hd__a211o_4
X_82263_ _82263_/CLK _80522_/Y _82263_/Q sky130_fd_sc_hd__dfxtp_4
X_67197_ _67197_/A _67196_/X _67197_/Y sky130_fd_sc_hd__nand2_4
X_84002_ _81755_/CLK _84002_/D _84002_/Q sky130_fd_sc_hd__dfxtp_4
X_81214_ _84981_/CLK _74868_/X _48915_/A sky130_fd_sc_hd__dfxtp_4
X_54162_ _54149_/A _47344_/A _54162_/Y sky130_fd_sc_hd__nand2_4
X_66148_ _66145_/X _65967_/B _66147_/X _66148_/Y sky130_fd_sc_hd__nand3_4
X_51374_ _51364_/A _50862_/B _51374_/Y sky130_fd_sc_hd__nand2_4
X_82194_ _82386_/CLK _82194_/D _82194_/Q sky130_fd_sc_hd__dfxtp_4
X_53113_ _53133_/A _53113_/B _53107_/C _53113_/D _53113_/X sky130_fd_sc_hd__and4_4
X_50325_ _86223_/Q _50316_/X _50324_/Y _50325_/Y sky130_fd_sc_hd__o21ai_4
X_81145_ _81197_/CLK _75008_/A _81145_/Q sky130_fd_sc_hd__dfxtp_4
X_54093_ _53434_/A _47221_/A _54093_/Y sky130_fd_sc_hd__nand2_4
X_58970_ _58970_/A _58973_/B _58970_/Y sky130_fd_sc_hd__nand2_4
X_66079_ _66123_/A _66004_/B _84158_/Q _66079_/X sky130_fd_sc_hd__and3_4
X_57921_ _57912_/Y _57758_/X _57917_/X _57920_/X _84940_/D sky130_fd_sc_hd__a22oi_4
X_53044_ _53048_/A _53063_/B _53058_/C _53044_/D _53044_/X sky130_fd_sc_hd__and4_4
X_69907_ _87545_/Q _66608_/A _68348_/X _69906_/X _69907_/X sky130_fd_sc_hd__a211o_4
X_50256_ _50256_/A _50918_/A sky130_fd_sc_hd__buf_2
X_85953_ _85953_/CLK _51751_/Y _85953_/Q sky130_fd_sc_hd__dfxtp_4
X_81076_ _81087_/CLK _75889_/A _81076_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_7_34_0_CLK clkbuf_7_35_0_CLK/A clkbuf_8_69_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_84904_ _84903_/CLK _58223_/Y _63376_/B sky130_fd_sc_hd__dfxtp_4
X_80027_ _60107_/C _64088_/C _80027_/X sky130_fd_sc_hd__xor2_4
X_57852_ _57711_/X _57852_/X sky130_fd_sc_hd__buf_2
X_69838_ _69897_/A _69838_/B _69838_/Y sky130_fd_sc_hd__nor2_4
X_50187_ _51286_/A _50187_/X sky130_fd_sc_hd__buf_2
X_85884_ _85884_/CLK _85884_/D _65501_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_174_0_CLK clkbuf_7_87_0_CLK/X clkbuf_8_174_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_56803_ _56803_/A _57170_/B sky130_fd_sc_hd__buf_2
X_87623_ _87883_/CLK _42975_/Y _66861_/B sky130_fd_sc_hd__dfxtp_4
X_84835_ _84835_/CLK _84835_/D _64467_/C sky130_fd_sc_hd__dfxtp_4
X_57783_ _68342_/A _69182_/A sky130_fd_sc_hd__buf_2
X_69769_ _69765_/X _69767_/X _69768_/X _69772_/A sky130_fd_sc_hd__a21o_4
X_54995_ _54250_/A _55011_/A sky130_fd_sc_hd__buf_2
X_71800_ _71783_/Y _71800_/Y sky130_fd_sc_hd__inv_2
X_59522_ _59571_/B _59544_/A sky130_fd_sc_hd__buf_2
X_56734_ _56674_/X _57149_/D sky130_fd_sc_hd__buf_2
X_87554_ _88060_/CLK _43158_/Y _73198_/A sky130_fd_sc_hd__dfxtp_4
X_41960_ _42013_/A _41960_/X sky130_fd_sc_hd__buf_2
X_53946_ _53951_/A _53946_/B _53946_/Y sky130_fd_sc_hd__nand2_4
X_72780_ _72744_/X _86208_/Q _72746_/X _72779_/X _72780_/X sky130_fd_sc_hd__a211o_4
X_84766_ _84766_/CLK _59142_/Y _84766_/Q sky130_fd_sc_hd__dfxtp_4
X_81978_ _82234_/CLK _81978_/D _81978_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_290_0_CLK clkbuf_9_291_0_CLK/A clkbuf_9_290_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_7_49_0_CLK clkbuf_6_24_0_CLK/X clkbuf_8_99_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_86505_ _86505_/CLK _86505_/D _86505_/Q sky130_fd_sc_hd__dfxtp_4
X_40911_ _40911_/A _40911_/Y sky130_fd_sc_hd__inv_2
X_71731_ _71729_/A _71313_/X _71724_/X _71731_/Y sky130_fd_sc_hd__nand3_4
X_59453_ _84728_/Q _59454_/A sky130_fd_sc_hd__inv_2
X_83717_ _83721_/CLK _70720_/Y _83717_/Q sky130_fd_sc_hd__dfxtp_4
X_56665_ _56664_/Y _56665_/Y sky130_fd_sc_hd__inv_2
X_80929_ _80928_/CLK _84105_/Q _80929_/Q sky130_fd_sc_hd__dfxtp_4
X_87485_ _88001_/CLK _43315_/X _87485_/Q sky130_fd_sc_hd__dfxtp_4
X_41891_ _41967_/A _41891_/X sky130_fd_sc_hd__buf_2
X_53877_ _53848_/A _53877_/B _53877_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_189_0_CLK clkbuf_7_94_0_CLK/X clkbuf_9_378_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_84697_ _84329_/CLK _59804_/X _80455_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_184_0_CLK clkbuf_9_92_0_CLK/X _81282_/CLK sky130_fd_sc_hd__clkbuf_1
X_58404_ _58388_/X _83369_/Q _58403_/Y _84857_/D sky130_fd_sc_hd__o21a_4
X_43630_ _87334_/Q _68695_/B sky130_fd_sc_hd__inv_2
X_55616_ _55608_/X _55613_/X _55615_/X _55616_/X sky130_fd_sc_hd__a21o_4
X_74450_ _74448_/Y _72107_/X _74449_/Y _83064_/D sky130_fd_sc_hd__a21boi_4
X_86436_ _86436_/CLK _49183_/Y _65357_/B sky130_fd_sc_hd__dfxtp_4
X_52828_ _52824_/Y _52809_/X _52827_/X _52828_/Y sky130_fd_sc_hd__a21oi_4
X_40842_ _48904_/A _40842_/X sky130_fd_sc_hd__buf_2
X_71662_ _71660_/A _71256_/B _71660_/C _71662_/Y sky130_fd_sc_hd__nand3_4
X_83648_ _82774_/CLK _70965_/Y _83648_/Q sky130_fd_sc_hd__dfxtp_4
X_59384_ _59380_/Y _59383_/Y _59351_/X _59384_/X sky130_fd_sc_hd__a21o_4
X_56596_ _56596_/A _72652_/C sky130_fd_sc_hd__buf_2
X_73401_ _73353_/A _85864_/Q _73401_/X sky130_fd_sc_hd__and2_4
X_70613_ _70719_/A _70613_/B _70620_/C _70594_/X _70613_/Y sky130_fd_sc_hd__nand4_4
X_58335_ _58335_/A _58335_/Y sky130_fd_sc_hd__inv_2
X_43561_ _43217_/A _43561_/X sky130_fd_sc_hd__buf_2
X_55547_ _55477_/A _85144_/Q _55547_/X sky130_fd_sc_hd__and2_4
X_74381_ _74381_/A _72113_/B _74366_/C _74381_/X sky130_fd_sc_hd__and3_4
X_86367_ _83721_/CLK _86367_/D _86367_/Q sky130_fd_sc_hd__dfxtp_4
X_40773_ _40585_/A _40773_/X sky130_fd_sc_hd__buf_2
X_52759_ _52753_/Y _52755_/X _52758_/X _52759_/Y sky130_fd_sc_hd__a21oi_4
X_71593_ _71581_/X _83445_/Q _71592_/Y _83445_/D sky130_fd_sc_hd__a21o_4
X_83579_ _86193_/CLK _71184_/Y _83579_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_112_0_CLK clkbuf_7_56_0_CLK/X clkbuf_8_112_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_45300_ _85159_/Q _45284_/X _45265_/X _45300_/X sky130_fd_sc_hd__o21a_4
X_76120_ _76117_/Y _76119_/Y _76121_/B sky130_fd_sc_hd__xor2_4
X_42512_ _42511_/Y _42512_/Y sky130_fd_sc_hd__inv_2
X_88106_ _88111_/CLK _41917_/Y _88106_/Q sky130_fd_sc_hd__dfxtp_4
X_73332_ _72908_/X _85579_/Q _72909_/X _73331_/X _73332_/X sky130_fd_sc_hd__a211o_4
X_85318_ _85317_/CLK _85318_/D _85318_/Q sky130_fd_sc_hd__dfxtp_4
X_46280_ _46280_/A _46326_/A sky130_fd_sc_hd__buf_2
X_70544_ _70543_/Y _71586_/A sky130_fd_sc_hd__buf_2
X_58266_ _58253_/X _83445_/Q _58265_/Y _84893_/D sky130_fd_sc_hd__o21a_4
X_55478_ _82995_/Q _55475_/X _44097_/X _55477_/X _55478_/X sky130_fd_sc_hd__a211o_4
X_43492_ _41721_/X _43484_/X _87394_/Q _43485_/X _43492_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_10_199_0_CLK clkbuf_9_99_0_CLK/X _84672_/CLK sky130_fd_sc_hd__clkbuf_1
X_86298_ _86297_/CLK _86298_/D _86298_/Q sky130_fd_sc_hd__dfxtp_4
X_45231_ _83020_/Q _45232_/A sky130_fd_sc_hd__inv_2
X_57217_ _57179_/A _57217_/B _57217_/Y sky130_fd_sc_hd__nand2_4
X_76051_ _76042_/Y _76049_/Y _76050_/Y _76051_/X sky130_fd_sc_hd__o21a_4
X_88037_ _88044_/CLK _88037_/D _88037_/Q sky130_fd_sc_hd__dfxtp_4
X_54429_ _54435_/A _54417_/B _54429_/C _46894_/Y _54429_/X sky130_fd_sc_hd__and4_4
X_42443_ _40542_/X _42434_/X _87861_/Q _42435_/X _87861_/D sky130_fd_sc_hd__a2bb2o_4
X_73263_ _73259_/X _73261_/X _73262_/X _73267_/A sky130_fd_sc_hd__a21o_4
X_85249_ _85249_/CLK _85249_/D _56287_/C sky130_fd_sc_hd__dfxtp_4
X_70475_ _71483_/B _70483_/B sky130_fd_sc_hd__buf_2
X_58197_ _84910_/Q _58198_/A sky130_fd_sc_hd__buf_2
X_75002_ _81143_/D _75003_/B _75002_/Y sky130_fd_sc_hd__nor2_4
X_72214_ _72214_/A _72214_/Y sky130_fd_sc_hd__inv_2
X_45162_ _55836_/B _45131_/X _45161_/X _45162_/X sky130_fd_sc_hd__o21a_4
X_57148_ _57147_/X _85072_/D sky130_fd_sc_hd__inv_2
X_42374_ _42373_/X _42374_/X sky130_fd_sc_hd__buf_2
X_73194_ _72725_/A _73194_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_127_0_CLK clkbuf_7_63_0_CLK/X clkbuf_9_255_0_CLK/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_122_0_CLK clkbuf_9_61_0_CLK/X _84287_/CLK sky130_fd_sc_hd__clkbuf_1
X_44113_ _44112_/X _44113_/X sky130_fd_sc_hd__buf_2
X_79810_ _79782_/X _79785_/Y _79795_/X _79798_/Y _79810_/X sky130_fd_sc_hd__o22a_4
X_41325_ _41186_/A _41325_/X sky130_fd_sc_hd__buf_2
X_72145_ _72143_/X _85375_/Q _72144_/X _72145_/Y sky130_fd_sc_hd__o21ai_4
X_49970_ _49967_/Y _49951_/X _49969_/X _49970_/Y sky130_fd_sc_hd__a21oi_4
X_45093_ _55879_/B _45044_/X _45079_/X _45093_/X sky130_fd_sc_hd__o21a_4
X_57079_ _57319_/D _57318_/D sky130_fd_sc_hd__buf_2
Xclkbuf_10_752_0_CLK clkbuf_9_376_0_CLK/X _87260_/CLK sky130_fd_sc_hd__clkbuf_1
X_48921_ _48920_/Y _48922_/B sky130_fd_sc_hd__buf_2
X_44044_ _44043_/X _44044_/X sky130_fd_sc_hd__buf_2
X_79741_ _84220_/Q _83268_/Q _79741_/X sky130_fd_sc_hd__xor2_4
X_41256_ _41186_/A _41280_/B sky130_fd_sc_hd__buf_2
X_60090_ _59971_/X _60003_/Y _60092_/B _60087_/Y _60089_/Y _84664_/D
+ sky130_fd_sc_hd__a41oi_4
X_72076_ _72073_/Y _72033_/X _72075_/Y _83290_/D sky130_fd_sc_hd__a21boi_4
X_76953_ _76953_/A _76953_/B _76951_/A _76957_/C sky130_fd_sc_hd__nand3_4
Xclkbuf_9_243_0_CLK clkbuf_9_243_0_CLK/A clkbuf_9_243_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_71027_ _71173_/A _71030_/B _71030_/C _71018_/D _71027_/Y sky130_fd_sc_hd__nand4_4
X_75904_ _84502_/Q _84374_/Q _75904_/X sky130_fd_sc_hd__xor2_4
X_48852_ _86470_/Q _48836_/X _48851_/Y _48852_/Y sky130_fd_sc_hd__o21ai_4
X_79672_ _79670_/X _79677_/B _79672_/Y sky130_fd_sc_hd__xnor2_4
X_41187_ _81715_/Q _41197_/B _41187_/X sky130_fd_sc_hd__or2_4
X_76884_ _81676_/Q _76884_/B _76884_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_10_137_0_CLK clkbuf_9_68_0_CLK/X _81260_/CLK sky130_fd_sc_hd__clkbuf_1
X_47803_ _47803_/A _53253_/D sky130_fd_sc_hd__buf_2
X_78623_ _78623_/A _78623_/B _78640_/B sky130_fd_sc_hd__nand2_4
X_75835_ _75793_/B _75832_/X _75834_/X _75836_/B sky130_fd_sc_hd__a21boi_4
Xclkbuf_10_767_0_CLK clkbuf_9_383_0_CLK/X _87544_/CLK sky130_fd_sc_hd__clkbuf_1
X_48783_ _48793_/A _50466_/B _48783_/Y sky130_fd_sc_hd__nand2_4
X_45995_ _45981_/X _45995_/X sky130_fd_sc_hd__buf_2
X_62800_ _62679_/X _62834_/B sky130_fd_sc_hd__buf_2
X_47734_ _54907_/B _53213_/B sky130_fd_sc_hd__buf_2
X_78554_ _78554_/A _78554_/B _78555_/A sky130_fd_sc_hd__nor2_4
X_44946_ _55960_/B _44882_/X _44884_/X _44946_/X sky130_fd_sc_hd__o21a_4
X_63780_ _61762_/X _63738_/B _63738_/C _63738_/D _63780_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_9_258_0_CLK clkbuf_9_259_0_CLK/A clkbuf_9_258_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_75766_ _75766_/A _75765_/Y _80887_/D sky130_fd_sc_hd__xnor2_4
X_60992_ _60910_/B _60992_/X sky130_fd_sc_hd__buf_2
X_72978_ _72978_/A _72978_/X sky130_fd_sc_hd__buf_2
X_77505_ _82229_/Q _77505_/Y sky130_fd_sc_hd__inv_2
X_62731_ _62731_/A _63081_/A _62704_/C _62717_/X _62731_/X sky130_fd_sc_hd__and4_4
X_74717_ _71266_/A _74739_/B sky130_fd_sc_hd__buf_2
X_47665_ _47660_/Y _47651_/X _47664_/X _86611_/D sky130_fd_sc_hd__a21oi_4
X_71929_ _57010_/Y _71917_/X _71928_/Y _83325_/D sky130_fd_sc_hd__o21ai_4
X_78485_ _78484_/Y _78485_/Y sky130_fd_sc_hd__inv_2
X_44877_ _56192_/C _45604_/B _44876_/X _44877_/Y sky130_fd_sc_hd__o21ai_4
X_75697_ _75685_/A _75692_/A _75697_/X sky130_fd_sc_hd__and2_4
X_49404_ _86393_/Q _49388_/X _49403_/Y _49404_/Y sky130_fd_sc_hd__o21ai_4
X_46616_ _46616_/A _46617_/A sky130_fd_sc_hd__buf_2
X_65450_ _65447_/Y _65448_/X _65449_/X _84200_/D sky130_fd_sc_hd__a21o_4
X_77436_ _77415_/X _77435_/Y _77436_/Y sky130_fd_sc_hd__nand2_4
X_43828_ _41134_/X _43817_/X _87247_/Q _43818_/X _43828_/X sky130_fd_sc_hd__a2bb2o_4
X_74648_ _56613_/A _74641_/X _74647_/Y _83001_/D sky130_fd_sc_hd__a21boi_4
X_62662_ _62646_/B _62664_/B sky130_fd_sc_hd__buf_2
X_47596_ _47592_/Y _47555_/X _47595_/X _86618_/D sky130_fd_sc_hd__a21oi_4
X_64401_ _64377_/X _64401_/B _64391_/X _64401_/X sky130_fd_sc_hd__and3_4
X_49335_ _48535_/A _49352_/A sky130_fd_sc_hd__buf_2
X_61613_ _61613_/A _61613_/Y sky130_fd_sc_hd__inv_2
X_46547_ _46547_/A _50858_/B _46547_/Y sky130_fd_sc_hd__nand2_4
X_65381_ _65381_/A _65381_/B _65381_/X sky130_fd_sc_hd__and2_4
X_77367_ _77376_/A _77376_/B _77367_/X sky130_fd_sc_hd__xor2_4
X_43759_ _40955_/X _43752_/X _69179_/B _43753_/X _87280_/D sky130_fd_sc_hd__a2bb2o_4
X_62593_ _62395_/X _62593_/X sky130_fd_sc_hd__buf_2
X_74579_ _45108_/A _74568_/X _74578_/X _74579_/Y sky130_fd_sc_hd__o21ai_4
X_67120_ _68057_/A _67120_/X sky130_fd_sc_hd__buf_2
X_79106_ _82657_/Q _82529_/D _79107_/A sky130_fd_sc_hd__xor2_4
X_64332_ _64304_/A _64303_/X _84959_/Q _64318_/D _64332_/X sky130_fd_sc_hd__and4_4
X_76318_ _76311_/A _76296_/A _76319_/A sky130_fd_sc_hd__nor2_4
X_49266_ _86421_/Q _49255_/X _49265_/Y _49266_/Y sky130_fd_sc_hd__o21ai_4
X_61544_ _61544_/A _61544_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_705_0_CLK clkbuf_9_352_0_CLK/X _86814_/CLK sky130_fd_sc_hd__clkbuf_1
X_46478_ _46491_/A _50827_/B _46478_/Y sky130_fd_sc_hd__nand2_4
X_77298_ _77295_/X _77296_/Y _77297_/Y _77301_/A sky130_fd_sc_hd__a21oi_4
X_48217_ _50270_/A _48201_/B _48195_/X _48217_/X sky130_fd_sc_hd__and3_4
X_67051_ _67048_/X _67050_/X _67026_/X _67051_/X sky130_fd_sc_hd__a21o_4
X_79037_ _79027_/B _79027_/A _79037_/C _79044_/A sky130_fd_sc_hd__nand3_4
X_45429_ _44887_/X _45429_/X sky130_fd_sc_hd__buf_2
X_64263_ _64263_/A _64287_/A sky130_fd_sc_hd__buf_2
X_76249_ _76245_/Y _76247_/Y _76248_/Y _76254_/A sky130_fd_sc_hd__o21ai_4
X_49197_ _49156_/X _50721_/B _49197_/Y sky130_fd_sc_hd__nand2_4
X_61475_ _72176_/A _61476_/A sky130_fd_sc_hd__buf_2
X_66002_ _66002_/A _66003_/A sky130_fd_sc_hd__buf_2
X_63214_ _63288_/A _64420_/B _63165_/X _63192_/D _63214_/X sky130_fd_sc_hd__and4_4
X_48148_ _48801_/A _48148_/B _48148_/X sky130_fd_sc_hd__and2_4
X_60426_ _60417_/A _60441_/B _60473_/B _60383_/A _60427_/A sky130_fd_sc_hd__and4_4
X_64194_ _62186_/X _64182_/B _64182_/C _64182_/D _64194_/Y sky130_fd_sc_hd__nand4_4
X_63145_ _60606_/X _63146_/C sky130_fd_sc_hd__buf_2
X_60357_ _60477_/A _60319_/X _79605_/A _60357_/Y sky130_fd_sc_hd__nor3_4
X_48079_ _47981_/X _48079_/B _48079_/X sky130_fd_sc_hd__and2_4
X_50110_ _50106_/A _72014_/B _50110_/X sky130_fd_sc_hd__and2_4
X_51090_ _51087_/Y _51065_/X _51089_/X _86076_/D sky130_fd_sc_hd__a21oi_4
X_67953_ _68640_/A _67953_/X sky130_fd_sc_hd__buf_2
X_63076_ _60458_/X _63077_/D sky130_fd_sc_hd__buf_2
X_79939_ _84925_/Q _65855_/C _79939_/Y sky130_fd_sc_hd__nor2_4
X_60288_ _62644_/A _60251_/A _60288_/C _60288_/X sky130_fd_sc_hd__and3_4
X_50041_ _50039_/Y _50029_/X _50040_/X _86276_/D sky130_fd_sc_hd__a21oi_4
X_66904_ _87429_/Q _66878_/X _66879_/X _66903_/X _66904_/X sky130_fd_sc_hd__a211o_4
X_62027_ _62027_/A _62027_/X sky130_fd_sc_hd__buf_2
X_82950_ _82774_/CLK _82758_/Q _82950_/Q sky130_fd_sc_hd__dfxtp_4
X_67884_ _67881_/X _67883_/X _67858_/X _67887_/A sky130_fd_sc_hd__a21o_4
X_81901_ _81989_/CLK _77390_/X _82277_/D sky130_fd_sc_hd__dfxtp_4
X_69623_ _72859_/A _68394_/A _68741_/X _69622_/Y _69623_/X sky130_fd_sc_hd__a211o_4
X_66835_ _66769_/A _88200_/Q _66835_/X sky130_fd_sc_hd__and2_4
X_82881_ _82368_/CLK _78303_/B _82881_/Q sky130_fd_sc_hd__dfxtp_4
X_53800_ _53900_/A _53801_/B sky130_fd_sc_hd__buf_2
X_84620_ _84620_/CLK _60370_/Y _79553_/A sky130_fd_sc_hd__dfxtp_4
X_69554_ _88020_/Q _69424_/X _69465_/X _69553_/X _69554_/X sky130_fd_sc_hd__a211o_4
X_81832_ _82084_/CLK _81864_/Q _77305_/A sky130_fd_sc_hd__dfxtp_4
X_54780_ _54672_/X _54798_/C sky130_fd_sc_hd__buf_2
X_66766_ _87435_/Q _66762_/X _66764_/X _66765_/X _66766_/X sky130_fd_sc_hd__a211o_4
X_51992_ _51982_/X _53516_/B _51992_/Y sky130_fd_sc_hd__nand2_4
X_63978_ _60920_/A _64040_/C sky130_fd_sc_hd__buf_2
X_68505_ _68452_/A _87246_/Q _68505_/X sky130_fd_sc_hd__and2_4
X_53731_ _53750_/A _48602_/Y _53731_/Y sky130_fd_sc_hd__nand2_4
X_65717_ _65859_/A _65717_/X sky130_fd_sc_hd__buf_2
X_84551_ _84292_/CLK _84551_/D _76999_/A sky130_fd_sc_hd__dfxtp_4
X_50943_ _50938_/X _51807_/B _50943_/Y sky130_fd_sc_hd__nand2_4
X_62929_ _62923_/Y _62924_/X _62928_/Y _58344_/A _62650_/X _62929_/Y
+ sky130_fd_sc_hd__o32ai_4
X_81763_ _88116_/CLK _75982_/X _48697_/A sky130_fd_sc_hd__dfxtp_4
X_69485_ _69485_/A _69485_/X sky130_fd_sc_hd__buf_2
X_66697_ _69582_/A _66697_/X sky130_fd_sc_hd__buf_2
X_83502_ _84228_/CLK _83502_/D _83502_/Q sky130_fd_sc_hd__dfxtp_4
X_56450_ _56377_/X _56454_/B _56450_/C _56450_/Y sky130_fd_sc_hd__nand3_4
X_80714_ _80681_/CLK _75900_/X _80682_/D sky130_fd_sc_hd__dfxtp_4
X_68436_ _65976_/A _68436_/X sky130_fd_sc_hd__buf_2
X_87270_ _87782_/CLK _43783_/Y _69318_/B sky130_fd_sc_hd__dfxtp_4
X_53662_ _53755_/A _53662_/X sky130_fd_sc_hd__buf_2
X_65648_ _65533_/X _65646_/Y _65647_/Y _65648_/Y sky130_fd_sc_hd__o21ai_4
X_84482_ _84481_/CLK _61426_/Y _79150_/B sky130_fd_sc_hd__dfxtp_4
X_50874_ _50857_/X _51389_/B _50874_/Y sky130_fd_sc_hd__nand2_4
X_81694_ _81695_/CLK _80228_/X _76755_/A sky130_fd_sc_hd__dfxtp_4
X_55401_ _55399_/X _55181_/B _55400_/Y _55403_/A sky130_fd_sc_hd__a21o_4
X_86221_ _85599_/CLK _86221_/D _86221_/Q sky130_fd_sc_hd__dfxtp_4
X_52613_ _85786_/Q _52601_/X _52612_/Y _52613_/Y sky130_fd_sc_hd__o21ai_4
X_83433_ _83372_/CLK _71627_/X _83433_/Q sky130_fd_sc_hd__dfxtp_4
X_56381_ _56458_/A _56363_/B _56381_/C _56381_/Y sky130_fd_sc_hd__nand3_4
X_80645_ _74767_/X _74709_/Y DATA_FROM_HASH[2] sky130_fd_sc_hd__ebufn_2
X_68367_ _68366_/X _43587_/Y _68367_/Y sky130_fd_sc_hd__nor2_4
X_53593_ _53601_/A _53593_/B _53593_/Y sky130_fd_sc_hd__nand2_4
X_65579_ _65438_/X _86199_/Q _65576_/X _65578_/X _65579_/X sky130_fd_sc_hd__a211o_4
X_58120_ _84923_/Q _79903_/A sky130_fd_sc_hd__inv_2
XPHY_205 sky130_fd_sc_hd__decap_3
X_55332_ _55317_/A _57414_/A _55332_/X sky130_fd_sc_hd__and2_4
X_67318_ _87924_/Q _67293_/X _67271_/X _67317_/X _67318_/X sky130_fd_sc_hd__a211o_4
X_86152_ _86155_/CLK _50696_/Y _86152_/Q sky130_fd_sc_hd__dfxtp_4
X_52544_ _52540_/Y _52541_/X _52543_/Y _52544_/Y sky130_fd_sc_hd__a21boi_4
XPHY_216 sky130_fd_sc_hd__decap_3
X_83364_ _83362_/CLK _83364_/D _83364_/Q sky130_fd_sc_hd__dfxtp_4
X_80576_ _84772_/Q _84164_/Q _80576_/Y sky130_fd_sc_hd__nand2_4
XPHY_227 sky130_fd_sc_hd__decap_3
X_68298_ _83989_/Q _68279_/X _68297_/X _68298_/X sky130_fd_sc_hd__a21bo_4
XPHY_238 sky130_fd_sc_hd__decap_3
X_85103_ _85103_/CLK _85103_/D _45673_/A sky130_fd_sc_hd__dfxtp_4
XPHY_249 sky130_fd_sc_hd__decap_3
X_58051_ _57947_/X _85705_/Q _57948_/X _58051_/X sky130_fd_sc_hd__o21a_4
X_82315_ _81195_/CLK _77065_/B _82315_/Q sky130_fd_sc_hd__dfxtp_4
X_55263_ _55264_/A _55264_/C _83321_/Q _55263_/X sky130_fd_sc_hd__a21o_4
X_67249_ _87927_/Q _67176_/X _67153_/X _67248_/X _67249_/X sky130_fd_sc_hd__a211o_4
X_86083_ _85764_/CLK _51052_/Y _86083_/Q sky130_fd_sc_hd__dfxtp_4
X_52475_ _52473_/Y _52462_/X _52474_/Y _52475_/Y sky130_fd_sc_hd__a21boi_4
X_83295_ _85538_/CLK _72050_/Y _83295_/Q sky130_fd_sc_hd__dfxtp_4
X_57002_ _56758_/X _56730_/X _56740_/X _56994_/D _57003_/B _57004_/B
+ sky130_fd_sc_hd__a41oi_4
X_54214_ _54212_/Y _54197_/X _54213_/X _85483_/D sky130_fd_sc_hd__a21oi_4
X_85034_ _85034_/CLK _57330_/Y _57326_/B sky130_fd_sc_hd__dfxtp_4
X_51426_ _51410_/X _51421_/X _51438_/C _52954_/D _51426_/X sky130_fd_sc_hd__and4_4
X_70260_ _70260_/A _70260_/B _70260_/C _70260_/D _70260_/X sky130_fd_sc_hd__and4_4
X_82246_ _82436_/CLK _82246_/D _82246_/Q sky130_fd_sc_hd__dfxtp_4
X_55194_ _55188_/X _55193_/X _83749_/Q _55196_/A sky130_fd_sc_hd__a21o_4
Xclkbuf_opt_26_CLK _86505_/CLK _86186_/CLK sky130_fd_sc_hd__clkbuf_16
X_54145_ _49793_/A _54254_/A sky130_fd_sc_hd__buf_2
X_51357_ _51355_/Y _51339_/X _51356_/X _51357_/Y sky130_fd_sc_hd__a21oi_4
X_82177_ _82177_/CLK _65916_/C _82177_/Q sky130_fd_sc_hd__dfxtp_4
X_70191_ _70169_/X _83843_/Q _70190_/X _70191_/X sky130_fd_sc_hd__a21o_4
X_41110_ _40989_/A _41110_/X sky130_fd_sc_hd__buf_2
X_50308_ _50308_/A _74509_/C _50247_/X _50308_/X sky130_fd_sc_hd__and3_4
X_81128_ _81125_/CLK _81128_/D _40727_/A sky130_fd_sc_hd__dfxtp_4
X_42090_ _42083_/X _42077_/X _41004_/X _88039_/Q _42078_/X _42090_/Y
+ sky130_fd_sc_hd__o32ai_4
X_58953_ _58953_/A _59090_/B _58953_/Y sky130_fd_sc_hd__nor2_4
X_54076_ _54074_/Y _54060_/X _54075_/Y _85510_/D sky130_fd_sc_hd__a21boi_4
X_51288_ _64874_/B _51285_/X _51287_/Y _51288_/Y sky130_fd_sc_hd__o21ai_4
X_86985_ _82538_/CLK _44726_/Y _44725_/A sky130_fd_sc_hd__dfxtp_4
X_41041_ _40946_/A _41041_/X sky130_fd_sc_hd__buf_2
X_53027_ _52754_/A _53111_/A sky130_fd_sc_hd__buf_2
X_57904_ _57903_/X _85493_/Q _57849_/X _57904_/X sky130_fd_sc_hd__o21a_4
X_50239_ _50213_/X _50240_/A sky130_fd_sc_hd__buf_2
X_73950_ _73850_/X _86225_/Q _73948_/X _73949_/X _73950_/X sky130_fd_sc_hd__a211o_4
X_85936_ _86096_/CLK _51845_/Y _85936_/Q sky130_fd_sc_hd__dfxtp_4
X_81059_ _81059_/CLK _81091_/Q _75085_/B sky130_fd_sc_hd__dfxtp_4
X_58884_ _58879_/Y _58881_/Y _58883_/X _58884_/X sky130_fd_sc_hd__a21o_4
X_72901_ _72739_/X _72901_/X sky130_fd_sc_hd__buf_2
X_57835_ _57824_/X _85498_/Q _57736_/X _57835_/X sky130_fd_sc_hd__o21a_4
X_73881_ _73854_/X _85620_/Q _73782_/X _73880_/X _73881_/X sky130_fd_sc_hd__a211o_4
X_85867_ _86506_/CLK _52213_/Y _85867_/Q sky130_fd_sc_hd__dfxtp_4
X_44800_ _41436_/Y _44788_/X _86947_/Q _44789_/X _86947_/D sky130_fd_sc_hd__a2bb2o_4
X_75620_ _75640_/A _75609_/Y _75620_/Y sky130_fd_sc_hd__nor2_4
X_87606_ _87348_/CLK _87606_/D _67259_/B sky130_fd_sc_hd__dfxtp_4
X_72832_ _43119_/Y _72830_/X _72799_/X _72831_/Y _72832_/X sky130_fd_sc_hd__a211o_4
X_84818_ _84877_/CLK _84818_/D _84818_/Q sky130_fd_sc_hd__dfxtp_4
X_45780_ _57199_/A _45354_/X _45395_/X _45780_/X sky130_fd_sc_hd__o21a_4
X_57766_ _44019_/A _64567_/A sky130_fd_sc_hd__buf_2
X_54978_ _54927_/A _54978_/X sky130_fd_sc_hd__buf_2
X_42992_ _42992_/A _42992_/Y sky130_fd_sc_hd__inv_2
X_85798_ _86119_/CLK _85798_/D _65298_/B sky130_fd_sc_hd__dfxtp_4
X_59505_ _64295_/C _63448_/B sky130_fd_sc_hd__buf_2
X_56717_ _57416_/A _57416_/C _56764_/B _56717_/Y sky130_fd_sc_hd__a21oi_4
X_44731_ _86982_/Q _44731_/Y sky130_fd_sc_hd__inv_2
X_75551_ _80800_/Q _75551_/B _80768_/D sky130_fd_sc_hd__xnor2_4
X_87537_ _87544_/CLK _43209_/Y _87537_/Q sky130_fd_sc_hd__dfxtp_4
X_53929_ _53929_/A _53949_/A sky130_fd_sc_hd__buf_2
X_41943_ _41932_/X _41927_/X _40682_/X _73963_/A _41928_/X _41944_/A
+ sky130_fd_sc_hd__o32ai_4
X_72763_ _72738_/X _72764_/C _72762_/X _72763_/X sky130_fd_sc_hd__a21o_4
X_84749_ _86665_/CLK _84749_/D _84749_/Q sky130_fd_sc_hd__dfxtp_4
X_57697_ _57696_/X _57697_/X sky130_fd_sc_hd__buf_2
X_74502_ _74500_/Y _74492_/X _74501_/X _74502_/Y sky130_fd_sc_hd__a21oi_4
X_47450_ _83729_/Q _47451_/A sky130_fd_sc_hd__inv_2
X_71714_ _71823_/A _71713_/Y _71714_/Y sky130_fd_sc_hd__nor2_4
X_59436_ _64526_/B _59436_/Y sky130_fd_sc_hd__inv_2
X_78270_ _82684_/Q _78270_/B _78270_/X sky130_fd_sc_hd__xor2_4
X_44662_ _44662_/A _87012_/D sky130_fd_sc_hd__inv_2
X_56648_ _55491_/A _55490_/X _55676_/B _56972_/A sky130_fd_sc_hd__a21bo_4
X_75482_ _75477_/X _75480_/Y _75478_/Y _75482_/Y sky130_fd_sc_hd__nand3_4
X_87468_ _87708_/CLK _87468_/D _87468_/Q sky130_fd_sc_hd__dfxtp_4
X_41874_ _41873_/Y _88115_/D sky130_fd_sc_hd__inv_2
X_72694_ _70236_/C _72686_/X _72693_/Y _83187_/D sky130_fd_sc_hd__a21bo_4
X_46401_ _46401_/A _46408_/A sky130_fd_sc_hd__buf_2
X_77221_ _77219_/B _77219_/A _77223_/A sky130_fd_sc_hd__nand2_4
X_43613_ _43613_/A _43613_/Y sky130_fd_sc_hd__inv_2
X_74433_ _74413_/X _48514_/A _74433_/Y sky130_fd_sc_hd__nand2_4
X_86419_ _86422_/CLK _86419_/D _86419_/Q sky130_fd_sc_hd__dfxtp_4
X_40825_ _40783_/X _82293_/Q _40824_/X _40826_/A sky130_fd_sc_hd__o21a_4
X_47381_ _47375_/Y _47364_/X _47380_/X _47381_/Y sky130_fd_sc_hd__a21oi_4
X_59367_ _59231_/X _85411_/Q _59366_/X _59367_/Y sky130_fd_sc_hd__o21ai_4
X_71645_ _59500_/Y _71628_/A _71644_/Y _71645_/Y sky130_fd_sc_hd__o21ai_4
X_56579_ _56568_/X _56578_/X _55599_/B _56572_/X _85150_/D sky130_fd_sc_hd__a2bb2o_4
X_44593_ _44529_/A _44593_/X sky130_fd_sc_hd__buf_2
X_87399_ _86932_/CLK _87399_/D _87399_/Q sky130_fd_sc_hd__dfxtp_4
X_49120_ _49018_/X _48618_/Y _49119_/Y _49121_/A sky130_fd_sc_hd__a21o_4
X_46332_ _46327_/Y _46258_/X _46331_/Y _46332_/Y sky130_fd_sc_hd__a21boi_4
X_58318_ _58310_/X _83456_/Q _58317_/Y _84880_/D sky130_fd_sc_hd__o21a_4
X_77152_ _77152_/A _77152_/B _77152_/X sky130_fd_sc_hd__xor2_4
X_43544_ _43544_/A _43544_/Y sky130_fd_sc_hd__inv_2
X_74364_ _83081_/Q _72066_/X _74363_/Y _74364_/Y sky130_fd_sc_hd__o21ai_4
X_40756_ _40756_/A _40756_/X sky130_fd_sc_hd__buf_2
X_59298_ _59294_/Y _59296_/Y _59297_/X _59298_/X sky130_fd_sc_hd__a21o_4
X_71576_ _70570_/Y _71576_/X sky130_fd_sc_hd__buf_2
X_76103_ _76103_/A _76102_/Y _76104_/B sky130_fd_sc_hd__xor2_4
X_49051_ _49047_/Y _49038_/X _49050_/X _49051_/Y sky130_fd_sc_hd__a21oi_4
X_73315_ _73313_/X _73301_/X _73303_/X _73315_/Y sky130_fd_sc_hd__nand3_4
X_46263_ _46526_/A _46349_/A sky130_fd_sc_hd__buf_2
X_70527_ _57682_/Y _70500_/Y _70526_/Y _70527_/Y sky130_fd_sc_hd__o21ai_4
X_58249_ _58219_/X _58246_/Y _58248_/Y _84898_/D sky130_fd_sc_hd__a21oi_4
X_77083_ _77073_/A _77077_/A _77086_/B _77083_/X sky130_fd_sc_hd__and3_4
X_43475_ _43425_/X _43475_/X sky130_fd_sc_hd__buf_2
X_74295_ _74297_/A _74297_/B _56003_/B _74295_/Y sky130_fd_sc_hd__nand3_4
X_40687_ _40835_/A _40687_/X sky130_fd_sc_hd__buf_2
X_48002_ _83545_/Q _53535_/B sky130_fd_sc_hd__inv_2
X_45214_ _85293_/Q _45194_/X _45153_/X _45214_/X sky130_fd_sc_hd__o21a_4
X_76034_ _76024_/A _76028_/A _76028_/B _76034_/X sky130_fd_sc_hd__and3_4
X_42426_ _42417_/X _42410_/X _40501_/X _87869_/Q _42411_/X _42427_/A
+ sky130_fd_sc_hd__o32ai_4
X_61260_ _61260_/A _61260_/X sky130_fd_sc_hd__buf_2
X_73246_ _83159_/Q _73193_/X _73245_/Y _83159_/D sky130_fd_sc_hd__a21o_4
X_70458_ _70457_/X _70458_/X sky130_fd_sc_hd__buf_2
X_46194_ _46143_/D _46222_/B _46128_/D _46133_/C _46195_/D sky130_fd_sc_hd__nand4_4
Xclkbuf_10_691_0_CLK clkbuf_9_345_0_CLK/X _87636_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_opt_17_CLK _85535_/CLK _85556_/CLK sky130_fd_sc_hd__clkbuf_16
X_60211_ _60211_/A _60309_/D _60212_/A sky130_fd_sc_hd__nand2_4
X_45145_ _45127_/X _61509_/B _45144_/X _45145_/Y sky130_fd_sc_hd__o21ai_4
X_42357_ _42304_/X _42357_/X sky130_fd_sc_hd__buf_2
X_61191_ _72543_/A _61234_/A sky130_fd_sc_hd__buf_2
X_73177_ _87555_/Q _72758_/X _73177_/Y sky130_fd_sc_hd__nor2_4
X_70389_ _70366_/X _74527_/A _70375_/C _70389_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_9_182_0_CLK clkbuf_8_91_0_CLK/X clkbuf_9_182_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_41308_ _41253_/A _41308_/X sky130_fd_sc_hd__buf_2
X_60142_ _79936_/B _79937_/A sky130_fd_sc_hd__inv_2
X_72128_ _59326_/X _72128_/B _72128_/Y sky130_fd_sc_hd__nor2_4
X_49953_ _49973_/A _49943_/B _49953_/C _53165_/D _49953_/X sky130_fd_sc_hd__and4_4
X_45076_ _56494_/C _45060_/X _45040_/X _45076_/X sky130_fd_sc_hd__o21a_4
X_42288_ _41552_/X _42271_/X _87938_/Q _42272_/X _87938_/D sky130_fd_sc_hd__a2bb2o_4
X_77985_ _82078_/Q _77999_/A sky130_fd_sc_hd__inv_2
X_48904_ _48904_/A _48976_/A sky130_fd_sc_hd__buf_2
X_44027_ _44247_/A _69654_/A sky130_fd_sc_hd__buf_2
X_79724_ _79720_/X _79724_/B _79724_/X sky130_fd_sc_hd__xor2_4
X_64950_ _64947_/X _64949_/X _64851_/X _64953_/A sky130_fd_sc_hd__a21o_4
X_41239_ _40999_/A _41239_/X sky130_fd_sc_hd__buf_2
X_72059_ _71978_/A _72059_/X sky130_fd_sc_hd__buf_2
X_76936_ _81503_/Q _76933_/Y _76935_/X _76936_/Y sky130_fd_sc_hd__o21ai_4
X_60073_ _60072_/Y _60073_/Y sky130_fd_sc_hd__inv_2
X_49884_ _49893_/A _49884_/B _49893_/C _53099_/D _49884_/X sky130_fd_sc_hd__and4_4
X_63901_ _64334_/B _63920_/B _63840_/C _63920_/D _63901_/Y sky130_fd_sc_hd__nand4_4
X_48835_ _48832_/Y _48813_/X _48834_/X _86474_/D sky130_fd_sc_hd__a21oi_4
X_79655_ _84211_/Q _83259_/Q _79655_/Y sky130_fd_sc_hd__nand2_4
X_64881_ _64826_/A _85847_/Q _64881_/X sky130_fd_sc_hd__and2_4
X_76867_ _76857_/Y _76867_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_9_197_0_CLK clkbuf_8_98_0_CLK/X clkbuf_9_197_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_66620_ _66617_/X _66619_/X _66547_/X _66620_/X sky130_fd_sc_hd__a21o_4
X_78606_ _78599_/X _78605_/Y _82774_/D sky130_fd_sc_hd__xor2_4
X_63832_ _63823_/X _63810_/X _63825_/Y _63828_/Y _63831_/X _63832_/X
+ sky130_fd_sc_hd__a41o_4
X_75818_ _75818_/A _75817_/Y _75821_/A sky130_fd_sc_hd__nor2_4
X_48766_ _50447_/A _48766_/B _48786_/C _48766_/X sky130_fd_sc_hd__and3_4
X_79586_ _79586_/A _79585_/Y _79587_/B sky130_fd_sc_hd__nand2_4
X_45978_ _40407_/Y _45974_/X _86830_/Q _45976_/X _45978_/X sky130_fd_sc_hd__a2bb2o_4
X_76798_ _76784_/Y _76785_/Y _81488_/Q _81360_/D _76798_/X sky130_fd_sc_hd__a2bb2o_4
X_47717_ _54898_/B _53205_/B sky130_fd_sc_hd__buf_2
X_66551_ _64706_/A _69183_/A sky130_fd_sc_hd__buf_2
X_78537_ _78533_/X _78536_/X _78561_/B sky130_fd_sc_hd__xor2_4
X_44929_ _85183_/Q _44882_/X _44884_/X _44929_/X sky130_fd_sc_hd__o21a_4
X_75749_ _80918_/Q _75751_/A sky130_fd_sc_hd__inv_2
X_63763_ _63733_/X _64184_/C sky130_fd_sc_hd__buf_2
X_60975_ _64191_/D _61012_/A sky130_fd_sc_hd__buf_2
X_48697_ _48697_/A _48697_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_9_120_0_CLK clkbuf_8_60_0_CLK/X clkbuf_9_120_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_65502_ _65438_/X _86204_/Q _65182_/X _65501_/X _65502_/X sky130_fd_sc_hd__a211o_4
X_62714_ _60362_/A _62727_/A sky130_fd_sc_hd__buf_2
X_69270_ _81400_/D _69230_/X _69269_/X _83936_/D sky130_fd_sc_hd__a21bo_4
X_47648_ _54859_/B _53167_/B sky130_fd_sc_hd__buf_2
X_66482_ _66475_/X _66244_/Y _66481_/Y _66482_/Y sky130_fd_sc_hd__o21ai_4
X_78468_ _78475_/A _78467_/Y _82765_/D sky130_fd_sc_hd__xnor2_4
X_63694_ _63484_/A _63694_/B _63672_/C _60682_/A _63694_/X sky130_fd_sc_hd__and4_4
X_68221_ _68097_/A _68221_/X sky130_fd_sc_hd__buf_2
X_65433_ _65399_/X _65431_/Y _65432_/Y _65433_/Y sky130_fd_sc_hd__o21ai_4
X_77419_ _77403_/B _77417_/X _77418_/X _77419_/Y sky130_fd_sc_hd__a21boi_4
X_62645_ _60271_/X _62646_/B sky130_fd_sc_hd__buf_2
X_47579_ _47595_/A _47595_/B _47595_/C _53129_/D _47579_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_644_0_CLK clkbuf_9_322_0_CLK/X _86935_/CLK sky130_fd_sc_hd__clkbuf_1
X_78399_ _78397_/Y _78369_/B _78398_/X _78400_/B sky130_fd_sc_hd__o21ai_4
X_49318_ _52533_/A _49317_/X _49312_/C _49318_/X sky130_fd_sc_hd__and3_4
X_80430_ _80423_/A _80423_/B _80430_/Y sky130_fd_sc_hd__nand2_4
X_68152_ _66965_/X _66967_/X _68129_/X _68152_/Y sky130_fd_sc_hd__a21oi_4
X_65364_ _65285_/A _86020_/Q _65364_/X sky130_fd_sc_hd__and2_4
X_50590_ _50575_/A _48944_/B _50590_/Y sky130_fd_sc_hd__nand2_4
X_62576_ _62556_/A _61640_/A _62576_/C _62548_/D _62576_/X sky130_fd_sc_hd__and4_4
Xclkbuf_9_135_0_CLK clkbuf_8_67_0_CLK/X clkbuf_9_135_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_67103_ _66625_/A _67131_/A sky130_fd_sc_hd__buf_2
X_64315_ _64315_/A _64316_/B sky130_fd_sc_hd__buf_2
Xclkbuf_9_62_0_CLK clkbuf_9_63_0_CLK/A clkbuf_9_62_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_49249_ _49263_/A _53983_/B _49249_/Y sky130_fd_sc_hd__nand2_4
X_61527_ _61340_/A _61542_/C sky130_fd_sc_hd__buf_2
X_80361_ _80361_/A _80361_/B _80362_/A sky130_fd_sc_hd__and2_4
X_68083_ _68371_/A _88148_/Q _68083_/X sky130_fd_sc_hd__and2_4
X_65295_ _65292_/Y _65195_/X _65294_/X _84207_/D sky130_fd_sc_hd__a21o_4
X_82100_ _82349_/CLK _77488_/B _82100_/Q sky130_fd_sc_hd__dfxtp_4
X_67034_ _87936_/Q _66935_/X _67032_/X _67033_/X _67034_/X sky130_fd_sc_hd__a211o_4
X_52260_ _85857_/Q _52239_/X _52259_/Y _52260_/Y sky130_fd_sc_hd__o21ai_4
X_64246_ _64223_/A _64246_/B _64223_/C _64246_/X sky130_fd_sc_hd__and3_4
X_83080_ _86525_/CLK _74372_/Y _83080_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_659_0_CLK clkbuf_9_329_0_CLK/X _87421_/CLK sky130_fd_sc_hd__clkbuf_1
X_80292_ _80292_/A _80292_/B _80296_/A sky130_fd_sc_hd__nand2_4
X_61458_ _61302_/A _72561_/C sky130_fd_sc_hd__buf_2
X_51211_ _51211_/A _51212_/A sky130_fd_sc_hd__buf_2
X_82031_ _81985_/CLK _77850_/B _81999_/D sky130_fd_sc_hd__dfxtp_4
X_60409_ _60408_/X _60482_/A sky130_fd_sc_hd__buf_2
X_52191_ _85871_/Q _52178_/X _52190_/Y _52191_/Y sky130_fd_sc_hd__o21ai_4
X_64177_ _61685_/A _64177_/B _64189_/D _64177_/D _64181_/A sky130_fd_sc_hd__nand4_4
X_61389_ _72550_/C _61390_/D sky130_fd_sc_hd__buf_2
Xclkbuf_9_77_0_CLK clkbuf_8_38_0_CLK/X clkbuf_9_77_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_51142_ _51160_/A _51121_/B _51141_/X _52835_/D _51142_/X sky130_fd_sc_hd__and4_4
X_63128_ _63126_/Y _63127_/X _63114_/X _63128_/Y sky130_fd_sc_hd__a21oi_4
X_68985_ _87078_/Q _68818_/X _68819_/X _68984_/X _68985_/X sky130_fd_sc_hd__a211o_4
X_51073_ _51101_/A _51073_/X sky130_fd_sc_hd__buf_2
X_67936_ _68028_/A _87706_/Q _67936_/X sky130_fd_sc_hd__and2_4
X_55950_ _85213_/Q _55641_/A _55610_/X _55949_/X _55950_/X sky130_fd_sc_hd__a211o_4
X_63059_ _60523_/A _63059_/X sky130_fd_sc_hd__buf_2
X_86770_ _86770_/CLK _46158_/Y _86770_/Q sky130_fd_sc_hd__dfxtp_4
X_83982_ _82629_/CLK _83982_/D _83982_/Q sky130_fd_sc_hd__dfxtp_4
X_50024_ _72427_/B _50012_/X _50023_/Y _50024_/Y sky130_fd_sc_hd__o21ai_4
X_54901_ _54910_/A _54910_/B _54910_/C _53207_/D _54901_/X sky130_fd_sc_hd__and4_4
X_85721_ _84746_/CLK _52972_/Y _85721_/Q sky130_fd_sc_hd__dfxtp_4
X_82933_ _82933_/CLK _78270_/X _46389_/A sky130_fd_sc_hd__dfxtp_4
X_55881_ _55881_/A _55880_/X _55882_/A sky130_fd_sc_hd__and2_4
X_67867_ _87901_/Q _67770_/X _67865_/X _67866_/X _67867_/X sky130_fd_sc_hd__a211o_4
X_57620_ _57618_/Y _57592_/X _57619_/X _57620_/Y sky130_fd_sc_hd__a21oi_4
X_69606_ _87568_/Q _69368_/X _68552_/X _69605_/X _69606_/X sky130_fd_sc_hd__a211o_4
X_54832_ _54828_/Y _54830_/X _54831_/X _85370_/D sky130_fd_sc_hd__a21oi_4
X_66818_ _87945_/Q _66816_/X _66794_/X _66817_/X _66818_/X sky130_fd_sc_hd__a211o_4
X_85652_ _85651_/CLK _85652_/D _85652_/Q sky130_fd_sc_hd__dfxtp_4
X_82864_ _82859_/CLK _78174_/B _82864_/Q sky130_fd_sc_hd__dfxtp_4
X_67798_ _68389_/A _68429_/A sky130_fd_sc_hd__buf_2
X_84603_ _84603_/CLK _60544_/X _79143_/A sky130_fd_sc_hd__dfxtp_4
X_57551_ _46290_/A _72017_/A sky130_fd_sc_hd__buf_2
X_81815_ _81304_/CLK _81815_/D _81815_/Q sky130_fd_sc_hd__dfxtp_4
X_69537_ _87010_/Q _69414_/X _69430_/X _69536_/X _69537_/X sky130_fd_sc_hd__a211o_4
X_88371_ _87859_/CLK _88371_/D _88371_/Q sky130_fd_sc_hd__dfxtp_4
X_54763_ _54758_/X _47481_/A _54763_/Y sky130_fd_sc_hd__nand2_4
X_66749_ _87436_/Q _66678_/X _66747_/X _66748_/X _66749_/X sky130_fd_sc_hd__a211o_4
X_85583_ _86193_/CLK _53712_/Y _85583_/Q sky130_fd_sc_hd__dfxtp_4
X_51975_ _51961_/X _47924_/B _51975_/Y sky130_fd_sc_hd__nand2_4
X_82795_ _82797_/CLK _82827_/Q _78434_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_15_0_CLK clkbuf_8_7_0_CLK/X clkbuf_9_15_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_56502_ _56074_/X _56499_/X _56501_/Y _56502_/Y sky130_fd_sc_hd__o21ai_4
X_87322_ _87577_/CLK _87322_/D _74145_/A sky130_fd_sc_hd__dfxtp_4
X_53714_ _85582_/Q _53687_/X _53713_/Y _53714_/Y sky130_fd_sc_hd__o21ai_4
X_84534_ _84534_/CLK _84534_/D _84534_/Q sky130_fd_sc_hd__dfxtp_4
X_50926_ _50932_/A _51791_/B _50926_/Y sky130_fd_sc_hd__nand2_4
X_57482_ _56910_/X _57400_/X _56915_/Y _57485_/A sky130_fd_sc_hd__nand3_4
X_69468_ _64713_/A _69468_/X sky130_fd_sc_hd__buf_2
X_81746_ _81746_/CLK _76040_/B _81746_/Q sky130_fd_sc_hd__dfxtp_4
X_54694_ _54693_/X _54694_/X sky130_fd_sc_hd__buf_2
X_59221_ _59219_/X _85743_/Q _59220_/X _59221_/X sky130_fd_sc_hd__o21a_4
X_56433_ _56431_/A _56433_/B _85195_/Q _56433_/Y sky130_fd_sc_hd__nand3_4
X_68419_ _73599_/A _68384_/X _68385_/X _68418_/Y _68419_/X sky130_fd_sc_hd__a211o_4
X_87253_ _87253_/CLK _87253_/D _69544_/B sky130_fd_sc_hd__dfxtp_4
X_53645_ _53778_/A _52123_/B _53645_/Y sky130_fd_sc_hd__nand2_4
X_84465_ _84469_/CLK _61625_/Y _79133_/B sky130_fd_sc_hd__dfxtp_4
X_50857_ _50505_/A _50857_/X sky130_fd_sc_hd__buf_2
X_81677_ _81260_/CLK _80045_/X _81677_/Q sky130_fd_sc_hd__dfxtp_4
X_69399_ _57716_/A _69399_/X sky130_fd_sc_hd__buf_2
X_86204_ _85884_/CLK _50422_/Y _86204_/Q sky130_fd_sc_hd__dfxtp_4
X_40610_ _40610_/A _40610_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_3_0_CLK clkbuf_9_3_0_CLK/A clkbuf_9_3_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_59152_ _58864_/A _59152_/X sky130_fd_sc_hd__buf_2
X_71430_ _71432_/A _71432_/B _70778_/A _71432_/D _71430_/X sky130_fd_sc_hd__and4_4
X_83416_ _83415_/CLK _83416_/D _83416_/Q sky130_fd_sc_hd__dfxtp_4
X_56364_ _56164_/X _56284_/X _56363_/Y _85220_/D sky130_fd_sc_hd__o21ai_4
X_80628_ _80613_/X _80614_/X _80627_/Y _80629_/B sky130_fd_sc_hd__a21boi_4
X_41590_ _40518_/B _41624_/B _41590_/X sky130_fd_sc_hd__or2_4
X_87184_ _83753_/CLK _87184_/D _43957_/B sky130_fd_sc_hd__dfxtp_4
X_53576_ _53573_/Y _53574_/X _53575_/Y _85610_/D sky130_fd_sc_hd__a21boi_4
X_84396_ _84396_/CLK _62617_/Y _62616_/C sky130_fd_sc_hd__dfxtp_4
X_50788_ _50787_/X _52482_/B _50788_/Y sky130_fd_sc_hd__nand2_4
X_58103_ _58065_/X _85701_/Q _58089_/X _58103_/X sky130_fd_sc_hd__o21a_4
X_55315_ _45681_/A _55311_/X _55312_/X _55314_/X _55315_/X sky130_fd_sc_hd__a211o_4
X_86135_ _85527_/CLK _50780_/Y _86135_/Q sky130_fd_sc_hd__dfxtp_4
X_40541_ _40463_/X _81155_/Q _40540_/X _40541_/Y sky130_fd_sc_hd__o21ai_4
X_52527_ _65144_/B _52516_/X _52526_/Y _52527_/Y sky130_fd_sc_hd__o21ai_4
X_59083_ _58858_/X _85434_/Q _59082_/X _59083_/Y sky130_fd_sc_hd__o21ai_4
X_71361_ _71366_/A _71351_/X _70782_/A _71363_/D _71361_/X sky130_fd_sc_hd__and4_4
X_83347_ _83763_/CLK _83347_/D _83347_/Q sky130_fd_sc_hd__dfxtp_4
X_56295_ _56350_/A _56296_/A sky130_fd_sc_hd__buf_2
X_80559_ _80559_/A _80559_/B _80560_/B sky130_fd_sc_hd__xor2_4
X_73100_ _73101_/B _73101_/C _73099_/X _73100_/X sky130_fd_sc_hd__a21o_4
X_58034_ _57939_/X _85995_/Q _58033_/X _58034_/Y sky130_fd_sc_hd__o21ai_4
X_70312_ _70249_/X _70328_/D sky130_fd_sc_hd__buf_2
X_43260_ _43162_/A _43260_/X sky130_fd_sc_hd__buf_2
X_55246_ _55276_/A _57199_/A _55246_/X sky130_fd_sc_hd__and2_4
X_86066_ _85748_/CLK _86066_/D _86066_/Q sky130_fd_sc_hd__dfxtp_4
X_74080_ _73378_/A _74080_/X sky130_fd_sc_hd__buf_2
X_40472_ _82320_/Q _40471_/X _40472_/X sky130_fd_sc_hd__or2_4
X_52458_ _52436_/A _53978_/B _52458_/Y sky130_fd_sc_hd__nand2_4
X_83278_ _83278_/CLK _83278_/D _83278_/Q sky130_fd_sc_hd__dfxtp_4
X_71292_ _71291_/Y _71308_/A sky130_fd_sc_hd__buf_2
X_42211_ _41328_/X _42209_/X _87979_/Q _42210_/X _42211_/X sky130_fd_sc_hd__a2bb2o_4
X_85017_ _85049_/CLK _85017_/D _57397_/B sky130_fd_sc_hd__dfxtp_4
X_73031_ _45896_/X _73031_/X sky130_fd_sc_hd__buf_2
X_51409_ _86015_/Q _51402_/X _51408_/Y _51409_/Y sky130_fd_sc_hd__o21ai_4
X_70243_ _70239_/A _70239_/B _83184_/Q _70239_/D _70243_/X sky130_fd_sc_hd__and4_4
X_82229_ _81839_/CLK _82261_/Q _82229_/Q sky130_fd_sc_hd__dfxtp_4
X_43191_ _43047_/X _53944_/A _40899_/X _43190_/Y _43142_/X _87546_/D
+ sky130_fd_sc_hd__o32ai_4
X_55177_ _55177_/A _55176_/Y _55177_/Y sky130_fd_sc_hd__nor2_4
X_52389_ _52618_/A _52496_/A sky130_fd_sc_hd__buf_2
X_42142_ _42096_/A _42142_/X sky130_fd_sc_hd__buf_2
X_54128_ _54127_/X _54123_/B _54118_/X _52963_/D _54128_/X sky130_fd_sc_hd__and4_4
X_70174_ _70134_/X _70233_/A sky130_fd_sc_hd__buf_2
X_59985_ _59985_/A _59985_/X sky130_fd_sc_hd__buf_2
X_46950_ _46903_/A _46981_/C sky130_fd_sc_hd__buf_2
X_42073_ _41912_/A _42073_/X sky130_fd_sc_hd__buf_2
X_58936_ _58858_/X _85444_/Q _58935_/X _58936_/Y sky130_fd_sc_hd__o21ai_4
X_54059_ _85513_/Q _54018_/X _54058_/Y _54059_/Y sky130_fd_sc_hd__o21ai_4
X_77770_ _77780_/B _81927_/D _77773_/A sky130_fd_sc_hd__xnor2_4
X_74982_ _81140_/D _74989_/C _74982_/Y sky130_fd_sc_hd__nand2_4
X_86968_ _87188_/CLK _44762_/Y _86968_/Q sky130_fd_sc_hd__dfxtp_4
X_45901_ _45884_/Y _45898_/X _46159_/A _45900_/Y _45901_/X sky130_fd_sc_hd__a211o_4
X_41024_ _40931_/A _41024_/X sky130_fd_sc_hd__buf_2
X_76721_ _76707_/X _76708_/A _76721_/X sky130_fd_sc_hd__and2_4
X_73933_ _73933_/A _73932_/X _73933_/Y sky130_fd_sc_hd__nand2_4
X_85919_ _85920_/CLK _51942_/Y _65932_/B sky130_fd_sc_hd__dfxtp_4
X_46881_ _58921_/A _46859_/X _46880_/Y _46881_/Y sky130_fd_sc_hd__o21ai_4
X_58867_ _58867_/A _59090_/B _58867_/Y sky130_fd_sc_hd__nor2_4
X_86899_ _80664_/CLK _86899_/D _64353_/B sky130_fd_sc_hd__dfxtp_4
X_48620_ _48563_/X _48077_/A _48619_/Y _48621_/A sky130_fd_sc_hd__o21ai_4
X_79440_ _79416_/A _79416_/B _79429_/A _79428_/Y _79440_/X sky130_fd_sc_hd__o22a_4
X_57818_ _84948_/Q _57691_/X _57810_/X _57817_/X _84948_/D sky130_fd_sc_hd__a2bb2oi_4
X_45832_ _45832_/A _45832_/B _45832_/Y sky130_fd_sc_hd__nand2_4
X_76652_ _81682_/Q _76652_/Y sky130_fd_sc_hd__inv_2
X_73864_ _73864_/A _73864_/B _73864_/X sky130_fd_sc_hd__xor2_4
X_58798_ _58796_/X _86095_/Q _58797_/X _58798_/Y sky130_fd_sc_hd__o21ai_4
X_75603_ _75600_/X _75602_/Y _75604_/B sky130_fd_sc_hd__xor2_4
X_48551_ _48550_/Y _48551_/X sky130_fd_sc_hd__buf_2
X_72815_ _73306_/A _73516_/A sky130_fd_sc_hd__buf_2
X_79371_ _84804_/Q _66433_/C _79373_/A sky130_fd_sc_hd__xor2_4
X_45763_ _62083_/D _61611_/A sky130_fd_sc_hd__buf_2
X_57749_ _57739_/X _85726_/Q _44252_/X _57749_/X sky130_fd_sc_hd__o21a_4
X_76583_ _76583_/A _76583_/Y sky130_fd_sc_hd__inv_2
X_42975_ _42975_/A _42975_/Y sky130_fd_sc_hd__inv_2
X_73795_ _73795_/A _73624_/X _73795_/Y sky130_fd_sc_hd__nor2_4
X_47502_ _47502_/A _53084_/D sky130_fd_sc_hd__buf_2
X_78322_ _78320_/Y _82786_/Q _78321_/Y _78324_/B sky130_fd_sc_hd__a21bo_4
X_44714_ _44714_/A _44714_/X sky130_fd_sc_hd__buf_2
X_75534_ _75533_/Y _75535_/B sky130_fd_sc_hd__inv_2
X_41926_ _41878_/A _42024_/A sky130_fd_sc_hd__buf_2
X_60760_ _60715_/X _60761_/B sky130_fd_sc_hd__buf_2
X_48482_ _48515_/A _48482_/B _48482_/Y sky130_fd_sc_hd__nand2_4
X_72746_ _73351_/A _72746_/X sky130_fd_sc_hd__buf_2
X_45694_ _45690_/X _45693_/Y _45678_/X _45694_/X sky130_fd_sc_hd__a21o_4
X_47433_ _47444_/A _53046_/B _47433_/Y sky130_fd_sc_hd__nand2_4
X_59419_ _59419_/A _59421_/A sky130_fd_sc_hd__buf_2
X_78253_ _78241_/X _78253_/B _82496_/Q _78254_/A sky130_fd_sc_hd__nand3_4
X_44645_ _41050_/A _44618_/X _87019_/Q _44619_/X _44645_/X sky130_fd_sc_hd__a2bb2o_4
X_75465_ _75506_/C _75465_/Y sky130_fd_sc_hd__inv_2
X_41857_ _40538_/X _41847_/X _88118_/Q _41848_/X _88118_/D sky130_fd_sc_hd__a2bb2o_4
X_60691_ _60690_/X _60727_/A sky130_fd_sc_hd__inv_2
X_72677_ _72683_/A _72683_/B _55360_/X _72677_/Y sky130_fd_sc_hd__nand3_4
X_77204_ _77202_/B _82012_/Q _82300_/D _77204_/Y sky130_fd_sc_hd__nand3_4
X_62430_ _62501_/A _62490_/C sky130_fd_sc_hd__buf_2
X_74416_ _74416_/A _74395_/X _74421_/C _74416_/X sky130_fd_sc_hd__and3_4
X_40808_ _82872_/Q _40779_/B _40808_/X sky130_fd_sc_hd__or2_4
X_47364_ _47414_/A _47364_/X sky130_fd_sc_hd__buf_2
X_71628_ _71628_/A _71628_/X sky130_fd_sc_hd__buf_2
X_78184_ _78183_/A _82489_/Q _78191_/C sky130_fd_sc_hd__nand2_4
X_44576_ _44575_/Y _44576_/Y sky130_fd_sc_hd__inv_2
X_75396_ _75396_/A _75393_/Y _75396_/C _75401_/A sky130_fd_sc_hd__or3_4
X_41788_ _41788_/A _41788_/Y sky130_fd_sc_hd__inv_2
X_49103_ _49096_/Y _49086_/X _49102_/X _86444_/D sky130_fd_sc_hd__a21oi_4
X_46315_ _46421_/A _51261_/B _46315_/Y sky130_fd_sc_hd__nand2_4
X_77135_ _77141_/B _77141_/C _77135_/Y sky130_fd_sc_hd__nand2_4
X_43527_ _40391_/X _43513_/X _87375_/Q _43514_/X _87375_/D sky130_fd_sc_hd__a2bb2o_4
X_62361_ _61448_/X _62420_/B _62233_/C _62334_/D _62361_/Y sky130_fd_sc_hd__nand4_4
X_74347_ _74351_/A _74342_/X _55773_/D _74347_/Y sky130_fd_sc_hd__nand3_4
X_40739_ _40739_/A _40739_/X sky130_fd_sc_hd__buf_2
X_47295_ _47330_/A _47311_/B _47321_/C _52967_/D _47295_/X sky130_fd_sc_hd__and4_4
X_71559_ _70670_/A _71553_/B _71558_/X _71559_/Y sky130_fd_sc_hd__nor3_4
X_64100_ _64116_/A _64087_/X _64100_/C _64100_/Y sky130_fd_sc_hd__nor3_4
X_49034_ _83610_/Q _53856_/B sky130_fd_sc_hd__inv_2
X_61312_ _61312_/A _61313_/A sky130_fd_sc_hd__buf_2
X_46246_ _86753_/Q _44736_/X _46245_/X _46247_/A sky130_fd_sc_hd__o21ai_4
XPHY_580 sky130_fd_sc_hd__decap_3
X_65080_ _44150_/X _86735_/Q _64980_/X _65079_/X _65080_/X sky130_fd_sc_hd__a211o_4
X_77066_ _77066_/A _82284_/D _77073_/A sky130_fd_sc_hd__xor2_4
X_43458_ _43458_/A _43458_/Y sky130_fd_sc_hd__inv_2
X_62292_ _60084_/A _62631_/D sky130_fd_sc_hd__buf_2
X_74278_ _74278_/A _74278_/B _74278_/Y sky130_fd_sc_hd__nand2_4
XPHY_591 sky130_fd_sc_hd__decap_3
X_64031_ _64025_/Y _64027_/Y _64029_/Y _64030_/Y _64031_/X sky130_fd_sc_hd__and4_4
X_76017_ _81712_/D _76036_/C _76024_/A sky130_fd_sc_hd__xor2_4
X_42409_ _42408_/Y _87877_/D sky130_fd_sc_hd__inv_2
X_61243_ _61097_/X _64456_/C _61117_/X _61243_/Y sky130_fd_sc_hd__o21ai_4
X_73229_ _69808_/B _57377_/X _73055_/X _73228_/Y _73229_/X sky130_fd_sc_hd__a211o_4
X_46177_ _66517_/B _72527_/A sky130_fd_sc_hd__buf_2
X_43389_ _41437_/X _43386_/X _87447_/Q _43388_/X _43389_/X sky130_fd_sc_hd__a2bb2o_4
X_45128_ _64378_/B _61499_/B sky130_fd_sc_hd__buf_2
X_61174_ _61165_/A _61165_/B _61174_/C _61174_/Y sky130_fd_sc_hd__nor3_4
X_60125_ _60125_/A _60214_/B _84658_/Q _60125_/Y sky130_fd_sc_hd__nor3_4
X_49936_ _49955_/A _53148_/B _49936_/Y sky130_fd_sc_hd__nand2_4
X_45059_ _80670_/Q _45284_/A sky130_fd_sc_hd__buf_2
X_68770_ _69178_/A _68770_/X sky130_fd_sc_hd__buf_2
X_65982_ _65824_/X _84988_/Q _65707_/X _65981_/X _65982_/X sky130_fd_sc_hd__a211o_4
X_77968_ _77980_/A _77967_/Y _77968_/X sky130_fd_sc_hd__and2_4
X_67721_ _67715_/X _67720_/X _67619_/X _67726_/A sky130_fd_sc_hd__a21o_4
X_79707_ _79694_/X _79705_/X _79706_/X _79707_/Y sky130_fd_sc_hd__a21oi_4
X_64933_ _64930_/X _64932_/X _64807_/X _64933_/X sky130_fd_sc_hd__a21o_4
X_60056_ _60056_/A _60059_/B sky130_fd_sc_hd__inv_2
X_76919_ _76931_/B _76919_/Y sky130_fd_sc_hd__inv_2
X_49867_ _49865_/Y _49844_/X _49866_/X _49867_/Y sky130_fd_sc_hd__a21oi_4
X_77899_ _82069_/Q _77899_/Y sky130_fd_sc_hd__inv_2
X_48818_ _52204_/A _48829_/B _48814_/C _48818_/X sky130_fd_sc_hd__and3_4
X_79638_ _79636_/X _79646_/B _79638_/Y sky130_fd_sc_hd__xnor2_4
X_67652_ _67675_/A _67652_/B _67652_/X sky130_fd_sc_hd__and2_4
X_64864_ _64991_/A _64864_/X sky130_fd_sc_hd__buf_2
X_49798_ _49825_/A _49798_/X sky130_fd_sc_hd__buf_2
X_66603_ _87378_/Q _66571_/X _66574_/X _66602_/X _66603_/X sky130_fd_sc_hd__a211o_4
X_63815_ _63765_/A _64257_/A _63765_/C _63815_/X sky130_fd_sc_hd__and3_4
X_48749_ _48747_/Y _48734_/X _48748_/X _48749_/Y sky130_fd_sc_hd__a21oi_4
X_67583_ _87465_/Q _67512_/X _67581_/X _67582_/X _67583_/X sky130_fd_sc_hd__a211o_4
X_79569_ _79569_/A _79569_/B _79569_/Y sky130_fd_sc_hd__nand2_4
X_64795_ _64615_/X _85530_/Q _64642_/X _64794_/X _64795_/X sky130_fd_sc_hd__a211o_4
X_81600_ _81473_/CLK _65449_/C _76942_/B sky130_fd_sc_hd__dfxtp_4
X_69322_ _69322_/A _88294_/Q _69322_/X sky130_fd_sc_hd__and2_4
X_66534_ _66534_/A _69633_/A sky130_fd_sc_hd__buf_2
X_51760_ _51814_/A _51782_/B sky130_fd_sc_hd__buf_2
X_63746_ _63743_/X _63744_/X _63745_/Y _84297_/D sky130_fd_sc_hd__a21oi_4
X_82580_ _82580_/CLK _82612_/Q _78203_/A sky130_fd_sc_hd__dfxtp_4
X_60958_ _60953_/X _60954_/X _60957_/Y _60958_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_10_583_0_CLK clkbuf_9_291_0_CLK/X _80931_/CLK sky130_fd_sc_hd__clkbuf_1
X_50711_ _50709_/Y _50699_/X _50710_/Y _86149_/D sky130_fd_sc_hd__a21boi_4
X_81531_ _81703_/CLK _76522_/B _81531_/Q sky130_fd_sc_hd__dfxtp_4
X_69253_ _69253_/A _88299_/Q _69253_/X sky130_fd_sc_hd__and2_4
X_66465_ _66463_/Y _66449_/X _66464_/X _84118_/D sky130_fd_sc_hd__a21o_4
X_51691_ _51697_/A _53213_/B _51691_/Y sky130_fd_sc_hd__nand2_4
X_63677_ _61656_/A _63600_/X _63661_/C _63661_/D _63677_/Y sky130_fd_sc_hd__nand4_4
X_60889_ _60879_/D _60889_/X sky130_fd_sc_hd__buf_2
X_68204_ _67277_/X _67280_/X _68173_/X _68204_/Y sky130_fd_sc_hd__a21oi_4
X_53430_ _53427_/Y _53408_/X _53429_/X _85635_/D sky130_fd_sc_hd__a21oi_4
X_65416_ _65782_/A _65416_/X sky130_fd_sc_hd__buf_2
X_84250_ _84250_/CLK _64398_/X _79722_/B sky130_fd_sc_hd__dfxtp_4
X_50642_ _50627_/X _50133_/B _50642_/Y sky130_fd_sc_hd__nand2_4
X_62628_ _62269_/X _84906_/Q _62628_/C _62219_/X _62628_/X sky130_fd_sc_hd__and4_4
X_81462_ _81482_/CLK _76838_/B _81462_/Q sky130_fd_sc_hd__dfxtp_4
X_69184_ _69027_/A _88304_/Q _69184_/X sky130_fd_sc_hd__and2_4
X_66396_ _66393_/Y _66377_/X _66395_/Y _84131_/D sky130_fd_sc_hd__a21o_4
X_83201_ _83835_/CLK _83201_/D _83201_/Q sky130_fd_sc_hd__dfxtp_4
X_80413_ _80413_/A _80413_/B _80413_/X sky130_fd_sc_hd__xor2_4
X_68135_ _68121_/X _66837_/Y _68128_/X _68134_/Y _68135_/X sky130_fd_sc_hd__a211o_4
X_53361_ _85648_/Q _53351_/X _53360_/Y _53361_/Y sky130_fd_sc_hd__o21ai_4
X_65347_ _65529_/A _65347_/X sky130_fd_sc_hd__buf_2
X_84181_ _83508_/CLK _65746_/X _84181_/Q sky130_fd_sc_hd__dfxtp_4
X_50573_ _50580_/A _71970_/B _50573_/Y sky130_fd_sc_hd__nand2_4
X_81393_ _81351_/CLK _81393_/D _76949_/B sky130_fd_sc_hd__dfxtp_4
X_62559_ _60056_/A _62097_/X _59936_/X _58184_/A _62559_/Y sky130_fd_sc_hd__a22oi_4
Xclkbuf_10_598_0_CLK clkbuf_9_299_0_CLK/X _83906_/CLK sky130_fd_sc_hd__clkbuf_1
X_55100_ _55118_/A _47780_/A _55100_/Y sky130_fd_sc_hd__nand2_4
X_52312_ _52299_/A _48982_/X _52312_/Y sky130_fd_sc_hd__nand2_4
X_83132_ _83133_/CLK _83132_/D _83132_/Q sky130_fd_sc_hd__dfxtp_4
X_56080_ _56100_/A _56086_/B _56080_/C _56080_/Y sky130_fd_sc_hd__nand3_4
X_80344_ _84751_/Q _84143_/Q _80344_/X sky130_fd_sc_hd__or2_4
X_68066_ _69747_/A _68066_/X sky130_fd_sc_hd__buf_2
X_53292_ _51843_/A _53293_/B sky130_fd_sc_hd__buf_2
X_65278_ _65271_/X _65276_/X _65277_/X _65281_/A sky130_fd_sc_hd__a21o_4
X_55031_ _55017_/X _55030_/X _55026_/C _55031_/D _55031_/X sky130_fd_sc_hd__and4_4
X_67017_ _66947_/X _67005_/Y _66910_/X _67016_/Y _67017_/X sky130_fd_sc_hd__a211o_4
X_52243_ _48680_/A _52248_/B _52223_/C _52243_/X sky130_fd_sc_hd__and3_4
X_64229_ _64440_/A _64229_/X sky130_fd_sc_hd__buf_2
X_83063_ _85581_/CLK _83063_/D _83063_/Q sky130_fd_sc_hd__dfxtp_4
X_87940_ _88386_/CLK _42285_/Y _87940_/Q sky130_fd_sc_hd__dfxtp_4
X_80275_ _80273_/Y _80274_/Y _80275_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_521_0_CLK clkbuf_9_260_0_CLK/X _81431_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_12_0_CLK clkbuf_5_6_0_CLK/X clkbuf_6_12_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_82014_ _82139_/CLK _82046_/Q _77200_/A sky130_fd_sc_hd__dfxtp_4
X_52174_ _85874_/Q _52152_/X _52173_/Y _52174_/Y sky130_fd_sc_hd__o21ai_4
X_87871_ _82888_/CLK _87871_/D _87871_/Q sky130_fd_sc_hd__dfxtp_4
X_51125_ _51115_/A _51121_/B _51115_/C _52818_/D _51125_/X sky130_fd_sc_hd__and4_4
X_86822_ _87077_/CLK _45998_/X _86822_/Q sky130_fd_sc_hd__dfxtp_4
X_59770_ _59770_/A _65044_/A sky130_fd_sc_hd__buf_2
X_56982_ _57019_/A _56982_/X sky130_fd_sc_hd__buf_2
X_68968_ _87483_/Q _68870_/X _68871_/X _68967_/X _68968_/X sky130_fd_sc_hd__a211o_4
X_58721_ _58721_/A _58764_/B sky130_fd_sc_hd__buf_2
X_51056_ _51056_/A _51045_/B _51045_/C _52746_/D _51056_/X sky130_fd_sc_hd__and4_4
X_55933_ _55930_/X _55932_/X _55615_/A _55936_/A sky130_fd_sc_hd__a21o_4
X_67919_ _67992_/A _88155_/Q _67919_/X sky130_fd_sc_hd__and2_4
X_86753_ _86753_/CLK _46247_/Y _86753_/Q sky130_fd_sc_hd__dfxtp_4
X_83965_ _83967_/CLK _68690_/X _80821_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_536_0_CLK clkbuf_9_268_0_CLK/X _81412_/CLK sky130_fd_sc_hd__clkbuf_1
X_68899_ _87486_/Q _68870_/X _68871_/X _68898_/X _68899_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_6_27_0_CLK clkbuf_6_27_0_CLK/A clkbuf_7_55_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_50007_ _50001_/A _53219_/B _50007_/Y sky130_fd_sc_hd__nand2_4
X_85704_ _85704_/CLK _85704_/D _85704_/Q sky130_fd_sc_hd__dfxtp_4
X_70930_ _70905_/A _70863_/C _70925_/X _70913_/A _70930_/Y sky130_fd_sc_hd__nand4_4
X_58652_ _58639_/Y _58624_/X _58647_/X _58651_/X _84811_/D sky130_fd_sc_hd__a22oi_4
X_82916_ _82368_/CLK _78144_/X _82916_/Q sky130_fd_sc_hd__dfxtp_4
X_55864_ _55830_/X _56083_/C _55854_/X _55863_/X _55864_/X sky130_fd_sc_hd__and4_4
X_86684_ _86686_/CLK _86684_/D _59057_/A sky130_fd_sc_hd__dfxtp_4
X_83896_ _82299_/CLK _83896_/D _81968_/D sky130_fd_sc_hd__dfxtp_4
X_57603_ _46542_/X _57603_/X sky130_fd_sc_hd__buf_2
X_54815_ _85373_/Q _54812_/X _54814_/Y _54815_/Y sky130_fd_sc_hd__o21ai_4
X_85635_ _85635_/CLK _85635_/D _85635_/Q sky130_fd_sc_hd__dfxtp_4
X_70861_ _51791_/B _70855_/X _70860_/Y _70861_/Y sky130_fd_sc_hd__o21ai_4
X_58583_ _58580_/Y _58582_/Y _58105_/X _58583_/X sky130_fd_sc_hd__a21o_4
X_82847_ _82152_/CLK _82847_/D _82847_/Q sky130_fd_sc_hd__dfxtp_4
X_55795_ _85196_/Q _55747_/X _55300_/X _55794_/X _55795_/X sky130_fd_sc_hd__a211o_4
X_72600_ _72576_/A _72535_/A _59829_/X _72600_/Y sky130_fd_sc_hd__a21oi_4
X_57534_ _84984_/Q _57527_/X _57533_/Y _57534_/Y sky130_fd_sc_hd__o21ai_4
X_88354_ _86998_/CLK _88354_/D _88354_/Q sky130_fd_sc_hd__dfxtp_4
X_42760_ _41272_/X _42757_/X _69076_/B _42759_/X _87734_/D sky130_fd_sc_hd__a2bb2o_4
X_54746_ _85385_/Q _54729_/X _54745_/Y _54746_/Y sky130_fd_sc_hd__o21ai_4
X_85566_ _85566_/CLK _53802_/Y _85566_/Q sky130_fd_sc_hd__dfxtp_4
X_73580_ _88370_/Q _72769_/B _73007_/A _73580_/X sky130_fd_sc_hd__o21a_4
X_51958_ _47886_/A _51352_/B _51958_/C _51958_/X sky130_fd_sc_hd__and3_4
X_70792_ _52869_/B _70761_/A _70791_/Y _70792_/Y sky130_fd_sc_hd__o21ai_4
X_82778_ _82206_/CLK _82778_/D _82778_/Q sky130_fd_sc_hd__dfxtp_4
X_87305_ _88327_/CLK _87305_/D _87305_/Q sky130_fd_sc_hd__dfxtp_4
X_41711_ _41672_/X _41673_/X _41710_/X _88164_/Q _41668_/X _41712_/A
+ sky130_fd_sc_hd__o32ai_4
X_84517_ _84498_/CLK _84517_/D _84517_/Q sky130_fd_sc_hd__dfxtp_4
X_72531_ _72597_/B _72535_/B _72597_/C _72531_/Y sky130_fd_sc_hd__nand3_4
X_50909_ _50907_/Y _50902_/X _50908_/X _86109_/D sky130_fd_sc_hd__a21oi_4
X_57465_ _57465_/A _56872_/Y _57465_/X sky130_fd_sc_hd__or2_4
X_81729_ _81346_/CLK _81729_/D _41114_/A sky130_fd_sc_hd__dfxtp_4
X_42691_ _42687_/X _42688_/X _41087_/X _87768_/Q _42673_/X _42692_/A
+ sky130_fd_sc_hd__o32ai_4
X_88285_ _87011_/CLK _41060_/X _88285_/Q sky130_fd_sc_hd__dfxtp_4
X_54677_ _54594_/X _54682_/A sky130_fd_sc_hd__buf_2
X_85497_ _83745_/CLK _54138_/Y _85497_/Q sky130_fd_sc_hd__dfxtp_4
X_51889_ _51875_/A _51026_/B _51889_/Y sky130_fd_sc_hd__nand2_4
X_59204_ _80441_/A _59204_/Y sky130_fd_sc_hd__inv_2
X_44430_ _44430_/A _87113_/D sky130_fd_sc_hd__inv_2
X_56416_ _56418_/A _56418_/B _85202_/Q _56416_/Y sky130_fd_sc_hd__nand3_4
X_75250_ _80782_/Q _75249_/Y _75250_/X sky130_fd_sc_hd__xor2_4
X_41642_ _41588_/X _81759_/Q _41641_/X _41642_/Y sky130_fd_sc_hd__o21ai_4
X_87236_ _87758_/CLK _87236_/D _87236_/Q sky130_fd_sc_hd__dfxtp_4
X_53628_ _53656_/A _74373_/B _53628_/Y sky130_fd_sc_hd__nand2_4
X_72462_ _86596_/Q _72401_/B _72462_/Y sky130_fd_sc_hd__nor2_4
X_84448_ _84449_/CLK _61883_/Y _78071_/B sky130_fd_sc_hd__dfxtp_4
X_57396_ _57394_/X _56607_/X _85018_/Q _57395_/X _85018_/D sky130_fd_sc_hd__a2bb2o_4
X_74201_ _74191_/Y _74201_/B _74201_/Y sky130_fd_sc_hd__xnor2_4
X_71413_ _70689_/A _71411_/B _71411_/C _71413_/Y sky130_fd_sc_hd__nor3_4
X_59135_ _58877_/A _59135_/X sky130_fd_sc_hd__buf_2
X_44361_ _44361_/A _44361_/Y sky130_fd_sc_hd__inv_2
X_56347_ _56347_/A _56358_/A sky130_fd_sc_hd__buf_2
X_87167_ _87417_/CLK _87167_/D _87167_/Q sky130_fd_sc_hd__dfxtp_4
X_75181_ _75167_/B _75162_/A _75162_/B _75181_/Y sky130_fd_sc_hd__a21boi_4
X_41573_ _41533_/X _82315_/Q _41572_/X _41573_/X sky130_fd_sc_hd__o21a_4
X_53559_ _85613_/Q _53556_/X _53558_/Y _53559_/Y sky130_fd_sc_hd__o21ai_4
X_72393_ _83259_/Q _72381_/X _72385_/X _72392_/X _83259_/D sky130_fd_sc_hd__a2bb2oi_4
X_84379_ _84375_/CLK _84379_/D _62825_/C sky130_fd_sc_hd__dfxtp_4
X_46100_ _46111_/A _46099_/X _46094_/X _46101_/A sky130_fd_sc_hd__nor3_4
X_43312_ _43312_/A _87487_/D sky130_fd_sc_hd__inv_2
X_74132_ _73588_/A _66256_/B _74132_/X sky130_fd_sc_hd__and2_4
X_86118_ _86118_/CLK _86118_/D _86118_/Q sky130_fd_sc_hd__dfxtp_4
X_40524_ _40523_/Y _40524_/X sky130_fd_sc_hd__buf_2
X_47080_ _86672_/Q _47050_/X _47079_/Y _47080_/Y sky130_fd_sc_hd__o21ai_4
X_59066_ _59029_/A _86363_/Q _59066_/Y sky130_fd_sc_hd__nor2_4
X_71344_ _71344_/A _71344_/X sky130_fd_sc_hd__buf_2
X_44292_ _44292_/A _72498_/B sky130_fd_sc_hd__buf_2
X_56278_ _56278_/A _57223_/D sky130_fd_sc_hd__buf_2
X_87098_ _87011_/CLK _44461_/Y _87098_/Q sky130_fd_sc_hd__dfxtp_4
X_46031_ _41468_/Y _46029_/X _86804_/Q _46030_/X _46031_/X sky130_fd_sc_hd__a2bb2o_4
X_58017_ _58703_/A _58017_/X sky130_fd_sc_hd__buf_2
X_55229_ _55129_/A _85060_/Q _55229_/X sky130_fd_sc_hd__and2_4
X_43243_ _43243_/A _87521_/D sky130_fd_sc_hd__inv_2
X_74063_ _74022_/X _66214_/B _74063_/X sky130_fd_sc_hd__and2_4
X_78940_ _78940_/A _78942_/A sky130_fd_sc_hd__inv_2
X_86049_ _85535_/CLK _51239_/Y _64572_/B sky130_fd_sc_hd__dfxtp_4
X_40455_ _47825_/A _40783_/A sky130_fd_sc_hd__buf_2
X_71275_ _53193_/B _71265_/X _71274_/Y _83551_/D sky130_fd_sc_hd__o21ai_4
X_73014_ _73011_/X _73013_/X _72812_/X _73018_/A sky130_fd_sc_hd__a21o_4
X_70226_ _70224_/X _83831_/Q _70225_/X _83831_/D sky130_fd_sc_hd__a21o_4
X_43174_ _43174_/A _43174_/Y sky130_fd_sc_hd__inv_2
X_78871_ _82842_/Q _82554_/Q _78896_/A sky130_fd_sc_hd__xnor2_4
X_40386_ _40381_/X _81182_/Q _40385_/X _40386_/Y sky130_fd_sc_hd__o21ai_4
X_42125_ _51719_/A _42125_/X sky130_fd_sc_hd__buf_2
X_77822_ _77822_/A _77822_/B _77822_/Y sky130_fd_sc_hd__nand2_4
X_70157_ _70157_/A _70157_/X sky130_fd_sc_hd__buf_2
X_47982_ _47982_/A _47973_/B _47982_/X sky130_fd_sc_hd__or2_4
X_59968_ _59968_/A _59968_/B _59968_/X sky130_fd_sc_hd__and2_4
X_49721_ _49716_/X _52936_/B _49721_/Y sky130_fd_sc_hd__nand2_4
X_46933_ _54449_/D _52758_/D sky130_fd_sc_hd__buf_2
X_58919_ _58698_/A _58920_/A sky130_fd_sc_hd__buf_2
X_42056_ _42056_/A _42056_/Y sky130_fd_sc_hd__inv_2
X_77753_ _77745_/Y _77753_/B _77754_/B sky130_fd_sc_hd__xor2_4
X_74965_ _80763_/Q _74965_/B _74971_/B sky130_fd_sc_hd__xor2_4
X_70088_ _83853_/Q _70085_/X _70087_/X _70088_/X sky130_fd_sc_hd__a21bo_4
X_59899_ _43969_/A _59899_/B _43969_/B _59899_/D _59899_/X sky130_fd_sc_hd__and4_4
X_41007_ _41007_/A _41007_/B _41007_/X sky130_fd_sc_hd__or2_4
X_76704_ _76698_/Y _76699_/X _76703_/Y _76704_/Y sky130_fd_sc_hd__a21oi_4
X_49652_ _49651_/X _49642_/B _49629_/X _52867_/D _49652_/X sky130_fd_sc_hd__and4_4
X_61930_ _61711_/X _61949_/A sky130_fd_sc_hd__buf_2
X_73916_ _44705_/A _73916_/B _73916_/Y sky130_fd_sc_hd__nor2_4
X_46864_ _86695_/Q _46859_/X _46863_/Y _46864_/Y sky130_fd_sc_hd__o21ai_4
X_77684_ _77662_/Y _77695_/B _77693_/C _77688_/A sky130_fd_sc_hd__o21a_4
X_74896_ _81130_/D _80842_/Q _74905_/A sky130_fd_sc_hd__xor2_4
X_48603_ _48602_/Y _50508_/B sky130_fd_sc_hd__buf_2
X_79423_ _79417_/Y _79422_/Y _82840_/D sky130_fd_sc_hd__xor2_4
X_45815_ _56887_/B _45798_/X _45743_/X _45815_/X sky130_fd_sc_hd__o21a_4
X_76635_ _76635_/A _76634_/Y _76635_/X sky130_fd_sc_hd__xor2_4
X_61861_ _84881_/Q _61861_/X sky130_fd_sc_hd__buf_2
X_49583_ _49571_/X _49561_/B _49577_/C _52797_/D _49583_/X sky130_fd_sc_hd__and4_4
X_73847_ _73843_/X _73846_/X _73799_/X _73866_/B sky130_fd_sc_hd__a21o_4
X_46795_ _52677_/B _50987_/B sky130_fd_sc_hd__buf_2
X_63600_ _63478_/A _63600_/X sky130_fd_sc_hd__buf_2
X_60812_ _60732_/C _60711_/X _60722_/A _60812_/Y sky130_fd_sc_hd__o21ai_4
X_48534_ _48528_/Y _48517_/X _48533_/X _86514_/D sky130_fd_sc_hd__a21oi_4
X_79354_ _79350_/X _79353_/Y _79354_/X sky130_fd_sc_hd__xor2_4
X_45746_ _74679_/B _45746_/B _45746_/Y sky130_fd_sc_hd__nand2_4
X_64580_ _64621_/A _64580_/B _64580_/X sky130_fd_sc_hd__and2_4
X_76566_ _76566_/A _76584_/D _76566_/Y sky130_fd_sc_hd__nand2_4
X_42958_ _40391_/X _42950_/X _66676_/B _42951_/X _87631_/D sky130_fd_sc_hd__a2bb2o_4
X_61792_ _58232_/X _61728_/X _61756_/X _61790_/X _61791_/X _61792_/X
+ sky130_fd_sc_hd__a41o_4
X_73778_ _68595_/B _73777_/X _73656_/X _73778_/X sky130_fd_sc_hd__o21a_4
X_78305_ _78305_/A _78304_/Y _78309_/A sky130_fd_sc_hd__nand2_4
X_63531_ _63527_/Y _63516_/X _63530_/Y _63531_/Y sky130_fd_sc_hd__a21oi_4
X_75517_ _80703_/Q _80959_/D _75517_/Y sky130_fd_sc_hd__nand2_4
X_41909_ _46450_/A _50256_/A _41909_/B1 _41909_/Y sky130_fd_sc_hd__a21oi_4
X_48465_ _50443_/A _48489_/B _48476_/C _48465_/X sky130_fd_sc_hd__and3_4
X_60743_ _60694_/B _60739_/X _63648_/B _60743_/X sky130_fd_sc_hd__o21a_4
X_72729_ _41980_/Y _72723_/X _72725_/X _72728_/Y _72729_/X sky130_fd_sc_hd__a211o_4
X_79285_ _79278_/X _79285_/B _79285_/Y sky130_fd_sc_hd__nand2_4
X_45677_ _85039_/Q _45675_/X _45676_/X _45677_/Y sky130_fd_sc_hd__o21ai_4
X_76497_ _76513_/B _76513_/D _76497_/X sky130_fd_sc_hd__and2_4
X_42889_ _42874_/X _42875_/X _41631_/X _87667_/Q _42881_/X _42889_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47416_ _81805_/Q _47417_/A sky130_fd_sc_hd__inv_2
X_66250_ _66125_/X _86217_/Q _66180_/X _66249_/X _66250_/X sky130_fd_sc_hd__a211o_4
X_78236_ _82583_/Q _82495_/Q _78236_/Y sky130_fd_sc_hd__nand2_4
X_44628_ _44622_/X _44623_/X _41003_/X _87027_/Q _44625_/X _44628_/Y
+ sky130_fd_sc_hd__o32ai_4
X_63462_ _63488_/A _61861_/X _63462_/X sky130_fd_sc_hd__and2_4
X_75448_ _75446_/X _75448_/B _75467_/A sky130_fd_sc_hd__and2_4
X_48396_ _74381_/A _53636_/A sky130_fd_sc_hd__buf_2
X_60674_ _60660_/A _60804_/B sky130_fd_sc_hd__buf_2
X_65201_ _65225_/A _85834_/Q _65201_/X sky130_fd_sc_hd__and2_4
X_62413_ _62411_/X _62412_/X _84412_/Q _62413_/Y sky130_fd_sc_hd__nor3_4
X_47347_ _81812_/Q _47348_/A sky130_fd_sc_hd__inv_2
X_66181_ _66181_/A _85902_/Q _66181_/X sky130_fd_sc_hd__and2_4
X_78167_ _78167_/A _78166_/Y _78168_/B sky130_fd_sc_hd__xor2_4
X_44559_ _44547_/X _44548_/X _40849_/X _87055_/Q _44549_/X _44560_/A
+ sky130_fd_sc_hd__o32ai_4
X_63393_ _63390_/Y _63391_/X _63392_/Y _63393_/Y sky130_fd_sc_hd__a21oi_4
X_75379_ _75375_/Y _75377_/Y _75378_/Y _75383_/B sky130_fd_sc_hd__o21a_4
X_65132_ _65002_/A _86253_/Q _65132_/X sky130_fd_sc_hd__and2_4
X_77118_ _77118_/A _77118_/B _77118_/X sky130_fd_sc_hd__xor2_4
X_62344_ _62269_/A _62344_/X sky130_fd_sc_hd__buf_2
X_47278_ _54125_/B _52959_/B sky130_fd_sc_hd__buf_2
X_78098_ _78087_/Y _78098_/Y sky130_fd_sc_hd__inv_2
X_49017_ _64951_/B _49003_/X _49016_/Y _49017_/Y sky130_fd_sc_hd__o21ai_4
X_46229_ _40335_/B _46091_/Y _46162_/A _46096_/D _46228_/Y _46229_/Y
+ sky130_fd_sc_hd__a41oi_4
X_69940_ _69525_/X _69527_/X _69939_/X _69940_/Y sky130_fd_sc_hd__a21oi_4
X_65063_ _65058_/X _65062_/X _64989_/X _65063_/X sky130_fd_sc_hd__a21o_4
X_77049_ _82089_/Q _77049_/B _77049_/X sky130_fd_sc_hd__xor2_4
X_62275_ _62362_/A _62272_/Y _62273_/Y _62274_/Y _62275_/Y sky130_fd_sc_hd__nand4_4
X_64014_ _60879_/B _64029_/C sky130_fd_sc_hd__buf_2
X_61226_ _64419_/B _61226_/X sky130_fd_sc_hd__buf_2
X_80060_ _84663_/Q _64037_/C _80060_/X sky130_fd_sc_hd__xor2_4
X_69871_ _64615_/A _42604_/Y _69871_/Y sky130_fd_sc_hd__nor2_4
X_68822_ _68817_/X _68821_/X _68822_/Y sky130_fd_sc_hd__nand2_4
X_61157_ _61165_/A _61138_/B _84517_/Q _61157_/Y sky130_fd_sc_hd__nor3_4
X_60108_ _60078_/X _60079_/Y _59962_/A _60100_/Y _60107_/Y _60108_/Y
+ sky130_fd_sc_hd__a41oi_4
X_49919_ _72192_/B _49906_/X _49918_/Y _49919_/Y sky130_fd_sc_hd__o21ai_4
X_68753_ _67816_/A _69233_/A sky130_fd_sc_hd__buf_2
X_65965_ _57770_/A _86557_/Q _65965_/X sky130_fd_sc_hd__and2_4
X_61088_ _65044_/A _61414_/A sky130_fd_sc_hd__buf_2
X_67704_ _87460_/Q _67628_/X _67702_/X _67703_/X _67704_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_4_2_1_CLK clkbuf_4_2_1_CLK/A clkbuf_4_2_1_CLK/X sky130_fd_sc_hd__clkbuf_1
X_52930_ _52903_/X _52944_/A sky130_fd_sc_hd__buf_2
X_64916_ _64767_/A _85813_/Q _64916_/X sky130_fd_sc_hd__and2_4
X_60039_ _59974_/Y _59951_/D _60049_/A sky130_fd_sc_hd__nand2_4
X_83750_ _83753_/CLK _70556_/X _83750_/Q sky130_fd_sc_hd__dfxtp_4
X_80962_ _80962_/CLK _80962_/D _80950_/D sky130_fd_sc_hd__dfxtp_4
X_68684_ _69035_/A _68684_/X sky130_fd_sc_hd__buf_2
X_65896_ _65896_/A _86498_/Q _65896_/X sky130_fd_sc_hd__and2_4
X_82701_ _81190_/CLK _78909_/X _78793_/A sky130_fd_sc_hd__dfxtp_4
X_67635_ _87155_/Q _67585_/X _67633_/X _67634_/X _67635_/X sky130_fd_sc_hd__a211o_4
X_52861_ _52853_/A _52853_/B _52853_/C _52861_/D _52861_/X sky130_fd_sc_hd__and4_4
X_64847_ _64616_/A _64948_/A sky130_fd_sc_hd__buf_2
X_83681_ _83681_/CLK _70861_/Y _83681_/Q sky130_fd_sc_hd__dfxtp_4
X_80893_ _80991_/CLK _75824_/Y _80893_/Q sky130_fd_sc_hd__dfxtp_4
X_54600_ _54600_/A _47195_/A _54600_/Y sky130_fd_sc_hd__nand2_4
X_85420_ _85645_/CLK _54560_/Y _85420_/Q sky130_fd_sc_hd__dfxtp_4
X_51812_ _51796_/A _51812_/B _51812_/Y sky130_fd_sc_hd__nand2_4
X_82632_ _87671_/CLK _82632_/D _78865_/B sky130_fd_sc_hd__dfxtp_4
X_55580_ _55580_/A _55580_/B _55580_/X sky130_fd_sc_hd__and2_4
X_67566_ _67522_/X _67555_/Y _67507_/X _67565_/Y _67566_/X sky130_fd_sc_hd__a211o_4
X_52792_ _52684_/A _52792_/X sky130_fd_sc_hd__buf_2
X_64778_ _64778_/A _85819_/Q _64778_/X sky130_fd_sc_hd__and2_4
X_69305_ _69305_/A _87271_/Q _69305_/X sky130_fd_sc_hd__and2_4
X_54531_ _54509_/A _54526_/B _54509_/C _47074_/A _54531_/X sky130_fd_sc_hd__and4_4
X_66517_ _66338_/X _66517_/B _66340_/X _66517_/Y sky130_fd_sc_hd__nand3_4
X_85351_ _85351_/CLK _85351_/D _85351_/Q sky130_fd_sc_hd__dfxtp_4
X_51743_ _51738_/Y _51719_/X _51742_/X _51743_/Y sky130_fd_sc_hd__a21oi_4
X_63729_ _60930_/C _64190_/D sky130_fd_sc_hd__buf_2
X_82563_ _82563_/CLK _82595_/Q _82563_/Q sky130_fd_sc_hd__dfxtp_4
X_67497_ _67497_/A _87660_/Q _67497_/X sky130_fd_sc_hd__and2_4
XPHY_14 sky130_fd_sc_hd__decap_3
XPHY_25 sky130_fd_sc_hd__decap_3
X_84302_ _84358_/CLK _63681_/Y _80323_/B sky130_fd_sc_hd__dfxtp_4
X_81514_ _81514_/CLK _81514_/D _81514_/Q sky130_fd_sc_hd__dfxtp_4
X_57250_ _56960_/X _85051_/Q _57249_/X _57250_/Y sky130_fd_sc_hd__nor3_4
X_69236_ _69236_/A _69236_/B _69236_/X sky130_fd_sc_hd__and2_4
XPHY_36 sky130_fd_sc_hd__decap_3
X_88070_ _87814_/CLK _42017_/Y _73106_/A sky130_fd_sc_hd__dfxtp_4
X_54462_ _54453_/X _54440_/B _54471_/C _46952_/A _54462_/X sky130_fd_sc_hd__and4_4
X_66448_ _60110_/X _65031_/Y _66447_/Y _66448_/Y sky130_fd_sc_hd__o21ai_4
X_85282_ _82979_/CLK _56178_/Y _55741_/B sky130_fd_sc_hd__dfxtp_4
X_51674_ _51672_/Y _51667_/X _51673_/X _85967_/D sky130_fd_sc_hd__a21oi_4
XPHY_47 sky130_fd_sc_hd__decap_3
X_82494_ _82503_/CLK _82494_/D _78228_/B sky130_fd_sc_hd__dfxtp_4
XPHY_58 sky130_fd_sc_hd__decap_3
XPHY_69 sky130_fd_sc_hd__decap_3
X_56201_ _56200_/X _56192_/B _85278_/Q _56201_/Y sky130_fd_sc_hd__nand3_4
X_87021_ _87026_/CLK _87021_/D _87021_/Q sky130_fd_sc_hd__dfxtp_4
X_53413_ _85638_/Q _53404_/X _53412_/Y _53413_/Y sky130_fd_sc_hd__o21ai_4
X_84233_ _85346_/CLK _64610_/X _84233_/Q sky130_fd_sc_hd__dfxtp_4
X_50625_ _50623_/Y _50619_/X _50624_/Y _86165_/D sky130_fd_sc_hd__a21boi_4
X_57181_ _56814_/A _57153_/B _57180_/Y _85067_/D sky130_fd_sc_hd__a21o_4
X_81445_ _81412_/CLK _81445_/D _81445_/Q sky130_fd_sc_hd__dfxtp_4
X_69167_ _69164_/X _69166_/X _69116_/X _69167_/X sky130_fd_sc_hd__a21o_4
X_54393_ _85450_/Q _54376_/X _54392_/Y _54393_/Y sky130_fd_sc_hd__o21ai_4
X_66379_ _66433_/A _66415_/B _84134_/Q _66379_/X sky130_fd_sc_hd__and3_4
X_56132_ _56112_/X _56130_/X _56131_/Y _85291_/D sky130_fd_sc_hd__o21ai_4
X_68118_ _68097_/X _66743_/Y _68110_/X _68117_/Y _68118_/X sky130_fd_sc_hd__a211o_4
X_53344_ _53342_/Y _53328_/X _53343_/X _53344_/Y sky130_fd_sc_hd__a21oi_4
X_84164_ _84166_/CLK _65989_/X _84164_/Q sky130_fd_sc_hd__dfxtp_4
X_50556_ _50556_/A _50556_/B _50556_/Y sky130_fd_sc_hd__nand2_4
X_81376_ _81473_/CLK _81376_/D _81376_/Q sky130_fd_sc_hd__dfxtp_4
X_69098_ _69607_/A _69098_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_460_0_CLK clkbuf_9_230_0_CLK/X _85974_/CLK sky130_fd_sc_hd__clkbuf_1
X_83115_ _83115_/CLK _83115_/D _83115_/Q sky130_fd_sc_hd__dfxtp_4
X_80327_ _84750_/Q _84142_/Q _80327_/Y sky130_fd_sc_hd__nand2_4
X_56063_ _74312_/C _55997_/X _56063_/Y sky130_fd_sc_hd__xnor2_4
X_68049_ _68049_/A _68049_/B _68049_/Y sky130_fd_sc_hd__nand2_4
X_53275_ _53271_/Y _53272_/X _53274_/X _85664_/D sky130_fd_sc_hd__a21oi_4
X_84095_ _80928_/CLK _66827_/X _80919_/D sky130_fd_sc_hd__dfxtp_4
X_50487_ _52194_/A _50492_/B _50497_/C _50487_/X sky130_fd_sc_hd__and3_4
X_55014_ _55012_/Y _54998_/X _55013_/X _55014_/Y sky130_fd_sc_hd__a21oi_4
X_52226_ _85864_/Q _52214_/X _52225_/Y _52226_/Y sky130_fd_sc_hd__o21ai_4
X_71060_ _71058_/A _71082_/B _71055_/C _71060_/Y sky130_fd_sc_hd__nand3_4
X_83046_ _83046_/CLK _74526_/Y _83046_/Q sky130_fd_sc_hd__dfxtp_4
X_87923_ _87671_/CLK _42322_/Y _87923_/Q sky130_fd_sc_hd__dfxtp_4
X_80258_ _80257_/Y _80259_/B sky130_fd_sc_hd__inv_2
X_70011_ _68823_/A _70011_/X sky130_fd_sc_hd__buf_2
X_59822_ _59756_/A _59822_/X sky130_fd_sc_hd__buf_2
X_52157_ _52155_/Y _52145_/X _52156_/X _52157_/Y sky130_fd_sc_hd__a21oi_4
X_87854_ _86984_/CLK _87854_/D _68490_/A sky130_fd_sc_hd__dfxtp_4
X_80189_ _80189_/A _80198_/A _80189_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_475_0_CLK clkbuf_9_237_0_CLK/X _86381_/CLK sky130_fd_sc_hd__clkbuf_1
X_51108_ _86072_/Q _51101_/X _51107_/Y _51108_/Y sky130_fd_sc_hd__o21ai_4
X_86805_ _87888_/CLK _86805_/D _86805_/Q sky130_fd_sc_hd__dfxtp_4
X_59753_ _72584_/C _59753_/B _60312_/C _60312_/D _59753_/Y sky130_fd_sc_hd__nand4_4
X_52088_ _52086_/Y _52066_/X _52087_/Y _85891_/D sky130_fd_sc_hd__a21boi_4
X_56965_ _56949_/X _56634_/X _45582_/A _56989_/A _85109_/D sky130_fd_sc_hd__a2bb2o_4
X_87785_ _87789_/CLK _87785_/D _87785_/Q sky130_fd_sc_hd__dfxtp_4
X_84997_ _86855_/CLK _57478_/Y _57473_/B sky130_fd_sc_hd__dfxtp_4
X_58704_ _58605_/X _85942_/Q _58679_/X _58704_/X sky130_fd_sc_hd__o21a_4
X_43930_ _41416_/X _43928_/X _87195_/Q _43929_/X _87195_/D sky130_fd_sc_hd__a2bb2o_4
X_51039_ _51039_/A _51039_/X sky130_fd_sc_hd__buf_2
X_55916_ _45046_/A _55607_/A _44099_/X _55915_/X _55916_/X sky130_fd_sc_hd__a211o_4
X_74750_ _74764_/A _74804_/A sky130_fd_sc_hd__buf_2
X_86736_ _86736_/CLK _46454_/Y _86736_/Q sky130_fd_sc_hd__dfxtp_4
X_71962_ _71957_/A _48887_/Y _71962_/Y sky130_fd_sc_hd__nand2_4
X_59684_ _59642_/X _59684_/X sky130_fd_sc_hd__buf_2
X_83948_ _83973_/CLK _83948_/D _80804_/D sky130_fd_sc_hd__dfxtp_4
X_56896_ _46155_/X _55208_/B _56895_/X _44137_/A _56897_/B sky130_fd_sc_hd__a211o_4
X_73701_ _87341_/Q _73701_/B _73701_/Y sky130_fd_sc_hd__nor2_4
X_70913_ _70913_/A _70914_/D sky130_fd_sc_hd__buf_2
X_58635_ _58635_/A _58868_/A sky130_fd_sc_hd__buf_2
X_43861_ _41230_/X _43842_/X _68920_/B _43843_/X _43861_/X sky130_fd_sc_hd__a2bb2o_4
X_55847_ _56233_/C _55489_/A _55469_/X _55846_/X _55847_/X sky130_fd_sc_hd__a211o_4
X_86667_ _86351_/CLK _47134_/Y _59270_/A sky130_fd_sc_hd__dfxtp_4
X_74681_ _74680_/Y _82987_/D sky130_fd_sc_hd__inv_2
X_71893_ _70716_/A _71893_/X sky130_fd_sc_hd__buf_2
X_83879_ _82557_/CLK _69987_/X _82559_/D sky130_fd_sc_hd__dfxtp_4
X_45600_ _45600_/A _45617_/B _45600_/Y sky130_fd_sc_hd__nor2_4
X_76420_ _76387_/A _76403_/B _76400_/X _76420_/X sky130_fd_sc_hd__and3_4
X_42812_ _42812_/A _87706_/D sky130_fd_sc_hd__inv_2
X_73632_ _72978_/X _74244_/B sky130_fd_sc_hd__buf_2
X_85618_ _85630_/CLK _53534_/Y _85618_/Q sky130_fd_sc_hd__dfxtp_4
X_46580_ _82916_/Q _46579_/X _46580_/X sky130_fd_sc_hd__or2_4
X_70844_ _70871_/A _70846_/B _70849_/C _70860_/D _70844_/Y sky130_fd_sc_hd__nand4_4
X_58566_ _86721_/Q _58614_/B _58566_/Y sky130_fd_sc_hd__nor2_4
X_43792_ _43790_/X _43781_/X _41036_/X _87265_/Q _43791_/X _43792_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55778_ _55775_/X _55777_/X _44110_/X _55778_/X sky130_fd_sc_hd__a21o_4
X_86598_ _85959_/CLK _86598_/D _86598_/Q sky130_fd_sc_hd__dfxtp_4
X_45531_ _45511_/X _61430_/A _45530_/X _45531_/Y sky130_fd_sc_hd__o21ai_4
X_57517_ _57514_/Y _57515_/X _57516_/Y _84988_/D sky130_fd_sc_hd__a21boi_4
X_76351_ _76350_/X _76353_/B sky130_fd_sc_hd__inv_2
X_42743_ _42743_/A _51949_/A sky130_fd_sc_hd__buf_2
X_88337_ _88337_/CLK _88337_/D _69597_/B sky130_fd_sc_hd__dfxtp_4
X_54729_ _54729_/A _54729_/X sky130_fd_sc_hd__buf_2
X_73563_ _73497_/A _65908_/B _73563_/X sky130_fd_sc_hd__and2_4
X_85549_ _86256_/CLK _53885_/Y _85549_/Q sky130_fd_sc_hd__dfxtp_4
X_70775_ _70867_/A _70779_/B _70791_/C _70791_/D _70775_/Y sky130_fd_sc_hd__nand4_4
X_58497_ _84834_/Q _58498_/A sky130_fd_sc_hd__inv_2
Xclkbuf_10_413_0_CLK clkbuf_9_206_0_CLK/X _85335_/CLK sky130_fd_sc_hd__clkbuf_1
X_75302_ _75298_/X _75301_/X _75309_/A sky130_fd_sc_hd__xor2_4
X_48250_ _66101_/B _48241_/X _48249_/Y _48250_/Y sky130_fd_sc_hd__o21ai_4
X_72514_ _72514_/A _72607_/C sky130_fd_sc_hd__buf_2
X_79070_ _79065_/Y _79070_/B _79071_/B sky130_fd_sc_hd__xor2_4
X_45462_ _45458_/X _45461_/X _45446_/X _45462_/X sky130_fd_sc_hd__a21o_4
X_57448_ _57448_/A _57463_/B _57448_/X sky130_fd_sc_hd__or2_4
X_76282_ _76282_/A _76276_/X _76282_/C _76283_/A sky130_fd_sc_hd__nand3_4
X_88268_ _88268_/CLK _41154_/X _68549_/B sky130_fd_sc_hd__dfxtp_4
X_42674_ _42665_/X _42666_/X _41045_/X _87776_/Q _42673_/X _42674_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73494_ _73494_/A _73493_/X _73494_/Y sky130_fd_sc_hd__nand2_4
X_47201_ _47201_/A _51220_/D sky130_fd_sc_hd__buf_2
X_78021_ _78021_/A _82176_/Q _78021_/C _78022_/A sky130_fd_sc_hd__nand3_4
X_44413_ _44454_/A _44413_/X sky130_fd_sc_hd__buf_2
X_75233_ _75212_/Y _75233_/B _75233_/X sky130_fd_sc_hd__or2_4
X_87219_ _88180_/CLK _87219_/D _87219_/Q sky130_fd_sc_hd__dfxtp_4
X_41625_ _41588_/X _40546_/A _41624_/X _41625_/Y sky130_fd_sc_hd__o21ai_4
X_48181_ _50048_/A _50232_/B _48181_/Y sky130_fd_sc_hd__nand2_4
X_72445_ _72381_/A _72445_/X sky130_fd_sc_hd__buf_2
X_45393_ _45393_/A _45393_/Y sky130_fd_sc_hd__inv_2
X_57379_ _45886_/X _45882_/A _45898_/X _73916_/B _44038_/X _57379_/Y
+ sky130_fd_sc_hd__a41oi_4
X_88199_ _88133_/CLK _41522_/Y _66857_/B sky130_fd_sc_hd__dfxtp_4
X_47132_ _54565_/D _52872_/D sky130_fd_sc_hd__buf_2
X_59118_ _59118_/A _59068_/B _59118_/Y sky130_fd_sc_hd__nor2_4
X_44344_ _41697_/X _44326_/X _87155_/Q _44327_/X _87155_/D sky130_fd_sc_hd__a2bb2o_4
X_75164_ _75133_/Y _75147_/Y _75164_/Y sky130_fd_sc_hd__nand2_4
X_41556_ _41555_/Y _41556_/X sky130_fd_sc_hd__buf_2
X_72376_ _72373_/Y _72375_/Y _72292_/X _72376_/X sky130_fd_sc_hd__a21o_4
X_60390_ _60473_/C _60399_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_428_0_CLK clkbuf_9_214_0_CLK/X _84119_/CLK sky130_fd_sc_hd__clkbuf_1
X_74115_ _57605_/B _74115_/B _74116_/B sky130_fd_sc_hd__xor2_4
X_40507_ _40506_/Y _40507_/X sky130_fd_sc_hd__buf_2
X_47063_ _47063_/A _52833_/B _47063_/Y sky130_fd_sc_hd__nand2_4
X_59049_ _59048_/X _85661_/Q _59010_/X _59049_/X sky130_fd_sc_hd__o21a_4
X_71327_ _71335_/A _71335_/B _70472_/X _71327_/Y sky130_fd_sc_hd__nand3_4
X_44275_ _44274_/X _57327_/B sky130_fd_sc_hd__buf_2
X_79972_ _84927_/Q _84175_/Q _79972_/Y sky130_fd_sc_hd__nand2_4
X_75095_ _80676_/Q _80932_/D _75096_/A sky130_fd_sc_hd__nor2_4
X_41487_ _41457_/A _41487_/X sky130_fd_sc_hd__buf_2
X_46014_ _45981_/X _46014_/X sky130_fd_sc_hd__buf_2
X_43226_ _43162_/A _43226_/X sky130_fd_sc_hd__buf_2
X_62060_ _59699_/A _62060_/X sky130_fd_sc_hd__buf_2
X_74046_ _57590_/B _74046_/B _74046_/X sky130_fd_sc_hd__xor2_4
X_78923_ _78921_/Y _78923_/B _78931_/B sky130_fd_sc_hd__xor2_4
X_40438_ _82325_/Q _40907_/B _40438_/X sky130_fd_sc_hd__or2_4
X_71258_ _71258_/A _71232_/B _71141_/B _71258_/Y sky130_fd_sc_hd__nand3_4
X_61011_ _60963_/X _61010_/Y _60999_/X _76989_/A _60898_/X _84541_/D
+ sky130_fd_sc_hd__o32a_4
X_70209_ _70209_/A _70209_/X sky130_fd_sc_hd__buf_2
X_43157_ _43146_/X _43149_/X _40854_/X _73198_/A _43154_/X _43158_/A
+ sky130_fd_sc_hd__o32ai_4
X_78854_ _78874_/A _78854_/B _78854_/Y sky130_fd_sc_hd__nor2_4
X_40369_ _40368_/X _81183_/Q _40369_/X sky130_fd_sc_hd__or2_4
X_71189_ _71137_/A _71189_/B _71190_/A sky130_fd_sc_hd__nor2_4
X_42108_ _42099_/X _42094_/X _41045_/X _88032_/Q _42096_/X _42109_/A
+ sky130_fd_sc_hd__o32ai_4
X_77805_ _82154_/Q _77805_/B _77805_/X sky130_fd_sc_hd__xor2_4
X_47965_ _47946_/A _47965_/B _47965_/X sky130_fd_sc_hd__and2_4
X_43088_ _43085_/X _43086_/X _40712_/X _43087_/Y _43058_/X _43088_/Y
+ sky130_fd_sc_hd__o32ai_4
X_78785_ _82528_/Q _78784_/A _82496_/D sky130_fd_sc_hd__xnor2_4
X_75997_ _81333_/Q _81421_/Q _76005_/B sky130_fd_sc_hd__or2_4
X_49704_ _59376_/B _49687_/X _49703_/Y _49704_/Y sky130_fd_sc_hd__o21ai_4
X_46916_ _82946_/Q _46916_/Y sky130_fd_sc_hd__inv_2
X_42039_ _42028_/X _42024_/X _40885_/X _73320_/A _42025_/X _42040_/A
+ sky130_fd_sc_hd__o32ai_4
X_65750_ _65735_/A _86476_/Q _65750_/X sky130_fd_sc_hd__and2_4
X_77736_ _82259_/Q _77736_/Y sky130_fd_sc_hd__inv_2
X_62962_ _62960_/X _62942_/X _62961_/Y _84366_/D sky130_fd_sc_hd__a21oi_4
X_74948_ _74958_/A _74959_/A _74949_/B sky130_fd_sc_hd__xor2_4
X_47896_ _47892_/Y _47846_/X _47895_/X _47896_/Y sky130_fd_sc_hd__a21oi_4
X_64701_ _64619_/A _64701_/X sky130_fd_sc_hd__buf_2
X_49635_ _86351_/Q _49632_/X _49634_/Y _49635_/Y sky130_fd_sc_hd__o21ai_4
X_61913_ _61960_/A _61960_/B _78069_/B _61913_/Y sky130_fd_sc_hd__nor3_4
X_46847_ _46846_/Y _52709_/D sky130_fd_sc_hd__buf_2
X_65681_ _65757_/A _65681_/X sky130_fd_sc_hd__buf_2
X_77667_ _77665_/X _77639_/Y _77667_/C _77667_/X sky130_fd_sc_hd__and3_4
X_62893_ _62893_/A _62893_/X sky130_fd_sc_hd__buf_2
X_74879_ _74879_/A _74879_/B _81216_/D sky130_fd_sc_hd__xor2_4
X_67420_ _67062_/X _67517_/A sky130_fd_sc_hd__buf_2
X_79406_ _79404_/X _79405_/X _79419_/B sky130_fd_sc_hd__xnor2_4
X_64632_ _64599_/X _83312_/Q _64600_/X _64631_/X _64632_/X sky130_fd_sc_hd__a211o_4
X_76618_ _76593_/Y _76597_/B _76595_/Y _76618_/X sky130_fd_sc_hd__o21a_4
X_49566_ _49564_/Y _49541_/X _49565_/X _86364_/D sky130_fd_sc_hd__a21oi_4
X_61844_ _84722_/Q _61844_/X sky130_fd_sc_hd__buf_2
X_46778_ _46778_/A _52667_/B sky130_fd_sc_hd__inv_2
X_77598_ _77584_/A _77584_/B _77583_/A _77606_/A sky130_fd_sc_hd__o21a_4
X_48517_ _48651_/A _48517_/X sky130_fd_sc_hd__buf_2
X_67351_ _67347_/X _67350_/X _67113_/X _67351_/Y sky130_fd_sc_hd__a21oi_4
X_79337_ _79324_/X _79335_/X _79336_/X _79337_/Y sky130_fd_sc_hd__a21oi_4
X_64563_ _64665_/A _64696_/A sky130_fd_sc_hd__buf_2
X_45729_ _45726_/X _45728_/Y _45714_/X _45729_/Y sky130_fd_sc_hd__a21oi_4
X_76549_ _81372_/Q _76548_/X _81340_/D sky130_fd_sc_hd__xor2_4
X_49497_ _49444_/A _49502_/A sky130_fd_sc_hd__buf_2
X_61775_ _59730_/A _61776_/D sky130_fd_sc_hd__buf_2
X_66302_ _66225_/X _84966_/Q _66118_/X _66301_/X _66303_/B sky130_fd_sc_hd__a211o_4
Xclkbuf_8_40_0_CLK clkbuf_8_41_0_CLK/A clkbuf_8_40_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_63514_ _59407_/A _63491_/B _63514_/C _63491_/D _63514_/Y sky130_fd_sc_hd__nand4_4
X_48448_ _48448_/A _48449_/A sky130_fd_sc_hd__inv_2
X_60726_ _60725_/Y _60726_/Y sky130_fd_sc_hd__inv_2
X_67282_ _67141_/X _67268_/Y _67269_/X _67281_/Y _67282_/X sky130_fd_sc_hd__a211o_4
X_79268_ _79266_/X _79276_/B _79268_/Y sky130_fd_sc_hd__xnor2_4
X_64494_ _64494_/A _64494_/B _64207_/A _64494_/X sky130_fd_sc_hd__and3_4
X_69021_ _69021_/A _74186_/A _69021_/X sky130_fd_sc_hd__and2_4
X_66233_ _66230_/Y _66205_/X _66232_/X _84147_/D sky130_fd_sc_hd__a21o_4
X_78219_ _78228_/A _78228_/B _78225_/A sky130_fd_sc_hd__xor2_4
X_63445_ _63434_/X _63435_/X _63438_/X _63442_/X _63444_/Y _63445_/Y
+ sky130_fd_sc_hd__o41ai_4
X_48379_ _48379_/A _74373_/B sky130_fd_sc_hd__inv_2
X_60657_ _60713_/A _63540_/A sky130_fd_sc_hd__buf_2
X_79199_ _79197_/Y _79198_/Y _79203_/A sky130_fd_sc_hd__nand2_4
X_50410_ _50432_/A _48391_/X _50410_/Y sky130_fd_sc_hd__nand2_4
X_81230_ _81227_/CLK _81038_/Q _81230_/Q sky130_fd_sc_hd__dfxtp_4
X_66164_ _66164_/A _66164_/B _66164_/C _66164_/Y sky130_fd_sc_hd__nor3_4
X_51390_ _86019_/Q _51387_/X _51389_/Y _51390_/Y sky130_fd_sc_hd__o21ai_4
X_63376_ _63400_/A _63376_/B _63400_/C _63376_/X sky130_fd_sc_hd__and3_4
X_60588_ _60588_/A _60588_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_55_0_CLK clkbuf_8_55_0_CLK/A clkbuf_8_55_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_65115_ _64946_/A _65115_/B _65115_/X sky130_fd_sc_hd__and2_4
X_50341_ _50317_/X _50341_/B _50341_/Y sky130_fd_sc_hd__nand2_4
X_62327_ _62033_/A _62327_/X sky130_fd_sc_hd__buf_2
X_81161_ _81125_/CLK _74895_/B _41584_/A sky130_fd_sc_hd__dfxtp_4
X_66095_ _65990_/X _86228_/Q _66021_/X _66094_/X _66095_/X sky130_fd_sc_hd__a211o_4
X_80112_ _80121_/A _80121_/B _80112_/Y sky130_fd_sc_hd__xnor2_4
X_53060_ _53040_/X _53060_/B _53060_/Y sky130_fd_sc_hd__nand2_4
X_65046_ _84217_/Q _65047_/C sky130_fd_sc_hd__inv_2
X_69923_ _69877_/A _69923_/B _69923_/X sky130_fd_sc_hd__and2_4
X_50272_ _50251_/X _47924_/B _50272_/Y sky130_fd_sc_hd__nand2_4
X_62258_ _59931_/X _61780_/X _62257_/X _62258_/X sky130_fd_sc_hd__a21o_4
X_81092_ _82084_/CLK _79563_/Y _81092_/Q sky130_fd_sc_hd__dfxtp_4
X_52011_ _50308_/A _51972_/X _51958_/C _52011_/X sky130_fd_sc_hd__and3_4
X_61209_ _64303_/A _64234_/B sky130_fd_sc_hd__buf_2
X_80043_ _80025_/Y _80043_/B _80043_/X sky130_fd_sc_hd__or2_4
X_84920_ _84905_/CLK _84920_/D _58149_/A sky130_fd_sc_hd__dfxtp_4
X_69854_ _44573_/A _66550_/X _66552_/X _69853_/X _69855_/B sky130_fd_sc_hd__a211o_4
X_62189_ _63348_/A _59700_/Y _61695_/A _59840_/A _62189_/X sky130_fd_sc_hd__a2bb2o_4
X_68805_ _87586_/Q _68757_/X _68731_/X _68804_/Y _68805_/X sky130_fd_sc_hd__a211o_4
X_84851_ _83438_/CLK _84851_/D _84851_/Q sky130_fd_sc_hd__dfxtp_4
X_69785_ _69785_/A _69785_/B _69785_/Y sky130_fd_sc_hd__nand2_4
X_66997_ _66642_/A _66997_/X sky130_fd_sc_hd__buf_2
X_83802_ _83820_/CLK _70309_/X _74729_/A sky130_fd_sc_hd__dfxtp_4
X_56750_ _56593_/A _56750_/B _56749_/X _56750_/Y sky130_fd_sc_hd__nand3_4
X_68736_ _86993_/Q _68707_/X _68630_/X _68735_/X _68736_/X sky130_fd_sc_hd__a211o_4
X_87570_ _83153_/CLK _87570_/D _43115_/A sky130_fd_sc_hd__dfxtp_4
X_53962_ _85533_/Q _53940_/X _53961_/Y _53962_/Y sky130_fd_sc_hd__o21ai_4
X_65948_ _65859_/X _85630_/Q _65860_/X _65947_/X _65948_/X sky130_fd_sc_hd__a211o_4
X_84782_ _83438_/CLK _84782_/D _84782_/Q sky130_fd_sc_hd__dfxtp_4
X_81994_ _81994_/CLK _81994_/D _77050_/A sky130_fd_sc_hd__dfxtp_4
X_55701_ _55701_/A _74284_/C sky130_fd_sc_hd__buf_2
X_86521_ _83584_/CLK _48453_/Y _72993_/B sky130_fd_sc_hd__dfxtp_4
X_52913_ _52911_/Y _52892_/X _52912_/X _52913_/Y sky130_fd_sc_hd__a21oi_4
X_83733_ _86317_/CLK _83733_/D _47410_/A sky130_fd_sc_hd__dfxtp_4
X_56681_ _83327_/Q _56684_/C sky130_fd_sc_hd__buf_2
X_80945_ _80968_/CLK _80945_/D _80945_/Q sky130_fd_sc_hd__dfxtp_4
X_68667_ _57803_/A _68669_/A sky130_fd_sc_hd__buf_2
X_53893_ _50677_/A _53875_/B _53888_/C _53893_/X sky130_fd_sc_hd__and3_4
X_65879_ _65876_/X _85571_/Q _65669_/X _65878_/X _65879_/X sky130_fd_sc_hd__a211o_4
X_58420_ _84852_/Q _58421_/A sky130_fd_sc_hd__inv_2
X_55632_ _45416_/A _55605_/X _44101_/A _55631_/X _55632_/X sky130_fd_sc_hd__a211o_4
X_67618_ _57776_/A _68442_/A sky130_fd_sc_hd__buf_2
X_86452_ _85535_/CLK _49023_/Y _64951_/B sky130_fd_sc_hd__dfxtp_4
X_52844_ _85744_/Q _52821_/X _52843_/Y _52844_/Y sky130_fd_sc_hd__o21ai_4
X_83664_ _86089_/CLK _83664_/D _46850_/A sky130_fd_sc_hd__dfxtp_4
X_80876_ _80849_/CLK _75667_/B _80876_/Q sky130_fd_sc_hd__dfxtp_4
X_68598_ _68479_/A _68599_/A sky130_fd_sc_hd__buf_2
X_85403_ _85499_/CLK _54653_/Y _85403_/Q sky130_fd_sc_hd__dfxtp_4
X_58351_ _84871_/Q _58352_/A sky130_fd_sc_hd__buf_2
X_82615_ _82711_/CLK _79001_/B _82615_/Q sky130_fd_sc_hd__dfxtp_4
X_55563_ _55826_/A _55836_/A sky130_fd_sc_hd__buf_2
X_86383_ _86384_/CLK _86383_/D _58800_/B sky130_fd_sc_hd__dfxtp_4
X_67549_ _67546_/X _67548_/X _67502_/X _67555_/A sky130_fd_sc_hd__a21o_4
X_52775_ _52775_/A _52775_/B _52775_/C _52775_/D _52775_/X sky130_fd_sc_hd__and4_4
X_83595_ _86749_/CLK _71132_/Y _49184_/A sky130_fd_sc_hd__dfxtp_4
X_57302_ _57302_/A _57302_/Y sky130_fd_sc_hd__inv_2
X_88122_ _87865_/CLK _88122_/D _67183_/B sky130_fd_sc_hd__dfxtp_4
X_54514_ _54518_/A _53336_/B _54514_/Y sky130_fd_sc_hd__nand2_4
X_85334_ _85334_/CLK _55019_/Y _85334_/Q sky130_fd_sc_hd__dfxtp_4
X_51726_ _51709_/X _51721_/X _51715_/C _53249_/D _51726_/X sky130_fd_sc_hd__and4_4
X_70560_ _70533_/X _83749_/Q _70559_/Y _83749_/D sky130_fd_sc_hd__a21o_4
X_58282_ _58341_/A _58282_/X sky130_fd_sc_hd__buf_2
X_82546_ _82541_/CLK _83866_/Q _82546_/Q sky130_fd_sc_hd__dfxtp_4
X_55494_ _45582_/A _55492_/X _44047_/X _55493_/Y _55494_/X sky130_fd_sc_hd__a211o_4
X_57233_ _57327_/B _57326_/C sky130_fd_sc_hd__buf_2
X_69219_ _88045_/Q _69217_/X _68976_/X _69218_/X _69219_/X sky130_fd_sc_hd__a211o_4
X_88053_ _88324_/CLK _42062_/Y _88053_/Q sky130_fd_sc_hd__dfxtp_4
X_54445_ _54443_/Y _54422_/X _54444_/X _85441_/D sky130_fd_sc_hd__a21oi_4
X_85265_ _83025_/CLK _56236_/Y _85265_/Q sky130_fd_sc_hd__dfxtp_4
X_51657_ _52593_/A _51657_/X sky130_fd_sc_hd__buf_2
X_70491_ HASH_ADDR[0] _70491_/Y sky130_fd_sc_hd__inv_2
X_82477_ _82570_/CLK _78469_/X _78103_/B sky130_fd_sc_hd__dfxtp_4
X_87004_ _83139_/CLK _87004_/D _44675_/A sky130_fd_sc_hd__dfxtp_4
X_41410_ _41410_/A _41410_/Y sky130_fd_sc_hd__inv_2
X_72230_ _72228_/X _85976_/Q _72229_/X _72230_/Y sky130_fd_sc_hd__o21ai_4
X_84216_ _84228_/CLK _84216_/D _84216_/Q sky130_fd_sc_hd__dfxtp_4
X_50608_ _86168_/Q _50563_/X _50607_/Y _50608_/Y sky130_fd_sc_hd__o21ai_4
X_81428_ _81428_/CLK _81460_/Q _76058_/B sky130_fd_sc_hd__dfxtp_4
X_57164_ _57170_/B _56808_/A _57155_/D _57129_/Y _57164_/X sky130_fd_sc_hd__and4_4
X_42390_ _40391_/X _42388_/X _87887_/Q _42389_/X _87887_/D sky130_fd_sc_hd__a2bb2o_4
X_54376_ _54376_/A _54376_/X sky130_fd_sc_hd__buf_2
X_85196_ _80670_/CLK _85196_/D _85196_/Q sky130_fd_sc_hd__dfxtp_4
X_51588_ _51580_/A _51603_/B _51603_/C _53113_/D _51588_/X sky130_fd_sc_hd__and4_4
X_56115_ _56131_/A _56115_/B _85293_/Q _56115_/Y sky130_fd_sc_hd__nand3_4
X_41341_ _41340_/X _41341_/X sky130_fd_sc_hd__buf_2
X_53327_ _85654_/Q _53324_/X _53326_/Y _53327_/Y sky130_fd_sc_hd__o21ai_4
X_72161_ _57790_/X _72162_/B sky130_fd_sc_hd__buf_2
X_84147_ _84231_/CLK _84147_/D _80397_/B sky130_fd_sc_hd__dfxtp_4
X_50539_ _48667_/A _50552_/B _50552_/C _50539_/X sky130_fd_sc_hd__and3_4
X_57095_ _56561_/X _57087_/X _56931_/X _45386_/A _57192_/A _85089_/D
+ sky130_fd_sc_hd__a32o_4
X_81359_ _81492_/CLK _81359_/D _76343_/A sky130_fd_sc_hd__dfxtp_4
X_71112_ _71003_/A _71112_/X sky130_fd_sc_hd__buf_2
X_44060_ _44059_/X _44060_/X sky130_fd_sc_hd__buf_2
X_56046_ _55907_/X _55914_/X _74306_/C sky130_fd_sc_hd__and2_4
X_41272_ _41271_/Y _41272_/X sky130_fd_sc_hd__buf_2
X_53258_ _53256_/Y _53242_/X _53257_/X _85667_/D sky130_fd_sc_hd__a21oi_4
X_72092_ _72091_/X _53917_/B _72092_/Y sky130_fd_sc_hd__nand2_4
X_84078_ _84014_/CLK _67235_/X _84078_/Q sky130_fd_sc_hd__dfxtp_4
X_43011_ _40548_/X _51934_/A _87604_/Q _42634_/A _87604_/D sky130_fd_sc_hd__a2bb2o_4
X_52209_ _52207_/Y _52117_/X _52208_/Y _85868_/D sky130_fd_sc_hd__a21boi_4
X_71043_ _71041_/X _70588_/A _71276_/C _71039_/D _71043_/Y sky130_fd_sc_hd__nand4_4
X_83029_ _85269_/CLK _83029_/D _45094_/A sky130_fd_sc_hd__dfxtp_4
X_87906_ _87394_/CLK _42354_/X _87906_/Q sky130_fd_sc_hd__dfxtp_4
X_75920_ _84518_/Q _84390_/Q _75920_/X sky130_fd_sc_hd__xor2_4
X_53189_ _53189_/A _53189_/X sky130_fd_sc_hd__buf_2
X_59805_ _59805_/A _59805_/Y sky130_fd_sc_hd__inv_2
X_75851_ _81104_/Q _75851_/B _75867_/A sky130_fd_sc_hd__xnor2_4
X_87837_ _87588_/CLK _42516_/Y _74071_/A sky130_fd_sc_hd__dfxtp_4
X_57997_ _45926_/X _57997_/X sky130_fd_sc_hd__buf_2
X_74802_ _83848_/Q _74735_/X _74799_/X _74800_/X _74801_/X _74802_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_47750_ _47744_/Y _47745_/X _47749_/X _86602_/D sky130_fd_sc_hd__a21oi_4
X_59736_ _59842_/A _59737_/A sky130_fd_sc_hd__buf_2
X_78570_ _78569_/B _78569_/C _78569_/A _78574_/C sky130_fd_sc_hd__o21ai_4
X_44962_ _44957_/Y _44961_/Y _44889_/X _44962_/X sky130_fd_sc_hd__a21o_4
X_56948_ _44214_/X _56584_/X _85117_/Q _56947_/X _85117_/D sky130_fd_sc_hd__a2bb2o_4
X_75782_ _75771_/Y _75775_/Y _75782_/Y sky130_fd_sc_hd__nor2_4
X_87768_ _87520_/CLK _42692_/Y _87768_/Q sky130_fd_sc_hd__dfxtp_4
X_72994_ _72978_/X _83073_/Q _72992_/X _72993_/X _72994_/X sky130_fd_sc_hd__a211o_4
X_46701_ _54314_/B _46701_/X sky130_fd_sc_hd__buf_2
X_77521_ _77502_/A _77514_/A _77521_/Y sky130_fd_sc_hd__nor2_4
X_43913_ _43913_/A _87202_/D sky130_fd_sc_hd__inv_2
X_74733_ _83826_/Q _74716_/X _74720_/X _74730_/Y _74732_/X _80643_/A
+ sky130_fd_sc_hd__a2111o_4
X_86719_ _86398_/CLK _86719_/D _86719_/Q sky130_fd_sc_hd__dfxtp_4
X_47681_ _86609_/Q _47666_/X _47680_/Y _47681_/Y sky130_fd_sc_hd__o21ai_4
X_71945_ _74523_/A _71001_/C _71349_/D _71945_/D _71945_/Y sky130_fd_sc_hd__nand4_4
X_59667_ _59824_/B _59668_/B sky130_fd_sc_hd__buf_2
X_44893_ _44892_/X _44894_/B sky130_fd_sc_hd__buf_2
X_56879_ _56645_/Y _56860_/X _83330_/Q _56880_/B sky130_fd_sc_hd__nand3_4
X_87699_ _87888_/CLK _42825_/X _66535_/B sky130_fd_sc_hd__dfxtp_4
X_49420_ _49420_/A _49420_/B _49420_/C _46716_/X _49420_/X sky130_fd_sc_hd__and4_4
X_46632_ _46627_/Y _46598_/X _46631_/X _86720_/D sky130_fd_sc_hd__a21oi_4
X_58618_ _58618_/A _58618_/X sky130_fd_sc_hd__buf_2
X_77452_ _77452_/A _77451_/X _82193_/D sky130_fd_sc_hd__xnor2_4
X_43844_ _41179_/X _43842_/X _87238_/Q _43843_/X _43844_/X sky130_fd_sc_hd__a2bb2o_4
X_74664_ _74664_/A _74664_/Y sky130_fd_sc_hd__inv_2
X_71876_ _70543_/Y _71883_/B _71873_/X _71874_/D _71876_/Y sky130_fd_sc_hd__nor4_4
X_59598_ _59598_/A _59544_/A _59544_/B _59544_/D _60630_/C sky130_fd_sc_hd__nand4_4
Xclkbuf_10_352_0_CLK clkbuf_9_176_0_CLK/X _83736_/CLK sky130_fd_sc_hd__clkbuf_1
X_76403_ _76400_/X _76403_/B _76406_/A sky130_fd_sc_hd__nand2_4
X_49351_ _49349_/Y _48194_/X _49350_/Y _86404_/D sky130_fd_sc_hd__a21boi_4
X_73615_ _72874_/A _73641_/A sky130_fd_sc_hd__buf_2
X_46563_ _83781_/Q _54077_/B sky130_fd_sc_hd__inv_2
X_70827_ _70358_/X _70827_/B _70827_/C _70828_/A sky130_fd_sc_hd__nor3_4
X_58549_ _58334_/X _58546_/Y _58548_/Y _58549_/Y sky130_fd_sc_hd__a21oi_4
X_77383_ _77382_/B _77381_/Y _77382_/A _77383_/Y sky130_fd_sc_hd__o21ai_4
X_43775_ _43756_/A _43776_/A sky130_fd_sc_hd__buf_2
X_74595_ _45199_/A _74582_/X _74594_/X _83022_/D sky130_fd_sc_hd__o21ai_4
X_40987_ _40941_/A _40987_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_982_0_CLK clkbuf_9_491_0_CLK/X _85837_/CLK sky130_fd_sc_hd__clkbuf_1
X_48302_ _48193_/X _48302_/X sky130_fd_sc_hd__buf_2
X_79122_ _79122_/A _79122_/B _82499_/D sky130_fd_sc_hd__nand2_4
X_45514_ _45506_/X _45510_/X _45513_/Y _45514_/Y sky130_fd_sc_hd__a21oi_4
X_76334_ _76330_/Y _76331_/Y _76333_/Y _76336_/A sky130_fd_sc_hd__or3_4
X_42726_ _41179_/X _42717_/X _87750_/Q _42718_/X _87750_/D sky130_fd_sc_hd__a2bb2o_4
X_49282_ _71959_/A _49283_/B sky130_fd_sc_hd__buf_2
X_61560_ _61541_/A _61560_/B _61541_/C _61560_/Y sky130_fd_sc_hd__nand3_4
X_73546_ _73367_/A _73546_/X sky130_fd_sc_hd__buf_2
X_46494_ _81196_/Q _46495_/B sky130_fd_sc_hd__inv_2
X_70758_ _70758_/A _70758_/B _70758_/C _70764_/A sky130_fd_sc_hd__nor3_4
Xclkbuf_9_473_0_CLK clkbuf_8_236_0_CLK/X clkbuf_9_473_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_48233_ _48193_/X _48233_/X sky130_fd_sc_hd__buf_2
X_60511_ _79149_/A _60246_/X _60586_/D _60510_/Y _60511_/Y sky130_fd_sc_hd__a2bb2oi_4
X_79053_ _79053_/A _79053_/B _79054_/A sky130_fd_sc_hd__nand2_4
X_45445_ _55596_/B _45412_/X _45443_/X _45444_/Y _45445_/X sky130_fd_sc_hd__a211o_4
X_76265_ _76261_/X _76262_/Y _76264_/Y _76267_/A sky130_fd_sc_hd__a21o_4
X_42657_ _42657_/A _42657_/Y sky130_fd_sc_hd__inv_2
X_73477_ _73359_/X _83053_/Q _73406_/X _73476_/X _73477_/X sky130_fd_sc_hd__a211o_4
X_61491_ _61482_/A _61490_/X _61482_/C _61491_/Y sky130_fd_sc_hd__nand3_4
X_70689_ _70689_/A _70692_/B _70692_/C _70689_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_10_367_0_CLK clkbuf_9_183_0_CLK/X _85700_/CLK sky130_fd_sc_hd__clkbuf_1
X_78004_ _78006_/B _78004_/Y sky130_fd_sc_hd__inv_2
X_75216_ _75216_/A _75216_/Y sky130_fd_sc_hd__inv_2
X_63230_ _63230_/A _63316_/B _63295_/C _63267_/D _63230_/X sky130_fd_sc_hd__or4_4
X_41608_ _41607_/X _41608_/X sky130_fd_sc_hd__buf_2
X_48164_ _48164_/A _57489_/B _48163_/X _48164_/Y sky130_fd_sc_hd__nand3_4
X_60442_ _60399_/B _60583_/A _60442_/C _60445_/A sky130_fd_sc_hd__nor3_4
X_72428_ _72428_/A _72428_/B _72428_/Y sky130_fd_sc_hd__nor2_4
X_45376_ _56458_/C _45326_/X _45375_/X _45376_/Y sky130_fd_sc_hd__o21ai_4
X_76196_ _76194_/Y _76196_/B _76192_/X _76196_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_997_0_CLK clkbuf_9_498_0_CLK/X _85884_/CLK sky130_fd_sc_hd__clkbuf_1
X_42588_ _42588_/A _42588_/Y sky130_fd_sc_hd__inv_2
X_47115_ _47115_/A _47116_/A sky130_fd_sc_hd__inv_2
X_44327_ _40509_/X _44327_/X sky130_fd_sc_hd__buf_2
X_63161_ _63161_/A _63113_/B _63161_/C _63149_/X _63161_/X sky130_fd_sc_hd__or4_4
X_75147_ _75144_/Y _75146_/Y _75147_/Y sky130_fd_sc_hd__nor2_4
X_41539_ _41538_/Y _41539_/Y sky130_fd_sc_hd__inv_2
X_60373_ _79538_/A _60323_/X _60372_/Y _60337_/Y _60373_/X sky130_fd_sc_hd__o22a_4
X_72359_ _72287_/X _85325_/Q _72324_/X _72359_/X sky130_fd_sc_hd__o21a_4
X_48095_ _48461_/A _48449_/B sky130_fd_sc_hd__buf_2
Xclkbuf_9_488_0_CLK clkbuf_9_489_0_CLK/A clkbuf_9_488_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_62112_ _61627_/B _62161_/B _62128_/C _62011_/X _62112_/Y sky130_fd_sc_hd__nand4_4
X_47046_ _47046_/A _47047_/A sky130_fd_sc_hd__inv_2
X_44258_ _44258_/A _44256_/A _44258_/Y sky130_fd_sc_hd__nor2_4
X_79955_ _79957_/B _79957_/C _79955_/Y sky130_fd_sc_hd__nand2_4
X_63092_ _58177_/Y _63081_/B _63081_/C _63092_/D _63092_/X sky130_fd_sc_hd__or4_4
X_75078_ _75075_/Y _75077_/Y _75078_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_920_0_CLK clkbuf_9_460_0_CLK/X _87068_/CLK sky130_fd_sc_hd__clkbuf_1
X_43209_ _43209_/A _43209_/Y sky130_fd_sc_hd__inv_2
X_66920_ _66823_/A _66920_/B _66920_/X sky130_fd_sc_hd__and2_4
X_62043_ _61568_/B _61995_/X _62010_/X _62011_/X _62047_/C sky130_fd_sc_hd__nand4_4
X_74029_ _74027_/X _74028_/Y _73982_/X _74029_/X sky130_fd_sc_hd__a21o_4
X_78906_ _78894_/Y _78898_/Y _78900_/A _78906_/Y sky130_fd_sc_hd__a21boi_4
X_44189_ _72806_/A _44189_/X sky130_fd_sc_hd__buf_2
X_79886_ _79871_/X _79873_/B _79885_/Y _79886_/Y sky130_fd_sc_hd__a21boi_4
Xclkbuf_9_411_0_CLK clkbuf_9_411_0_CLK/A clkbuf_9_411_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_66851_ _66534_/A _66851_/X sky130_fd_sc_hd__buf_2
X_78837_ _78834_/X _78837_/B _78838_/B sky130_fd_sc_hd__xor2_4
X_48997_ _48946_/X _48485_/A _48996_/Y _48998_/A sky130_fd_sc_hd__a21o_4
Xclkbuf_10_305_0_CLK clkbuf_9_152_0_CLK/X _83362_/CLK sky130_fd_sc_hd__clkbuf_1
X_65802_ _65888_/A _65802_/B _65802_/C _65802_/Y sky130_fd_sc_hd__nor3_4
X_69570_ _66547_/A _69570_/X sky130_fd_sc_hd__buf_2
X_47948_ _47840_/A _47948_/X sky130_fd_sc_hd__buf_2
X_66782_ _66760_/A _87690_/Q _66782_/X sky130_fd_sc_hd__and2_4
X_78768_ _78767_/Y _78769_/B sky130_fd_sc_hd__inv_2
X_63994_ _63912_/X _63994_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_935_0_CLK clkbuf_9_467_0_CLK/X _87285_/CLK sky130_fd_sc_hd__clkbuf_1
X_68521_ _88109_/Q _68069_/X _68439_/X _68520_/Y _68521_/X sky130_fd_sc_hd__a211o_4
X_65733_ _64828_/A _65733_/X sky130_fd_sc_hd__buf_2
X_77719_ _77710_/A _77709_/X _77717_/A _77723_/C sky130_fd_sc_hd__nand3_4
X_62945_ _58287_/Y _60337_/C _62945_/Y sky130_fd_sc_hd__nor2_4
X_47879_ _47866_/Y _47846_/X _47878_/X _86590_/D sky130_fd_sc_hd__a21oi_4
X_78699_ _78697_/X _78722_/A _78700_/A sky130_fd_sc_hd__and2_4
Xclkbuf_9_426_0_CLK clkbuf_9_427_0_CLK/A clkbuf_9_426_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_49618_ _86354_/Q _49606_/X _49617_/Y _49618_/Y sky130_fd_sc_hd__o21ai_4
X_68452_ _68452_/A _87248_/Q _68452_/X sky130_fd_sc_hd__and2_4
X_80730_ _81048_/CLK _75916_/X _80730_/Q sky130_fd_sc_hd__dfxtp_4
X_65664_ _65664_/A _65663_/Y _65664_/Y sky130_fd_sc_hd__nand2_4
X_50890_ _50918_/A _50908_/A sky130_fd_sc_hd__buf_2
X_62876_ _58483_/A _62841_/X _60309_/C _60202_/A _62876_/Y sky130_fd_sc_hd__nand4_4
X_67403_ _67305_/X _67387_/Y _67390_/X _67402_/Y _67403_/X sky130_fd_sc_hd__a211o_4
X_64615_ _64615_/A _64615_/X sky130_fd_sc_hd__buf_2
X_49549_ _49561_/A _49537_/B _49548_/X _52763_/D _49549_/X sky130_fd_sc_hd__and4_4
X_61827_ _61839_/A _61839_/B _61839_/C _63079_/B _61827_/X sky130_fd_sc_hd__and4_4
X_80661_ _80657_/CLK _80661_/D _46087_/A sky130_fd_sc_hd__dfxtp_4
X_68383_ _45924_/A _68384_/A sky130_fd_sc_hd__buf_2
X_65595_ _64666_/A _65595_/X sky130_fd_sc_hd__buf_2
X_82400_ _82965_/CLK _82208_/Q _82400_/Q sky130_fd_sc_hd__dfxtp_4
X_67334_ _87987_/Q _67236_/X _67284_/X _67333_/X _67334_/X sky130_fd_sc_hd__a211o_4
X_52560_ _65335_/B _52549_/X _52559_/Y _52560_/Y sky130_fd_sc_hd__o21ai_4
X_64546_ _64546_/A _64225_/B _64546_/C _64546_/X sky130_fd_sc_hd__and3_4
X_83380_ _83380_/CLK _71776_/X _83380_/Q sky130_fd_sc_hd__dfxtp_4
X_61758_ _58225_/X _61728_/X _61756_/X _59591_/A _61757_/X _61758_/X
+ sky130_fd_sc_hd__a41o_4
X_80592_ _80581_/X _80592_/Y sky130_fd_sc_hd__inv_2
XPHY_409 sky130_fd_sc_hd__decap_3
X_51511_ _51539_/A _51511_/X sky130_fd_sc_hd__buf_2
X_82331_ _87086_/CLK _77182_/B _82331_/Q sky130_fd_sc_hd__dfxtp_4
X_60709_ _60694_/B _60696_/Y _60708_/Y _60709_/X sky130_fd_sc_hd__o21a_4
X_67265_ _67260_/X _67263_/X _67264_/X _67268_/A sky130_fd_sc_hd__a21o_4
X_52491_ _64974_/B _52470_/X _52490_/Y _52491_/Y sky130_fd_sc_hd__o21ai_4
X_64477_ _61238_/C _64457_/C _64475_/Y _64477_/D _64477_/Y sky130_fd_sc_hd__nand4_4
X_61689_ _61682_/Y _61684_/Y _61334_/A _61685_/Y _61688_/Y _61689_/X
+ sky130_fd_sc_hd__a41o_4
X_69004_ _69004_/A _69004_/B _69004_/X sky130_fd_sc_hd__and2_4
X_54230_ _54230_/A _53060_/B _54230_/Y sky130_fd_sc_hd__nand2_4
X_66216_ _66216_/A _64633_/B _66216_/C _66216_/Y sky130_fd_sc_hd__nand3_4
X_85050_ _85050_/CLK _85050_/D _45504_/A sky130_fd_sc_hd__dfxtp_4
X_51442_ _51170_/A _51467_/C sky130_fd_sc_hd__buf_2
X_63428_ _63400_/A _84900_/Q _63463_/C _63428_/X sky130_fd_sc_hd__and3_4
X_82262_ _82253_/CLK _82262_/D _82262_/Q sky130_fd_sc_hd__dfxtp_4
X_67196_ _87109_/Q _67193_/X _67194_/X _67195_/X _67196_/X sky130_fd_sc_hd__a211o_4
X_84001_ _81755_/CLK _68250_/X _84001_/Q sky130_fd_sc_hd__dfxtp_4
X_81213_ _82288_/CLK _81213_/D _46302_/A sky130_fd_sc_hd__dfxtp_4
X_54161_ _54159_/Y _54144_/X _54160_/X _85493_/D sky130_fd_sc_hd__a21oi_4
X_66147_ _57761_/X _84977_/Q _65950_/X _66146_/X _66147_/X sky130_fd_sc_hd__a211o_4
X_51373_ _51371_/Y _51366_/X _51372_/X _51373_/Y sky130_fd_sc_hd__a21oi_4
X_63359_ _58403_/A _63370_/A _63359_/Y sky130_fd_sc_hd__nor2_4
X_82193_ _82386_/CLK _82193_/D _82193_/Q sky130_fd_sc_hd__dfxtp_4
X_53112_ _53112_/A _53133_/A sky130_fd_sc_hd__buf_2
X_50324_ _50317_/X _48024_/B _50324_/Y sky130_fd_sc_hd__nand2_4
X_81144_ _81197_/CLK _80768_/Q _40639_/A sky130_fd_sc_hd__dfxtp_4
X_54092_ _54090_/Y _54051_/X _54091_/X _54092_/Y sky130_fd_sc_hd__a21oi_4
X_66078_ _65969_/A _66123_/A sky130_fd_sc_hd__buf_2
X_53043_ _53069_/A _53063_/B sky130_fd_sc_hd__buf_2
X_57920_ _57781_/X _57918_/Y _57919_/Y _57893_/X _57795_/X _57920_/X
+ sky130_fd_sc_hd__o32a_4
X_65029_ _64924_/A _65029_/B _65029_/X sky130_fd_sc_hd__and2_4
X_69906_ _69906_/A _87289_/Q _69906_/X sky130_fd_sc_hd__and2_4
X_50255_ _54043_/B _50475_/B sky130_fd_sc_hd__buf_2
X_85952_ _85471_/CLK _85952_/D _85952_/Q sky130_fd_sc_hd__dfxtp_4
X_81075_ _81070_/CLK _81107_/Q _81075_/Q sky130_fd_sc_hd__dfxtp_4
X_80026_ _84932_/Q _84180_/Q _80026_/X sky130_fd_sc_hd__xor2_4
X_84903_ _84903_/CLK _58227_/Y _58225_/A sky130_fd_sc_hd__dfxtp_4
X_57851_ _57811_/X _85401_/Q _57850_/X _57851_/Y sky130_fd_sc_hd__o21ai_4
X_69837_ _69751_/A _69837_/X sky130_fd_sc_hd__buf_2
X_50186_ _50063_/A _51286_/A sky130_fd_sc_hd__buf_2
X_85883_ _86490_/CLK _52131_/Y _65519_/B sky130_fd_sc_hd__dfxtp_4
X_56802_ _56755_/X _57140_/B _56759_/X _83322_/Q _56803_/A sky130_fd_sc_hd__and4_4
X_87622_ _87883_/CLK _42978_/Y _87622_/Q sky130_fd_sc_hd__dfxtp_4
X_84834_ _84308_/CLK _84834_/D _84834_/Q sky130_fd_sc_hd__dfxtp_4
X_57782_ _68714_/A _68342_/A sky130_fd_sc_hd__buf_2
X_69768_ _69768_/A _69768_/X sky130_fd_sc_hd__buf_2
X_54994_ _55072_/A _54994_/X sky130_fd_sc_hd__buf_2
X_59521_ _59521_/A _59571_/B sky130_fd_sc_hd__buf_2
X_56733_ _56739_/A _56733_/X sky130_fd_sc_hd__buf_2
X_68719_ _87493_/Q _68472_/A _68545_/X _68718_/X _68719_/X sky130_fd_sc_hd__a211o_4
X_87553_ _87553_/CLK _43160_/Y _73228_/A sky130_fd_sc_hd__dfxtp_4
X_53945_ _53943_/Y _53892_/X _53944_/Y _85537_/D sky130_fd_sc_hd__a21oi_4
X_84765_ _84760_/CLK _84765_/D _59143_/A sky130_fd_sc_hd__dfxtp_4
X_81977_ _82234_/CLK _83905_/Q _81977_/Q sky130_fd_sc_hd__dfxtp_4
X_69699_ _73033_/A _44299_/A _68933_/X _69698_/Y _69699_/X sky130_fd_sc_hd__a211o_4
X_86504_ _86500_/CLK _48646_/Y _86504_/Q sky130_fd_sc_hd__dfxtp_4
X_40910_ _40870_/X _40871_/X _40909_/X _69923_/B _40867_/X _40911_/A
+ sky130_fd_sc_hd__o32ai_4
X_71730_ _58236_/Y _71718_/X _71729_/Y _83396_/D sky130_fd_sc_hd__o21ai_4
X_83716_ _83716_/CLK _70723_/Y _83716_/Q sky130_fd_sc_hd__dfxtp_4
X_59452_ _59442_/X _83465_/Q _59451_/Y _59452_/X sky130_fd_sc_hd__o21a_4
X_56664_ _56593_/A _83329_/Q _56663_/X _56664_/Y sky130_fd_sc_hd__nand3_4
X_80928_ _80928_/CLK _84104_/Q _75852_/A sky130_fd_sc_hd__dfxtp_4
X_87484_ _87484_/CLK _87484_/D _87484_/Q sky130_fd_sc_hd__dfxtp_4
X_41890_ _41881_/A _41967_/A sky130_fd_sc_hd__buf_2
X_53876_ _53873_/Y _53829_/X _53875_/X _53876_/Y sky130_fd_sc_hd__a21oi_4
X_84696_ _84713_/CLK _84696_/D _80442_/A sky130_fd_sc_hd__dfxtp_4
X_58403_ _58403_/A _58403_/B _58403_/Y sky130_fd_sc_hd__nand2_4
X_55615_ _55615_/A _55615_/X sky130_fd_sc_hd__buf_2
X_86435_ _86436_/CLK _86435_/D _65392_/B sky130_fd_sc_hd__dfxtp_4
X_40841_ _40840_/Y _88325_/D sky130_fd_sc_hd__inv_2
X_52827_ _52818_/A _52831_/B _52818_/C _52827_/D _52827_/X sky130_fd_sc_hd__and4_4
X_59383_ _59381_/X _86050_/Q _59382_/X _59383_/Y sky130_fd_sc_hd__o21ai_4
X_71661_ _58518_/Y _71649_/X _71660_/Y _83421_/D sky130_fd_sc_hd__o21ai_4
X_83647_ _86422_/CLK _70968_/Y _83647_/Q sky130_fd_sc_hd__dfxtp_4
X_56595_ _56595_/A _56595_/B _56596_/A sky130_fd_sc_hd__and2_4
X_80859_ _83974_/CLK _80891_/Q _75032_/B sky130_fd_sc_hd__dfxtp_4
X_73400_ _44581_/Y _73006_/X _73399_/Y _73412_/C sky130_fd_sc_hd__a21o_4
X_70612_ _70611_/X _70620_/C sky130_fd_sc_hd__buf_2
X_58334_ _58334_/A _58334_/X sky130_fd_sc_hd__buf_2
X_55546_ _55543_/X _55545_/X _55516_/X _55546_/X sky130_fd_sc_hd__a21o_4
X_43560_ _53443_/A _43560_/X sky130_fd_sc_hd__buf_2
X_74380_ _83078_/Q _74377_/X _74379_/Y _74380_/Y sky130_fd_sc_hd__o21ai_4
X_86366_ _83716_/CLK _86366_/D _86366_/Q sky130_fd_sc_hd__dfxtp_4
X_40772_ _40771_/X _40754_/X _88338_/Q _40756_/X _40772_/X sky130_fd_sc_hd__a2bb2o_4
X_52758_ _52775_/A _52746_/B _52746_/C _52758_/D _52758_/X sky130_fd_sc_hd__and4_4
X_71592_ _70558_/X _71590_/B _71582_/X _71592_/Y sky130_fd_sc_hd__nor3_4
X_83578_ _83313_/CLK _71186_/Y _83578_/Q sky130_fd_sc_hd__dfxtp_4
X_88105_ _87595_/CLK _88105_/D _88105_/Q sky130_fd_sc_hd__dfxtp_4
X_42511_ _42495_/X _42496_/X _40702_/X _87839_/Q _42506_/X _42511_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73331_ _73381_/A _86475_/Q _73331_/X sky130_fd_sc_hd__and2_4
X_85317_ _85317_/CLK _55109_/Y _85317_/Q sky130_fd_sc_hd__dfxtp_4
X_51709_ _52593_/A _51709_/X sky130_fd_sc_hd__buf_2
X_70543_ DATA_TO_HASH[6] _70543_/Y sky130_fd_sc_hd__inv_2
X_82529_ _82529_/CLK _82529_/D _78798_/A sky130_fd_sc_hd__dfxtp_4
X_58265_ _58264_/Y _58268_/B _58265_/Y sky130_fd_sc_hd__nand2_4
X_43491_ _41715_/X _43484_/X _87395_/Q _43485_/X _87395_/D sky130_fd_sc_hd__a2bb2o_4
X_55477_ _55477_/A _85139_/Q _55477_/X sky130_fd_sc_hd__and2_4
X_86297_ _86297_/CLK _49933_/Y _72220_/B sky130_fd_sc_hd__dfxtp_4
X_52689_ _52770_/A _52694_/B sky130_fd_sc_hd__buf_2
X_45230_ _56124_/C _45194_/X _45229_/X _45230_/X sky130_fd_sc_hd__o21a_4
X_57216_ _57215_/X _57665_/A _57196_/Y _57216_/Y sky130_fd_sc_hd__nand3_4
X_76050_ _81339_/Q _76041_/B _76050_/Y sky130_fd_sc_hd__nand2_4
X_42442_ _40538_/X _42434_/X _87862_/Q _42435_/X _87862_/D sky130_fd_sc_hd__a2bb2o_4
X_88036_ _88036_/CLK _42101_/Y _88036_/Q sky130_fd_sc_hd__dfxtp_4
X_54428_ _54401_/A _54429_/C sky130_fd_sc_hd__buf_2
X_73262_ _73262_/A _73262_/X sky130_fd_sc_hd__buf_2
X_85248_ _85248_/CLK _85248_/D _55976_/B sky130_fd_sc_hd__dfxtp_4
X_70474_ _58350_/Y _70458_/X _70473_/Y _70474_/Y sky130_fd_sc_hd__o21ai_4
X_58196_ _58196_/A _58196_/Y sky130_fd_sc_hd__inv_2
X_75001_ _75001_/A _75000_/X _75001_/Y sky130_fd_sc_hd__nand2_4
X_72213_ _83274_/Q _72115_/X _72206_/X _72212_/X _72213_/Y sky130_fd_sc_hd__a2bb2oi_4
X_45161_ _45237_/A _45161_/X sky130_fd_sc_hd__buf_2
X_57147_ _57121_/X _57145_/Y _57146_/Y _57147_/X sky130_fd_sc_hd__a21bo_4
X_42373_ _50523_/A _42373_/X sky130_fd_sc_hd__buf_2
X_54359_ _54356_/Y _54338_/X _54358_/X _85457_/D sky130_fd_sc_hd__a21oi_4
X_73193_ _73193_/A _73193_/X sky130_fd_sc_hd__buf_2
X_85179_ _85277_/CLK _85179_/D _55931_/B sky130_fd_sc_hd__dfxtp_4
X_44112_ _44111_/X _44112_/X sky130_fd_sc_hd__buf_2
X_41324_ _41143_/A _41324_/X sky130_fd_sc_hd__buf_2
X_72144_ _59346_/X _85343_/Q _72120_/X _72144_/X sky130_fd_sc_hd__o21a_4
X_45092_ _45089_/Y _45091_/Y _45063_/X _45092_/X sky130_fd_sc_hd__a21o_4
X_57078_ _45842_/Y _56943_/X _57076_/X _57077_/Y _85092_/D sky130_fd_sc_hd__a22oi_4
X_48920_ _48920_/A _48920_/Y sky130_fd_sc_hd__inv_2
X_44043_ _55133_/A _44043_/X sky130_fd_sc_hd__buf_2
X_56029_ _56169_/A _56029_/X sky130_fd_sc_hd__buf_2
X_79740_ _64997_/C _72286_/Y _79739_/Y _79740_/X sky130_fd_sc_hd__o21a_4
X_41255_ _41143_/A _41255_/X sky130_fd_sc_hd__buf_2
X_72075_ _72075_/A _53902_/B _72075_/Y sky130_fd_sc_hd__nand2_4
X_76952_ _76948_/Y _76952_/B _76957_/A sky130_fd_sc_hd__nand2_4
X_71026_ _71026_/A _71030_/C sky130_fd_sc_hd__buf_2
X_75903_ _75903_/A _84373_/Q _75903_/X sky130_fd_sc_hd__xor2_4
X_48851_ _48851_/A _48851_/B _48851_/Y sky130_fd_sc_hd__nand2_4
X_79671_ _79671_/A _84245_/Q _79677_/B sky130_fd_sc_hd__xor2_4
X_41186_ _41186_/A _41197_/B sky130_fd_sc_hd__buf_2
X_76883_ _76873_/Y _76874_/Y _76882_/Y _76888_/C sky130_fd_sc_hd__o21a_4
X_47802_ _81220_/Q _47803_/A sky130_fd_sc_hd__inv_2
X_78622_ _78640_/C _78621_/Y _78626_/A sky130_fd_sc_hd__nand2_4
X_75834_ _75821_/B _75821_/A _75810_/C _75810_/B _75833_/Y _75834_/X
+ sky130_fd_sc_hd__o41a_4
X_48782_ _48837_/A _48793_/A sky130_fd_sc_hd__buf_2
X_45994_ _45980_/A _45994_/X sky130_fd_sc_hd__buf_2
X_47733_ _83547_/Q _54907_/B sky130_fd_sc_hd__inv_2
X_59719_ _59713_/Y _59688_/X _59689_/Y _59717_/Y _59718_/Y _59719_/Y
+ sky130_fd_sc_hd__a41oi_4
X_78553_ _78554_/A _78554_/B _78552_/Y _78557_/B sky130_fd_sc_hd__o21a_4
X_44945_ _45827_/B _44945_/X sky130_fd_sc_hd__buf_2
X_75765_ _75759_/B _75759_/A _75764_/Y _75765_/Y sky130_fd_sc_hd__a21oi_4
X_72977_ _42002_/Y _72771_/A _72889_/X _72976_/Y _72977_/X sky130_fd_sc_hd__a211o_4
X_60991_ _60961_/X _60987_/Y _60935_/X _60989_/X _60990_/X _84544_/D
+ sky130_fd_sc_hd__o41a_4
X_77504_ _77486_/Y _77487_/Y _77488_/Y _77512_/A sky130_fd_sc_hd__o21a_4
Xclkbuf_10_291_0_CLK clkbuf_9_145_0_CLK/X _84360_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_7_103_0_CLK clkbuf_6_51_0_CLK/X clkbuf_8_207_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_74716_ _74716_/A _71846_/A _70758_/C _70730_/X _74716_/X sky130_fd_sc_hd__and4_4
X_62730_ _62847_/A _62731_/A sky130_fd_sc_hd__buf_2
X_47664_ _47655_/A _47692_/B _47692_/C _53177_/D _47664_/X sky130_fd_sc_hd__and4_4
X_71928_ _74527_/A _70979_/C _71940_/C _71928_/D _71928_/Y sky130_fd_sc_hd__nand4_4
X_78484_ _78472_/A _82670_/D _78484_/Y sky130_fd_sc_hd__nand2_4
X_44876_ _56287_/C _44874_/X _44875_/X _44876_/X sky130_fd_sc_hd__o21a_4
X_75696_ _75696_/A _75695_/Y _75696_/X sky130_fd_sc_hd__xor2_4
X_49403_ _49410_/A _51791_/B _49403_/Y sky130_fd_sc_hd__nand2_4
X_46615_ _46614_/X _46647_/B sky130_fd_sc_hd__buf_2
X_77435_ _77416_/A _77435_/Y sky130_fd_sc_hd__inv_2
X_43827_ _41130_/X _43817_/X _87248_/Q _43818_/X _43827_/X sky130_fd_sc_hd__a2bb2o_4
X_62661_ _62678_/A _60273_/X _61744_/X _62661_/Y sky130_fd_sc_hd__nand3_4
X_74647_ _74642_/X _45527_/A _74647_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_73_0_CLK clkbuf_9_36_0_CLK/X _86869_/CLK sky130_fd_sc_hd__clkbuf_1
X_47595_ _47595_/A _47595_/B _47595_/C _53139_/D _47595_/X sky130_fd_sc_hd__and4_4
X_71859_ _71859_/A _71857_/B _71851_/X _71857_/D _71859_/Y sky130_fd_sc_hd__nor4_4
X_64400_ _63562_/A _61226_/X _64400_/Y sky130_fd_sc_hd__nor2_4
X_61612_ _84842_/Q _61323_/B _61613_/A sky130_fd_sc_hd__or2_4
X_49334_ _48163_/X _49334_/X sky130_fd_sc_hd__buf_2
X_46546_ _54069_/B _50858_/B sky130_fd_sc_hd__buf_2
X_65380_ _65607_/A _65548_/B sky130_fd_sc_hd__buf_2
X_77366_ _77353_/A _82091_/D _77360_/C _77387_/A sky130_fd_sc_hd__a21boi_4
X_43758_ _43757_/Y _87281_/D sky130_fd_sc_hd__inv_2
X_62592_ _62585_/X _62589_/Y _62591_/X _84870_/Q _62572_/X _62592_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74578_ _74575_/X _74569_/X _56073_/Y _74570_/X _74578_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_7_118_0_CLK clkbuf_6_59_0_CLK/X clkbuf_8_237_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_79105_ _82833_/Q _82545_/Q _82529_/D sky130_fd_sc_hd__xor2_4
X_64331_ _59399_/A _64316_/B _64331_/Y sky130_fd_sc_hd__nor2_4
X_76317_ _76313_/X _76317_/B _76325_/A sky130_fd_sc_hd__xnor2_4
X_42709_ _42709_/A _42709_/Y sky130_fd_sc_hd__inv_2
X_49265_ _49261_/A _49265_/B _49265_/Y sky130_fd_sc_hd__nand2_4
X_61543_ _58438_/A _61563_/B _61563_/C _61514_/D _61544_/A sky130_fd_sc_hd__nand4_4
X_73529_ _72730_/X _73529_/X sky130_fd_sc_hd__buf_2
X_46477_ _52522_/B _50827_/B sky130_fd_sc_hd__buf_2
X_77297_ _77285_/C _77279_/Y _77297_/Y sky130_fd_sc_hd__nand2_4
X_43689_ _40802_/X _43685_/X _72947_/A _43686_/X _43689_/X sky130_fd_sc_hd__a2bb2o_4
X_48216_ _86554_/Q _48188_/X _48215_/Y _48216_/Y sky130_fd_sc_hd__o21ai_4
X_67050_ _87423_/Q _66997_/X _66998_/X _67049_/X _67050_/X sky130_fd_sc_hd__a211o_4
X_79036_ _79031_/B _79029_/Y _79037_/C sky130_fd_sc_hd__nand2_4
X_45428_ _45424_/X _45427_/X _45361_/X _45428_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_10_88_0_CLK clkbuf_9_44_0_CLK/X _84408_/CLK sky130_fd_sc_hd__clkbuf_1
X_64262_ _64248_/A _64248_/B _84717_/Q _64262_/X sky130_fd_sc_hd__and3_4
X_76248_ _81641_/Q _76248_/Y sky130_fd_sc_hd__inv_2
X_61474_ _61413_/A _61518_/A sky130_fd_sc_hd__buf_2
X_49196_ _53936_/B _50721_/B sky130_fd_sc_hd__buf_2
X_66001_ _65700_/X _65999_/Y _66000_/Y _66001_/Y sky130_fd_sc_hd__o21ai_4
X_63213_ _60452_/X _63288_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_234_0_CLK clkbuf_8_235_0_CLK/A clkbuf_9_469_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_48147_ _48134_/X _82915_/Q _48146_/X _48148_/B sky130_fd_sc_hd__o21ai_4
X_60425_ _60420_/A _60441_/B sky130_fd_sc_hd__buf_2
X_45359_ _56454_/C _45326_/X _45358_/X _45359_/Y sky130_fd_sc_hd__o21ai_4
X_64193_ _64189_/Y _64190_/Y _64191_/Y _64193_/D _64193_/X sky130_fd_sc_hd__and4_4
X_76179_ _76174_/Y _76177_/Y _76178_/Y _76179_/Y sky130_fd_sc_hd__a21oi_4
X_63144_ _60503_/X _63144_/X sky130_fd_sc_hd__buf_2
X_48078_ _48075_/X _82922_/Q _48077_/X _48079_/B sky130_fd_sc_hd__o21ai_4
X_60356_ _60355_/Y _60356_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_11_0_CLK clkbuf_9_5_0_CLK/X _85244_/CLK sky130_fd_sc_hd__clkbuf_1
X_47029_ _47029_/A _47029_/B _47029_/C _52811_/D _47029_/X sky130_fd_sc_hd__and4_4
Xclkbuf_9_350_0_CLK clkbuf_9_351_0_CLK/A clkbuf_9_350_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_67952_ _87961_/Q _67950_/X _67879_/X _67951_/X _67952_/X sky130_fd_sc_hd__a211o_4
X_63075_ _63038_/A _64284_/B _63085_/C _63085_/D _63075_/X sky130_fd_sc_hd__and4_4
X_79938_ _79936_/Y _79937_/Y _79942_/A sky130_fd_sc_hd__nand2_4
X_60287_ _79797_/A _59822_/X _60284_/Y _60286_/X _60287_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_8_249_0_CLK clkbuf_8_249_0_CLK/A clkbuf_9_499_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_244_0_CLK clkbuf_9_122_0_CLK/X _84583_/CLK sky130_fd_sc_hd__clkbuf_1
X_50040_ _50050_/A _50040_/B _51750_/C _53253_/D _50040_/X sky130_fd_sc_hd__and4_4
X_66903_ _66902_/X _86792_/Q _66903_/X sky130_fd_sc_hd__and2_4
X_62026_ _61558_/B _61995_/X _62010_/X _62011_/X _62026_/Y sky130_fd_sc_hd__nand4_4
X_67883_ _87388_/Q _67834_/X _67835_/X _67882_/X _67883_/X sky130_fd_sc_hd__a211o_4
X_79869_ _64663_/C _83279_/Q _79869_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_874_0_CLK clkbuf_9_437_0_CLK/X _86235_/CLK sky130_fd_sc_hd__clkbuf_1
X_81900_ _82104_/CLK _77375_/X _82276_/D sky130_fd_sc_hd__dfxtp_4
X_69622_ _69908_/A _69622_/B _69622_/Y sky130_fd_sc_hd__nor2_4
X_66834_ _66717_/A _66834_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_26_0_CLK clkbuf_9_13_0_CLK/X _85138_/CLK sky130_fd_sc_hd__clkbuf_1
X_82880_ _82368_/CLK _82472_/Q _82880_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_365_0_CLK clkbuf_9_365_0_CLK/A clkbuf_9_365_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_69553_ _69956_/A _69553_/B _69553_/X sky130_fd_sc_hd__and2_4
X_81831_ _81859_/CLK _81863_/Q _77294_/A sky130_fd_sc_hd__dfxtp_4
X_66765_ _66664_/X _66765_/B _66765_/X sky130_fd_sc_hd__and2_4
X_51991_ _73827_/B _51960_/X _51990_/Y _51991_/Y sky130_fd_sc_hd__o21ai_4
X_63977_ _63975_/X _63913_/X _63976_/Y _63977_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_259_0_CLK clkbuf_9_129_0_CLK/X _84877_/CLK sky130_fd_sc_hd__clkbuf_1
X_68504_ _68757_/A _68504_/X sky130_fd_sc_hd__buf_2
X_53730_ _53755_/A _53750_/A sky130_fd_sc_hd__buf_2
X_65716_ _65623_/X _86190_/Q _65517_/X _65715_/X _65716_/X sky130_fd_sc_hd__a211o_4
X_84550_ _84293_/CLK _60932_/Y _60931_/C sky130_fd_sc_hd__dfxtp_4
X_50942_ _50940_/Y _50928_/X _50941_/X _50942_/Y sky130_fd_sc_hd__a21oi_4
X_62928_ _60337_/A _62949_/B _62928_/C _62928_/D _62928_/Y sky130_fd_sc_hd__nand4_4
X_81762_ _86582_/CLK _81762_/D _81762_/Q sky130_fd_sc_hd__dfxtp_4
X_69484_ _69481_/X _69483_/X _69385_/X _69484_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_10_889_0_CLK clkbuf_9_444_0_CLK/X _86045_/CLK sky130_fd_sc_hd__clkbuf_1
X_66696_ _66693_/X _66695_/X _66696_/Y sky130_fd_sc_hd__nand2_4
X_83501_ _83498_/CLK _71433_/X _83501_/Q sky130_fd_sc_hd__dfxtp_4
X_68435_ _83975_/Q _68338_/X _68434_/X _68435_/X sky130_fd_sc_hd__a21bo_4
X_80713_ _80679_/CLK _75899_/X _80681_/D sky130_fd_sc_hd__dfxtp_4
X_53661_ _53661_/A _53755_/A sky130_fd_sc_hd__buf_2
X_65647_ _64990_/X _65647_/B _64993_/X _65647_/Y sky130_fd_sc_hd__nand3_4
X_84481_ _84481_/CLK _61435_/Y _61434_/C sky130_fd_sc_hd__dfxtp_4
X_50873_ _50871_/Y _50243_/X _50872_/Y _50873_/Y sky130_fd_sc_hd__a21boi_4
X_62859_ _62681_/X _62859_/X sky130_fd_sc_hd__buf_2
X_81693_ _81269_/CLK _80211_/X _81693_/Q sky130_fd_sc_hd__dfxtp_4
X_55400_ _55400_/A _55400_/Y sky130_fd_sc_hd__inv_2
X_86220_ _86570_/CLK _86220_/D _86220_/Q sky130_fd_sc_hd__dfxtp_4
X_52612_ _52624_/A _46685_/A _52612_/Y sky130_fd_sc_hd__nand2_4
X_83432_ _83431_/CLK _71633_/Y _83432_/Q sky130_fd_sc_hd__dfxtp_4
X_56380_ _56005_/X _56378_/X _56379_/Y _56380_/Y sky130_fd_sc_hd__o21ai_4
X_80644_ _80644_/A _74708_/Y DATA_FROM_HASH[1] sky130_fd_sc_hd__ebufn_2
X_68366_ _57803_/A _68366_/X sky130_fd_sc_hd__buf_2
X_53592_ _53589_/Y _53574_/X _53591_/Y _85607_/D sky130_fd_sc_hd__a21boi_4
X_65578_ _65731_/A _73040_/B _65578_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_812_0_CLK clkbuf_9_406_0_CLK/X _82859_/CLK sky130_fd_sc_hd__clkbuf_1
X_55331_ _55329_/Y _55330_/X _55356_/A sky130_fd_sc_hd__nand2_4
X_67317_ _67248_/A _87668_/Q _67317_/X sky130_fd_sc_hd__and2_4
X_86151_ _85542_/CLK _86151_/D _86151_/Q sky130_fd_sc_hd__dfxtp_4
X_52543_ _52542_/X _50850_/B _52543_/Y sky130_fd_sc_hd__nand2_4
XPHY_206 sky130_fd_sc_hd__decap_3
X_64529_ _64522_/Y _64528_/X _60074_/X _64529_/Y sky130_fd_sc_hd__o21ai_4
X_83363_ _83362_/CLK _83363_/D _83363_/Q sky130_fd_sc_hd__dfxtp_4
X_80575_ _80570_/Y _80574_/Y _82268_/D sky130_fd_sc_hd__xor2_4
X_68297_ _68272_/X _67815_/Y _68287_/X _68296_/Y _68297_/X sky130_fd_sc_hd__a211o_4
XPHY_217 sky130_fd_sc_hd__decap_3
XPHY_228 sky130_fd_sc_hd__decap_3
XPHY_239 sky130_fd_sc_hd__decap_3
X_85102_ _85039_/CLK _85102_/D _85102_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_303_0_CLK clkbuf_9_303_0_CLK/A clkbuf_9_303_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_58050_ _57983_/X _85385_/Q _58049_/X _58050_/Y sky130_fd_sc_hd__o21ai_4
X_82314_ _81179_/CLK _77060_/B _82314_/Q sky130_fd_sc_hd__dfxtp_4
X_67248_ _67248_/A _67248_/B _67248_/X sky130_fd_sc_hd__and2_4
X_55262_ _82985_/Q _44059_/A _55140_/X _55261_/X _55264_/C sky130_fd_sc_hd__a211o_4
X_86082_ _85764_/CLK _51057_/Y _86082_/Q sky130_fd_sc_hd__dfxtp_4
X_52474_ _52468_/A _53993_/B _52474_/Y sky130_fd_sc_hd__nand2_4
X_83294_ _85536_/CLK _83294_/D _83294_/Q sky130_fd_sc_hd__dfxtp_4
X_57001_ _57001_/A _85103_/D sky130_fd_sc_hd__inv_2
X_54213_ _54208_/X _54191_/B _54209_/C _53048_/D _54213_/X sky130_fd_sc_hd__and4_4
X_85033_ _83335_/CLK _85033_/D _85033_/Q sky130_fd_sc_hd__dfxtp_4
X_51425_ _86012_/Q _51402_/X _51424_/Y _51425_/Y sky130_fd_sc_hd__o21ai_4
X_82245_ _82263_/CLK _80322_/X _82245_/Q sky130_fd_sc_hd__dfxtp_4
X_55193_ _82989_/Q _55190_/X _44095_/A _55192_/X _55193_/X sky130_fd_sc_hd__a211o_4
X_67179_ _67133_/A _67179_/B _67179_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_827_0_CLK clkbuf_9_413_0_CLK/X _82369_/CLK sky130_fd_sc_hd__clkbuf_1
X_54144_ _53436_/X _54144_/X sky130_fd_sc_hd__buf_2
X_51356_ _51306_/X _51356_/B _51356_/X sky130_fd_sc_hd__and2_4
X_70190_ _70200_/A _70200_/B _83203_/Q _70200_/D _70190_/X sky130_fd_sc_hd__and4_4
X_82176_ _84115_/CLK _84168_/Q _82176_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_318_0_CLK clkbuf_9_318_0_CLK/A clkbuf_9_318_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_50307_ _86226_/Q _50238_/X _50306_/Y _50307_/Y sky130_fd_sc_hd__o21ai_4
X_81127_ _81125_/CLK _81127_/D _40732_/A sky130_fd_sc_hd__dfxtp_4
X_58952_ _58941_/A _86371_/Q _58952_/Y sky130_fd_sc_hd__nor2_4
X_54075_ _53801_/B _54075_/B _54075_/Y sky130_fd_sc_hd__nand2_4
X_51287_ _51296_/A _50777_/B _51287_/Y sky130_fd_sc_hd__nand2_4
X_86984_ _86984_/CLK _86984_/D _44727_/A sky130_fd_sc_hd__dfxtp_4
X_41040_ _40999_/A _41040_/X sky130_fd_sc_hd__buf_2
X_53026_ _85710_/Q _53010_/X _53025_/Y _53026_/Y sky130_fd_sc_hd__o21ai_4
X_57903_ _58605_/A _57903_/X sky130_fd_sc_hd__buf_2
X_50238_ _50464_/A _50238_/X sky130_fd_sc_hd__buf_2
X_85935_ _86096_/CLK _51852_/Y _85935_/Q sky130_fd_sc_hd__dfxtp_4
X_81058_ _81059_/CLK _81090_/Q _81058_/Q sky130_fd_sc_hd__dfxtp_4
X_58883_ _59053_/A _58883_/X sky130_fd_sc_hd__buf_2
Xclkbuf_5_3_0_CLK clkbuf_5_2_0_CLK/A clkbuf_6_7_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_72900_ _72892_/B _72900_/X sky130_fd_sc_hd__buf_2
X_80009_ _80000_/A _79999_/X _80011_/B sky130_fd_sc_hd__or2_4
X_57834_ _57801_/X _57832_/Y _57833_/Y _57822_/X _57809_/X _57834_/X
+ sky130_fd_sc_hd__o32a_4
X_50169_ _50169_/A _50169_/B _50169_/Y sky130_fd_sc_hd__nand2_4
X_73880_ _73829_/X _66097_/B _73880_/X sky130_fd_sc_hd__and2_4
X_85866_ _85866_/CLK _85866_/D _85866_/Q sky130_fd_sc_hd__dfxtp_4
X_87605_ _87348_/CLK _87605_/D _67285_/B sky130_fd_sc_hd__dfxtp_4
X_72831_ _72831_/A _72924_/B _72831_/Y sky130_fd_sc_hd__nor2_4
X_84817_ _84815_/CLK _84817_/D _84817_/Q sky130_fd_sc_hd__dfxtp_4
X_57765_ _57760_/X _85405_/Q _57764_/X _57765_/Y sky130_fd_sc_hd__o21ai_4
X_42991_ _42984_/X _42985_/X _40491_/X _87615_/Q _42463_/A _42992_/A
+ sky130_fd_sc_hd__o32ai_4
X_54977_ _85342_/Q _54967_/X _54976_/Y _54977_/Y sky130_fd_sc_hd__o21ai_4
X_85797_ _85800_/CLK _85797_/D _65335_/B sky130_fd_sc_hd__dfxtp_4
X_59504_ _59504_/A _59504_/Y sky130_fd_sc_hd__inv_2
X_44730_ _44730_/A _44730_/Y sky130_fd_sc_hd__inv_2
X_56716_ _56715_/Y _57416_/C sky130_fd_sc_hd__buf_2
X_75550_ _75551_/B _75550_/Y sky130_fd_sc_hd__inv_2
X_87536_ _88087_/CLK _43210_/X _87536_/Q sky130_fd_sc_hd__dfxtp_4
X_41942_ _41937_/X _41919_/X _40678_/X _41941_/Y _41939_/X _88099_/D
+ sky130_fd_sc_hd__o32ai_4
X_53928_ _85540_/Q _53921_/X _53927_/Y _53928_/Y sky130_fd_sc_hd__o21ai_4
X_72762_ _48357_/Y _72762_/B _72762_/X sky130_fd_sc_hd__xor2_4
X_84748_ _84760_/CLK _59363_/Y _84748_/Q sky130_fd_sc_hd__dfxtp_4
X_57696_ _58805_/A _57696_/X sky130_fd_sc_hd__buf_2
X_74501_ _74501_/A _74501_/B _74501_/C _74501_/X sky130_fd_sc_hd__and3_4
X_71713_ _70700_/A _70700_/B _71713_/Y sky130_fd_sc_hd__nand2_4
X_59435_ _59417_/X _83342_/Q _59434_/Y _84734_/D sky130_fd_sc_hd__o21a_4
X_56647_ _45893_/C _44292_/A _46173_/X _56647_/A4 _56646_/Y _56647_/X
+ sky130_fd_sc_hd__a41o_4
X_44661_ _44658_/X _44659_/X _41086_/X _87012_/Q _44660_/X _44662_/A
+ sky130_fd_sc_hd__o32ai_4
X_75481_ _75477_/X _75478_/Y _75480_/Y _75481_/X sky130_fd_sc_hd__a21o_4
X_87467_ _86934_/CLK _87467_/D _87467_/Q sky130_fd_sc_hd__dfxtp_4
X_41873_ _57491_/B _50731_/A _40560_/X _73552_/A _41872_/X _41873_/Y
+ sky130_fd_sc_hd__o32ai_4
X_53859_ _53857_/Y _53838_/X _53858_/Y _85554_/D sky130_fd_sc_hd__a21boi_4
X_72693_ _72697_/A _72697_/B _55423_/B _72693_/Y sky130_fd_sc_hd__nand3_4
X_84679_ _84396_/CLK _84679_/D _59982_/C sky130_fd_sc_hd__dfxtp_4
X_46400_ _46259_/A _46401_/A sky130_fd_sc_hd__buf_2
X_77220_ _82112_/Q _77220_/B _77220_/X sky130_fd_sc_hd__xor2_4
X_43612_ _40604_/X _43609_/X _68468_/B _43611_/X _43613_/A sky130_fd_sc_hd__a2bb2o_4
X_86418_ _85516_/CLK _49284_/Y _86418_/Q sky130_fd_sc_hd__dfxtp_4
X_74432_ _74429_/Y _74430_/X _74431_/X _74432_/Y sky130_fd_sc_hd__a21oi_4
X_40824_ _82869_/Q _40847_/B _40824_/X sky130_fd_sc_hd__or2_4
X_47380_ _47380_/A _47408_/B _47377_/X _53015_/D _47380_/X sky130_fd_sc_hd__and4_4
X_59366_ _59292_/X _85635_/Q _59365_/X _59366_/X sky130_fd_sc_hd__o21a_4
X_71644_ _71637_/A _71232_/B _71644_/C _71644_/Y sky130_fd_sc_hd__nand3_4
X_44592_ _44591_/Y _44592_/Y sky130_fd_sc_hd__inv_2
X_56578_ _56577_/Y _56578_/X sky130_fd_sc_hd__buf_2
X_87398_ _87150_/CLK _87398_/D _87398_/Q sky130_fd_sc_hd__dfxtp_4
X_46331_ _46288_/A _52454_/B _46331_/Y sky130_fd_sc_hd__nand2_4
X_58317_ _58317_/A _58326_/B _58317_/Y sky130_fd_sc_hd__nand2_4
X_77151_ _77151_/A _77151_/B _77152_/B sky130_fd_sc_hd__xnor2_4
X_43543_ _43542_/X _43523_/X _40440_/X _87367_/Q _43528_/X _43544_/A
+ sky130_fd_sc_hd__o32ai_4
X_55529_ _55534_/A _55529_/B _55529_/X sky130_fd_sc_hd__and2_4
X_74363_ _72068_/A _48357_/Y _74363_/Y sky130_fd_sc_hd__nand2_4
X_86349_ _86351_/CLK _49647_/Y _59244_/B sky130_fd_sc_hd__dfxtp_4
X_40755_ _40755_/A _40756_/A sky130_fd_sc_hd__buf_2
X_59297_ _59297_/A _59297_/X sky130_fd_sc_hd__buf_2
X_71575_ _71556_/Y _58336_/B _71574_/Y _83451_/D sky130_fd_sc_hd__a21o_4
X_76102_ _76094_/A _76099_/B _76093_/A _76102_/Y sky130_fd_sc_hd__o21ai_4
X_49050_ _50645_/A _50645_/B _48917_/X _49050_/X sky130_fd_sc_hd__o21a_4
X_73314_ _73301_/X _73303_/X _73313_/X _73314_/X sky130_fd_sc_hd__a21o_4
X_70526_ _70526_/A _74533_/A _70962_/C _70526_/Y sky130_fd_sc_hd__nand3_4
X_46262_ _46348_/A _46262_/X sky130_fd_sc_hd__buf_2
X_77082_ _81998_/Q _81910_/Q _77096_/A sky130_fd_sc_hd__xor2_4
X_58248_ _58248_/A _58248_/B _58248_/Y sky130_fd_sc_hd__nor2_4
X_43474_ _43474_/A _87404_/D sky130_fd_sc_hd__inv_2
X_74294_ _70275_/C _74288_/X _74293_/Y _74294_/X sky130_fd_sc_hd__a21bo_4
X_40686_ _40686_/A _40835_/A sky130_fd_sc_hd__buf_2
X_48001_ _48731_/A _48004_/A sky130_fd_sc_hd__buf_2
X_45213_ _45208_/Y _45211_/Y _45212_/X _45213_/X sky130_fd_sc_hd__a21o_4
X_76033_ _81714_/D _76042_/B _76047_/A sky130_fd_sc_hd__xor2_4
X_88019_ _87249_/CLK _88019_/D _88019_/Q sky130_fd_sc_hd__dfxtp_4
X_42425_ _40497_/X _42414_/X _87870_/Q _42415_/X _87870_/D sky130_fd_sc_hd__a2bb2o_4
X_73245_ _73243_/X _73244_/Y _73221_/X _73245_/Y sky130_fd_sc_hd__a21oi_4
X_46193_ _46207_/B _46217_/C _46222_/B sky130_fd_sc_hd__and2_4
X_70457_ _70455_/Y _71462_/B _70457_/X sky130_fd_sc_hd__and2_4
X_58179_ _64292_/A _58217_/B _58179_/Y sky130_fd_sc_hd__nand2_4
X_60210_ _60189_/A _60309_/D sky130_fd_sc_hd__buf_2
X_45144_ _45219_/A _45144_/X sky130_fd_sc_hd__buf_2
X_42356_ _42290_/A _42356_/X sky130_fd_sc_hd__buf_2
X_61190_ _61188_/B _61190_/X sky130_fd_sc_hd__buf_2
X_73176_ _69776_/Y _73195_/A _72889_/X _73175_/Y _73176_/X sky130_fd_sc_hd__a211o_4
X_70388_ _70997_/A _74527_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_80_0_CLK clkbuf_7_81_0_CLK/A clkbuf_7_80_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_41307_ _41181_/A _41307_/X sky130_fd_sc_hd__buf_2
X_72127_ _83281_/Q _72115_/X _72119_/X _72126_/X _72127_/Y sky130_fd_sc_hd__a2bb2oi_4
X_60141_ _59913_/X _60011_/X _60100_/Y _60141_/Y sky130_fd_sc_hd__a21boi_4
X_49952_ _46308_/A _49973_/A sky130_fd_sc_hd__buf_2
X_45075_ _56221_/C _45073_/X _45074_/X _45075_/Y sky130_fd_sc_hd__o21ai_4
X_42287_ _42287_/A _87939_/D sky130_fd_sc_hd__inv_2
X_77984_ _77984_/A _77983_/Y _77984_/Y sky130_fd_sc_hd__nand2_4
X_48903_ _48903_/A _48908_/A sky130_fd_sc_hd__buf_2
X_44026_ _44006_/X _44025_/X _44026_/Y sky130_fd_sc_hd__nand2_4
X_79723_ _79721_/X _79722_/X _79724_/B sky130_fd_sc_hd__xnor2_4
X_41238_ _41237_/Y _88252_/D sky130_fd_sc_hd__inv_2
X_60072_ _60056_/A _59931_/A _60072_/Y sky130_fd_sc_hd__nor2_4
X_72058_ _83293_/Q _72001_/X _72057_/Y _72058_/Y sky130_fd_sc_hd__o21ai_4
X_76935_ _76918_/A _76918_/B _76906_/A _76934_/Y _76935_/X sky130_fd_sc_hd__a2bb2o_4
X_49883_ _58135_/B _49880_/X _49882_/Y _49883_/Y sky130_fd_sc_hd__o21ai_4
X_63900_ _58511_/A _63900_/B _63900_/C _63900_/D _63903_/B sky130_fd_sc_hd__nand4_4
X_71009_ _49320_/B _70983_/A _71008_/Y _71009_/Y sky130_fd_sc_hd__o21ai_4
X_48834_ _52218_/A _48849_/B _48849_/C _48834_/X sky130_fd_sc_hd__and3_4
X_79654_ _79651_/X _79653_/Y _79654_/Y sky130_fd_sc_hd__xnor2_4
X_41169_ _41168_/Y _41169_/X sky130_fd_sc_hd__buf_2
X_64880_ _64876_/X _64712_/B _64879_/X _64880_/Y sky130_fd_sc_hd__nand3_4
X_76866_ _76849_/A _76862_/A _76866_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_7_95_0_CLK clkbuf_7_95_0_CLK/A clkbuf_7_95_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_78605_ _78601_/Y _78581_/B _78604_/X _78605_/Y sky130_fd_sc_hd__o21ai_4
X_63831_ _63831_/A _64272_/A _63765_/C _63831_/X sky130_fd_sc_hd__and3_4
X_75817_ _75817_/A _75817_/B _75817_/Y sky130_fd_sc_hd__xnor2_4
X_48765_ _48790_/A _48786_/C sky130_fd_sc_hd__buf_2
X_79585_ _84206_/Q _83254_/Q _79585_/Y sky130_fd_sc_hd__nand2_4
X_45977_ _40403_/Y _45974_/X _86831_/Q _45976_/X _45977_/X sky130_fd_sc_hd__a2bb2o_4
X_76797_ _76773_/Y _81360_/D sky130_fd_sc_hd__inv_2
X_47716_ _47716_/A _54898_/B sky130_fd_sc_hd__inv_2
X_66550_ _69457_/A _66550_/X sky130_fd_sc_hd__buf_2
X_78536_ _78534_/Y _78536_/B _78536_/X sky130_fd_sc_hd__xor2_4
X_44928_ _56198_/C _44911_/X _44927_/X _44928_/Y sky130_fd_sc_hd__o21ai_4
X_63762_ _61330_/X _63781_/B _63781_/C _63761_/X _63762_/Y sky130_fd_sc_hd__nand4_4
X_75748_ _81013_/Q _75748_/B _75748_/X sky130_fd_sc_hd__xor2_4
X_60974_ _60928_/X _64191_/D sky130_fd_sc_hd__buf_2
X_48696_ _86499_/Q _48669_/X _48695_/Y _48696_/Y sky130_fd_sc_hd__o21ai_4
X_65501_ _65184_/A _65501_/B _65501_/X sky130_fd_sc_hd__and2_4
X_62713_ _62949_/B _62713_/X sky130_fd_sc_hd__buf_2
X_47647_ _83628_/Q _54859_/B sky130_fd_sc_hd__inv_2
X_66481_ _65215_/X _66476_/B _65217_/X _66481_/Y sky130_fd_sc_hd__nand3_4
X_78467_ _78475_/B _78453_/B _78466_/X _78467_/Y sky130_fd_sc_hd__o21ai_4
X_44859_ _44857_/X _44844_/X _41772_/X _67988_/B _44858_/X _44860_/A
+ sky130_fd_sc_hd__o32ai_4
X_63693_ _63688_/Y _63679_/X _63692_/Y _84301_/D sky130_fd_sc_hd__a21oi_4
X_75679_ _75666_/A _75674_/A _75679_/X sky130_fd_sc_hd__and2_4
X_68220_ _68160_/A _68220_/X sky130_fd_sc_hd__buf_2
X_65432_ _64595_/X _65340_/X _64604_/X _65432_/Y sky130_fd_sc_hd__nand3_4
X_77418_ _77381_/A _77382_/X _77417_/B _77418_/X sky130_fd_sc_hd__a21o_4
X_62644_ _62644_/A _62644_/X sky130_fd_sc_hd__buf_2
X_47578_ _47578_/A _53129_/D sky130_fd_sc_hd__buf_2
X_78398_ _78365_/A _78379_/A _78380_/A _78398_/X sky130_fd_sc_hd__a21o_4
X_49317_ _71959_/A _49317_/X sky130_fd_sc_hd__buf_2
X_68151_ _82066_/D _68140_/X _68150_/X _68151_/X sky130_fd_sc_hd__a21bo_4
X_46529_ _46525_/X _49129_/A _46528_/X _51360_/B sky130_fd_sc_hd__o21ai_4
X_65363_ _65718_/A _65363_/X sky130_fd_sc_hd__buf_2
X_77349_ _77319_/X _77347_/Y _77348_/X _77349_/X sky130_fd_sc_hd__o21a_4
X_62575_ _62573_/Y _62540_/X _62574_/Y _84400_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_7_33_0_CLK clkbuf_6_16_0_CLK/X clkbuf_8_67_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_67102_ _67099_/X _67101_/X _67102_/Y sky130_fd_sc_hd__nand2_4
X_64314_ _64314_/A _64314_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_173_0_CLK clkbuf_7_86_0_CLK/X clkbuf_9_347_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_49248_ _49215_/A _49263_/A sky130_fd_sc_hd__buf_2
X_61526_ _72528_/A _61542_/B sky130_fd_sc_hd__buf_2
X_80360_ _80358_/Y _80360_/B _80350_/B _80361_/B sky130_fd_sc_hd__nand3_4
X_68082_ _68079_/X _68081_/X _68033_/X _68082_/X sky130_fd_sc_hd__a21o_4
X_65294_ _65268_/A _65294_/B _65294_/C _65294_/X sky130_fd_sc_hd__and3_4
X_67033_ _67057_/A _67033_/B _67033_/X sky130_fd_sc_hd__and2_4
X_79019_ _82745_/Q _79019_/B _82713_/D sky130_fd_sc_hd__xor2_4
X_64245_ _64273_/A _64273_/B _63400_/B _64221_/X _64245_/X sky130_fd_sc_hd__and4_4
X_49179_ _49179_/A _49161_/B _49179_/Y sky130_fd_sc_hd__nor2_4
X_61457_ _61454_/X _61455_/X _61456_/Y _61457_/Y sky130_fd_sc_hd__a21oi_4
X_80291_ _84748_/Q _84140_/Q _80292_/B sky130_fd_sc_hd__nand2_4
X_51210_ _51074_/A _51211_/A sky130_fd_sc_hd__buf_2
X_82030_ _81985_/CLK _77843_/B _81998_/D sky130_fd_sc_hd__dfxtp_4
X_60408_ _60408_/A _60406_/X _60408_/C _60408_/X sky130_fd_sc_hd__and3_4
X_52190_ _52210_/A _48561_/B _52190_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_7_48_0_CLK clkbuf_6_24_0_CLK/X clkbuf_8_97_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_64176_ _64174_/X _64129_/X _64175_/Y _64176_/Y sky130_fd_sc_hd__a21oi_4
X_61388_ _61377_/A _61387_/X _61377_/C _61388_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_8_188_0_CLK clkbuf_7_94_0_CLK/X clkbuf_8_188_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_51141_ _51141_/A _51141_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_183_0_CLK clkbuf_9_91_0_CLK/X _83322_/CLK sky130_fd_sc_hd__clkbuf_1
X_63127_ _63127_/A _63113_/B _63103_/C _63092_/D _63127_/X sky130_fd_sc_hd__or4_4
X_60339_ _60317_/A _60319_/X _79658_/A _60339_/Y sky130_fd_sc_hd__nor3_4
X_68984_ _69027_/A _68984_/B _68984_/X sky130_fd_sc_hd__and2_4
X_51072_ _51070_/Y _51065_/X _51071_/X _51072_/Y sky130_fd_sc_hd__a21oi_4
X_67935_ _68479_/A _68028_/A sky130_fd_sc_hd__buf_2
X_63058_ _79467_/A _63008_/X _63057_/Y _63058_/X sky130_fd_sc_hd__a21o_4
X_83981_ _82629_/CLK _83981_/D _82629_/D sky130_fd_sc_hd__dfxtp_4
X_50023_ _50027_/A _53236_/B _50023_/Y sky130_fd_sc_hd__nand2_4
X_54900_ _54900_/A _54910_/B sky130_fd_sc_hd__buf_2
X_62009_ _61549_/X _62007_/X _61967_/C _62008_/X _62015_/B sky130_fd_sc_hd__nand4_4
X_85720_ _85718_/CLK _85720_/D _85720_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_111_0_CLK clkbuf_7_55_0_CLK/X clkbuf_9_222_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_82932_ _82931_/CLK _78261_/X _82932_/Q sky130_fd_sc_hd__dfxtp_4
X_55880_ _45094_/A _55531_/X _55533_/X _55879_/X _55880_/X sky130_fd_sc_hd__a211o_4
X_67866_ _67817_/X _87645_/Q _67866_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_198_0_CLK clkbuf_9_99_0_CLK/X _84273_/CLK sky130_fd_sc_hd__clkbuf_1
X_69605_ _69605_/A _72831_/A _69605_/X sky130_fd_sc_hd__and2_4
X_54831_ _54825_/A _54843_/B _54831_/C _53139_/D _54831_/X sky130_fd_sc_hd__and4_4
X_66817_ _66795_/A _66817_/B _66817_/X sky130_fd_sc_hd__and2_4
X_85651_ _85651_/CLK _53344_/Y _85651_/Q sky130_fd_sc_hd__dfxtp_4
X_82863_ _82859_/CLK _78177_/B _82863_/Q sky130_fd_sc_hd__dfxtp_4
X_67797_ _87456_/Q _67751_/X _67702_/X _67796_/X _67797_/X sky130_fd_sc_hd__a211o_4
X_84602_ _84477_/CLK _60548_/Y _79142_/A sky130_fd_sc_hd__dfxtp_4
X_57550_ _46542_/X _57550_/X sky130_fd_sc_hd__buf_2
X_81814_ _81689_/CLK _81622_/Q _81814_/Q sky130_fd_sc_hd__dfxtp_4
X_69536_ _44022_/X _69536_/B _69536_/X sky130_fd_sc_hd__and2_4
X_88370_ _86982_/CLK _40575_/Y _88370_/Q sky130_fd_sc_hd__dfxtp_4
X_54762_ _54760_/Y _54747_/X _54761_/X _85383_/D sky130_fd_sc_hd__a21oi_4
X_66748_ _66819_/A _86799_/Q _66748_/X sky130_fd_sc_hd__and2_4
X_85582_ _86506_/CLK _53717_/Y _85582_/Q sky130_fd_sc_hd__dfxtp_4
X_51974_ _51971_/Y _51951_/X _51973_/X _85914_/D sky130_fd_sc_hd__a21oi_4
X_82794_ _82797_/CLK _82826_/Q _78418_/A sky130_fd_sc_hd__dfxtp_4
X_56501_ _56510_/A _56507_/B _56501_/C _56501_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_8_126_0_CLK clkbuf_7_63_0_CLK/X clkbuf_9_253_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_87321_ _87577_/CLK _87321_/D _74166_/A sky130_fd_sc_hd__dfxtp_4
X_53713_ _53713_/A _48572_/A _53713_/Y sky130_fd_sc_hd__nand2_4
X_84533_ _84538_/CLK _84533_/D _76981_/A sky130_fd_sc_hd__dfxtp_4
X_50925_ _50922_/Y _50902_/X _50924_/X _86106_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_121_0_CLK clkbuf_9_60_0_CLK/X _84293_/CLK sky130_fd_sc_hd__clkbuf_1
X_81745_ _82642_/CLK _81745_/D _41369_/A sky130_fd_sc_hd__dfxtp_4
X_57481_ _57481_/A _84996_/D sky130_fd_sc_hd__inv_2
X_69467_ _88027_/Q _69424_/X _69465_/X _69466_/X _69467_/X sky130_fd_sc_hd__a211o_4
X_54693_ _54284_/A _54693_/X sky130_fd_sc_hd__buf_2
X_66679_ _66602_/A _86834_/Q _66679_/X sky130_fd_sc_hd__and2_4
X_59220_ _58847_/A _59220_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_751_0_CLK clkbuf_9_375_0_CLK/X _87758_/CLK sky130_fd_sc_hd__clkbuf_1
X_56432_ _56121_/X _56426_/X _56431_/Y _85196_/D sky130_fd_sc_hd__o21ai_4
X_68418_ _69001_/A _68418_/B _68418_/Y sky130_fd_sc_hd__nor2_4
X_87252_ _87766_/CLK _87252_/D _69555_/B sky130_fd_sc_hd__dfxtp_4
X_53644_ _85596_/Q _53610_/X _53643_/Y _53644_/Y sky130_fd_sc_hd__o21ai_4
X_84464_ _84469_/CLK _61635_/Y _79132_/B sky130_fd_sc_hd__dfxtp_4
X_50856_ _50213_/X _50856_/X sky130_fd_sc_hd__buf_2
X_81676_ _81660_/CLK _80036_/X _81676_/Q sky130_fd_sc_hd__dfxtp_4
X_69398_ _87520_/Q _69261_/X _69396_/X _69397_/X _69398_/X sky130_fd_sc_hd__a211o_4
X_86203_ _86203_/CLK _86203_/D _86203_/Q sky130_fd_sc_hd__dfxtp_4
X_59151_ _59148_/Y _59150_/Y _58939_/X _59151_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_9_242_0_CLK clkbuf_9_243_0_CLK/A clkbuf_9_242_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_83415_ _83415_/CLK _83415_/D _83415_/Q sky130_fd_sc_hd__dfxtp_4
X_80627_ _84776_/Q _84168_/Q _80627_/Y sky130_fd_sc_hd__nand2_4
X_56363_ _56360_/A _56363_/B _55722_/B _56363_/Y sky130_fd_sc_hd__nand3_4
X_68349_ _69178_/A _69906_/A sky130_fd_sc_hd__buf_2
X_87183_ _87183_/CLK _44200_/Y _43983_/A sky130_fd_sc_hd__dfxtp_4
X_53575_ _53565_/A _57609_/B _53575_/Y sky130_fd_sc_hd__nand2_4
X_84395_ _84396_/CLK _62627_/Y _84395_/Q sky130_fd_sc_hd__dfxtp_4
X_50787_ _50718_/A _50787_/X sky130_fd_sc_hd__buf_2
X_58102_ _58085_/X _85381_/Q _58101_/X _58102_/Y sky130_fd_sc_hd__o21ai_4
X_55314_ _55323_/A _85135_/Q _55314_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_136_0_CLK clkbuf_9_68_0_CLK/X _81296_/CLK sky130_fd_sc_hd__clkbuf_1
X_86134_ _85527_/CLK _86134_/D _86134_/Q sky130_fd_sc_hd__dfxtp_4
X_40540_ _82307_/Q _40467_/B _40540_/X sky130_fd_sc_hd__or2_4
X_52526_ _52518_/A _52526_/B _52526_/Y sky130_fd_sc_hd__nand2_4
X_59082_ _58934_/X _85658_/Q _59081_/X _59082_/X sky130_fd_sc_hd__o21a_4
X_71360_ _71344_/X _83526_/Q _71359_/X _71360_/X sky130_fd_sc_hd__a21o_4
X_83346_ _82251_/CLK _83346_/D _83346_/Q sky130_fd_sc_hd__dfxtp_4
X_56294_ _56284_/X _56016_/X _56293_/Y _56294_/Y sky130_fd_sc_hd__o21ai_4
X_80558_ _84771_/Q _84163_/Q _80560_/A sky130_fd_sc_hd__xor2_4
Xclkbuf_10_766_0_CLK clkbuf_9_383_0_CLK/X _87782_/CLK sky130_fd_sc_hd__clkbuf_1
X_58033_ _57966_/X _85707_/Q _58020_/X _58033_/X sky130_fd_sc_hd__o21a_4
X_70311_ _70247_/X _70328_/B sky130_fd_sc_hd__buf_2
X_55245_ _55245_/A _55276_/A sky130_fd_sc_hd__buf_2
X_86065_ _85748_/CLK _51151_/Y _86065_/Q sky130_fd_sc_hd__dfxtp_4
X_52457_ _85818_/Q _52438_/X _52456_/Y _52457_/Y sky130_fd_sc_hd__o21ai_4
X_40471_ _40947_/A _40471_/X sky130_fd_sc_hd__buf_2
X_71291_ _71287_/Y _71291_/Y sky130_fd_sc_hd__inv_2
X_83277_ _83278_/CLK _83277_/D _72165_/A sky130_fd_sc_hd__dfxtp_4
X_80489_ _80489_/A _80489_/B _80489_/X sky130_fd_sc_hd__or2_4
Xclkbuf_9_257_0_CLK clkbuf_8_128_0_CLK/X clkbuf_9_257_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_42210_ _42162_/A _42210_/X sky130_fd_sc_hd__buf_2
X_73030_ _44127_/X _73030_/X sky130_fd_sc_hd__buf_2
X_85016_ _85049_/CLK _85016_/D _85016_/Q sky130_fd_sc_hd__dfxtp_4
X_51408_ _51403_/X _52936_/B _51408_/Y sky130_fd_sc_hd__nand2_4
X_70242_ _70238_/X _74804_/B _70241_/X _83825_/D sky130_fd_sc_hd__a21o_4
X_82228_ _82515_/CLK _82260_/Q _82228_/Q sky130_fd_sc_hd__dfxtp_4
X_43190_ _43190_/A _43190_/Y sky130_fd_sc_hd__inv_2
X_55176_ _85132_/Q _55176_/Y sky130_fd_sc_hd__inv_2
X_52388_ _65247_/B _52372_/X _52387_/Y _52388_/Y sky130_fd_sc_hd__o21ai_4
X_42141_ _42077_/A _42141_/X sky130_fd_sc_hd__buf_2
X_54127_ _53418_/X _54127_/X sky130_fd_sc_hd__buf_2
X_51339_ _51793_/A _51339_/X sky130_fd_sc_hd__buf_2
X_70173_ _70232_/A _70183_/B sky130_fd_sc_hd__buf_2
X_82159_ _84197_/CLK _84151_/Q _82159_/Q sky130_fd_sc_hd__dfxtp_4
X_59984_ _59976_/A _62576_/C sky130_fd_sc_hd__buf_2
X_58935_ _58934_/X _85924_/Q _58793_/X _58935_/X sky130_fd_sc_hd__o21a_4
X_54058_ _54020_/A _54058_/B _54058_/Y sky130_fd_sc_hd__nand2_4
X_42072_ _51719_/A _42072_/X sky130_fd_sc_hd__buf_2
X_74981_ _74987_/B _74987_/C _74981_/Y sky130_fd_sc_hd__nand2_4
X_86967_ _86934_/CLK _86967_/D _86967_/Q sky130_fd_sc_hd__dfxtp_4
X_45900_ _42447_/C _45893_/B _45893_/C _45900_/Y sky130_fd_sc_hd__nor3_4
X_41023_ _41022_/Y _88292_/D sky130_fd_sc_hd__inv_2
X_53009_ _53006_/Y _53001_/X _53008_/X _53009_/Y sky130_fd_sc_hd__a21oi_4
X_76720_ _76708_/A _76707_/X _76720_/X sky130_fd_sc_hd__or2_4
X_85918_ _86558_/CLK _85918_/D _73636_/B sky130_fd_sc_hd__dfxtp_4
X_73932_ _73930_/X _84978_/Q _45885_/X _73931_/X _73932_/X sky130_fd_sc_hd__a211o_4
X_46880_ _46860_/X _51037_/B _46880_/Y sky130_fd_sc_hd__nand2_4
X_58866_ _58941_/A _86378_/Q _58866_/Y sky130_fd_sc_hd__nor2_4
X_86898_ _86887_/CLK _45112_/Y _64364_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_704_0_CLK clkbuf_9_352_0_CLK/X _86784_/CLK sky130_fd_sc_hd__clkbuf_1
X_45831_ _82981_/Q _45832_/A sky130_fd_sc_hd__inv_2
X_57817_ _57813_/Y _57816_/Y _57718_/X _57817_/X sky130_fd_sc_hd__a21o_4
X_76651_ _76650_/Y _81682_/Q _76651_/Y sky130_fd_sc_hd__nand2_4
X_73863_ _73863_/A _73863_/B _73864_/B sky130_fd_sc_hd__nand2_4
X_85849_ _85558_/CLK _85849_/D _64826_/B sky130_fd_sc_hd__dfxtp_4
X_58797_ _58714_/X _85775_/Q _58716_/X _58797_/X sky130_fd_sc_hd__o21a_4
X_75602_ _75601_/Y _75588_/Y _75595_/A _75602_/Y sky130_fd_sc_hd__o21ai_4
X_48550_ _48550_/A _48550_/Y sky130_fd_sc_hd__inv_2
X_72814_ _72814_/A _73306_/A sky130_fd_sc_hd__buf_2
X_79370_ _58738_/Y _66435_/Y _79369_/Y _79374_/A sky130_fd_sc_hd__o21a_4
X_45762_ _45759_/X _45761_/Y _45714_/X _45762_/Y sky130_fd_sc_hd__a21oi_4
X_57748_ _46224_/X _85406_/Q _57747_/X _57748_/Y sky130_fd_sc_hd__o21ai_4
X_76582_ _76614_/A _76614_/C _76583_/A sky130_fd_sc_hd__and2_4
X_42974_ _42970_/X _42971_/X _40440_/X _66861_/B _42954_/X _42975_/A
+ sky130_fd_sc_hd__o32ai_4
X_73794_ _70106_/Y _73697_/X _73793_/X _73794_/Y sky130_fd_sc_hd__o21ai_4
X_47501_ _47501_/A _47502_/A sky130_fd_sc_hd__inv_2
X_78321_ _78312_/A _82658_/D _78321_/Y sky130_fd_sc_hd__nand2_4
X_44713_ _41936_/A _44713_/X sky130_fd_sc_hd__buf_2
X_75533_ _75530_/Y _75533_/B _75531_/Y _75533_/Y sky130_fd_sc_hd__nand3_4
X_87519_ _87273_/CLK _43249_/X _87519_/Q sky130_fd_sc_hd__dfxtp_4
X_41925_ _41925_/A _88103_/D sky130_fd_sc_hd__inv_2
X_48481_ _73073_/A _48482_/B sky130_fd_sc_hd__buf_2
X_72745_ _72745_/A _73351_/A sky130_fd_sc_hd__buf_2
X_45693_ _85038_/Q _45675_/X _45692_/X _45693_/Y sky130_fd_sc_hd__o21ai_4
X_57679_ _84955_/Q _57680_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_719_0_CLK clkbuf_9_359_0_CLK/X _87757_/CLK sky130_fd_sc_hd__clkbuf_1
X_47432_ _47431_/Y _53046_/B sky130_fd_sc_hd__buf_2
X_59418_ _84738_/Q _59419_/A sky130_fd_sc_hd__inv_2
X_78252_ _78252_/A _78241_/X _78252_/C _78252_/X sky130_fd_sc_hd__and3_4
X_44644_ _44644_/A _44644_/Y sky130_fd_sc_hd__inv_2
X_75464_ _75462_/X _75507_/A _75506_/C sky130_fd_sc_hd__and2_4
X_41856_ _41856_/A _88119_/D sky130_fd_sc_hd__inv_2
X_60690_ _60686_/X _60689_/Y _60690_/X sky130_fd_sc_hd__and2_4
X_72676_ _83194_/Q _72672_/X _72675_/Y _72676_/X sky130_fd_sc_hd__a21bo_4
X_77203_ _77188_/X _77203_/B _77205_/A sky130_fd_sc_hd__or2_4
X_74415_ _83071_/Q _74412_/X _74414_/Y _74415_/Y sky130_fd_sc_hd__o21ai_4
X_40807_ _40806_/X _40793_/X _88331_/Q _40794_/X _40807_/X sky130_fd_sc_hd__a2bb2o_4
X_47363_ _47363_/A _47414_/A sky130_fd_sc_hd__buf_2
X_71627_ _71625_/Y _83433_/Q _71626_/Y _71627_/X sky130_fd_sc_hd__a21o_4
X_59349_ _59311_/X _85733_/Q _59334_/X _59349_/X sky130_fd_sc_hd__o21a_4
X_78183_ _78183_/A _82489_/Q _78191_/B sky130_fd_sc_hd__or2_4
X_44575_ _44565_/X _44567_/X _40885_/X _87049_/Q _44568_/X _44575_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75395_ _75394_/Y _75396_/C sky130_fd_sc_hd__inv_2
X_41787_ _41753_/X _41754_/X _41786_/X _88149_/Q _41736_/X _41788_/A
+ sky130_fd_sc_hd__o32ai_4
X_49102_ _52370_/A _49113_/B _49091_/C _49102_/X sky130_fd_sc_hd__and3_4
X_46314_ _46313_/Y _51261_/B sky130_fd_sc_hd__buf_2
X_77134_ _77134_/A _82293_/D _77141_/C sky130_fd_sc_hd__nand2_4
X_43526_ _40387_/X _43513_/X _87376_/Q _43514_/X _43526_/X sky130_fd_sc_hd__a2bb2o_4
X_62360_ _59896_/X _62420_/B sky130_fd_sc_hd__buf_2
X_74346_ _83090_/Q _74340_/X _74345_/Y _83090_/D sky130_fd_sc_hd__a21bo_4
X_40738_ _40731_/X _82854_/Q _40737_/X _40739_/A sky130_fd_sc_hd__o21ai_4
X_47294_ _47294_/A _52967_/D sky130_fd_sc_hd__buf_2
X_71558_ _71164_/B _71558_/X sky130_fd_sc_hd__buf_2
X_49033_ _49027_/Y _48985_/X _49032_/X _86451_/D sky130_fd_sc_hd__a21oi_4
X_61311_ _72529_/C _72506_/C sky130_fd_sc_hd__buf_2
X_46245_ _44803_/A _46241_/X _46244_/Y _46245_/X sky130_fd_sc_hd__o21a_4
X_70509_ _70511_/A _70940_/B _70508_/X _70509_/Y sky130_fd_sc_hd__nand3_4
XPHY_570 sky130_fd_sc_hd__decap_3
X_77065_ _77065_/A _77065_/B _77065_/X sky130_fd_sc_hd__xor2_4
X_43457_ _43449_/X _43452_/X _41621_/X _87413_/Q _43456_/X _43458_/A
+ sky130_fd_sc_hd__o32ai_4
X_74277_ _72730_/X _84962_/Q _74021_/X _74276_/X _74278_/B sky130_fd_sc_hd__a211o_4
X_62291_ _62572_/A _62634_/A sky130_fd_sc_hd__buf_2
XPHY_581 sky130_fd_sc_hd__decap_3
X_40669_ _40669_/A _88357_/D sky130_fd_sc_hd__inv_2
X_71489_ _71488_/X _71422_/C _70483_/B _71489_/X sky130_fd_sc_hd__and3_4
XPHY_592 sky130_fd_sc_hd__decap_3
X_76016_ _81519_/Q _81743_/D _81768_/D sky130_fd_sc_hd__xor2_4
X_64030_ _62005_/A _64046_/B _64046_/C _64016_/D _64030_/Y sky130_fd_sc_hd__nand4_4
X_42408_ _42401_/X _42397_/X _40452_/X _87877_/Q _42398_/X _42408_/Y
+ sky130_fd_sc_hd__o32ai_4
X_61242_ _75902_/A _60979_/X _61163_/Y _61241_/X _61242_/Y sky130_fd_sc_hd__a2bb2oi_4
X_73228_ _73228_/A _73228_/B _73228_/Y sky130_fd_sc_hd__nor2_4
X_46176_ _46174_/X _46175_/Y _46158_/B _86767_/D sky130_fd_sc_hd__o21ai_4
X_43388_ _43397_/A _43388_/X sky130_fd_sc_hd__buf_2
X_45127_ _45350_/A _45127_/X sky130_fd_sc_hd__buf_2
X_42339_ _42330_/X _42319_/X _41688_/X _87913_/Q _42320_/X _42340_/A
+ sky130_fd_sc_hd__o32ai_4
X_61173_ _61173_/A _61173_/Y sky130_fd_sc_hd__inv_2
X_73159_ _72870_/X _86194_/Q _72905_/X _73158_/X _73159_/X sky130_fd_sc_hd__a211o_4
X_60124_ _59852_/A _60214_/B sky130_fd_sc_hd__buf_2
X_49935_ _49854_/A _49955_/A sky130_fd_sc_hd__buf_2
X_45058_ _56219_/C _44998_/X _45057_/X _45058_/Y sky130_fd_sc_hd__o21ai_4
X_65981_ _65980_/X _73689_/B _65981_/X sky130_fd_sc_hd__and2_4
X_77967_ _77960_/Y _77967_/B _77967_/C _77967_/Y sky130_fd_sc_hd__nand3_4
X_44009_ _57686_/A _44247_/A sky130_fd_sc_hd__buf_2
X_67720_ _87395_/Q _67717_/X _67718_/X _67719_/X _67720_/X sky130_fd_sc_hd__a211o_4
X_79706_ _79692_/Y _79689_/Y _79706_/X sky130_fd_sc_hd__and2_4
X_64932_ _64858_/X _85557_/Q _64859_/X _64931_/X _64932_/X sky130_fd_sc_hd__a211o_4
X_60055_ _60055_/A _60056_/A sky130_fd_sc_hd__buf_2
X_76918_ _76918_/A _76918_/B _76931_/B sky130_fd_sc_hd__xor2_4
X_49866_ _49851_/A _49884_/B _49862_/C _53078_/D _49866_/X sky130_fd_sc_hd__and4_4
X_77898_ _82164_/Q _82036_/D _82132_/D sky130_fd_sc_hd__xor2_4
X_48817_ _86477_/Q _48809_/X _48816_/Y _48817_/Y sky130_fd_sc_hd__o21ai_4
X_67651_ _68402_/A _67651_/X sky130_fd_sc_hd__buf_2
X_79637_ _60346_/C _79637_/B _79646_/B sky130_fd_sc_hd__xor2_4
X_64863_ _44170_/A _64991_/A sky130_fd_sc_hd__buf_2
X_76849_ _76849_/A _76854_/A sky130_fd_sc_hd__inv_2
X_49797_ _49792_/Y _49787_/X _49796_/X _86322_/D sky130_fd_sc_hd__a21oi_4
X_66602_ _66602_/A _66602_/B _66602_/X sky130_fd_sc_hd__and2_4
X_63814_ _61376_/X _63781_/B _63814_/C _63761_/X _63814_/Y sky130_fd_sc_hd__nand4_4
X_48748_ _52135_/A _48766_/B _48761_/C _48748_/X sky130_fd_sc_hd__and3_4
X_67582_ _67582_/A _87209_/Q _67582_/X sky130_fd_sc_hd__and2_4
X_79568_ _79567_/Y _79568_/B _79569_/B sky130_fd_sc_hd__nand2_4
X_64794_ _64769_/A _64794_/B _64794_/X sky130_fd_sc_hd__and2_4
X_69321_ _69223_/A _69322_/A sky130_fd_sc_hd__buf_2
X_66533_ _66565_/A _66534_/A sky130_fd_sc_hd__buf_2
X_78519_ _78519_/A _78519_/B _82768_/D sky130_fd_sc_hd__xor2_4
X_63745_ _63701_/A _63701_/B _63745_/C _63745_/Y sky130_fd_sc_hd__nor3_4
X_48679_ _48623_/A _48894_/C sky130_fd_sc_hd__buf_2
X_60957_ _63781_/C _60957_/B _60957_/Y sky130_fd_sc_hd__nor2_4
X_79499_ _84815_/Q _84135_/Q _79499_/Y sky130_fd_sc_hd__nand2_4
X_50710_ _50695_/A _50710_/B _50710_/Y sky130_fd_sc_hd__nand2_4
X_81530_ _82053_/CLK _81542_/Q _81530_/Q sky130_fd_sc_hd__dfxtp_4
X_69252_ _69247_/X _69250_/X _69251_/X _69255_/A sky130_fd_sc_hd__a21o_4
X_66464_ _66433_/A _66419_/X _84118_/Q _66464_/X sky130_fd_sc_hd__and3_4
X_51690_ _51687_/Y _51667_/X _51689_/X _85964_/D sky130_fd_sc_hd__a21oi_4
X_63676_ _61649_/B _63609_/X _63674_/X _63675_/X _63676_/X sky130_fd_sc_hd__a211o_4
X_60888_ _60863_/X _60888_/Y sky130_fd_sc_hd__inv_2
X_68203_ _82053_/D _68200_/X _68202_/X _68203_/X sky130_fd_sc_hd__a21bo_4
Xclkbuf_10_1023_0_CLK clkbuf_9_511_0_CLK/X _86500_/CLK sky130_fd_sc_hd__clkbuf_1
X_65415_ _65412_/X _65414_/X _65287_/X _65415_/X sky130_fd_sc_hd__a21o_4
X_50641_ _50637_/Y _50619_/X _50640_/Y _50641_/Y sky130_fd_sc_hd__a21boi_4
X_62627_ _62625_/Y _62593_/X _62626_/Y _62627_/Y sky130_fd_sc_hd__a21oi_4
X_81461_ _81461_/CLK _76826_/B _81461_/Q sky130_fd_sc_hd__dfxtp_4
X_69183_ _69183_/A _69183_/X sky130_fd_sc_hd__buf_2
X_66395_ _66389_/A _66389_/B _66395_/C _66395_/Y sky130_fd_sc_hd__nor3_4
X_83200_ _83843_/CLK _83200_/D _70198_/C sky130_fd_sc_hd__dfxtp_4
X_80412_ _84757_/Q _80419_/B _80412_/X sky130_fd_sc_hd__xor2_4
X_68134_ _66844_/X _66846_/X _68133_/X _68134_/Y sky130_fd_sc_hd__a21oi_4
X_53360_ _53353_/A _53360_/B _53360_/Y sky130_fd_sc_hd__nand2_4
X_65346_ _65198_/X _65333_/Y _65345_/Y _65346_/Y sky130_fd_sc_hd__o21ai_4
X_84180_ _84194_/CLK _84180_/D _84180_/Q sky130_fd_sc_hd__dfxtp_4
X_50572_ _50572_/A _50580_/A sky130_fd_sc_hd__buf_2
X_62558_ _62557_/Y _59945_/Y _84785_/Q _59931_/A _62558_/X sky130_fd_sc_hd__a2bb2o_4
X_81392_ _81473_/CLK _83928_/Q _76929_/B sky130_fd_sc_hd__dfxtp_4
X_52311_ _52308_/Y _52289_/X _52310_/X _85848_/D sky130_fd_sc_hd__a21oi_4
X_83131_ _83561_/CLK _73915_/Y _70113_/A sky130_fd_sc_hd__dfxtp_4
X_61509_ _61499_/A _61509_/B _61459_/X _61509_/Y sky130_fd_sc_hd__nand3_4
X_80343_ _80347_/A _80347_/B _80343_/X sky130_fd_sc_hd__xor2_4
X_68065_ _81475_/D _68040_/X _68064_/X _68065_/X sky130_fd_sc_hd__a21bo_4
X_53291_ _85660_/Q _53268_/X _53290_/Y _53291_/Y sky130_fd_sc_hd__o21ai_4
X_65277_ _64851_/A _65277_/X sky130_fd_sc_hd__buf_2
X_62489_ _62236_/A _62566_/B sky130_fd_sc_hd__buf_2
X_55030_ _54927_/A _55030_/X sky130_fd_sc_hd__buf_2
X_67016_ _67010_/X _67012_/X _67015_/X _67016_/Y sky130_fd_sc_hd__a21oi_4
X_52242_ _85861_/Q _52239_/X _52241_/Y _52242_/Y sky130_fd_sc_hd__o21ai_4
X_64228_ _59454_/A _64226_/X _64227_/Y _64228_/Y sky130_fd_sc_hd__o21ai_4
X_83062_ _85571_/CLK _74460_/Y _83062_/Q sky130_fd_sc_hd__dfxtp_4
X_80274_ _84747_/Q _84139_/Q _80274_/Y sky130_fd_sc_hd__nand2_4
X_82013_ _82009_/CLK _82013_/D _77194_/A sky130_fd_sc_hd__dfxtp_4
X_52173_ _52168_/A _48788_/B _52173_/Y sky130_fd_sc_hd__nand2_4
X_64159_ _64155_/Y _64159_/B _64157_/Y _64159_/D _64159_/X sky130_fd_sc_hd__and4_4
X_87870_ _88128_/CLK _87870_/D _87870_/Q sky130_fd_sc_hd__dfxtp_4
X_51124_ _86069_/Q _51101_/X _51123_/Y _51124_/Y sky130_fd_sc_hd__o21ai_4
X_86821_ _88245_/CLK _86821_/D _66975_/B sky130_fd_sc_hd__dfxtp_4
X_56981_ _56696_/A _44220_/B _56980_/Y _85105_/D sky130_fd_sc_hd__a21oi_4
X_68967_ _69011_/A _87227_/Q _68967_/X sky130_fd_sc_hd__and2_4
X_58720_ _58659_/A _58720_/B _58720_/Y sky130_fd_sc_hd__nor2_4
X_51055_ _50973_/A _51056_/A sky130_fd_sc_hd__buf_2
X_55932_ _56392_/C _55641_/A _55610_/X _55931_/X _55932_/X sky130_fd_sc_hd__a211o_4
X_67918_ _67913_/X _67916_/X _67917_/X _67918_/X sky130_fd_sc_hd__a21o_4
X_86752_ _85535_/CLK _86752_/D _86752_/Q sky130_fd_sc_hd__dfxtp_4
X_83964_ _81994_/CLK _68712_/X _83964_/Q sky130_fd_sc_hd__dfxtp_4
X_68898_ _68759_/A _68898_/B _68898_/X sky130_fd_sc_hd__and2_4
X_50006_ _50002_/Y _50003_/X _50005_/X _86283_/D sky130_fd_sc_hd__a21oi_4
X_85703_ _85700_/CLK _85703_/D _85703_/Q sky130_fd_sc_hd__dfxtp_4
X_58651_ _58631_/X _58648_/Y _58649_/Y _58650_/X _58636_/X _58651_/X
+ sky130_fd_sc_hd__o32a_4
X_82915_ _86582_/CLK _78139_/X _82915_/Q sky130_fd_sc_hd__dfxtp_4
X_55863_ _55862_/X _55863_/X sky130_fd_sc_hd__buf_2
X_67849_ _86954_/Q _67825_/X _67755_/X _67848_/X _67849_/X sky130_fd_sc_hd__a211o_4
X_86683_ _86361_/CLK _46982_/Y _59068_/A sky130_fd_sc_hd__dfxtp_4
X_83895_ _82299_/CLK _83895_/D _81967_/D sky130_fd_sc_hd__dfxtp_4
X_57602_ _57600_/Y _57592_/X _57601_/X _84971_/D sky130_fd_sc_hd__a21oi_4
X_54814_ _54823_/A _47561_/Y _54814_/Y sky130_fd_sc_hd__nand2_4
X_85634_ _86655_/CLK _53440_/Y _85634_/Q sky130_fd_sc_hd__dfxtp_4
X_70860_ _70860_/A _71088_/C _70863_/C _70860_/D _70860_/Y sky130_fd_sc_hd__nand4_4
X_58582_ _58140_/X _86112_/Q _58581_/X _58582_/Y sky130_fd_sc_hd__o21ai_4
X_82846_ _81019_/CLK _82846_/D _82814_/D sky130_fd_sc_hd__dfxtp_4
X_55794_ _55794_/A _85164_/Q _55794_/X sky130_fd_sc_hd__and2_4
X_57533_ _57528_/X _53501_/B _57533_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_690_0_CLK clkbuf_9_345_0_CLK/X _86914_/CLK sky130_fd_sc_hd__clkbuf_1
X_69519_ _81382_/D _69504_/X _69518_/X _83918_/D sky130_fd_sc_hd__a21bo_4
X_88353_ _87859_/CLK _88353_/D _88353_/Q sky130_fd_sc_hd__dfxtp_4
X_54745_ _54731_/X _47451_/A _54745_/Y sky130_fd_sc_hd__nand2_4
X_85565_ _85561_/CLK _85565_/D _85565_/Q sky130_fd_sc_hd__dfxtp_4
X_51957_ _51956_/X _51958_/C sky130_fd_sc_hd__buf_2
X_70791_ _70903_/A _70791_/B _70791_/C _70791_/D _70791_/Y sky130_fd_sc_hd__nand4_4
X_82777_ _82206_/CLK _82777_/D _82777_/Q sky130_fd_sc_hd__dfxtp_4
X_87304_ _87820_/CLK _43697_/X _73056_/A sky130_fd_sc_hd__dfxtp_4
X_41710_ _41709_/X _41710_/X sky130_fd_sc_hd__buf_2
X_72530_ _72530_/A _72569_/A sky130_fd_sc_hd__buf_2
X_84516_ _84498_/CLK _84516_/D _61165_/C sky130_fd_sc_hd__dfxtp_4
X_50908_ _50908_/A _50919_/B _50897_/X _51772_/D _50908_/X sky130_fd_sc_hd__and4_4
Xclkbuf_9_181_0_CLK clkbuf_8_90_0_CLK/X clkbuf_9_181_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_81728_ _84079_/CLK _81728_/D _41119_/A sky130_fd_sc_hd__dfxtp_4
X_57464_ _57441_/X _83335_/Q _57463_/X _57464_/X sky130_fd_sc_hd__o21a_4
X_88284_ _87011_/CLK _88284_/D _88284_/Q sky130_fd_sc_hd__dfxtp_4
X_42690_ _42689_/Y _87769_/D sky130_fd_sc_hd__inv_2
X_54676_ _54729_/A _54676_/X sky130_fd_sc_hd__buf_2
X_85496_ _83745_/CLK _85496_/D _85496_/Q sky130_fd_sc_hd__dfxtp_4
X_51888_ _51885_/Y _51877_/X _51887_/X _51888_/Y sky130_fd_sc_hd__a21oi_4
X_59203_ _84761_/Q _59129_/X _59195_/X _59202_/X _84761_/D sky130_fd_sc_hd__a2bb2oi_4
X_56415_ _56079_/X _56409_/X _56414_/Y _85203_/D sky130_fd_sc_hd__o21ai_4
X_87235_ _87235_/CLK _43850_/X _87235_/Q sky130_fd_sc_hd__dfxtp_4
X_41641_ _82911_/Q _41624_/B _41641_/X sky130_fd_sc_hd__or2_4
X_53627_ _54067_/A _53656_/A sky130_fd_sc_hd__buf_2
X_72461_ _72461_/A _72461_/B _72461_/Y sky130_fd_sc_hd__nor2_4
X_84447_ _84452_/CLK _61900_/Y _78070_/B sky130_fd_sc_hd__dfxtp_4
X_50839_ _50957_/A _50839_/X sky130_fd_sc_hd__buf_2
X_57395_ _57380_/X _57395_/X sky130_fd_sc_hd__buf_2
X_81659_ _81279_/CLK _76728_/A _81659_/Q sky130_fd_sc_hd__dfxtp_4
X_74200_ _53593_/B _74200_/B _74201_/B sky130_fd_sc_hd__xor2_4
X_59134_ _59115_/X _59130_/Y _59131_/Y _59133_/X _59119_/X _59134_/X
+ sky130_fd_sc_hd__o32a_4
X_71412_ _71396_/Y _83508_/Q _71411_/Y _71412_/X sky130_fd_sc_hd__a21o_4
X_44360_ _44350_/X _44351_/X _41735_/X _87147_/Q _44353_/X _44361_/A
+ sky130_fd_sc_hd__o32ai_4
X_56346_ _56130_/X _56337_/X _56345_/Y _85227_/D sky130_fd_sc_hd__o21ai_4
X_75180_ _75180_/A _75179_/Y _75182_/A sky130_fd_sc_hd__nor2_4
X_87166_ _81746_/CLK _87166_/D _87166_/Q sky130_fd_sc_hd__dfxtp_4
X_53558_ _53622_/A _57590_/B _53558_/Y sky130_fd_sc_hd__nand2_4
X_41572_ _41572_/A _41563_/B _41572_/X sky130_fd_sc_hd__or2_4
X_72392_ _72388_/Y _72391_/Y _72344_/X _72392_/X sky130_fd_sc_hd__a21o_4
X_84378_ _84507_/CLK _84378_/D _84378_/Q sky130_fd_sc_hd__dfxtp_4
X_43311_ _43296_/X _43305_/X _41220_/X _87487_/Q _43308_/X _43312_/A
+ sky130_fd_sc_hd__o32ai_4
X_74131_ _74128_/X _74130_/X _74085_/X _74134_/A sky130_fd_sc_hd__a21o_4
X_86117_ _86121_/CLK _50869_/Y _86117_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_196_0_CLK clkbuf_8_98_0_CLK/X clkbuf_9_196_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_40523_ _40463_/X _81159_/Q _40522_/X _40523_/Y sky130_fd_sc_hd__o21ai_4
X_52509_ _50812_/A _52509_/B _52498_/C _52509_/X sky130_fd_sc_hd__and3_4
X_71343_ _71343_/A _71344_/A sky130_fd_sc_hd__inv_2
X_59065_ _84772_/Q _59043_/X _59058_/X _59064_/X _84772_/D sky130_fd_sc_hd__a2bb2oi_4
X_83329_ _83337_/CLK _83329_/D _83329_/Q sky130_fd_sc_hd__dfxtp_4
X_44291_ _44290_/X _44292_/A sky130_fd_sc_hd__buf_2
X_56277_ _56277_/A _56279_/A sky130_fd_sc_hd__inv_2
X_87097_ _88272_/CLK _44462_/X _87097_/Q sky130_fd_sc_hd__dfxtp_4
X_53489_ _53487_/Y _53455_/X _53488_/Y _85627_/D sky130_fd_sc_hd__a21boi_4
X_46030_ _45975_/X _46030_/X sky130_fd_sc_hd__buf_2
X_58016_ _58010_/X _58012_/Y _58013_/Y _57899_/X _58015_/X _58016_/X
+ sky130_fd_sc_hd__o32a_4
X_43242_ _43241_/X _43229_/X _41036_/X _87521_/Q _43232_/X _43243_/A
+ sky130_fd_sc_hd__o32ai_4
X_55228_ _55218_/Y _55226_/Y _55227_/Y _55228_/Y sky130_fd_sc_hd__o21ai_4
X_74062_ _74059_/X _74061_/X _74019_/X _74065_/A sky130_fd_sc_hd__a21o_4
X_86048_ _85536_/CLK _51243_/Y _64617_/B sky130_fd_sc_hd__dfxtp_4
X_40454_ _40454_/A _40454_/Y sky130_fd_sc_hd__inv_2
X_71274_ _71173_/A _71276_/B _71276_/C _71276_/D _71274_/Y sky130_fd_sc_hd__nand4_4
X_73013_ _72959_/X _85592_/Q _72839_/X _73012_/X _73013_/X sky130_fd_sc_hd__a211o_4
X_70225_ _70229_/A _70229_/B _70225_/C _70229_/D _70225_/X sky130_fd_sc_hd__and4_4
X_55159_ _55159_/A _85130_/Q _55159_/X sky130_fd_sc_hd__and2_4
X_43173_ _43162_/X _43167_/X _40885_/X _73323_/A _43172_/X _43174_/A
+ sky130_fd_sc_hd__o32ai_4
X_78870_ _78870_/A _78886_/A sky130_fd_sc_hd__inv_2
X_40385_ _82334_/Q _40385_/B _40385_/X sky130_fd_sc_hd__or2_4
X_42124_ _42124_/A _88024_/D sky130_fd_sc_hd__inv_2
X_77821_ _82059_/Q _77818_/Y _77820_/X _77822_/B sky130_fd_sc_hd__o21ai_4
X_70156_ _70155_/X _70157_/A sky130_fd_sc_hd__buf_2
X_47981_ _47857_/X _47981_/X sky130_fd_sc_hd__buf_2
X_59967_ _59966_/Y _59935_/A _59985_/A _59968_/B sky130_fd_sc_hd__a21o_4
X_87999_ _88001_/CLK _42172_/Y _87999_/Q sky130_fd_sc_hd__dfxtp_4
X_49720_ _49718_/Y _49706_/X _49719_/X _86336_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_643_0_CLK clkbuf_9_321_0_CLK/X _87653_/CLK sky130_fd_sc_hd__clkbuf_1
X_46932_ _82400_/Q _54449_/D sky130_fd_sc_hd__inv_2
X_42055_ _42052_/X _42043_/X _40914_/X _73462_/A _42044_/X _42056_/A
+ sky130_fd_sc_hd__o32ai_4
X_58918_ _58918_/A _58918_/X sky130_fd_sc_hd__buf_2
X_77752_ _77752_/A _77758_/A _77753_/B sky130_fd_sc_hd__nand2_4
X_74964_ _80946_/Q _74964_/B _74964_/X sky130_fd_sc_hd__xor2_4
X_70087_ _69603_/X _69937_/Y _70081_/X _70086_/Y _70087_/X sky130_fd_sc_hd__a211o_4
X_59898_ _59898_/A _60058_/B sky130_fd_sc_hd__buf_2
X_41006_ _41005_/Y _41006_/Y sky130_fd_sc_hd__inv_2
X_76703_ _76703_/A _76703_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_9_134_0_CLK clkbuf_8_67_0_CLK/X clkbuf_9_134_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_49651_ _49571_/A _49651_/X sky130_fd_sc_hd__buf_2
X_73915_ _70117_/A _73818_/X _73914_/X _73915_/Y sky130_fd_sc_hd__o21ai_4
X_46863_ _46860_/X _51026_/B _46863_/Y sky130_fd_sc_hd__nand2_4
X_58849_ _58796_/X _86091_/Q _58848_/X _58849_/Y sky130_fd_sc_hd__o21ai_4
X_77683_ _77687_/B _77688_/B sky130_fd_sc_hd__inv_2
Xclkbuf_9_61_0_CLK clkbuf_9_61_0_CLK/A clkbuf_9_61_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_74895_ _80937_/Q _74895_/B _81186_/D sky130_fd_sc_hd__xor2_4
X_48602_ _48602_/A _48602_/Y sky130_fd_sc_hd__inv_2
X_79422_ _79401_/B _79418_/X _79421_/Y _79422_/Y sky130_fd_sc_hd__a21oi_4
X_45814_ _45810_/X _45813_/X _45757_/X _45814_/X sky130_fd_sc_hd__a21o_4
X_76634_ _76620_/X _81664_/Q _76633_/Y _76634_/Y sky130_fd_sc_hd__a21oi_4
X_49582_ _86361_/Q _49579_/X _49581_/Y _49582_/Y sky130_fd_sc_hd__o21ai_4
X_61860_ _61427_/B _61843_/B _61860_/C _61860_/D _61860_/Y sky130_fd_sc_hd__nand4_4
X_73846_ _68672_/B _73597_/X _73772_/X _73845_/Y _73846_/X sky130_fd_sc_hd__a211o_4
X_46794_ _46794_/A _52677_/B sky130_fd_sc_hd__inv_2
Xclkbuf_10_658_0_CLK clkbuf_9_329_0_CLK/X _87671_/CLK sky130_fd_sc_hd__clkbuf_1
X_48533_ _48533_/A _48500_/X _48533_/C _48533_/X sky130_fd_sc_hd__and3_4
X_60811_ _60684_/X _60692_/X _60737_/Y _60809_/Y _60810_/Y _84561_/D
+ sky130_fd_sc_hd__a41oi_4
X_79353_ _79351_/X _79360_/B _79353_/Y sky130_fd_sc_hd__xnor2_4
X_45745_ _45745_/A _74679_/B sky130_fd_sc_hd__inv_2
X_76565_ _76563_/X _76566_/A sky130_fd_sc_hd__inv_2
X_42957_ _40387_/X _42950_/X _87632_/Q _42951_/X _42957_/X sky130_fd_sc_hd__a2bb2o_4
X_61791_ _61839_/A _61791_/B _61732_/X _63051_/B _61791_/X sky130_fd_sc_hd__and4_4
X_73777_ _72899_/A _73777_/X sky130_fd_sc_hd__buf_2
X_70989_ _70944_/A _70990_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_149_0_CLK clkbuf_8_74_0_CLK/X clkbuf_9_149_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_78304_ _78306_/C _78304_/Y sky130_fd_sc_hd__inv_2
X_63530_ _63554_/A _63554_/B _84316_/Q _63530_/Y sky130_fd_sc_hd__nor3_4
X_75516_ _80703_/Q _80959_/D _75516_/Y sky130_fd_sc_hd__nor2_4
X_41908_ _41902_/A _50256_/A sky130_fd_sc_hd__buf_2
X_48464_ _48464_/A _50443_/A sky130_fd_sc_hd__buf_2
X_72728_ _72728_/A _72769_/B _72728_/Y sky130_fd_sc_hd__nor2_4
X_60742_ _63370_/A _63648_/B sky130_fd_sc_hd__buf_2
Xclkbuf_9_76_0_CLK clkbuf_8_38_0_CLK/X clkbuf_9_76_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_79284_ _79281_/X _79283_/Y _82827_/D sky130_fd_sc_hd__xnor2_4
X_45676_ _57419_/A _45357_/X _45339_/X _45676_/X sky130_fd_sc_hd__o21a_4
X_76496_ _76491_/X _76494_/Y _76492_/Y _76513_/D sky130_fd_sc_hd__nand3_4
X_42888_ _41626_/X _42886_/X _87668_/Q _42887_/X _87668_/D sky130_fd_sc_hd__a2bb2o_4
X_47415_ _47556_/A _47415_/X sky130_fd_sc_hd__buf_2
X_78235_ _82583_/Q _82495_/Q _78235_/Y sky130_fd_sc_hd__nor2_4
X_44627_ _44627_/A _44627_/Y sky130_fd_sc_hd__inv_2
X_63461_ _63398_/A _63488_/A sky130_fd_sc_hd__buf_2
X_75447_ _75443_/Y _75445_/Y _75442_/Y _75448_/B sky130_fd_sc_hd__o21ai_4
X_41839_ _41802_/A _41839_/X sky130_fd_sc_hd__buf_2
X_48395_ _48043_/X _48914_/B _48394_/Y _74381_/A sky130_fd_sc_hd__o21ai_4
X_60673_ _72250_/A _60673_/X sky130_fd_sc_hd__buf_2
X_72659_ _72687_/A _72668_/A sky130_fd_sc_hd__buf_2
X_65200_ _64667_/A _65225_/A sky130_fd_sc_hd__buf_2
X_62412_ _62179_/X _62412_/X sky130_fd_sc_hd__buf_2
X_47346_ _57919_/A _47332_/X _47345_/Y _47346_/Y sky130_fd_sc_hd__o21ai_4
X_66180_ _66180_/A _66180_/X sky130_fd_sc_hd__buf_2
X_78166_ _78166_/A _78165_/X _78166_/Y sky130_fd_sc_hd__nand2_4
X_44558_ _44554_/X _44555_/X _40845_/A _44556_/Y _44557_/X _87056_/D
+ sky130_fd_sc_hd__o32ai_4
X_63392_ _63305_/X _63392_/B _63392_/C _63392_/Y sky130_fd_sc_hd__nor3_4
X_75378_ _75381_/B _75378_/Y sky130_fd_sc_hd__inv_2
X_65131_ _64999_/X _86157_/Q _65127_/X _65130_/X _65131_/X sky130_fd_sc_hd__a211o_4
X_77117_ _77111_/X _77126_/A _77118_/B sky130_fd_sc_hd__xor2_4
X_43509_ _41768_/X _43498_/X _87385_/Q _43499_/X _43509_/X sky130_fd_sc_hd__a2bb2o_4
X_74329_ _74342_/A _74338_/B sky130_fd_sc_hd__buf_2
X_62343_ _62339_/Y _62327_/X _62342_/Y _84417_/D sky130_fd_sc_hd__a21oi_4
X_47277_ _83387_/Q _54125_/B sky130_fd_sc_hd__inv_2
X_78097_ _82565_/Q _78103_/B _78100_/A sky130_fd_sc_hd__xnor2_4
X_44489_ _44481_/X _44482_/X _41219_/X _87083_/Q _44484_/X _44489_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49016_ _49007_/A _49015_/X _49016_/Y sky130_fd_sc_hd__nand2_4
X_46228_ _46228_/A _46090_/Y _46214_/C _46214_/D _46228_/Y sky130_fd_sc_hd__nand4_4
X_65062_ _65059_/X _85552_/Q _65060_/X _65061_/X _65062_/X sky130_fd_sc_hd__a211o_4
X_77048_ _77045_/X _77048_/B _77049_/B sky130_fd_sc_hd__xor2_4
X_62274_ _61376_/X _59898_/A _62233_/C _62597_/D _62274_/Y sky130_fd_sc_hd__nand4_4
X_64013_ _64412_/C _63934_/X _64091_/C _64027_/D _64013_/Y sky130_fd_sc_hd__nand4_4
X_61225_ _64361_/A _61128_/A _64221_/A _64419_/B sky130_fd_sc_hd__nand3_4
X_46159_ _46159_/A _46159_/X sky130_fd_sc_hd__buf_2
X_69870_ _70012_/A _69870_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_14_0_CLK clkbuf_8_7_0_CLK/X clkbuf_9_14_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_68821_ _87085_/Q _68818_/X _68819_/X _68820_/X _68821_/X sky130_fd_sc_hd__a211o_4
X_61156_ _61271_/A _61176_/B _61195_/A _61156_/X sky130_fd_sc_hd__a21o_4
X_78999_ _78993_/B _78993_/A _78998_/Y _78999_/Y sky130_fd_sc_hd__a21oi_4
X_60107_ _60125_/A _60103_/B _60107_/C _60107_/Y sky130_fd_sc_hd__nor3_4
X_49918_ _49928_/A _53131_/B _49918_/Y sky130_fd_sc_hd__nand2_4
X_68752_ _68749_/X _68751_/X _68477_/X _68752_/Y sky130_fd_sc_hd__a21oi_4
X_65964_ _66391_/A _65967_/B sky130_fd_sc_hd__buf_2
X_61087_ _61070_/X _61122_/B sky130_fd_sc_hd__buf_2
Xclkbuf_9_2_0_CLK clkbuf_9_3_0_CLK/A clkbuf_9_2_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_67703_ _67678_/X _87204_/Q _67703_/X sky130_fd_sc_hd__and2_4
X_64915_ _64561_/A _64915_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_29_0_CLK clkbuf_9_29_0_CLK/A clkbuf_9_29_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_60038_ _60027_/X _59995_/X _72584_/C _60038_/Y sky130_fd_sc_hd__o21ai_4
X_49849_ _58058_/B _49825_/X _49848_/Y _49849_/Y sky130_fd_sc_hd__o21ai_4
X_80961_ _80961_/CLK _80961_/D _75076_/B sky130_fd_sc_hd__dfxtp_4
X_68683_ _68389_/A _69035_/A sky130_fd_sc_hd__buf_2
X_65895_ _64611_/A _65896_/A sky130_fd_sc_hd__buf_2
X_82700_ _84115_/CLK _82700_/D _82700_/Q sky130_fd_sc_hd__dfxtp_4
X_67634_ _67539_/X _67634_/B _67634_/X sky130_fd_sc_hd__and2_4
X_52860_ _85741_/Q _52848_/X _52859_/Y _52860_/Y sky130_fd_sc_hd__o21ai_4
X_64846_ _64615_/A _64846_/X sky130_fd_sc_hd__buf_2
X_83680_ _83681_/CLK _70864_/Y _46700_/A sky130_fd_sc_hd__dfxtp_4
X_80892_ _80740_/CLK _80892_/D _80892_/Q sky130_fd_sc_hd__dfxtp_4
X_51811_ _51808_/Y _51793_/X _51810_/X _51811_/Y sky130_fd_sc_hd__a21oi_4
X_82631_ _88180_/CLK _83983_/Q _78857_/B sky130_fd_sc_hd__dfxtp_4
X_67565_ _67562_/X _67564_/X _67423_/X _67565_/Y sky130_fd_sc_hd__a21oi_4
X_52791_ _52788_/Y _52783_/X _52790_/X _52791_/Y sky130_fd_sc_hd__a21oi_4
X_64777_ _64777_/A _64778_/A sky130_fd_sc_hd__buf_2
X_61989_ _62002_/A _62002_/B _78064_/B _61989_/Y sky130_fd_sc_hd__nor3_4
X_69304_ _45915_/X _69305_/A sky130_fd_sc_hd__buf_2
X_54530_ _54475_/A _54530_/X sky130_fd_sc_hd__buf_2
X_85350_ _85959_/CLK _54938_/Y _85350_/Q sky130_fd_sc_hd__dfxtp_4
X_66516_ _82723_/D _79165_/B sky130_fd_sc_hd__inv_2
X_51742_ _52588_/A _51721_/X _54286_/C _53261_/D _51742_/X sky130_fd_sc_hd__and4_4
X_63728_ _64012_/A _63731_/D sky130_fd_sc_hd__buf_2
X_82562_ _82595_/CLK _82562_/D _78083_/A sky130_fd_sc_hd__dfxtp_4
X_67496_ _67495_/X _67496_/X sky130_fd_sc_hd__buf_2
XPHY_15 sky130_fd_sc_hd__decap_3
X_84301_ _84299_/CLK _84301_/D _80310_/B sky130_fd_sc_hd__dfxtp_4
XPHY_26 sky130_fd_sc_hd__decap_3
X_81513_ _82067_/CLK _81513_/D _75971_/A sky130_fd_sc_hd__dfxtp_4
X_69235_ _88044_/Q _69121_/X _69232_/X _69234_/X _69235_/X sky130_fd_sc_hd__a211o_4
X_54461_ _85438_/Q _54457_/X _54460_/Y _54461_/Y sky130_fd_sc_hd__o21ai_4
X_66447_ _66145_/X _66397_/X _66147_/X _66447_/Y sky130_fd_sc_hd__nand3_4
X_85281_ _85249_/CLK _85281_/D _56192_/C sky130_fd_sc_hd__dfxtp_4
X_51673_ _51657_/X _51684_/B _51684_/C _53196_/D _51673_/X sky130_fd_sc_hd__and4_4
XPHY_37 sky130_fd_sc_hd__decap_3
X_63659_ _63697_/A _58187_/A _63537_/C _63659_/X sky130_fd_sc_hd__and3_4
X_82493_ _82702_/CLK _82493_/D _78213_/B sky130_fd_sc_hd__dfxtp_4
XPHY_48 sky130_fd_sc_hd__decap_3
XPHY_59 sky130_fd_sc_hd__decap_3
X_56200_ _56255_/A _56200_/X sky130_fd_sc_hd__buf_2
X_87020_ _87026_/CLK _44644_/Y _87020_/Q sky130_fd_sc_hd__dfxtp_4
X_53412_ _53405_/X _54587_/B _53412_/Y sky130_fd_sc_hd__nand2_4
X_84232_ _85346_/CLK _84232_/D _81024_/D sky130_fd_sc_hd__dfxtp_4
X_50624_ _50624_/A _53844_/B _50624_/Y sky130_fd_sc_hd__nand2_4
X_81444_ _81412_/CLK _76674_/X _81412_/D sky130_fd_sc_hd__dfxtp_4
X_57180_ _57178_/Y _57179_/Y _57112_/X _57180_/Y sky130_fd_sc_hd__a21oi_4
X_69166_ _87537_/Q _68958_/X _69113_/X _69165_/X _69166_/X sky130_fd_sc_hd__a211o_4
X_54392_ _54378_/A _52700_/B _54392_/Y sky130_fd_sc_hd__nand2_4
X_66378_ _65307_/A _66433_/A sky130_fd_sc_hd__buf_2
X_56131_ _56131_/A _56140_/B _85291_/Q _56131_/Y sky130_fd_sc_hd__nand3_4
X_68117_ _66750_/X _66753_/X _68062_/X _68117_/Y sky130_fd_sc_hd__a21oi_4
X_53343_ _53339_/A _53330_/B _53330_/C _52831_/D _53343_/X sky130_fd_sc_hd__and4_4
X_65329_ _65325_/X _65328_/X _65277_/X _65333_/A sky130_fd_sc_hd__a21o_4
X_84163_ _84166_/CLK _66005_/X _84163_/Q sky130_fd_sc_hd__dfxtp_4
X_50555_ _86178_/Q _50499_/X _50554_/Y _50555_/Y sky130_fd_sc_hd__o21ai_4
X_81375_ _81362_/CLK _76933_/Y _81375_/Q sky130_fd_sc_hd__dfxtp_4
X_69097_ _87989_/Q _69007_/X _69051_/X _69096_/X _69097_/X sky130_fd_sc_hd__a211o_4
X_83114_ _83145_/CLK _83114_/D _70133_/A sky130_fd_sc_hd__dfxtp_4
X_56062_ _56058_/X _56060_/X _56061_/Y _85303_/D sky130_fd_sc_hd__o21ai_4
X_80326_ _80325_/X _80326_/X sky130_fd_sc_hd__buf_2
X_68048_ _86945_/Q _68023_/X _68024_/X _68047_/X _68049_/B sky130_fd_sc_hd__a211o_4
X_53274_ _51914_/A _53274_/B _53293_/C _52758_/D _53274_/X sky130_fd_sc_hd__and4_4
X_84094_ _80928_/CLK _66849_/X _80918_/D sky130_fd_sc_hd__dfxtp_4
X_50486_ _86191_/Q _50464_/X _50485_/Y _50486_/Y sky130_fd_sc_hd__o21ai_4
X_55013_ _55013_/A _55026_/B _55013_/C _55013_/D _55013_/X sky130_fd_sc_hd__and4_4
X_52225_ _52220_/A _48843_/B _52225_/Y sky130_fd_sc_hd__nand2_4
X_83045_ _83046_/CLK _74528_/Y _47031_/A sky130_fd_sc_hd__dfxtp_4
X_87922_ _87922_/CLK _87922_/D _87922_/Q sky130_fd_sc_hd__dfxtp_4
X_80257_ _80257_/A _80256_/X _80257_/Y sky130_fd_sc_hd__xnor2_4
X_70010_ _70048_/A _70010_/X sky130_fd_sc_hd__buf_2
X_59821_ _59805_/Y _59840_/A _59820_/Y _80422_/A _59814_/X _84694_/D
+ sky130_fd_sc_hd__o32a_4
X_52156_ _52156_/A _52140_/X _52156_/C _52156_/X sky130_fd_sc_hd__and3_4
X_87853_ _87068_/CLK _42474_/Y _73699_/A sky130_fd_sc_hd__dfxtp_4
X_80188_ _80184_/Y _80187_/Y _80198_/B sky130_fd_sc_hd__xor2_4
X_69999_ _69640_/Y _69916_/X _69984_/X _69998_/Y _69999_/X sky130_fd_sc_hd__a211o_4
X_51107_ _51112_/A _52799_/B _51107_/Y sky130_fd_sc_hd__nand2_4
X_86804_ _87995_/CLK _46031_/X _86804_/Q sky130_fd_sc_hd__dfxtp_4
X_59752_ _59752_/A _60312_/D sky130_fd_sc_hd__buf_2
X_52087_ _52083_/A _50385_/B _52087_/Y sky130_fd_sc_hd__nand2_4
X_56964_ _56940_/Y _56989_/A sky130_fd_sc_hd__buf_2
X_87784_ _87544_/CLK _42657_/Y _87784_/Q sky130_fd_sc_hd__dfxtp_4
X_84996_ _85005_/CLK _84996_/D _84996_/Q sky130_fd_sc_hd__dfxtp_4
X_58703_ _58703_/A _58703_/X sky130_fd_sc_hd__buf_2
X_51038_ _86085_/Q _51020_/X _51037_/Y _51038_/Y sky130_fd_sc_hd__o21ai_4
X_55915_ _55949_/A _55915_/B _55915_/X sky130_fd_sc_hd__and2_4
X_86735_ _86127_/CLK _86735_/D _86735_/Q sky130_fd_sc_hd__dfxtp_4
X_71961_ _71958_/Y _57592_/X _71960_/X _71961_/Y sky130_fd_sc_hd__a21oi_4
X_59683_ _59683_/A _59687_/C sky130_fd_sc_hd__inv_2
X_83947_ _83973_/CLK _83947_/D _80803_/D sky130_fd_sc_hd__dfxtp_4
X_56895_ _56893_/Y _56894_/Y _45888_/A _56895_/X sky130_fd_sc_hd__o21a_4
X_73700_ _41899_/Y _73529_/X _73698_/X _73699_/Y _73700_/X sky130_fd_sc_hd__a211o_4
X_58634_ _58634_/A _58649_/B _58634_/Y sky130_fd_sc_hd__nor2_4
X_70912_ _70908_/A _70913_/A sky130_fd_sc_hd__inv_2
X_43860_ _43859_/Y _87230_/D sky130_fd_sc_hd__inv_2
X_55846_ _44079_/X _55846_/B _55846_/X sky130_fd_sc_hd__and2_4
X_74680_ _74675_/X _56814_/A _74679_/Y _74680_/Y sky130_fd_sc_hd__o21ai_4
X_86666_ _86351_/CLK _86666_/D _86666_/Q sky130_fd_sc_hd__dfxtp_4
X_71892_ _71891_/Y _71892_/X sky130_fd_sc_hd__buf_2
X_83878_ _82558_/CLK _83878_/D _82558_/D sky130_fd_sc_hd__dfxtp_4
X_42811_ _42795_/X _42796_/X _41424_/X _87706_/Q _42805_/X _42812_/A
+ sky130_fd_sc_hd__o32ai_4
X_73631_ _73626_/X _73630_/X _56549_/X _73646_/B sky130_fd_sc_hd__a21o_4
X_85617_ _85630_/CLK _85617_/D _85617_/Q sky130_fd_sc_hd__dfxtp_4
X_70843_ _70862_/A _70860_/D sky130_fd_sc_hd__buf_2
X_58565_ _58676_/A _58614_/B sky130_fd_sc_hd__buf_2
X_82829_ _82462_/CLK _82829_/D _82829_/Q sky130_fd_sc_hd__dfxtp_4
X_43791_ _43776_/A _43791_/X sky130_fd_sc_hd__buf_2
X_55777_ _85194_/Q _55272_/X _55300_/X _55776_/X _55777_/X sky130_fd_sc_hd__a211o_4
X_86597_ _85957_/CLK _47796_/Y _72447_/A sky130_fd_sc_hd__dfxtp_4
X_52989_ _52997_/A _52997_/B _52997_/C _52989_/D _52989_/X sky130_fd_sc_hd__and4_4
X_45530_ _45452_/A _45530_/X sky130_fd_sc_hd__buf_2
X_57516_ _57497_/A _48207_/X _57516_/Y sky130_fd_sc_hd__nand2_4
X_76350_ _76330_/Y _76331_/Y _76332_/Y _76350_/X sky130_fd_sc_hd__o21a_4
X_88336_ _88337_/CLK _88336_/D _69612_/B sky130_fd_sc_hd__dfxtp_4
X_42742_ _42741_/Y _87742_/D sky130_fd_sc_hd__inv_2
X_54728_ _54724_/Y _54720_/X _54727_/X _54728_/Y sky130_fd_sc_hd__a21oi_4
X_73562_ _73378_/X _86241_/Q _73446_/X _73561_/X _73562_/X sky130_fd_sc_hd__a211o_4
X_85548_ _85837_/CLK _85548_/D _85548_/Q sky130_fd_sc_hd__dfxtp_4
X_70774_ _70862_/A _70791_/D sky130_fd_sc_hd__buf_2
X_58496_ _58492_/X _58493_/Y _58495_/Y _84835_/D sky130_fd_sc_hd__a21oi_4
X_75301_ _75299_/Y _75301_/B _75301_/X sky130_fd_sc_hd__xor2_4
X_72513_ _72512_/X _72513_/Y sky130_fd_sc_hd__inv_2
X_45461_ _55585_/B _45412_/X _45443_/X _45460_/Y _45461_/X sky130_fd_sc_hd__a211o_4
X_57447_ _57447_/A _57447_/Y sky130_fd_sc_hd__inv_2
X_76281_ _76281_/A _76282_/A sky130_fd_sc_hd__inv_2
X_88267_ _88267_/CLK _88267_/D _88267_/Q sky130_fd_sc_hd__dfxtp_4
X_54659_ _54655_/Y _54638_/X _54658_/X _85402_/D sky130_fd_sc_hd__a21oi_4
X_42673_ _42580_/A _42673_/X sky130_fd_sc_hd__buf_2
X_73493_ _44595_/Y _73491_/X _73492_/Y _73493_/X sky130_fd_sc_hd__a21o_4
X_85479_ _84926_/CLK _54238_/Y _85479_/Q sky130_fd_sc_hd__dfxtp_4
X_47200_ _82372_/Q _47201_/A sky130_fd_sc_hd__inv_2
X_78020_ _78021_/A _78021_/C _82176_/Q _78020_/Y sky130_fd_sc_hd__a21oi_4
X_44412_ _44363_/X _44412_/X sky130_fd_sc_hd__buf_2
X_75232_ _75223_/Y _75245_/A _75242_/A sky130_fd_sc_hd__xor2_4
X_87218_ _82906_/CLK _87218_/D _87218_/Q sky130_fd_sc_hd__dfxtp_4
X_41624_ _41624_/A _41624_/B _41624_/X sky130_fd_sc_hd__or2_4
X_48180_ _48174_/Y _48175_/X _48179_/Y _48180_/Y sky130_fd_sc_hd__a21boi_4
X_72444_ _83254_/Q _72381_/X _72438_/X _72443_/X _72444_/Y sky130_fd_sc_hd__a2bb2oi_4
X_45392_ _55635_/B _45388_/X _45390_/X _45391_/Y _45392_/X sky130_fd_sc_hd__a211o_4
X_57378_ _57377_/X _73916_/B sky130_fd_sc_hd__buf_2
X_88198_ _88201_/CLK _88198_/D _88198_/Q sky130_fd_sc_hd__dfxtp_4
X_47131_ _82379_/Q _54565_/D sky130_fd_sc_hd__inv_2
X_59117_ _59117_/A _86359_/Q _59117_/Y sky130_fd_sc_hd__nor2_4
X_44343_ _41693_/X _44326_/X _87156_/Q _44327_/X _87156_/D sky130_fd_sc_hd__a2bb2o_4
X_56329_ _56085_/X _56321_/X _56328_/Y _56329_/Y sky130_fd_sc_hd__o21ai_4
X_75163_ _75162_/X _75163_/X sky130_fd_sc_hd__buf_2
X_87149_ _87149_/CLK _44358_/X _87149_/Q sky130_fd_sc_hd__dfxtp_4
X_41555_ _41548_/X _82319_/Q _41554_/X _41555_/Y sky130_fd_sc_hd__o21ai_4
X_72375_ _72327_/X _85964_/Q _72374_/X _72375_/Y sky130_fd_sc_hd__o21ai_4
X_74114_ _74111_/X _74114_/B _74115_/B sky130_fd_sc_hd__nand2_4
X_40506_ _40504_/X _82314_/Q _40505_/X _40506_/Y sky130_fd_sc_hd__o21ai_4
X_59048_ _58877_/A _59048_/X sky130_fd_sc_hd__buf_2
X_47062_ _53345_/B _52833_/B sky130_fd_sc_hd__buf_2
X_71326_ _71196_/A _71335_/B sky130_fd_sc_hd__buf_2
X_44274_ _44120_/Y _44010_/A _72896_/B _44274_/D _44274_/X sky130_fd_sc_hd__and4_4
X_75094_ _80771_/Q _81027_/D _75094_/X sky130_fd_sc_hd__xor2_4
X_79971_ _84927_/Q _84175_/Q _79971_/X sky130_fd_sc_hd__or2_4
X_41486_ _41486_/A _41486_/X sky130_fd_sc_hd__buf_2
X_46013_ _40556_/A _46013_/X sky130_fd_sc_hd__buf_2
X_43225_ _40986_/X _43216_/X _87529_/Q _43218_/X _43225_/X sky130_fd_sc_hd__a2bb2o_4
X_78922_ _82847_/Q _82559_/Q _78923_/B sky130_fd_sc_hd__xnor2_4
X_74045_ _74045_/A _74045_/B _74046_/B sky130_fd_sc_hd__nand2_4
X_40437_ _44733_/A _40437_/X sky130_fd_sc_hd__buf_2
X_71257_ _50260_/B _71239_/A _71256_/Y _71257_/Y sky130_fd_sc_hd__o21ai_4
X_61010_ _60998_/X _60992_/X _60905_/Y _61010_/Y sky130_fd_sc_hd__o21ai_4
X_70208_ _70195_/X _74773_/C _70207_/X _83837_/D sky130_fd_sc_hd__a21o_4
Xclkbuf_10_582_0_CLK clkbuf_9_291_0_CLK/X _83973_/CLK sky130_fd_sc_hd__clkbuf_1
X_43156_ _43156_/A _43156_/Y sky130_fd_sc_hd__inv_2
X_78853_ _78865_/B _78852_/X _78866_/A sky130_fd_sc_hd__xnor2_4
X_40368_ _40420_/A _40368_/X sky130_fd_sc_hd__buf_2
X_71188_ _71191_/A _71189_/B sky130_fd_sc_hd__buf_2
X_42107_ _42106_/Y _88033_/D sky130_fd_sc_hd__inv_2
X_77804_ _77795_/X _77817_/A _77805_/B sky130_fd_sc_hd__xor2_4
X_70139_ _70139_/A _70139_/B _70139_/C _70139_/D _70154_/A sky130_fd_sc_hd__and4_4
X_47964_ _47904_/X _46389_/A _47963_/X _47965_/B sky130_fd_sc_hd__o21ai_4
X_43087_ _87581_/Q _43087_/Y sky130_fd_sc_hd__inv_2
X_78784_ _78784_/A _78784_/Y sky130_fd_sc_hd__inv_2
X_75996_ _81516_/Q _81740_/D _75996_/X sky130_fd_sc_hd__xor2_4
X_49703_ _49699_/A _52918_/B _49703_/Y sky130_fd_sc_hd__nand2_4
X_46915_ _46915_/A _46915_/X sky130_fd_sc_hd__buf_2
X_42038_ _42035_/X _42010_/X _40881_/X _42036_/Y _42037_/X _88062_/D
+ sky130_fd_sc_hd__o32ai_4
X_77735_ _77734_/Y _82259_/Q _78045_/A sky130_fd_sc_hd__nand2_4
X_62961_ _62988_/A _62988_/B _84366_/Q _62961_/Y sky130_fd_sc_hd__nor3_4
X_74947_ _74947_/A _74946_/X _74959_/A sky130_fd_sc_hd__nand2_4
X_47895_ _47887_/A _47895_/B _47895_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_597_0_CLK clkbuf_9_298_0_CLK/X _81928_/CLK sky130_fd_sc_hd__clkbuf_1
X_64700_ _64696_/X _85533_/Q _64697_/X _64699_/X _64700_/X sky130_fd_sc_hd__a211o_4
X_49634_ _49638_/A _52850_/B _49634_/Y sky130_fd_sc_hd__nand2_4
X_61912_ _61901_/X _61906_/X _61911_/Y _84742_/Q _61895_/X _61912_/Y
+ sky130_fd_sc_hd__o32ai_4
X_46846_ _82953_/Q _46846_/Y sky130_fd_sc_hd__inv_2
X_65680_ _65680_/A _65757_/A sky130_fd_sc_hd__buf_2
X_77666_ _77666_/A _77666_/B _77667_/C sky130_fd_sc_hd__or2_4
X_74878_ _74897_/B _74878_/B _74879_/B sky130_fd_sc_hd__xnor2_4
X_62892_ _62885_/X _62886_/X _62888_/Y _62889_/Y _62891_/X _62892_/X
+ sky130_fd_sc_hd__a41o_4
X_79405_ _84351_/Q _79405_/B _79405_/X sky130_fd_sc_hd__xor2_4
X_64631_ _64684_/A _86464_/Q _64631_/X sky130_fd_sc_hd__and2_4
X_76617_ _76614_/C _76602_/Y _76614_/B _76624_/B sky130_fd_sc_hd__a21bo_4
X_49565_ _49561_/A _49561_/B _49548_/X _52779_/D _49565_/X sky130_fd_sc_hd__and4_4
X_73829_ _73709_/X _73829_/X sky130_fd_sc_hd__buf_2
X_61843_ _61417_/B _61843_/B _61795_/C _61778_/X _61843_/Y sky130_fd_sc_hd__nand4_4
X_46777_ _46772_/Y _46751_/X _46776_/X _86705_/D sky130_fd_sc_hd__a21oi_4
X_77597_ _81946_/Q _82202_/D _81914_/D sky130_fd_sc_hd__xor2_4
X_43989_ _43985_/X _43988_/X _43989_/Y sky130_fd_sc_hd__nand2_4
X_48516_ _86515_/Q _48478_/X _48515_/Y _48516_/Y sky130_fd_sc_hd__o21ai_4
X_67350_ _87167_/Q _67348_/X _67278_/X _67349_/X _67350_/X sky130_fd_sc_hd__a211o_4
X_79336_ _79322_/Y _79336_/B _79336_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_520_0_CLK clkbuf_9_260_0_CLK/X _81433_/CLK sky130_fd_sc_hd__clkbuf_1
X_45728_ _45728_/A _45746_/B _45728_/Y sky130_fd_sc_hd__nand2_4
X_64562_ _45924_/A _64665_/A sky130_fd_sc_hd__buf_2
X_76548_ _76548_/A _76547_/Y _76548_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_6_11_0_CLK clkbuf_5_5_0_CLK/X clkbuf_7_23_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_49496_ _49496_/A _49496_/X sky130_fd_sc_hd__buf_2
X_61774_ _62185_/B _61794_/B sky130_fd_sc_hd__buf_2
X_66301_ _66326_/A _66301_/B _66301_/X sky130_fd_sc_hd__and2_4
X_63513_ _61479_/B _63487_/X _63511_/X _63512_/X _63513_/X sky130_fd_sc_hd__a211o_4
X_60725_ _60725_/A _60725_/B _60725_/Y sky130_fd_sc_hd__nor2_4
X_48447_ _72993_/B _48419_/X _48446_/Y _48447_/Y sky130_fd_sc_hd__o21ai_4
X_67281_ _67277_/X _67280_/X _67255_/X _67281_/Y sky130_fd_sc_hd__a21oi_4
X_79267_ _79267_/A _79267_/B _79276_/B sky130_fd_sc_hd__xor2_4
X_45659_ _45659_/A _45659_/Y sky130_fd_sc_hd__inv_2
X_76479_ _76474_/X _76479_/B _76479_/C _76513_/C sky130_fd_sc_hd__nand3_4
X_64493_ _64363_/A _64363_/B _58187_/A _61145_/X _64493_/X sky130_fd_sc_hd__and4_4
X_69020_ _83951_/Q _68954_/X _69019_/X _83951_/D sky130_fd_sc_hd__a21bo_4
X_66232_ _66231_/X _66151_/B _80397_/B _66232_/X sky130_fd_sc_hd__and3_4
X_78218_ _82677_/Q _78218_/B _78218_/X sky130_fd_sc_hd__xor2_4
X_63444_ _64282_/A _63465_/B _63465_/C _63465_/D _63444_/Y sky130_fd_sc_hd__nand4_4
X_48378_ _48370_/Y _48302_/X _48377_/X _48378_/Y sky130_fd_sc_hd__a21oi_4
X_60656_ _60702_/C _60713_/A sky130_fd_sc_hd__buf_2
X_79198_ _79198_/A _79198_/B _79198_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_535_0_CLK clkbuf_9_267_0_CLK/X _81507_/CLK sky130_fd_sc_hd__clkbuf_1
X_47329_ _47329_/A _52989_/D sky130_fd_sc_hd__buf_2
X_66163_ _84152_/Q _66164_/C sky130_fd_sc_hd__inv_2
Xclkbuf_6_26_0_CLK clkbuf_6_27_0_CLK/A clkbuf_6_26_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_78149_ _82571_/Q _82483_/Q _78149_/Y sky130_fd_sc_hd__nand2_4
X_63375_ _63375_/A _63400_/A sky130_fd_sc_hd__buf_2
X_60587_ _79133_/A _60577_/X _60586_/X _60563_/X _60587_/Y sky130_fd_sc_hd__a2bb2oi_4
X_65114_ _65112_/Y _65070_/X _65113_/X _65114_/X sky130_fd_sc_hd__a21o_4
X_50340_ _50336_/Y _50313_/X _50339_/X _86221_/D sky130_fd_sc_hd__a21oi_4
X_62326_ _62315_/X _62322_/Y _62325_/X _58177_/A _62300_/X _62326_/Y
+ sky130_fd_sc_hd__o32ai_4
X_81160_ _81160_/CLK _74890_/B _40518_/B sky130_fd_sc_hd__dfxtp_4
X_66094_ _65992_/A _66094_/B _66094_/X sky130_fd_sc_hd__and2_4
X_80111_ _60064_/C _80111_/B _80121_/B sky130_fd_sc_hd__xor2_4
X_65045_ _65045_/A _65047_/B sky130_fd_sc_hd__buf_2
X_69922_ _69919_/X _69921_/X _68470_/X _69922_/X sky130_fd_sc_hd__a21o_4
X_50271_ _50269_/Y _50243_/X _50270_/X _50271_/Y sky130_fd_sc_hd__a21oi_4
X_62257_ _62478_/A _59995_/A _64246_/B _60025_/X _62257_/X sky130_fd_sc_hd__and4_4
X_81091_ _82084_/CLK _79893_/X _81091_/Q sky130_fd_sc_hd__dfxtp_4
X_52010_ _85906_/Q _51945_/X _52009_/Y _52010_/Y sky130_fd_sc_hd__o21ai_4
X_61208_ _61195_/A _61207_/X _61086_/X _61208_/Y sky130_fd_sc_hd__o21ai_4
X_80042_ _80042_/A _80041_/Y _80052_/B sky130_fd_sc_hd__xor2_4
X_69853_ _69853_/A _88318_/Q _69853_/X sky130_fd_sc_hd__and2_4
X_62188_ _61715_/A _62188_/B _62188_/C _62187_/Y _62188_/Y sky130_fd_sc_hd__nand4_4
X_68804_ _68366_/X _43641_/Y _68804_/Y sky130_fd_sc_hd__nor2_4
X_84850_ _84732_/CLK _84850_/D _84850_/Q sky130_fd_sc_hd__dfxtp_4
X_61139_ _60933_/X _61238_/B _61110_/Y _61131_/Y _61138_/Y _61139_/Y
+ sky130_fd_sc_hd__a41oi_4
X_69784_ _87055_/Q _69664_/X _69665_/X _69783_/X _69785_/B sky130_fd_sc_hd__a211o_4
X_66996_ _87873_/Q _66994_/X _66926_/X _66995_/X _66996_/X sky130_fd_sc_hd__a211o_4
X_83801_ _83819_/CLK _70314_/X _74808_/B sky130_fd_sc_hd__dfxtp_4
X_68735_ _68735_/A _68735_/B _68735_/X sky130_fd_sc_hd__and2_4
X_53961_ _53942_/A _46295_/A _53961_/Y sky130_fd_sc_hd__nand2_4
X_65947_ _65934_/X _73638_/B _65947_/X sky130_fd_sc_hd__and2_4
X_84781_ _83438_/CLK _84781_/D _58983_/A sky130_fd_sc_hd__dfxtp_4
X_81993_ _81989_/CLK _81993_/D _77054_/A sky130_fd_sc_hd__dfxtp_4
X_55700_ _55700_/A _55700_/B _55701_/A sky130_fd_sc_hd__and2_4
X_86520_ _83584_/CLK _86520_/D _73016_/B sky130_fd_sc_hd__dfxtp_4
X_52912_ _52895_/A _52916_/B _52900_/C _51220_/D _52912_/X sky130_fd_sc_hd__and4_4
X_83732_ _84930_/CLK _83732_/D _83732_/Q sky130_fd_sc_hd__dfxtp_4
X_56680_ _56680_/A _56684_/B sky130_fd_sc_hd__buf_2
X_80944_ _80849_/CLK _80944_/D _80944_/Q sky130_fd_sc_hd__dfxtp_4
X_68666_ _69146_/A _68666_/X sky130_fd_sc_hd__buf_2
X_53892_ _53773_/A _53892_/X sky130_fd_sc_hd__buf_2
X_65878_ _65878_/A _86467_/Q _65878_/X sky130_fd_sc_hd__and2_4
X_55631_ _44085_/C _85152_/Q _55631_/X sky130_fd_sc_hd__and2_4
X_67617_ _87463_/Q _67594_/X _67595_/X _67616_/X _67617_/X sky130_fd_sc_hd__a211o_4
X_86451_ _85555_/CLK _86451_/D _64992_/B sky130_fd_sc_hd__dfxtp_4
X_52843_ _52843_/A _52843_/B _52843_/Y sky130_fd_sc_hd__nand2_4
X_64829_ _64829_/A _64829_/X sky130_fd_sc_hd__buf_2
X_83663_ _83663_/CLK _83663_/D _46861_/A sky130_fd_sc_hd__dfxtp_4
X_80875_ _80754_/CLK _75655_/B _80875_/Q sky130_fd_sc_hd__dfxtp_4
X_68597_ _68597_/A _68596_/X _68597_/Y sky130_fd_sc_hd__nand2_4
X_85402_ _83745_/CLK _85402_/D _85402_/Q sky130_fd_sc_hd__dfxtp_4
X_58350_ _58350_/A _58350_/Y sky130_fd_sc_hd__inv_2
X_82614_ _82617_/CLK _78994_/B _82614_/Q sky130_fd_sc_hd__dfxtp_4
X_55562_ _55559_/X _55561_/X _44113_/X _55562_/X sky130_fd_sc_hd__a21o_4
X_67548_ _87466_/Q _67476_/X _67477_/X _67547_/X _67548_/X sky130_fd_sc_hd__a211o_4
X_86382_ _86384_/CLK _86382_/D _58804_/B sky130_fd_sc_hd__dfxtp_4
X_52774_ _85757_/Q _52765_/X _52773_/Y _52774_/Y sky130_fd_sc_hd__o21ai_4
X_83594_ _83594_/CLK _71134_/Y _49195_/A sky130_fd_sc_hd__dfxtp_4
X_57301_ _57280_/X _57297_/X _57298_/Y _57300_/Y _57302_/A sky130_fd_sc_hd__a211o_4
X_88121_ _88121_/CLK _88121_/D _67206_/B sky130_fd_sc_hd__dfxtp_4
X_54513_ _54486_/A _54518_/A sky130_fd_sc_hd__buf_2
X_85333_ _83627_/CLK _55027_/Y _85333_/Q sky130_fd_sc_hd__dfxtp_4
X_51725_ _85957_/Q _51701_/X _51724_/Y _51725_/Y sky130_fd_sc_hd__o21ai_4
X_58281_ _58271_/X _83409_/Q _58280_/Y _58281_/X sky130_fd_sc_hd__o21a_4
X_82545_ _83133_/CLK _82545_/D _82545_/Q sky130_fd_sc_hd__dfxtp_4
X_55493_ _44061_/X _45581_/Y _55493_/Y sky130_fd_sc_hd__nor2_4
X_67479_ _87405_/Q _67476_/X _67477_/X _67478_/X _67479_/X sky130_fd_sc_hd__a211o_4
X_57232_ _55211_/B _57192_/A _57230_/Y _57231_/X _85058_/D sky130_fd_sc_hd__a211o_4
X_69218_ _69191_/A _69218_/B _69218_/X sky130_fd_sc_hd__and2_4
X_88052_ _88085_/CLK _42064_/Y _42063_/A sky130_fd_sc_hd__dfxtp_4
X_54444_ _54435_/A _54440_/B _54429_/C _46924_/Y _54444_/X sky130_fd_sc_hd__and4_4
X_85264_ _85167_/CLK _85264_/D _85264_/Q sky130_fd_sc_hd__dfxtp_4
X_51656_ _52620_/A _52593_/A sky130_fd_sc_hd__buf_2
X_70490_ _58372_/Y _70458_/X _70489_/Y _83762_/D sky130_fd_sc_hd__o21ai_4
X_82476_ _82498_/CLK _78454_/X _78088_/B sky130_fd_sc_hd__dfxtp_4
X_87003_ _86984_/CLK _44678_/Y _87003_/Q sky130_fd_sc_hd__dfxtp_4
X_84215_ _84220_/CLK _84215_/D _84215_/Q sky130_fd_sc_hd__dfxtp_4
X_50607_ _50607_/A _52307_/B _50607_/Y sky130_fd_sc_hd__nand2_4
X_57163_ _57170_/A _56737_/X _57163_/C _57156_/X _57163_/Y sky130_fd_sc_hd__nand4_4
X_81427_ _83926_/CLK _81459_/Q _76041_/B sky130_fd_sc_hd__dfxtp_4
X_69149_ _45915_/X _69755_/A sky130_fd_sc_hd__buf_2
X_54375_ _54034_/A _54376_/A sky130_fd_sc_hd__buf_2
X_85195_ _80671_/CLK _85195_/D _85195_/Q sky130_fd_sc_hd__dfxtp_4
X_51587_ _51694_/A _51603_/B sky130_fd_sc_hd__buf_2
X_56114_ _56114_/A _56114_/X sky130_fd_sc_hd__buf_2
X_41340_ _41242_/X _82903_/Q _41339_/X _41340_/X sky130_fd_sc_hd__o21a_4
X_53326_ _53332_/A _47023_/Y _53326_/Y sky130_fd_sc_hd__nand2_4
X_72160_ _59238_/X _72160_/B _72160_/Y sky130_fd_sc_hd__nor2_4
X_84146_ _84231_/CLK _84146_/D _66247_/C sky130_fd_sc_hd__dfxtp_4
X_50538_ _50538_/A _50552_/C sky130_fd_sc_hd__buf_2
X_57094_ _57093_/Y _57192_/A sky130_fd_sc_hd__buf_2
X_81358_ _81492_/CLK _81358_/D _81358_/Q sky130_fd_sc_hd__dfxtp_4
X_71111_ _50674_/B _71095_/A _71110_/Y _71111_/Y sky130_fd_sc_hd__o21ai_4
X_56045_ _55997_/X _74312_/C _74310_/C _56044_/X _56045_/Y sky130_fd_sc_hd__nand4_4
X_80309_ _80308_/B _80309_/Y sky130_fd_sc_hd__inv_2
X_41271_ _41255_/X _81124_/Q _41270_/X _41271_/Y sky130_fd_sc_hd__o21ai_4
X_53257_ _53243_/X _51747_/A _53266_/C _53257_/D _53257_/X sky130_fd_sc_hd__and4_4
X_72091_ _72052_/A _72091_/X sky130_fd_sc_hd__buf_2
X_84077_ _82067_/CLK _67258_/X _80901_/D sky130_fd_sc_hd__dfxtp_4
X_50469_ _50469_/A _50492_/B _50497_/C _50469_/X sky130_fd_sc_hd__and3_4
X_81289_ _81603_/CLK _76977_/X _81257_/D sky130_fd_sc_hd__dfxtp_4
X_43010_ _40542_/X _51934_/A _67285_/B _42634_/A _87605_/D sky130_fd_sc_hd__a2bb2o_4
X_52208_ _52188_/A _50503_/B _52208_/Y sky130_fd_sc_hd__nand2_4
X_71042_ _71026_/A _71276_/C sky130_fd_sc_hd__buf_2
X_83028_ _85269_/CLK _74579_/Y _45107_/A sky130_fd_sc_hd__dfxtp_4
X_87905_ _87646_/CLK _87905_/D _87905_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_9_0_CLK clkbuf_8_9_0_CLK/A clkbuf_8_9_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_53188_ _85680_/Q _53172_/X _53187_/Y _53188_/Y sky130_fd_sc_hd__o21ai_4
X_59804_ _80455_/A _59803_/X _59631_/Y _59804_/X sky130_fd_sc_hd__a21bo_4
X_52139_ _52139_/A _52198_/A sky130_fd_sc_hd__buf_2
X_75850_ _75850_/A _75849_/Y _75850_/Y sky130_fd_sc_hd__nand2_4
X_87836_ _87834_/CLK _87836_/D _42518_/A sky130_fd_sc_hd__dfxtp_4
X_57996_ _84933_/Q _57996_/Y sky130_fd_sc_hd__inv_2
X_74801_ _71266_/X _74801_/B _71846_/A _70500_/B _74801_/X sky130_fd_sc_hd__and4_4
X_59735_ _65515_/A _59842_/A sky130_fd_sc_hd__buf_2
X_44961_ _85213_/Q _44945_/X _44960_/X _44961_/Y sky130_fd_sc_hd__o21ai_4
X_56947_ _56940_/Y _56947_/X sky130_fd_sc_hd__buf_2
X_75781_ _75769_/Y _75781_/Y sky130_fd_sc_hd__inv_2
X_87767_ _87767_/CLK _42693_/X _69521_/B sky130_fd_sc_hd__dfxtp_4
X_72993_ _73186_/A _72993_/B _72993_/X sky130_fd_sc_hd__and2_4
X_84979_ _86549_/CLK _84979_/D _84979_/Q sky130_fd_sc_hd__dfxtp_4
X_46700_ _46700_/A _54314_/B sky130_fd_sc_hd__inv_2
X_77520_ _77516_/X _77520_/B _77520_/X sky130_fd_sc_hd__xor2_4
X_43912_ _43895_/X _43902_/X _41376_/X _67752_/B _43897_/X _43913_/A
+ sky130_fd_sc_hd__o32ai_4
X_74732_ _70192_/Y _70692_/C _83834_/Q _74731_/X _74732_/X sky130_fd_sc_hd__a2bb2o_4
X_86718_ _86398_/CLK _46648_/Y _58601_/A sky130_fd_sc_hd__dfxtp_4
X_47680_ _47696_/A _53183_/B _47680_/Y sky130_fd_sc_hd__nand2_4
X_71944_ _71942_/Y _83320_/Q _71943_/Y _71944_/X sky130_fd_sc_hd__a21o_4
X_59666_ _59666_/A _59687_/B sky130_fd_sc_hd__inv_2
X_44892_ _44891_/X _44892_/X sky130_fd_sc_hd__buf_2
X_56878_ _56877_/X _56878_/Y sky130_fd_sc_hd__inv_2
X_87698_ _87950_/CLK _42826_/X _87698_/Q sky130_fd_sc_hd__dfxtp_4
X_46631_ _46670_/A _46647_/B _46659_/C _51756_/D _46631_/X sky130_fd_sc_hd__and4_4
X_58617_ _58591_/X _85469_/Q _58616_/X _58617_/Y sky130_fd_sc_hd__o21ai_4
X_77451_ _77433_/Y _77439_/Y _77431_/Y _77451_/X sky130_fd_sc_hd__o21a_4
X_43843_ _43802_/A _43843_/X sky130_fd_sc_hd__buf_2
X_55829_ _55802_/X _55811_/X _56108_/A _55828_/X _55830_/A sky130_fd_sc_hd__and4_4
X_74663_ _82992_/Q _74641_/X _74662_/Y _74664_/A sky130_fd_sc_hd__o21ai_4
X_86649_ _86647_/CLK _86649_/D _57846_/A sky130_fd_sc_hd__dfxtp_4
X_71875_ _71871_/X _83345_/Q _71874_/Y _71875_/X sky130_fd_sc_hd__a21o_4
X_59597_ _59557_/X _59564_/B _59544_/D _60630_/A sky130_fd_sc_hd__nand3_4
X_76402_ _76401_/X _76403_/B sky130_fd_sc_hd__inv_2
X_49350_ _48917_/X _52565_/B _49350_/Y sky130_fd_sc_hd__nand2_4
X_73614_ _73614_/A _73614_/X sky130_fd_sc_hd__buf_2
X_70826_ _52918_/B _70802_/A _70825_/Y _83690_/D sky130_fd_sc_hd__o21ai_4
X_46562_ _46557_/Y _46523_/X _46561_/Y _86726_/D sky130_fd_sc_hd__a21boi_4
X_58548_ _58548_/A _58548_/B _58548_/Y sky130_fd_sc_hd__nor2_4
X_77382_ _77382_/A _77382_/B _77381_/Y _77382_/X sky130_fd_sc_hd__or3_4
X_43774_ _43774_/A _43774_/X sky130_fd_sc_hd__buf_2
X_74594_ _74591_/X _74583_/X _56109_/A _74584_/X _74594_/X sky130_fd_sc_hd__a211o_4
X_40986_ _40985_/Y _40986_/X sky130_fd_sc_hd__buf_2
X_48301_ _86539_/Q _48263_/X _48300_/Y _48301_/Y sky130_fd_sc_hd__o21ai_4
X_79121_ _78804_/B _82498_/D sky130_fd_sc_hd__inv_2
X_45513_ _45511_/X _61421_/A _45452_/X _45513_/Y sky130_fd_sc_hd__o21ai_4
X_76333_ _76332_/Y _76333_/Y sky130_fd_sc_hd__inv_2
X_88319_ _88056_/CLK _88319_/D _69842_/B sky130_fd_sc_hd__dfxtp_4
X_42725_ _42725_/A _42725_/Y sky130_fd_sc_hd__inv_2
X_49281_ _49405_/A _49281_/X sky130_fd_sc_hd__buf_2
X_73545_ _73543_/X _73532_/X _73534_/X _73545_/Y sky130_fd_sc_hd__nand3_4
X_46493_ _48606_/A _46493_/X sky130_fd_sc_hd__buf_2
X_70757_ _70416_/Y _70758_/C sky130_fd_sc_hd__buf_2
X_58479_ _58467_/X _58476_/Y _58478_/Y _84839_/D sky130_fd_sc_hd__a21oi_4
X_48232_ _86551_/Q _48188_/X _48231_/Y _48232_/Y sky130_fd_sc_hd__o21ai_4
X_60510_ _63252_/B _60570_/B _60627_/A _60626_/A _60509_/Y _60510_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_79052_ _79053_/B _79053_/A _79055_/A sky130_fd_sc_hd__nor2_4
X_45444_ _45444_/A _45397_/X _45444_/Y sky130_fd_sc_hd__nor2_4
X_76264_ _76264_/A _76264_/Y sky130_fd_sc_hd__inv_2
X_42656_ _42647_/X _42648_/X _40994_/X _87784_/Q _42637_/X _42657_/A
+ sky130_fd_sc_hd__o32ai_4
X_61490_ _84820_/Q _61490_/X sky130_fd_sc_hd__buf_2
X_73476_ _73476_/A _86501_/Q _73476_/X sky130_fd_sc_hd__and2_4
X_70688_ _71887_/A _70689_/A sky130_fd_sc_hd__buf_2
X_78003_ _78003_/A _78003_/Y sky130_fd_sc_hd__inv_2
X_75215_ _75212_/Y _75233_/B _75216_/A sky130_fd_sc_hd__xor2_4
X_41607_ _40567_/A _41607_/X sky130_fd_sc_hd__buf_2
X_60441_ _60439_/X _60441_/B _60440_/X _60442_/C sky130_fd_sc_hd__and3_4
X_72427_ _72414_/X _72427_/B _72427_/Y sky130_fd_sc_hd__nor2_4
X_48163_ _48186_/A _48163_/X sky130_fd_sc_hd__buf_2
X_45375_ _55738_/B _45357_/X _45339_/X _45375_/X sky130_fd_sc_hd__o21a_4
X_76195_ _76192_/X _76196_/B _76194_/Y _76195_/X sky130_fd_sc_hd__a21o_4
X_42587_ _42573_/X _42574_/X _40854_/X _69790_/A _42580_/X _42588_/A
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_4_1_1_CLK clkbuf_4_1_0_CLK/X clkbuf_5_2_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_47114_ _47110_/Y _47081_/X _47113_/X _86669_/D sky130_fd_sc_hd__a21oi_4
X_44326_ _40409_/X _44326_/X sky130_fd_sc_hd__buf_2
X_63160_ _60489_/X _63161_/C sky130_fd_sc_hd__buf_2
X_75146_ _75145_/Y _75146_/Y sky130_fd_sc_hd__inv_2
X_41538_ _41489_/X _41490_/X _41536_/X _66932_/B _41537_/X _41538_/Y
+ sky130_fd_sc_hd__o32ai_4
X_48094_ _48094_/A _48642_/B sky130_fd_sc_hd__inv_2
X_60372_ _60331_/D _60331_/B _60224_/Y _60371_/X _57703_/X _60372_/Y
+ sky130_fd_sc_hd__o32ai_4
X_72358_ _72358_/A _72358_/X sky130_fd_sc_hd__buf_2
X_62111_ _59692_/Y _62161_/B sky130_fd_sc_hd__buf_2
X_47045_ _46903_/A _47048_/C sky130_fd_sc_hd__buf_2
X_71309_ _71196_/A _71314_/B sky130_fd_sc_hd__buf_2
X_44257_ _43948_/B _44254_/X _44227_/Y _44218_/X _44258_/A sky130_fd_sc_hd__o22a_4
X_63091_ _60508_/A _63092_/D sky130_fd_sc_hd__buf_2
X_75077_ _75076_/Y _75077_/Y sky130_fd_sc_hd__inv_2
X_79954_ _84926_/Q _84174_/Q _79957_/C sky130_fd_sc_hd__nand2_4
X_41469_ _41468_/Y _41469_/X sky130_fd_sc_hd__buf_2
X_72289_ _72264_/X _85363_/Q _72288_/X _72289_/Y sky130_fd_sc_hd__o21ai_4
X_62042_ _61570_/B _62007_/X _62149_/C _62008_/X _62047_/B sky130_fd_sc_hd__nand4_4
X_43208_ _43196_/X _43207_/X _40950_/X _87537_/Q _43172_/X _43209_/A
+ sky130_fd_sc_hd__o32ai_4
X_74028_ _74026_/X _74028_/B _74028_/C _74028_/Y sky130_fd_sc_hd__nand3_4
X_78905_ _78892_/B _82508_/D sky130_fd_sc_hd__inv_2
X_44188_ _72720_/A _72806_/A sky130_fd_sc_hd__buf_2
X_79885_ _81024_/D _83280_/Q _79885_/Y sky130_fd_sc_hd__nand2_4
X_43139_ _43100_/X _43110_/X _40814_/X _73036_/A _43121_/X _43140_/A
+ sky130_fd_sc_hd__o32ai_4
X_66850_ _66971_/A _66850_/X sky130_fd_sc_hd__buf_2
X_78836_ _78835_/Y _78830_/A _78829_/A _78837_/B sky130_fd_sc_hd__o21ai_4
X_48996_ _48996_/A _49009_/B _48996_/Y sky130_fd_sc_hd__nor2_4
X_65801_ _84177_/Q _65802_/C sky130_fd_sc_hd__inv_2
X_47947_ _47942_/Y _47903_/X _47946_/X _47947_/Y sky130_fd_sc_hd__a21oi_4
X_66781_ _80921_/D _66734_/X _66780_/X _84097_/D sky130_fd_sc_hd__a21bo_4
X_78767_ _78764_/Y _78767_/B _78765_/Y _78767_/Y sky130_fd_sc_hd__nand3_4
X_75979_ _75963_/C _75975_/Y _75978_/Y _75980_/B sky130_fd_sc_hd__o21a_4
X_63993_ _63985_/X _63969_/X _63987_/Y _63990_/Y _63992_/X _63993_/X
+ sky130_fd_sc_hd__a41o_4
X_68520_ _66053_/A _68520_/B _68520_/Y sky130_fd_sc_hd__nor2_4
X_65732_ _65654_/X _86189_/Q _65576_/X _65731_/X _65732_/X sky130_fd_sc_hd__a211o_4
X_77718_ _77718_/A _77718_/B _77723_/A sky130_fd_sc_hd__nand2_4
X_62944_ _62941_/X _62942_/X _62943_/Y _84368_/D sky130_fd_sc_hd__a21oi_4
X_47878_ _48196_/A _49312_/C _53697_/C _47878_/X sky130_fd_sc_hd__and3_4
X_78698_ _78693_/X _78696_/Y _78694_/Y _78722_/A sky130_fd_sc_hd__nand3_4
X_49617_ _49607_/X _52833_/B _49617_/Y sky130_fd_sc_hd__nand2_4
X_68451_ _68451_/A _68452_/A sky130_fd_sc_hd__buf_2
X_46829_ _46828_/Y _52698_/D sky130_fd_sc_hd__buf_2
X_65663_ _65659_/X _65663_/B _65662_/X _65663_/Y sky130_fd_sc_hd__nand3_4
X_77649_ _77648_/Y _77650_/B sky130_fd_sc_hd__inv_2
X_62875_ _60335_/Y _62875_/X sky130_fd_sc_hd__buf_2
X_67402_ _67397_/X _67400_/X _67401_/X _67402_/Y sky130_fd_sc_hd__a21oi_4
X_64614_ _65117_/A _64615_/A sky130_fd_sc_hd__buf_2
X_61826_ _59605_/Y _61839_/C sky130_fd_sc_hd__buf_2
X_49548_ _49548_/A _49548_/X sky130_fd_sc_hd__buf_2
X_80660_ _80657_/CLK _74826_/Y _46111_/B sky130_fd_sc_hd__dfxtp_4
X_68382_ _88114_/Q _68377_/X _68379_/X _68381_/Y _68382_/X sky130_fd_sc_hd__a211o_4
X_65594_ _65591_/X _65593_/X _65457_/X _65599_/A sky130_fd_sc_hd__a21o_4
X_79319_ _79309_/X _79311_/B _79318_/Y _79336_/B sky130_fd_sc_hd__a21boi_4
X_67333_ _67333_/A _67333_/B _67333_/X sky130_fd_sc_hd__and2_4
X_64545_ _64545_/A _64545_/B _64545_/C _64545_/X sky130_fd_sc_hd__and3_4
X_49479_ _49467_/A _49500_/B _49467_/C _52694_/D _49479_/X sky130_fd_sc_hd__and4_4
X_61757_ _61730_/X _61791_/B _61732_/X _63030_/B _61757_/X sky130_fd_sc_hd__and4_4
X_80591_ _80617_/A _80601_/A sky130_fd_sc_hd__inv_2
X_51510_ _51508_/Y _51503_/X _51509_/X _85997_/D sky130_fd_sc_hd__a21oi_4
X_82330_ _82284_/CLK _77178_/B _82330_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_474_0_CLK clkbuf_9_237_0_CLK/X _86701_/CLK sky130_fd_sc_hd__clkbuf_1
X_60708_ _60712_/B _60694_/C _60711_/A _60660_/A _60708_/Y sky130_fd_sc_hd__nand4_4
X_67264_ _67025_/X _67264_/X sky130_fd_sc_hd__buf_2
X_52490_ _52476_/A _46411_/A _52490_/Y sky130_fd_sc_hd__nand2_4
X_64476_ _61232_/X _61607_/B _61207_/X _64477_/D sky130_fd_sc_hd__nand3_4
X_61688_ _61688_/A _61688_/Y sky130_fd_sc_hd__inv_2
X_69003_ _69000_/X _69002_/X _68390_/X _69003_/X sky130_fd_sc_hd__a21o_4
X_66215_ _57761_/X _84972_/Q _65309_/X _66214_/X _66216_/C sky130_fd_sc_hd__a211o_4
X_51441_ _86009_/Q _51429_/X _51440_/Y _51441_/Y sky130_fd_sc_hd__o21ai_4
X_63427_ _63427_/A _61811_/X _63427_/X sky130_fd_sc_hd__and2_4
X_82261_ _82253_/CLK _82261_/D _82261_/Q sky130_fd_sc_hd__dfxtp_4
X_60639_ _60639_/A _61075_/C sky130_fd_sc_hd__buf_2
X_67195_ _67149_/A _88185_/Q _67195_/X sky130_fd_sc_hd__and2_4
X_84000_ _81755_/CLK _68253_/X _82648_/D sky130_fd_sc_hd__dfxtp_4
X_81212_ _82284_/CLK _74853_/X _46318_/A sky130_fd_sc_hd__dfxtp_4
X_54160_ _54160_/A _54160_/B _54146_/X _52993_/D _54160_/X sky130_fd_sc_hd__and4_4
X_66146_ _66011_/X _86545_/Q _66146_/X sky130_fd_sc_hd__and2_4
X_51372_ _51367_/X _51372_/B _51372_/X sky130_fd_sc_hd__and2_4
X_63358_ _63357_/X _63358_/X sky130_fd_sc_hd__buf_2
X_82192_ _82386_/CLK _82192_/D _82192_/Q sky130_fd_sc_hd__dfxtp_4
X_53111_ _53111_/A _53111_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_489_0_CLK clkbuf_9_244_0_CLK/X _85961_/CLK sky130_fd_sc_hd__clkbuf_1
X_50323_ _50319_/Y _50299_/X _50322_/Y _86224_/D sky130_fd_sc_hd__a21boi_4
X_62309_ _61399_/X _62309_/B _62309_/C _62211_/D _62310_/D sky130_fd_sc_hd__nand4_4
X_81143_ _86758_/CLK _81143_/D _40644_/A sky130_fd_sc_hd__dfxtp_4
X_54091_ _54091_/A _54043_/B _51749_/X _54091_/X sky130_fd_sc_hd__and3_4
X_66077_ _66068_/X _65599_/Y _66076_/Y _66077_/Y sky130_fd_sc_hd__o21ai_4
X_63289_ _60502_/Y _63289_/X sky130_fd_sc_hd__buf_2
X_53042_ _85708_/Q _53038_/X _53041_/Y _53042_/Y sky130_fd_sc_hd__o21ai_4
X_69905_ _83888_/Q _69894_/X _69904_/X _69905_/X sky130_fd_sc_hd__a21bo_4
X_65028_ _64772_/A _65028_/X sky130_fd_sc_hd__buf_2
X_50254_ _74458_/A _54043_/B sky130_fd_sc_hd__buf_2
X_85951_ _85514_/CLK _51762_/Y _85951_/Q sky130_fd_sc_hd__dfxtp_4
X_81074_ _81074_/CLK _75574_/A _75299_/A sky130_fd_sc_hd__dfxtp_4
X_80025_ _80019_/A _80018_/X _80024_/Y _80025_/Y sky130_fd_sc_hd__a21boi_4
X_84902_ _84360_/CLK _84902_/D _63400_/B sky130_fd_sc_hd__dfxtp_4
X_57850_ _57824_/X _85497_/Q _57849_/X _57850_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_10_412_0_CLK clkbuf_9_206_0_CLK/X _85334_/CLK sky130_fd_sc_hd__clkbuf_1
X_69836_ _73273_/A _69833_/X _69617_/X _69835_/Y _69836_/X sky130_fd_sc_hd__a211o_4
X_50185_ _50113_/A _50185_/X sky130_fd_sc_hd__buf_2
X_85882_ _85879_/CLK _52136_/Y _72957_/B sky130_fd_sc_hd__dfxtp_4
X_56801_ _56800_/X _56801_/X sky130_fd_sc_hd__buf_2
X_87621_ _88394_/CLK _87621_/D _87621_/Q sky130_fd_sc_hd__dfxtp_4
X_84833_ _84714_/CLK _58503_/Y _64307_/C sky130_fd_sc_hd__dfxtp_4
X_57781_ _58631_/A _57781_/X sky130_fd_sc_hd__buf_2
X_69767_ _88068_/Q _69751_/X _69088_/X _69766_/Y _69767_/X sky130_fd_sc_hd__a211o_4
X_54993_ _54990_/Y _54971_/X _54992_/X _54993_/Y sky130_fd_sc_hd__a21oi_4
X_66979_ _88386_/Q _66954_/X _66955_/X _66978_/X _66979_/X sky130_fd_sc_hd__a211o_4
X_59520_ _59520_/A _59536_/A sky130_fd_sc_hd__buf_2
X_56732_ _57023_/A _56732_/X sky130_fd_sc_hd__buf_2
X_68718_ _69906_/A _68718_/B _68718_/X sky130_fd_sc_hd__and2_4
X_87552_ _87814_/CLK _43164_/Y _73252_/A sky130_fd_sc_hd__dfxtp_4
X_53944_ _53944_/A _57491_/B _53944_/C _53944_/Y sky130_fd_sc_hd__nor3_4
X_84764_ _84760_/CLK _59171_/Y _59159_/A sky130_fd_sc_hd__dfxtp_4
X_81976_ _81928_/CLK _81976_/D _77775_/B sky130_fd_sc_hd__dfxtp_4
X_69698_ _64696_/A _69698_/B _69698_/Y sky130_fd_sc_hd__nor2_4
X_86503_ _86499_/CLK _48658_/Y _86503_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_427_0_CLK clkbuf_9_213_0_CLK/X _83238_/CLK sky130_fd_sc_hd__clkbuf_1
X_59451_ _59450_/Y _59444_/X _59451_/Y sky130_fd_sc_hd__nand2_4
X_83715_ _85436_/CLK _70725_/Y _46975_/A sky130_fd_sc_hd__dfxtp_4
X_56663_ _56663_/A _56663_/X sky130_fd_sc_hd__buf_2
X_80927_ _81169_/CLK _80927_/D _80927_/Q sky130_fd_sc_hd__dfxtp_4
X_68649_ _68649_/A _68649_/X sky130_fd_sc_hd__buf_2
X_87483_ _87484_/CLK _87483_/D _87483_/Q sky130_fd_sc_hd__dfxtp_4
X_53875_ _52355_/A _53875_/B _53806_/C _53875_/X sky130_fd_sc_hd__and3_4
X_84695_ _84355_/CLK _84695_/D _80433_/A sky130_fd_sc_hd__dfxtp_4
X_58402_ _84857_/Q _58403_/A sky130_fd_sc_hd__inv_2
X_55614_ _44115_/A _55615_/A sky130_fd_sc_hd__buf_2
X_86434_ _83594_/CLK _86434_/D _86434_/Q sky130_fd_sc_hd__dfxtp_4
X_40840_ _40835_/X _40836_/X _40839_/X _69756_/B _40832_/X _40840_/Y
+ sky130_fd_sc_hd__o32ai_4
X_52826_ _52852_/A _52831_/B sky130_fd_sc_hd__buf_2
X_83646_ _86422_/CLK _83646_/D _83646_/Q sky130_fd_sc_hd__dfxtp_4
X_59382_ _59311_/X _85730_/Q _59334_/X _59382_/X sky130_fd_sc_hd__o21a_4
X_71660_ _71660_/A _71228_/B _71660_/C _71660_/Y sky130_fd_sc_hd__nand3_4
X_56594_ _55504_/Y _56629_/B sky130_fd_sc_hd__buf_2
X_80858_ _80740_/CLK _80890_/Q _75016_/B sky130_fd_sc_hd__dfxtp_4
X_70611_ _70773_/A _70611_/X sky130_fd_sc_hd__buf_2
X_58333_ _56995_/X _58334_/A sky130_fd_sc_hd__buf_2
X_55545_ _57254_/B _55510_/X _55512_/X _55544_/Y _55545_/X sky130_fd_sc_hd__a211o_4
X_86365_ _83716_/CLK _49562_/Y _59044_/B sky130_fd_sc_hd__dfxtp_4
X_40771_ _40770_/Y _40771_/X sky130_fd_sc_hd__buf_2
X_52757_ _52757_/A _52775_/A sky130_fd_sc_hd__buf_2
X_71591_ _71581_/X _83446_/Q _71590_/Y _83446_/D sky130_fd_sc_hd__a21o_4
X_83577_ _86505_/CLK _83577_/D _48538_/A sky130_fd_sc_hd__dfxtp_4
X_80789_ _80813_/CLK _75754_/Y _75358_/A sky130_fd_sc_hd__dfxtp_4
X_42510_ _42486_/X _42501_/X _40696_/X _42509_/Y _42489_/X _42510_/Y
+ sky130_fd_sc_hd__o32ai_4
X_88104_ _88104_/CLK _88104_/D _41922_/A sky130_fd_sc_hd__dfxtp_4
X_73330_ _72870_/X _86187_/Q _72905_/X _73329_/X _73330_/X sky130_fd_sc_hd__a211o_4
X_85316_ _85346_/CLK _55113_/Y _85316_/Q sky130_fd_sc_hd__dfxtp_4
X_51708_ _85960_/Q _51701_/X _51707_/Y _51708_/Y sky130_fd_sc_hd__o21ai_4
X_70542_ _70533_/X _83753_/Q _70541_/Y _70542_/X sky130_fd_sc_hd__a21o_4
X_58264_ _58264_/A _58264_/Y sky130_fd_sc_hd__inv_2
X_82528_ _82529_/CLK _79101_/Y _82528_/Q sky130_fd_sc_hd__dfxtp_4
X_43490_ _43490_/A _87396_/D sky130_fd_sc_hd__inv_2
X_55476_ _55826_/A _55477_/A sky130_fd_sc_hd__buf_2
X_86296_ _86297_/CLK _49939_/Y _72232_/B sky130_fd_sc_hd__dfxtp_4
X_52688_ _52688_/A _52770_/A sky130_fd_sc_hd__buf_2
X_57215_ _56893_/B _56877_/X _56860_/X _57215_/X sky130_fd_sc_hd__a21o_4
X_88035_ _87789_/CLK _42102_/X _88035_/Q sky130_fd_sc_hd__dfxtp_4
X_42441_ _42440_/Y _87863_/D sky130_fd_sc_hd__inv_2
X_54427_ _54399_/A _54435_/A sky130_fd_sc_hd__buf_2
X_73261_ _73210_/X _85582_/Q _73092_/X _73260_/X _73261_/X sky130_fd_sc_hd__a211o_4
X_85247_ _85184_/CLK _56294_/Y _85247_/Q sky130_fd_sc_hd__dfxtp_4
X_51639_ _51639_/A _51639_/X sky130_fd_sc_hd__buf_2
X_70473_ _71323_/A _71500_/C _70472_/X _70473_/Y sky130_fd_sc_hd__nand3_4
X_58195_ _58191_/X _58192_/Y _58194_/Y _58195_/Y sky130_fd_sc_hd__a21oi_4
X_82459_ _83520_/CLK _79151_/X _82427_/D sky130_fd_sc_hd__dfxtp_4
X_75000_ _74986_/X _74994_/X _75000_/X sky130_fd_sc_hd__and2_4
X_72212_ _72208_/Y _72211_/Y _72201_/X _72212_/X sky130_fd_sc_hd__a21o_4
X_45160_ _45152_/X _45157_/Y _45159_/Y _45160_/Y sky130_fd_sc_hd__a21oi_4
X_57146_ _57416_/A _57158_/C _57416_/C _57146_/Y sky130_fd_sc_hd__nand3_4
X_42372_ _42371_/Y _87896_/D sky130_fd_sc_hd__inv_2
X_54358_ _54362_/A _54362_/B _54362_/C _46774_/Y _54358_/X sky130_fd_sc_hd__and4_4
X_73192_ _83161_/Q _73079_/X _73191_/X _73192_/X sky130_fd_sc_hd__a21o_4
X_85178_ _85241_/CLK _56486_/Y _85178_/Q sky130_fd_sc_hd__dfxtp_4
X_44111_ _44110_/X _44111_/X sky130_fd_sc_hd__buf_2
X_53309_ _53298_/A _53309_/B _53309_/Y sky130_fd_sc_hd__nand2_4
X_41323_ _41322_/Y _41323_/Y sky130_fd_sc_hd__inv_2
X_72143_ _57759_/X _72143_/X sky130_fd_sc_hd__buf_2
X_84129_ _85346_/CLK _84129_/D _84129_/Q sky130_fd_sc_hd__dfxtp_4
X_45091_ _56407_/C _45027_/X _45090_/X _45091_/Y sky130_fd_sc_hd__o21ai_4
X_57077_ _56903_/X _57075_/Y _57077_/Y sky130_fd_sc_hd__nand2_4
X_54289_ _85469_/Q _54266_/X _54288_/Y _54289_/Y sky130_fd_sc_hd__o21ai_4
X_44042_ _80665_/Q _55133_/A sky130_fd_sc_hd__inv_2
X_56028_ _55688_/X _56026_/X _56027_/Y _85309_/D sky130_fd_sc_hd__o21ai_4
X_41254_ _41250_/X _41251_/X _68984_/B _41253_/X _88250_/D sky130_fd_sc_hd__a2bb2o_4
X_72074_ _71993_/A _72075_/A sky130_fd_sc_hd__buf_2
X_76951_ _76951_/A _76952_/B sky130_fd_sc_hd__inv_2
X_71025_ _70773_/A _71026_/A sky130_fd_sc_hd__buf_2
X_75902_ _75902_/A _84372_/Q _75902_/X sky130_fd_sc_hd__xor2_4
X_48850_ _48848_/Y _48840_/X _48849_/X _48850_/Y sky130_fd_sc_hd__a21oi_4
X_79670_ _84213_/Q _72357_/A _79670_/X sky130_fd_sc_hd__xor2_4
X_41185_ _40947_/A _41186_/A sky130_fd_sc_hd__buf_2
X_76882_ _76881_/C _81498_/Q _81370_/D _76882_/Y sky130_fd_sc_hd__nand3_4
X_47801_ _47661_/A _50886_/C sky130_fd_sc_hd__buf_2
X_78621_ _78621_/A _78621_/Y sky130_fd_sc_hd__inv_2
X_75833_ _75815_/A _75820_/A _75821_/A _75833_/Y sky130_fd_sc_hd__a21oi_4
X_87819_ _87821_/CLK _87819_/D _87819_/Q sky130_fd_sc_hd__dfxtp_4
X_48781_ _48781_/A _48781_/X sky130_fd_sc_hd__buf_2
X_45993_ _45992_/Y _86824_/D sky130_fd_sc_hd__inv_2
X_57979_ _84935_/Q _57896_/X _57973_/X _57978_/X _84935_/D sky130_fd_sc_hd__a2bb2oi_4
X_47732_ _47728_/Y _47698_/X _47731_/X _86604_/D sky130_fd_sc_hd__a21oi_4
X_59718_ _59696_/A _59711_/B _80568_/A _59718_/Y sky130_fd_sc_hd__nor3_4
X_78552_ _78552_/A _78552_/Y sky130_fd_sc_hd__inv_2
X_44944_ _85278_/Q _44911_/X _44943_/X _44944_/Y sky130_fd_sc_hd__o21ai_4
X_75764_ _75751_/A _75750_/Y _75764_/Y sky130_fd_sc_hd__nor2_4
X_60990_ _60969_/X _60835_/X _84544_/Q _60990_/X sky130_fd_sc_hd__or3_4
X_72976_ _87819_/Q _72894_/X _72976_/Y sky130_fd_sc_hd__nor2_4
X_77503_ _81940_/Q _82196_/D _81908_/D sky130_fd_sc_hd__xor2_4
X_74715_ MACRO_RD_SELECT _74715_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_8_54_0_CLK clkbuf_8_55_0_CLK/A clkbuf_8_54_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_47663_ _47663_/A _53177_/D sky130_fd_sc_hd__buf_2
X_71927_ _56721_/A _71917_/X _71926_/Y _83326_/D sky130_fd_sc_hd__o21ai_4
X_59649_ _59649_/A _59628_/A _59743_/B _59649_/Y sky130_fd_sc_hd__nor3_4
X_78483_ _82510_/Q _82766_/D _78483_/X sky130_fd_sc_hd__xor2_4
X_44875_ _80671_/Q _44875_/X sky130_fd_sc_hd__buf_2
X_75695_ _81120_/Q _75695_/B _75695_/Y sky130_fd_sc_hd__xnor2_4
X_49402_ _49400_/Y _49378_/X _49401_/X _86394_/D sky130_fd_sc_hd__a21oi_4
X_46614_ _46892_/A _46614_/X sky130_fd_sc_hd__buf_2
X_77434_ _77416_/X _77434_/B _77434_/Y sky130_fd_sc_hd__nor2_4
X_43826_ _43826_/A _87249_/D sky130_fd_sc_hd__inv_2
X_62660_ _62886_/A _62660_/X sky130_fd_sc_hd__buf_2
X_74646_ _74638_/X _56607_/A _83002_/Q _74645_/X _83002_/D sky130_fd_sc_hd__a2bb2o_4
X_47594_ _47594_/A _53139_/D sky130_fd_sc_hd__buf_2
X_71858_ _71848_/X _83351_/Q _71857_/Y _83351_/D sky130_fd_sc_hd__a21o_4
X_49333_ _49331_/Y _49326_/X _49332_/Y _49333_/Y sky130_fd_sc_hd__a21boi_4
X_61611_ _61611_/A _61611_/B _61611_/C _61572_/D _61611_/Y sky130_fd_sc_hd__nand4_4
X_46545_ _46545_/A _54069_/B sky130_fd_sc_hd__inv_2
X_70809_ _70809_/A _70942_/B sky130_fd_sc_hd__buf_2
X_77365_ _81931_/Q _82187_/D _81899_/D sky130_fd_sc_hd__xor2_4
X_43757_ _43005_/X _43563_/X _40950_/X _69165_/B _43756_/X _43757_/Y
+ sky130_fd_sc_hd__o32ai_4
X_62591_ _61649_/B _62548_/C _62507_/X _62548_/B _62590_/X _62591_/X
+ sky130_fd_sc_hd__a41o_4
X_74577_ _45095_/A _74568_/X _74576_/X _83029_/D sky130_fd_sc_hd__o21ai_4
X_40969_ _40968_/X _40941_/X _69224_/B _40942_/X _40969_/X sky130_fd_sc_hd__a2bb2o_4
X_71789_ _58186_/Y _71784_/X _71788_/Y _83376_/D sky130_fd_sc_hd__o21ai_4
X_79104_ _79109_/A _79109_/B _79104_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_69_0_CLK clkbuf_8_69_0_CLK/A clkbuf_8_69_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_64330_ _79784_/B _64314_/X _64329_/X _84256_/D sky130_fd_sc_hd__a21o_4
X_76316_ _76316_/A _76315_/X _76317_/B sky130_fd_sc_hd__xor2_4
X_42708_ _42687_/X _42688_/X _41139_/X _87758_/Q _42700_/X _42709_/A
+ sky130_fd_sc_hd__o32ai_4
X_61542_ _61542_/A _61542_/B _61542_/C _61512_/X _61542_/Y sky130_fd_sc_hd__nand4_4
X_49264_ _49262_/Y _49247_/X _49263_/Y _49264_/Y sky130_fd_sc_hd__a21boi_4
X_73528_ _42063_/Y _72974_/X _73393_/X _73527_/Y _73528_/X sky130_fd_sc_hd__a211o_4
X_46476_ _46476_/A _52522_/B sky130_fd_sc_hd__inv_2
X_77296_ _77296_/A _77312_/A _77294_/Y _77296_/Y sky130_fd_sc_hd__nand3_4
X_43688_ _40798_/X _43685_/X _72924_/A _43686_/X _87309_/D sky130_fd_sc_hd__a2bb2o_4
X_48215_ _48190_/A _50268_/B _48215_/Y sky130_fd_sc_hd__nand2_4
X_79035_ _82747_/Q _79035_/B _79035_/X sky130_fd_sc_hd__xor2_4
X_45427_ _45425_/Y _45412_/X _45396_/X _45426_/Y _45427_/X sky130_fd_sc_hd__a211o_4
X_64261_ _64275_/A _63049_/B _64223_/C _64261_/X sky130_fd_sc_hd__and3_4
X_76247_ _76251_/C _76247_/Y sky130_fd_sc_hd__inv_2
X_42639_ _42639_/A _42639_/Y sky130_fd_sc_hd__inv_2
X_49195_ _49195_/A _53936_/B sky130_fd_sc_hd__inv_2
X_61473_ _61460_/Y _61463_/Y _61464_/X _61468_/Y _61472_/Y _61473_/X
+ sky130_fd_sc_hd__a41o_4
X_73459_ _73445_/Y _73458_/X _73460_/B sky130_fd_sc_hd__xnor2_4
X_66000_ _65523_/X _66062_/B _65526_/X _66000_/Y sky130_fd_sc_hd__nand3_4
X_63212_ _58383_/A _63190_/X _63175_/X _58259_/A _63176_/X _63212_/Y
+ sky130_fd_sc_hd__o32ai_4
X_48146_ _48146_/A _48136_/B _48146_/X sky130_fd_sc_hd__or2_4
X_60424_ _60376_/X _60399_/Y _60414_/Y _60532_/A _60423_/X _60424_/X
+ sky130_fd_sc_hd__o41a_4
X_45358_ _55715_/B _45357_/X _45339_/X _45358_/X sky130_fd_sc_hd__o21a_4
X_64192_ _62629_/A _64192_/B _64192_/C _64192_/D _64193_/D sky130_fd_sc_hd__nand4_4
X_76178_ _76161_/Y _76159_/Y _76178_/Y sky130_fd_sc_hd__nand2_4
X_44309_ _44308_/X _57470_/B sky130_fd_sc_hd__buf_2
X_75129_ _75129_/A _75129_/Y sky130_fd_sc_hd__inv_2
X_63143_ _63097_/A _64353_/B _63108_/C _63121_/D _63143_/X sky130_fd_sc_hd__and4_4
X_48077_ _48077_/A _48086_/B _48077_/X sky130_fd_sc_hd__or2_4
X_60355_ _59552_/C _60407_/C _60132_/A _60355_/Y sky130_fd_sc_hd__nand3_4
X_45289_ _56145_/C _45269_/X _45229_/X _45289_/X sky130_fd_sc_hd__o21a_4
X_47028_ _54503_/D _52811_/D sky130_fd_sc_hd__buf_2
X_63074_ _58424_/Y _63073_/X _63059_/X _59471_/A _63060_/X _63074_/Y
+ sky130_fd_sc_hd__o32ai_4
X_67951_ _67972_/A _87705_/Q _67951_/X sky130_fd_sc_hd__and2_4
X_79937_ _79937_/A _79937_/B _79937_/Y sky130_fd_sc_hd__nand2_4
X_60286_ _60273_/X _60259_/A _60285_/Y _60286_/X sky130_fd_sc_hd__a21o_4
X_66902_ _68614_/A _66902_/X sky130_fd_sc_hd__buf_2
X_62025_ _61560_/B _62007_/X _61967_/C _62008_/X _62025_/Y sky130_fd_sc_hd__nand4_4
X_79868_ _79875_/B _79868_/B _79868_/X sky130_fd_sc_hd__xor2_4
X_67882_ _67955_/A _86920_/Q _67882_/X sky130_fd_sc_hd__and2_4
X_69621_ _57803_/A _69908_/A sky130_fd_sc_hd__buf_2
X_66833_ _69457_/A _66833_/X sky130_fd_sc_hd__buf_2
X_78819_ _78817_/Y _78818_/Y _78820_/B sky130_fd_sc_hd__nand2_4
X_48979_ _48979_/A _48940_/B _48928_/C _48979_/X sky130_fd_sc_hd__and3_4
X_79799_ _79795_/X _79798_/Y _79799_/X sky130_fd_sc_hd__xor2_4
X_69552_ _83915_/Q _69504_/X _69551_/X _69552_/X sky130_fd_sc_hd__a21bo_4
X_81830_ _82211_/CLK _81862_/Q _77279_/A sky130_fd_sc_hd__dfxtp_4
X_66764_ _66879_/A _66764_/X sky130_fd_sc_hd__buf_2
X_51990_ _51961_/X _48236_/B _51990_/Y sky130_fd_sc_hd__nand2_4
X_63976_ _63960_/A _63960_/B _80102_/B _63976_/Y sky130_fd_sc_hd__nor3_4
X_68503_ _88014_/Q _68402_/X _68501_/X _68502_/X _68503_/X sky130_fd_sc_hd__a211o_4
X_65715_ _65777_/A _85870_/Q _65715_/X sky130_fd_sc_hd__and2_4
X_50941_ _50941_/A _50941_/B _50948_/C _46716_/X _50941_/X sky130_fd_sc_hd__and4_4
X_62927_ _62927_/A _62926_/B _84785_/Q _62928_/D sky130_fd_sc_hd__nand3_4
X_81761_ _81412_/CLK _76150_/X _41286_/A sky130_fd_sc_hd__dfxtp_4
X_69483_ _87514_/Q _69356_/X _69371_/X _69482_/X _69483_/X sky130_fd_sc_hd__a211o_4
X_66695_ _87130_/Q _66593_/X _66594_/X _66694_/X _66695_/X sky130_fd_sc_hd__a211o_4
X_83500_ _84223_/CLK _83500_/D _83500_/Q sky130_fd_sc_hd__dfxtp_4
X_80712_ _80681_/CLK _75898_/X _80680_/D sky130_fd_sc_hd__dfxtp_4
X_68434_ _68376_/X _66524_/B _68424_/Y _68433_/Y _68434_/X sky130_fd_sc_hd__a211o_4
X_53660_ _53687_/A _53660_/X sky130_fd_sc_hd__buf_2
X_65646_ _65646_/A _65645_/X _65646_/Y sky130_fd_sc_hd__nand2_4
X_84480_ _84481_/CLK _61446_/Y _79148_/B sky130_fd_sc_hd__dfxtp_4
X_50872_ _50228_/X _52565_/B _50872_/Y sky130_fd_sc_hd__nand2_4
X_62858_ _62646_/B _62858_/X sky130_fd_sc_hd__buf_2
X_81692_ _81695_/CLK _80202_/X _81692_/Q sky130_fd_sc_hd__dfxtp_4
X_52611_ _52609_/Y _52592_/X _52610_/X _52611_/Y sky130_fd_sc_hd__a21oi_4
X_83431_ _83431_/CLK _71636_/Y _59484_/A sky130_fd_sc_hd__dfxtp_4
X_61809_ _61387_/X _61794_/B _61809_/C _61776_/D _61809_/Y sky130_fd_sc_hd__nand4_4
X_80643_ _80643_/A _74715_/Y DATA_FROM_HASH[0] sky130_fd_sc_hd__ebufn_2
X_68365_ _68757_/A _68365_/X sky130_fd_sc_hd__buf_2
X_65577_ _64903_/A _65731_/A sky130_fd_sc_hd__buf_2
X_53591_ _53604_/A _50368_/B _53591_/Y sky130_fd_sc_hd__nand2_4
X_62789_ _62789_/A _63139_/A _62744_/X _62789_/D _62789_/X sky130_fd_sc_hd__and4_4
X_55330_ _55328_/C _55384_/A _55316_/X _55330_/X sky130_fd_sc_hd__a21bo_4
X_67316_ _67316_/A _67315_/X _67316_/Y sky130_fd_sc_hd__nand2_4
X_86150_ _85542_/CLK _50705_/Y _86150_/Q sky130_fd_sc_hd__dfxtp_4
X_52542_ _52319_/A _52542_/X sky130_fd_sc_hd__buf_2
X_64528_ _64523_/X _64524_/X _64525_/X _64527_/Y _64521_/X _64528_/X
+ sky130_fd_sc_hd__o41a_4
X_83362_ _83362_/CLK _71822_/X _83362_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_207 sky130_fd_sc_hd__decap_3
X_80574_ _80554_/Y _80571_/X _80573_/X _80574_/Y sky130_fd_sc_hd__a21boi_4
X_68296_ _67824_/X _67827_/X _68295_/X _68296_/Y sky130_fd_sc_hd__a21oi_4
XPHY_218 sky130_fd_sc_hd__decap_3
X_85101_ _85037_/CLK _85101_/D _85101_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_229 sky130_fd_sc_hd__decap_3
X_82313_ _82335_/CLK _77049_/B _82313_/Q sky130_fd_sc_hd__dfxtp_4
X_55261_ _55252_/A _85129_/Q _55261_/X sky130_fd_sc_hd__and2_4
X_67247_ _67247_/A _67246_/X _67247_/Y sky130_fd_sc_hd__nand2_4
X_86081_ _85761_/CLK _51062_/Y _86081_/Q sky130_fd_sc_hd__dfxtp_4
X_52473_ _85815_/Q _52470_/X _52472_/Y _52473_/Y sky130_fd_sc_hd__o21ai_4
X_64459_ _58393_/Y _61082_/X _61179_/A _64203_/B _64459_/Y sky130_fd_sc_hd__nor4_4
X_83293_ _83304_/CLK _83293_/D _83293_/Q sky130_fd_sc_hd__dfxtp_4
X_57000_ _56966_/X _57153_/A _56999_/Y _57001_/A sky130_fd_sc_hd__o21ai_4
X_54212_ _85483_/Q _54193_/X _54211_/Y _54212_/Y sky130_fd_sc_hd__o21ai_4
X_85032_ _83335_/CLK _57344_/Y _57340_/B sky130_fd_sc_hd__dfxtp_4
X_51424_ _51403_/X _52950_/B _51424_/Y sky130_fd_sc_hd__nand2_4
X_82244_ _82263_/CLK _82244_/D _82244_/Q sky130_fd_sc_hd__dfxtp_4
X_67178_ _87866_/Q _67176_/X _67153_/X _67177_/X _67178_/X sky130_fd_sc_hd__a211o_4
X_55192_ _55192_/A _85133_/Q _55192_/X sky130_fd_sc_hd__and2_4
X_54143_ _85496_/Q _54140_/X _54142_/Y _54143_/Y sky130_fd_sc_hd__o21ai_4
X_66129_ _66054_/X _73927_/B _66129_/X sky130_fd_sc_hd__and2_4
X_51355_ _86026_/Q _51332_/X _51354_/Y _51355_/Y sky130_fd_sc_hd__o21ai_4
X_82175_ _82575_/CLK _84167_/Q _78006_/B sky130_fd_sc_hd__dfxtp_4
X_50306_ _50240_/A _50306_/B _50306_/Y sky130_fd_sc_hd__nand2_4
X_81126_ _80835_/CLK _81126_/D _40737_/A sky130_fd_sc_hd__dfxtp_4
X_58951_ _58948_/Y _58950_/Y _58939_/X _58951_/X sky130_fd_sc_hd__a21o_4
X_54074_ _85510_/Q _54067_/X _54073_/Y _54074_/Y sky130_fd_sc_hd__o21ai_4
X_51286_ _51286_/A _51296_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_351_0_CLK clkbuf_9_175_0_CLK/X _85748_/CLK sky130_fd_sc_hd__clkbuf_1
X_86983_ _86998_/CLK _44730_/Y _74119_/A sky130_fd_sc_hd__dfxtp_4
X_57902_ _58876_/A _58605_/A sky130_fd_sc_hd__buf_2
X_53025_ _53025_/A _53025_/B _53025_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_981_0_CLK clkbuf_9_490_0_CLK/X _85555_/CLK sky130_fd_sc_hd__clkbuf_1
X_50237_ _50505_/A _50464_/A sky130_fd_sc_hd__buf_2
X_85934_ _86096_/CLK _51856_/Y _85934_/Q sky130_fd_sc_hd__dfxtp_4
X_81057_ _85335_/CLK _81057_/D _81057_/Q sky130_fd_sc_hd__dfxtp_4
X_58882_ _58882_/A _59053_/A sky130_fd_sc_hd__buf_2
X_80008_ _80004_/X _80007_/Y _80008_/X sky130_fd_sc_hd__xor2_4
X_57833_ _86650_/Q _57833_/B _57833_/Y sky130_fd_sc_hd__nor2_4
X_69819_ _81967_/D _69763_/X _69818_/X _83895_/D sky130_fd_sc_hd__a21bo_4
Xclkbuf_9_472_0_CLK clkbuf_8_236_0_CLK/X clkbuf_9_472_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_50168_ _50165_/Y _50166_/X _50167_/X _86251_/D sky130_fd_sc_hd__a21oi_4
X_85865_ _85865_/CLK _85865_/D _85865_/Q sky130_fd_sc_hd__dfxtp_4
X_87604_ _87348_/CLK _87604_/D _87604_/Q sky130_fd_sc_hd__dfxtp_4
X_72830_ _72829_/X _72830_/X sky130_fd_sc_hd__buf_2
X_84816_ _84815_/CLK _58584_/Y _84816_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_366_0_CLK clkbuf_9_183_0_CLK/X _85990_/CLK sky130_fd_sc_hd__clkbuf_1
X_57764_ _57761_/X _85501_/Q _57763_/X _57764_/X sky130_fd_sc_hd__o21a_4
X_42990_ _40485_/X _42962_/X _87616_/Q _42963_/X _87616_/D sky130_fd_sc_hd__a2bb2o_4
X_50099_ _50103_/A _52307_/B _50099_/Y sky130_fd_sc_hd__nand2_4
X_54976_ _54985_/A _47552_/A _54976_/Y sky130_fd_sc_hd__nand2_4
X_85796_ _85507_/CLK _85796_/D _65360_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_996_0_CLK clkbuf_9_498_0_CLK/X _85596_/CLK sky130_fd_sc_hd__clkbuf_1
X_59503_ _46159_/X _59500_/Y _59502_/Y _59503_/Y sky130_fd_sc_hd__a21oi_4
X_56715_ _57270_/A _56713_/X _56714_/Y _56715_/Y sky130_fd_sc_hd__o21ai_4
X_87535_ _87544_/CLK _87535_/D _87535_/Q sky130_fd_sc_hd__dfxtp_4
X_41941_ _41941_/A _41941_/Y sky130_fd_sc_hd__inv_2
X_53927_ _53951_/A _49176_/A _53927_/Y sky130_fd_sc_hd__nand2_4
X_72761_ _72754_/X _72761_/B _72762_/B sky130_fd_sc_hd__nand2_4
X_84747_ _84760_/CLK _84747_/D _84747_/Q sky130_fd_sc_hd__dfxtp_4
X_57695_ _57694_/X _58805_/A sky130_fd_sc_hd__buf_2
X_81959_ _82339_/CLK _81959_/D _77919_/B sky130_fd_sc_hd__dfxtp_4
X_74500_ _83053_/Q _46250_/X _74499_/Y _74500_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_487_0_CLK clkbuf_9_486_0_CLK/A clkbuf_9_487_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_71712_ _71711_/Y _71712_/Y sky130_fd_sc_hd__inv_2
X_59434_ _59433_/Y _59424_/B _59434_/Y sky130_fd_sc_hd__nand2_4
X_44660_ _44714_/A _44660_/X sky130_fd_sc_hd__buf_2
X_56646_ _45957_/A _56645_/Y _56646_/Y sky130_fd_sc_hd__nor2_4
X_75480_ _75479_/X _75480_/Y sky130_fd_sc_hd__inv_2
X_87466_ _87708_/CLK _87466_/D _87466_/Q sky130_fd_sc_hd__dfxtp_4
X_41872_ _41872_/A _41872_/X sky130_fd_sc_hd__buf_2
X_53858_ _53844_/A _53858_/B _53858_/Y sky130_fd_sc_hd__nand2_4
X_72692_ _83188_/Q _72686_/X _72691_/Y _72692_/X sky130_fd_sc_hd__a21bo_4
X_84678_ _84396_/CLK _84678_/D _80215_/A sky130_fd_sc_hd__dfxtp_4
X_43611_ _43611_/A _43611_/X sky130_fd_sc_hd__buf_2
X_74431_ _74431_/A _74420_/X _74425_/X _74431_/X sky130_fd_sc_hd__and3_4
X_86417_ _86422_/CLK _49290_/Y _65029_/B sky130_fd_sc_hd__dfxtp_4
X_52809_ _52783_/A _52809_/X sky130_fd_sc_hd__buf_2
X_40823_ _40820_/X _40821_/X _88328_/Q _40822_/X _40823_/X sky130_fd_sc_hd__a2bb2o_4
X_59365_ _59081_/A _59365_/X sky130_fd_sc_hd__buf_2
X_71643_ _59497_/Y _71628_/X _71642_/Y _71643_/Y sky130_fd_sc_hd__o21ai_4
X_83629_ _83630_/CLK _71034_/Y _83629_/Q sky130_fd_sc_hd__dfxtp_4
X_44591_ _44588_/X _44589_/X _40914_/X _87043_/Q _44590_/X _44591_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56577_ _72641_/C _56558_/X _56577_/Y sky130_fd_sc_hd__xnor2_4
X_87397_ _87397_/CLK _43488_/Y _87397_/Q sky130_fd_sc_hd__dfxtp_4
X_53789_ _48894_/A _53806_/B _53774_/C _53789_/X sky130_fd_sc_hd__and3_4
X_46330_ _46330_/A _52454_/B sky130_fd_sc_hd__buf_2
X_58316_ _84880_/Q _58317_/A sky130_fd_sc_hd__inv_2
X_77150_ _77146_/B _77154_/A _77149_/Y _77151_/B sky130_fd_sc_hd__a21boi_4
X_43542_ _40363_/X _43542_/X sky130_fd_sc_hd__buf_2
X_55528_ _55477_/A _55534_/A sky130_fd_sc_hd__buf_2
X_86348_ _86351_/CLK _86348_/D _59256_/B sky130_fd_sc_hd__dfxtp_4
X_74362_ _83082_/Q _72699_/X _74361_/Y _74362_/X sky130_fd_sc_hd__a21bo_4
X_40754_ _40793_/A _40754_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_410_0_CLK clkbuf_9_411_0_CLK/A clkbuf_9_410_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_59296_ _59208_/X _86057_/Q _59295_/X _59296_/Y sky130_fd_sc_hd__o21ai_4
X_71574_ _71865_/A _71583_/B _71574_/C _71574_/Y sky130_fd_sc_hd__nor3_4
X_76101_ _81723_/D _76109_/B _76103_/A sky130_fd_sc_hd__xor2_4
X_73313_ _48593_/A _73313_/B _73313_/X sky130_fd_sc_hd__xor2_4
X_46261_ _48631_/A _46348_/A sky130_fd_sc_hd__buf_2
X_70525_ _57678_/Y _70500_/Y _70524_/Y _83755_/D sky130_fd_sc_hd__o21ai_4
X_58247_ _84898_/Q _58248_/A sky130_fd_sc_hd__buf_2
X_77081_ _82093_/Q _77081_/B _77081_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_10_304_0_CLK clkbuf_9_152_0_CLK/X _83495_/CLK sky130_fd_sc_hd__clkbuf_1
X_43473_ _43472_/X _43452_/X _41667_/X _87404_/Q _43456_/X _43474_/A
+ sky130_fd_sc_hd__o32ai_4
X_55459_ _55454_/X _45599_/Y _55459_/Y sky130_fd_sc_hd__nor2_4
X_74293_ _74297_/A _74297_/B _55966_/X _74293_/Y sky130_fd_sc_hd__nand3_4
X_86279_ _85959_/CLK _50026_/Y _72427_/B sky130_fd_sc_hd__dfxtp_4
X_40685_ _40685_/A _88354_/D sky130_fd_sc_hd__inv_2
X_48000_ _48755_/A _48731_/A sky130_fd_sc_hd__buf_2
X_45212_ _45212_/A _45212_/X sky130_fd_sc_hd__buf_2
X_76032_ _76032_/A _81745_/D _76032_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_10_934_0_CLK clkbuf_9_467_0_CLK/X _88086_/CLK sky130_fd_sc_hd__clkbuf_1
X_88018_ _87260_/CLK _88018_/D _88018_/Q sky130_fd_sc_hd__dfxtp_4
X_42424_ _42424_/A _87871_/D sky130_fd_sc_hd__inv_2
X_73244_ _73242_/X _73230_/X _73232_/Y _73244_/Y sky130_fd_sc_hd__nand3_4
X_70456_ _70694_/A HASH_ADDR[4] _70412_/X _71462_/B sky130_fd_sc_hd__nor3_4
X_46192_ _46164_/A _46092_/X _46217_/C sky130_fd_sc_hd__nor2_4
X_58178_ _58177_/Y _64292_/A sky130_fd_sc_hd__buf_2
X_45143_ _64392_/B _61509_/B sky130_fd_sc_hd__buf_2
X_57129_ _57129_/A _57129_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_9_425_0_CLK clkbuf_9_424_0_CLK/A clkbuf_9_425_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_42355_ _41727_/X _42342_/X _87905_/Q _42343_/X _87905_/D sky130_fd_sc_hd__a2bb2o_4
X_73175_ _73175_/A _44127_/X _73175_/Y sky130_fd_sc_hd__nor2_4
X_70387_ _70387_/A _70997_/A sky130_fd_sc_hd__buf_2
X_41306_ _41305_/Y _41306_/X sky130_fd_sc_hd__buf_2
X_60140_ _60078_/X _60063_/Y _60045_/Y _60138_/Y _60139_/Y _60140_/Y
+ sky130_fd_sc_hd__a41oi_4
X_72126_ _72122_/Y _72125_/Y _59351_/X _72126_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_10_319_0_CLK clkbuf_9_159_0_CLK/X _85379_/CLK sky130_fd_sc_hd__clkbuf_1
X_49951_ _49924_/A _49951_/X sky130_fd_sc_hd__buf_2
X_45074_ _56317_/C _45056_/X _45012_/X _45074_/X sky130_fd_sc_hd__o21a_4
X_42286_ _42279_/X _42275_/X _41545_/X _87939_/Q _42276_/X _42287_/A
+ sky130_fd_sc_hd__o32ai_4
X_77983_ _77983_/A _77983_/B _77983_/C _77983_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_949_0_CLK clkbuf_9_474_0_CLK/X _86218_/CLK sky130_fd_sc_hd__clkbuf_1
X_48902_ _64658_/B _48896_/X _48901_/Y _48902_/Y sky130_fd_sc_hd__o21ai_4
X_44025_ _44025_/A _44025_/X sky130_fd_sc_hd__buf_2
X_79722_ _79722_/A _79722_/B _79722_/X sky130_fd_sc_hd__xor2_4
X_41237_ _41205_/X _41206_/X _41234_/X _88252_/Q _41236_/X _41237_/Y
+ sky130_fd_sc_hd__o32ai_4
X_76934_ _76934_/A _76934_/Y sky130_fd_sc_hd__inv_2
X_60071_ _60011_/X _59995_/X _61277_/C _60070_/Y _60071_/X sky130_fd_sc_hd__a211o_4
X_72057_ _72040_/A _49083_/A _72057_/Y sky130_fd_sc_hd__nand2_4
X_49882_ _49901_/A _53095_/B _49882_/Y sky130_fd_sc_hd__nand2_4
X_71008_ _71055_/A _71066_/B _71001_/C _71008_/Y sky130_fd_sc_hd__nand3_4
X_48833_ _48833_/A _48849_/B sky130_fd_sc_hd__buf_2
X_79653_ _79645_/B _79639_/X _79652_/X _79653_/Y sky130_fd_sc_hd__a21boi_4
X_41168_ _41143_/X _40648_/A _41167_/X _41168_/Y sky130_fd_sc_hd__o21ai_4
X_76865_ _81498_/Q _81370_/D _76910_/A sky130_fd_sc_hd__xor2_4
X_78604_ _78591_/A _78602_/Y _78603_/Y _78604_/X sky130_fd_sc_hd__a21bo_4
X_63830_ _64184_/A _63831_/A sky130_fd_sc_hd__buf_2
X_75816_ _80925_/Q _75818_/A sky130_fd_sc_hd__inv_2
X_48764_ _73042_/B _48754_/X _48763_/Y _48764_/Y sky130_fd_sc_hd__o21ai_4
X_79584_ _79584_/A _79586_/A sky130_fd_sc_hd__buf_2
X_45976_ _45975_/X _45976_/X sky130_fd_sc_hd__buf_2
X_41099_ _41098_/X _41065_/X _69536_/B _41066_/X _88278_/D sky130_fd_sc_hd__a2bb2o_4
X_76796_ _76785_/Y _81361_/D sky130_fd_sc_hd__inv_2
X_47715_ _47620_/X _47715_/X sky130_fd_sc_hd__buf_2
X_78535_ _78547_/A _82674_/D _78536_/B sky130_fd_sc_hd__xor2_4
X_44927_ _85247_/Q _44874_/X _44926_/X _44927_/X sky130_fd_sc_hd__o21a_4
X_63761_ _63761_/A _63761_/X sky130_fd_sc_hd__buf_2
X_75747_ _75747_/A _75747_/B _75748_/B sky130_fd_sc_hd__xor2_4
X_48695_ _48695_/A _48695_/B _48695_/Y sky130_fd_sc_hd__nand2_4
X_60973_ _60901_/B _61012_/C sky130_fd_sc_hd__buf_2
X_72959_ _73257_/A _72959_/X sky130_fd_sc_hd__buf_2
X_65500_ _64757_/X _65548_/B _64760_/X _65512_/A sky130_fd_sc_hd__nand3_4
X_62712_ _58237_/X _62689_/X _62708_/X _62699_/X _62711_/X _62712_/Y
+ sky130_fd_sc_hd__a41oi_4
X_47646_ _47642_/Y _47602_/X _47645_/X _86613_/D sky130_fd_sc_hd__a21oi_4
X_66480_ _66477_/Y _66449_/X _66479_/Y _66480_/X sky130_fd_sc_hd__a21o_4
X_78466_ _78466_/A _78466_/B _78466_/X sky130_fd_sc_hd__or2_4
X_44858_ _43896_/X _44858_/X sky130_fd_sc_hd__buf_2
X_63692_ _63701_/A _63701_/B _80310_/B _63692_/Y sky130_fd_sc_hd__nor3_4
X_75678_ _75678_/A _75677_/Y _75685_/A sky130_fd_sc_hd__xor2_4
X_65431_ _65427_/X _65431_/B _65431_/Y sky130_fd_sc_hd__nand2_4
X_77417_ _77417_/A _77417_/B _77417_/X sky130_fd_sc_hd__xor2_4
X_43809_ _40554_/X _43810_/A sky130_fd_sc_hd__buf_2
X_74629_ _74675_/A _74694_/A sky130_fd_sc_hd__buf_2
X_62643_ _60239_/B _62924_/C sky130_fd_sc_hd__buf_2
X_47577_ _81244_/Q _47578_/A sky130_fd_sc_hd__inv_2
X_78397_ _78369_/A _78397_/B _78397_/Y sky130_fd_sc_hd__nand2_4
X_44789_ _44650_/A _44789_/X sky130_fd_sc_hd__buf_2
X_49316_ _49405_/A _49316_/X sky130_fd_sc_hd__buf_2
X_68150_ _68144_/X _66934_/Y _68148_/X _68149_/Y _68150_/X sky130_fd_sc_hd__a211o_4
X_46528_ _46528_/A _46527_/X _46528_/X sky130_fd_sc_hd__or2_4
X_65362_ _65859_/A _65362_/X sky130_fd_sc_hd__buf_2
X_77348_ _77316_/B _77334_/A _77333_/A _77348_/X sky130_fd_sc_hd__o21a_4
X_62574_ _62551_/X _62553_/X _84400_/Q _62574_/Y sky130_fd_sc_hd__nor3_4
X_67101_ _87113_/Q _67074_/X _67075_/X _67100_/X _67101_/X sky130_fd_sc_hd__a211o_4
X_64313_ _79797_/B _64255_/X _64312_/X _64313_/X sky130_fd_sc_hd__a21o_4
X_49247_ _49247_/A _49247_/X sky130_fd_sc_hd__buf_2
X_61525_ _61334_/A _61525_/X sky130_fd_sc_hd__buf_2
X_68081_ _87380_/Q _67987_/X _68053_/X _68080_/X _68081_/X sky130_fd_sc_hd__a211o_4
X_65293_ _64789_/A _65294_/B sky130_fd_sc_hd__buf_2
X_46459_ _46459_/A _46459_/B _46459_/X sky130_fd_sc_hd__or2_4
X_77279_ _77279_/A _82086_/D _77279_/Y sky130_fd_sc_hd__nand2_4
X_67032_ _66794_/A _67032_/X sky130_fd_sc_hd__buf_2
X_79018_ _79018_/A _79017_/Y _79019_/B sky130_fd_sc_hd__xnor2_4
X_64244_ _64303_/A _64273_/B sky130_fd_sc_hd__buf_2
X_49178_ _65357_/B _49153_/X _49177_/Y _49178_/Y sky130_fd_sc_hd__o21ai_4
X_61456_ _61434_/A _61434_/B _84479_/Q _61456_/Y sky130_fd_sc_hd__nor3_4
X_80290_ _59354_/Y _66332_/C _80292_/A sky130_fd_sc_hd__nand2_4
Xclkbuf_5_19_0_CLK clkbuf_4_9_1_CLK/X clkbuf_6_39_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_48129_ _48125_/Y _48109_/X _48128_/X _86565_/D sky130_fd_sc_hd__a21oi_4
X_60407_ _60407_/A _61293_/B _60407_/C _60408_/C sky130_fd_sc_hd__and3_4
X_64175_ _64187_/A _64187_/B _79921_/A _64175_/Y sky130_fd_sc_hd__nor3_4
X_61387_ _84852_/Q _61387_/X sky130_fd_sc_hd__buf_2
X_51140_ _86066_/Q _51128_/X _51139_/Y _51140_/Y sky130_fd_sc_hd__o21ai_4
X_63126_ _63119_/Y _63121_/X _63122_/X _63124_/X _63125_/X _63126_/Y
+ sky130_fd_sc_hd__o41ai_4
X_60338_ _79671_/A _60323_/X _60334_/Y _60337_/Y _60338_/X sky130_fd_sc_hd__o22a_4
X_68983_ _69223_/A _69027_/A sky130_fd_sc_hd__buf_2
X_51071_ _51056_/A _51071_/B _51071_/C _52763_/D _51071_/X sky130_fd_sc_hd__and4_4
X_67934_ _67934_/A _67933_/X _67934_/Y sky130_fd_sc_hd__nand2_4
X_63057_ _63052_/Y _63054_/X _63056_/X _63057_/Y sky130_fd_sc_hd__a21oi_4
X_60269_ _60268_/Y _60259_/A _79817_/A _59868_/X _84643_/D sky130_fd_sc_hd__a2bb2o_4
X_83980_ _82629_/CLK _83980_/D _82628_/D sky130_fd_sc_hd__dfxtp_4
X_50022_ _50019_/Y _50003_/X _50021_/X _86280_/D sky130_fd_sc_hd__a21oi_4
X_62008_ _61856_/A _62008_/X sky130_fd_sc_hd__buf_2
X_82931_ _82931_/CLK _78257_/X _82931_/Q sky130_fd_sc_hd__dfxtp_4
X_67865_ _68651_/A _67865_/X sky130_fd_sc_hd__buf_2
X_69604_ _69733_/A _69604_/X sky130_fd_sc_hd__buf_2
X_54830_ _54882_/A _54830_/X sky130_fd_sc_hd__buf_2
X_66816_ _69582_/A _66816_/X sky130_fd_sc_hd__buf_2
X_85650_ _85651_/CLK _85650_/D _85650_/Q sky130_fd_sc_hd__dfxtp_4
X_82862_ _82859_/CLK _82862_/D _40864_/A sky130_fd_sc_hd__dfxtp_4
X_67796_ _67891_/A _87200_/Q _67796_/X sky130_fd_sc_hd__and2_4
X_84601_ _84333_/CLK _84601_/D _79141_/A sky130_fd_sc_hd__dfxtp_4
X_81813_ _81259_/CLK _81813_/D _81813_/Q sky130_fd_sc_hd__dfxtp_4
X_69535_ _69532_/X _69534_/X _69346_/X _69535_/X sky130_fd_sc_hd__a21o_4
X_54761_ _54775_/A _54755_/B _54775_/C _47474_/A _54761_/X sky130_fd_sc_hd__and4_4
X_66747_ _66628_/X _66747_/X sky130_fd_sc_hd__buf_2
X_85581_ _85581_/CLK _53721_/Y _85581_/Q sky130_fd_sc_hd__dfxtp_4
X_51973_ _50270_/A _51972_/X _51958_/C _51973_/X sky130_fd_sc_hd__and3_4
X_63959_ _63954_/X _63890_/X _63956_/Y _63957_/Y _63958_/X _63959_/X
+ sky130_fd_sc_hd__a41o_4
X_82793_ _82792_/CLK _82825_/Q _78405_/A sky130_fd_sc_hd__dfxtp_4
X_56500_ _56525_/A _56510_/A sky130_fd_sc_hd__buf_2
X_87320_ _87577_/CLK _87320_/D _74186_/A sky130_fd_sc_hd__dfxtp_4
X_53712_ _53710_/Y _53680_/X _53711_/X _53712_/Y sky130_fd_sc_hd__a21oi_4
X_84532_ _84538_/CLK _84532_/D _76980_/A sky130_fd_sc_hd__dfxtp_4
X_50924_ _50941_/A _50919_/B _50948_/C _51787_/D _50924_/X sky130_fd_sc_hd__and4_4
X_57480_ _57484_/A _56903_/X _57479_/X _57481_/A sky130_fd_sc_hd__o21ai_4
X_81744_ _88175_/CLK _81744_/D _41374_/A sky130_fd_sc_hd__dfxtp_4
X_69466_ _69302_/A _69466_/B _69466_/X sky130_fd_sc_hd__and2_4
X_54692_ _85395_/Q _54676_/X _54691_/Y _54692_/Y sky130_fd_sc_hd__o21ai_4
X_66678_ _69162_/A _66678_/X sky130_fd_sc_hd__buf_2
X_56431_ _56431_/A _56433_/B _85196_/Q _56431_/Y sky130_fd_sc_hd__nand3_4
X_68417_ _73595_/A _68414_/X _68379_/X _68416_/Y _68417_/X sky130_fd_sc_hd__a211o_4
X_87251_ _87776_/CLK _43821_/Y _87251_/Q sky130_fd_sc_hd__dfxtp_4
X_53643_ _53611_/X _74389_/B _53643_/Y sky130_fd_sc_hd__nand2_4
X_65629_ _65769_/A _86516_/Q _65629_/X sky130_fd_sc_hd__and2_4
X_84463_ _82452_/CLK _61647_/Y _79131_/B sky130_fd_sc_hd__dfxtp_4
X_50855_ _50853_/Y _50849_/X _50854_/Y _86120_/D sky130_fd_sc_hd__a21boi_4
X_81675_ _81275_/CLK _80023_/Y _76874_/A sky130_fd_sc_hd__dfxtp_4
X_69397_ _69288_/A _69397_/B _69397_/X sky130_fd_sc_hd__and2_4
X_86202_ _86490_/CLK _86202_/D _86202_/Q sky130_fd_sc_hd__dfxtp_4
X_59150_ _59085_/X _86069_/Q _59149_/X _59150_/Y sky130_fd_sc_hd__o21ai_4
X_83414_ _83414_/CLK _83414_/D _58480_/A sky130_fd_sc_hd__dfxtp_4
X_56362_ _56351_/A _56363_/B sky130_fd_sc_hd__buf_2
X_80626_ _84777_/Q _65916_/C _80629_/A sky130_fd_sc_hd__xor2_4
X_68348_ _68517_/A _68348_/X sky130_fd_sc_hd__buf_2
X_87182_ _87183_/CLK _87182_/D _44053_/A sky130_fd_sc_hd__dfxtp_4
X_53574_ _53696_/A _53574_/X sky130_fd_sc_hd__buf_2
X_84394_ _84393_/CLK _84394_/D _62636_/C sky130_fd_sc_hd__dfxtp_4
X_50786_ _86133_/Q _50775_/X _50785_/Y _50786_/Y sky130_fd_sc_hd__o21ai_4
X_58101_ _58100_/X _85477_/Q _58062_/X _58101_/X sky130_fd_sc_hd__o21a_4
X_55313_ _55317_/A _55323_/A sky130_fd_sc_hd__buf_2
X_86133_ _86424_/CLK _86133_/D _86133_/Q sky130_fd_sc_hd__dfxtp_4
X_52525_ _52523_/Y _52496_/X _52524_/X _52525_/Y sky130_fd_sc_hd__a21oi_4
X_59081_ _59081_/A _59081_/X sky130_fd_sc_hd__buf_2
X_83345_ _83338_/CLK _71875_/X _83345_/Q sky130_fd_sc_hd__dfxtp_4
X_80557_ _59078_/Y _66016_/Y _80556_/Y _80557_/X sky130_fd_sc_hd__o21a_4
X_56293_ _56368_/A _56270_/B _85247_/Q _56293_/Y sky130_fd_sc_hd__nand3_4
X_68279_ _68338_/A _68279_/X sky130_fd_sc_hd__buf_2
X_70310_ _70246_/A _70328_/A sky130_fd_sc_hd__buf_2
X_58032_ _58017_/X _85387_/Q _58031_/X _58032_/Y sky130_fd_sc_hd__o21ai_4
X_55244_ _55244_/A _55272_/A sky130_fd_sc_hd__buf_2
X_86064_ _85748_/CLK _51155_/Y _86064_/Q sky130_fd_sc_hd__dfxtp_4
X_40470_ _40469_/X _40410_/X _88387_/Q _40411_/X _40470_/X sky130_fd_sc_hd__a2bb2o_4
X_52456_ _52466_/A _53976_/B _52456_/Y sky130_fd_sc_hd__nand2_4
X_71290_ _71289_/Y _71290_/X sky130_fd_sc_hd__buf_2
X_83276_ _83278_/CLK _83276_/D _83276_/Q sky130_fd_sc_hd__dfxtp_4
X_80488_ _80480_/A _80471_/A _80488_/X sky130_fd_sc_hd__and2_4
X_85015_ _85013_/CLK _85015_/D _57401_/B sky130_fd_sc_hd__dfxtp_4
X_51407_ _51405_/Y _51229_/X _51406_/X _86016_/D sky130_fd_sc_hd__a21oi_4
X_70241_ _70239_/A _70239_/B _70241_/C _70239_/D _70241_/X sky130_fd_sc_hd__and4_4
X_82227_ _81094_/CLK _82259_/Q _77473_/A sky130_fd_sc_hd__dfxtp_4
X_55175_ _55174_/X _55177_/A sky130_fd_sc_hd__buf_2
X_52387_ _52373_/X _49135_/X _52387_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_7_102_0_CLK clkbuf_6_51_0_CLK/X clkbuf_8_205_0_CLK/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_290_0_CLK clkbuf_9_145_0_CLK/X _84921_/CLK sky130_fd_sc_hd__clkbuf_1
X_54126_ _85499_/Q _54113_/X _54125_/Y _54126_/Y sky130_fd_sc_hd__o21ai_4
X_42140_ _41134_/X _42137_/X _88015_/Q _42138_/X _88015_/D sky130_fd_sc_hd__a2bb2o_4
X_51338_ _51822_/A _51793_/A sky130_fd_sc_hd__buf_2
X_82158_ _84197_/CLK _84150_/Q _82158_/Q sky130_fd_sc_hd__dfxtp_4
X_70172_ _70154_/X _70232_/A sky130_fd_sc_hd__buf_2
X_59983_ _59881_/X _59971_/X _59979_/Y _59981_/Y _59982_/Y _84679_/D
+ sky130_fd_sc_hd__a41oi_4
Xclkbuf_10_72_0_CLK clkbuf_9_36_0_CLK/X _83013_/CLK sky130_fd_sc_hd__clkbuf_1
X_81109_ _81104_/CLK _79760_/X _81109_/Q sky130_fd_sc_hd__dfxtp_4
X_42071_ _42071_/A _42071_/Y sky130_fd_sc_hd__inv_2
X_58934_ _58641_/A _58934_/X sky130_fd_sc_hd__buf_2
X_54057_ _54055_/Y _54006_/X _54056_/Y _85514_/D sky130_fd_sc_hd__a21boi_4
X_51269_ _64780_/B _51259_/X _51268_/Y _51269_/Y sky130_fd_sc_hd__o21ai_4
X_74980_ _81141_/D _74980_/B _74987_/C sky130_fd_sc_hd__nand2_4
X_86966_ _87397_/CLK _86966_/D _86966_/Q sky130_fd_sc_hd__dfxtp_4
X_82089_ _82008_/CLK _82089_/D _82089_/Q sky130_fd_sc_hd__dfxtp_4
X_41022_ _40999_/X _41000_/X _41021_/X _88292_/Q _40995_/X _41022_/Y
+ sky130_fd_sc_hd__o32ai_4
X_53008_ _53019_/A _52997_/B _53019_/C _53008_/D _53008_/X sky130_fd_sc_hd__and4_4
X_73931_ _72758_/X _86546_/Q _73931_/X sky130_fd_sc_hd__and2_4
X_85917_ _86558_/CLK _51959_/Y _85917_/Q sky130_fd_sc_hd__dfxtp_4
X_58865_ _58749_/A _58941_/A sky130_fd_sc_hd__buf_2
Xclkbuf_7_117_0_CLK clkbuf_6_58_0_CLK/X clkbuf_8_235_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_86897_ _80664_/CLK _45130_/Y _64378_/B sky130_fd_sc_hd__dfxtp_4
X_45830_ _55207_/A _45798_/X _44889_/A _45830_/X sky130_fd_sc_hd__o21a_4
X_57816_ _57726_/X _86012_/Q _57815_/X _57816_/Y sky130_fd_sc_hd__o21ai_4
X_76650_ _81394_/Q _76650_/Y sky130_fd_sc_hd__inv_2
X_85848_ _85558_/CLK _85848_/D _64844_/B sky130_fd_sc_hd__dfxtp_4
X_73862_ _73786_/X _84981_/Q _73859_/X _73861_/X _73863_/B sky130_fd_sc_hd__a211o_4
X_58796_ _58796_/A _58796_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_87_0_CLK clkbuf_9_43_0_CLK/X _83248_/CLK sky130_fd_sc_hd__clkbuf_1
X_75601_ _75594_/Y _75601_/Y sky130_fd_sc_hd__inv_2
X_72813_ _72808_/X _72810_/X _72812_/X _72813_/X sky130_fd_sc_hd__a21o_4
X_45761_ _45761_/A _45746_/B _45761_/Y sky130_fd_sc_hd__nand2_4
X_57747_ _57705_/X _85502_/Q _57736_/X _57747_/X sky130_fd_sc_hd__o21a_4
X_76581_ _76576_/X _76579_/Y _76577_/Y _76614_/C sky130_fd_sc_hd__nand3_4
X_42973_ _42972_/Y _87624_/D sky130_fd_sc_hd__inv_2
X_54959_ _54955_/A _54955_/B _54255_/C _47532_/A _54959_/X sky130_fd_sc_hd__and4_4
Xclkbuf_8_233_0_CLK clkbuf_8_233_0_CLK/A clkbuf_9_467_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_73793_ _73791_/X _73792_/Y _73720_/X _73793_/X sky130_fd_sc_hd__a21o_4
X_85779_ _82956_/CLK _85779_/D _85779_/Q sky130_fd_sc_hd__dfxtp_4
X_47500_ _86628_/Q _47478_/X _47499_/Y _47500_/Y sky130_fd_sc_hd__o21ai_4
X_78320_ _78320_/A _78320_/Y sky130_fd_sc_hd__inv_2
X_44712_ _44528_/A _44712_/X sky130_fd_sc_hd__buf_2
X_75532_ _75530_/Y _75531_/Y _75533_/B _75535_/A sky130_fd_sc_hd__a21oi_4
X_87518_ _87520_/CLK _87518_/D _87518_/Q sky130_fd_sc_hd__dfxtp_4
X_41924_ _41894_/X _41879_/X _40656_/X _73842_/A _41882_/X _41925_/A
+ sky130_fd_sc_hd__o32ai_4
X_48480_ _83582_/Q _73073_/A sky130_fd_sc_hd__inv_2
X_72744_ _73257_/A _72744_/X sky130_fd_sc_hd__buf_2
X_45692_ _55317_/B _45357_/X _45691_/X _45692_/X sky130_fd_sc_hd__o21a_4
X_57678_ _83755_/Q _57678_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_10_0_CLK clkbuf_9_5_0_CLK/X _85213_/CLK sky130_fd_sc_hd__clkbuf_1
X_47431_ _83731_/Q _47431_/Y sky130_fd_sc_hd__inv_2
X_59417_ _58982_/A _59417_/X sky130_fd_sc_hd__buf_2
X_78251_ _78251_/A _78250_/Y _78263_/B sky130_fd_sc_hd__nor2_4
X_44643_ _44638_/X _44639_/X _41045_/A _87020_/Q _44640_/X _44644_/A
+ sky130_fd_sc_hd__o32ai_4
X_56629_ _72664_/C _56629_/B _56630_/A sky130_fd_sc_hd__xnor2_4
X_75463_ _75458_/X _75509_/A _75509_/C _75507_/A sky130_fd_sc_hd__nand3_4
X_41855_ _41839_/X _41841_/X _40532_/X _67245_/B _41835_/X _41856_/A
+ sky130_fd_sc_hd__o32ai_4
X_87449_ _87221_/CLK _87449_/D _87449_/Q sky130_fd_sc_hd__dfxtp_4
X_72675_ _72683_/A _72683_/B _55491_/X _72675_/Y sky130_fd_sc_hd__nand3_4
X_77202_ _77202_/A _77202_/B _77202_/C _77203_/B sky130_fd_sc_hd__nand3_4
X_74414_ _74413_/X _74414_/B _74414_/Y sky130_fd_sc_hd__nand2_4
X_40806_ _40806_/A _40806_/X sky130_fd_sc_hd__buf_2
X_47362_ _86642_/Q _47332_/X _47361_/Y _47362_/Y sky130_fd_sc_hd__o21ai_4
X_59348_ _59331_/X _85413_/Q _59347_/X _59348_/Y sky130_fd_sc_hd__o21ai_4
X_71626_ _71626_/A _71626_/B _71626_/C _71626_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_8_248_0_CLK clkbuf_8_249_0_CLK/A clkbuf_9_497_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_78182_ _78182_/A _78182_/B _78182_/X sky130_fd_sc_hd__xor2_4
X_44574_ _44554_/X _44555_/X _40881_/X _44573_/Y _44557_/X _44574_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75394_ _75393_/A _75393_/B _75394_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_243_0_CLK clkbuf_9_121_0_CLK/X _84454_/CLK sky130_fd_sc_hd__clkbuf_1
X_41786_ _41785_/X _41786_/X sky130_fd_sc_hd__buf_2
X_49101_ _71959_/A _49113_/B sky130_fd_sc_hd__buf_2
X_46313_ _46313_/A _46313_/Y sky130_fd_sc_hd__inv_2
X_77133_ _77134_/A _82293_/D _77141_/B sky130_fd_sc_hd__or2_4
X_43525_ _43524_/Y _87377_/D sky130_fd_sc_hd__inv_2
Xclkbuf_10_873_0_CLK clkbuf_9_436_0_CLK/X _84991_/CLK sky130_fd_sc_hd__clkbuf_1
X_74345_ _74351_/A _74342_/X _55801_/B _74345_/Y sky130_fd_sc_hd__nand3_4
X_40737_ _40737_/A _40765_/B _40737_/X sky130_fd_sc_hd__or2_4
X_47293_ _81818_/Q _47294_/A sky130_fd_sc_hd__inv_2
X_59279_ _59275_/Y _59277_/Y _59278_/X _59279_/X sky130_fd_sc_hd__a21o_4
X_71557_ _71556_/Y _71557_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_25_0_CLK clkbuf_9_12_0_CLK/X _85186_/CLK sky130_fd_sc_hd__clkbuf_1
X_49032_ _49022_/A _53854_/B _49032_/X sky130_fd_sc_hd__and2_4
X_61310_ _61686_/A _72529_/C sky130_fd_sc_hd__buf_2
X_46244_ _44803_/A _46242_/Y _46623_/A _46244_/Y sky130_fd_sc_hd__nand3_4
XPHY_560 sky130_fd_sc_hd__decap_3
X_70508_ _70966_/A _70508_/X sky130_fd_sc_hd__buf_2
X_77064_ _77067_/B _77063_/Y _77065_/B sky130_fd_sc_hd__xnor2_4
X_43456_ _43528_/A _43456_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_364_0_CLK clkbuf_9_365_0_CLK/A clkbuf_9_364_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_62290_ _59931_/X _61811_/X _62289_/X _62290_/X sky130_fd_sc_hd__a21o_4
X_74276_ _74022_/X _86530_/Q _74276_/X sky130_fd_sc_hd__and2_4
XPHY_571 sky130_fd_sc_hd__decap_3
X_40668_ _40635_/X _40638_/X _40667_/X _68735_/B _40612_/X _40669_/A
+ sky130_fd_sc_hd__o32ai_4
X_71488_ _71291_/Y _71488_/X sky130_fd_sc_hd__buf_2
XPHY_582 sky130_fd_sc_hd__decap_3
XPHY_593 sky130_fd_sc_hd__decap_3
X_76015_ _76015_/A _76015_/B _81743_/D sky130_fd_sc_hd__xnor2_4
X_42407_ _42407_/A _42407_/Y sky130_fd_sc_hd__inv_2
X_61241_ _61241_/A _61147_/Y _61241_/X sky130_fd_sc_hd__and2_4
X_73227_ _73227_/A _73228_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_258_0_CLK clkbuf_9_129_0_CLK/X _84250_/CLK sky130_fd_sc_hd__clkbuf_1
X_70439_ _48236_/B _70422_/X _70438_/Y _83774_/D sky130_fd_sc_hd__o21ai_4
X_46175_ _46162_/X _46170_/C _46107_/A _46164_/A _46094_/X _46175_/Y
+ sky130_fd_sc_hd__a2111oi_4
X_43387_ _43217_/A _43397_/A sky130_fd_sc_hd__buf_2
X_40599_ _40599_/A _40599_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_888_0_CLK clkbuf_9_444_0_CLK/X _86246_/CLK sky130_fd_sc_hd__clkbuf_1
X_45126_ _45121_/X _45124_/Y _45125_/X _45126_/Y sky130_fd_sc_hd__a21oi_4
X_42338_ _41681_/X _42325_/X _87914_/Q _42326_/X _87914_/D sky130_fd_sc_hd__a2bb2o_4
X_61172_ _61172_/A _64211_/C _61112_/X _61205_/A _61173_/A sky130_fd_sc_hd__and4_4
X_73158_ _73495_/A _85874_/Q _73158_/X sky130_fd_sc_hd__and2_4
X_60123_ _60122_/Y _60123_/Y sky130_fd_sc_hd__inv_2
X_72109_ _72106_/Y _72107_/X _72108_/Y _83283_/D sky130_fd_sc_hd__a21boi_4
Xclkbuf_9_379_0_CLK clkbuf_9_378_0_CLK/A clkbuf_9_379_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_49934_ _49906_/A _49934_/X sky130_fd_sc_hd__buf_2
X_45057_ _85239_/Q _45056_/X _45012_/X _45057_/X sky130_fd_sc_hd__o21a_4
X_42269_ _42269_/A _42269_/Y sky130_fd_sc_hd__inv_2
X_65980_ _65673_/A _65980_/X sky130_fd_sc_hd__buf_2
X_77966_ _77960_/Y _77967_/C _77967_/B _77980_/A sky130_fd_sc_hd__a21o_4
X_73089_ _87059_/Q _45904_/X _73088_/X _73101_/C sky130_fd_sc_hd__o21ai_4
X_44008_ _44008_/A _57686_/A sky130_fd_sc_hd__buf_2
X_79705_ _79689_/Y _79692_/Y _79705_/X sky130_fd_sc_hd__or2_4
X_64931_ _64804_/A _64931_/B _64931_/X sky130_fd_sc_hd__and2_4
X_60054_ _62198_/B _59985_/A _59943_/X _59910_/X _60055_/A sky130_fd_sc_hd__and4_4
X_76917_ _76917_/A _76917_/B _76918_/B sky130_fd_sc_hd__xnor2_4
Xclkbuf_10_811_0_CLK clkbuf_9_405_0_CLK/X _82558_/CLK sky130_fd_sc_hd__clkbuf_1
X_49865_ _58096_/B _49853_/X _49864_/Y _49865_/Y sky130_fd_sc_hd__o21ai_4
X_77897_ _77902_/A _77902_/B _82036_/D sky130_fd_sc_hd__xor2_4
X_48816_ _48831_/A _48816_/B _48816_/Y sky130_fd_sc_hd__nand2_4
X_67650_ _66560_/X _68402_/A sky130_fd_sc_hd__buf_2
X_79636_ _84210_/Q _72394_/A _79636_/X sky130_fd_sc_hd__xor2_4
X_64862_ _64857_/X _64861_/X _64807_/X _64862_/X sky130_fd_sc_hd__a21o_4
X_76848_ _76846_/Y _76847_/Y _76849_/A sky130_fd_sc_hd__xor2_4
Xclkbuf_9_302_0_CLK clkbuf_9_303_0_CLK/A clkbuf_9_302_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_49796_ _49807_/A _49802_/B _49795_/X _53008_/D _49796_/X sky130_fd_sc_hd__and4_4
X_66601_ _68721_/A _66602_/A sky130_fd_sc_hd__buf_2
X_63813_ _63972_/A _63814_/C sky130_fd_sc_hd__buf_2
X_48747_ _72960_/B _48730_/X _48746_/Y _48747_/Y sky130_fd_sc_hd__o21ai_4
X_67581_ _67226_/A _67581_/X sky130_fd_sc_hd__buf_2
X_79567_ _79566_/B _79567_/Y sky130_fd_sc_hd__inv_2
X_45959_ _44104_/Y _45927_/X _45959_/X sky130_fd_sc_hd__or2_4
X_64793_ _64666_/X _86138_/Q _64766_/X _64792_/X _64793_/X sky130_fd_sc_hd__a211o_4
X_76779_ _76765_/Y _76766_/Y _81486_/Q _81358_/D _76779_/X sky130_fd_sc_hd__a2bb2o_4
X_69320_ _69317_/X _69319_/X _69251_/X _69320_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_10_826_0_CLK clkbuf_9_413_0_CLK/X _82942_/CLK sky130_fd_sc_hd__clkbuf_1
X_66532_ _44019_/A _66565_/A sky130_fd_sc_hd__buf_2
X_78518_ _78482_/B _78513_/Y _78517_/Y _78519_/B sky130_fd_sc_hd__a21oi_4
X_63744_ _63578_/A _63744_/X sky130_fd_sc_hd__buf_2
X_48678_ _74501_/A _48680_/A sky130_fd_sc_hd__buf_2
X_60956_ _63972_/A _63781_/C sky130_fd_sc_hd__buf_2
X_79498_ _79505_/B _79498_/B _82847_/D sky130_fd_sc_hd__xor2_4
X_69251_ _57716_/A _69251_/X sky130_fd_sc_hd__buf_2
X_47629_ _47655_/A _47645_/B _47614_/X _53155_/D _47629_/X sky130_fd_sc_hd__and4_4
Xclkbuf_9_317_0_CLK clkbuf_8_158_0_CLK/X clkbuf_9_317_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_66463_ _66411_/X _66189_/Y _66462_/Y _66463_/Y sky130_fd_sc_hd__o21ai_4
X_78449_ _78448_/X _78475_/B sky130_fd_sc_hd__inv_2
X_63675_ _63697_/A _84910_/Q _63537_/C _63675_/X sky130_fd_sc_hd__and3_4
X_60887_ _60882_/X _60984_/A _60901_/A _60901_/B _61036_/C sky130_fd_sc_hd__nor4_4
X_68202_ _68196_/X _67247_/Y _68189_/X _68201_/Y _68202_/X sky130_fd_sc_hd__a211o_4
X_65414_ _65362_/X _85506_/Q _65363_/X _65413_/X _65414_/X sky130_fd_sc_hd__a211o_4
X_50640_ _50640_/A _53858_/B _50640_/Y sky130_fd_sc_hd__nand2_4
X_62626_ _62653_/A _62653_/B _84395_/Q _62626_/Y sky130_fd_sc_hd__nor3_4
X_81460_ _81461_/CLK _76819_/B _81460_/Q sky130_fd_sc_hd__dfxtp_4
X_69182_ _69182_/A _69182_/X sky130_fd_sc_hd__buf_2
X_66394_ _84131_/Q _66395_/C sky130_fd_sc_hd__inv_2
X_80411_ _80401_/A _80400_/X _80410_/Y _80411_/Y sky130_fd_sc_hd__a21boi_4
Xclkbuf_5_2_0_CLK clkbuf_5_2_0_CLK/A clkbuf_6_5_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_68133_ _68106_/A _68133_/X sky130_fd_sc_hd__buf_2
X_65345_ _65339_/X _65340_/X _65344_/X _65345_/Y sky130_fd_sc_hd__nand3_4
X_50571_ _86175_/Q _50499_/X _50570_/Y _50571_/Y sky130_fd_sc_hd__o21ai_4
X_62557_ _62557_/A _62557_/Y sky130_fd_sc_hd__inv_2
X_81391_ _83926_/CLK _81391_/D _76917_/B sky130_fd_sc_hd__dfxtp_4
X_52310_ _48979_/A _52310_/B _52291_/C _52310_/X sky130_fd_sc_hd__and3_4
X_83130_ _83561_/CLK _83130_/D _83130_/Q sky130_fd_sc_hd__dfxtp_4
X_61508_ _61506_/X _61455_/X _61507_/Y _84475_/D sky130_fd_sc_hd__a21oi_4
X_80342_ _80341_/Y _80350_/A sky130_fd_sc_hd__inv_2
X_68064_ _67948_/X _68049_/Y _67983_/X _68063_/Y _68064_/X sky130_fd_sc_hd__a211o_4
X_53290_ _53276_/A _54469_/B _53290_/Y sky130_fd_sc_hd__nand2_4
X_65276_ _65272_/X _85511_/Q _65146_/X _65275_/X _65276_/X sky130_fd_sc_hd__a211o_4
X_62488_ _62487_/X _62022_/A _62628_/C _62219_/X _62488_/X sky130_fd_sc_hd__and4_4
X_67015_ _67014_/X _67015_/X sky130_fd_sc_hd__buf_2
X_52241_ _52250_/A _48673_/B _52241_/Y sky130_fd_sc_hd__nand2_4
X_64227_ _64250_/A _84856_/Q _64250_/C _64227_/Y sky130_fd_sc_hd__nand3_4
X_83061_ _85581_/CLK _83061_/D _83061_/Q sky130_fd_sc_hd__dfxtp_4
X_61439_ _61429_/A _61438_/X _61429_/C _61439_/Y sky130_fd_sc_hd__nand3_4
X_80273_ _59364_/Y _66345_/C _80273_/Y sky130_fd_sc_hd__nand2_4
X_82012_ _82139_/CLK _82044_/Q _82012_/Q sky130_fd_sc_hd__dfxtp_4
X_52172_ _52169_/Y _52170_/X _52171_/X _52172_/Y sky130_fd_sc_hd__a21oi_4
X_64158_ _58201_/X _64158_/B _64158_/C _64192_/D _64159_/D sky130_fd_sc_hd__nand4_4
X_51123_ _51112_/A _52813_/B _51123_/Y sky130_fd_sc_hd__nand2_4
X_63109_ _63088_/A _84832_/Q _63087_/X _63077_/D _63109_/X sky130_fd_sc_hd__and4_4
X_86820_ _87077_/CLK _86820_/D _86820_/Q sky130_fd_sc_hd__dfxtp_4
X_56980_ _56978_/Y _56979_/Y _56930_/X _56980_/Y sky130_fd_sc_hd__a21oi_4
X_68966_ _87995_/Q _68895_/X _68916_/X _68965_/X _68966_/X sky130_fd_sc_hd__a211o_4
X_64089_ _64084_/Y _64073_/X _64088_/Y _84276_/D sky130_fd_sc_hd__a21oi_4
X_51054_ _86082_/Q _51047_/X _51053_/Y _51054_/Y sky130_fd_sc_hd__o21ai_4
X_67917_ _68429_/A _67917_/X sky130_fd_sc_hd__buf_2
X_55931_ _55947_/A _55931_/B _55931_/X sky130_fd_sc_hd__and2_4
X_86751_ _85535_/CLK _46278_/Y _86751_/Q sky130_fd_sc_hd__dfxtp_4
X_83963_ _80991_/CLK _83963_/D _83963_/Q sky130_fd_sc_hd__dfxtp_4
X_68897_ _87998_/Q _68895_/X _68800_/X _68896_/X _68897_/X sky130_fd_sc_hd__a211o_4
X_50005_ _50025_/A _49994_/X _50005_/C _53217_/D _50005_/X sky130_fd_sc_hd__and4_4
X_85702_ _85700_/CLK _85702_/D _85702_/Q sky130_fd_sc_hd__dfxtp_4
X_58650_ _58007_/A _58650_/X sky130_fd_sc_hd__buf_2
X_82914_ _82925_/CLK _78128_/X _48157_/B sky130_fd_sc_hd__dfxtp_4
X_55862_ _55859_/X _55862_/B _55862_/X sky130_fd_sc_hd__and2_4
X_67848_ _67873_/A _67848_/B _67848_/X sky130_fd_sc_hd__and2_4
X_86682_ _86361_/CLK _86682_/D _59090_/A sky130_fd_sc_hd__dfxtp_4
X_83894_ _82558_/CLK _69830_/X _81966_/D sky130_fd_sc_hd__dfxtp_4
X_57601_ _48067_/A _57619_/B _71960_/C _57601_/X sky130_fd_sc_hd__and3_4
X_54813_ _54758_/A _54823_/A sky130_fd_sc_hd__buf_2
X_85633_ _83161_/CLK _85633_/D _85633_/Q sky130_fd_sc_hd__dfxtp_4
X_58581_ _58571_/X _85792_/Q _58089_/X _58581_/X sky130_fd_sc_hd__o21a_4
X_82845_ _82975_/CLK _82845_/D _82845_/Q sky130_fd_sc_hd__dfxtp_4
X_67779_ _67775_/X _67778_/X _67637_/X _67779_/Y sky130_fd_sc_hd__a21oi_4
X_55793_ _85260_/Q _55177_/A _44045_/X _55792_/X _55793_/X sky130_fd_sc_hd__a211o_4
X_57532_ _57530_/Y _57515_/X _57531_/Y _84985_/D sky130_fd_sc_hd__a21boi_4
X_69518_ _69505_/X _69515_/Y _69516_/X _69517_/Y _69518_/X sky130_fd_sc_hd__a211o_4
X_88352_ _88363_/CLK _40697_/X _88352_/Q sky130_fd_sc_hd__dfxtp_4
X_54744_ _54742_/Y _54720_/X _54743_/X _54744_/Y sky130_fd_sc_hd__a21oi_4
X_85564_ _85561_/CLK _53811_/Y _85564_/Q sky130_fd_sc_hd__dfxtp_4
X_51956_ _50537_/A _51956_/X sky130_fd_sc_hd__buf_2
X_70790_ _70790_/A _70903_/A sky130_fd_sc_hd__buf_2
X_82776_ _82774_/CLK _82776_/D _82968_/D sky130_fd_sc_hd__dfxtp_4
X_87303_ _87813_/CLK _87303_/D _87303_/Q sky130_fd_sc_hd__dfxtp_4
X_84515_ _84503_/CLK _84515_/D _84515_/Q sky130_fd_sc_hd__dfxtp_4
X_50907_ _86109_/Q _50882_/X _50906_/Y _50907_/Y sky130_fd_sc_hd__o21ai_4
X_57463_ _84999_/Q _57463_/B _57463_/X sky130_fd_sc_hd__or2_4
X_81727_ _84014_/CLK _81727_/D _81727_/Q sky130_fd_sc_hd__dfxtp_4
X_69449_ _68923_/X _68925_/X _69418_/X _69449_/Y sky130_fd_sc_hd__a21oi_4
X_88283_ _88283_/CLK _41071_/X _69472_/B sky130_fd_sc_hd__dfxtp_4
X_54675_ _54670_/Y _54666_/X _54674_/X _85399_/D sky130_fd_sc_hd__a21oi_4
X_85495_ _85492_/CLK _85495_/D _85495_/Q sky130_fd_sc_hd__dfxtp_4
X_51887_ _51887_/A _51870_/B _51870_/C _52716_/D _51887_/X sky130_fd_sc_hd__and4_4
X_59202_ _59198_/Y _59201_/Y _59140_/X _59202_/X sky130_fd_sc_hd__a21o_4
X_56414_ _56418_/A _56418_/B _56414_/C _56414_/Y sky130_fd_sc_hd__nand3_4
X_87234_ _87235_/CLK _87234_/D _68793_/B sky130_fd_sc_hd__dfxtp_4
X_53626_ _53687_/A _53626_/X sky130_fd_sc_hd__buf_2
X_41640_ _41636_/X _41638_/X _67365_/B _41639_/X _88178_/D sky130_fd_sc_hd__a2bb2o_4
X_72460_ _72457_/Y _72459_/Y _57718_/A _72460_/X sky130_fd_sc_hd__a21o_4
X_84446_ _84452_/CLK _61914_/Y _78069_/B sky130_fd_sc_hd__dfxtp_4
X_50838_ _51010_/A _50957_/A sky130_fd_sc_hd__buf_2
X_81658_ _81680_/CLK _81690_/Q _81658_/Q sky130_fd_sc_hd__dfxtp_4
X_57394_ _57465_/A _57394_/X sky130_fd_sc_hd__buf_2
X_59133_ _59133_/A _59133_/X sky130_fd_sc_hd__buf_2
X_71411_ _71411_/A _71411_/B _71411_/C _71411_/Y sky130_fd_sc_hd__nor3_4
X_80609_ _80601_/A _80600_/Y _80608_/X _80610_/B sky130_fd_sc_hd__o21ai_4
X_56345_ _56345_/A _56345_/B _55783_/B _56345_/Y sky130_fd_sc_hd__nand3_4
X_41571_ _41570_/X _41530_/X _67087_/B _41531_/X _88190_/D sky130_fd_sc_hd__a2bb2o_4
X_87165_ _86941_/CLK _87165_/D _87165_/Q sky130_fd_sc_hd__dfxtp_4
X_53557_ _54067_/A _53622_/A sky130_fd_sc_hd__buf_2
X_72391_ _72352_/X _85963_/Q _72390_/X _72391_/Y sky130_fd_sc_hd__o21ai_4
X_84377_ _84507_/CLK _62854_/Y _75907_/B sky130_fd_sc_hd__dfxtp_4
X_50769_ _50764_/A _53983_/B _50769_/Y sky130_fd_sc_hd__nand2_4
X_81589_ _81351_/CLK _84189_/Q _81589_/Q sky130_fd_sc_hd__dfxtp_4
X_43310_ _43309_/Y _87488_/D sky130_fd_sc_hd__inv_2
Xclkbuf_7_94_0_CLK clkbuf_7_95_0_CLK/A clkbuf_7_94_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_74130_ _74106_/X _85609_/Q _74107_/X _74129_/X _74130_/X sky130_fd_sc_hd__a211o_4
X_86116_ _85507_/CLK _50873_/Y _86116_/Q sky130_fd_sc_hd__dfxtp_4
X_40522_ _82311_/Q _40467_/B _40522_/X sky130_fd_sc_hd__or2_4
X_52508_ _52309_/A _52509_/B sky130_fd_sc_hd__buf_2
X_59064_ _59060_/Y _59063_/Y _59053_/X _59064_/X sky130_fd_sc_hd__a21o_4
X_71342_ _71137_/B _71342_/B _71343_/A sky130_fd_sc_hd__nor2_4
X_83328_ _83337_/CLK _83328_/D _83328_/Q sky130_fd_sc_hd__dfxtp_4
X_56276_ _56171_/A _56275_/X _56171_/C _56277_/A sky130_fd_sc_hd__nand3_4
X_44290_ _44228_/X _44290_/X sky130_fd_sc_hd__buf_2
X_87096_ _88268_/CLK _87096_/D _87096_/Q sky130_fd_sc_hd__dfxtp_4
X_53488_ _53458_/A _53488_/B _53488_/Y sky130_fd_sc_hd__nand2_4
X_58015_ _58701_/A _58015_/X sky130_fd_sc_hd__buf_2
X_43241_ _43162_/A _43241_/X sky130_fd_sc_hd__buf_2
X_74061_ _74016_/X _85612_/Q _56933_/X _74060_/X _74061_/X sky130_fd_sc_hd__a211o_4
X_55227_ _55227_/A _83315_/Q _55225_/X _55227_/Y sky130_fd_sc_hd__nand3_4
X_86047_ _85535_/CLK _51248_/Y _64643_/B sky130_fd_sc_hd__dfxtp_4
X_40453_ _40437_/X _40443_/X _40452_/X _88389_/Q _40447_/X _40454_/A
+ sky130_fd_sc_hd__o32ai_4
X_52439_ _52185_/A _52466_/A sky130_fd_sc_hd__buf_2
X_83259_ _86282_/CLK _83259_/D _83259_/Q sky130_fd_sc_hd__dfxtp_4
X_71273_ _70638_/A _71276_/D sky130_fd_sc_hd__buf_2
X_73012_ _73093_/A _73012_/B _73012_/X sky130_fd_sc_hd__and2_4
X_70224_ _70238_/A _70224_/X sky130_fd_sc_hd__buf_2
X_43172_ _43121_/A _43172_/X sky130_fd_sc_hd__buf_2
X_55158_ _55158_/A _55172_/A sky130_fd_sc_hd__buf_2
X_40384_ _46317_/A _40385_/B sky130_fd_sc_hd__buf_2
X_42123_ _42120_/X _42116_/X _41087_/X _88024_/Q _42117_/X _42124_/A
+ sky130_fd_sc_hd__o32ai_4
X_54109_ _54245_/A _54217_/A sky130_fd_sc_hd__buf_2
X_77820_ _77806_/Y _77807_/Y _82058_/Q _77819_/Y _77820_/X sky130_fd_sc_hd__a2bb2o_4
X_70155_ _70127_/X _70134_/X _70154_/X _70155_/X sky130_fd_sc_hd__and3_4
X_47980_ _73904_/B _47948_/X _47979_/Y _47980_/Y sky130_fd_sc_hd__o21ai_4
X_55089_ _55093_/A _47762_/Y _55089_/Y sky130_fd_sc_hd__nand2_4
X_59966_ _59917_/X _59909_/Y _59966_/Y sky130_fd_sc_hd__nor2_4
X_87998_ _87748_/CLK _42175_/Y _87998_/Q sky130_fd_sc_hd__dfxtp_4
X_46931_ _86688_/Q _46908_/X _46930_/Y _46931_/Y sky130_fd_sc_hd__o21ai_4
X_42054_ _42053_/Y _42054_/Y sky130_fd_sc_hd__inv_2
X_58917_ _84790_/Q _58871_/X _58911_/X _58916_/X _84790_/D sky130_fd_sc_hd__a2bb2oi_4
X_77751_ _77747_/X _77751_/B _77751_/C _77758_/A sky130_fd_sc_hd__nand3_4
X_74963_ _74971_/A _74963_/B _74964_/B sky130_fd_sc_hd__xor2_4
X_70086_ _69057_/X _69060_/X _69156_/X _70086_/Y sky130_fd_sc_hd__a21oi_4
X_86949_ _88215_/CLK _86949_/D _86949_/Q sky130_fd_sc_hd__dfxtp_4
X_59897_ _59896_/X _59898_/A sky130_fd_sc_hd__buf_2
X_41005_ _40999_/X _41000_/X _41004_/X _88295_/Q _40995_/X _41005_/Y
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_7_32_0_CLK clkbuf_6_16_0_CLK/X clkbuf_8_65_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_76702_ _76699_/X _76700_/Y _76701_/X _76703_/A sky130_fd_sc_hd__a21oi_4
X_49650_ _49570_/A _49650_/X sky130_fd_sc_hd__buf_2
X_73914_ _73912_/X _73913_/Y _73839_/X _73914_/X sky130_fd_sc_hd__a21o_4
X_46862_ _52718_/B _51026_/B sky130_fd_sc_hd__buf_2
X_58848_ _58846_/X _85771_/Q _58847_/X _58848_/X sky130_fd_sc_hd__o21a_4
X_77682_ _77680_/X _77693_/D _77687_/B sky130_fd_sc_hd__and2_4
X_74894_ _74894_/A _74893_/Y _74895_/B sky130_fd_sc_hd__xor2_4
Xclkbuf_8_172_0_CLK clkbuf_7_86_0_CLK/X clkbuf_9_345_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_48601_ _48595_/Y _48403_/X _48600_/Y _86508_/D sky130_fd_sc_hd__a21boi_4
X_79421_ _79408_/X _79419_/X _79420_/X _79421_/Y sky130_fd_sc_hd__a21oi_4
X_45813_ _45811_/Y _45632_/X _45616_/X _45812_/Y _45813_/X sky130_fd_sc_hd__a211o_4
X_76633_ _76633_/A _76633_/Y sky130_fd_sc_hd__inv_2
X_49581_ _49580_/X _52794_/B _49581_/Y sky130_fd_sc_hd__nand2_4
X_73845_ _73845_/A _73873_/B _73845_/Y sky130_fd_sc_hd__nor2_4
X_46793_ _46789_/Y _46751_/X _46792_/X _86703_/D sky130_fd_sc_hd__a21oi_4
X_58779_ _58699_/A _86384_/Q _58779_/Y sky130_fd_sc_hd__nor2_4
X_48532_ _52175_/A _48533_/A sky130_fd_sc_hd__buf_2
X_60810_ _60792_/A _60810_/B _60810_/C _60810_/Y sky130_fd_sc_hd__nor3_4
X_79352_ _84346_/Q _79352_/B _79360_/B sky130_fd_sc_hd__xor2_4
X_45744_ _85131_/Q _45709_/X _45743_/X _45744_/X sky130_fd_sc_hd__o21a_4
X_76564_ _76562_/Y _76563_/X _76564_/X sky130_fd_sc_hd__xor2_4
X_42956_ _42955_/Y _87633_/D sky130_fd_sc_hd__inv_2
X_61790_ _61948_/A _61790_/X sky130_fd_sc_hd__buf_2
X_73776_ _72973_/B _73776_/X sky130_fd_sc_hd__buf_2
X_70988_ _51316_/B _70983_/X _70987_/Y _70988_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_7_47_0_CLK clkbuf_7_47_0_CLK/A clkbuf_8_95_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_78303_ _82593_/Q _78303_/B _78306_/C sky130_fd_sc_hd__xnor2_4
X_75515_ _81087_/Q _75519_/A sky130_fd_sc_hd__inv_2
X_41907_ _51719_/A _41907_/X sky130_fd_sc_hd__buf_2
X_48463_ _48372_/X _82360_/Q _48462_/Y _48464_/A sky130_fd_sc_hd__o21ai_4
X_60741_ _63436_/A _63370_/A sky130_fd_sc_hd__buf_2
X_72727_ _72795_/A _72769_/B sky130_fd_sc_hd__buf_2
X_79283_ _79275_/B _79292_/B _79282_/X _79283_/Y sky130_fd_sc_hd__a21boi_4
X_45675_ _45252_/A _45675_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_187_0_CLK clkbuf_7_93_0_CLK/X clkbuf_9_375_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_76495_ _76491_/X _76492_/Y _76494_/Y _76513_/B sky130_fd_sc_hd__a21o_4
X_42887_ _42832_/A _42887_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_182_0_CLK clkbuf_9_91_0_CLK/X _83325_/CLK sky130_fd_sc_hd__clkbuf_1
X_47414_ _47414_/A _47414_/X sky130_fd_sc_hd__buf_2
X_78234_ _78234_/A _78233_/X _78234_/Y sky130_fd_sc_hd__nand2_4
X_44626_ _44622_/X _44623_/X _40994_/A _87028_/Q _44625_/X _44627_/A
+ sky130_fd_sc_hd__o32ai_4
X_75446_ _75442_/Y _75443_/Y _75445_/Y _75446_/X sky130_fd_sc_hd__or3_4
X_63460_ _58535_/Y _63436_/X _61430_/A _63437_/X _63460_/X sky130_fd_sc_hd__a2bb2o_4
X_41838_ _40485_/X _41813_/X _67028_/B _41814_/X _41838_/X sky130_fd_sc_hd__a2bb2o_4
X_48394_ _48044_/A _47869_/A _48394_/Y sky130_fd_sc_hd__nand2_4
X_60672_ _78080_/A _60323_/X _60647_/Y _60671_/Y _84585_/D sky130_fd_sc_hd__o22a_4
X_72658_ _72630_/X _72658_/X sky130_fd_sc_hd__buf_2
X_62411_ _62120_/A _62411_/X sky130_fd_sc_hd__buf_2
X_47345_ _47333_/X _52995_/B _47345_/Y sky130_fd_sc_hd__nand2_4
X_71609_ _70543_/Y _70573_/B _70568_/D _71606_/X _71609_/Y sky130_fd_sc_hd__nor4_4
X_78165_ _78165_/A _78162_/C _78165_/X sky130_fd_sc_hd__and2_4
X_44557_ _44533_/A _44557_/X sky130_fd_sc_hd__buf_2
X_63391_ _63516_/A _63391_/X sky130_fd_sc_hd__buf_2
X_75377_ _75376_/Y _75377_/Y sky130_fd_sc_hd__inv_2
X_41769_ _41768_/X _41750_/X _88153_/Q _41751_/X _88153_/D sky130_fd_sc_hd__a2bb2o_4
X_72589_ _79352_/B _72445_/X _72587_/Y _72588_/Y _83226_/D sky130_fd_sc_hd__a2bb2oi_4
Xclkbuf_opt_6_CLK _83248_/CLK _84838_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_8_110_0_CLK clkbuf_7_55_0_CLK/X clkbuf_9_220_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_65130_ _65155_/A _65130_/B _65130_/X sky130_fd_sc_hd__and2_4
X_77116_ _77113_/Y _77115_/X _77126_/A sky130_fd_sc_hd__nand2_4
X_43508_ _43507_/Y _87386_/D sky130_fd_sc_hd__inv_2
X_62342_ _62342_/A _62341_/X _76993_/B _62342_/Y sky130_fd_sc_hd__nor3_4
X_74328_ _72704_/A _74338_/A sky130_fd_sc_hd__buf_2
X_47276_ _47270_/Y _47271_/X _47275_/X _47276_/Y sky130_fd_sc_hd__a21oi_4
X_78096_ _82660_/Q _78096_/B _78096_/Y sky130_fd_sc_hd__xnor2_4
Xclkbuf_10_197_0_CLK clkbuf_9_98_0_CLK/X _84660_/CLK sky130_fd_sc_hd__clkbuf_1
X_44488_ _44488_/A _44488_/Y sky130_fd_sc_hd__inv_2
X_49015_ _53848_/B _49015_/X sky130_fd_sc_hd__buf_2
X_46227_ _46227_/A _46227_/Y sky130_fd_sc_hd__inv_2
X_65061_ _65012_/A _65061_/B _65061_/X sky130_fd_sc_hd__and2_4
XPHY_390 sky130_fd_sc_hd__decap_3
X_77047_ _77047_/A _77047_/B _77048_/B sky130_fd_sc_hd__nand2_4
X_43439_ _43439_/A _43439_/Y sky130_fd_sc_hd__inv_2
X_62273_ _62632_/A _63410_/B _62319_/C _62273_/Y sky130_fd_sc_hd__nand3_4
X_74259_ _48141_/A _74259_/B _74259_/X sky130_fd_sc_hd__xor2_4
X_64012_ _64012_/A _64091_/C sky130_fd_sc_hd__buf_2
X_61224_ _61220_/Y _61149_/X _61221_/Y _61190_/X _61223_/Y _84504_/D
+ sky130_fd_sc_hd__a41oi_4
X_46158_ _46158_/A _46158_/B _46158_/C _46158_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_8_125_0_CLK clkbuf_7_62_0_CLK/X clkbuf_9_251_0_CLK/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_120_0_CLK clkbuf_9_60_0_CLK/X _84292_/CLK sky130_fd_sc_hd__clkbuf_1
X_45109_ _45106_/X _45108_/Y _45049_/X _45109_/Y sky130_fd_sc_hd__a21oi_4
X_68820_ _68938_/A _68820_/B _68820_/X sky130_fd_sc_hd__and2_4
X_61155_ _61140_/X _61271_/A sky130_fd_sc_hd__buf_2
X_46089_ _46089_/A _46151_/B _46089_/C _46143_/A _46112_/A sky130_fd_sc_hd__nand4_4
Xclkbuf_10_750_0_CLK clkbuf_9_375_0_CLK/X _87748_/CLK sky130_fd_sc_hd__clkbuf_1
X_78998_ _78998_/A _78998_/B _78998_/Y sky130_fd_sc_hd__nor2_4
X_60106_ _60105_/X _60125_/A sky130_fd_sc_hd__buf_2
X_49917_ _49913_/Y _49897_/X _49916_/X _49917_/Y sky130_fd_sc_hd__a21oi_4
X_68751_ _44705_/A _68394_/X _68421_/X _68750_/X _68751_/X sky130_fd_sc_hd__a211o_4
X_65963_ _58602_/A _66391_/A sky130_fd_sc_hd__buf_2
X_61086_ _61085_/X _61086_/X sky130_fd_sc_hd__buf_2
X_77949_ _77945_/Y _77933_/B _77948_/Y _77950_/B sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_241_0_CLK clkbuf_8_120_0_CLK/X clkbuf_9_241_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_67702_ _67226_/A _67702_/X sky130_fd_sc_hd__buf_2
X_64914_ _64912_/Y _64814_/X _64913_/X _84222_/D sky130_fd_sc_hd__a21o_4
X_60037_ _72564_/A _72604_/B sky130_fd_sc_hd__buf_2
X_49848_ _49827_/X _53060_/B _49848_/Y sky130_fd_sc_hd__nand2_4
X_68682_ _87495_/Q _68626_/X _68601_/X _68681_/X _68682_/X sky130_fd_sc_hd__a211o_4
X_80960_ _81996_/CLK _75554_/B _80960_/Q sky130_fd_sc_hd__dfxtp_4
X_65894_ _65891_/X _65893_/X _65809_/X _65894_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_10_135_0_CLK clkbuf_9_67_0_CLK/X _83787_/CLK sky130_fd_sc_hd__clkbuf_1
X_67633_ _68370_/A _67633_/X sky130_fd_sc_hd__buf_2
X_79619_ _79619_/A _79619_/B _79620_/A sky130_fd_sc_hd__and2_4
Xclkbuf_10_765_0_CLK clkbuf_9_382_0_CLK/X _88056_/CLK sky130_fd_sc_hd__clkbuf_1
X_64845_ _64666_/X _86168_/Q _64766_/X _64844_/X _64845_/X sky130_fd_sc_hd__a211o_4
X_49779_ _49779_/A _49802_/B _49789_/C _52993_/D _49779_/X sky130_fd_sc_hd__and4_4
X_80891_ _80991_/CLK _80891_/D _80891_/Q sky130_fd_sc_hd__dfxtp_4
X_51810_ _51805_/A _51794_/B _51810_/C _46728_/X _51810_/X sky130_fd_sc_hd__and4_4
X_82630_ _82629_/CLK _83982_/Q _78840_/A sky130_fd_sc_hd__dfxtp_4
X_67564_ _87158_/Q _67467_/X _67516_/X _67563_/X _67564_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_9_256_0_CLK clkbuf_8_128_0_CLK/X clkbuf_9_256_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_52790_ _52784_/X _52775_/B _52789_/X _52790_/D _52790_/X sky130_fd_sc_hd__and4_4
X_64776_ _64776_/A _64776_/X sky130_fd_sc_hd__buf_2
X_61988_ _61979_/X _61982_/X _61987_/Y _84849_/Q _61973_/X _61988_/Y
+ sky130_fd_sc_hd__o32ai_4
X_69303_ _88039_/Q _69162_/X _69202_/X _69302_/X _69303_/X sky130_fd_sc_hd__a211o_4
X_66515_ _66512_/Y _59756_/X _66514_/Y _84108_/D sky130_fd_sc_hd__a21o_4
X_51741_ _54317_/A _54286_/C sky130_fd_sc_hd__buf_2
X_63727_ _60879_/D _64012_/A sky130_fd_sc_hd__buf_2
X_82561_ _82558_/CLK _83881_/Q _82561_/Q sky130_fd_sc_hd__dfxtp_4
X_60939_ _64180_/C _60957_/B sky130_fd_sc_hd__inv_2
X_67495_ _60109_/A _67495_/X sky130_fd_sc_hd__buf_2
X_84300_ _84299_/CLK _63702_/Y _80293_/A sky130_fd_sc_hd__dfxtp_4
X_81512_ _84020_/CLK _81512_/D _81512_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_16 sky130_fd_sc_hd__decap_3
X_69234_ _69234_/A _87788_/Q _69234_/X sky130_fd_sc_hd__and2_4
X_54460_ _54478_/A _54460_/B _54460_/Y sky130_fd_sc_hd__nand2_4
X_66446_ _66442_/Y _66414_/X _66445_/Y _66446_/X sky130_fd_sc_hd__a21o_4
X_85280_ _85184_/CLK _56197_/Y _56196_/C sky130_fd_sc_hd__dfxtp_4
X_51672_ _85967_/Q _51647_/X _51671_/Y _51672_/Y sky130_fd_sc_hd__o21ai_4
XPHY_27 sky130_fd_sc_hd__decap_3
X_63658_ _63375_/A _63697_/A sky130_fd_sc_hd__buf_2
X_82492_ _82491_/CLK _82492_/D _82492_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_38 sky130_fd_sc_hd__decap_3
XPHY_49 sky130_fd_sc_hd__decap_3
X_53411_ _53407_/Y _53408_/X _53410_/X _53411_/Y sky130_fd_sc_hd__a21oi_4
X_84231_ _84231_/CLK _84231_/D _64663_/C sky130_fd_sc_hd__dfxtp_4
X_50623_ _86165_/Q _50594_/X _50622_/Y _50623_/Y sky130_fd_sc_hd__o21ai_4
X_62609_ _62288_/X _62285_/X _64535_/B _62609_/D _62609_/X sky130_fd_sc_hd__and4_4
X_81443_ _84079_/CLK _81443_/D _81443_/Q sky130_fd_sc_hd__dfxtp_4
X_69165_ _69755_/A _69165_/B _69165_/X sky130_fd_sc_hd__and2_4
X_54391_ _54389_/Y _54366_/X _54390_/X _85451_/D sky130_fd_sc_hd__a21oi_4
X_66377_ _66377_/A _66377_/X sky130_fd_sc_hd__buf_2
X_63589_ _63556_/X _63582_/X _63583_/X _63587_/X _63588_/Y _63589_/Y
+ sky130_fd_sc_hd__o41ai_4
X_56130_ _56130_/A _56130_/X sky130_fd_sc_hd__buf_2
X_68116_ _84035_/Q _68101_/X _68115_/X _68116_/X sky130_fd_sc_hd__a21bo_4
X_53342_ _85651_/Q _53324_/X _53341_/Y _53342_/Y sky130_fd_sc_hd__o21ai_4
X_65328_ _65272_/X _85541_/Q _65326_/X _65327_/X _65328_/X sky130_fd_sc_hd__a211o_4
X_84162_ _84161_/CLK _84162_/D _84162_/Q sky130_fd_sc_hd__dfxtp_4
X_50554_ _50575_/A _48872_/B _50554_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_703_0_CLK clkbuf_9_351_0_CLK/X _87950_/CLK sky130_fd_sc_hd__clkbuf_1
X_81374_ _83926_/CLK _76934_/Y _81374_/Q sky130_fd_sc_hd__dfxtp_4
X_69096_ _69134_/A _87733_/Q _69096_/X sky130_fd_sc_hd__and2_4
X_83113_ _83846_/CLK _74285_/X _70267_/C sky130_fd_sc_hd__dfxtp_4
X_56061_ _56052_/A _56052_/B _55900_/B _56061_/Y sky130_fd_sc_hd__nand3_4
X_80325_ _84750_/Q _84142_/Q _80325_/X sky130_fd_sc_hd__or2_4
X_68047_ _68025_/A _68047_/B _68047_/X sky130_fd_sc_hd__and2_4
X_53273_ _53302_/A _53293_/C sky130_fd_sc_hd__buf_2
X_65259_ _65172_/X _86120_/Q _65256_/X _65258_/X _65259_/X sky130_fd_sc_hd__a211o_4
X_84093_ _81507_/CLK _84093_/D _80917_/D sky130_fd_sc_hd__dfxtp_4
X_50485_ _50465_/X _48561_/B _50485_/Y sky130_fd_sc_hd__nand2_4
X_55012_ _85335_/Q _54994_/X _55011_/Y _55012_/Y sky130_fd_sc_hd__o21ai_4
X_52224_ _52221_/Y _52203_/X _52223_/X _85865_/D sky130_fd_sc_hd__a21oi_4
X_83044_ _83046_/CLK _74530_/Y _83044_/Q sky130_fd_sc_hd__dfxtp_4
X_87921_ _87922_/CLK _87921_/D _87921_/Q sky130_fd_sc_hd__dfxtp_4
X_80256_ _80253_/X _80256_/B _80256_/X sky130_fd_sc_hd__xor2_4
Xclkbuf_10_718_0_CLK clkbuf_9_359_0_CLK/X _88006_/CLK sky130_fd_sc_hd__clkbuf_1
X_59820_ _59743_/B _59680_/A _72381_/A _59820_/Y sky130_fd_sc_hd__o21ai_4
X_52155_ _85878_/Q _52152_/X _52154_/Y _52155_/Y sky130_fd_sc_hd__o21ai_4
X_87852_ _88104_/CLK _42476_/Y _42475_/A sky130_fd_sc_hd__dfxtp_4
X_80187_ _80187_/A _80186_/X _80187_/Y sky130_fd_sc_hd__xnor2_4
X_69998_ _68497_/X _68499_/X _69925_/X _69998_/Y sky130_fd_sc_hd__a21oi_4
X_51106_ _51104_/Y _51093_/X _51105_/X _51106_/Y sky130_fd_sc_hd__a21oi_4
X_86803_ _87073_/CLK _46034_/Y _86803_/Q sky130_fd_sc_hd__dfxtp_4
X_59751_ _59751_/A _60312_/C sky130_fd_sc_hd__buf_2
Xclkbuf_9_209_0_CLK clkbuf_8_104_0_CLK/X clkbuf_9_209_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_52086_ _66334_/B _52075_/X _52085_/Y _52086_/Y sky130_fd_sc_hd__o21ai_4
X_56963_ _56949_/X _56630_/X _45572_/A _56947_/X _85110_/D sky130_fd_sc_hd__a2bb2o_4
X_68949_ _68994_/A _88252_/Q _68949_/X sky130_fd_sc_hd__and2_4
X_87783_ _87544_/CLK _42660_/Y _87783_/Q sky130_fd_sc_hd__dfxtp_4
X_84995_ _85005_/CLK _57485_/X _55219_/B sky130_fd_sc_hd__dfxtp_4
X_58702_ _58696_/X _58699_/Y _58700_/Y _58603_/X _58701_/X _58702_/X
+ sky130_fd_sc_hd__o32a_4
X_51037_ _51022_/A _51037_/B _51037_/Y sky130_fd_sc_hd__nand2_4
X_55914_ _83033_/Q _55617_/X _44099_/X _55913_/X _55914_/X sky130_fd_sc_hd__a211o_4
X_86734_ _86414_/CLK _86734_/D _86734_/Q sky130_fd_sc_hd__dfxtp_4
X_71960_ _48884_/A _71959_/X _71960_/C _71960_/X sky130_fd_sc_hd__and3_4
X_83946_ _83973_/CLK _83946_/D _80802_/D sky130_fd_sc_hd__dfxtp_4
X_59682_ _59836_/D _59664_/C _59664_/A _59683_/A sky130_fd_sc_hd__nor3_4
X_56894_ _56849_/X _56894_/Y sky130_fd_sc_hd__inv_2
X_70911_ _70925_/A _70914_/C sky130_fd_sc_hd__buf_2
X_58633_ _58659_/A _58633_/B _58633_/Y sky130_fd_sc_hd__nor2_4
X_55845_ _56088_/A _55845_/B _55842_/X _55844_/X _56083_/C sky130_fd_sc_hd__and4_4
X_86665_ _86665_/CLK _47156_/Y _86665_/Q sky130_fd_sc_hd__dfxtp_4
X_71891_ _70530_/Y _71137_/B _71891_/Y sky130_fd_sc_hd__nor2_4
X_83877_ _82557_/CLK _69997_/X _82557_/D sky130_fd_sc_hd__dfxtp_4
X_42810_ _41416_/X _42802_/X _67901_/B _42803_/X _42810_/X sky130_fd_sc_hd__a2bb2o_4
X_73630_ _43032_/Y _73627_/X _73464_/X _73629_/Y _73630_/X sky130_fd_sc_hd__a211o_4
X_85616_ _86576_/CLK _85616_/D _85616_/Q sky130_fd_sc_hd__dfxtp_4
X_70842_ _51765_/B _70831_/X _70841_/Y _70842_/Y sky130_fd_sc_hd__o21ai_4
X_58564_ _58576_/A _86401_/Q _58564_/Y sky130_fd_sc_hd__nor2_4
X_82828_ _82828_/CLK _82828_/D _82828_/Q sky130_fd_sc_hd__dfxtp_4
X_55776_ _55794_/A _85162_/Q _55776_/X sky130_fd_sc_hd__and2_4
X_43790_ _43774_/A _43790_/X sky130_fd_sc_hd__buf_2
X_86596_ _85955_/CLK _86596_/D _86596_/Q sky130_fd_sc_hd__dfxtp_4
X_52988_ _53069_/A _52997_/B sky130_fd_sc_hd__buf_2
X_57515_ _46399_/A _57515_/X sky130_fd_sc_hd__buf_2
X_88335_ _88327_/CLK _88335_/D _69627_/B sky130_fd_sc_hd__dfxtp_4
X_54727_ _54748_/A _54734_/B _54748_/C _47417_/A _54727_/X sky130_fd_sc_hd__and4_4
X_42741_ _42739_/X _42740_/X _41225_/X _68896_/B _42732_/X _42741_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73561_ _73583_/A _73561_/B _73561_/X sky130_fd_sc_hd__and2_4
X_85547_ _85547_/CLK _53894_/Y _85547_/Q sky130_fd_sc_hd__dfxtp_4
X_51939_ _53259_/A _50232_/B _51939_/Y sky130_fd_sc_hd__nand2_4
X_82759_ _82961_/CLK _82759_/D _82759_/Q sky130_fd_sc_hd__dfxtp_4
X_70773_ _70773_/A _70862_/A sky130_fd_sc_hd__buf_2
X_58495_ _58495_/A _58502_/B _58495_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_4_9_0_CLK clkbuf_4_9_0_CLK/A clkbuf_4_9_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_75300_ _80690_/Q _80990_/Q _75301_/B sky130_fd_sc_hd__xor2_4
X_72512_ _72506_/Y _72510_/Y _59654_/X _61281_/C _72511_/Y _72512_/X
+ sky130_fd_sc_hd__a41o_4
X_45460_ _45460_/A _45397_/X _45460_/Y sky130_fd_sc_hd__nor2_4
X_57446_ _57440_/X _57444_/X _57445_/Y _57447_/A sky130_fd_sc_hd__o21ai_4
X_76280_ _76276_/X _76282_/C _76281_/A _76293_/A sky130_fd_sc_hd__a21boi_4
X_88266_ _88268_/CLK _88266_/D _68607_/B sky130_fd_sc_hd__dfxtp_4
X_42672_ _42672_/A _42672_/Y sky130_fd_sc_hd__inv_2
X_54658_ _54667_/A _54674_/B _54644_/X _47294_/A _54658_/X sky130_fd_sc_hd__and4_4
X_73492_ _88310_/Q _73153_/X _72901_/X _73492_/Y sky130_fd_sc_hd__o21ai_4
X_85478_ _84926_/CLK _85478_/D _85478_/Q sky130_fd_sc_hd__dfxtp_4
X_44411_ _41525_/X _44394_/X _87122_/Q _44395_/X _87122_/D sky130_fd_sc_hd__a2bb2o_4
X_75231_ _75230_/X _75245_/A sky130_fd_sc_hd__buf_2
X_41623_ _41623_/A _41623_/Y sky130_fd_sc_hd__inv_2
X_87217_ _87408_/CLK _87217_/D _67395_/B sky130_fd_sc_hd__dfxtp_4
X_53609_ _53607_/Y _53603_/X _53608_/Y _85603_/D sky130_fd_sc_hd__a21boi_4
X_72443_ _72440_/Y _72442_/Y _57779_/X _72443_/X sky130_fd_sc_hd__a21o_4
X_84429_ _84430_/CLK _62156_/Y _78052_/B sky130_fd_sc_hd__dfxtp_4
X_45391_ _85121_/Q _44892_/X _45391_/Y sky130_fd_sc_hd__nor2_4
X_57377_ _57376_/X _57377_/X sky130_fd_sc_hd__buf_2
X_88197_ _87686_/CLK _88197_/D _88197_/Q sky130_fd_sc_hd__dfxtp_4
X_54589_ _54481_/A _54589_/X sky130_fd_sc_hd__buf_2
X_59116_ _58698_/A _59117_/A sky130_fd_sc_hd__buf_2
X_47130_ _47130_/A _47133_/B sky130_fd_sc_hd__buf_2
X_44342_ _44341_/Y _44342_/Y sky130_fd_sc_hd__inv_2
X_56328_ _56332_/A _56335_/B _55846_/B _56328_/Y sky130_fd_sc_hd__nand3_4
X_87148_ _88158_/CLK _87148_/D _87148_/Q sky130_fd_sc_hd__dfxtp_4
X_75162_ _75162_/A _75162_/B _75162_/X sky130_fd_sc_hd__and2_4
X_41554_ _81167_/Q _41584_/B _41554_/X sky130_fd_sc_hd__or2_4
X_72374_ _72361_/X _85676_/Q _72362_/X _72374_/X sky130_fd_sc_hd__o21a_4
X_74113_ _73566_/X _84970_/Q _74087_/X _74112_/X _74114_/B sky130_fd_sc_hd__a211o_4
X_40505_ _40416_/A _81162_/Q _40505_/X sky130_fd_sc_hd__or2_4
X_47061_ _83042_/Q _53345_/B sky130_fd_sc_hd__inv_2
X_59047_ _59027_/X _59044_/Y _59045_/Y _59046_/X _59031_/X _59047_/X
+ sky130_fd_sc_hd__o32a_4
X_71325_ _71337_/A _71335_/A sky130_fd_sc_hd__buf_2
X_44273_ _72739_/A _44272_/X _44273_/Y sky130_fd_sc_hd__nor2_4
X_56259_ _56263_/A _56263_/B _85256_/Q _56259_/Y sky130_fd_sc_hd__nand3_4
X_79970_ _60136_/C _84271_/Q _79973_/A sky130_fd_sc_hd__xor2_4
X_75093_ _75092_/X _81027_/D sky130_fd_sc_hd__buf_2
X_41485_ _41484_/Y _41485_/X sky130_fd_sc_hd__buf_2
X_87079_ _88006_/CLK _44500_/Y _87079_/Q sky130_fd_sc_hd__dfxtp_4
X_46012_ _40506_/Y _46007_/X _67133_/B _46008_/X _86815_/D sky130_fd_sc_hd__a2bb2o_4
X_43224_ _40982_/X _43216_/X _87530_/Q _43218_/X _43224_/X sky130_fd_sc_hd__a2bb2o_4
X_74044_ _73907_/X _84973_/Q _74021_/X _74043_/X _74045_/B sky130_fd_sc_hd__a211o_4
X_78921_ _78921_/A _78921_/Y sky130_fd_sc_hd__inv_2
X_40436_ _40686_/A _44733_/A sky130_fd_sc_hd__buf_2
X_71256_ _71258_/A _71256_/B _71141_/B _71256_/Y sky130_fd_sc_hd__nand3_4
X_70207_ _70214_/A _70214_/B _83197_/Q _70204_/X _70207_/X sky130_fd_sc_hd__and4_4
X_43155_ _43146_/X _43149_/X _40849_/X _87555_/Q _43154_/X _43156_/A
+ sky130_fd_sc_hd__o32ai_4
X_78852_ _82840_/Q _82552_/Q _78852_/X sky130_fd_sc_hd__xor2_4
X_40367_ _40629_/A _40420_/A sky130_fd_sc_hd__buf_2
X_71187_ _70491_/Y _70827_/C _70696_/B _70578_/A _71191_/A sky130_fd_sc_hd__nand4_4
X_42106_ _42099_/X _42094_/X _41036_/X _88033_/Q _42096_/X _42106_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77803_ _77798_/Y _77766_/Y _77802_/Y _77817_/A sky130_fd_sc_hd__o21ai_4
X_70138_ _83529_/Q _83177_/Q _83520_/Q _83168_/Q _70139_/D sky130_fd_sc_hd__a22oi_4
X_47963_ _47963_/A _47963_/B _47963_/X sky130_fd_sc_hd__or2_4
X_59949_ _59943_/X _59950_/C sky130_fd_sc_hd__buf_2
X_43086_ _43189_/A _43086_/X sky130_fd_sc_hd__buf_2
X_78783_ _78783_/A _78782_/Y _78784_/A sky130_fd_sc_hd__nand2_4
Xclkbuf_10_1022_0_CLK clkbuf_9_511_0_CLK/X _86505_/CLK sky130_fd_sc_hd__clkbuf_1
X_75995_ _76005_/A _75994_/Y _81740_/D sky130_fd_sc_hd__xor2_4
X_49702_ _49700_/Y _49677_/X _49701_/X _49702_/Y sky130_fd_sc_hd__a21oi_4
X_46914_ _86690_/Q _46908_/X _46913_/Y _46914_/Y sky130_fd_sc_hd__o21ai_4
X_42037_ _42000_/A _42037_/X sky130_fd_sc_hd__buf_2
X_77734_ _77737_/B _77734_/Y sky130_fd_sc_hd__inv_2
X_74946_ _74937_/Y _74944_/Y _74945_/Y _74946_/X sky130_fd_sc_hd__o21a_4
X_62960_ _62956_/Y _62886_/X _62957_/Y _62958_/Y _62959_/X _62960_/X
+ sky130_fd_sc_hd__a41o_4
X_70069_ _68940_/Y _68823_/X _70056_/X _70068_/Y _70069_/X sky130_fd_sc_hd__a211o_4
X_47894_ _46578_/X _82940_/Q _47893_/X _47895_/B sky130_fd_sc_hd__o21ai_4
X_49633_ _49580_/A _49638_/A sky130_fd_sc_hd__buf_2
X_61911_ _61879_/A _61907_/Y _61908_/Y _61910_/Y _61911_/Y sky130_fd_sc_hd__nand4_4
X_46845_ _46845_/A _46845_/X sky130_fd_sc_hd__buf_2
X_77665_ _77665_/A _77625_/X _77665_/X sky130_fd_sc_hd__or2_4
X_62891_ _62847_/X _63244_/A _62911_/C _62967_/D _62891_/X sky130_fd_sc_hd__and4_4
X_74877_ _74872_/Y _74897_/A _74876_/Y _74878_/B sky130_fd_sc_hd__a21boi_4
X_79404_ _84807_/Q _66420_/C _79404_/X sky130_fd_sc_hd__xor2_4
X_64630_ _64625_/X _64628_/X _64629_/X _64630_/X sky130_fd_sc_hd__a21o_4
X_76616_ _76615_/Y _76616_/B _76616_/X sky130_fd_sc_hd__or2_4
X_49564_ _86364_/Q _49551_/X _49563_/Y _49564_/Y sky130_fd_sc_hd__o21ai_4
X_61842_ _61842_/A _61843_/B sky130_fd_sc_hd__buf_2
X_73828_ _73731_/X _86230_/Q _73804_/X _73827_/X _73828_/X sky130_fd_sc_hd__a211o_4
X_46776_ _46784_/A _46784_/B _46784_/C _46775_/X _46776_/X sky130_fd_sc_hd__and4_4
X_77596_ _77596_/A _77596_/B _82202_/D sky130_fd_sc_hd__xor2_4
X_43988_ _43986_/Y _43954_/X _43945_/A _43987_/Y _43988_/X sky130_fd_sc_hd__a211o_4
X_48515_ _48515_/A _50466_/B _48515_/Y sky130_fd_sc_hd__nand2_4
X_79335_ _79336_/B _79322_/Y _79335_/X sky130_fd_sc_hd__or2_4
X_45727_ _45727_/A _45728_/A sky130_fd_sc_hd__inv_2
X_64561_ _64561_/A _64561_/X sky130_fd_sc_hd__buf_2
X_76547_ _76516_/Y _76543_/X _76546_/X _76547_/Y sky130_fd_sc_hd__a21boi_4
X_42939_ _41768_/X _42930_/X _87641_/Q _42931_/X _87641_/D sky130_fd_sc_hd__a2bb2o_4
X_49495_ _49492_/Y _49487_/X _49494_/X _86377_/D sky130_fd_sc_hd__a21oi_4
X_61773_ _58228_/X _61728_/X _61756_/X _59591_/A _61772_/X _61773_/X
+ sky130_fd_sc_hd__a41o_4
X_73759_ _73711_/A _66024_/B _73759_/X sky130_fd_sc_hd__and2_4
X_66300_ _66297_/X _66299_/X _66240_/X _66300_/X sky130_fd_sc_hd__a21o_4
X_63512_ _63512_/A _84957_/Q _63476_/C _63512_/X sky130_fd_sc_hd__and3_4
X_48446_ _48469_/A _52137_/B _48446_/Y sky130_fd_sc_hd__nand2_4
X_60724_ _60724_/A _60724_/B _60624_/X _60725_/B sky130_fd_sc_hd__nand3_4
X_67280_ _87106_/Q _67230_/X _67278_/X _67279_/X _67280_/X sky130_fd_sc_hd__a211o_4
X_79266_ _84794_/Q _84114_/Q _79266_/X sky130_fd_sc_hd__xor2_4
X_45658_ _45650_/X _45655_/Y _45657_/Y _45658_/Y sky130_fd_sc_hd__a21oi_4
X_64492_ _58348_/A _64511_/B _64492_/Y sky130_fd_sc_hd__nor2_4
X_76478_ _76474_/X _76479_/C _76479_/B _76478_/X sky130_fd_sc_hd__a21o_4
X_66231_ _65969_/A _66231_/X sky130_fd_sc_hd__buf_2
X_78217_ _78214_/Y _78217_/B _78218_/B sky130_fd_sc_hd__xor2_4
X_44609_ _44588_/X _44589_/X _40959_/A _87035_/Q _44590_/X _44609_/Y
+ sky130_fd_sc_hd__o32ai_4
X_63443_ _63443_/A _63465_/C sky130_fd_sc_hd__buf_2
X_75429_ _75413_/A _75413_/B _75411_/Y _75430_/A sky130_fd_sc_hd__o21a_4
X_60655_ _60655_/A _60702_/C sky130_fd_sc_hd__buf_2
X_48377_ _52103_/A _48364_/X _48354_/X _48377_/X sky130_fd_sc_hd__and3_4
X_79197_ _79196_/Y _79197_/B _79197_/Y sky130_fd_sc_hd__nand2_4
X_45589_ _82997_/Q _45401_/X _45588_/X _45589_/Y sky130_fd_sc_hd__o21ai_4
X_47328_ _81814_/Q _47329_/A sky130_fd_sc_hd__inv_2
X_66162_ _66068_/X _65694_/Y _66161_/Y _66162_/Y sky130_fd_sc_hd__o21ai_4
X_78148_ _82571_/Q _82483_/Q _78148_/Y sky130_fd_sc_hd__nor2_4
X_63374_ _63374_/A _61744_/X _63374_/X sky130_fd_sc_hd__and2_4
X_60586_ _60586_/A _60413_/X _60435_/C _60586_/D _60586_/X sky130_fd_sc_hd__and4_4
X_65113_ _65196_/A _65268_/B _84214_/Q _65113_/X sky130_fd_sc_hd__and3_4
X_62325_ _61417_/B _62278_/X _60027_/A _62323_/X _62324_/X _62325_/X
+ sky130_fd_sc_hd__a41o_4
X_47259_ _47259_/A _47260_/A sky130_fd_sc_hd__inv_2
X_66093_ _66090_/Y _66065_/X _66092_/Y _66093_/X sky130_fd_sc_hd__a21o_4
X_78079_ _84584_/Q _78079_/B _78079_/X sky130_fd_sc_hd__xor2_4
X_80110_ _84940_/Q _84188_/Q _80121_/A sky130_fd_sc_hd__xor2_4
X_65044_ _65044_/A _65045_/A sky130_fd_sc_hd__buf_2
X_69921_ _73440_/A _68467_/X _68385_/X _69920_/Y _69921_/X sky130_fd_sc_hd__a211o_4
X_50270_ _50270_/A _74509_/C _50247_/X _50270_/X sky130_fd_sc_hd__and3_4
X_62256_ _62194_/A _58228_/X _62244_/C _62244_/D _62256_/X sky130_fd_sc_hd__and4_4
X_81090_ _83905_/CLK _81090_/D _81090_/Q sky130_fd_sc_hd__dfxtp_4
X_61207_ _64223_/C _61207_/X sky130_fd_sc_hd__buf_2
X_80041_ _80039_/X _80046_/B _80041_/Y sky130_fd_sc_hd__xnor2_4
X_69852_ _69849_/X _69851_/X _69570_/X _69852_/X sky130_fd_sc_hd__a21o_4
X_62187_ _62186_/X _59761_/A _62187_/C _59761_/B _62187_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_9_180_0_CLK clkbuf_8_90_0_CLK/X clkbuf_9_180_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_68803_ _73963_/A _68778_/X _68800_/X _68802_/Y _68803_/X sky130_fd_sc_hd__a211o_4
X_61138_ _61165_/A _61138_/B _84518_/Q _61138_/Y sky130_fd_sc_hd__nor3_4
X_69783_ _69770_/A _88323_/Q _69783_/X sky130_fd_sc_hd__and2_4
X_66995_ _66972_/X _66995_/B _66995_/X sky130_fd_sc_hd__and2_4
X_83800_ _83819_/CLK _70316_/X _74794_/B sky130_fd_sc_hd__dfxtp_4
X_68734_ _68729_/X _68733_/X _68684_/X _68734_/X sky130_fd_sc_hd__a21o_4
X_53960_ _53958_/Y _53948_/X _53959_/Y _85534_/D sky130_fd_sc_hd__a21boi_4
X_65946_ _64714_/X _86238_/Q _65904_/X _65945_/X _65946_/X sky130_fd_sc_hd__a211o_4
X_61069_ _57686_/A _59598_/A _44003_/A _60232_/Y _59551_/A _61070_/C
+ sky130_fd_sc_hd__o41a_4
X_84780_ _83464_/CLK _84780_/D _58987_/A sky130_fd_sc_hd__dfxtp_4
X_81992_ _81989_/CLK _81992_/D _81992_/Q sky130_fd_sc_hd__dfxtp_4
X_52911_ _85732_/Q _52902_/X _52910_/Y _52911_/Y sky130_fd_sc_hd__o21ai_4
X_83731_ _84930_/CLK _83731_/D _83731_/Q sky130_fd_sc_hd__dfxtp_4
X_80943_ _81195_/CLK _80943_/D _74940_/A sky130_fd_sc_hd__dfxtp_4
X_68665_ _64636_/A _69146_/A sky130_fd_sc_hd__buf_2
X_53891_ _85547_/Q _53869_/X _53890_/Y _53891_/Y sky130_fd_sc_hd__o21ai_4
X_65877_ _65877_/A _65878_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_195_0_CLK clkbuf_8_97_0_CLK/X clkbuf_9_195_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_55630_ _55626_/X _55629_/X _44118_/B _55630_/X sky130_fd_sc_hd__a21o_4
X_67616_ _67615_/X _67616_/B _67616_/X sky130_fd_sc_hd__and2_4
X_86450_ _83303_/CLK _86450_/D _86450_/Q sky130_fd_sc_hd__dfxtp_4
X_52842_ _52838_/Y _52839_/X _52841_/X _52842_/Y sky130_fd_sc_hd__a21oi_4
X_64828_ _64828_/A _64828_/X sky130_fd_sc_hd__buf_2
X_83662_ _85447_/CLK _70922_/Y _83662_/Q sky130_fd_sc_hd__dfxtp_4
X_80874_ _80754_/CLK _75648_/B _80874_/Q sky130_fd_sc_hd__dfxtp_4
X_68596_ _86998_/Q _68570_/X _68571_/X _68595_/X _68596_/X sky130_fd_sc_hd__a211o_4
X_85401_ _83745_/CLK _85401_/D _85401_/Q sky130_fd_sc_hd__dfxtp_4
X_82613_ _82518_/CLK _78982_/B _82613_/Q sky130_fd_sc_hd__dfxtp_4
X_55561_ _85051_/Q _55522_/X _55523_/X _55560_/Y _55561_/X sky130_fd_sc_hd__a211o_4
X_67547_ _67572_/A _87210_/Q _67547_/X sky130_fd_sc_hd__and2_4
X_86381_ _86381_/CLK _86381_/D _86381_/Q sky130_fd_sc_hd__dfxtp_4
X_52773_ _52773_/A _52773_/B _52773_/Y sky130_fd_sc_hd__nand2_4
X_64759_ _64836_/A _64759_/B _64759_/X sky130_fd_sc_hd__and2_4
X_83593_ _83589_/CLK _71142_/Y _83593_/Q sky130_fd_sc_hd__dfxtp_4
X_57300_ _57299_/Y _57300_/Y sky130_fd_sc_hd__inv_2
X_88120_ _88376_/CLK _88120_/D _67218_/B sky130_fd_sc_hd__dfxtp_4
X_54512_ _54540_/A _54512_/X sky130_fd_sc_hd__buf_2
X_85332_ _85332_/CLK _85332_/D _85332_/Q sky130_fd_sc_hd__dfxtp_4
X_51724_ _51717_/A _53246_/B _51724_/Y sky130_fd_sc_hd__nand2_4
X_58280_ _58279_/Y _58280_/B _58280_/Y sky130_fd_sc_hd__nand2_4
X_82544_ _83141_/CLK _82544_/D _82544_/Q sky130_fd_sc_hd__dfxtp_4
X_55492_ _55342_/X _55492_/X sky130_fd_sc_hd__buf_2
X_67478_ _67381_/A _86937_/Q _67478_/X sky130_fd_sc_hd__and2_4
X_57231_ _56927_/A _57086_/X _56927_/C _57231_/X sky130_fd_sc_hd__and3_4
X_69217_ _69315_/A _69217_/X sky130_fd_sc_hd__buf_2
X_88051_ _88084_/CLK _88051_/D _88051_/Q sky130_fd_sc_hd__dfxtp_4
X_54443_ _85441_/Q _54431_/X _54442_/Y _54443_/Y sky130_fd_sc_hd__o21ai_4
X_66429_ _66389_/A _66402_/B _66429_/C _66429_/Y sky130_fd_sc_hd__nor3_4
X_85263_ _85198_/CLK _85263_/D _85263_/Q sky130_fd_sc_hd__dfxtp_4
X_51655_ _50256_/A _52620_/A sky130_fd_sc_hd__buf_2
X_82475_ _82563_/CLK _78444_/X _78091_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_642_0_CLK clkbuf_9_321_0_CLK/X _86932_/CLK sky130_fd_sc_hd__clkbuf_1
X_87002_ _86998_/CLK _87002_/D _87002_/Q sky130_fd_sc_hd__dfxtp_4
X_84214_ _84220_/CLK _65114_/X _84214_/Q sky130_fd_sc_hd__dfxtp_4
X_50606_ _50604_/Y _50577_/X _50605_/Y _86169_/D sky130_fd_sc_hd__a21boi_4
X_57162_ _57007_/X _57158_/C _57162_/Y sky130_fd_sc_hd__nand2_4
X_81426_ _81461_/CLK _81426_/D _76042_/B sky130_fd_sc_hd__dfxtp_4
X_69148_ _88050_/Q _68883_/X _68884_/X _69147_/X _69148_/X sky130_fd_sc_hd__a211o_4
X_54374_ _54370_/Y _54366_/X _54373_/X _85454_/D sky130_fd_sc_hd__a21oi_4
X_85194_ _80670_/CLK _85194_/D _85194_/Q sky130_fd_sc_hd__dfxtp_4
X_51586_ _52688_/A _51694_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_133_0_CLK clkbuf_8_66_0_CLK/X clkbuf_9_133_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_56113_ _55811_/X _55802_/X _56114_/A sky130_fd_sc_hd__xnor2_4
Xclkbuf_9_60_0_CLK clkbuf_9_61_0_CLK/A clkbuf_9_60_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_53325_ _53352_/A _53332_/A sky130_fd_sc_hd__buf_2
X_84145_ _84231_/CLK _84145_/D _84145_/Q sky130_fd_sc_hd__dfxtp_4
X_50537_ _50537_/A _50538_/A sky130_fd_sc_hd__buf_2
X_81357_ _81428_/CLK _81357_/D _76312_/A sky130_fd_sc_hd__dfxtp_4
X_69079_ _87478_/Q _68989_/X _69010_/X _69078_/X _69079_/X sky130_fd_sc_hd__a211o_4
X_57093_ _45885_/X _45890_/X _56935_/X _57092_/X _44184_/A _57093_/Y
+ sky130_fd_sc_hd__a41oi_4
X_71110_ _71101_/X _71064_/B _70890_/D _71110_/Y sky130_fd_sc_hd__nand3_4
X_56044_ _56043_/X _56044_/X sky130_fd_sc_hd__buf_2
X_80308_ _80308_/A _80308_/B _80308_/Y sky130_fd_sc_hd__nand2_4
X_41270_ _41096_/B _41280_/B _41270_/X sky130_fd_sc_hd__or2_4
X_53256_ _85667_/Q _51929_/X _53255_/Y _53256_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_657_0_CLK clkbuf_9_328_0_CLK/X _87417_/CLK sky130_fd_sc_hd__clkbuf_1
X_72090_ _71985_/A _72090_/X sky130_fd_sc_hd__buf_2
X_84076_ _84074_/CLK _84076_/D _80900_/D sky130_fd_sc_hd__dfxtp_4
X_50468_ _50510_/A _50497_/C sky130_fd_sc_hd__buf_2
X_81288_ _81288_/CLK _76976_/X _81256_/D sky130_fd_sc_hd__dfxtp_4
X_52207_ _85868_/Q _52184_/X _52206_/Y _52207_/Y sky130_fd_sc_hd__o21ai_4
X_71041_ _70824_/A _71041_/X sky130_fd_sc_hd__buf_2
X_83027_ _85177_/CLK _74581_/Y _45122_/A sky130_fd_sc_hd__dfxtp_4
X_87904_ _87646_/CLK _87904_/D _87904_/Q sky130_fd_sc_hd__dfxtp_4
X_80239_ _80233_/A _80232_/X _80238_/Y _80239_/Y sky130_fd_sc_hd__a21boi_4
X_53187_ _53187_/A _53187_/B _53187_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_148_0_CLK clkbuf_8_74_0_CLK/X clkbuf_9_148_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_50399_ _86208_/Q _50333_/X _50398_/Y _50399_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_75_0_CLK clkbuf_8_37_0_CLK/X clkbuf_9_75_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_59803_ _59802_/X _59803_/X sky130_fd_sc_hd__buf_2
X_52138_ _85881_/Q _52125_/X _52137_/Y _52138_/Y sky130_fd_sc_hd__o21ai_4
X_87835_ _87288_/CLK _87835_/D _68955_/A sky130_fd_sc_hd__dfxtp_4
X_57995_ _57980_/Y _57981_/X _57988_/X _57994_/X _84934_/D sky130_fd_sc_hd__a22oi_4
X_74800_ _70586_/X _83832_/Q _74753_/X _74800_/X sky130_fd_sc_hd__and3_4
X_59734_ _45923_/X _65515_/A sky130_fd_sc_hd__buf_2
X_44960_ _55949_/B _44882_/X _44959_/X _44960_/X sky130_fd_sc_hd__o21a_4
X_52069_ _52065_/Y _52066_/X _52068_/Y _85895_/D sky130_fd_sc_hd__a21boi_4
X_56946_ _44214_/X _56578_/X _45440_/A _56943_/X _85118_/D sky130_fd_sc_hd__a2bb2o_4
X_75780_ _75778_/Y _75779_/Y _75784_/A sky130_fd_sc_hd__xor2_4
X_87766_ _87766_/CLK _87766_/D _69531_/B sky130_fd_sc_hd__dfxtp_4
X_72992_ _72880_/A _72992_/X sky130_fd_sc_hd__buf_2
X_84978_ _86238_/CLK _84978_/D _84978_/Q sky130_fd_sc_hd__dfxtp_4
X_43911_ _41371_/X _43907_/X _67729_/B _43908_/X _87203_/D sky130_fd_sc_hd__a2bb2o_4
X_74731_ _74731_/A _70630_/B _71735_/C _74731_/X sky130_fd_sc_hd__and3_4
X_86717_ _86398_/CLK _86717_/D _86717_/Q sky130_fd_sc_hd__dfxtp_4
X_71943_ _71586_/A _71930_/B _71598_/C _71943_/Y sky130_fd_sc_hd__nor3_4
X_59665_ _59665_/A _59666_/A sky130_fd_sc_hd__buf_2
X_83929_ _83932_/CLK _83929_/D _81393_/D sky130_fd_sc_hd__dfxtp_4
X_44891_ _45387_/A _44891_/X sky130_fd_sc_hd__buf_2
X_56877_ _56876_/X _56877_/X sky130_fd_sc_hd__buf_2
X_87697_ _87950_/CLK _87697_/D _66626_/B sky130_fd_sc_hd__dfxtp_4
X_58616_ _58605_/X _85949_/Q _58568_/X _58616_/X sky130_fd_sc_hd__o21a_4
X_46630_ _54275_/D _51756_/D sky130_fd_sc_hd__buf_2
X_77450_ _77442_/X _77449_/X _77452_/A sky130_fd_sc_hd__xnor2_4
X_43842_ _43842_/A _43842_/X sky130_fd_sc_hd__buf_2
X_74662_ _57416_/A _57416_/C _74656_/X _74662_/Y sky130_fd_sc_hd__nand3_4
X_55828_ _55825_/X _55827_/X _55828_/X sky130_fd_sc_hd__and2_4
X_86648_ _86008_/CLK _86648_/D _86648_/Q sky130_fd_sc_hd__dfxtp_4
X_71874_ _70534_/Y _71883_/B _71873_/X _71874_/D _71874_/Y sky130_fd_sc_hd__nor4_4
X_59596_ _59622_/A _60182_/A _60174_/C sky130_fd_sc_hd__nor2_4
X_76401_ _76396_/X _76400_/C _76391_/X _76401_/X sky130_fd_sc_hd__o21a_4
X_73613_ _73608_/X _73611_/X _73612_/X _73618_/A sky130_fd_sc_hd__a21o_4
X_46561_ _46531_/A _54075_/B _46561_/Y sky130_fd_sc_hd__nand2_4
X_70825_ _71219_/A _71066_/B _70703_/X _70825_/Y sky130_fd_sc_hd__nand3_4
X_58547_ _58547_/A _58548_/A sky130_fd_sc_hd__buf_2
X_77381_ _77381_/A _77381_/Y sky130_fd_sc_hd__inv_2
X_43773_ _40986_/X _43770_/X _69274_/B _43772_/X _43773_/X sky130_fd_sc_hd__a2bb2o_4
X_55759_ _56444_/C _55177_/A _55300_/X _55758_/X _55759_/X sky130_fd_sc_hd__a211o_4
X_74593_ _45182_/A _74582_/X _74592_/X _74593_/Y sky130_fd_sc_hd__o21ai_4
X_86579_ _86578_/CLK _47985_/Y _73904_/B sky130_fd_sc_hd__dfxtp_4
X_40985_ _40504_/X _82295_/Q _40984_/X _40985_/Y sky130_fd_sc_hd__o21ai_4
X_48300_ _48264_/X _52047_/B _48300_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_13_0_CLK clkbuf_8_6_0_CLK/X clkbuf_9_13_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_79120_ _79053_/A _82525_/D sky130_fd_sc_hd__inv_2
X_45512_ _63089_/B _61421_/A sky130_fd_sc_hd__buf_2
X_76332_ _76332_/A _81563_/Q _76332_/Y sky130_fd_sc_hd__nand2_4
X_42724_ _42721_/X _42723_/X _41174_/X _87751_/Q _42700_/X _42725_/A
+ sky130_fd_sc_hd__o32ai_4
X_88318_ _87063_/CLK _40882_/X _88318_/Q sky130_fd_sc_hd__dfxtp_4
X_49280_ _86418_/Q _49204_/X _49279_/Y _49280_/Y sky130_fd_sc_hd__o21ai_4
X_73544_ _73532_/X _73534_/X _73543_/X _73544_/X sky130_fd_sc_hd__a21o_4
X_46492_ _86732_/Q _46474_/X _46491_/Y _46492_/Y sky130_fd_sc_hd__o21ai_4
X_70756_ _53135_/B _70740_/A _70755_/Y _83706_/D sky130_fd_sc_hd__o21ai_4
X_58478_ _58478_/A _58474_/B _58478_/Y sky130_fd_sc_hd__nor2_4
X_48231_ _48190_/A _48231_/B _48231_/Y sky130_fd_sc_hd__nand2_4
X_79051_ _82829_/Q _79051_/B _79053_/A sky130_fd_sc_hd__xnor2_4
X_45443_ _45395_/X _45443_/X sky130_fd_sc_hd__buf_2
X_57429_ _57429_/A _85006_/D sky130_fd_sc_hd__inv_2
X_76263_ _76248_/Y _76245_/Y _76251_/C _76264_/A sky130_fd_sc_hd__o21a_4
X_88249_ _88247_/CLK _88249_/D _88249_/Q sky130_fd_sc_hd__dfxtp_4
X_42655_ _40986_/X _42652_/X _87785_/Q _42653_/X _87785_/D sky130_fd_sc_hd__a2bb2o_4
X_73475_ _73471_/X _73474_/X _72949_/X _73478_/A sky130_fd_sc_hd__a21o_4
X_70687_ _70664_/A _47497_/A _70686_/Y _70687_/X sky130_fd_sc_hd__a21o_4
X_78002_ _78002_/A _78001_/Y _78003_/A sky130_fd_sc_hd__xor2_4
Xclkbuf_9_1_0_CLK clkbuf_8_0_0_CLK/X clkbuf_9_1_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_75214_ _81068_/Q _75214_/B _75233_/B sky130_fd_sc_hd__xnor2_4
X_41606_ _41605_/X _41606_/X sky130_fd_sc_hd__buf_2
X_48162_ _48162_/A _48186_/A sky130_fd_sc_hd__buf_2
X_60440_ _60440_/A _60440_/X sky130_fd_sc_hd__buf_2
X_72426_ _83256_/Q _72381_/X _72418_/X _72425_/X _72426_/Y sky130_fd_sc_hd__a2bb2oi_4
X_45374_ _56280_/C _44880_/X _45373_/X _45374_/Y sky130_fd_sc_hd__o21ai_4
X_76194_ _76168_/B _76179_/Y _76181_/A _76194_/Y sky130_fd_sc_hd__o21ai_4
X_42586_ _42585_/Y _42586_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_9_28_0_CLK clkbuf_9_29_0_CLK/A clkbuf_9_28_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_47113_ _47113_/A _47082_/X _47091_/X _52861_/D _47113_/X sky130_fd_sc_hd__and4_4
X_44325_ _41647_/X _40543_/X _87164_/Q _40544_/X _87164_/D sky130_fd_sc_hd__a2bb2o_4
X_75145_ _75143_/Y _75141_/X _75145_/C _75145_/Y sky130_fd_sc_hd__nand3_4
X_41537_ _41235_/X _41537_/X sky130_fd_sc_hd__buf_2
X_72357_ _72357_/A _72357_/Y sky130_fd_sc_hd__inv_2
X_48093_ _86568_/Q _48049_/X _48092_/Y _48093_/Y sky130_fd_sc_hd__o21ai_4
X_60371_ _60371_/A _60371_/X sky130_fd_sc_hd__buf_2
X_62110_ _61629_/B _62007_/X _62149_/C _62008_/X _62110_/Y sky130_fd_sc_hd__nand4_4
X_47044_ _86676_/Q _47004_/X _47043_/Y _47044_/Y sky130_fd_sc_hd__o21ai_4
X_71308_ _71308_/A _71500_/A sky130_fd_sc_hd__buf_2
X_44256_ _44256_/A _44255_/X _87177_/D sky130_fd_sc_hd__nor2_4
X_63090_ _63084_/Y _63085_/X _63088_/X _63089_/X _63067_/X _63090_/Y
+ sky130_fd_sc_hd__o41ai_4
X_75076_ _75072_/Y _75076_/B _75074_/B _75076_/Y sky130_fd_sc_hd__nand3_4
X_79953_ _79952_/X _79957_/B sky130_fd_sc_hd__buf_2
X_41468_ _41449_/X _82335_/Q _41467_/X _41468_/Y sky130_fd_sc_hd__o21ai_4
X_72288_ _72287_/X _85331_/Q _72225_/X _72288_/X sky130_fd_sc_hd__o21a_4
X_43207_ _43167_/A _43207_/X sky130_fd_sc_hd__buf_2
X_62041_ _61966_/A _62149_/C sky130_fd_sc_hd__buf_2
X_78904_ _78902_/Y _78903_/Y _78908_/A sky130_fd_sc_hd__xor2_4
X_74027_ _74028_/B _74028_/C _74026_/X _74027_/X sky130_fd_sc_hd__a21o_4
X_40419_ _40418_/X _40410_/X _88394_/Q _40411_/X _88394_/D sky130_fd_sc_hd__a2bb2o_4
X_71239_ _71239_/A _71239_/X sky130_fd_sc_hd__buf_2
X_44187_ _44187_/A _72720_/A sky130_fd_sc_hd__buf_2
X_79884_ _84233_/Q _83281_/Q _79887_/A sky130_fd_sc_hd__xor2_4
X_41399_ _41336_/X _41399_/X sky130_fd_sc_hd__buf_2
X_43138_ _43129_/X _43130_/X _40810_/X _43137_/Y _43127_/X _87562_/D
+ sky130_fd_sc_hd__o32ai_4
X_78835_ _78828_/Y _78835_/Y sky130_fd_sc_hd__inv_2
X_48995_ _48995_/A _49022_/A sky130_fd_sc_hd__buf_2
X_65800_ _65789_/X _65233_/Y _65799_/Y _65800_/Y sky130_fd_sc_hd__o21ai_4
X_47946_ _47946_/A _48234_/A _47946_/X sky130_fd_sc_hd__and2_4
X_43069_ _43053_/X _43054_/X _40673_/X _43068_/Y _43058_/X _43069_/Y
+ sky130_fd_sc_hd__o32ai_4
X_66780_ _66757_/X _66771_/Y _66672_/X _66779_/Y _66780_/X sky130_fd_sc_hd__a211o_4
X_78766_ _78764_/Y _78765_/Y _78767_/B _78769_/A sky130_fd_sc_hd__a21oi_4
X_63992_ _64053_/A _59421_/A _63958_/C _63992_/X sky130_fd_sc_hd__and3_4
X_75978_ _75976_/A _75976_/B _75977_/Y _75978_/Y sky130_fd_sc_hd__a21oi_4
X_65731_ _65731_/A _85869_/Q _65731_/X sky130_fd_sc_hd__and2_4
X_77717_ _77717_/A _77718_/B sky130_fd_sc_hd__inv_2
X_62943_ _62930_/A _62930_/B _62943_/C _62943_/Y sky130_fd_sc_hd__nor3_4
X_74929_ _74912_/X _74923_/A _74923_/B _74929_/X sky130_fd_sc_hd__and3_4
X_47877_ _47877_/A _53697_/C sky130_fd_sc_hd__buf_2
X_78697_ _78693_/X _78694_/Y _78696_/Y _78697_/X sky130_fd_sc_hd__a21o_4
X_49616_ _49613_/Y _49596_/X _49615_/X _49616_/Y sky130_fd_sc_hd__a21oi_4
X_68450_ _68450_/A _68450_/X sky130_fd_sc_hd__buf_2
X_46828_ _82955_/Q _46828_/Y sky130_fd_sc_hd__inv_2
X_65662_ _65660_/X _83066_/Q _65568_/X _65661_/X _65662_/X sky130_fd_sc_hd__a211o_4
X_77648_ _77648_/A _81949_/Q _77648_/C _77648_/Y sky130_fd_sc_hd__nand3_4
X_62874_ _62872_/X _62838_/X _62873_/Y _84375_/D sky130_fd_sc_hd__a21oi_4
X_67401_ _67014_/X _67401_/X sky130_fd_sc_hd__buf_2
X_64613_ _45924_/A _65117_/A sky130_fd_sc_hd__buf_2
X_49547_ _86367_/Q _49524_/X _49546_/Y _49547_/Y sky130_fd_sc_hd__o21ai_4
X_61825_ _59684_/X _61839_/B sky130_fd_sc_hd__buf_2
X_68381_ _44149_/A _68380_/Y _68381_/Y sky130_fd_sc_hd__nor2_4
X_46759_ _46733_/A _46758_/X _46759_/Y sky130_fd_sc_hd__nand2_4
X_65593_ _65453_/X _85590_/Q _65470_/X _65592_/X _65593_/X sky130_fd_sc_hd__a211o_4
X_77579_ _81945_/Q _82201_/D _81913_/D sky130_fd_sc_hd__xor2_4
X_67332_ _67093_/X _67333_/A sky130_fd_sc_hd__buf_2
X_79318_ _84798_/Q _84118_/Q _79318_/Y sky130_fd_sc_hd__nand2_4
X_64544_ _64234_/A _64234_/B _64544_/C _64221_/X _64544_/X sky130_fd_sc_hd__and4_4
X_49478_ _49451_/A _49500_/B sky130_fd_sc_hd__buf_2
X_80590_ _80608_/A _80608_/B _80617_/A sky130_fd_sc_hd__xor2_4
X_61756_ _61755_/X _61756_/X sky130_fd_sc_hd__buf_2
X_48429_ _74396_/A _48744_/A sky130_fd_sc_hd__buf_2
X_60707_ _60359_/A _60707_/X sky130_fd_sc_hd__buf_2
X_67263_ _87350_/Q _67239_/X _67240_/X _67262_/X _67263_/X sky130_fd_sc_hd__a211o_4
X_79249_ _79247_/X _79248_/Y _79250_/A sky130_fd_sc_hd__and2_4
X_64475_ _64474_/X _61169_/X _84834_/Q _64475_/Y sky130_fd_sc_hd__nand3_4
X_61687_ _58370_/A _72555_/B _61317_/X _72563_/B _61688_/A sky130_fd_sc_hd__nand4_4
X_69002_ _88089_/Q _68384_/X _68745_/X _69001_/Y _69002_/X sky130_fd_sc_hd__a211o_4
X_66214_ _66011_/X _66214_/B _66214_/X sky130_fd_sc_hd__and2_4
X_51440_ _51430_/X _52969_/B _51440_/Y sky130_fd_sc_hd__nand2_4
X_63426_ _63426_/A _63426_/X sky130_fd_sc_hd__buf_2
X_82260_ _82463_/CLK _80493_/X _82260_/Q sky130_fd_sc_hd__dfxtp_4
X_60638_ _61286_/A _60616_/B _60509_/Y _60638_/Y sky130_fd_sc_hd__nor3_4
X_67194_ _66717_/A _67194_/X sky130_fd_sc_hd__buf_2
X_81211_ _81211_/CLK _74849_/X _48947_/A sky130_fd_sc_hd__dfxtp_4
X_66145_ _66142_/X _66144_/X _65937_/X _66145_/X sky130_fd_sc_hd__a21o_4
X_51371_ _65275_/B _51362_/X _51370_/Y _51371_/Y sky130_fd_sc_hd__o21ai_4
X_63357_ _63356_/X _63357_/X sky130_fd_sc_hd__buf_2
X_82191_ _84945_/CLK _82191_/D _82191_/Q sky130_fd_sc_hd__dfxtp_4
X_60569_ _60435_/C _60562_/Y _60567_/Y _60476_/Y _60568_/Y _60569_/Y
+ sky130_fd_sc_hd__a41oi_4
X_53110_ _85695_/Q _53093_/X _53109_/Y _53110_/Y sky130_fd_sc_hd__o21ai_4
X_50322_ _50356_/A _50322_/B _50322_/Y sky130_fd_sc_hd__nand2_4
X_62308_ _62249_/A _59501_/X _62632_/C _62310_/C sky130_fd_sc_hd__nand3_4
X_81142_ _86758_/CLK _80766_/Q _40648_/A sky130_fd_sc_hd__dfxtp_4
X_54090_ _85506_/Q _54035_/X _54089_/Y _54090_/Y sky130_fd_sc_hd__o21ai_4
X_66076_ _66073_/X _65967_/B _66075_/X _66076_/Y sky130_fd_sc_hd__nand3_4
X_63288_ _63288_/A _64494_/B _63312_/C _63237_/X _63288_/X sky130_fd_sc_hd__and4_4
X_53041_ _53040_/X _53041_/B _53041_/Y sky130_fd_sc_hd__nand2_4
X_65027_ _65024_/X _65026_/X _64851_/X _65031_/A sky130_fd_sc_hd__a21o_4
X_69904_ _69832_/X _69902_/Y _69870_/X _69903_/Y _69904_/X sky130_fd_sc_hd__a211o_4
X_50253_ _86237_/Q _50250_/X _50252_/Y _50253_/Y sky130_fd_sc_hd__o21ai_4
X_62239_ _61329_/B _62628_/C _60027_/A _60011_/X _62238_/X _62239_/X
+ sky130_fd_sc_hd__a41o_4
X_85950_ _82394_/CLK _51769_/Y _85950_/Q sky130_fd_sc_hd__dfxtp_4
X_81073_ _81070_/CLK _81105_/Q _75287_/A sky130_fd_sc_hd__dfxtp_4
X_80024_ _84931_/Q _84179_/Q _80024_/Y sky130_fd_sc_hd__nand2_4
X_84901_ _84727_/CLK _58235_/X _58232_/A sky130_fd_sc_hd__dfxtp_4
X_69835_ _69791_/A _69835_/B _69835_/Y sky130_fd_sc_hd__nor2_4
X_50184_ _50182_/Y _50166_/X _50183_/X _50184_/Y sky130_fd_sc_hd__a21oi_4
X_85881_ _85879_/CLK _85881_/D _85881_/Q sky130_fd_sc_hd__dfxtp_4
X_56800_ _56808_/A _56800_/X sky130_fd_sc_hd__buf_2
X_87620_ _88394_/CLK _87620_/D _87620_/Q sky130_fd_sc_hd__dfxtp_4
X_84832_ _84714_/CLK _84832_/D _84832_/Q sky130_fd_sc_hd__dfxtp_4
X_57780_ _57765_/Y _57775_/Y _57779_/X _57780_/X sky130_fd_sc_hd__a21o_4
X_69766_ _69766_/A _42583_/Y _69766_/Y sky130_fd_sc_hd__nor2_4
X_54992_ _55013_/A _54978_/X _54974_/C _47586_/A _54992_/X sky130_fd_sc_hd__and4_4
X_66978_ _66956_/A _66978_/B _66978_/X sky130_fd_sc_hd__and2_4
X_56731_ _57140_/B _57023_/A sky130_fd_sc_hd__buf_2
X_68717_ _88005_/Q _68715_/X _68540_/X _68716_/X _68717_/X sky130_fd_sc_hd__a211o_4
X_87551_ _87553_/CLK _87551_/D _73275_/A sky130_fd_sc_hd__dfxtp_4
X_53943_ _85537_/Q _53940_/X _53942_/Y _53943_/Y sky130_fd_sc_hd__o21ai_4
X_65929_ _65929_/A _65970_/B sky130_fd_sc_hd__buf_2
X_84763_ _84766_/CLK _84763_/D _84763_/Q sky130_fd_sc_hd__dfxtp_4
X_81975_ _81975_/CLK _81975_/D _81975_/Q sky130_fd_sc_hd__dfxtp_4
X_69697_ _87817_/Q _69698_/B sky130_fd_sc_hd__inv_2
X_86502_ _86499_/CLK _48668_/Y _86502_/Q sky130_fd_sc_hd__dfxtp_4
X_83714_ _83716_/CLK _70728_/Y _46983_/A sky130_fd_sc_hd__dfxtp_4
X_59450_ _84729_/Q _59450_/Y sky130_fd_sc_hd__inv_2
X_56662_ _56661_/Y _83328_/Q _83327_/Q _56682_/A _56663_/A sky130_fd_sc_hd__and4_4
X_80926_ _81169_/CLK _84102_/Q _80926_/Q sky130_fd_sc_hd__dfxtp_4
X_68648_ _67388_/X _68649_/A sky130_fd_sc_hd__buf_2
X_87482_ _87235_/CLK _87482_/D _87482_/Q sky130_fd_sc_hd__dfxtp_4
X_53874_ _53874_/A _53875_/B sky130_fd_sc_hd__buf_2
X_84694_ _84299_/CLK _84694_/D _80422_/A sky130_fd_sc_hd__dfxtp_4
X_58401_ _58388_/X _83346_/Q _58400_/Y _58401_/X sky130_fd_sc_hd__o21a_4
X_55613_ _45426_/A _55641_/A _55611_/X _55612_/Y _55613_/X sky130_fd_sc_hd__a211o_4
X_86433_ _86246_/CLK _49211_/Y _64580_/B sky130_fd_sc_hd__dfxtp_4
X_52825_ _52688_/A _52852_/A sky130_fd_sc_hd__buf_2
X_59381_ _59286_/A _59381_/X sky130_fd_sc_hd__buf_2
X_83645_ _86422_/CLK _83645_/D _46385_/A sky130_fd_sc_hd__dfxtp_4
X_56593_ _56593_/A _73078_/A sky130_fd_sc_hd__buf_2
X_80857_ _80991_/CLK _80889_/Q _75008_/B sky130_fd_sc_hd__dfxtp_4
X_68579_ _68576_/X _68578_/X _68558_/X _68579_/X sky130_fd_sc_hd__a21o_4
X_70610_ _70627_/A _70773_/A sky130_fd_sc_hd__buf_2
X_58332_ _58328_/X _83452_/Q _58331_/Y _84876_/D sky130_fd_sc_hd__o21a_4
X_55544_ _55498_/X _45519_/Y _55544_/Y sky130_fd_sc_hd__nor2_4
X_86364_ _83716_/CLK _86364_/D _86364_/Q sky130_fd_sc_hd__dfxtp_4
X_40770_ _40731_/X _82304_/Q _40769_/X _40770_/Y sky130_fd_sc_hd__o21ai_4
X_52756_ _52620_/A _52757_/A sky130_fd_sc_hd__buf_2
X_71590_ _71859_/A _71590_/B _71582_/X _71590_/Y sky130_fd_sc_hd__nor3_4
X_83576_ _86499_/CLK _71198_/Y _48550_/A sky130_fd_sc_hd__dfxtp_4
X_80788_ _80813_/CLK _80788_/D _75346_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_581_0_CLK clkbuf_9_290_0_CLK/X _81065_/CLK sky130_fd_sc_hd__clkbuf_1
X_88103_ _88111_/CLK _88103_/D _73842_/A sky130_fd_sc_hd__dfxtp_4
X_85315_ _85315_/CLK _55117_/Y _85315_/Q sky130_fd_sc_hd__dfxtp_4
X_51707_ _51717_/A _53232_/B _51707_/Y sky130_fd_sc_hd__nand2_4
X_70541_ _71626_/A _70692_/B _70538_/X _70550_/D _70541_/Y sky130_fd_sc_hd__nor4_4
X_58263_ _58253_/X _83446_/Q _58262_/Y _84894_/D sky130_fd_sc_hd__o21a_4
X_82527_ _82743_/CLK _82527_/D _78767_/B sky130_fd_sc_hd__dfxtp_4
X_55475_ _55468_/X _55475_/X sky130_fd_sc_hd__buf_2
X_86295_ _86611_/CLK _86295_/D _86295_/Q sky130_fd_sc_hd__dfxtp_4
X_52687_ _85773_/Q _52684_/X _52686_/Y _52687_/Y sky130_fd_sc_hd__o21ai_4
X_57214_ _57214_/A _85062_/D sky130_fd_sc_hd__inv_2
X_42440_ _42439_/X _42430_/X _40532_/X _87863_/Q _41967_/A _42440_/Y
+ sky130_fd_sc_hd__o32ai_4
X_88034_ _88034_/CLK _88034_/D _88034_/Q sky130_fd_sc_hd__dfxtp_4
X_54426_ _85444_/Q _54404_/X _54425_/Y _54426_/Y sky130_fd_sc_hd__o21ai_4
X_73260_ _73260_/A _86478_/Q _73260_/X sky130_fd_sc_hd__and2_4
X_85246_ _85248_/CLK _56297_/Y _55958_/B sky130_fd_sc_hd__dfxtp_4
X_51638_ _85973_/Q _51621_/X _51637_/Y _51638_/Y sky130_fd_sc_hd__o21ai_4
X_70472_ _71054_/A _70472_/X sky130_fd_sc_hd__buf_2
X_82458_ _82833_/CLK _82458_/D _82458_/Q sky130_fd_sc_hd__dfxtp_4
X_58194_ _58194_/A _58184_/B _58194_/Y sky130_fd_sc_hd__nor2_4
X_72211_ _72209_/X _85978_/Q _72210_/X _72211_/Y sky130_fd_sc_hd__o21ai_4
X_57145_ _56997_/X _45659_/A _57144_/X _57145_/Y sky130_fd_sc_hd__o21ai_4
X_81409_ _81587_/CLK _83945_/Q _76785_/B sky130_fd_sc_hd__dfxtp_4
X_42371_ _42350_/X _42369_/X _41773_/X _87896_/Q _42370_/X _42371_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54357_ _54329_/A _54362_/B sky130_fd_sc_hd__buf_2
X_73191_ _73190_/X _73191_/B _73191_/X sky130_fd_sc_hd__and2_4
X_85177_ _85177_/CLK _85177_/D _56488_/C sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_596_0_CLK clkbuf_9_298_0_CLK/X _83905_/CLK sky130_fd_sc_hd__clkbuf_1
X_51569_ _85986_/Q _51566_/X _51568_/Y _51569_/Y sky130_fd_sc_hd__o21ai_4
X_82389_ _84766_/CLK _82389_/D _82389_/Q sky130_fd_sc_hd__dfxtp_4
X_44110_ _44109_/X _44110_/X sky130_fd_sc_hd__buf_2
X_41322_ _41239_/X _41241_/X _41321_/X _88236_/Q _41236_/X _41322_/Y
+ sky130_fd_sc_hd__o32ai_4
X_53308_ _53306_/Y _53301_/X _53307_/X _53308_/Y sky130_fd_sc_hd__a21oi_4
X_72142_ _72137_/X _72139_/Y _72140_/Y _59342_/X _72141_/X _72142_/X
+ sky130_fd_sc_hd__o32a_4
X_84128_ _84161_/CLK _66416_/X _66415_/C sky130_fd_sc_hd__dfxtp_4
X_45090_ _55876_/B _45060_/X _45040_/X _45090_/X sky130_fd_sc_hd__o21a_4
X_57076_ _57075_/Y _56903_/X _56952_/A _57076_/X sky130_fd_sc_hd__o21a_4
X_54288_ _54288_/A _46650_/A _54288_/Y sky130_fd_sc_hd__nand2_4
X_56027_ _56023_/A _56017_/B _56027_/C _56027_/Y sky130_fd_sc_hd__nand3_4
X_44041_ _44160_/A _87187_/Q _44041_/Y sky130_fd_sc_hd__nand2_4
X_53239_ _53237_/Y _53215_/X _53238_/X _85671_/D sky130_fd_sc_hd__a21oi_4
X_41253_ _41253_/A _41253_/X sky130_fd_sc_hd__buf_2
X_72073_ _83290_/Q _72051_/X _72072_/Y _72073_/Y sky130_fd_sc_hd__o21ai_4
X_76950_ _81505_/Q _76949_/X _76951_/A sky130_fd_sc_hd__xor2_4
X_84059_ _82648_/CLK _67687_/X _84059_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_6_10_0_CLK clkbuf_5_5_0_CLK/X clkbuf_7_21_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_75901_ _75901_/A _84371_/Q _75901_/X sky130_fd_sc_hd__xor2_4
X_71024_ _70588_/A _71030_/B sky130_fd_sc_hd__buf_2
X_41184_ _41143_/A _41184_/X sky130_fd_sc_hd__buf_2
X_76881_ _76870_/Y _76910_/A _76881_/C _76888_/A sky130_fd_sc_hd__nand3_4
X_47800_ _86596_/Q _47760_/X _47799_/Y _47800_/Y sky130_fd_sc_hd__o21ai_4
X_78620_ _78615_/X _78618_/Y _78610_/X _78621_/A sky130_fd_sc_hd__o21a_4
X_75832_ _75793_/A _75832_/B _75800_/A _75823_/C _75832_/X sky130_fd_sc_hd__and4_4
X_87818_ _83158_/CLK _42565_/Y _87818_/Q sky130_fd_sc_hd__dfxtp_4
X_48780_ _48778_/Y _48760_/X _48779_/X _48780_/Y sky130_fd_sc_hd__a21oi_4
X_57978_ _57975_/Y _57977_/Y _57909_/X _57978_/X sky130_fd_sc_hd__a21o_4
X_45992_ _45980_/X _45987_/X _40451_/X _86824_/Q _45982_/X _45992_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47731_ _47758_/A _47739_/B _47749_/C _53211_/D _47731_/X sky130_fd_sc_hd__and4_4
X_59717_ _59716_/Y _59717_/Y sky130_fd_sc_hd__inv_2
X_78551_ _78551_/A _78554_/B sky130_fd_sc_hd__inv_2
X_44943_ _55958_/B _44874_/X _44926_/X _44943_/X sky130_fd_sc_hd__o21a_4
X_56929_ _85122_/Q _56753_/A _56928_/Y _56929_/X sky130_fd_sc_hd__a21o_4
X_87749_ _87749_/CLK _87749_/D _87749_/Q sky130_fd_sc_hd__dfxtp_4
X_75763_ _75761_/Y _75762_/Y _75766_/A sky130_fd_sc_hd__xor2_4
Xclkbuf_10_534_0_CLK clkbuf_9_267_0_CLK/X _83932_/CLK sky130_fd_sc_hd__clkbuf_1
X_72975_ _88331_/Q _72974_/X _56548_/X _72975_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_6_25_0_CLK clkbuf_6_25_0_CLK/A clkbuf_7_50_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_77502_ _77502_/A _77501_/Y _82196_/D sky130_fd_sc_hd__xor2_4
X_74714_ MACRO_RD_SELECT _74714_/Y sky130_fd_sc_hd__inv_2
X_47662_ _47662_/A _47663_/A sky130_fd_sc_hd__inv_2
X_71926_ _70383_/X _70979_/C _71940_/C _71928_/D _71926_/Y sky130_fd_sc_hd__nand4_4
X_59648_ _59648_/A _59743_/B sky130_fd_sc_hd__buf_2
X_78482_ _78482_/A _78482_/B _82766_/D sky130_fd_sc_hd__xnor2_4
X_44874_ _45197_/A _44874_/X sky130_fd_sc_hd__buf_2
X_75694_ _75694_/A _75696_/A sky130_fd_sc_hd__inv_2
X_49401_ _49397_/A _49420_/B _49408_/C _51787_/D _49401_/X sky130_fd_sc_hd__and4_4
X_46613_ _53097_/A _46892_/A sky130_fd_sc_hd__buf_2
X_77433_ _77433_/A _77433_/Y sky130_fd_sc_hd__inv_2
X_43825_ _43810_/X _43824_/X _41125_/X _68427_/B _43811_/X _43826_/A
+ sky130_fd_sc_hd__o32ai_4
X_74645_ _74691_/A _74645_/X sky130_fd_sc_hd__buf_2
X_47593_ _81242_/Q _47594_/A sky130_fd_sc_hd__inv_2
X_71857_ _71857_/A _71857_/B _71851_/X _71857_/D _71857_/Y sky130_fd_sc_hd__nor4_4
X_59579_ _59579_/A _59657_/A sky130_fd_sc_hd__inv_2
X_49332_ _49327_/X _50854_/B _49332_/Y sky130_fd_sc_hd__nand2_4
X_61610_ _61608_/X _61609_/X _61619_/C _61610_/Y sky130_fd_sc_hd__nand3_4
X_70808_ _52881_/B _70802_/X _70807_/Y _70808_/Y sky130_fd_sc_hd__o21ai_4
X_46544_ _46366_/A _46547_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_549_0_CLK clkbuf_9_274_0_CLK/X _81514_/CLK sky130_fd_sc_hd__clkbuf_1
X_77364_ _77362_/X _77363_/Y _82187_/D sky130_fd_sc_hd__xor2_4
X_43756_ _43756_/A _43756_/X sky130_fd_sc_hd__buf_2
X_62590_ _62570_/A _62140_/X _62601_/C _62623_/D _62590_/X sky130_fd_sc_hd__and4_4
X_74576_ _74575_/X _74569_/X _56069_/Y _74570_/X _74576_/X sky130_fd_sc_hd__a211o_4
X_40968_ _40968_/A _40968_/X sky130_fd_sc_hd__buf_2
X_71788_ _71235_/A _71246_/B _71785_/X _71788_/Y sky130_fd_sc_hd__nand3_4
X_79103_ _79102_/X _79109_/B sky130_fd_sc_hd__inv_2
X_76315_ _76328_/A _81518_/D _76315_/X sky130_fd_sc_hd__xor2_4
X_42707_ _41134_/X _42695_/X _68480_/B _42696_/X _42707_/X sky130_fd_sc_hd__a2bb2o_4
X_49263_ _49263_/A _52478_/B _49263_/Y sky130_fd_sc_hd__nand2_4
X_61541_ _61541_/A _61541_/B _61541_/C _61541_/Y sky130_fd_sc_hd__nand3_4
X_73527_ _73527_/A _72732_/B _73527_/Y sky130_fd_sc_hd__nor2_4
X_46475_ _46623_/A _46491_/A sky130_fd_sc_hd__buf_2
X_70739_ _70755_/A _70740_/A sky130_fd_sc_hd__buf_2
X_77295_ _77296_/A _77294_/Y _77312_/A _77295_/X sky130_fd_sc_hd__a21o_4
X_43687_ _40792_/X _43685_/X _87310_/Q _43686_/X _87310_/D sky130_fd_sc_hd__a2bb2o_4
X_40899_ _40898_/Y _40899_/X sky130_fd_sc_hd__buf_2
X_48214_ _48211_/Y _48175_/X _48213_/Y _48214_/Y sky130_fd_sc_hd__a21boi_4
X_79034_ _79034_/A _79033_/Y _79035_/B sky130_fd_sc_hd__xnor2_4
X_45426_ _45426_/A _45397_/X _45426_/Y sky130_fd_sc_hd__nor2_4
X_64260_ _64377_/A _64275_/A sky130_fd_sc_hd__buf_2
X_76246_ _81257_/Q _81513_/D _76251_/C sky130_fd_sc_hd__nand2_4
X_42638_ _42614_/X _42615_/X _40950_/X _87793_/Q _42637_/X _42639_/A
+ sky130_fd_sc_hd__o32ai_4
X_73458_ _48660_/A _73457_/Y _73458_/X sky130_fd_sc_hd__xor2_4
X_49194_ _49187_/Y _49189_/X _49193_/X _86435_/D sky130_fd_sc_hd__a21oi_4
X_61472_ _61471_/Y _61472_/Y sky130_fd_sc_hd__inv_2
X_63211_ _79330_/A _63189_/X _63210_/Y _63211_/X sky130_fd_sc_hd__a21o_4
X_48145_ _50105_/A _48801_/A sky130_fd_sc_hd__buf_2
X_60423_ _60513_/A _60513_/B _79157_/A _60423_/X sky130_fd_sc_hd__or3_4
X_72409_ _72389_/X _85673_/Q _72308_/X _72409_/X sky130_fd_sc_hd__o21a_4
X_45357_ _45284_/A _45357_/X sky130_fd_sc_hd__buf_2
X_64191_ _84882_/Q _64191_/B _63731_/D _64191_/D _64191_/Y sky130_fd_sc_hd__nand4_4
X_76177_ _76171_/Y _76175_/Y _76176_/Y _76177_/Y sky130_fd_sc_hd__o21ai_4
X_42569_ _42547_/A _42569_/X sky130_fd_sc_hd__buf_2
X_73389_ _48627_/A _73388_/Y _73389_/X sky130_fd_sc_hd__xor2_4
X_44308_ _44308_/A _44308_/X sky130_fd_sc_hd__buf_2
X_63142_ _58551_/A _63131_/X _63117_/X _58326_/A _63118_/X _63142_/Y
+ sky130_fd_sc_hd__o32ai_4
X_75128_ _75113_/A _81061_/Q _75113_/C _75129_/A sky130_fd_sc_hd__a21boi_4
X_48076_ _47972_/A _48086_/B sky130_fd_sc_hd__buf_2
X_60354_ _60353_/Y _60122_/Y _60350_/A _79615_/A _60341_/X _84624_/D
+ sky130_fd_sc_hd__o32a_4
X_45288_ _45283_/Y _45286_/Y _45287_/X _45288_/X sky130_fd_sc_hd__a21o_4
X_47027_ _82390_/Q _54503_/D sky130_fd_sc_hd__inv_2
X_44239_ _44239_/A _44256_/A sky130_fd_sc_hd__buf_2
X_67950_ _69747_/A _67950_/X sky130_fd_sc_hd__buf_2
X_75059_ _75055_/Y _75059_/B _75059_/X sky130_fd_sc_hd__xor2_4
X_79936_ _79935_/Y _79936_/B _79936_/Y sky130_fd_sc_hd__nand2_4
X_63073_ _63010_/A _63073_/X sky130_fd_sc_hd__buf_2
X_60285_ _60285_/A _64386_/A _60285_/Y sky130_fd_sc_hd__nand2_4
X_66901_ _87941_/Q _66875_/X _66807_/X _66900_/X _66901_/X sky130_fd_sc_hd__a211o_4
X_62024_ _61736_/A _62142_/A sky130_fd_sc_hd__buf_2
X_67881_ _87900_/Q _67831_/X _67879_/X _67880_/X _67881_/X sky130_fd_sc_hd__a211o_4
X_79867_ _79859_/A _79858_/Y _79866_/X _79868_/B sky130_fd_sc_hd__o21ai_4
X_69620_ _72855_/A _44299_/A _69617_/X _69619_/Y _69620_/X sky130_fd_sc_hd__a211o_4
X_66832_ _66829_/X _66831_/X _66787_/X _66832_/X sky130_fd_sc_hd__a21o_4
X_78818_ _79122_/A _79122_/B _78818_/C _78818_/Y sky130_fd_sc_hd__nand3_4
X_48978_ _48978_/A _48979_/A sky130_fd_sc_hd__buf_2
X_79798_ _79796_/X _79798_/B _79798_/Y sky130_fd_sc_hd__xnor2_4
X_69551_ _69505_/X _46199_/X _69549_/Y _69550_/Y _69551_/X sky130_fd_sc_hd__a211o_4
X_47929_ _47925_/Y _47903_/X _47928_/X _86585_/D sky130_fd_sc_hd__a21oi_4
X_66763_ _68347_/A _66879_/A sky130_fd_sc_hd__buf_2
X_78749_ _78749_/A _78749_/Y sky130_fd_sc_hd__inv_2
X_63975_ _63968_/Y _63969_/X _63971_/Y _63973_/Y _63974_/X _63975_/X
+ sky130_fd_sc_hd__a41o_4
X_68502_ _68553_/A _87758_/Q _68502_/X sky130_fd_sc_hd__and2_4
X_65714_ _65712_/Y _65681_/X _65713_/X _84183_/D sky130_fd_sc_hd__a21o_4
X_50940_ _86103_/Q _50936_/X _50939_/Y _50940_/Y sky130_fd_sc_hd__o21ai_4
X_62926_ _61618_/X _62926_/B _60255_/B _60228_/A _62928_/C sky130_fd_sc_hd__nand4_4
X_81760_ _81783_/CLK _76142_/B _41634_/B sky130_fd_sc_hd__dfxtp_4
X_69482_ _69383_/A _87258_/Q _69482_/X sky130_fd_sc_hd__and2_4
X_66694_ _66669_/A _66694_/B _66694_/X sky130_fd_sc_hd__and2_4
X_68433_ _68430_/X _68432_/X _68331_/X _68433_/Y sky130_fd_sc_hd__a21oi_4
X_80711_ _80679_/CLK _75897_/X _80679_/D sky130_fd_sc_hd__dfxtp_4
X_65645_ _65596_/X _83067_/Q _65540_/X _65644_/X _65645_/X sky130_fd_sc_hd__a211o_4
X_50871_ _86116_/Q _50856_/X _50870_/Y _50871_/Y sky130_fd_sc_hd__o21ai_4
X_62857_ _62869_/A _62812_/B _61997_/X _62857_/Y sky130_fd_sc_hd__nand3_4
X_81691_ _81632_/CLK _80191_/Y _76728_/A sky130_fd_sc_hd__dfxtp_4
X_52610_ _52614_/A _52605_/X _52622_/C _50919_/D _52610_/X sky130_fd_sc_hd__and4_4
X_83430_ _83431_/CLK _71638_/Y _83430_/Q sky130_fd_sc_hd__dfxtp_4
X_61808_ _59668_/B _61809_/C sky130_fd_sc_hd__buf_2
X_80642_ _80642_/HI THREAD_COUNT[3] sky130_fd_sc_hd__conb_1
X_68364_ _68392_/A _68757_/A sky130_fd_sc_hd__buf_2
X_53590_ _53793_/A _53604_/A sky130_fd_sc_hd__buf_2
X_65576_ _64902_/A _65576_/X sky130_fd_sc_hd__buf_2
X_62788_ _62847_/A _62789_/A sky130_fd_sc_hd__buf_2
Xclkbuf_8_8_0_CLK clkbuf_8_9_0_CLK/A clkbuf_8_8_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_67315_ _88372_/Q _67311_/X _67313_/X _67314_/X _67315_/X sky130_fd_sc_hd__a211o_4
X_52541_ _52486_/A _52541_/X sky130_fd_sc_hd__buf_2
X_64527_ _58985_/A _64226_/X _64526_/Y _64527_/Y sky130_fd_sc_hd__o21ai_4
X_83361_ _83756_/CLK _83361_/D _83361_/Q sky130_fd_sc_hd__dfxtp_4
X_61739_ _61842_/A _62149_/B sky130_fd_sc_hd__buf_2
X_80573_ _80557_/X _80561_/B _80572_/X _80573_/X sky130_fd_sc_hd__a21o_4
X_68295_ _68737_/A _68295_/X sky130_fd_sc_hd__buf_2
XPHY_208 sky130_fd_sc_hd__decap_3
XPHY_219 sky130_fd_sc_hd__decap_3
X_85100_ _85100_/CLK _57022_/Y _45719_/A sky130_fd_sc_hd__dfxtp_4
X_82312_ _80835_/CLK _77044_/B _82312_/Q sky130_fd_sc_hd__dfxtp_4
X_55260_ _55257_/X _55259_/X _55138_/X _55264_/A sky130_fd_sc_hd__a21o_4
X_86080_ _85761_/CLK _86080_/D _86080_/Q sky130_fd_sc_hd__dfxtp_4
X_67246_ _88375_/Q _67193_/X _67194_/X _67245_/X _67246_/X sky130_fd_sc_hd__a211o_4
X_52472_ _52476_/A _46367_/Y _52472_/Y sky130_fd_sc_hd__nand2_4
X_64458_ _64223_/A _64458_/B _64545_/C _64458_/X sky130_fd_sc_hd__and3_4
X_83292_ _85538_/CLK _72065_/Y _83292_/Q sky130_fd_sc_hd__dfxtp_4
X_54211_ _54215_/A _47431_/Y _54211_/Y sky130_fd_sc_hd__nand2_4
X_85031_ _85031_/CLK _57351_/Y _57349_/B sky130_fd_sc_hd__dfxtp_4
X_51423_ _51419_/Y _51420_/X _51422_/X _51423_/Y sky130_fd_sc_hd__a21oi_4
X_63409_ _63471_/A _63410_/D sky130_fd_sc_hd__buf_2
X_82243_ _81859_/CLK _80287_/X _82243_/Q sky130_fd_sc_hd__dfxtp_4
X_55191_ _55711_/A _55192_/A sky130_fd_sc_hd__buf_2
X_67177_ _67131_/A _87610_/Q _67177_/X sky130_fd_sc_hd__and2_4
X_64389_ _59421_/A _64418_/B _64389_/Y sky130_fd_sc_hd__nor2_4
X_54142_ _54149_/A _47306_/A _54142_/Y sky130_fd_sc_hd__nand2_4
X_66128_ _66125_/X _86226_/Q _66021_/X _66127_/X _66128_/X sky130_fd_sc_hd__a211o_4
X_51354_ _51350_/A _49320_/B _51354_/Y sky130_fd_sc_hd__nand2_4
X_82174_ _82575_/CLK _84166_/Q _77994_/A sky130_fd_sc_hd__dfxtp_4
X_50305_ _50303_/Y _50299_/X _50304_/Y _86227_/D sky130_fd_sc_hd__a21boi_4
X_81125_ _81125_/CLK _81125_/D _40741_/A sky130_fd_sc_hd__dfxtp_4
X_58950_ _58796_/X _86083_/Q _58949_/X _58950_/Y sky130_fd_sc_hd__o21ai_4
X_54073_ _54068_/X _54073_/B _54073_/Y sky130_fd_sc_hd__nand2_4
X_66059_ _65980_/X _86551_/Q _66059_/X sky130_fd_sc_hd__and2_4
X_51285_ _51259_/A _51285_/X sky130_fd_sc_hd__buf_2
X_86982_ _86982_/CLK _86982_/D _86982_/Q sky130_fd_sc_hd__dfxtp_4
X_53024_ _53022_/Y _53001_/X _53023_/X _53024_/Y sky130_fd_sc_hd__a21oi_4
X_57901_ _64713_/A _58876_/A sky130_fd_sc_hd__buf_2
X_50236_ _50595_/A _50505_/A sky130_fd_sc_hd__buf_2
X_85933_ _86091_/CLK _51861_/Y _85933_/Q sky130_fd_sc_hd__dfxtp_4
X_81056_ _85332_/CLK _75550_/Y _81056_/Q sky130_fd_sc_hd__dfxtp_4
X_58881_ _58787_/X _86089_/Q _58880_/X _58881_/Y sky130_fd_sc_hd__o21ai_4
X_80007_ _80005_/X _80006_/X _80007_/Y sky130_fd_sc_hd__xnor2_4
X_57832_ _57806_/X _57832_/B _57832_/Y sky130_fd_sc_hd__nor2_4
X_69818_ _69746_/X _69813_/Y _69815_/X _69817_/Y _69818_/X sky130_fd_sc_hd__a211o_4
X_50167_ _50677_/A _51256_/B _50147_/C _50167_/X sky130_fd_sc_hd__and3_4
X_85864_ _85859_/CLK _85864_/D _85864_/Q sky130_fd_sc_hd__dfxtp_4
X_87603_ _88108_/CLK _87603_/D _73554_/A sky130_fd_sc_hd__dfxtp_4
X_84815_ _84815_/CLK _84815_/D _84815_/Q sky130_fd_sc_hd__dfxtp_4
X_57763_ _58793_/A _57763_/X sky130_fd_sc_hd__buf_2
X_69749_ _68587_/X _69749_/B _69749_/Y sky130_fd_sc_hd__nor2_4
X_50098_ _50096_/Y _50092_/X _50097_/X _86265_/D sky130_fd_sc_hd__a21oi_4
X_54975_ _54970_/Y _54971_/X _54974_/X _54975_/Y sky130_fd_sc_hd__a21oi_4
X_85795_ _86736_/CLK _85795_/D _65375_/B sky130_fd_sc_hd__dfxtp_4
X_59502_ _59501_/X _58532_/X _59502_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_4_0_1_CLK clkbuf_4_0_1_CLK/A clkbuf_4_0_1_CLK/X sky130_fd_sc_hd__clkbuf_1
X_56714_ _45890_/X _44228_/X _56663_/X _56714_/Y sky130_fd_sc_hd__a21oi_4
X_87534_ _88084_/CLK _87534_/D _87534_/Q sky130_fd_sc_hd__dfxtp_4
X_41940_ _41937_/X _41919_/X _40673_/X _41938_/Y _41939_/X _88100_/D
+ sky130_fd_sc_hd__o32ai_4
X_53926_ _53924_/Y _53914_/X _53925_/Y _85541_/D sky130_fd_sc_hd__a21boi_4
X_72760_ _72755_/X _83081_/Q _45885_/X _72759_/X _72761_/B sky130_fd_sc_hd__a211o_4
X_84746_ _84746_/CLK _59385_/Y _84746_/Q sky130_fd_sc_hd__dfxtp_4
X_57694_ _64601_/A _57694_/X sky130_fd_sc_hd__buf_2
X_81958_ _82301_/CLK _83886_/Q _81958_/Q sky130_fd_sc_hd__dfxtp_4
X_71711_ _71711_/A _70698_/B _71711_/Y sky130_fd_sc_hd__nor2_4
X_59433_ _59433_/A _59433_/Y sky130_fd_sc_hd__inv_2
X_80909_ _84087_/CLK _84085_/Q _80909_/Q sky130_fd_sc_hd__dfxtp_4
X_56645_ _83332_/Q _56645_/Y sky130_fd_sc_hd__inv_2
X_87465_ _87210_/CLK _87465_/D _87465_/Q sky130_fd_sc_hd__dfxtp_4
X_41871_ _41880_/A _41872_/A sky130_fd_sc_hd__buf_2
X_53857_ _85554_/Q _53846_/X _53856_/Y _53857_/Y sky130_fd_sc_hd__o21ai_4
X_72691_ _72697_/A _72697_/B _55200_/C _72691_/Y sky130_fd_sc_hd__nand3_4
X_84677_ _84393_/CLK _84677_/D _59992_/C sky130_fd_sc_hd__dfxtp_4
X_81889_ _82436_/CLK _78080_/X _81857_/D sky130_fd_sc_hd__dfxtp_4
X_43610_ _43610_/A _68468_/B sky130_fd_sc_hd__inv_2
X_74430_ _74492_/A _74430_/X sky130_fd_sc_hd__buf_2
X_86416_ _86414_/CLK _86416_/D _65054_/B sky130_fd_sc_hd__dfxtp_4
X_40822_ _40756_/A _40822_/X sky130_fd_sc_hd__buf_2
X_52808_ _85750_/Q _52792_/X _52807_/Y _52808_/Y sky130_fd_sc_hd__o21ai_4
X_71642_ _71637_/A _71256_/B _71644_/C _71642_/Y sky130_fd_sc_hd__nand3_4
X_59364_ _84747_/Q _59364_/Y sky130_fd_sc_hd__inv_2
X_83628_ _83627_/CLK _83628_/D _83628_/Q sky130_fd_sc_hd__dfxtp_4
X_44590_ _44549_/A _44590_/X sky130_fd_sc_hd__buf_2
X_56576_ _56568_/X _56575_/X _55622_/B _56572_/X _85151_/D sky130_fd_sc_hd__a2bb2o_4
X_87396_ _87144_/CLK _87396_/D _87396_/Q sky130_fd_sc_hd__dfxtp_4
X_53788_ _53733_/A _53806_/B sky130_fd_sc_hd__buf_2
X_58315_ _58310_/X _83457_/Q _58314_/Y _58315_/X sky130_fd_sc_hd__o21a_4
X_55527_ _55507_/X _55527_/X sky130_fd_sc_hd__buf_2
X_43541_ _43540_/Y _87368_/D sky130_fd_sc_hd__inv_2
X_74361_ _45954_/X _58334_/A _56167_/A _74361_/Y sky130_fd_sc_hd__nand3_4
X_86347_ _86351_/CLK _86347_/D _86347_/Q sky130_fd_sc_hd__dfxtp_4
X_52739_ _52744_/A _52739_/B _52739_/Y sky130_fd_sc_hd__nand2_4
X_40753_ _40753_/A _40753_/X sky130_fd_sc_hd__buf_2
X_71573_ _71556_/Y _83452_/Q _71572_/Y _71573_/X sky130_fd_sc_hd__a21o_4
X_59295_ _59219_/X _85737_/Q _59220_/X _59295_/X sky130_fd_sc_hd__o21a_4
X_83559_ _86592_/CLK _71249_/Y _83559_/Q sky130_fd_sc_hd__dfxtp_4
X_76100_ _81530_/Q _76100_/B _76100_/X sky130_fd_sc_hd__xor2_4
X_73312_ _73312_/A _73311_/X _73313_/B sky130_fd_sc_hd__nand2_4
X_46260_ _46347_/A _46288_/A sky130_fd_sc_hd__buf_2
X_70524_ _70526_/A _70954_/B _70962_/C _70524_/Y sky130_fd_sc_hd__nand3_4
X_58246_ _58246_/A _58246_/Y sky130_fd_sc_hd__inv_2
X_77080_ _77080_/A _77079_/Y _77081_/B sky130_fd_sc_hd__xor2_4
X_43472_ _43518_/A _43472_/X sky130_fd_sc_hd__buf_2
X_55458_ _55457_/X _55458_/X sky130_fd_sc_hd__buf_2
X_74292_ _70273_/A _74288_/X _74291_/Y _74292_/X sky130_fd_sc_hd__a21bo_4
X_86278_ _85957_/CLK _86278_/D _72436_/B sky130_fd_sc_hd__dfxtp_4
X_40684_ _40635_/X _40638_/X _40682_/X _88354_/Q _40683_/X _40685_/A
+ sky130_fd_sc_hd__o32ai_4
X_45211_ _85197_/Q _45176_/X _45210_/X _45211_/Y sky130_fd_sc_hd__o21ai_4
X_76031_ _76031_/A _76030_/Y _81745_/D sky130_fd_sc_hd__xor2_4
X_42423_ _42417_/X _42410_/X _40491_/X _87871_/Q _42411_/X _42424_/A
+ sky130_fd_sc_hd__o32ai_4
X_88017_ _87776_/CLK _42135_/Y _88017_/Q sky130_fd_sc_hd__dfxtp_4
X_54409_ _54407_/Y _54394_/X _54408_/X _85448_/D sky130_fd_sc_hd__a21oi_4
X_73243_ _73230_/X _73232_/Y _73242_/X _73243_/X sky130_fd_sc_hd__a21o_4
X_85229_ _85192_/CLK _85229_/D _56341_/C sky130_fd_sc_hd__dfxtp_4
X_46191_ _86762_/Q _46125_/A _46196_/A sky130_fd_sc_hd__or2_4
X_70455_ _70454_/Y _70455_/Y sky130_fd_sc_hd__inv_2
X_58177_ _58177_/A _58177_/Y sky130_fd_sc_hd__inv_2
X_55389_ _56719_/A _56719_/B _55388_/Y _55389_/Y sky130_fd_sc_hd__a21oi_4
X_45142_ _45139_/X _45141_/Y _45125_/X _45142_/Y sky130_fd_sc_hd__a21oi_4
X_57128_ _83334_/Q _83333_/Q _56675_/X _56876_/X _57129_/A sky130_fd_sc_hd__nand4_4
X_42354_ _41721_/X _42342_/X _87906_/Q _42343_/X _42354_/X sky130_fd_sc_hd__a2bb2o_4
X_73174_ _88323_/Q _72731_/X _56548_/X _73174_/Y sky130_fd_sc_hd__o21ai_4
X_70386_ DATA_TO_HASH[3] _70387_/A sky130_fd_sc_hd__buf_2
X_41305_ _41290_/X _82909_/Q _41304_/X _41305_/Y sky130_fd_sc_hd__o21ai_4
X_72125_ _59381_/X _85985_/Q _72124_/X _72125_/Y sky130_fd_sc_hd__o21ai_4
X_49950_ _86293_/Q _49934_/X _49949_/Y _49950_/Y sky130_fd_sc_hd__o21ai_4
X_45073_ _45297_/A _45073_/X sky130_fd_sc_hd__buf_2
X_57059_ _57057_/X _57058_/Y _56953_/X _57059_/Y sky130_fd_sc_hd__a21oi_4
X_42285_ _42284_/Y _42285_/Y sky130_fd_sc_hd__inv_2
X_77982_ _77983_/A _77983_/C _77983_/B _77984_/A sky130_fd_sc_hd__a21o_4
X_48901_ _48901_/A _48901_/B _48901_/Y sky130_fd_sc_hd__nand2_4
X_44024_ _44024_/A _64629_/A _57736_/A _58834_/A _44025_/A sky130_fd_sc_hd__and4_4
X_79721_ _84218_/Q _83266_/Q _79721_/X sky130_fd_sc_hd__xor2_4
X_41236_ _41235_/X _41236_/X sky130_fd_sc_hd__buf_2
X_60070_ _60069_/Y _60070_/Y sky130_fd_sc_hd__inv_2
X_72056_ _72054_/Y _72033_/X _72055_/Y _83294_/D sky130_fd_sc_hd__a21boi_4
X_76933_ _76918_/B _76933_/Y sky130_fd_sc_hd__inv_2
X_49881_ _49854_/A _49901_/A sky130_fd_sc_hd__buf_2
X_71007_ _51350_/B _70983_/A _71006_/Y _71007_/Y sky130_fd_sc_hd__o21ai_4
X_48832_ _86474_/Q _48809_/X _48831_/Y _48832_/Y sky130_fd_sc_hd__o21ai_4
X_79652_ _79652_/A _79638_/Y _79652_/X sky130_fd_sc_hd__or2_4
X_41167_ _81718_/Q _41145_/B _41167_/X sky130_fd_sc_hd__or2_4
X_76864_ _81674_/Q _76864_/B _81370_/D sky130_fd_sc_hd__xor2_4
Xclkbuf_10_473_0_CLK clkbuf_9_236_0_CLK/X _83666_/CLK sky130_fd_sc_hd__clkbuf_1
X_78603_ _78591_/A _78602_/Y _78575_/B _78603_/Y sky130_fd_sc_hd__o21ai_4
X_75815_ _75815_/A _75815_/Y sky130_fd_sc_hd__inv_2
X_48763_ _48777_/A _48763_/B _48763_/Y sky130_fd_sc_hd__nand2_4
X_79583_ _84206_/Q _83254_/Q _79584_/A sky130_fd_sc_hd__or2_4
X_45975_ _43605_/A _45975_/X sky130_fd_sc_hd__buf_2
X_41098_ _41098_/A _41098_/X sky130_fd_sc_hd__buf_2
X_76795_ _76781_/Y _76794_/X _76795_/Y sky130_fd_sc_hd__nand2_4
X_47714_ _47714_/A _47714_/X sky130_fd_sc_hd__buf_2
X_78534_ _82802_/Q _78534_/Y sky130_fd_sc_hd__inv_2
X_44926_ _45237_/A _44926_/X sky130_fd_sc_hd__buf_2
X_63760_ _61744_/X _63738_/B _63738_/C _63738_/D _63760_/Y sky130_fd_sc_hd__nand4_4
X_75746_ _75734_/A _75733_/Y _75745_/X _75747_/B sky130_fd_sc_hd__o21ai_4
X_48694_ _48694_/A _48695_/B sky130_fd_sc_hd__buf_2
X_72958_ _72806_/X _86202_/Q _72955_/X _72957_/X _72958_/X sky130_fd_sc_hd__a211o_4
X_60972_ _60921_/X _60934_/X _63781_/C _60972_/X sky130_fd_sc_hd__and3_4
X_62711_ _62711_/A _64276_/C _62676_/C _62657_/X _62711_/X sky130_fd_sc_hd__and4_4
X_47645_ _47655_/A _47645_/B _47614_/X _53165_/D _47645_/X sky130_fd_sc_hd__and4_4
X_71909_ _56645_/Y _71891_/Y _71908_/Y _71909_/Y sky130_fd_sc_hd__o21ai_4
X_78465_ _78465_/A _78464_/X _78475_/A sky130_fd_sc_hd__xor2_4
X_44857_ _45980_/A _44857_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_488_0_CLK clkbuf_9_244_0_CLK/X _86600_/CLK sky130_fd_sc_hd__clkbuf_1
X_63691_ _63849_/A _63701_/B sky130_fd_sc_hd__buf_2
X_75677_ _81118_/Q _75677_/B _75677_/Y sky130_fd_sc_hd__xnor2_4
X_72889_ _73351_/A _72889_/X sky130_fd_sc_hd__buf_2
X_65430_ _65428_/X _83081_/Q _65407_/X _65429_/X _65431_/B sky130_fd_sc_hd__a211o_4
X_77416_ _77416_/A _77415_/X _77416_/X sky130_fd_sc_hd__xor2_4
X_43808_ _43808_/A _87257_/D sky130_fd_sc_hd__inv_2
X_62642_ _60325_/B _62642_/B _62642_/Y sky130_fd_sc_hd__nand2_4
X_74628_ _74627_/Y _74675_/A sky130_fd_sc_hd__buf_2
X_47576_ _47530_/A _47595_/A sky130_fd_sc_hd__buf_2
X_78396_ _78395_/X _78400_/A sky130_fd_sc_hd__buf_2
X_44788_ _44803_/A _44788_/X sky130_fd_sc_hd__buf_2
X_49315_ _86411_/Q _49300_/X _49314_/Y _49315_/Y sky130_fd_sc_hd__o21ai_4
X_46527_ _47972_/A _46527_/X sky130_fd_sc_hd__buf_2
X_65361_ _65334_/X _86116_/Q _65256_/X _65360_/X _65361_/X sky130_fd_sc_hd__a211o_4
X_77347_ _77334_/Y _77316_/B _77316_/A _77347_/Y sky130_fd_sc_hd__nand3_4
X_43739_ _51337_/A _48759_/A sky130_fd_sc_hd__buf_2
X_74559_ _56863_/X _74559_/X sky130_fd_sc_hd__buf_2
X_62573_ _62565_/X _62569_/Y _62571_/X _84872_/Q _62572_/X _62573_/Y
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_10_411_0_CLK clkbuf_9_205_0_CLK/X _83520_/CLK sky130_fd_sc_hd__clkbuf_1
X_67100_ _67028_/A _67100_/B _67100_/X sky130_fd_sc_hd__and2_4
X_64312_ _64301_/Y _64311_/X _64269_/X _64312_/X sky130_fd_sc_hd__o21a_4
X_49246_ _86425_/Q _49222_/X _49245_/Y _49246_/Y sky130_fd_sc_hd__o21ai_4
X_61524_ _61482_/A _61522_/X _61541_/C _61524_/Y sky130_fd_sc_hd__nand3_4
X_68080_ _68405_/A _86912_/Q _68080_/X sky130_fd_sc_hd__and2_4
X_46458_ _86735_/Q _46430_/X _46457_/Y _46458_/Y sky130_fd_sc_hd__o21ai_4
X_65292_ _64915_/X _65281_/Y _65291_/Y _65292_/Y sky130_fd_sc_hd__o21ai_4
X_77278_ _77279_/A _82086_/D _77278_/X sky130_fd_sc_hd__or2_4
X_67031_ _66910_/A _67031_/X sky130_fd_sc_hd__buf_2
X_79017_ _82648_/Q _82520_/D _79016_/Y _79017_/Y sky130_fd_sc_hd__a21oi_4
X_45409_ _45409_/A _44892_/X _45409_/Y sky130_fd_sc_hd__nor2_4
X_64243_ _64243_/A _64273_/A sky130_fd_sc_hd__buf_2
X_76229_ _76233_/C _76229_/Y sky130_fd_sc_hd__inv_2
X_61455_ _61394_/A _61455_/X sky130_fd_sc_hd__buf_2
X_49177_ _49156_/X _50712_/B _49177_/Y sky130_fd_sc_hd__nand2_4
X_46389_ _46389_/A _46380_/B _46389_/X sky130_fd_sc_hd__or2_4
X_60406_ _60636_/B _60406_/B _60512_/A _60406_/X sky130_fd_sc_hd__and3_4
X_48128_ _48138_/A _48337_/A _48128_/X sky130_fd_sc_hd__and2_4
X_64174_ _64170_/X _63741_/X _64171_/Y _64172_/Y _64173_/X _64174_/X
+ sky130_fd_sc_hd__a41o_4
X_61386_ _61375_/A _61386_/B _61375_/C _61386_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_10_426_0_CLK clkbuf_9_213_0_CLK/X _82792_/CLK sky130_fd_sc_hd__clkbuf_1
X_63125_ _63020_/A _63125_/X sky130_fd_sc_hd__buf_2
X_48059_ _48054_/Y _48055_/X _48058_/X _86572_/D sky130_fd_sc_hd__a21oi_4
X_60337_ _60337_/A _60284_/A _60337_/C _60337_/D _60337_/Y sky130_fd_sc_hd__nand4_4
X_68982_ _68978_/X _68981_/X _68773_/X _68982_/X sky130_fd_sc_hd__a21o_4
X_51070_ _86079_/Q _51047_/X _51069_/Y _51070_/Y sky130_fd_sc_hd__o21ai_4
X_67933_ _87142_/Q _67906_/X _67908_/X _67932_/X _67933_/X sky130_fd_sc_hd__a211o_4
X_63056_ _63231_/A _63056_/X sky130_fd_sc_hd__buf_2
X_79919_ _58108_/A _84172_/Q _79919_/Y sky130_fd_sc_hd__nand2_4
X_60268_ _60268_/A _60267_/X _60268_/C _60268_/Y sky130_fd_sc_hd__nand3_4
X_50021_ _50025_/A _50040_/B _50025_/C _53234_/D _50021_/X sky130_fd_sc_hd__and4_4
X_62007_ _61842_/A _62007_/X sky130_fd_sc_hd__buf_2
X_82930_ _82925_/CLK _78247_/X _82930_/Q sky130_fd_sc_hd__dfxtp_4
X_67864_ _66673_/X _68651_/A sky130_fd_sc_hd__buf_2
X_60199_ _60168_/A _60199_/X sky130_fd_sc_hd__buf_2
X_69603_ _64732_/A _69603_/X sky130_fd_sc_hd__buf_2
X_66815_ _66815_/A _66814_/X _66815_/Y sky130_fd_sc_hd__nand2_4
X_82861_ _82859_/CLK _78154_/B _82861_/Q sky130_fd_sc_hd__dfxtp_4
X_67795_ _68451_/A _67891_/A sky130_fd_sc_hd__buf_2
X_84600_ _84606_/CLK _60561_/Y _79140_/A sky130_fd_sc_hd__dfxtp_4
X_81812_ _81811_/CLK _81620_/Q _81812_/Q sky130_fd_sc_hd__dfxtp_4
X_69534_ _87510_/Q _69468_/X _69343_/X _69533_/X _69534_/X sky130_fd_sc_hd__a211o_4
X_54760_ _85383_/Q _54757_/X _54759_/Y _54760_/Y sky130_fd_sc_hd__o21ai_4
X_66746_ _87948_/Q _66697_/X _66675_/X _66745_/X _66746_/X sky130_fd_sc_hd__a211o_4
X_85580_ _83572_/CLK _53727_/Y _85580_/Q sky130_fd_sc_hd__dfxtp_4
X_51972_ _51265_/A _51972_/X sky130_fd_sc_hd__buf_2
X_63958_ _63942_/A _59411_/A _63958_/C _63958_/X sky130_fd_sc_hd__and3_4
X_82792_ _82792_/CLK _82824_/Q _82792_/Q sky130_fd_sc_hd__dfxtp_4
X_53711_ _52194_/A _53720_/B _53734_/C _53711_/X sky130_fd_sc_hd__and3_4
X_84531_ _84531_/CLK _84531_/D _84531_/Q sky130_fd_sc_hd__dfxtp_4
X_50923_ _50952_/A _50948_/C sky130_fd_sc_hd__buf_2
X_62909_ _61593_/B _62858_/X _62859_/X _62908_/X _62909_/Y sky130_fd_sc_hd__nand4_4
X_81743_ _88175_/CLK _81743_/D _81743_/Q sky130_fd_sc_hd__dfxtp_4
X_69465_ _68617_/A _69465_/X sky130_fd_sc_hd__buf_2
X_54691_ _54682_/A _47352_/A _54691_/Y sky130_fd_sc_hd__nand2_4
X_66677_ _87887_/Q _66562_/X _66675_/X _66676_/X _66677_/X sky130_fd_sc_hd__a211o_4
X_63889_ _63883_/Y _63884_/Y _63885_/Y _63888_/Y _63889_/X sky130_fd_sc_hd__and4_4
X_56430_ _56114_/X _56426_/X _56429_/Y _56430_/Y sky130_fd_sc_hd__o21ai_4
X_68416_ _44149_/A _68415_/Y _68416_/Y sky130_fd_sc_hd__nor2_4
X_87250_ _87260_/CLK _43822_/X _87250_/Q sky130_fd_sc_hd__dfxtp_4
X_53642_ _53639_/Y _53603_/X _53641_/Y _53642_/Y sky130_fd_sc_hd__a21boi_4
X_65628_ _65625_/X _65627_/X _65566_/X _65628_/X sky130_fd_sc_hd__a21o_4
X_84462_ _82436_/CLK _84462_/D _79130_/B sky130_fd_sc_hd__dfxtp_4
X_50854_ _50845_/A _50854_/B _50854_/Y sky130_fd_sc_hd__nand2_4
X_81674_ _81671_/CLK _81674_/D _81674_/Q sky130_fd_sc_hd__dfxtp_4
X_69396_ _66540_/A _69396_/X sky130_fd_sc_hd__buf_2
X_86201_ _86490_/CLK _86201_/D _86201_/Q sky130_fd_sc_hd__dfxtp_4
X_83413_ _83761_/CLK _71681_/Y _83413_/Q sky130_fd_sc_hd__dfxtp_4
X_56361_ _56159_/X _56350_/X _56360_/Y _85221_/D sky130_fd_sc_hd__o21ai_4
X_80625_ _80625_/A _63365_/C _80625_/X sky130_fd_sc_hd__xor2_4
X_68347_ _68347_/A _68517_/A sky130_fd_sc_hd__buf_2
X_87181_ _87169_/CLK _44215_/X _44067_/B sky130_fd_sc_hd__dfxtp_4
X_53573_ _85610_/Q _53540_/X _53572_/Y _53573_/Y sky130_fd_sc_hd__o21ai_4
X_65559_ _65559_/A _65559_/B _65559_/C _65559_/X sky130_fd_sc_hd__and3_4
X_84393_ _84393_/CLK _62654_/Y _75923_/B sky130_fd_sc_hd__dfxtp_4
X_50785_ _50777_/A _49265_/B _50785_/Y sky130_fd_sc_hd__nand2_4
X_58100_ _58605_/A _58100_/X sky130_fd_sc_hd__buf_2
X_55312_ _44095_/X _55312_/X sky130_fd_sc_hd__buf_2
X_86132_ _85527_/CLK _86132_/D _86132_/Q sky130_fd_sc_hd__dfxtp_4
X_52524_ _52524_/A _52509_/B _52498_/C _52524_/X sky130_fd_sc_hd__and3_4
X_59080_ _64776_/A _59081_/A sky130_fd_sc_hd__buf_2
X_83344_ _83491_/CLK _71877_/X _83344_/Q sky130_fd_sc_hd__dfxtp_4
X_56292_ _56005_/X _56290_/X _56291_/Y _85248_/D sky130_fd_sc_hd__o21ai_4
X_80556_ _80547_/X _80549_/B _80556_/Y sky130_fd_sc_hd__nand2_4
X_68278_ _83994_/Q _68259_/X _68277_/X _68278_/X sky130_fd_sc_hd__a21bo_4
X_58031_ _58030_/X _85483_/Q _57962_/X _58031_/X sky130_fd_sc_hd__o21a_4
X_55243_ _55243_/A _55243_/B _56889_/B _55288_/B sky130_fd_sc_hd__nand3_4
X_67229_ _67224_/X _67228_/X _67204_/X _67229_/X sky130_fd_sc_hd__a21o_4
X_86063_ _85745_/CLK _51161_/Y _86063_/Q sky130_fd_sc_hd__dfxtp_4
X_52455_ _52453_/Y _52430_/X _52454_/Y _52455_/Y sky130_fd_sc_hd__a21boi_4
X_83275_ _83275_/CLK _83275_/D _83275_/Q sky130_fd_sc_hd__dfxtp_4
X_80487_ _80487_/A _80487_/Y sky130_fd_sc_hd__inv_2
X_85014_ _85049_/CLK _57403_/X _85014_/Q sky130_fd_sc_hd__dfxtp_4
X_51406_ _51220_/A _51230_/X _51225_/C _52934_/D _51406_/X sky130_fd_sc_hd__and4_4
X_70240_ _70238_/X _83826_/Q _70239_/X _83826_/D sky130_fd_sc_hd__a21o_4
X_82226_ _81094_/CLK _82258_/Q _77455_/A sky130_fd_sc_hd__dfxtp_4
X_55174_ _55244_/A _55174_/X sky130_fd_sc_hd__buf_2
X_52386_ _52384_/Y _52364_/X _52385_/X _52386_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_8_53_0_CLK clkbuf_8_53_0_CLK/A clkbuf_8_53_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_54125_ _54134_/A _54125_/B _54125_/Y sky130_fd_sc_hd__nand2_4
X_51337_ _51337_/A _51822_/A sky130_fd_sc_hd__buf_2
X_70171_ _70231_/A _70183_/A sky130_fd_sc_hd__buf_2
X_82157_ _84175_/CLK _80419_/B _82157_/Q sky130_fd_sc_hd__dfxtp_4
X_59982_ _59873_/A _59873_/B _59982_/C _59982_/Y sky130_fd_sc_hd__nor3_4
X_81108_ _81087_/CLK _79751_/X _75889_/A sky130_fd_sc_hd__dfxtp_4
X_42070_ _42052_/X _42043_/X _40959_/X _88047_/Q _42044_/X _42071_/A
+ sky130_fd_sc_hd__o32ai_4
X_54056_ _54031_/A _49322_/B _54056_/Y sky130_fd_sc_hd__nand2_4
X_58933_ _84788_/Q _79180_/A sky130_fd_sc_hd__inv_2
X_51268_ _51280_/A _50757_/B _51268_/Y sky130_fd_sc_hd__nand2_4
X_86965_ _86965_/CLK _44770_/Y _86965_/Q sky130_fd_sc_hd__dfxtp_4
X_82088_ _81970_/CLK _82132_/Q _82088_/Q sky130_fd_sc_hd__dfxtp_4
X_41021_ _41021_/A _41021_/X sky130_fd_sc_hd__buf_2
X_53007_ _53062_/A _53019_/C sky130_fd_sc_hd__buf_2
X_50219_ _50655_/A _50219_/X sky130_fd_sc_hd__buf_2
X_73930_ _72894_/X _73930_/X sky130_fd_sc_hd__buf_2
X_85916_ _86560_/CLK _85916_/D _65972_/B sky130_fd_sc_hd__dfxtp_4
X_81039_ _81038_/CLK _81039_/D _81039_/Q sky130_fd_sc_hd__dfxtp_4
X_58864_ _58864_/A _58864_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_68_0_CLK clkbuf_8_69_0_CLK/A clkbuf_8_68_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_51199_ _51184_/X _52889_/B _51199_/Y sky130_fd_sc_hd__nand2_4
X_86896_ _86896_/CLK _45146_/Y _64392_/B sky130_fd_sc_hd__dfxtp_4
X_57815_ _57739_/X _85724_/Q _57814_/X _57815_/X sky130_fd_sc_hd__o21a_4
X_73861_ _73954_/A _66087_/B _73861_/X sky130_fd_sc_hd__and2_4
X_85847_ _83303_/CLK _52316_/Y _85847_/Q sky130_fd_sc_hd__dfxtp_4
X_58795_ _58740_/X _85455_/Q _58794_/X _58795_/Y sky130_fd_sc_hd__o21ai_4
X_75600_ _75607_/B _75891_/A _75600_/X sky130_fd_sc_hd__xor2_4
X_72812_ _73067_/A _72812_/X sky130_fd_sc_hd__buf_2
X_45760_ _82986_/Q _45761_/A sky130_fd_sc_hd__inv_2
X_57746_ _46213_/X _57744_/Y _57745_/Y _57700_/X _57703_/X _57746_/X
+ sky130_fd_sc_hd__o32a_4
X_76580_ _76576_/X _76577_/Y _76579_/Y _76614_/A sky130_fd_sc_hd__a21o_4
X_42972_ _42970_/X _42971_/X _40432_/X _87624_/Q _42954_/X _42972_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54958_ _85345_/Q _54249_/X _54957_/Y _54958_/Y sky130_fd_sc_hd__o21ai_4
X_73792_ _73790_/X _73792_/B _73779_/Y _73792_/Y sky130_fd_sc_hd__nand3_4
X_85778_ _85778_/CLK _52662_/Y _85778_/Q sky130_fd_sc_hd__dfxtp_4
X_44711_ _44707_/X _44708_/X _40678_/A _44709_/Y _44710_/X _86991_/D
+ sky130_fd_sc_hd__o32ai_4
X_75531_ _75528_/B _75528_/A _75531_/Y sky130_fd_sc_hd__nand2_4
X_87517_ _87767_/CLK _87517_/D _87517_/Q sky130_fd_sc_hd__dfxtp_4
X_41923_ _41887_/X _41919_/X _40650_/X _41922_/Y _41891_/X _88104_/D
+ sky130_fd_sc_hd__o32ai_4
X_53909_ _85544_/Q _53896_/X _53908_/Y _53909_/Y sky130_fd_sc_hd__o21ai_4
X_72743_ _44514_/Y _56275_/X _72742_/Y _72764_/C sky130_fd_sc_hd__a21o_4
X_84729_ _83402_/CLK _59452_/X _84729_/Q sky130_fd_sc_hd__dfxtp_4
X_45691_ _45265_/A _45691_/X sky130_fd_sc_hd__buf_2
X_57677_ _57650_/A _57677_/X sky130_fd_sc_hd__buf_2
X_54889_ _54889_/A _54910_/C sky130_fd_sc_hd__buf_2
X_47430_ _47525_/A _47444_/A sky130_fd_sc_hd__buf_2
X_59416_ _59394_/X _83483_/Q _59415_/Y _84739_/D sky130_fd_sc_hd__o21a_4
X_78250_ _78250_/A _78250_/Y sky130_fd_sc_hd__inv_2
X_56628_ _56626_/X _56553_/Y _56627_/Y _56628_/Y sky130_fd_sc_hd__a21oi_4
X_44642_ _44642_/A _87021_/D sky130_fd_sc_hd__inv_2
X_75462_ _75458_/X _75509_/C _75509_/A _75462_/X sky130_fd_sc_hd__a21o_4
X_87448_ _87221_/CLK _43385_/X _87448_/Q sky130_fd_sc_hd__dfxtp_4
X_41854_ _40528_/X _41847_/X _67218_/B _41848_/X _88120_/D sky130_fd_sc_hd__a2bb2o_4
X_72674_ _72688_/A _72683_/B sky130_fd_sc_hd__buf_2
X_77201_ _77202_/A _77184_/X _77202_/B _77202_/C _77201_/Y sky130_fd_sc_hd__nand4_4
X_74413_ _46280_/A _74413_/X sky130_fd_sc_hd__buf_2
X_40805_ _40773_/X _82297_/Q _40804_/X _40806_/A sky130_fd_sc_hd__o21ai_4
X_47361_ _47333_/X _53005_/B _47361_/Y sky130_fd_sc_hd__nand2_4
X_59347_ _59346_/X _85637_/Q _59308_/X _59347_/X sky130_fd_sc_hd__o21a_4
X_71625_ _71628_/A _71625_/Y sky130_fd_sc_hd__inv_2
X_78181_ _78191_/A _78192_/A _78182_/B sky130_fd_sc_hd__xor2_4
X_44573_ _44573_/A _44573_/Y sky130_fd_sc_hd__inv_2
X_56559_ _55624_/X _56564_/B sky130_fd_sc_hd__buf_2
X_75393_ _75393_/A _75393_/B _75393_/Y sky130_fd_sc_hd__nor2_4
X_41785_ _40385_/B _82883_/Q _41784_/X _41785_/X sky130_fd_sc_hd__o21a_4
X_87379_ _87993_/CLK _43521_/X _87379_/Q sky130_fd_sc_hd__dfxtp_4
X_49100_ _48499_/A _71959_/A sky130_fd_sc_hd__buf_2
X_46312_ _46297_/Y _46300_/X _46311_/X _86749_/D sky130_fd_sc_hd__a21oi_4
X_77132_ _82100_/Q _77132_/B _77132_/X sky130_fd_sc_hd__xor2_4
X_43524_ _43518_/X _43523_/X _40371_/X _87377_/Q _43506_/X _43524_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74344_ _70328_/C _74340_/X _74343_/Y _83091_/D sky130_fd_sc_hd__a21bo_4
X_40736_ _40736_/A _40765_/B sky130_fd_sc_hd__buf_2
X_59278_ _59053_/A _59278_/X sky130_fd_sc_hd__buf_2
X_47292_ _47198_/X _47330_/A sky130_fd_sc_hd__buf_2
X_71556_ _71556_/A _71556_/Y sky130_fd_sc_hd__inv_2
X_49031_ _49031_/A _53854_/B sky130_fd_sc_hd__buf_2
X_46243_ _46290_/A _46623_/A sky130_fd_sc_hd__buf_2
X_70507_ _71170_/A _70966_/A sky130_fd_sc_hd__buf_2
X_58229_ _58229_/A _58229_/Y sky130_fd_sc_hd__inv_2
XPHY_550 sky130_fd_sc_hd__decap_3
X_77063_ _77068_/A _77067_/A _77062_/Y _77063_/Y sky130_fd_sc_hd__a21boi_4
X_43455_ _43020_/A _43528_/A sky130_fd_sc_hd__buf_2
X_74275_ _74272_/X _74274_/X _74019_/X _74278_/A sky130_fd_sc_hd__a21o_4
XPHY_561 sky130_fd_sc_hd__decap_3
X_40667_ _40667_/A _40667_/X sky130_fd_sc_hd__buf_2
X_71487_ _71487_/A _71487_/X sky130_fd_sc_hd__buf_2
XPHY_572 sky130_fd_sc_hd__decap_3
XPHY_583 sky130_fd_sc_hd__decap_3
X_76014_ _76009_/Y _76010_/A _76013_/Y _76015_/B sky130_fd_sc_hd__a21boi_4
X_42406_ _42401_/X _42397_/X _40446_/X _87878_/Q _42398_/X _42407_/A
+ sky130_fd_sc_hd__o32ai_4
XPHY_594 sky130_fd_sc_hd__decap_3
X_61240_ _61198_/X _61107_/X _61230_/C _61241_/A sky130_fd_sc_hd__nand3_4
X_73226_ _69804_/Y _73224_/X _73194_/X _73225_/Y _73226_/X sky130_fd_sc_hd__a211o_4
X_46174_ _46162_/X _46173_/X _46166_/C _46174_/X sky130_fd_sc_hd__and3_4
X_70438_ _70442_/A _70947_/B _70431_/C _70438_/Y sky130_fd_sc_hd__nand3_4
X_43386_ _43396_/A _43386_/X sky130_fd_sc_hd__buf_2
X_40598_ _40755_/A _40599_/A sky130_fd_sc_hd__buf_2
X_45125_ _44972_/X _45125_/X sky130_fd_sc_hd__buf_2
X_42337_ _42337_/A _87915_/D sky130_fd_sc_hd__inv_2
X_61171_ _64250_/C _64211_/C sky130_fd_sc_hd__buf_2
X_73157_ _72757_/A _73495_/A sky130_fd_sc_hd__buf_2
X_70369_ _70361_/Y _70370_/A sky130_fd_sc_hd__buf_2
X_60122_ _60122_/A _60267_/A _60122_/C _60122_/Y sky130_fd_sc_hd__nand3_4
X_72108_ _74391_/A _50719_/B _72108_/Y sky130_fd_sc_hd__nand2_4
X_49933_ _49929_/Y _49924_/X _49932_/X _49933_/Y sky130_fd_sc_hd__a21oi_4
X_45056_ _45197_/A _45056_/X sky130_fd_sc_hd__buf_2
X_42268_ _42252_/X _42243_/X _41498_/X _87948_/Q _42244_/X _42269_/A
+ sky130_fd_sc_hd__o32ai_4
X_77965_ _77965_/A _77967_/B sky130_fd_sc_hd__inv_2
X_73088_ _69725_/B _73086_/X _73087_/X _73088_/X sky130_fd_sc_hd__o21a_4
X_44007_ HASH_EN _44010_/A sky130_fd_sc_hd__buf_2
X_79704_ _79704_/A _79704_/B _79704_/X sky130_fd_sc_hd__and2_4
X_41219_ _41042_/X _81709_/Q _41218_/X _41219_/X sky130_fd_sc_hd__o21a_4
X_64930_ _64817_/X _86165_/Q _64927_/X _64929_/X _64930_/X sky130_fd_sc_hd__a211o_4
X_60053_ _72584_/C _60053_/X sky130_fd_sc_hd__buf_2
X_72039_ _72037_/Y _72033_/X _72038_/Y _72039_/Y sky130_fd_sc_hd__a21boi_4
X_76916_ _81503_/Q _76918_/A sky130_fd_sc_hd__inv_2
X_49864_ _49864_/A _53076_/B _49864_/Y sky130_fd_sc_hd__nand2_4
X_42199_ _41878_/A _42199_/X sky130_fd_sc_hd__buf_2
X_77896_ _77880_/B _77893_/X _77895_/Y _77902_/B sky130_fd_sc_hd__a21oi_4
Xclkbuf_3_7_1_CLK clkbuf_3_7_0_CLK/X clkbuf_3_7_1_CLK/X sky130_fd_sc_hd__clkbuf_1
X_48815_ _48812_/Y _48813_/X _48814_/X _48815_/Y sky130_fd_sc_hd__a21oi_4
X_79635_ _79630_/A _79629_/X _79634_/Y _79652_/A sky130_fd_sc_hd__a21boi_4
X_64861_ _64858_/X _85528_/Q _64859_/X _64860_/X _64861_/X sky130_fd_sc_hd__a211o_4
X_76847_ _76847_/A _76847_/B _76847_/Y sky130_fd_sc_hd__xnor2_4
X_49795_ _49794_/X _49795_/X sky130_fd_sc_hd__buf_2
X_66600_ _66553_/X _68721_/A sky130_fd_sc_hd__buf_2
X_63812_ _61796_/X _63860_/B _63738_/C _63860_/D _63812_/Y sky130_fd_sc_hd__nand4_4
X_48746_ _48737_/A _48435_/B _48746_/Y sky130_fd_sc_hd__nand2_4
X_67580_ _87977_/Q _67533_/X _67508_/X _67579_/X _67580_/X sky130_fd_sc_hd__a211o_4
X_79566_ _79566_/A _79566_/B _79569_/A sky130_fd_sc_hd__nand2_4
X_45958_ _44216_/X _44217_/X _44153_/X _45950_/B _45958_/X sky130_fd_sc_hd__a211o_4
X_64792_ _64767_/A _85818_/Q _64792_/X sky130_fd_sc_hd__and2_4
X_76778_ _76755_/Y _81358_/D sky130_fd_sc_hd__inv_2
X_66531_ _69245_/A _66531_/X sky130_fd_sc_hd__buf_2
X_78517_ _78497_/X _78515_/Y _78516_/Y _78517_/Y sky130_fd_sc_hd__a21oi_4
X_44909_ _44890_/X _44902_/X _44908_/Y _44909_/Y sky130_fd_sc_hd__a21oi_4
X_63743_ _63732_/X _63736_/X _63738_/Y _63739_/Y _63742_/Y _63743_/X
+ sky130_fd_sc_hd__a41o_4
X_75729_ _75723_/B _75723_/A _75728_/Y _75730_/B sky130_fd_sc_hd__a21oi_4
X_60955_ _60915_/X _63972_/A sky130_fd_sc_hd__buf_2
X_48677_ _48652_/X _82341_/Q _48676_/Y _74501_/A sky130_fd_sc_hd__o21ai_4
X_79497_ _79489_/A _79488_/Y _79496_/X _79498_/B sky130_fd_sc_hd__o21ai_4
X_45889_ _45889_/A _45893_/B sky130_fd_sc_hd__buf_2
X_69250_ _87531_/Q _69044_/X _69248_/X _69249_/X _69250_/X sky130_fd_sc_hd__a211o_4
X_47628_ _55013_/D _53155_/D sky130_fd_sc_hd__buf_2
X_66462_ _65107_/X _66476_/B _65110_/X _66462_/Y sky130_fd_sc_hd__nand3_4
X_78448_ _78466_/A _78466_/B _78448_/X sky130_fd_sc_hd__xor2_4
X_63674_ _63696_/A _62140_/X _63674_/X sky130_fd_sc_hd__and2_4
X_60886_ _60996_/B _60901_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_350_0_CLK clkbuf_9_175_0_CLK/X _85651_/CLK sky130_fd_sc_hd__clkbuf_1
X_68201_ _67252_/X _67254_/X _68173_/X _68201_/Y sky130_fd_sc_hd__a21oi_4
X_65413_ _65285_/A _65413_/B _65413_/X sky130_fd_sc_hd__and2_4
X_62625_ _62618_/X _62622_/Y _62624_/X _84867_/Q _62212_/A _62625_/Y
+ sky130_fd_sc_hd__o32ai_4
X_69181_ _69177_/X _69180_/X _69025_/X _69181_/X sky130_fd_sc_hd__a21o_4
X_47559_ _47530_/X _47595_/B _47519_/X _53118_/D _47559_/X sky130_fd_sc_hd__and4_4
X_66393_ _66282_/X _65999_/Y _66392_/Y _66393_/Y sky130_fd_sc_hd__o21ai_4
X_78379_ _78379_/A _78380_/B sky130_fd_sc_hd__inv_2
Xclkbuf_10_980_0_CLK clkbuf_9_490_0_CLK/X _85557_/CLK sky130_fd_sc_hd__clkbuf_1
X_80410_ _84756_/Q _84148_/Q _80410_/Y sky130_fd_sc_hd__nand2_4
X_68132_ _82071_/D _68120_/X _68131_/X _68132_/X sky130_fd_sc_hd__a21bo_4
X_65344_ _65342_/X _86725_/Q _65239_/X _65343_/X _65344_/X sky130_fd_sc_hd__a211o_4
X_50570_ _50575_/A _48901_/B _50570_/Y sky130_fd_sc_hd__nand2_4
X_62556_ _62556_/A _63280_/B _59977_/A _62548_/D _62556_/X sky130_fd_sc_hd__and4_4
X_81390_ _83926_/CLK _81390_/D _76907_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_471_0_CLK clkbuf_9_471_0_CLK/A clkbuf_9_471_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_61507_ _61518_/A _61518_/B _84475_/Q _61507_/Y sky130_fd_sc_hd__nor3_4
X_49229_ _64710_/B _49204_/X _49228_/Y _49229_/Y sky130_fd_sc_hd__o21ai_4
X_80341_ _80324_/A _80326_/X _80327_/Y _80341_/Y sky130_fd_sc_hd__a21boi_4
X_68063_ _68056_/X _68061_/X _68062_/X _68063_/Y sky130_fd_sc_hd__a21oi_4
X_65275_ _65403_/A _65275_/B _65275_/X sky130_fd_sc_hd__and2_4
X_62487_ _62269_/A _62487_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_365_0_CLK clkbuf_9_182_0_CLK/X _85704_/CLK sky130_fd_sc_hd__clkbuf_1
X_67014_ _67013_/X _67014_/X sky130_fd_sc_hd__buf_2
X_52240_ _52215_/A _52250_/A sky130_fd_sc_hd__buf_2
X_64226_ _64249_/A _64226_/X sky130_fd_sc_hd__buf_2
X_83060_ _83562_/CLK _83060_/D _83060_/Q sky130_fd_sc_hd__dfxtp_4
X_61438_ _84824_/Q _61438_/X sky130_fd_sc_hd__buf_2
X_80272_ _80636_/A _80270_/X _80271_/Y _80288_/A sky130_fd_sc_hd__a21boi_4
Xclkbuf_10_995_0_CLK clkbuf_9_497_0_CLK/X _85593_/CLK sky130_fd_sc_hd__clkbuf_1
X_82011_ _82139_/CLK _82043_/Q _82011_/Q sky130_fd_sc_hd__dfxtp_4
X_52171_ _50469_/A _52194_/B _52182_/C _52171_/X sky130_fd_sc_hd__and3_4
X_64157_ _64524_/B _64179_/B _64179_/C _64179_/D _64157_/Y sky130_fd_sc_hd__nand4_4
X_61369_ _61368_/Y _61369_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_9_486_0_CLK clkbuf_9_486_0_CLK/A clkbuf_9_486_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_51122_ _51118_/Y _51119_/X _51121_/X _51122_/Y sky130_fd_sc_hd__a21oi_4
X_63108_ _63097_/A _64320_/B _63108_/C _63085_/D _63108_/X sky130_fd_sc_hd__and4_4
X_68965_ _68987_/A _87739_/Q _68965_/X sky130_fd_sc_hd__and2_4
X_64088_ _64116_/A _64087_/X _64088_/C _64088_/Y sky130_fd_sc_hd__nor3_4
X_51053_ _51058_/A _46912_/X _51053_/Y sky130_fd_sc_hd__nand2_4
X_55930_ _56208_/C _55605_/X _44090_/B _55929_/X _55930_/X sky130_fd_sc_hd__a211o_4
X_67916_ _87387_/Q _67868_/X _67821_/X _67915_/X _67916_/X sky130_fd_sc_hd__a211o_4
X_63039_ _63039_/A _64248_/C _63028_/X _63014_/D _63039_/X sky130_fd_sc_hd__and4_4
X_86750_ _85822_/CLK _46289_/Y _86750_/Q sky130_fd_sc_hd__dfxtp_4
X_83962_ _80991_/CLK _83962_/D _80818_/D sky130_fd_sc_hd__dfxtp_4
X_68896_ _68779_/A _68896_/B _68896_/X sky130_fd_sc_hd__and2_4
X_50004_ _46308_/A _50025_/A sky130_fd_sc_hd__buf_2
X_85701_ _85700_/CLK _53079_/Y _85701_/Q sky130_fd_sc_hd__dfxtp_4
X_82913_ _81195_/CLK _78307_/X _82913_/Q sky130_fd_sc_hd__dfxtp_4
X_55861_ _45122_/A _55522_/X _55532_/X _55860_/X _55862_/B sky130_fd_sc_hd__a211o_4
X_86681_ _86361_/CLK _86681_/D _59094_/A sky130_fd_sc_hd__dfxtp_4
X_67847_ _67844_/X _67846_/X _67799_/X _67847_/X sky130_fd_sc_hd__a21o_4
X_83893_ _82299_/CLK _83893_/D _83893_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_303_0_CLK clkbuf_9_151_0_CLK/X _84321_/CLK sky130_fd_sc_hd__clkbuf_1
X_57600_ _84971_/Q _57562_/X _57599_/Y _57600_/Y sky130_fd_sc_hd__o21ai_4
X_54812_ _54892_/A _54812_/X sky130_fd_sc_hd__buf_2
X_85632_ _86592_/CLK _53459_/Y _85632_/Q sky130_fd_sc_hd__dfxtp_4
X_58580_ _58085_/X _85472_/Q _58579_/X _58580_/Y sky130_fd_sc_hd__o21ai_4
X_82844_ _82748_/CLK _82844_/D _82844_/Q sky130_fd_sc_hd__dfxtp_4
X_55792_ _55711_/X _85228_/Q _55792_/X sky130_fd_sc_hd__and2_4
X_67778_ _87149_/Q _67706_/X _67755_/X _67777_/X _67778_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_933_0_CLK clkbuf_9_466_0_CLK/X _87045_/CLK sky130_fd_sc_hd__clkbuf_1
X_57531_ _57531_/A _50275_/B _57531_/Y sky130_fd_sc_hd__nand2_4
X_69517_ _69036_/X _69038_/X _69500_/X _69517_/Y sky130_fd_sc_hd__a21oi_4
X_88351_ _87859_/CLK _40704_/Y _88351_/Q sky130_fd_sc_hd__dfxtp_4
X_54743_ _54748_/A _54755_/B _54748_/C _54743_/D _54743_/X sky130_fd_sc_hd__and4_4
X_66729_ _88397_/Q _66633_/X _66682_/X _66728_/X _66729_/X sky130_fd_sc_hd__a211o_4
X_85563_ _83310_/CLK _53815_/Y _85563_/Q sky130_fd_sc_hd__dfxtp_4
X_51955_ _85917_/Q _51945_/X _51954_/Y _51955_/Y sky130_fd_sc_hd__o21ai_4
X_82775_ _82965_/CLK _82775_/D _82967_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_424_0_CLK clkbuf_9_424_0_CLK/A clkbuf_9_424_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_87302_ _87553_/CLK _87302_/D _43703_/A sky130_fd_sc_hd__dfxtp_4
X_84514_ _84498_/CLK _84514_/D _61174_/C sky130_fd_sc_hd__dfxtp_4
X_50906_ _50906_/A _51770_/B _50906_/Y sky130_fd_sc_hd__nand2_4
X_57462_ _57461_/Y _85000_/D sky130_fd_sc_hd__inv_2
X_81726_ _84020_/CLK _81726_/D _81726_/Q sky130_fd_sc_hd__dfxtp_4
X_69448_ _69445_/X _69448_/B _69448_/Y sky130_fd_sc_hd__nand2_4
X_88282_ _87026_/CLK _41078_/Y _69486_/B sky130_fd_sc_hd__dfxtp_4
X_54674_ _54674_/A _54674_/B _54674_/C _47320_/A _54674_/X sky130_fd_sc_hd__and4_4
X_85494_ _85492_/CLK _85494_/D _85494_/Q sky130_fd_sc_hd__dfxtp_4
X_51886_ _51804_/A _51887_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_318_0_CLK clkbuf_9_159_0_CLK/X _85381_/CLK sky130_fd_sc_hd__clkbuf_1
X_59201_ _59177_/X _86065_/Q _59200_/X _59201_/Y sky130_fd_sc_hd__o21ai_4
X_56413_ _56074_/X _56409_/X _56412_/Y _85204_/D sky130_fd_sc_hd__o21ai_4
X_87233_ _87748_/CLK _87233_/D _68815_/B sky130_fd_sc_hd__dfxtp_4
X_53625_ _53623_/Y _53619_/X _53624_/X _53625_/Y sky130_fd_sc_hd__a21oi_4
X_84445_ _84452_/CLK _84445_/D _78068_/B sky130_fd_sc_hd__dfxtp_4
X_50837_ _86123_/Q _50820_/X _50836_/Y _50837_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_948_0_CLK clkbuf_9_474_0_CLK/X _84970_/CLK sky130_fd_sc_hd__clkbuf_1
X_57393_ _56600_/X _57391_/Y _57392_/Y _57393_/Y sky130_fd_sc_hd__a21oi_4
X_81657_ _81697_/CLK _76707_/A _81657_/Q sky130_fd_sc_hd__dfxtp_4
X_69379_ _69329_/X _68798_/Y _69325_/X _69378_/Y _69379_/X sky130_fd_sc_hd__a211o_4
X_59132_ _58602_/A _59133_/A sky130_fd_sc_hd__buf_2
X_71410_ _71397_/X _83509_/Q _71409_/Y _83509_/D sky130_fd_sc_hd__a21o_4
X_56344_ _56121_/X _56337_/X _56343_/Y _56344_/Y sky130_fd_sc_hd__o21ai_4
X_80608_ _80608_/A _80608_/B _80608_/X sky130_fd_sc_hd__or2_4
X_87164_ _86941_/CLK _87164_/D _87164_/Q sky130_fd_sc_hd__dfxtp_4
X_41570_ _41569_/Y _41570_/X sky130_fd_sc_hd__buf_2
X_53556_ _53687_/A _53556_/X sky130_fd_sc_hd__buf_2
X_72390_ _72389_/X _85675_/Q _72308_/X _72390_/X sky130_fd_sc_hd__o21a_4
X_84376_ _84507_/CLK _84376_/D _62864_/C sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_439_0_CLK clkbuf_9_438_0_CLK/A clkbuf_9_439_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_50768_ _50768_/A _50768_/X sky130_fd_sc_hd__buf_2
X_81588_ _84087_/CLK _84188_/Q _76819_/A sky130_fd_sc_hd__dfxtp_4
X_86115_ _86736_/CLK _50877_/Y _86115_/Q sky130_fd_sc_hd__dfxtp_4
X_40521_ _40520_/X _40508_/X _88378_/Q _40510_/X _40521_/X sky130_fd_sc_hd__a2bb2o_4
X_52507_ _65049_/B _52422_/X _52506_/Y _52507_/Y sky130_fd_sc_hd__o21ai_4
X_59063_ _59061_/X _86076_/Q _59062_/X _59063_/Y sky130_fd_sc_hd__o21ai_4
X_71341_ _71485_/B _71342_/B sky130_fd_sc_hd__buf_2
X_83327_ _83333_/CLK _83327_/D _83327_/Q sky130_fd_sc_hd__dfxtp_4
X_56275_ _56274_/X _56275_/X sky130_fd_sc_hd__buf_2
X_80539_ _80539_/A _84321_/Q _80540_/B sky130_fd_sc_hd__xor2_4
X_87095_ _88267_/CLK _87095_/D _87095_/Q sky130_fd_sc_hd__dfxtp_4
X_53487_ _85627_/Q _53476_/X _53486_/Y _53487_/Y sky130_fd_sc_hd__o21ai_4
X_50699_ _50577_/A _50699_/X sky130_fd_sc_hd__buf_2
X_58014_ _58635_/A _58701_/A sky130_fd_sc_hd__buf_2
X_43240_ _41032_/X _43216_/X _87522_/Q _43218_/X _87522_/D sky130_fd_sc_hd__a2bb2o_4
X_55226_ _55227_/A _55225_/X _83315_/Q _55226_/Y sky130_fd_sc_hd__a21oi_4
X_74060_ _73972_/X _66211_/B _74060_/X sky130_fd_sc_hd__and2_4
X_86046_ _85535_/CLK _51252_/Y _64670_/B sky130_fd_sc_hd__dfxtp_4
X_40452_ _40451_/X _40452_/X sky130_fd_sc_hd__buf_2
X_52438_ _52438_/A _52438_/X sky130_fd_sc_hd__buf_2
X_71272_ _53187_/B _71265_/X _71271_/Y _83552_/D sky130_fd_sc_hd__o21ai_4
X_83258_ _81227_/CLK _83258_/D _72394_/A sky130_fd_sc_hd__dfxtp_4
X_73011_ _72806_/X _86200_/Q _72955_/X _73010_/X _73011_/X sky130_fd_sc_hd__a211o_4
X_70223_ _70337_/A _70238_/A sky130_fd_sc_hd__buf_2
X_82209_ _82965_/CLK _82209_/D _82209_/Q sky130_fd_sc_hd__dfxtp_4
X_43171_ _43046_/X _43125_/X _40881_/X _43170_/Y _43142_/X _43171_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55157_ _44058_/A _55157_/X sky130_fd_sc_hd__buf_2
X_40383_ _40586_/A _46317_/A sky130_fd_sc_hd__buf_2
X_52369_ _52247_/A _52369_/X sky130_fd_sc_hd__buf_2
X_83189_ _83188_/CLK _83189_/D _70229_/C sky130_fd_sc_hd__dfxtp_4
X_42122_ _42122_/A _88025_/D sky130_fd_sc_hd__inv_2
X_54108_ _43013_/X _54245_/A sky130_fd_sc_hd__buf_2
X_70154_ _70154_/A _70144_/X _70149_/X _70153_/Y _70154_/X sky130_fd_sc_hd__and4_4
X_55088_ _55086_/Y _55076_/X _55087_/X _85321_/D sky130_fd_sc_hd__a21oi_4
X_59965_ _59923_/Y _59943_/A _59880_/X _59884_/X _59927_/A _59968_/A
+ sky130_fd_sc_hd__a41o_4
X_87997_ _88001_/CLK _42176_/X _87997_/Q sky130_fd_sc_hd__dfxtp_4
X_46930_ _46948_/A _52752_/B _46930_/Y sky130_fd_sc_hd__nand2_4
X_58916_ _58913_/Y _58915_/Y _58883_/X _58916_/X sky130_fd_sc_hd__a21o_4
X_54039_ _46471_/A _53964_/B _53969_/C _54039_/X sky130_fd_sc_hd__and3_4
X_42053_ _42052_/X _42043_/X _40909_/X _73438_/A _42044_/X _42053_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77750_ _77747_/X _77751_/C _77751_/B _77752_/A sky130_fd_sc_hd__a21o_4
X_74962_ _74959_/Y _74962_/B _74963_/B sky130_fd_sc_hd__nand2_4
X_70085_ _70048_/A _70085_/X sky130_fd_sc_hd__buf_2
X_86948_ _88215_/CLK _86948_/D _86948_/Q sky130_fd_sc_hd__dfxtp_4
X_59896_ _62288_/A _59896_/X sky130_fd_sc_hd__buf_2
X_41004_ _41003_/X _41004_/X sky130_fd_sc_hd__buf_2
X_76701_ _81351_/D _76691_/A _76701_/X sky130_fd_sc_hd__and2_4
X_73913_ _73911_/X _73913_/B _73913_/C _73913_/Y sky130_fd_sc_hd__nand3_4
X_46861_ _46861_/A _52718_/B sky130_fd_sc_hd__inv_2
X_58847_ _58847_/A _58847_/X sky130_fd_sc_hd__buf_2
X_77681_ _77676_/X _77679_/Y _77677_/Y _77693_/D sky130_fd_sc_hd__nand3_4
X_74893_ _74888_/A _74900_/A _74893_/Y sky130_fd_sc_hd__nand2_4
X_86879_ _86878_/CLK _45407_/Y _61714_/A sky130_fd_sc_hd__dfxtp_4
X_48600_ _48557_/A _50503_/B _48600_/Y sky130_fd_sc_hd__nand2_4
X_79420_ _79419_/B _79419_/A _79420_/X sky130_fd_sc_hd__and2_4
X_45812_ _57468_/A _45740_/B _45812_/Y sky130_fd_sc_hd__nor2_4
X_76632_ _76620_/A _81548_/Q _76633_/A sky130_fd_sc_hd__nand2_4
X_49580_ _49580_/A _49580_/X sky130_fd_sc_hd__buf_2
X_73844_ _72852_/X _73873_/B sky130_fd_sc_hd__buf_2
X_46792_ _46784_/A _46784_/B _46784_/C _46791_/X _46792_/X sky130_fd_sc_hd__and4_4
X_58778_ _58769_/Y _58739_/X _58774_/X _58777_/X _84801_/D sky130_fd_sc_hd__a22oi_4
X_48531_ _40585_/A _48529_/Y _48530_/Y _52175_/A sky130_fd_sc_hd__a21o_4
X_79351_ _84802_/Q _84122_/Q _79351_/X sky130_fd_sc_hd__xor2_4
X_57729_ _57725_/Y _57728_/Y _57718_/X _57729_/X sky130_fd_sc_hd__a21o_4
X_45743_ _45651_/A _45743_/X sky130_fd_sc_hd__buf_2
X_76563_ _76548_/A _76547_/Y _76541_/B _76563_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_5_18_0_CLK clkbuf_4_9_1_CLK/X clkbuf_6_37_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_42955_ _42944_/X _42945_/X _40371_/X _66616_/B _42954_/X _42955_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73775_ _73771_/X _73774_/X _73679_/X _73792_/B sky130_fd_sc_hd__a21o_4
X_70987_ _70976_/A _71073_/B _70990_/C _70987_/Y sky130_fd_sc_hd__nand3_4
X_78302_ _78302_/A _78302_/B _78305_/A sky130_fd_sc_hd__nand2_4
X_75514_ _75514_/A _75513_/X _75514_/X sky130_fd_sc_hd__xor2_4
X_41906_ _51584_/A _51719_/A sky130_fd_sc_hd__buf_2
X_48462_ _48976_/B _48485_/B _48462_/Y sky130_fd_sc_hd__nand2_4
X_60740_ _60662_/A _60711_/A _60632_/X _60702_/C _63436_/A sky130_fd_sc_hd__nand4_4
X_72726_ _72978_/A _72795_/A sky130_fd_sc_hd__buf_2
X_79282_ _79282_/A _79268_/Y _79282_/X sky130_fd_sc_hd__or2_4
X_45674_ _45672_/Y _45596_/X _45644_/X _45673_/Y _45674_/X sky130_fd_sc_hd__a211o_4
X_76494_ _76494_/A _76494_/Y sky130_fd_sc_hd__inv_2
X_42886_ _42820_/X _42886_/X sky130_fd_sc_hd__buf_2
X_47413_ _86637_/Q _47382_/X _47412_/Y _47413_/Y sky130_fd_sc_hd__o21ai_4
X_78233_ _78225_/A _78230_/A _78233_/X sky130_fd_sc_hd__and2_4
X_44625_ _44714_/A _44625_/X sky130_fd_sc_hd__buf_2
X_75445_ _75445_/A _75445_/Y sky130_fd_sc_hd__inv_2
X_41837_ _41837_/A _88129_/D sky130_fd_sc_hd__inv_2
X_60671_ _60671_/A _60671_/B _60671_/C _60671_/Y sky130_fd_sc_hd__nand3_4
X_48393_ _72843_/B _48350_/X _48392_/Y _48393_/Y sky130_fd_sc_hd__o21ai_4
X_72657_ _70198_/C _72645_/X _72656_/Y _83200_/D sky130_fd_sc_hd__a21bo_4
X_62410_ _62399_/X _62406_/Y _62409_/X _84740_/Q _62367_/X _62410_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47344_ _47344_/A _52995_/B sky130_fd_sc_hd__buf_2
X_71608_ _71604_/X _83441_/Q _71607_/Y _83441_/D sky130_fd_sc_hd__a21o_4
X_78164_ _78154_/X _78145_/A _82860_/D _78165_/A sky130_fd_sc_hd__nand3_4
X_44556_ _44556_/A _44556_/Y sky130_fd_sc_hd__inv_2
X_63390_ _63368_/X _63384_/X _63385_/X _63388_/X _63389_/Y _63390_/Y
+ sky130_fd_sc_hd__o41ai_4
X_75376_ _75376_/A _75376_/B _75376_/Y sky130_fd_sc_hd__nand2_4
X_41768_ _41767_/Y _41768_/X sky130_fd_sc_hd__buf_2
X_72588_ _72528_/Y _72607_/B _72597_/C _72583_/C _72525_/A _72588_/Y
+ sky130_fd_sc_hd__a32oi_4
X_77115_ _77115_/A _77112_/C _77115_/X sky130_fd_sc_hd__and2_4
X_43507_ _43495_/X _43503_/X _41762_/X _87386_/Q _43506_/X _43507_/Y
+ sky130_fd_sc_hd__o32ai_4
X_62341_ _62179_/X _62341_/X sky130_fd_sc_hd__buf_2
X_74327_ _72943_/A _74327_/X sky130_fd_sc_hd__buf_2
X_40719_ _40793_/A _40719_/X sky130_fd_sc_hd__buf_2
X_47275_ _47246_/X _47311_/B _47234_/X _52954_/D _47275_/X sky130_fd_sc_hd__and4_4
X_71539_ _70673_/A _71622_/D _71546_/C _71539_/Y sky130_fd_sc_hd__nor3_4
X_78095_ _78096_/B _78095_/Y sky130_fd_sc_hd__inv_2
X_44487_ _44481_/X _44482_/X _41213_/X _87084_/Q _44484_/X _44488_/A
+ sky130_fd_sc_hd__o32ai_4
X_41699_ _40620_/X _41699_/B _41699_/X sky130_fd_sc_hd__or2_4
X_49014_ _83612_/Q _53848_/B sky130_fd_sc_hd__inv_2
X_46226_ _46222_/Y _58151_/A _46225_/Y _46227_/A sky130_fd_sc_hd__nand3_4
X_65060_ _64829_/A _65060_/X sky130_fd_sc_hd__buf_2
XPHY_380 sky130_fd_sc_hd__decap_3
X_77046_ _81992_/Q _82280_/D _77047_/B sky130_fd_sc_hd__nand2_4
X_43438_ _43422_/X _43426_/X _41574_/X _87421_/Q _43434_/X _43439_/A
+ sky130_fd_sc_hd__o32ai_4
X_62272_ _61378_/A _62631_/B _62631_/C _62225_/X _62272_/Y sky130_fd_sc_hd__nand4_4
X_74258_ _74258_/A _74258_/B _74259_/B sky130_fd_sc_hd__nand2_4
XPHY_391 sky130_fd_sc_hd__decap_3
X_64011_ _63206_/B _63947_/B _64040_/C _64025_/D _64011_/Y sky130_fd_sc_hd__nand4_4
X_73209_ _72720_/A _73355_/A sky130_fd_sc_hd__buf_2
X_61223_ _61234_/A _61250_/B _61223_/C _61223_/Y sky130_fd_sc_hd__nor3_4
X_46157_ _46120_/A _46120_/B _86770_/Q _46158_/C sky130_fd_sc_hd__nand3_4
X_43369_ _43369_/A _87456_/D sky130_fd_sc_hd__inv_2
X_74189_ _88344_/Q _72865_/X _72982_/X _74189_/Y sky130_fd_sc_hd__o21ai_4
X_45108_ _45108_/A _45067_/B _45108_/Y sky130_fd_sc_hd__nand2_4
X_61154_ _61176_/B _61151_/Y _61272_/B _61154_/X sky130_fd_sc_hd__o21a_4
X_46088_ _46188_/A _46143_/A sky130_fd_sc_hd__inv_2
X_78997_ _78997_/A _78997_/B _79000_/A sky130_fd_sc_hd__xor2_4
X_60105_ _65515_/A _60105_/X sky130_fd_sc_hd__buf_2
X_49916_ _49904_/A _49915_/X _49904_/C _53129_/D _49916_/X sky130_fd_sc_hd__and4_4
X_45039_ _56216_/C _44998_/X _45038_/X _45039_/Y sky130_fd_sc_hd__o21ai_4
X_68750_ _68750_/A _68750_/B _68750_/X sky130_fd_sc_hd__and2_4
X_65962_ _65958_/X _65960_/X _65961_/X _65962_/X sky130_fd_sc_hd__a21o_4
X_77948_ _82073_/Q _77946_/Y _77947_/X _77948_/Y sky130_fd_sc_hd__o21ai_4
X_61085_ _64249_/A _61085_/X sky130_fd_sc_hd__buf_2
X_67701_ _87972_/Q _67651_/X _67625_/X _67700_/X _67701_/X sky130_fd_sc_hd__a211o_4
X_64913_ _64637_/X _64913_/B _84222_/Q _64913_/X sky130_fd_sc_hd__and3_4
X_60036_ _60036_/A _72564_/A sky130_fd_sc_hd__buf_2
X_49847_ _49842_/Y _49844_/X _49846_/X _86313_/D sky130_fd_sc_hd__a21oi_4
X_68681_ _68604_/A _68681_/B _68681_/X sky130_fd_sc_hd__and2_4
X_65893_ _65859_/X _85570_/Q _65860_/X _65892_/X _65893_/X sky130_fd_sc_hd__a211o_4
X_77879_ _77879_/A _77878_/Y _77880_/B sky130_fd_sc_hd__nand2_4
X_67632_ _46210_/A _68370_/A sky130_fd_sc_hd__buf_2
X_79618_ _79616_/Y _79603_/Y _79609_/A _79619_/B sky130_fd_sc_hd__nand3_4
X_64844_ _64767_/A _64844_/B _64844_/X sky130_fd_sc_hd__and2_4
X_49778_ _49861_/A _49802_/B sky130_fd_sc_hd__buf_2
X_80890_ _80740_/CLK _80890_/D _80890_/Q sky130_fd_sc_hd__dfxtp_4
X_48729_ _48726_/Y _48156_/X _48728_/X _86494_/D sky130_fd_sc_hd__a21oi_4
X_79549_ _65373_/C _79549_/B _79549_/Y sky130_fd_sc_hd__nand2_4
X_67563_ _67539_/X _67563_/B _67563_/X sky130_fd_sc_hd__and2_4
X_64775_ _64775_/A _64775_/B _64775_/Y sky130_fd_sc_hd__nand2_4
X_61987_ _61957_/A _61983_/Y _61984_/Y _61986_/Y _61987_/Y sky130_fd_sc_hd__nand4_4
X_69302_ _69302_/A _87783_/Q _69302_/X sky130_fd_sc_hd__and2_4
X_66514_ _66445_/A _66514_/B _66514_/C _66514_/Y sky130_fd_sc_hd__nor3_4
Xclkbuf_7_101_0_CLK clkbuf_6_50_0_CLK/X clkbuf_8_203_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_51740_ _54400_/A _54317_/A sky130_fd_sc_hd__buf_2
X_63726_ _61301_/X _64192_/B _64192_/C _64189_/D _63726_/Y sky130_fd_sc_hd__nand4_4
X_82560_ _86988_/CLK _82560_/D _82560_/Q sky130_fd_sc_hd__dfxtp_4
X_60938_ _60938_/A _60938_/Y sky130_fd_sc_hd__inv_2
X_67494_ _81499_/D _67449_/X _67493_/X _84067_/D sky130_fd_sc_hd__a21bo_4
X_81511_ _84020_/CLK _81511_/D _81511_/Q sky130_fd_sc_hd__dfxtp_4
X_69233_ _69233_/A _69234_/A sky130_fd_sc_hd__buf_2
X_66445_ _66445_/A _66402_/B _66445_/C _66445_/Y sky130_fd_sc_hd__nor3_4
XPHY_17 sky130_fd_sc_hd__decap_3
X_51671_ _51671_/A _53193_/B _51671_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_71_0_CLK clkbuf_9_35_0_CLK/X _80664_/CLK sky130_fd_sc_hd__clkbuf_1
X_63657_ _63657_/A _62113_/X _63657_/X sky130_fd_sc_hd__and2_4
X_82491_ _82491_/CLK _82491_/D _82491_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_28 sky130_fd_sc_hd__decap_3
X_60869_ _60930_/A _64191_/B sky130_fd_sc_hd__buf_2
XPHY_39 sky130_fd_sc_hd__decap_3
X_53410_ _53397_/A _53402_/B _53410_/C _52895_/D _53410_/X sky130_fd_sc_hd__and4_4
X_84230_ _84150_/CLK _64690_/X _84230_/Q sky130_fd_sc_hd__dfxtp_4
X_50622_ _50597_/A _49006_/X _50622_/Y sky130_fd_sc_hd__nand2_4
X_81442_ _84079_/CLK _76649_/B _81442_/Q sky130_fd_sc_hd__dfxtp_4
X_62608_ _62269_/X _58207_/A _62618_/C _62608_/D _62608_/X sky130_fd_sc_hd__and4_4
X_69164_ _88049_/Q _69162_/X _68884_/X _69163_/X _69164_/X sky130_fd_sc_hd__a211o_4
X_54390_ _54395_/A _54395_/B _54395_/C _46828_/Y _54390_/X sky130_fd_sc_hd__and4_4
X_66376_ _66366_/X _64675_/Y _66375_/Y _66376_/Y sky130_fd_sc_hd__o21ai_4
X_63588_ _58442_/A _63541_/B _63575_/C _63541_/D _63588_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_7_116_0_CLK clkbuf_6_58_0_CLK/X clkbuf_8_233_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_68115_ _68088_/X _66720_/Y _68110_/X _68114_/Y _68115_/X sky130_fd_sc_hd__a211o_4
X_53341_ _53332_/A _47053_/A _53341_/Y sky130_fd_sc_hd__nand2_4
X_65327_ _65403_/A _65327_/B _65327_/X sky130_fd_sc_hd__and2_4
X_84161_ _84161_/CLK _84161_/D _84161_/Q sky130_fd_sc_hd__dfxtp_4
X_50553_ _50550_/Y _50551_/X _50552_/X _50553_/Y sky130_fd_sc_hd__a21oi_4
X_62539_ _62529_/X _62536_/Y _62538_/X _84843_/Q _62511_/X _62539_/Y
+ sky130_fd_sc_hd__o32ai_4
X_81373_ _81265_/CLK _81373_/D _81373_/Q sky130_fd_sc_hd__dfxtp_4
X_69095_ _68649_/A _69095_/X sky130_fd_sc_hd__buf_2
X_83112_ _83846_/CLK _83112_/D _83112_/Q sky130_fd_sc_hd__dfxtp_4
X_80324_ _80324_/A _80324_/Y sky130_fd_sc_hd__inv_2
X_68046_ _68043_/X _68045_/X _67977_/X _68049_/A sky130_fd_sc_hd__a21o_4
X_56060_ _56059_/Y _56060_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_86_0_CLK clkbuf_9_43_0_CLK/X _84892_/CLK sky130_fd_sc_hd__clkbuf_1
X_53272_ _51823_/A _53272_/X sky130_fd_sc_hd__buf_2
X_65258_ _65258_/A _85800_/Q _65258_/X sky130_fd_sc_hd__and2_4
X_84092_ _81507_/CLK _84092_/D _80916_/D sky130_fd_sc_hd__dfxtp_4
X_50484_ _50482_/Y _50474_/X _50483_/Y _50484_/Y sky130_fd_sc_hd__a21boi_4
X_55011_ _55011_/A _47623_/A _55011_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_232_0_CLK clkbuf_8_233_0_CLK/A clkbuf_8_232_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_52223_ _48841_/A _52198_/X _52223_/C _52223_/X sky130_fd_sc_hd__and3_4
X_87920_ _87473_/CLK _87920_/D _87920_/Q sky130_fd_sc_hd__dfxtp_4
X_64209_ _61117_/X _61169_/X _59477_/A _64209_/Y sky130_fd_sc_hd__nand3_4
X_83043_ _85428_/CLK _74532_/Y _47052_/A sky130_fd_sc_hd__dfxtp_4
X_80255_ _80242_/A _80241_/X _80254_/Y _80256_/B sky130_fd_sc_hd__a21boi_4
X_65189_ _64602_/A _65753_/A sky130_fd_sc_hd__buf_2
X_52154_ _52168_/A _48482_/B _52154_/Y sky130_fd_sc_hd__nand2_4
X_87851_ _87851_/CLK _42479_/Y _73750_/A sky130_fd_sc_hd__dfxtp_4
X_80186_ _80186_/A _84291_/Q _80186_/X sky130_fd_sc_hd__xor2_4
X_69997_ _82557_/D _69988_/X _69996_/Y _69997_/X sky130_fd_sc_hd__a21bo_4
X_51105_ _51084_/A _51115_/B _51110_/C _52797_/D _51105_/X sky130_fd_sc_hd__and4_4
X_86802_ _87484_/CLK _46035_/X _86802_/Q sky130_fd_sc_hd__dfxtp_4
X_59750_ _59755_/A _72584_/C sky130_fd_sc_hd__buf_2
X_52085_ _52121_/A _50383_/B _52085_/Y sky130_fd_sc_hd__nand2_4
X_56962_ _56626_/X _56952_/A _56961_/Y _85111_/D sky130_fd_sc_hd__a21oi_4
X_68948_ _69485_/A _68948_/X sky130_fd_sc_hd__buf_2
X_87782_ _87782_/CLK _42662_/Y _87782_/Q sky130_fd_sc_hd__dfxtp_4
X_84994_ _85100_/CLK _84994_/D _84994_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_247_0_CLK clkbuf_8_247_0_CLK/A clkbuf_9_495_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_242_0_CLK clkbuf_9_121_0_CLK/X _84452_/CLK sky130_fd_sc_hd__clkbuf_1
X_58701_ _58701_/A _58701_/X sky130_fd_sc_hd__buf_2
X_51036_ _51032_/Y _51011_/X _51035_/X _86086_/D sky130_fd_sc_hd__a21oi_4
X_55913_ _55620_/A _55913_/B _55913_/X sky130_fd_sc_hd__and2_4
X_86733_ _86733_/CLK _46488_/Y _86733_/Q sky130_fd_sc_hd__dfxtp_4
X_59681_ _59681_/A _59836_/D sky130_fd_sc_hd__buf_2
X_83945_ _83973_/CLK _83945_/D _83945_/Q sky130_fd_sc_hd__dfxtp_4
X_56893_ _56859_/X _56893_/B _56893_/Y sky130_fd_sc_hd__nor2_4
X_68879_ _68874_/X _68877_/X _68878_/X _68879_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_872_0_CLK clkbuf_9_436_0_CLK/X _86587_/CLK sky130_fd_sc_hd__clkbuf_1
X_70910_ _70866_/A _70914_/B sky130_fd_sc_hd__buf_2
X_58632_ _58749_/A _58659_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_24_0_CLK clkbuf_9_12_0_CLK/X _85249_/CLK sky130_fd_sc_hd__clkbuf_1
X_55844_ _45168_/A _55572_/X _44098_/X _55843_/X _55844_/X sky130_fd_sc_hd__a211o_4
X_86664_ _86665_/CLK _47164_/Y _86664_/Q sky130_fd_sc_hd__dfxtp_4
X_71890_ _71870_/Y _83338_/Q _71889_/Y _83338_/D sky130_fd_sc_hd__a21o_4
X_83876_ _82557_/CLK _83876_/D _82556_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_363_0_CLK clkbuf_9_363_0_CLK/A clkbuf_9_363_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_88403_ _87373_/CLK _88403_/D _88403_/Q sky130_fd_sc_hd__dfxtp_4
X_85615_ _83544_/CLK _85615_/D _85615_/Q sky130_fd_sc_hd__dfxtp_4
X_70841_ _70869_/A _70846_/B _70849_/C _70841_/D _70841_/Y sky130_fd_sc_hd__nand4_4
X_58563_ _58559_/X _83354_/Q _58562_/Y _84818_/D sky130_fd_sc_hd__o21a_4
X_82827_ _82462_/CLK _82827_/D _82827_/Q sky130_fd_sc_hd__dfxtp_4
X_55775_ _56253_/C _55747_/X _55165_/X _55774_/X _55775_/X sky130_fd_sc_hd__a211o_4
X_86595_ _85955_/CLK _86595_/D _86595_/Q sky130_fd_sc_hd__dfxtp_4
X_52987_ _85718_/Q _52984_/X _52986_/Y _52987_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_257_0_CLK clkbuf_9_128_0_CLK/X _84849_/CLK sky130_fd_sc_hd__clkbuf_1
X_57514_ _84988_/Q _57493_/X _57513_/Y _57514_/Y sky130_fd_sc_hd__o21ai_4
X_88334_ _84970_/CLK _88334_/D _88334_/Q sky130_fd_sc_hd__dfxtp_4
X_42740_ _42723_/A _42740_/X sky130_fd_sc_hd__buf_2
X_54726_ _54672_/X _54748_/C sky130_fd_sc_hd__buf_2
X_73560_ _72757_/A _73583_/A sky130_fd_sc_hd__buf_2
X_85546_ _86145_/CLK _85546_/D _85546_/Q sky130_fd_sc_hd__dfxtp_4
X_51938_ _51933_/Y _51934_/X _51937_/Y _85920_/D sky130_fd_sc_hd__a21boi_4
X_70772_ _70772_/A _70791_/C sky130_fd_sc_hd__buf_2
X_58494_ _64467_/C _58495_/A sky130_fd_sc_hd__buf_2
X_82758_ _82774_/CLK _82758_/D _82758_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_887_0_CLK clkbuf_9_443_0_CLK/X _85818_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_39_0_CLK clkbuf_9_19_0_CLK/X _85089_/CLK sky130_fd_sc_hd__clkbuf_1
X_72511_ _72592_/A _61414_/A _79513_/B _72511_/Y sky130_fd_sc_hd__nor3_4
X_81709_ _81755_/CLK _81333_/Q _81709_/Q sky130_fd_sc_hd__dfxtp_4
X_57445_ _57029_/A _57445_/B _56812_/X _57445_/Y sky130_fd_sc_hd__nand3_4
X_88265_ _88268_/CLK _88265_/D _68631_/B sky130_fd_sc_hd__dfxtp_4
X_42671_ _42665_/X _42666_/X _41036_/X _69381_/B _42658_/X _42672_/A
+ sky130_fd_sc_hd__o32ai_4
X_54657_ _54656_/X _54674_/B sky130_fd_sc_hd__buf_2
X_85477_ _84926_/CLK _54248_/Y _85477_/Q sky130_fd_sc_hd__dfxtp_4
X_73491_ _72899_/A _73491_/X sky130_fd_sc_hd__buf_2
X_51869_ _51843_/A _51870_/B sky130_fd_sc_hd__buf_2
X_82689_ _81216_/CLK _78793_/A _78309_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_378_0_CLK clkbuf_9_378_0_CLK/A clkbuf_9_378_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_44410_ _44410_/A _87123_/D sky130_fd_sc_hd__inv_2
X_87216_ _87408_/CLK _87216_/D _87216_/Q sky130_fd_sc_hd__dfxtp_4
X_75230_ _75228_/X _75230_/B _75230_/X sky130_fd_sc_hd__and2_4
X_41622_ _41611_/X _41613_/X _41621_/X _88181_/Q _41608_/X _41623_/A
+ sky130_fd_sc_hd__o32ai_4
X_53608_ _53604_/A _50385_/B _53608_/Y sky130_fd_sc_hd__nand2_4
X_72442_ _57697_/X _85958_/Q _72441_/X _72442_/Y sky130_fd_sc_hd__o21ai_4
X_84428_ _84426_/CLK _84428_/D _78051_/B sky130_fd_sc_hd__dfxtp_4
X_45390_ _45389_/X _45390_/X sky130_fd_sc_hd__buf_2
X_57376_ _73476_/A _57376_/X sky130_fd_sc_hd__buf_2
X_88196_ _88133_/CLK _41539_/Y _66932_/B sky130_fd_sc_hd__dfxtp_4
X_54588_ _85414_/Q _54567_/X _54587_/Y _54588_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_810_0_CLK clkbuf_9_405_0_CLK/X _82299_/CLK sky130_fd_sc_hd__clkbuf_1
X_59115_ _58918_/A _59115_/X sky130_fd_sc_hd__buf_2
X_44341_ _44330_/X _44331_/X _41688_/X _87157_/Q _44332_/X _44341_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56327_ _56079_/X _56321_/X _56326_/Y _85235_/D sky130_fd_sc_hd__o21ai_4
X_75161_ _75155_/Y _75161_/B _75159_/Y _75162_/B sky130_fd_sc_hd__nand3_4
X_87147_ _88164_/CLK _44361_/Y _87147_/Q sky130_fd_sc_hd__dfxtp_4
X_41553_ _41552_/X _41530_/X _88194_/Q _41531_/X _88194_/D sky130_fd_sc_hd__a2bb2o_4
X_53539_ _53536_/Y _53537_/X _53538_/X _85617_/D sky130_fd_sc_hd__a21oi_4
X_72373_ _57709_/X _85356_/Q _72372_/X _72373_/Y sky130_fd_sc_hd__o21ai_4
X_84359_ _84360_/CLK _63035_/X _79493_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_301_0_CLK clkbuf_8_150_0_CLK/X clkbuf_9_301_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_74112_ _73588_/A _66242_/B _74112_/X sky130_fd_sc_hd__and2_4
X_40504_ _40324_/X _40504_/X sky130_fd_sc_hd__buf_2
X_47060_ _47055_/Y _47035_/X _47059_/X _86675_/D sky130_fd_sc_hd__a21oi_4
X_71324_ _50358_/B _71320_/X _71323_/Y _71324_/Y sky130_fd_sc_hd__o21ai_4
X_59046_ _58603_/A _59046_/X sky130_fd_sc_hd__buf_2
X_44272_ _72838_/A _44272_/X sky130_fd_sc_hd__buf_2
X_56258_ _56245_/A _56263_/B sky130_fd_sc_hd__buf_2
X_87078_ _88267_/CLK _87078_/D _87078_/Q sky130_fd_sc_hd__dfxtp_4
X_75092_ _75090_/X _75107_/A _75092_/X sky130_fd_sc_hd__and2_4
X_41484_ _41481_/X _82332_/Q _41483_/X _41484_/Y sky130_fd_sc_hd__o21ai_4
X_46011_ _46011_/A _46011_/Y sky130_fd_sc_hd__inv_2
X_43223_ _43223_/A _87531_/D sky130_fd_sc_hd__inv_2
X_55209_ _82981_/Q _55190_/X _55172_/X _55208_/Y _55209_/X sky130_fd_sc_hd__a211o_4
X_74043_ _74022_/X _86541_/Q _74043_/X sky130_fd_sc_hd__and2_4
X_78920_ _82734_/Q _78920_/B _78920_/X sky130_fd_sc_hd__xor2_4
X_86029_ _86029_/CLK _86029_/D _65120_/B sky130_fd_sc_hd__dfxtp_4
X_40435_ _40435_/A _40686_/A sky130_fd_sc_hd__buf_2
X_71255_ _70819_/A _71256_/B sky130_fd_sc_hd__buf_2
X_56189_ _56186_/Y _56252_/A sky130_fd_sc_hd__buf_2
Xclkbuf_10_825_0_CLK clkbuf_9_412_0_CLK/X _82368_/CLK sky130_fd_sc_hd__clkbuf_1
X_70206_ _70195_/X _83838_/Q _70205_/X _70206_/X sky130_fd_sc_hd__a21o_4
X_43154_ _43121_/A _43154_/X sky130_fd_sc_hd__buf_2
X_78851_ _82727_/Q _78851_/B _78851_/X sky130_fd_sc_hd__xor2_4
X_40366_ _40365_/X _41061_/A sky130_fd_sc_hd__buf_2
X_71186_ _48788_/B _71164_/Y _71185_/Y _71186_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_316_0_CLK clkbuf_8_158_0_CLK/X clkbuf_9_316_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_42105_ _41032_/X _42103_/X _88034_/Q _42104_/X _88034_/D sky130_fd_sc_hd__a2bb2o_4
X_77802_ _77782_/Y _77796_/Y _77801_/X _77802_/Y sky130_fd_sc_hd__a21oi_4
X_70137_ _83521_/Q _83169_/Q _83504_/Q _83152_/Q _70139_/C sky130_fd_sc_hd__a22oi_4
X_47962_ _66084_/B _47948_/X _47961_/Y _47962_/Y sky130_fd_sc_hd__o21ai_4
X_43085_ _43129_/A _43085_/X sky130_fd_sc_hd__buf_2
X_59948_ _62198_/B _59950_/B sky130_fd_sc_hd__buf_2
X_78782_ _78782_/A _78778_/X _78782_/Y sky130_fd_sc_hd__nand2_4
X_75994_ _75990_/Y _75993_/X _75994_/Y sky130_fd_sc_hd__nand2_4
X_49701_ _49685_/A _49697_/B _49685_/C _51225_/D _49701_/X sky130_fd_sc_hd__and4_4
X_46913_ _46948_/A _46912_/X _46913_/Y sky130_fd_sc_hd__nand2_4
X_42036_ _42036_/A _42036_/Y sky130_fd_sc_hd__inv_2
X_77733_ _77730_/Y _77732_/Y _77725_/Y _77743_/A sky130_fd_sc_hd__a21oi_4
X_74945_ _81135_/D _74945_/B _74945_/Y sky130_fd_sc_hd__nand2_4
X_70068_ _69876_/X _69878_/X _68400_/X _70068_/Y sky130_fd_sc_hd__a21oi_4
X_47893_ _47893_/A _46579_/X _47893_/X sky130_fd_sc_hd__or2_4
Xclkbuf_5_1_0_CLK clkbuf_4_0_1_CLK/X clkbuf_6_3_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_59879_ _59579_/A _59585_/A _60174_/D sky130_fd_sc_hd__nor2_4
X_61910_ _61909_/X _61846_/B _61878_/C _61910_/D _61910_/Y sky130_fd_sc_hd__nand4_4
X_49632_ _49632_/A _49632_/X sky130_fd_sc_hd__buf_2
X_46844_ _46751_/A _46844_/X sky130_fd_sc_hd__buf_2
X_77664_ _77666_/A _77638_/Y _77664_/C _77639_/Y _77665_/A sky130_fd_sc_hd__nand4_4
X_62890_ _62717_/A _62967_/D sky130_fd_sc_hd__buf_2
X_74876_ _81126_/D _74869_/B _74876_/Y sky130_fd_sc_hd__nand2_4
X_79403_ _79395_/A _79395_/B _79402_/Y _79419_/A sky130_fd_sc_hd__a21boi_4
X_76615_ _76614_/X _76615_/Y sky130_fd_sc_hd__inv_2
X_49563_ _49558_/A _52777_/B _49563_/Y sky130_fd_sc_hd__nand2_4
X_61841_ _61419_/X _61794_/B _61809_/C _61776_/D _61847_/B sky130_fd_sc_hd__nand4_4
X_73827_ _73733_/A _73827_/B _73827_/X sky130_fd_sc_hd__and2_4
X_46775_ _46774_/Y _46775_/X sky130_fd_sc_hd__buf_2
X_77595_ _77593_/Y _77564_/B _77594_/X _77596_/B sky130_fd_sc_hd__o21ai_4
X_43987_ _43987_/A _43987_/B _43987_/Y sky130_fd_sc_hd__nor2_4
X_48514_ _48514_/A _50466_/B sky130_fd_sc_hd__buf_2
X_79334_ _79334_/A _79334_/B _79334_/X sky130_fd_sc_hd__and2_4
X_45726_ _85132_/Q _45709_/X _45651_/X _45726_/X sky130_fd_sc_hd__o21a_4
X_64560_ _64558_/Y _59655_/X _64559_/Y _64560_/Y sky130_fd_sc_hd__a21oi_4
X_76546_ _76519_/X _76544_/Y _76545_/Y _76546_/X sky130_fd_sc_hd__a21bo_4
X_42938_ _42937_/Y _87642_/D sky130_fd_sc_hd__inv_2
X_61772_ _61839_/A _61791_/B _61732_/X _63041_/B _61772_/X sky130_fd_sc_hd__and4_4
X_49494_ _49500_/A _49500_/B _49493_/X _52709_/D _49494_/X sky130_fd_sc_hd__and4_4
X_73758_ _73731_/X _86233_/Q _73683_/X _73757_/X _73758_/X sky130_fd_sc_hd__a211o_4
X_63511_ _63488_/A _61922_/X _63511_/X sky130_fd_sc_hd__and2_4
X_48445_ _74403_/B _52137_/B sky130_fd_sc_hd__buf_2
X_72709_ _72943_/A _72709_/X sky130_fd_sc_hd__buf_2
X_60723_ _60722_/Y _59755_/A _60696_/Y _60723_/X sky130_fd_sc_hd__and3_4
X_79265_ _79258_/X _79260_/B _79264_/Y _79282_/A sky130_fd_sc_hd__a21boi_4
X_45657_ _45591_/X _61528_/A _45608_/X _45657_/Y sky130_fd_sc_hd__o21ai_4
X_64491_ _64489_/Y _59655_/X _64490_/Y _84241_/D sky130_fd_sc_hd__a21oi_4
X_76477_ _76477_/A _76479_/B sky130_fd_sc_hd__inv_2
X_42869_ _42847_/X _42849_/X _41574_/X _67095_/B _42858_/X _42870_/A
+ sky130_fd_sc_hd__o32ai_4
X_73689_ _73641_/A _73689_/B _73689_/X sky130_fd_sc_hd__and2_4
X_66230_ _66179_/X _66228_/Y _66229_/Y _66230_/Y sky130_fd_sc_hd__o21ai_4
X_78216_ _78203_/A _82492_/Q _78215_/Y _78217_/B sky130_fd_sc_hd__a21oi_4
X_44608_ _40954_/Y _44602_/X _87036_/Q _44603_/X _44608_/X sky130_fd_sc_hd__a2bb2o_4
X_63442_ _61398_/B _63426_/X _63439_/X _63441_/X _63442_/X sky130_fd_sc_hd__a211o_4
X_75428_ _75427_/B _75427_/C _75423_/Y _75432_/C sky130_fd_sc_hd__o21ai_4
X_48376_ _74371_/A _52103_/A sky130_fd_sc_hd__buf_2
X_60654_ _63471_/A _60654_/X sky130_fd_sc_hd__buf_2
X_79196_ _79198_/B _79196_/Y sky130_fd_sc_hd__inv_2
X_45588_ _55499_/B _45507_/X _45429_/X _45588_/X sky130_fd_sc_hd__o21a_4
X_47327_ _47140_/A _47370_/C sky130_fd_sc_hd__buf_2
X_66161_ _66453_/A _66385_/B _66160_/X _66161_/Y sky130_fd_sc_hd__nand3_4
X_78147_ _78137_/Y _78146_/X _78147_/Y sky130_fd_sc_hd__nand2_4
X_63373_ _58409_/A _63370_/X _61338_/A _63372_/X _63373_/X sky130_fd_sc_hd__a2bb2o_4
X_44539_ _44539_/A _44539_/Y sky130_fd_sc_hd__inv_2
X_75359_ _75348_/Y _75349_/Y _75351_/A _75359_/X sky130_fd_sc_hd__o21a_4
X_60585_ _60583_/Y _60444_/Y _60584_/Y _79134_/A _60341_/X _60585_/X
+ sky130_fd_sc_hd__o32a_4
X_65112_ _60151_/X _65102_/Y _65111_/Y _65112_/Y sky130_fd_sc_hd__o21ai_4
X_62324_ _62597_/B _61844_/X _62237_/X _62280_/D _62324_/X sky130_fd_sc_hd__and4_4
X_47258_ _47254_/Y _47224_/X _47257_/X _86654_/D sky130_fd_sc_hd__a21oi_4
X_66092_ _66164_/A _65888_/B _66092_/C _66092_/Y sky130_fd_sc_hd__nor3_4
X_78078_ _60700_/C _78078_/B _78078_/X sky130_fd_sc_hd__xor2_4
X_46209_ _44244_/A _46210_/A sky130_fd_sc_hd__buf_2
X_65043_ _64915_/X _65031_/Y _65042_/Y _65043_/Y sky130_fd_sc_hd__o21ai_4
X_69920_ _57804_/A _43741_/Y _69920_/Y sky130_fd_sc_hd__nor2_4
X_77029_ _77036_/A _77036_/B _77034_/C sky130_fd_sc_hd__xor2_4
X_62255_ _62252_/Y _62253_/X _62254_/Y _62255_/Y sky130_fd_sc_hd__a21oi_4
X_47189_ _47189_/A _51214_/D sky130_fd_sc_hd__buf_2
X_61206_ _64274_/A _64223_/C sky130_fd_sc_hd__buf_2
X_80040_ _60103_/C _80040_/B _80046_/B sky130_fd_sc_hd__xor2_4
X_69851_ _42036_/A _69582_/X _69567_/X _69850_/Y _69851_/X sky130_fd_sc_hd__a211o_4
X_62186_ _62186_/A _62186_/X sky130_fd_sc_hd__buf_2
X_68802_ _69735_/A _68802_/B _68802_/Y sky130_fd_sc_hd__nor2_4
X_61137_ _72543_/A _61165_/A sky130_fd_sc_hd__buf_2
X_69782_ _69778_/X _69781_/X _69768_/X _69785_/A sky130_fd_sc_hd__a21o_4
X_66994_ _66758_/X _66994_/X sky130_fd_sc_hd__buf_2
X_68733_ _73895_/A _68626_/X _68731_/X _68732_/Y _68733_/X sky130_fd_sc_hd__a211o_4
X_65945_ _65932_/A _73636_/B _65945_/X sky130_fd_sc_hd__and2_4
X_61068_ _61066_/Y _61112_/A _64361_/A sky130_fd_sc_hd__and2_4
X_81991_ _81990_/CLK _81991_/D _77036_/A sky130_fd_sc_hd__dfxtp_4
X_52910_ _52910_/A _47195_/X _52910_/Y sky130_fd_sc_hd__nand2_4
X_60019_ _60079_/B _59922_/C _62556_/A _60019_/Y sky130_fd_sc_hd__o21ai_4
X_83730_ _84930_/CLK _70659_/Y _83730_/Q sky130_fd_sc_hd__dfxtp_4
X_80942_ _80818_/CLK _80986_/Q _74935_/A sky130_fd_sc_hd__dfxtp_4
X_68664_ _80822_/D _68586_/X _68663_/X _83966_/D sky130_fd_sc_hd__a21bo_4
Xclkbuf_7_93_0_CLK clkbuf_7_93_0_CLK/A clkbuf_7_93_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_53890_ _53871_/X _49106_/Y _53890_/Y sky130_fd_sc_hd__nand2_4
X_65876_ _65118_/A _65876_/X sky130_fd_sc_hd__buf_2
X_67615_ _66554_/X _67615_/X sky130_fd_sc_hd__buf_2
X_52841_ _52853_/A _52831_/B _52818_/C _52841_/D _52841_/X sky130_fd_sc_hd__and4_4
X_64827_ _64752_/X _86169_/Q _64716_/X _64826_/X _64827_/X sky130_fd_sc_hd__a211o_4
X_83661_ _83663_/CLK _83661_/D _83661_/Q sky130_fd_sc_hd__dfxtp_4
X_80873_ _80746_/CLK _75635_/B _80873_/Q sky130_fd_sc_hd__dfxtp_4
X_68595_ _68444_/A _68595_/B _68595_/X sky130_fd_sc_hd__and2_4
X_85400_ _83745_/CLK _54668_/Y _85400_/Q sky130_fd_sc_hd__dfxtp_4
X_82612_ _82518_/CLK _78975_/B _82612_/Q sky130_fd_sc_hd__dfxtp_4
X_55560_ _55475_/X _45488_/Y _55560_/Y sky130_fd_sc_hd__nor2_4
X_67546_ _87978_/Q _67473_/X _67524_/X _67545_/X _67546_/X sky130_fd_sc_hd__a211o_4
X_86380_ _86381_/CLK _49480_/Y _58830_/B sky130_fd_sc_hd__dfxtp_4
X_52772_ _52769_/Y _52755_/X _52771_/X _52772_/Y sky130_fd_sc_hd__a21oi_4
X_64758_ _45926_/X _64758_/X sky130_fd_sc_hd__buf_2
X_83592_ _83589_/CLK _83592_/D _83592_/Q sky130_fd_sc_hd__dfxtp_4
X_54511_ _54034_/A _54540_/A sky130_fd_sc_hd__buf_2
X_85331_ _85332_/CLK _85331_/D _85331_/Q sky130_fd_sc_hd__dfxtp_4
X_51723_ _51718_/Y _51719_/X _51722_/X _85958_/D sky130_fd_sc_hd__a21oi_4
X_63709_ _63368_/A _63703_/X _63704_/X _63707_/X _63708_/Y _63709_/Y
+ sky130_fd_sc_hd__o41ai_4
X_82543_ _82553_/CLK _82543_/D _82543_/Q sky130_fd_sc_hd__dfxtp_4
X_55491_ _55491_/A _55490_/X _55491_/X sky130_fd_sc_hd__and2_4
X_67477_ _67359_/X _67477_/X sky130_fd_sc_hd__buf_2
X_64689_ _64689_/A _64741_/B _64688_/Y _64689_/Y sky130_fd_sc_hd__nor3_4
X_57230_ _72484_/A _72710_/A _46173_/X _57223_/D _56923_/Y _57230_/Y
+ sky130_fd_sc_hd__a41oi_4
X_69216_ _69146_/A _69216_/X sky130_fd_sc_hd__buf_2
X_88050_ _88084_/CLK _88050_/D _88050_/Q sky130_fd_sc_hd__dfxtp_4
X_54442_ _54446_/A _54442_/B _54442_/Y sky130_fd_sc_hd__nand2_4
X_66428_ _84125_/Q _66429_/C sky130_fd_sc_hd__inv_2
X_85262_ _85198_/CLK _85262_/D _56243_/C sky130_fd_sc_hd__dfxtp_4
X_51654_ _85970_/Q _51647_/X _51653_/Y _51654_/Y sky130_fd_sc_hd__o21ai_4
X_82474_ _82595_/CLK _82474_/D _78083_/B sky130_fd_sc_hd__dfxtp_4
X_87001_ _83139_/CLK _44685_/Y _87001_/Q sky130_fd_sc_hd__dfxtp_4
X_84213_ _84228_/CLK _65143_/X _84213_/Q sky130_fd_sc_hd__dfxtp_4
X_50605_ _50580_/A _71998_/B _50605_/Y sky130_fd_sc_hd__nand2_4
X_57161_ _55320_/B _57106_/X _57160_/Y _57161_/Y sky130_fd_sc_hd__o21ai_4
X_81425_ _81333_/CLK _81425_/D _76027_/B sky130_fd_sc_hd__dfxtp_4
X_69147_ _69067_/A _69147_/B _69147_/X sky130_fd_sc_hd__and2_4
X_54373_ _54395_/A _54362_/B _54395_/C _46800_/Y _54373_/X sky130_fd_sc_hd__and4_4
X_66359_ _66318_/X _66319_/B _84138_/Q _66359_/X sky130_fd_sc_hd__and3_4
X_85193_ _85192_/CLK _56441_/Y _85193_/Q sky130_fd_sc_hd__dfxtp_4
X_51585_ _51639_/A _51585_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_31_0_CLK clkbuf_7_31_0_CLK/A clkbuf_8_63_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_56112_ _56142_/A _56112_/X sky130_fd_sc_hd__buf_2
X_53324_ _51900_/A _53324_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_171_0_CLK clkbuf_7_85_0_CLK/X clkbuf_9_343_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_84144_ _84175_/CLK _84144_/D _84144_/Q sky130_fd_sc_hd__dfxtp_4
X_50536_ _86182_/Q _50533_/X _50535_/Y _50536_/Y sky130_fd_sc_hd__o21ai_4
X_57092_ _73198_/B _57092_/X sky130_fd_sc_hd__buf_2
X_81356_ _81431_/CLK _76749_/Y _81356_/Q sky130_fd_sc_hd__dfxtp_4
X_69078_ _69011_/A _87222_/Q _69078_/X sky130_fd_sc_hd__and2_4
X_56043_ _55912_/X _55916_/X _56043_/X sky130_fd_sc_hd__and2_4
X_68029_ _87958_/Q _68006_/X _67984_/X _68028_/X _68029_/X sky130_fd_sc_hd__a211o_4
X_80307_ _80310_/B _80308_/A sky130_fd_sc_hd__inv_2
X_53255_ _53259_/A _53255_/B _53255_/Y sky130_fd_sc_hd__nand2_4
X_84075_ _84074_/CLK _84075_/D _80899_/D sky130_fd_sc_hd__dfxtp_4
X_50467_ _86195_/Q _50464_/X _50466_/Y _50467_/Y sky130_fd_sc_hd__o21ai_4
X_81287_ _81603_/CLK _76975_/X _81255_/D sky130_fd_sc_hd__dfxtp_4
X_52206_ _52185_/X _48820_/B _52206_/Y sky130_fd_sc_hd__nand2_4
X_71040_ _53174_/B _71013_/A _71039_/Y _71040_/Y sky130_fd_sc_hd__o21ai_4
X_83026_ _83025_/CLK _83026_/D _83026_/Q sky130_fd_sc_hd__dfxtp_4
X_87903_ _87898_/CLK _42360_/Y _87903_/Q sky130_fd_sc_hd__dfxtp_4
X_80238_ _84951_/Q _65466_/C _80238_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_7_46_0_CLK clkbuf_7_47_0_CLK/A clkbuf_8_93_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_53186_ _53184_/Y _53163_/X _53185_/X _85681_/D sky130_fd_sc_hd__a21oi_4
X_50398_ _50398_/A _48368_/X _50398_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_8_186_0_CLK clkbuf_7_93_0_CLK/X clkbuf_9_373_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_59802_ _70009_/A _59802_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_181_0_CLK clkbuf_9_90_0_CLK/X _83337_/CLK sky130_fd_sc_hd__clkbuf_1
X_52137_ _52127_/X _52137_/B _52137_/Y sky130_fd_sc_hd__nand2_4
X_87834_ _87834_/CLK _87834_/D _74143_/A sky130_fd_sc_hd__dfxtp_4
X_80169_ _80151_/Y _80169_/B _80169_/X sky130_fd_sc_hd__or2_4
X_57994_ _57989_/X _57991_/Y _57992_/Y _57893_/X _57993_/X _57994_/X
+ sky130_fd_sc_hd__o32a_4
X_59733_ _59754_/A _59731_/Y _59754_/C _59733_/Y sky130_fd_sc_hd__nand3_4
X_56945_ _44214_/X _56575_/X _85119_/Q _56943_/X _85119_/D sky130_fd_sc_hd__a2bb2o_4
X_52068_ _52083_/A _50368_/B _52068_/Y sky130_fd_sc_hd__nand2_4
X_87765_ _87766_/CLK _87765_/D _69542_/B sky130_fd_sc_hd__dfxtp_4
X_72991_ _72987_/X _72990_/X _72739_/X _72995_/A sky130_fd_sc_hd__a21o_4
X_84977_ _86238_/CLK _84977_/D _84977_/Q sky130_fd_sc_hd__dfxtp_4
X_43910_ _41367_/X _43907_/X _87204_/Q _43908_/X _43910_/X sky130_fd_sc_hd__a2bb2o_4
X_51019_ _51017_/Y _51011_/X _51018_/X _86089_/D sky130_fd_sc_hd__a21oi_4
X_86716_ _86398_/CLK _46671_/Y _58634_/A sky130_fd_sc_hd__dfxtp_4
X_74730_ _74722_/Y _74730_/B _74730_/C _74729_/Y _74730_/Y sky130_fd_sc_hd__nand4_4
X_83928_ _81473_/CLK _69380_/X _83928_/Q sky130_fd_sc_hd__dfxtp_4
X_71942_ _71938_/Y _71942_/Y sky130_fd_sc_hd__inv_2
X_59664_ _59664_/A _59679_/A _59664_/C _59754_/D _59665_/A sky130_fd_sc_hd__and4_4
X_44890_ _44877_/Y _44886_/Y _44889_/X _44890_/X sky130_fd_sc_hd__a21o_4
X_56876_ _83331_/Q _56876_/X sky130_fd_sc_hd__buf_2
X_87696_ _87952_/CLK _87696_/D _66651_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_196_0_CLK clkbuf_9_98_0_CLK/X _84668_/CLK sky130_fd_sc_hd__clkbuf_1
X_58615_ _58585_/X _58613_/Y _58614_/Y _58603_/X _58589_/X _58615_/X
+ sky130_fd_sc_hd__o32a_4
X_43841_ _43602_/X _43842_/A sky130_fd_sc_hd__buf_2
X_55827_ _45181_/A _55498_/X _44096_/X _55826_/X _55827_/X sky130_fd_sc_hd__a211o_4
X_74661_ _56696_/A _74641_/X _74660_/Y _82993_/D sky130_fd_sc_hd__a21boi_4
X_86647_ _86647_/CLK _86647_/D _86647_/Q sky130_fd_sc_hd__dfxtp_4
X_71873_ _71783_/C _71873_/X sky130_fd_sc_hd__buf_2
X_59595_ _45941_/A _44003_/A _59584_/C _60182_/A sky130_fd_sc_hd__nor3_4
X_83859_ _82541_/CLK _70066_/X _83859_/Q sky130_fd_sc_hd__dfxtp_4
X_76400_ _76391_/X _76396_/X _76400_/C _76400_/X sky130_fd_sc_hd__or3_4
X_73612_ _73262_/A _73612_/X sky130_fd_sc_hd__buf_2
X_70824_ _70824_/A _71066_/B sky130_fd_sc_hd__buf_2
X_46560_ _51376_/B _54075_/B sky130_fd_sc_hd__buf_2
X_58546_ _58546_/A _58546_/Y sky130_fd_sc_hd__inv_2
X_77380_ _77380_/A _82093_/D _77381_/A sky130_fd_sc_hd__nand2_4
X_43772_ _43802_/A _43772_/X sky130_fd_sc_hd__buf_2
X_55758_ _55192_/A _85159_/Q _55758_/X sky130_fd_sc_hd__and2_4
X_86578_ _86578_/CLK _47997_/Y _73927_/B sky130_fd_sc_hd__dfxtp_4
X_74592_ _74591_/X _74583_/X _56102_/X _74584_/X _74592_/X sky130_fd_sc_hd__a211o_4
X_40984_ _40937_/A _40984_/B _40984_/X sky130_fd_sc_hd__or2_4
Xclkbuf_8_124_0_CLK clkbuf_7_62_0_CLK/X clkbuf_8_124_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_45511_ _45668_/A _45511_/X sky130_fd_sc_hd__buf_2
X_76331_ _76332_/A _81563_/Q _76331_/Y sky130_fd_sc_hd__nor2_4
X_88317_ _88326_/CLK _40887_/Y _69865_/B sky130_fd_sc_hd__dfxtp_4
X_42723_ _42723_/A _42723_/X sky130_fd_sc_hd__buf_2
X_54709_ _54718_/A _47385_/Y _54709_/Y sky130_fd_sc_hd__nand2_4
X_73543_ _48704_/Y _73543_/B _73543_/X sky130_fd_sc_hd__xor2_4
X_85529_ _85529_/CLK _53984_/Y _85529_/Q sky130_fd_sc_hd__dfxtp_4
X_46491_ _46491_/A _50832_/B _46491_/Y sky130_fd_sc_hd__nand2_4
X_70755_ _70755_/A _70727_/A _70755_/Y sky130_fd_sc_hd__nand2_4
X_58477_ _64422_/C _58478_/A sky130_fd_sc_hd__buf_2
X_55689_ _55689_/A _55690_/A sky130_fd_sc_hd__buf_2
X_48230_ _48225_/Y _48226_/X _48229_/Y _86552_/D sky130_fd_sc_hd__a21boi_4
X_79050_ _82653_/Q _79053_/B sky130_fd_sc_hd__inv_2
X_45442_ _85022_/Q _55596_/B sky130_fd_sc_hd__inv_2
X_57428_ _57408_/X _57426_/X _57427_/Y _57429_/A sky130_fd_sc_hd__o21ai_4
X_76262_ _76260_/X _81642_/Q _76262_/Y sky130_fd_sc_hd__nand2_4
X_88248_ _88247_/CLK _41265_/X _88248_/Q sky130_fd_sc_hd__dfxtp_4
X_42654_ _40982_/X _42652_/X _87786_/Q _42653_/X _42654_/X sky130_fd_sc_hd__a2bb2o_4
X_73474_ _73355_/X _85573_/Q _73472_/X _73473_/X _73474_/X sky130_fd_sc_hd__a211o_4
X_70686_ _71411_/A _70692_/B _70692_/C _70686_/Y sky130_fd_sc_hd__nor3_4
X_78001_ _77993_/A _77993_/B _78000_/Y _78001_/Y sky130_fd_sc_hd__o21ai_4
X_75213_ _80684_/Q _80984_/Q _75214_/B sky130_fd_sc_hd__xor2_4
Xclkbuf_9_240_0_CLK clkbuf_8_120_0_CLK/X clkbuf_9_240_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_41605_ _41603_/X _40530_/B _41604_/X _41605_/X sky130_fd_sc_hd__o21a_4
X_72425_ _72421_/Y _72424_/Y _72344_/X _72425_/X sky130_fd_sc_hd__a21o_4
X_48161_ _48155_/Y _48156_/X _48160_/X _86562_/D sky130_fd_sc_hd__a21oi_4
X_45373_ _55736_/B _45354_/X _45311_/X _45373_/X sky130_fd_sc_hd__o21a_4
X_57359_ _57359_/A _85029_/Q _57249_/X _57359_/Y sky130_fd_sc_hd__nor3_4
X_76193_ _76193_/A _76188_/X _76193_/C _76196_/B sky130_fd_sc_hd__nand3_4
X_88179_ _87926_/CLK _88179_/D _67349_/B sky130_fd_sc_hd__dfxtp_4
X_42585_ _42573_/X _42574_/X _40849_/X _87811_/Q _42580_/X _42585_/Y
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_8_139_0_CLK clkbuf_7_69_0_CLK/X clkbuf_9_278_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_47112_ _54553_/D _52861_/D sky130_fd_sc_hd__buf_2
Xclkbuf_10_134_0_CLK clkbuf_9_67_0_CLK/X _83820_/CLK sky130_fd_sc_hd__clkbuf_1
X_44324_ _41643_/X _40543_/X _87165_/Q _40544_/X _87165_/D sky130_fd_sc_hd__a2bb2o_4
X_75144_ _75141_/X _75145_/C _75143_/Y _75144_/Y sky130_fd_sc_hd__a21oi_4
X_41536_ _41535_/X _41536_/X sky130_fd_sc_hd__buf_2
X_48092_ _48092_/A _50358_/B _48092_/Y sky130_fd_sc_hd__nand2_4
X_60370_ _60369_/X _60370_/Y sky130_fd_sc_hd__inv_2
X_72356_ _83262_/Q _72250_/X _72349_/X _72355_/X _83262_/D sky130_fd_sc_hd__a2bb2oi_4
Xclkbuf_10_764_0_CLK clkbuf_9_382_0_CLK/X _88044_/CLK sky130_fd_sc_hd__clkbuf_1
X_47043_ _47008_/A _51130_/B _47043_/Y sky130_fd_sc_hd__nand2_4
X_59029_ _59029_/A _86366_/Q _59029_/Y sky130_fd_sc_hd__nor2_4
X_71307_ _52036_/B _71290_/X _71306_/Y _71307_/Y sky130_fd_sc_hd__o21ai_4
X_44255_ _45950_/A _44227_/Y _44210_/X _43972_/B _44254_/X _44255_/X
+ sky130_fd_sc_hd__o32a_4
X_75075_ _75072_/Y _75074_/B _75076_/B _75075_/Y sky130_fd_sc_hd__a21oi_4
X_79952_ _84926_/Q _84174_/Q _79952_/X sky130_fd_sc_hd__or2_4
X_41467_ _81183_/Q _41459_/B _41467_/X sky130_fd_sc_hd__or2_4
X_72287_ _57711_/X _72287_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_255_0_CLK clkbuf_9_255_0_CLK/A clkbuf_9_255_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_43206_ _40939_/X _43180_/X _87538_/Q _43185_/X _43206_/X sky130_fd_sc_hd__a2bb2o_4
X_74026_ _53552_/B _74026_/B _74026_/X sky130_fd_sc_hd__xor2_4
X_62040_ _63611_/A _59825_/B _61572_/A _61981_/X _62040_/X sky130_fd_sc_hd__a2bb2o_4
X_78903_ _82845_/Q _78903_/B _78903_/Y sky130_fd_sc_hd__xnor2_4
X_40418_ _40417_/Y _40418_/X sky130_fd_sc_hd__buf_2
X_71238_ _71137_/A _71238_/B _71239_/A sky130_fd_sc_hd__nor2_4
X_44186_ _44186_/A _44185_/X _44186_/X sky130_fd_sc_hd__or2_4
X_79883_ _60214_/C _79883_/B _79883_/X sky130_fd_sc_hd__xor2_4
X_41398_ _41397_/X _41362_/X _67848_/B _41363_/X _88222_/D sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_10_149_0_CLK clkbuf_9_74_0_CLK/X _81696_/CLK sky130_fd_sc_hd__clkbuf_1
X_43137_ _43137_/A _43137_/Y sky130_fd_sc_hd__inv_2
X_78834_ _78841_/B _78833_/Y _78834_/X sky130_fd_sc_hd__xor2_4
X_40349_ _41869_/A _42447_/A sky130_fd_sc_hd__inv_2
X_71169_ _52137_/B _71165_/X _71168_/Y _71169_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_779_0_CLK clkbuf_9_389_0_CLK/X _82575_/CLK sky130_fd_sc_hd__clkbuf_1
X_48994_ _86454_/Q _48952_/X _48993_/Y _48994_/Y sky130_fd_sc_hd__o21ai_4
X_47945_ _51988_/A _48234_/A sky130_fd_sc_hd__buf_2
X_43068_ _43068_/A _43068_/Y sky130_fd_sc_hd__inv_2
X_78765_ _78761_/X _78762_/A _78765_/Y sky130_fd_sc_hd__nand2_4
X_63991_ _63734_/A _64053_/A sky130_fd_sc_hd__buf_2
X_75977_ _75969_/B _75977_/B _75977_/Y sky130_fd_sc_hd__nor2_4
X_42019_ _42018_/Y _88069_/D sky130_fd_sc_hd__inv_2
X_65730_ _65134_/X _65653_/B _65138_/X _65742_/A sky130_fd_sc_hd__nand3_4
X_77716_ _82125_/Q _77716_/B _77717_/A sky130_fd_sc_hd__xor2_4
X_62942_ _62893_/A _62942_/X sky130_fd_sc_hd__buf_2
X_74928_ _81134_/D _74928_/B _74942_/A sky130_fd_sc_hd__xor2_4
X_47876_ _47918_/A _47877_/A sky130_fd_sc_hd__buf_2
X_78696_ _78695_/X _78696_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_702_0_CLK clkbuf_9_351_0_CLK/X _87126_/CLK sky130_fd_sc_hd__clkbuf_1
X_49615_ _49610_/A _49614_/X _49615_/C _52831_/D _49615_/X sky130_fd_sc_hd__and4_4
X_46827_ _58853_/A _46813_/X _46826_/Y _46827_/Y sky130_fd_sc_hd__o21ai_4
X_65661_ _65769_/A _86514_/Q _65661_/X sky130_fd_sc_hd__and2_4
X_77647_ _77648_/A _77648_/C _81949_/Q _77650_/A sky130_fd_sc_hd__a21oi_4
X_62873_ _62894_/A _62852_/X _62873_/C _62873_/Y sky130_fd_sc_hd__nor3_4
X_74859_ _81123_/D _80835_/Q _74859_/Y sky130_fd_sc_hd__nand2_4
X_67400_ _86973_/Q _67348_/X _67398_/X _67399_/X _67400_/X sky130_fd_sc_hd__a211o_4
X_64612_ _64564_/X _86144_/Q _64566_/X _64611_/X _64612_/X sky130_fd_sc_hd__a211o_4
X_49546_ _49546_/A _52760_/B _49546_/Y sky130_fd_sc_hd__nand2_4
X_61824_ _61728_/A _61824_/X sky130_fd_sc_hd__buf_2
X_68380_ _68380_/A _68380_/Y sky130_fd_sc_hd__inv_2
X_46758_ _52658_/B _46758_/X sky130_fd_sc_hd__buf_2
X_65592_ _65592_/A _86486_/Q _65592_/X sky130_fd_sc_hd__and2_4
X_77578_ _77578_/A _77577_/Y _82201_/D sky130_fd_sc_hd__xor2_4
X_67331_ _67806_/A _67331_/X sky130_fd_sc_hd__buf_2
X_79317_ _79334_/B _79316_/Y _82830_/D sky130_fd_sc_hd__xor2_4
X_45709_ _45709_/A _45709_/X sky130_fd_sc_hd__buf_2
X_64543_ _58370_/A _64521_/X _64543_/Y sky130_fd_sc_hd__nor2_4
X_76529_ _76584_/A _76529_/B _81627_/D sky130_fd_sc_hd__xnor2_4
X_49477_ _58830_/B _49470_/X _49476_/Y _49477_/Y sky130_fd_sc_hd__o21ai_4
X_61755_ _61755_/A _61755_/X sky130_fd_sc_hd__buf_2
X_46689_ _46688_/Y _51787_/D sky130_fd_sc_hd__buf_2
Xclkbuf_10_717_0_CLK clkbuf_9_358_0_CLK/X _88263_/CLK sky130_fd_sc_hd__clkbuf_1
X_48428_ _48372_/X _82363_/Q _48427_/Y _74396_/A sky130_fd_sc_hd__o21ai_4
X_60706_ _60359_/X _60704_/Y _60694_/Y _60696_/Y _60705_/Y _60706_/Y
+ sky130_fd_sc_hd__a41oi_4
X_67262_ _67308_/A _86809_/Q _67262_/X sky130_fd_sc_hd__and2_4
X_79248_ _79246_/Y _79229_/Y _79248_/C _79248_/Y sky130_fd_sc_hd__nand3_4
X_64474_ _64474_/A _64474_/X sky130_fd_sc_hd__buf_2
X_61686_ _61686_/A _72555_/B sky130_fd_sc_hd__buf_2
Xclkbuf_9_208_0_CLK clkbuf_8_104_0_CLK/X clkbuf_9_208_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_69001_ _69001_/A _42528_/Y _69001_/Y sky130_fd_sc_hd__nor2_4
X_66213_ _66210_/X _66212_/X _65304_/X _66216_/A sky130_fd_sc_hd__a21o_4
X_63425_ _58421_/A _63370_/X _61390_/A _63372_/X _63425_/X sky130_fd_sc_hd__a2bb2o_4
X_48359_ _48392_/A _48358_/X _48359_/Y sky130_fd_sc_hd__nand2_4
X_60637_ _60637_/A _60642_/A sky130_fd_sc_hd__buf_2
X_67193_ _66953_/X _67193_/X sky130_fd_sc_hd__buf_2
X_79179_ _79175_/Y _79165_/Y _79173_/Y _79189_/A sky130_fd_sc_hd__a21oi_4
X_81210_ _84111_/CLK _75078_/Y _48959_/A sky130_fd_sc_hd__dfxtp_4
X_66144_ _64722_/X _85617_/Q _64724_/X _66143_/X _66144_/X sky130_fd_sc_hd__a211o_4
X_51370_ _51364_/A _50858_/B _51370_/Y sky130_fd_sc_hd__nand2_4
X_63356_ _60677_/A _63632_/A _60702_/C _63356_/X sky130_fd_sc_hd__and3_4
X_82190_ _84945_/CLK _82190_/D _82190_/Q sky130_fd_sc_hd__dfxtp_4
X_60568_ _60612_/A _60526_/B _79138_/A _60568_/Y sky130_fd_sc_hd__nor3_4
X_50321_ _50572_/A _50356_/A sky130_fd_sc_hd__buf_2
X_62307_ _61406_/A _62247_/X _62259_/X _62631_/D _62307_/Y sky130_fd_sc_hd__nand4_4
X_81141_ _86758_/CLK _81141_/D _40654_/A sky130_fd_sc_hd__dfxtp_4
X_66075_ _65308_/X _84982_/Q _65309_/X _66074_/X _66075_/X sky130_fd_sc_hd__a211o_4
X_63287_ _59427_/Y _63259_/X _63234_/X _58973_/A _63235_/X _63287_/Y
+ sky130_fd_sc_hd__o32ai_4
X_60499_ _60387_/A _60392_/A _60392_/C _60387_/C _60383_/A _60566_/A
+ sky130_fd_sc_hd__a41oi_4
X_53040_ _53147_/A _53040_/X sky130_fd_sc_hd__buf_2
X_65026_ _64846_/X _85521_/Q _64919_/X _65025_/X _65026_/X sky130_fd_sc_hd__a211o_4
X_69903_ _69484_/X _69487_/X _69816_/X _69903_/Y sky130_fd_sc_hd__a21oi_4
X_50252_ _50251_/X _51954_/B _50252_/Y sky130_fd_sc_hd__nand2_4
X_62238_ _62597_/B _61744_/X _62237_/X _62515_/C _62238_/X sky130_fd_sc_hd__and4_4
X_81072_ _81038_/CLK _81104_/Q _75267_/A sky130_fd_sc_hd__dfxtp_4
X_80023_ _80023_/A _80023_/B _80023_/Y sky130_fd_sc_hd__xnor2_4
X_84900_ _84727_/CLK _58239_/Y _84900_/Q sky130_fd_sc_hd__dfxtp_4
X_69834_ _87807_/Q _69835_/B sky130_fd_sc_hd__inv_2
Xclkbuf_4_8_0_CLK clkbuf_4_9_0_CLK/A clkbuf_4_8_1_CLK/A sky130_fd_sc_hd__clkbuf_1
X_50183_ _50131_/A _50183_/B _50183_/X sky130_fd_sc_hd__and2_4
X_62169_ _62065_/B _62063_/X _63703_/B _62183_/D _62169_/X sky130_fd_sc_hd__and4_4
X_85880_ _85879_/CLK _85880_/D _85880_/Q sky130_fd_sc_hd__dfxtp_4
X_84831_ _84960_/CLK _58512_/Y _64335_/C sky130_fd_sc_hd__dfxtp_4
X_69765_ _87556_/Q _69747_/X _68348_/X _69764_/X _69765_/X sky130_fd_sc_hd__a211o_4
X_54991_ _54888_/A _55013_/A sky130_fd_sc_hd__buf_2
X_66977_ _66974_/X _66976_/X _66905_/X _66977_/X sky130_fd_sc_hd__a21o_4
X_56730_ _56729_/X _56730_/X sky130_fd_sc_hd__buf_2
X_68716_ _68542_/X _87749_/Q _68716_/X sky130_fd_sc_hd__and2_4
X_87550_ _87820_/CLK _43171_/Y _43170_/A sky130_fd_sc_hd__dfxtp_4
X_53942_ _53942_/A _46242_/Y _53942_/Y sky130_fd_sc_hd__nand2_4
X_65928_ _65928_/A _65927_/Y _65928_/Y sky130_fd_sc_hd__nand2_4
X_84762_ _85485_/CLK _84762_/D _84762_/Q sky130_fd_sc_hd__dfxtp_4
X_69696_ _69696_/A _69696_/X sky130_fd_sc_hd__buf_2
X_81974_ _82234_/CLK _83902_/Q _81974_/Q sky130_fd_sc_hd__dfxtp_4
X_86501_ _86499_/CLK _48681_/Y _86501_/Q sky130_fd_sc_hd__dfxtp_4
X_83713_ _86303_/CLK _70741_/Y _47526_/A sky130_fd_sc_hd__dfxtp_4
X_80925_ _80928_/CLK _84101_/Q _80925_/Q sky130_fd_sc_hd__dfxtp_4
X_56661_ _56651_/Y _56655_/Y _56661_/C _56661_/Y sky130_fd_sc_hd__nor3_4
X_68647_ _68647_/A _68646_/X _68647_/Y sky130_fd_sc_hd__nand2_4
X_87481_ _87993_/CLK _87481_/D _87481_/Q sky130_fd_sc_hd__dfxtp_4
X_53873_ _85551_/Q _53869_/X _53872_/Y _53873_/Y sky130_fd_sc_hd__o21ai_4
X_65859_ _65859_/A _65859_/X sky130_fd_sc_hd__buf_2
X_84693_ _84713_/CLK _84693_/D _80413_/A sky130_fd_sc_hd__dfxtp_4
X_58400_ _58400_/A _58403_/B _58400_/Y sky130_fd_sc_hd__nand2_4
X_55612_ _55607_/A _45425_/Y _55612_/Y sky130_fd_sc_hd__nor2_4
X_86432_ _85535_/CLK _49217_/Y _86432_/Q sky130_fd_sc_hd__dfxtp_4
X_52824_ _85748_/Q _52821_/X _52823_/Y _52824_/Y sky130_fd_sc_hd__o21ai_4
X_59380_ _59331_/X _85410_/Q _59379_/X _59380_/Y sky130_fd_sc_hd__o21ai_4
X_83644_ _86422_/CLK _83644_/D _83644_/Q sky130_fd_sc_hd__dfxtp_4
X_56592_ _46233_/Y _56593_/A sky130_fd_sc_hd__buf_2
X_80856_ _80740_/CLK _80888_/Q _75020_/C sky130_fd_sc_hd__dfxtp_4
X_68578_ _87499_/Q _68504_/X _68450_/X _68577_/X _68578_/X sky130_fd_sc_hd__a211o_4
X_58331_ _58331_/A _58364_/B _58331_/Y sky130_fd_sc_hd__nand2_4
X_55543_ _85113_/Q _55510_/X _44048_/X _55542_/Y _55543_/X sky130_fd_sc_hd__a211o_4
X_67529_ _67526_/X _67528_/X _67502_/X _67532_/A sky130_fd_sc_hd__a21o_4
X_86363_ _83049_/CLK _86363_/D _86363_/Q sky130_fd_sc_hd__dfxtp_4
X_52755_ _52783_/A _52755_/X sky130_fd_sc_hd__buf_2
X_83575_ _86505_/CLK _71200_/Y _48559_/A sky130_fd_sc_hd__dfxtp_4
X_80787_ _80754_/CLK _80787_/D _75329_/A sky130_fd_sc_hd__dfxtp_4
X_88102_ _88108_/CLK _41930_/Y _88102_/Q sky130_fd_sc_hd__dfxtp_4
X_85314_ _85346_/CLK _85314_/D _85314_/Q sky130_fd_sc_hd__dfxtp_4
X_51706_ _51704_/Y _51693_/X _51705_/X _51706_/Y sky130_fd_sc_hd__a21oi_4
X_70540_ _71215_/C _70550_/D sky130_fd_sc_hd__buf_2
X_58262_ _58261_/Y _58268_/B _58262_/Y sky130_fd_sc_hd__nand2_4
X_82526_ _82624_/CLK _79090_/Y _78748_/A sky130_fd_sc_hd__dfxtp_4
X_55474_ _55471_/X _55473_/X _44112_/X _55474_/X sky130_fd_sc_hd__a21o_4
X_86294_ _86611_/CLK _49948_/Y _72251_/B sky130_fd_sc_hd__dfxtp_4
X_52686_ _52706_/A _52686_/B _52686_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_1021_0_CLK clkbuf_9_510_0_CLK/X _86499_/CLK sky130_fd_sc_hd__clkbuf_1
X_57213_ _57096_/Y _57209_/Y _57210_/Y _57212_/Y _57214_/A sky130_fd_sc_hd__a211o_4
X_88033_ _88036_/CLK _88033_/D _88033_/Q sky130_fd_sc_hd__dfxtp_4
X_54425_ _54425_/A _52732_/B _54425_/Y sky130_fd_sc_hd__nand2_4
X_85245_ _85244_/CLK _85245_/D _85245_/Q sky130_fd_sc_hd__dfxtp_4
X_51637_ _51627_/A _53161_/B _51637_/Y sky130_fd_sc_hd__nand2_4
X_70471_ _70466_/Y _83768_/Q _70470_/X _70471_/X sky130_fd_sc_hd__a21o_4
X_58193_ _62124_/B _58194_/A sky130_fd_sc_hd__buf_2
X_82457_ _82425_/CLK _79149_/X _82457_/Q sky130_fd_sc_hd__dfxtp_4
X_72210_ _72123_/X _85690_/Q _72146_/X _72210_/X sky130_fd_sc_hd__o21a_4
X_57144_ _57142_/X _57143_/X _45835_/A _57144_/X sky130_fd_sc_hd__a21o_4
X_81408_ _81351_/CLK _83944_/Q _76773_/B sky130_fd_sc_hd__dfxtp_4
X_54356_ _85457_/Q _54349_/X _54355_/Y _54356_/Y sky130_fd_sc_hd__o21ai_4
X_42370_ _41872_/A _42370_/X sky130_fd_sc_hd__buf_2
X_73190_ _73180_/Y _73189_/X _73190_/X sky130_fd_sc_hd__xor2_4
X_85176_ _85270_/CLK _85176_/D _85176_/Q sky130_fd_sc_hd__dfxtp_4
X_51568_ _51590_/A _53095_/B _51568_/Y sky130_fd_sc_hd__nand2_4
X_82388_ _85491_/CLK _82196_/Q _47046_/A sky130_fd_sc_hd__dfxtp_4
X_41321_ _41320_/X _41321_/X sky130_fd_sc_hd__buf_2
X_53307_ _53293_/A _53293_/B _53302_/X _52790_/D _53307_/X sky130_fd_sc_hd__and4_4
X_72141_ _72417_/A _72141_/X sky130_fd_sc_hd__buf_2
X_84127_ _84166_/CLK _84127_/D _66420_/C sky130_fd_sc_hd__dfxtp_4
X_50519_ _48841_/A _50526_/B _50526_/C _50519_/X sky130_fd_sc_hd__and3_4
X_57075_ _57075_/A _57075_/Y sky130_fd_sc_hd__inv_2
X_81339_ _81575_/CLK _81339_/D _81339_/Q sky130_fd_sc_hd__dfxtp_4
X_54287_ _54282_/Y _54285_/X _54286_/X _54287_/Y sky130_fd_sc_hd__a21oi_4
X_51499_ _51509_/A _51494_/B _51522_/C _53023_/D _51499_/X sky130_fd_sc_hd__and4_4
X_44040_ _60371_/A _44031_/X _57811_/A _59297_/A _44039_/X _44160_/A
+ sky130_fd_sc_hd__a41oi_4
X_56026_ _56025_/X _56026_/X sky130_fd_sc_hd__buf_2
X_41252_ _40755_/A _41253_/A sky130_fd_sc_hd__buf_2
X_53238_ _53217_/A _53244_/B _53222_/X _53238_/D _53238_/X sky130_fd_sc_hd__and4_4
X_72072_ _72053_/A _72072_/B _72072_/Y sky130_fd_sc_hd__nand2_4
X_84058_ _81461_/CLK _67712_/X _81490_/D sky130_fd_sc_hd__dfxtp_4
X_71023_ _70771_/A _71173_/A sky130_fd_sc_hd__buf_2
X_75900_ _61250_/C _62921_/C _75900_/X sky130_fd_sc_hd__xor2_4
X_83009_ _85075_/CLK _83009_/D _83009_/Q sky130_fd_sc_hd__dfxtp_4
X_41183_ _41179_/X _41181_/X _68708_/B _41182_/X _41183_/X sky130_fd_sc_hd__a2bb2o_4
X_53169_ _53195_/A _53169_/X sky130_fd_sc_hd__buf_2
X_76880_ _76874_/Y _76873_/Y _76881_/C sky130_fd_sc_hd__nand2_4
X_75831_ _75831_/A _75836_/A sky130_fd_sc_hd__inv_2
X_87817_ _88326_/CLK _42567_/Y _87817_/Q sky130_fd_sc_hd__dfxtp_4
X_45991_ _45991_/A _45991_/Y sky130_fd_sc_hd__inv_2
X_57977_ _57939_/X _85999_/Q _57976_/X _57977_/Y sky130_fd_sc_hd__o21ai_4
X_47730_ _47729_/Y _53211_/D sky130_fd_sc_hd__buf_2
X_59716_ _59716_/A _59716_/B _60132_/A _59716_/Y sky130_fd_sc_hd__nand3_4
X_78550_ _78549_/A _82675_/D _78551_/A sky130_fd_sc_hd__nand2_4
X_44942_ _44931_/X _44939_/X _44941_/Y _44942_/Y sky130_fd_sc_hd__a21oi_4
X_56928_ _44137_/A _56923_/Y _56927_/Y _56928_/Y sky130_fd_sc_hd__o21ai_4
X_75762_ _81095_/Q _80807_/Q _75762_/Y sky130_fd_sc_hd__xnor2_4
X_87748_ _87748_/CLK _87748_/D _68755_/B sky130_fd_sc_hd__dfxtp_4
X_72974_ _72722_/X _72974_/X sky130_fd_sc_hd__buf_2
X_77501_ _77465_/B _77498_/X _77500_/Y _77501_/Y sky130_fd_sc_hd__a21oi_4
X_74713_ MACRO_RD_SELECT _74713_/Y sky130_fd_sc_hd__inv_2
X_47661_ _47661_/A _47692_/C sky130_fd_sc_hd__buf_2
X_71925_ _70591_/A _71940_/C sky130_fd_sc_hd__buf_2
X_59647_ _59824_/B _59649_/A sky130_fd_sc_hd__buf_2
X_78481_ _78476_/Y _78453_/B _78480_/X _78482_/B sky130_fd_sc_hd__o21ai_4
X_44873_ _45193_/A _45197_/A sky130_fd_sc_hd__buf_2
X_56859_ _83333_/Q _56859_/X sky130_fd_sc_hd__buf_2
X_87679_ _87686_/CLK _42865_/Y _67047_/B sky130_fd_sc_hd__dfxtp_4
X_75693_ _81007_/Q _75693_/B _75693_/X sky130_fd_sc_hd__xor2_4
X_49400_ _86394_/Q _49388_/X _49399_/Y _49400_/Y sky130_fd_sc_hd__o21ai_4
X_46612_ _46612_/A _53097_/A sky130_fd_sc_hd__buf_2
X_77432_ _77430_/X _77431_/Y _77433_/A sky130_fd_sc_hd__and2_4
X_43824_ _43854_/A _43824_/X sky130_fd_sc_hd__buf_2
X_74644_ _56600_/A _74641_/X _74643_/Y _83003_/D sky130_fd_sc_hd__a21boi_4
X_47592_ _86618_/Q _47570_/X _47591_/Y _47592_/Y sky130_fd_sc_hd__o21ai_4
X_71856_ _71848_/X _83352_/Q _71855_/Y _83352_/D sky130_fd_sc_hd__a21o_4
X_59578_ _59577_/X _59579_/A sky130_fd_sc_hd__buf_2
X_49331_ _86408_/Q _49285_/X _49330_/Y _49331_/Y sky130_fd_sc_hd__o21ai_4
X_46543_ _46542_/X _46543_/X sky130_fd_sc_hd__buf_2
X_70807_ _70810_/A _70940_/B _70810_/C _70807_/Y sky130_fd_sc_hd__nand3_4
X_58529_ _58517_/X _58526_/Y _58528_/Y _84827_/D sky130_fd_sc_hd__a21oi_4
X_77363_ _77351_/B _77345_/A _77345_/B _77363_/Y sky130_fd_sc_hd__a21boi_4
X_43755_ _43591_/A _43756_/A sky130_fd_sc_hd__inv_2
X_74575_ _56863_/X _74575_/X sky130_fd_sc_hd__buf_2
X_40967_ _40931_/X _81723_/Q _40966_/X _40968_/A sky130_fd_sc_hd__o21ai_4
X_71787_ _58181_/Y _71784_/X _71786_/Y _83377_/D sky130_fd_sc_hd__o21ai_4
X_79102_ _79101_/Y _79086_/A _79102_/X sky130_fd_sc_hd__and2_4
X_76314_ _76314_/A _76316_/A sky130_fd_sc_hd__inv_2
X_42706_ _41130_/X _42695_/X _87760_/Q _42696_/X _42706_/X sky130_fd_sc_hd__a2bb2o_4
X_49262_ _86422_/Q _49255_/X _49261_/Y _49262_/Y sky130_fd_sc_hd__o21ai_4
X_73526_ _83147_/Q _73437_/X _73525_/Y _83147_/D sky130_fd_sc_hd__a21o_4
X_61540_ _84864_/Q _61541_/B sky130_fd_sc_hd__buf_2
X_46474_ _46719_/A _46474_/X sky130_fd_sc_hd__buf_2
X_70738_ _70755_/A _70738_/X sky130_fd_sc_hd__buf_2
X_77294_ _77294_/A _77294_/B _77294_/Y sky130_fd_sc_hd__nand2_4
X_43686_ _43673_/A _43686_/X sky130_fd_sc_hd__buf_2
X_40898_ _40817_/X _82280_/Q _40897_/X _40898_/Y sky130_fd_sc_hd__o21ai_4
X_48213_ _48184_/A _53488_/B _48213_/Y sky130_fd_sc_hd__nand2_4
X_79033_ _79027_/B _79027_/A _79032_/X _79033_/Y sky130_fd_sc_hd__a21oi_4
X_45425_ _85023_/Q _45425_/Y sky130_fd_sc_hd__inv_2
X_76245_ _81257_/Q _81513_/D _76245_/Y sky130_fd_sc_hd__nor2_4
X_42637_ _42580_/A _42637_/X sky130_fd_sc_hd__buf_2
X_49193_ _49173_/A _50719_/B _49193_/X sky130_fd_sc_hd__and2_4
X_61471_ _59403_/A _61484_/B _61484_/C _61452_/D _61471_/Y sky130_fd_sc_hd__nand4_4
X_73457_ _73457_/A _73456_/X _73457_/Y sky130_fd_sc_hd__nand2_4
X_70669_ _70669_/A _70676_/C sky130_fd_sc_hd__buf_2
X_63210_ _63207_/Y _63209_/X _63172_/X _63210_/Y sky130_fd_sc_hd__a21oi_4
X_60422_ _60422_/A _60513_/B sky130_fd_sc_hd__buf_2
X_48144_ _48144_/A _50105_/A sky130_fd_sc_hd__buf_2
X_72408_ _72305_/X _85353_/Q _72407_/X _72408_/Y sky130_fd_sc_hd__o21ai_4
X_45356_ _56270_/C _45297_/X _45355_/X _45356_/Y sky130_fd_sc_hd__o21ai_4
X_76176_ _76176_/A _76176_/Y sky130_fd_sc_hd__inv_2
X_64190_ _64190_/A _64190_/B _64189_/D _64190_/D _64190_/Y sky130_fd_sc_hd__nand4_4
X_42568_ _42554_/A _42568_/X sky130_fd_sc_hd__buf_2
X_73388_ _73384_/X _73387_/X _73388_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_194_0_CLK clkbuf_8_97_0_CLK/X clkbuf_9_194_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_44307_ _44120_/Y _44010_/A _74095_/B _44307_/D _44308_/A sky130_fd_sc_hd__and4_4
X_63141_ _79394_/A _63130_/X _63140_/Y _63141_/X sky130_fd_sc_hd__a21o_4
X_75127_ _75124_/X _81062_/Q _75127_/C _75143_/A sky130_fd_sc_hd__nand3_4
X_41519_ _41421_/X _82325_/Q _41518_/X _41519_/X sky130_fd_sc_hd__o21a_4
X_48075_ _48914_/A _48075_/X sky130_fd_sc_hd__buf_2
X_60353_ _60414_/B _60353_/B _59716_/B _60353_/Y sky130_fd_sc_hd__nand3_4
X_72339_ _59345_/X _72339_/X sky130_fd_sc_hd__buf_2
X_45287_ _45212_/A _45287_/X sky130_fd_sc_hd__buf_2
X_42499_ _42499_/A _68746_/B sky130_fd_sc_hd__inv_2
X_47026_ _59131_/A _47004_/X _47025_/Y _47026_/Y sky130_fd_sc_hd__o21ai_4
X_44238_ _57126_/A _44239_/A sky130_fd_sc_hd__buf_2
X_63072_ _63130_/A _63072_/X sky130_fd_sc_hd__buf_2
X_75058_ _75053_/B _75056_/X _75057_/Y _75059_/B sky130_fd_sc_hd__a21boi_4
X_79935_ _79937_/B _79935_/Y sky130_fd_sc_hd__inv_2
X_60284_ _60284_/A _60284_/B _60300_/C _60284_/Y sky130_fd_sc_hd__nand3_4
X_66900_ _66851_/X _66900_/B _66900_/X sky130_fd_sc_hd__and2_4
X_62023_ _63598_/A _59841_/X _61561_/A _61981_/X _62023_/X sky130_fd_sc_hd__a2bb2o_4
X_74009_ _74006_/X _74008_/X _73944_/X _74028_/B sky130_fd_sc_hd__a21o_4
X_44169_ _44244_/A _44170_/A sky130_fd_sc_hd__buf_2
X_67880_ _67901_/A _87644_/Q _67880_/X sky130_fd_sc_hd__and2_4
X_79866_ _79844_/X _79866_/B _79866_/X sky130_fd_sc_hd__or2_4
X_66831_ _87432_/Q _66762_/X _66764_/X _66830_/X _66831_/X sky130_fd_sc_hd__a211o_4
X_78817_ _78816_/Y _78817_/Y sky130_fd_sc_hd__inv_2
X_48977_ _48606_/X _81208_/Q _48976_/Y _48978_/A sky130_fd_sc_hd__o21ai_4
X_79797_ _79797_/A _79797_/B _79798_/B sky130_fd_sc_hd__xor2_4
Xclkbuf_10_641_0_CLK clkbuf_9_320_0_CLK/X _86934_/CLK sky130_fd_sc_hd__clkbuf_1
X_69550_ _69102_/X _69105_/X _69500_/X _69550_/Y sky130_fd_sc_hd__a21oi_4
X_47928_ _47887_/A _48221_/A _47928_/X sky130_fd_sc_hd__and2_4
X_66762_ _66642_/A _66762_/X sky130_fd_sc_hd__buf_2
X_78748_ _78748_/A _82782_/D _82494_/D sky130_fd_sc_hd__xor2_4
X_63974_ _63942_/A _59415_/A _63958_/C _63974_/X sky130_fd_sc_hd__and3_4
X_68501_ _68651_/A _68501_/X sky130_fd_sc_hd__buf_2
X_65713_ _65621_/A _65775_/B _65713_/C _65713_/X sky130_fd_sc_hd__and3_4
Xclkbuf_9_132_0_CLK clkbuf_8_66_0_CLK/X clkbuf_9_132_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_62925_ _62646_/B _62926_/B sky130_fd_sc_hd__buf_2
X_69481_ _88026_/Q _69368_/X _69478_/X _69480_/X _69481_/X sky130_fd_sc_hd__a211o_4
X_47859_ _82367_/Q _46579_/X _47859_/X sky130_fd_sc_hd__or2_4
X_66693_ _66690_/X _66692_/X _66667_/X _66693_/X sky130_fd_sc_hd__a21o_4
X_78679_ _78680_/A _78680_/B _78682_/B sky130_fd_sc_hd__nor2_4
X_68432_ _87101_/Q _68059_/X _68370_/X _68431_/X _68432_/X sky130_fd_sc_hd__a211o_4
X_80710_ _80679_/CLK _75896_/X _80710_/Q sky130_fd_sc_hd__dfxtp_4
X_65644_ _65474_/X _86515_/Q _65644_/X sky130_fd_sc_hd__and2_4
X_50870_ _50857_/X _50870_/B _50870_/Y sky130_fd_sc_hd__nand2_4
X_62856_ _63573_/A _60337_/D _62855_/Y _62856_/X sky130_fd_sc_hd__o21a_4
X_81690_ _81689_/CLK _80182_/X _81690_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_656_0_CLK clkbuf_9_328_0_CLK/X _87926_/CLK sky130_fd_sc_hd__clkbuf_1
X_61807_ _58237_/X _61728_/X _61756_/X _61790_/X _61806_/X _61807_/X
+ sky130_fd_sc_hd__a41o_4
X_49529_ _49527_/Y _49514_/X _49528_/X _49529_/Y sky130_fd_sc_hd__a21oi_4
X_80641_ _80641_/HI THREAD_COUNT[0] sky130_fd_sc_hd__conb_1
X_68363_ _73552_/A _68006_/X _68359_/X _68362_/Y _68363_/X sky130_fd_sc_hd__a211o_4
X_65575_ _64885_/X _65548_/B _64887_/X _65587_/A sky130_fd_sc_hd__nand3_4
X_62787_ _61461_/X _62743_/B _62742_/X _62834_/D _62787_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_9_147_0_CLK clkbuf_8_73_0_CLK/X clkbuf_9_147_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_67314_ _67266_/A _88116_/Q _67314_/X sky130_fd_sc_hd__and2_4
X_52540_ _65234_/B _52500_/X _52539_/Y _52540_/Y sky130_fd_sc_hd__o21ai_4
X_64526_ _64455_/X _64526_/B _61102_/X _64526_/Y sky130_fd_sc_hd__nand3_4
X_83360_ _83421_/CLK _83360_/D _83360_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_74_0_CLK clkbuf_8_37_0_CLK/X clkbuf_9_74_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_61738_ _59692_/Y _61842_/A sky130_fd_sc_hd__buf_2
X_80572_ _80550_/A _80549_/Y _80557_/X _80561_/B _80572_/X sky130_fd_sc_hd__o22a_4
X_68294_ _67013_/X _68737_/A sky130_fd_sc_hd__buf_2
XPHY_209 sky130_fd_sc_hd__decap_3
X_82311_ _82317_/CLK _77033_/B _82311_/Q sky130_fd_sc_hd__dfxtp_4
X_67245_ _67266_/A _67245_/B _67245_/X sky130_fd_sc_hd__and2_4
X_52471_ _52177_/A _52476_/A sky130_fd_sc_hd__buf_2
X_64457_ _64456_/Y _64457_/B _64457_/C _64457_/Y sky130_fd_sc_hd__nand3_4
X_83291_ _83304_/CLK _72071_/Y _83291_/Q sky130_fd_sc_hd__dfxtp_4
X_61669_ _61669_/A _61669_/Y sky130_fd_sc_hd__inv_2
X_54210_ _54206_/Y _54197_/X _54209_/X _85484_/D sky130_fd_sc_hd__a21oi_4
X_85030_ _85039_/CLK _85030_/D _45811_/A sky130_fd_sc_hd__dfxtp_4
X_51422_ _51410_/X _51421_/X _51438_/C _52948_/D _51422_/X sky130_fd_sc_hd__and4_4
X_63408_ _63403_/Y _63391_/X _63407_/Y _63408_/Y sky130_fd_sc_hd__a21oi_4
X_82242_ _84441_/CLK _80636_/Y _82242_/Q sky130_fd_sc_hd__dfxtp_4
X_55190_ _55710_/B _55190_/X sky130_fd_sc_hd__buf_2
X_67176_ _67055_/X _67176_/X sky130_fd_sc_hd__buf_2
X_64388_ _79733_/B _64373_/X _64387_/X _64388_/X sky130_fd_sc_hd__a21o_4
X_54141_ _54194_/A _54149_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_89_0_CLK clkbuf_9_88_0_CLK/A clkbuf_9_89_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_66127_ _66181_/A _85906_/Q _66127_/X sky130_fd_sc_hd__and2_4
X_51353_ _51351_/Y _51339_/X _51352_/X _86027_/D sky130_fd_sc_hd__a21oi_4
X_63339_ _59445_/A _60417_/A _60523_/A _58990_/Y _63060_/A _63339_/Y
+ sky130_fd_sc_hd__o32ai_4
X_82173_ _82047_/CLK _65970_/C _77983_/B sky130_fd_sc_hd__dfxtp_4
X_50304_ _50279_/X _48257_/B _50304_/Y sky130_fd_sc_hd__nand2_4
X_81124_ _81195_/CLK _81124_/D _81124_/Q sky130_fd_sc_hd__dfxtp_4
X_54072_ _54070_/Y _54060_/X _54071_/Y _54072_/Y sky130_fd_sc_hd__a21boi_4
X_66058_ _66051_/X _66056_/X _66057_/X _66061_/A sky130_fd_sc_hd__a21o_4
X_51284_ _51281_/Y _51263_/X _51283_/X _86040_/D sky130_fd_sc_hd__a21oi_4
X_86981_ _82538_/CLK _44737_/Y _86981_/Q sky130_fd_sc_hd__dfxtp_4
X_65009_ _58876_/A _65009_/X sky130_fd_sc_hd__buf_2
X_53023_ _53019_/A _53036_/B _53019_/C _53023_/D _53023_/X sky130_fd_sc_hd__and4_4
X_57900_ _57868_/X _57897_/Y _57898_/Y _57899_/X _57872_/X _57900_/X
+ sky130_fd_sc_hd__o32a_4
X_50235_ _50233_/Y _50227_/X _50234_/Y _50235_/Y sky130_fd_sc_hd__a21boi_4
X_85932_ _86091_/CLK _51866_/Y _85932_/Q sky130_fd_sc_hd__dfxtp_4
X_81055_ _85335_/CLK _75528_/X _81055_/Q sky130_fd_sc_hd__dfxtp_4
X_58880_ _58813_/X _85769_/Q _58838_/X _58880_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_9_12_0_CLK clkbuf_8_6_0_CLK/X clkbuf_9_12_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_80006_ _84658_/Q _64108_/C _80006_/X sky130_fd_sc_hd__xor2_4
X_57831_ _84947_/Q _57819_/X _57823_/X _57830_/X _57831_/Y sky130_fd_sc_hd__a2bb2oi_4
X_69817_ _69386_/X _69388_/X _69816_/X _69817_/Y sky130_fd_sc_hd__a21oi_4
X_50166_ _50092_/A _50166_/X sky130_fd_sc_hd__buf_2
X_85863_ _86500_/CLK _85863_/D _85863_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_609_0_CLK clkbuf_9_304_0_CLK/X _81125_/CLK sky130_fd_sc_hd__clkbuf_1
X_87602_ _88108_/CLK _43027_/Y _73577_/A sky130_fd_sc_hd__dfxtp_4
X_84814_ _82394_/CLK _84814_/D _84814_/Q sky130_fd_sc_hd__dfxtp_4
X_57762_ _57848_/A _58793_/A sky130_fd_sc_hd__buf_2
X_69748_ _87813_/Q _69749_/B sky130_fd_sc_hd__inv_2
X_50097_ _50069_/A _71998_/B _50097_/X sky130_fd_sc_hd__and2_4
X_54974_ _54964_/A _54955_/B _54974_/C _47548_/A _54974_/X sky130_fd_sc_hd__and4_4
X_85794_ _86122_/CLK _85794_/D _65411_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_0_0_CLK clkbuf_8_0_0_CLK/X clkbuf_9_0_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_59501_ _64286_/C _59501_/X sky130_fd_sc_hd__buf_2
X_56713_ _56713_/A _56684_/C _56682_/X _56674_/X _56713_/X sky130_fd_sc_hd__and4_4
Xclkbuf_9_27_0_CLK clkbuf_9_27_0_CLK/A clkbuf_9_27_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_87533_ _87533_/CLK _43219_/X _87533_/Q sky130_fd_sc_hd__dfxtp_4
X_53925_ _53902_/A _50710_/B _53925_/Y sky130_fd_sc_hd__nand2_4
X_84745_ _83438_/CLK _59389_/X _84745_/Q sky130_fd_sc_hd__dfxtp_4
X_57693_ _64717_/A _64601_/A sky130_fd_sc_hd__buf_2
X_81957_ _82339_/CLK _81957_/D _81957_/Q sky130_fd_sc_hd__dfxtp_4
X_69679_ _69674_/X _69677_/X _69678_/X _69679_/X sky130_fd_sc_hd__a21o_4
X_71710_ _70500_/D _71711_/A sky130_fd_sc_hd__buf_2
X_59432_ _59417_/X _83343_/Q _59431_/Y _84735_/D sky130_fd_sc_hd__o21a_4
X_56644_ _56636_/X _56643_/X _85139_/Q _56753_/A _85139_/D sky130_fd_sc_hd__a2bb2o_4
X_80908_ _83918_/CLK _84084_/Q _75656_/A sky130_fd_sc_hd__dfxtp_4
X_87464_ _87720_/CLK _87464_/D _87464_/Q sky130_fd_sc_hd__dfxtp_4
X_53856_ _53848_/A _53856_/B _53856_/Y sky130_fd_sc_hd__nand2_4
X_41870_ _40361_/A _41902_/A _41870_/B1 _41880_/A sky130_fd_sc_hd__a21o_4
X_72690_ _70229_/C _72686_/X _72689_/Y _83189_/D sky130_fd_sc_hd__a21bo_4
X_84676_ _84672_/CLK _84676_/D _80195_/A sky130_fd_sc_hd__dfxtp_4
X_81888_ _82531_/CLK _78079_/X _81888_/Q sky130_fd_sc_hd__dfxtp_4
X_86415_ _86127_/CLK _86415_/D _86415_/Q sky130_fd_sc_hd__dfxtp_4
X_40821_ _40793_/A _40821_/X sky130_fd_sc_hd__buf_2
X_52807_ _52803_/A _52807_/B _52807_/Y sky130_fd_sc_hd__nand2_4
X_71641_ _71641_/A _71644_/C sky130_fd_sc_hd__buf_2
X_83627_ _83627_/CLK _71040_/Y _47657_/A sky130_fd_sc_hd__dfxtp_4
X_59363_ _59354_/Y _59230_/X _59359_/X _59362_/X _59363_/Y sky130_fd_sc_hd__a22oi_4
X_56575_ _56574_/Y _56575_/X sky130_fd_sc_hd__buf_2
X_80839_ _80746_/CLK _80871_/Q _74875_/B sky130_fd_sc_hd__dfxtp_4
X_87395_ _87150_/CLK _87395_/D _87395_/Q sky130_fd_sc_hd__dfxtp_4
X_53787_ _85568_/Q _53784_/X _53786_/Y _53787_/Y sky130_fd_sc_hd__o21ai_4
X_50999_ _86092_/Q _50992_/X _50998_/Y _50999_/Y sky130_fd_sc_hd__o21ai_4
X_58314_ _58314_/A _58326_/B _58314_/Y sky130_fd_sc_hd__nand2_4
X_43540_ _43518_/X _43523_/X _40432_/X _87368_/Q _43528_/X _43540_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55526_ _55521_/X _55525_/X _44113_/X _55526_/X sky130_fd_sc_hd__a21o_4
X_74360_ _83083_/Q _72699_/X _74359_/Y _83083_/D sky130_fd_sc_hd__a21bo_4
X_86346_ _82381_/CLK _49665_/Y _86346_/Q sky130_fd_sc_hd__dfxtp_4
X_40752_ _40731_/X _40923_/A _40751_/X _40753_/A sky130_fd_sc_hd__o21ai_4
X_52738_ _52657_/A _52744_/A sky130_fd_sc_hd__buf_2
X_59294_ _59231_/X _85417_/Q _59293_/X _59294_/Y sky130_fd_sc_hd__o21ai_4
X_71572_ _71570_/X _71583_/B _71574_/C _71572_/Y sky130_fd_sc_hd__nor3_4
X_83558_ _86558_/CLK _83558_/D _83558_/Q sky130_fd_sc_hd__dfxtp_4
X_73311_ _73214_/X _83060_/Q _73238_/X _73310_/X _73311_/X sky130_fd_sc_hd__a211o_4
X_70523_ _57674_/Y _70500_/Y _70522_/Y _83756_/D sky130_fd_sc_hd__o21ai_4
X_58245_ _58219_/X _58240_/Y _58244_/Y _84899_/D sky130_fd_sc_hd__a21oi_4
XPHY_710 sky130_fd_sc_hd__decap_3
X_82509_ _82702_/CLK _82509_/D _78469_/A sky130_fd_sc_hd__dfxtp_4
X_55457_ _55301_/X _55457_/X sky130_fd_sc_hd__buf_2
X_43471_ _41663_/X _43465_/X _87405_/Q _43467_/X _87405_/D sky130_fd_sc_hd__a2bb2o_4
X_74291_ _74297_/A _74297_/B _55975_/X _74291_/Y sky130_fd_sc_hd__nand3_4
X_86277_ _85957_/CLK _86277_/D _86277_/Q sky130_fd_sc_hd__dfxtp_4
X_40683_ _40832_/A _40683_/X sky130_fd_sc_hd__buf_2
X_52669_ _52648_/X _52661_/B _52654_/C _46783_/X _52669_/X sky130_fd_sc_hd__and4_4
X_83489_ _83756_/CLK _83489_/D _83489_/Q sky130_fd_sc_hd__dfxtp_4
X_45210_ _56518_/C _45209_/X _45189_/X _45210_/X sky130_fd_sc_hd__o21a_4
X_76030_ _81712_/D _76036_/C _76029_/Y _76030_/Y sky130_fd_sc_hd__a21oi_4
X_88016_ _87260_/CLK _88016_/D _88016_/Q sky130_fd_sc_hd__dfxtp_4
X_42422_ _40485_/X _42414_/X _87872_/Q _42415_/X _87872_/D sky130_fd_sc_hd__a2bb2o_4
X_54408_ _54399_/X _54395_/B _54402_/C _46856_/A _54408_/X sky130_fd_sc_hd__and4_4
X_73242_ _48559_/Y _73241_/Y _73242_/X sky130_fd_sc_hd__xor2_4
X_85228_ _85192_/CLK _56344_/Y _85228_/Q sky130_fd_sc_hd__dfxtp_4
X_46190_ _46186_/X _74842_/B _46189_/Y _86763_/D sky130_fd_sc_hd__and3_4
X_70454_ _70758_/A _70827_/B _71287_/C _70609_/A _70454_/Y sky130_fd_sc_hd__nand4_4
X_58176_ _58171_/X _83491_/Q _58175_/Y _84915_/D sky130_fd_sc_hd__o21a_4
X_55388_ _55387_/X _55388_/Y sky130_fd_sc_hd__inv_2
X_45141_ _45141_/A _45182_/B _45141_/Y sky130_fd_sc_hd__nand2_4
X_57127_ _57158_/C _57153_/B sky130_fd_sc_hd__buf_2
X_42353_ _41715_/X _42342_/X _87907_/Q _42343_/X _87907_/D sky130_fd_sc_hd__a2bb2o_4
X_54339_ _54325_/A _54353_/B _54317_/X _46743_/Y _54339_/X sky130_fd_sc_hd__and4_4
X_73173_ _87055_/Q _73104_/B _73173_/Y sky130_fd_sc_hd__nor2_4
X_85159_ _83016_/CLK _56534_/Y _85159_/Q sky130_fd_sc_hd__dfxtp_4
X_70385_ _50862_/B _70364_/X _70384_/Y _70385_/Y sky130_fd_sc_hd__o21ai_4
X_41304_ _41304_/A _41292_/B _41304_/X sky130_fd_sc_hd__or2_4
X_72124_ _72123_/X _85697_/Q _59334_/X _72124_/X sky130_fd_sc_hd__o21a_4
X_45072_ _45064_/X _45068_/Y _45071_/Y _45072_/Y sky130_fd_sc_hd__a21oi_4
X_57058_ _56671_/X _57058_/B _57058_/Y sky130_fd_sc_hd__nand2_4
X_42284_ _42279_/X _42275_/X _41536_/X _87940_/Q _42276_/X _42284_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77981_ _77983_/A _77983_/C _77981_/Y sky130_fd_sc_hd__nand2_4
X_48900_ _48899_/Y _48901_/B sky130_fd_sc_hd__buf_2
X_44023_ _44022_/X _58834_/A sky130_fd_sc_hd__buf_2
X_56009_ _55928_/B _74310_/C sky130_fd_sc_hd__buf_2
X_79720_ _65047_/C _72313_/Y _79719_/Y _79720_/X sky130_fd_sc_hd__o21a_4
X_41235_ _40568_/A _41235_/X sky130_fd_sc_hd__buf_2
X_72055_ _72025_/A _53879_/B _72055_/Y sky130_fd_sc_hd__nand2_4
X_76932_ _76932_/A _76932_/Y sky130_fd_sc_hd__inv_2
X_49880_ _49906_/A _49880_/X sky130_fd_sc_hd__buf_2
X_71006_ _71055_/A _71064_/B _71001_/C _71006_/Y sky130_fd_sc_hd__nand3_4
X_48831_ _48831_/A _52216_/B _48831_/Y sky130_fd_sc_hd__nand2_4
X_79651_ _79647_/X _79664_/A _79651_/X sky130_fd_sc_hd__xor2_4
X_41166_ _41165_/X _41152_/X _68631_/B _41153_/X _88265_/D sky130_fd_sc_hd__a2bb2o_4
X_76863_ _81593_/Q _81465_/D _81561_/D sky130_fd_sc_hd__xor2_4
X_78602_ _78602_/A _78602_/Y sky130_fd_sc_hd__inv_2
X_75814_ _80796_/D _75807_/A _75815_/A sky130_fd_sc_hd__and2_4
X_48762_ _48758_/Y _48760_/X _48761_/X _86488_/D sky130_fd_sc_hd__a21oi_4
X_79582_ _79588_/A _79587_/A sky130_fd_sc_hd__inv_2
X_45974_ _45962_/X _45974_/X sky130_fd_sc_hd__buf_2
X_41097_ _41061_/X _40919_/B _41096_/X _41098_/A sky130_fd_sc_hd__o21ai_4
X_76794_ _76774_/X _76786_/X _76794_/X sky130_fd_sc_hd__and2_4
X_47713_ _47003_/A _47714_/A sky130_fd_sc_hd__buf_2
X_78533_ _78522_/Y _78526_/B _78525_/A _78533_/X sky130_fd_sc_hd__o21a_4
X_44925_ _80671_/Q _45237_/A sky130_fd_sc_hd__buf_2
X_75745_ _75735_/Y _75740_/B _75745_/X sky130_fd_sc_hd__or2_4
X_48693_ _48693_/A _48694_/A sky130_fd_sc_hd__inv_2
X_60971_ _60961_/X _60963_/X _60940_/Y _60968_/X _60970_/X _84547_/D
+ sky130_fd_sc_hd__o41a_4
X_72957_ _73132_/A _72957_/B _72957_/X sky130_fd_sc_hd__and2_4
X_62710_ _62979_/A _62711_/A sky130_fd_sc_hd__buf_2
X_47644_ _55026_/D _53165_/D sky130_fd_sc_hd__buf_2
X_71908_ _74529_/A _70710_/C _71902_/X _71928_/D _71908_/Y sky130_fd_sc_hd__nand4_4
X_78464_ _78464_/A _78464_/X sky130_fd_sc_hd__buf_2
X_44856_ _41767_/Y _44848_/X _67964_/B _44849_/X _86917_/D sky130_fd_sc_hd__a2bb2o_4
X_75676_ _80910_/Q _75678_/A sky130_fd_sc_hd__inv_2
X_63690_ _60422_/A _63849_/A sky130_fd_sc_hd__buf_2
X_72888_ _44189_/X _72888_/X sky130_fd_sc_hd__buf_2
X_77415_ _77415_/A _77415_/X sky130_fd_sc_hd__buf_2
X_43807_ _43790_/X _43797_/X _41082_/X _69494_/B _43791_/X _43808_/A
+ sky130_fd_sc_hd__o32ai_4
X_62641_ _62886_/A _62642_/B sky130_fd_sc_hd__buf_2
X_74627_ _44196_/A _45933_/Y _44037_/X _74627_/Y sky130_fd_sc_hd__a21oi_4
X_47575_ _72188_/A _47570_/X _47574_/Y _47575_/Y sky130_fd_sc_hd__o21ai_4
X_71839_ _71829_/X _71839_/B _70786_/A _70721_/A _71839_/X sky130_fd_sc_hd__and4_4
X_78395_ _78426_/C _78426_/B _78395_/X sky130_fd_sc_hd__and2_4
X_44787_ _46298_/A _44803_/A sky130_fd_sc_hd__buf_2
X_41999_ _88076_/Q _41999_/Y sky130_fd_sc_hd__inv_2
X_49314_ _49302_/A _51350_/B _49314_/Y sky130_fd_sc_hd__nand2_4
X_46526_ _46526_/A _47972_/A sky130_fd_sc_hd__buf_2
X_65360_ _65258_/A _65360_/B _65360_/X sky130_fd_sc_hd__and2_4
X_77346_ _77318_/A _77318_/B _77317_/X _77334_/Y _77346_/Y sky130_fd_sc_hd__nand4_4
X_43738_ _40903_/X _43736_/X _87289_/Q _43737_/X _43738_/X sky130_fd_sc_hd__a2bb2o_4
X_62572_ _62572_/A _62572_/X sky130_fd_sc_hd__buf_2
X_74558_ _44990_/A _74551_/X _74557_/X _74558_/Y sky130_fd_sc_hd__o21ai_4
X_64311_ _64304_/X _64305_/X _64307_/X _64310_/Y _64267_/X _64311_/X
+ sky130_fd_sc_hd__o41a_4
X_61523_ _61400_/X _61541_/C sky130_fd_sc_hd__buf_2
X_49245_ _49241_/A _49245_/B _49245_/Y sky130_fd_sc_hd__nand2_4
X_73509_ _73509_/A _73530_/B _73509_/Y sky130_fd_sc_hd__nor2_4
X_46457_ _46434_/A _51324_/B _46457_/Y sky130_fd_sc_hd__nand2_4
X_65291_ _65288_/X _65631_/B _65290_/X _65291_/Y sky130_fd_sc_hd__nand3_4
X_77277_ _77277_/A _77277_/B _81893_/D sky130_fd_sc_hd__xnor2_4
X_43669_ _43668_/X _87319_/D sky130_fd_sc_hd__inv_2
X_74489_ _74486_/Y _74463_/X _74488_/X _83056_/D sky130_fd_sc_hd__a21oi_4
X_67030_ _67027_/X _67030_/B _67030_/Y sky130_fd_sc_hd__nand2_4
X_79016_ _79010_/A _79010_/B _79016_/Y sky130_fd_sc_hd__nor2_4
X_45408_ _45408_/A _55625_/B sky130_fd_sc_hd__inv_2
X_64242_ _61368_/A _64219_/B _64242_/Y sky130_fd_sc_hd__nor2_4
X_76228_ _81256_/Q _81512_/D _76233_/C sky130_fd_sc_hd__nand2_4
X_49176_ _49176_/A _50712_/B sky130_fd_sc_hd__buf_2
X_61454_ _61447_/Y _61449_/Y _61403_/X _61451_/Y _61453_/Y _61454_/X
+ sky130_fd_sc_hd__a41o_4
X_46388_ _86741_/Q _46364_/X _46387_/Y _46388_/Y sky130_fd_sc_hd__o21ai_4
X_48127_ _48075_/X _46567_/A _48126_/X _48337_/A sky130_fd_sc_hd__o21ai_4
X_60405_ _60404_/Y _60410_/B sky130_fd_sc_hd__inv_2
X_45339_ _45265_/A _45339_/X sky130_fd_sc_hd__buf_2
X_64173_ _64184_/A _58364_/A _64173_/C _64173_/X sky130_fd_sc_hd__and3_4
X_76159_ _76159_/A _76158_/B _76159_/Y sky130_fd_sc_hd__nand2_4
X_61385_ _61383_/X _61349_/X _61384_/Y _61385_/Y sky130_fd_sc_hd__a21oi_4
X_63124_ _63100_/A _63124_/B _63079_/C _63124_/D _63124_/X sky130_fd_sc_hd__and4_4
X_48058_ _47981_/X _48058_/B _48058_/X sky130_fd_sc_hd__and2_4
X_60336_ _60335_/Y _60337_/D sky130_fd_sc_hd__buf_2
X_68981_ _87482_/Q _68792_/X _68979_/X _68980_/X _68981_/X sky130_fd_sc_hd__a211o_4
X_47009_ _86680_/Q _47004_/X _47008_/Y _47009_/Y sky130_fd_sc_hd__o21ai_4
X_67932_ _67909_/A _67932_/B _67932_/X sky130_fd_sc_hd__and2_4
X_63055_ _63055_/A _63231_/A sky130_fd_sc_hd__buf_2
X_79918_ _58108_/Y _65872_/C _79918_/Y sky130_fd_sc_hd__nand2_4
X_60267_ _60267_/A _60267_/X sky130_fd_sc_hd__buf_2
X_50020_ _49915_/A _50040_/B sky130_fd_sc_hd__buf_2
X_62006_ _63586_/A _59841_/X _61551_/A _61981_/X _62006_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_10_580_0_CLK clkbuf_9_290_0_CLK/X _83944_/CLK sky130_fd_sc_hd__clkbuf_1
X_67863_ _67863_/A _67863_/X sky130_fd_sc_hd__buf_2
X_79849_ _79875_/A _79859_/A sky130_fd_sc_hd__inv_2
X_60198_ _60198_/A _60198_/Y sky130_fd_sc_hd__inv_2
X_69602_ _81983_/D _69564_/X _69601_/X _83911_/D sky130_fd_sc_hd__a21bo_4
X_66814_ _88393_/Q _66715_/X _66717_/X _66813_/X _66814_/X sky130_fd_sc_hd__a211o_4
X_82860_ _82860_/CLK _82860_/D _82860_/Q sky130_fd_sc_hd__dfxtp_4
X_67794_ _87968_/Q _67770_/X _67748_/X _67793_/X _67794_/X sky130_fd_sc_hd__a211o_4
X_81811_ _81811_/CLK _81619_/Q _47355_/A sky130_fd_sc_hd__dfxtp_4
X_69533_ _69626_/A _87254_/Q _69533_/X sky130_fd_sc_hd__and2_4
X_66745_ _66795_/A _66745_/B _66745_/X sky130_fd_sc_hd__and2_4
X_51971_ _66006_/B _51945_/X _51970_/Y _51971_/Y sky130_fd_sc_hd__o21ai_4
X_63957_ _61490_/X _63908_/B _63894_/C _63908_/D _63957_/Y sky130_fd_sc_hd__nand4_4
X_82791_ _82792_/CLK _82823_/Q _78375_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_595_0_CLK clkbuf_9_297_0_CLK/X _81933_/CLK sky130_fd_sc_hd__clkbuf_1
X_53710_ _85583_/Q _53687_/X _53709_/Y _53710_/Y sky130_fd_sc_hd__o21ai_4
X_84530_ _84292_/CLK _61043_/X _84530_/Q sky130_fd_sc_hd__dfxtp_4
X_50922_ _86106_/Q _50910_/X _50921_/Y _50922_/Y sky130_fd_sc_hd__o21ai_4
X_62908_ _60274_/X _62908_/X sky130_fd_sc_hd__buf_2
X_81742_ _88175_/CLK _81742_/D _81742_/Q sky130_fd_sc_hd__dfxtp_4
X_69464_ _83922_/Q _69439_/X _69463_/X _69464_/X sky130_fd_sc_hd__a21bo_4
X_54690_ _54688_/Y _54666_/X _54689_/X _54690_/Y sky130_fd_sc_hd__a21oi_4
X_66676_ _66651_/A _66676_/B _66676_/X sky130_fd_sc_hd__and2_4
X_63888_ _57656_/X _63902_/B _63902_/C _63902_/D _63888_/Y sky130_fd_sc_hd__nand4_4
X_68415_ _87857_/Q _68415_/Y sky130_fd_sc_hd__inv_2
X_53641_ _53778_/A _52119_/B _53641_/Y sky130_fd_sc_hd__nand2_4
X_65627_ _65362_/X _85588_/Q _65363_/X _65626_/X _65627_/X sky130_fd_sc_hd__a211o_4
X_84461_ _82452_/CLK _61672_/Y _79129_/B sky130_fd_sc_hd__dfxtp_4
X_50853_ _86120_/Q _50804_/X _50852_/Y _50853_/Y sky130_fd_sc_hd__o21ai_4
X_62839_ _62792_/X _62839_/B _84378_/Q _62839_/Y sky130_fd_sc_hd__nor3_4
X_81673_ _81671_/CLK _80002_/X _81673_/Q sky130_fd_sc_hd__dfxtp_4
X_69395_ _88032_/Q _69315_/X _69393_/X _69394_/X _69395_/X sky130_fd_sc_hd__a211o_4
X_86200_ _85879_/CLK _86200_/D _86200_/Q sky130_fd_sc_hd__dfxtp_4
X_83412_ _83380_/CLK _71684_/X _83412_/Q sky130_fd_sc_hd__dfxtp_4
X_56360_ _56360_/A _56358_/B _55730_/B _56360_/Y sky130_fd_sc_hd__nand3_4
X_80624_ _80624_/A _80623_/X _80632_/A sky130_fd_sc_hd__nand2_4
X_68346_ _69645_/A _68472_/A sky130_fd_sc_hd__buf_2
X_87180_ _87183_/CLK _44220_/Y _87180_/Q sky130_fd_sc_hd__dfxtp_4
X_53572_ _53548_/A _57605_/B _53572_/Y sky130_fd_sc_hd__nand2_4
X_65558_ _65929_/A _65559_/B sky130_fd_sc_hd__buf_2
X_84392_ _84392_/CLK _62674_/Y _84392_/Q sky130_fd_sc_hd__dfxtp_4
X_50784_ _50782_/Y _50768_/X _50783_/Y _86134_/D sky130_fd_sc_hd__a21boi_4
X_55311_ _55305_/X _55311_/X sky130_fd_sc_hd__buf_2
X_86131_ _86424_/CLK _50798_/Y _86131_/Q sky130_fd_sc_hd__dfxtp_4
X_52523_ _65115_/B _52516_/X _52522_/Y _52523_/Y sky130_fd_sc_hd__o21ai_4
X_64509_ _64689_/A _64741_/B _79605_/B _64509_/Y sky130_fd_sc_hd__nor3_4
X_83343_ _83338_/CLK _71880_/X _83343_/Q sky130_fd_sc_hd__dfxtp_4
X_80555_ _80562_/B _80554_/Y _82266_/D sky130_fd_sc_hd__xor2_4
X_56291_ _56368_/A _56270_/B _55976_/B _56291_/Y sky130_fd_sc_hd__nand3_4
X_68277_ _68254_/X _67698_/Y _68268_/X _68276_/Y _68277_/X sky130_fd_sc_hd__a211o_4
X_65489_ _65592_/A _65489_/B _65489_/X sky130_fd_sc_hd__and2_4
X_58030_ _58605_/A _58030_/X sky130_fd_sc_hd__buf_2
X_55242_ _72712_/C _83317_/Q _55209_/X _56889_/B sky130_fd_sc_hd__nand3_4
X_67228_ _87416_/Q _67156_/X _67226_/X _67227_/X _67228_/X sky130_fd_sc_hd__a211o_4
X_86062_ _85745_/CLK _51166_/Y _86062_/Q sky130_fd_sc_hd__dfxtp_4
X_52454_ _52436_/A _52454_/B _52454_/Y sky130_fd_sc_hd__nand2_4
X_83274_ _86297_/CLK _72213_/Y _83274_/Q sky130_fd_sc_hd__dfxtp_4
X_80486_ _80482_/Y _80485_/Y _80487_/A sky130_fd_sc_hd__xor2_4
X_85013_ _85013_/CLK _85013_/D _45584_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_533_0_CLK clkbuf_9_266_0_CLK/X _83918_/CLK sky130_fd_sc_hd__clkbuf_1
X_51405_ _86016_/Q _51402_/X _51404_/Y _51405_/Y sky130_fd_sc_hd__o21ai_4
X_82225_ _82786_/CLK _82257_/Q _77443_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_6_24_0_CLK clkbuf_6_25_0_CLK/A clkbuf_6_24_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_55173_ _55125_/A _55244_/A sky130_fd_sc_hd__buf_2
X_67159_ _67155_/X _67158_/X _67085_/X _67159_/X sky130_fd_sc_hd__a21o_4
X_52385_ _52385_/A _52385_/B _52385_/X sky130_fd_sc_hd__and2_4
X_54124_ _54122_/Y _54117_/X _54123_/X _85500_/D sky130_fd_sc_hd__a21oi_4
X_51336_ _65120_/B _51332_/X _51335_/Y _51336_/Y sky130_fd_sc_hd__o21ai_4
X_70170_ _70127_/X _70231_/A sky130_fd_sc_hd__buf_2
X_82156_ _84220_/CLK _84148_/Q _82156_/Q sky130_fd_sc_hd__dfxtp_4
X_59981_ _59980_/X _59570_/A _59905_/B _59981_/Y sky130_fd_sc_hd__nor3_4
X_81107_ _81087_/CLK _79738_/Y _81107_/Q sky130_fd_sc_hd__dfxtp_4
X_58932_ _84789_/Q _58871_/X _58924_/X _58931_/X _84789_/D sky130_fd_sc_hd__a2bb2oi_4
X_54055_ _85514_/Q _54018_/X _54054_/Y _54055_/Y sky130_fd_sc_hd__o21ai_4
X_51267_ _51262_/Y _51263_/X _51266_/X _51267_/Y sky130_fd_sc_hd__a21oi_4
X_86964_ _88224_/CLK _86964_/D _86964_/Q sky130_fd_sc_hd__dfxtp_4
X_82087_ _82133_/CLK _77294_/B _82087_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_548_0_CLK clkbuf_9_274_0_CLK/X _81756_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_6_39_0_CLK clkbuf_6_39_0_CLK/A clkbuf_7_78_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_53006_ _85714_/Q _52984_/X _53005_/Y _53006_/Y sky130_fd_sc_hd__o21ai_4
X_41020_ _40991_/X _81714_/Q _41019_/X _41021_/A sky130_fd_sc_hd__o21a_4
X_50218_ _50218_/A _50655_/A sky130_fd_sc_hd__buf_2
X_85915_ _85915_/CLK _85915_/D _73707_/B sky130_fd_sc_hd__dfxtp_4
X_81038_ _81038_/CLK _75249_/Y _81038_/Q sky130_fd_sc_hd__dfxtp_4
X_58863_ _58860_/Y _58862_/Y _58761_/X _58863_/X sky130_fd_sc_hd__a21o_4
X_51198_ _51195_/Y _51175_/X _51197_/X _86056_/D sky130_fd_sc_hd__a21oi_4
X_86895_ _86896_/CLK _45160_/Y _64401_/B sky130_fd_sc_hd__dfxtp_4
X_57814_ _58020_/A _57814_/X sky130_fd_sc_hd__buf_2
X_50149_ _50153_/A _49073_/X _50149_/Y sky130_fd_sc_hd__nand2_4
X_73860_ _72874_/A _73954_/A sky130_fd_sc_hd__buf_2
X_85846_ _83303_/CLK _52321_/Y _64904_/B sky130_fd_sc_hd__dfxtp_4
X_58794_ _58756_/X _85935_/Q _58793_/X _58794_/X sky130_fd_sc_hd__o21a_4
X_72811_ _44131_/A _73067_/A sky130_fd_sc_hd__buf_2
X_57745_ _86654_/Q _57833_/B _57745_/Y sky130_fd_sc_hd__nor2_4
X_54957_ _54961_/A _47526_/Y _54957_/Y sky130_fd_sc_hd__nand2_4
X_42971_ _41992_/A _42971_/X sky130_fd_sc_hd__buf_2
X_73791_ _73792_/B _73779_/Y _73790_/X _73791_/X sky130_fd_sc_hd__a21o_4
X_85777_ _85778_/CLK _52666_/Y _85777_/Q sky130_fd_sc_hd__dfxtp_4
X_82989_ _83012_/CLK _74674_/X _82989_/Q sky130_fd_sc_hd__dfxtp_4
X_44710_ _44533_/A _44710_/X sky130_fd_sc_hd__buf_2
X_75530_ _75530_/A _75525_/X _75530_/Y sky130_fd_sc_hd__nand2_4
X_87516_ _87767_/CLK _87516_/D _87516_/Q sky130_fd_sc_hd__dfxtp_4
X_41922_ _41922_/A _41922_/Y sky130_fd_sc_hd__inv_2
X_53908_ _53898_/A _49135_/A _53908_/Y sky130_fd_sc_hd__nand2_4
X_84728_ _83402_/CLK _59455_/X _84728_/Q sky130_fd_sc_hd__dfxtp_4
X_72742_ _88339_/Q _56939_/X _72741_/X _72742_/Y sky130_fd_sc_hd__o21ai_4
X_45690_ _45688_/Y _45627_/X _45644_/X _45689_/Y _45690_/X sky130_fd_sc_hd__a211o_4
X_57676_ _45909_/X _57672_/X _57675_/Y _57676_/X sky130_fd_sc_hd__o21a_4
X_54888_ _54888_/A _54910_/A sky130_fd_sc_hd__buf_2
X_59415_ _59415_/A _59399_/B _59415_/Y sky130_fd_sc_hd__nand2_4
X_44641_ _44638_/X _44639_/X _41035_/X _87021_/Q _44640_/X _44642_/A
+ sky130_fd_sc_hd__o32ai_4
X_56627_ _56602_/X _56627_/B _56696_/B _56627_/Y sky130_fd_sc_hd__nor3_4
X_75461_ _75461_/A _75509_/A sky130_fd_sc_hd__inv_2
X_41853_ _40524_/X _41847_/X _67206_/B _41848_/X _88121_/D sky130_fd_sc_hd__a2bb2o_4
X_87447_ _87382_/CLK _43389_/X _87447_/Q sky130_fd_sc_hd__dfxtp_4
X_53839_ _53825_/A _72014_/B _53839_/Y sky130_fd_sc_hd__nand2_4
X_72673_ _72687_/A _72683_/A sky130_fd_sc_hd__buf_2
X_84659_ _84660_/CLK _84659_/D _84659_/Q sky130_fd_sc_hd__dfxtp_4
X_77200_ _77200_/A _82302_/D _77200_/X sky130_fd_sc_hd__xor2_4
X_74412_ _72001_/A _74412_/X sky130_fd_sc_hd__buf_2
X_40804_ _82873_/Q _40779_/B _40804_/X sky130_fd_sc_hd__or2_4
X_59346_ _59345_/X _59346_/X sky130_fd_sc_hd__buf_2
X_47360_ _47360_/A _53005_/B sky130_fd_sc_hd__buf_2
X_71624_ _71528_/X _71446_/X _71628_/A sky130_fd_sc_hd__nor2_4
X_78180_ _78176_/Y _78179_/X _78192_/A sky130_fd_sc_hd__nand2_4
X_44572_ _44571_/Y _44572_/Y sky130_fd_sc_hd__inv_2
X_56558_ _56557_/X _56558_/X sky130_fd_sc_hd__buf_2
X_75392_ _75392_/A _75396_/A sky130_fd_sc_hd__inv_2
X_87378_ _87995_/CLK _87378_/D _87378_/Q sky130_fd_sc_hd__dfxtp_4
X_41784_ _40414_/X _41784_/B _41784_/X sky130_fd_sc_hd__or2_4
X_46311_ _51256_/A _46428_/B _46428_/C _46311_/X sky130_fd_sc_hd__and3_4
X_77131_ _77141_/A _77142_/A _77132_/B sky130_fd_sc_hd__xor2_4
X_43523_ _43425_/X _43523_/X sky130_fd_sc_hd__buf_2
X_55509_ _45572_/A _55505_/X _55506_/X _55508_/Y _55509_/X sky130_fd_sc_hd__a211o_4
X_86329_ _86647_/CLK _86329_/D _86329_/Q sky130_fd_sc_hd__dfxtp_4
X_74343_ _74351_/A _74342_/X _55801_/C _74343_/Y sky130_fd_sc_hd__nand3_4
X_40735_ _40734_/X _40719_/X _69004_/B _40720_/X _40735_/X sky130_fd_sc_hd__a2bb2o_4
X_47291_ _86650_/Q _47286_/X _47290_/Y _47291_/Y sky130_fd_sc_hd__o21ai_4
X_59277_ _59177_/X _86059_/Q _59276_/X _59277_/Y sky130_fd_sc_hd__o21ai_4
X_71555_ _71602_/C _71164_/B _71556_/A sky130_fd_sc_hd__nor2_4
X_56489_ _56462_/X _56049_/Y _56488_/Y _85177_/D sky130_fd_sc_hd__o21ai_4
X_49030_ _49018_/X _48520_/A _49029_/Y _49031_/A sky130_fd_sc_hd__a21o_4
X_46242_ _46242_/A _46242_/Y sky130_fd_sc_hd__inv_2
XPHY_540 sky130_fd_sc_hd__decap_3
X_70506_ _70506_/A _71170_/A sky130_fd_sc_hd__buf_2
X_58228_ _63400_/B _58228_/X sky130_fd_sc_hd__buf_2
X_77062_ _77050_/A _81906_/Q _77062_/Y sky130_fd_sc_hd__nand2_4
X_43454_ _43454_/A _43454_/Y sky130_fd_sc_hd__inv_2
X_74274_ _74016_/X _85602_/Q _56933_/X _74273_/X _74274_/X sky130_fd_sc_hd__a211o_4
XPHY_551 sky130_fd_sc_hd__decap_3
X_40666_ _40601_/X _81139_/Q _40665_/X _40667_/A sky130_fd_sc_hd__o21a_4
X_71486_ _71486_/A _71487_/A sky130_fd_sc_hd__inv_2
XPHY_562 sky130_fd_sc_hd__decap_3
XPHY_573 sky130_fd_sc_hd__decap_3
X_76013_ _81710_/D _76013_/B _76013_/Y sky130_fd_sc_hd__nand2_4
X_42405_ _42405_/A _42405_/Y sky130_fd_sc_hd__inv_2
XPHY_584 sky130_fd_sc_hd__decap_3
X_73225_ _73225_/A _73196_/B _73225_/Y sky130_fd_sc_hd__nor2_4
X_70437_ _70994_/A _70947_/B sky130_fd_sc_hd__buf_2
X_46173_ _45904_/X _46173_/X sky130_fd_sc_hd__buf_2
X_58159_ _63044_/A _61368_/A sky130_fd_sc_hd__buf_2
XPHY_595 sky130_fd_sc_hd__decap_3
X_43385_ _41433_/X _43371_/X _87448_/Q _43372_/X _43385_/X sky130_fd_sc_hd__a2bb2o_4
X_40597_ _40565_/Y _40755_/A sky130_fd_sc_hd__buf_2
X_45124_ _45124_/A _45182_/B _45124_/Y sky130_fd_sc_hd__nand2_4
X_42336_ _42330_/X _42319_/X _41676_/X _87915_/Q _42320_/X _42337_/A
+ sky130_fd_sc_hd__o32ai_4
X_61170_ _61117_/X _61169_/X _59512_/X _61170_/Y sky130_fd_sc_hd__a21oi_4
X_73156_ _73156_/A _73155_/X _73156_/Y sky130_fd_sc_hd__nand2_4
X_70368_ _70984_/A _70368_/X sky130_fd_sc_hd__buf_2
X_60121_ _57689_/A _60267_/A sky130_fd_sc_hd__buf_2
X_72107_ _72083_/A _72107_/X sky130_fd_sc_hd__buf_2
X_49932_ _49925_/X _49915_/X _49953_/C _53144_/D _49932_/X sky130_fd_sc_hd__and4_4
X_45055_ _45043_/X _45050_/Y _45054_/Y _45055_/Y sky130_fd_sc_hd__a21oi_4
X_42267_ _42266_/Y _87949_/D sky130_fd_sc_hd__inv_2
X_77964_ _77964_/A _81948_/D _77965_/A sky130_fd_sc_hd__xor2_4
X_73087_ _73704_/A _73087_/X sky130_fd_sc_hd__buf_2
X_70299_ _70296_/X _70297_/X _83102_/Q _70301_/D _70299_/X sky130_fd_sc_hd__and4_4
X_44006_ _44005_/X _44006_/X sky130_fd_sc_hd__buf_2
X_79703_ _79702_/X _79703_/Y sky130_fd_sc_hd__inv_2
X_41218_ _41513_/A _40700_/A _41218_/X sky130_fd_sc_hd__or2_4
X_72038_ _72025_/A _53863_/A _72038_/Y sky130_fd_sc_hd__nand2_4
X_76915_ _76915_/A _81470_/D _81566_/D sky130_fd_sc_hd__xor2_4
X_60052_ _59971_/X _60049_/Y _60015_/Y _62203_/A _60051_/Y _84670_/D
+ sky130_fd_sc_hd__a41oi_4
X_49863_ _49860_/Y _49844_/X _49862_/X _49863_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_8_7_0_CLK clkbuf_8_7_0_CLK/A clkbuf_8_7_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_42198_ _41312_/X _42192_/X _87982_/Q _42193_/X _42198_/X sky130_fd_sc_hd__a2bb2o_4
X_77895_ _77884_/A _77883_/Y _77894_/X _77895_/Y sky130_fd_sc_hd__a21oi_4
X_48814_ _52199_/A _48829_/B _48814_/C _48814_/X sky130_fd_sc_hd__and3_4
X_79634_ _84209_/Q _83257_/Q _79634_/Y sky130_fd_sc_hd__nand2_4
X_41149_ _41149_/A _41145_/B _41149_/X sky130_fd_sc_hd__or2_4
X_64860_ _64804_/A _64860_/B _64860_/X sky130_fd_sc_hd__and2_4
X_76846_ _81496_/Q _76846_/Y sky130_fd_sc_hd__inv_2
X_49794_ _52679_/A _49794_/X sky130_fd_sc_hd__buf_2
X_63811_ _60984_/A _63860_/D sky130_fd_sc_hd__buf_2
X_48745_ _48742_/Y _48734_/X _48744_/X _86491_/D sky130_fd_sc_hd__a21oi_4
X_79565_ _79564_/Y _79565_/Y sky130_fd_sc_hd__inv_2
X_45957_ _45957_/A _74831_/A sky130_fd_sc_hd__buf_2
X_64791_ _64787_/Y _64662_/X _64790_/X _84227_/D sky130_fd_sc_hd__a21o_4
X_76777_ _76766_/Y _81359_/D sky130_fd_sc_hd__inv_2
X_73989_ _73989_/A _73250_/A _73989_/Y sky130_fd_sc_hd__nor2_4
X_66530_ _66563_/A _69245_/A sky130_fd_sc_hd__buf_2
X_78516_ _78491_/X _78492_/Y _78486_/Y _78516_/Y sky130_fd_sc_hd__a21boi_4
X_44908_ _61298_/B _44905_/X _44907_/X _44908_/Y sky130_fd_sc_hd__o21ai_4
X_63742_ _61323_/A _63741_/X _63742_/Y sky130_fd_sc_hd__nor2_4
X_75728_ _75715_/A _75714_/Y _75728_/Y sky130_fd_sc_hd__nor2_4
X_48676_ _48676_/A _48632_/B _48676_/Y sky130_fd_sc_hd__nand2_4
X_60954_ _60901_/A _60954_/X sky130_fd_sc_hd__buf_2
X_79496_ _79474_/Y _79496_/B _79496_/X sky130_fd_sc_hd__or2_4
X_45888_ _45888_/A _58517_/A sky130_fd_sc_hd__buf_2
X_47627_ _81239_/Q _55013_/D sky130_fd_sc_hd__inv_2
X_66461_ _66457_/Y _64532_/X _66460_/X _84119_/D sky130_fd_sc_hd__o21ai_4
X_78447_ _82796_/Q _78447_/B _78466_/B sky130_fd_sc_hd__xnor2_4
X_44839_ _45964_/A _44839_/X sky130_fd_sc_hd__buf_2
X_63673_ _59433_/Y _63626_/X _61655_/A _63627_/X _63673_/X sky130_fd_sc_hd__a2bb2o_4
X_75659_ _75659_/A _75659_/B _75660_/B sky130_fd_sc_hd__and2_4
X_60885_ _60879_/D _60996_/B sky130_fd_sc_hd__buf_2
X_68200_ _68160_/A _68200_/X sky130_fd_sc_hd__buf_2
X_65412_ _65334_/X _86114_/Q _65256_/X _65411_/X _65412_/X sky130_fd_sc_hd__a211o_4
X_62624_ _61682_/B _62548_/C _59987_/X _62548_/B _62623_/X _62624_/X
+ sky130_fd_sc_hd__a41o_4
X_69180_ _87536_/Q _69044_/X _68979_/X _69179_/X _69180_/X sky130_fd_sc_hd__a211o_4
X_47558_ _47558_/A _53118_/D sky130_fd_sc_hd__buf_2
X_66392_ _64782_/X _66417_/B _64785_/X _66392_/Y sky130_fd_sc_hd__nand3_4
X_78378_ _78378_/A _78374_/X _78375_/Y _78379_/A sky130_fd_sc_hd__nand3_4
X_68131_ _68097_/X _66815_/Y _68128_/X _68130_/Y _68131_/X sky130_fd_sc_hd__a211o_4
X_46509_ _46503_/Y _46445_/X _46508_/X _86731_/D sky130_fd_sc_hd__a21oi_4
X_65343_ _65289_/A _65343_/B _65343_/X sky130_fd_sc_hd__and2_4
X_77329_ _77328_/Y _82217_/Q _77325_/A _77329_/Y sky130_fd_sc_hd__nand3_4
X_62555_ _62550_/Y _62540_/X _62554_/Y _62555_/Y sky130_fd_sc_hd__a21oi_4
X_47489_ _47489_/A _47490_/A sky130_fd_sc_hd__inv_2
X_49228_ _49232_/A _46295_/X _49228_/Y sky130_fd_sc_hd__nand2_4
X_61506_ _61499_/Y _61501_/Y _61464_/X _61502_/Y _61505_/Y _61506_/X
+ sky130_fd_sc_hd__a41o_4
X_68062_ _68129_/A _68062_/X sky130_fd_sc_hd__buf_2
X_80340_ _80339_/X _82246_/D sky130_fd_sc_hd__inv_2
X_65274_ _65877_/A _65403_/A sky130_fd_sc_hd__buf_2
X_62486_ _62481_/Y _62467_/X _62485_/Y _84407_/D sky130_fd_sc_hd__a21oi_4
X_67013_ _45943_/A _67013_/X sky130_fd_sc_hd__buf_2
X_64225_ _64248_/A _64225_/B _64225_/C _64225_/X sky130_fd_sc_hd__and3_4
X_49159_ _49156_/X _50188_/B _49159_/Y sky130_fd_sc_hd__nand2_4
X_61437_ _61437_/A _61437_/B _61398_/C _61437_/Y sky130_fd_sc_hd__nand3_4
X_80271_ _84746_/Q _84138_/Q _80271_/Y sky130_fd_sc_hd__nand2_4
X_82010_ _82139_/CLK _82042_/Q _77170_/A sky130_fd_sc_hd__dfxtp_4
X_52170_ _52203_/A _52170_/X sky130_fd_sc_hd__buf_2
X_64156_ _58296_/A _64190_/B _64178_/C _64190_/D _64159_/B sky130_fd_sc_hd__nand4_4
X_61368_ _61368_/A _61368_/B _61368_/C _61368_/D _61368_/Y sky130_fd_sc_hd__nand4_4
X_51121_ _51115_/A _51121_/B _51115_/C _52811_/D _51121_/X sky130_fd_sc_hd__and4_4
X_63107_ _60466_/X _63108_/C sky130_fd_sc_hd__buf_2
X_60319_ _60525_/A _60319_/X sky130_fd_sc_hd__buf_2
X_68964_ _68961_/X _68963_/X _68846_/X _68964_/Y sky130_fd_sc_hd__a21oi_4
X_64087_ _64508_/A _64087_/X sky130_fd_sc_hd__buf_2
X_61299_ _61290_/X _61355_/A sky130_fd_sc_hd__buf_2
X_51052_ _51050_/Y _51039_/X _51051_/X _51052_/Y sky130_fd_sc_hd__a21oi_4
X_67915_ _67914_/X _67915_/B _67915_/X sky130_fd_sc_hd__and2_4
X_63038_ _63038_/A _64246_/B _63347_/C _60541_/B _63038_/X sky130_fd_sc_hd__and4_4
X_83961_ _83967_/CLK _83961_/D _83961_/Q sky130_fd_sc_hd__dfxtp_4
X_68895_ _69007_/A _68895_/X sky130_fd_sc_hd__buf_2
X_50003_ _40595_/X _50003_/X sky130_fd_sc_hd__buf_2
X_85700_ _85700_/CLK _85700_/D _85700_/Q sky130_fd_sc_hd__dfxtp_4
X_82912_ _87416_/CLK _78299_/B _82912_/Q sky130_fd_sc_hd__dfxtp_4
X_55860_ _55477_/A _56080_/C _55860_/X sky130_fd_sc_hd__and2_4
X_67846_ _87454_/Q _67751_/X _67821_/X _67845_/X _67846_/X sky130_fd_sc_hd__a211o_4
X_86680_ _86361_/CLK _86680_/D _86680_/Q sky130_fd_sc_hd__dfxtp_4
X_83892_ _87345_/CLK _83892_/D _81964_/D sky130_fd_sc_hd__dfxtp_4
X_54811_ _54806_/Y _54802_/X _54810_/X _54811_/Y sky130_fd_sc_hd__a21oi_4
X_85631_ _86592_/CLK _53463_/Y _85631_/Q sky130_fd_sc_hd__dfxtp_4
X_82843_ _82748_/CLK _82843_/D _82843_/Q sky130_fd_sc_hd__dfxtp_4
X_55791_ _55790_/X _55801_/C sky130_fd_sc_hd__buf_2
X_67777_ _67873_/A _88161_/Q _67777_/X sky130_fd_sc_hd__and2_4
X_64989_ _64729_/A _64989_/X sky130_fd_sc_hd__buf_2
X_57530_ _84985_/Q _57527_/X _57529_/Y _57530_/Y sky130_fd_sc_hd__o21ai_4
X_69516_ _69733_/A _69516_/X sky130_fd_sc_hd__buf_2
X_88350_ _87859_/CLK _40709_/Y _68892_/B sky130_fd_sc_hd__dfxtp_4
X_54742_ _85386_/Q _54729_/X _54741_/Y _54742_/Y sky130_fd_sc_hd__o21ai_4
X_66728_ _66728_/A _88141_/Q _66728_/X sky130_fd_sc_hd__and2_4
X_85562_ _85562_/CLK _53822_/Y _85562_/Q sky130_fd_sc_hd__dfxtp_4
X_51954_ _51947_/A _51954_/B _51954_/Y sky130_fd_sc_hd__nand2_4
X_82774_ _82774_/CLK _82774_/D _82966_/D sky130_fd_sc_hd__dfxtp_4
X_87301_ _87553_/CLK _87301_/D _87301_/Q sky130_fd_sc_hd__dfxtp_4
X_84513_ _84649_/CLK _84513_/D _84513_/Q sky130_fd_sc_hd__dfxtp_4
X_50905_ _50901_/Y _50902_/X _50904_/X _50905_/Y sky130_fd_sc_hd__a21oi_4
X_57461_ _57440_/X _57459_/X _57460_/Y _57461_/Y sky130_fd_sc_hd__o21ai_4
X_81725_ _80928_/CLK _81725_/D _81725_/Q sky130_fd_sc_hd__dfxtp_4
X_69447_ _87017_/Q _69277_/X _69278_/X _69446_/X _69448_/B sky130_fd_sc_hd__a211o_4
X_88281_ _88288_/CLK _41084_/Y _88281_/Q sky130_fd_sc_hd__dfxtp_4
X_54673_ _54672_/X _54674_/C sky130_fd_sc_hd__buf_2
X_66659_ _66655_/X _66657_/X _66658_/X _66659_/Y sky130_fd_sc_hd__a21oi_4
X_85493_ _85492_/CLK _85493_/D _85493_/Q sky130_fd_sc_hd__dfxtp_4
X_51885_ _85928_/Q _51873_/X _51884_/Y _51885_/Y sky130_fd_sc_hd__o21ai_4
X_59200_ _59199_/X _85745_/Q _59124_/X _59200_/X sky130_fd_sc_hd__o21a_4
X_56412_ _56418_/A _56418_/B _85204_/Q _56412_/Y sky130_fd_sc_hd__nand3_4
X_87232_ _87758_/CLK _43856_/Y _87232_/Q sky130_fd_sc_hd__dfxtp_4
X_53624_ _52103_/A _53620_/B _53620_/C _53624_/X sky130_fd_sc_hd__and3_4
X_84444_ _84452_/CLK _84444_/D _78067_/B sky130_fd_sc_hd__dfxtp_4
X_50836_ _50822_/A _51350_/B _50836_/Y sky130_fd_sc_hd__nand2_4
X_57392_ _57359_/A _57392_/B _57372_/X _57392_/Y sky130_fd_sc_hd__nor3_4
X_81656_ _81697_/CLK _81688_/Q _76470_/A sky130_fd_sc_hd__dfxtp_4
X_69378_ _69374_/X _69377_/X _69142_/X _69378_/Y sky130_fd_sc_hd__a21oi_4
X_59131_ _59131_/A _59068_/B _59131_/Y sky130_fd_sc_hd__nor2_4
X_56343_ _56345_/A _56345_/B _85228_/Q _56343_/Y sky130_fd_sc_hd__nand3_4
X_80607_ _80607_/A _80607_/B _80607_/X sky130_fd_sc_hd__xor2_4
X_68329_ _68319_/X _68005_/Y _68326_/X _68328_/Y _68329_/X sky130_fd_sc_hd__a211o_4
X_87163_ _88175_/CLK _87163_/D _87163_/Q sky130_fd_sc_hd__dfxtp_4
X_53555_ _53553_/Y _53537_/X _53554_/X _85614_/D sky130_fd_sc_hd__a21oi_4
X_84375_ _84375_/CLK _84375_/D _62873_/C sky130_fd_sc_hd__dfxtp_4
X_50767_ _86137_/Q _50742_/X _50766_/Y _50767_/Y sky130_fd_sc_hd__o21ai_4
X_81587_ _81587_/CLK _84187_/Q _76809_/A sky130_fd_sc_hd__dfxtp_4
X_86114_ _86121_/CLK _86114_/D _86114_/Q sky130_fd_sc_hd__dfxtp_4
X_40520_ _40519_/Y _40520_/X sky130_fd_sc_hd__buf_2
X_52506_ _52448_/A _46441_/Y _52506_/Y sky130_fd_sc_hd__nand2_4
X_59062_ _59013_/X _85756_/Q _59037_/X _59062_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_10_472_0_CLK clkbuf_9_236_0_CLK/X _86697_/CLK sky130_fd_sc_hd__clkbuf_1
X_71340_ _71462_/B _71485_/B sky130_fd_sc_hd__inv_2
X_83326_ _83322_/CLK _83326_/D _56682_/A sky130_fd_sc_hd__dfxtp_4
X_80538_ _84769_/Q _84161_/Q _80538_/X sky130_fd_sc_hd__xor2_4
X_56274_ _56273_/X _56274_/X sky130_fd_sc_hd__buf_2
X_87094_ _88268_/CLK _44468_/X _87094_/Q sky130_fd_sc_hd__dfxtp_4
X_53486_ _53478_/A _73717_/A _53486_/Y sky130_fd_sc_hd__nand2_4
X_50698_ _86151_/Q _50680_/X _50697_/Y _50698_/Y sky130_fd_sc_hd__o21ai_4
X_58013_ _86636_/Q _58039_/B _58013_/Y sky130_fd_sc_hd__nor2_4
X_55225_ _45861_/A _44058_/A _55140_/A _55224_/X _55225_/X sky130_fd_sc_hd__a211o_4
X_86045_ _86045_/CLK _51257_/Y _86045_/Q sky130_fd_sc_hd__dfxtp_4
X_40451_ _40421_/X _81171_/Q _40450_/X _40451_/X sky130_fd_sc_hd__o21a_4
X_52437_ _52435_/Y _52430_/X _52436_/Y _85823_/D sky130_fd_sc_hd__a21boi_4
X_71271_ _71171_/A _71276_/B _71276_/C _70656_/D _71271_/Y sky130_fd_sc_hd__nand4_4
X_83257_ _86282_/CLK _83257_/D _83257_/Q sky130_fd_sc_hd__dfxtp_4
X_80469_ _80457_/A _80456_/Y _80468_/X _80469_/X sky130_fd_sc_hd__a21o_4
X_73010_ _73132_/A _85880_/Q _73010_/X sky130_fd_sc_hd__and2_4
X_70222_ _70209_/X _83832_/Q _70221_/X _70222_/X sky130_fd_sc_hd__a21o_4
X_82208_ _82965_/CLK _82208_/D _82208_/Q sky130_fd_sc_hd__dfxtp_4
X_43170_ _43170_/A _43170_/Y sky130_fd_sc_hd__inv_2
X_55156_ _55151_/X _55155_/X _44108_/X _55156_/X sky130_fd_sc_hd__a21o_4
X_52368_ _65155_/B _52347_/X _52367_/Y _52368_/Y sky130_fd_sc_hd__o21ai_4
X_40382_ _40321_/A _40586_/A sky130_fd_sc_hd__buf_2
X_83188_ _83188_/CLK _72692_/X _83188_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_487_0_CLK clkbuf_9_243_0_CLK/X _86713_/CLK sky130_fd_sc_hd__clkbuf_1
X_54107_ _85502_/Q _53431_/X _54106_/Y _54107_/Y sky130_fd_sc_hd__o21ai_4
X_42121_ _42120_/X _42116_/X _41082_/X _88025_/Q _42117_/X _42122_/A
+ sky130_fd_sc_hd__o32ai_4
X_51319_ _51317_/Y _51313_/X _51318_/X _51319_/Y sky130_fd_sc_hd__a21oi_4
X_70153_ _70153_/A _70153_/Y sky130_fd_sc_hd__inv_2
X_82139_ _82139_/CLK _77958_/X _82095_/D sky130_fd_sc_hd__dfxtp_4
X_55087_ _55083_/A _55104_/B _55083_/C _47757_/A _55087_/X sky130_fd_sc_hd__and4_4
X_59964_ _59964_/A _59964_/Y sky130_fd_sc_hd__inv_2
X_52299_ _52299_/A _48955_/X _52299_/Y sky130_fd_sc_hd__nand2_4
X_87996_ _87487_/CLK _42178_/Y _87996_/Q sky130_fd_sc_hd__dfxtp_4
X_42052_ _42013_/A _42052_/X sky130_fd_sc_hd__buf_2
X_58915_ _58891_/X _86086_/Q _58914_/X _58915_/Y sky130_fd_sc_hd__o21ai_4
X_54038_ _85518_/Q _54035_/X _54037_/Y _54038_/Y sky130_fd_sc_hd__o21ai_4
X_74961_ _74960_/Y _74961_/B _74962_/B sky130_fd_sc_hd__and2_4
X_70084_ _83854_/Q _70067_/X _70083_/X _83854_/D sky130_fd_sc_hd__a21bo_4
X_86947_ _88215_/CLK _86947_/D _86947_/Q sky130_fd_sc_hd__dfxtp_4
X_59895_ _59881_/X _59884_/X _59927_/A _62288_/A sky130_fd_sc_hd__a21oi_4
X_41003_ _40429_/X _82293_/Q _41002_/X _41003_/X sky130_fd_sc_hd__o21a_4
X_76700_ _76692_/Y _76700_/Y sky130_fd_sc_hd__inv_2
X_73912_ _73913_/B _73913_/C _73911_/X _73912_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_10_410_0_CLK clkbuf_9_205_0_CLK/X _83521_/CLK sky130_fd_sc_hd__clkbuf_1
X_58846_ _58846_/A _58846_/X sky130_fd_sc_hd__buf_2
X_46860_ _46720_/A _46860_/X sky130_fd_sc_hd__buf_2
X_77680_ _77676_/X _77677_/Y _77679_/Y _77680_/X sky130_fd_sc_hd__a21o_4
X_74892_ _81128_/D _80840_/Q _74900_/A sky130_fd_sc_hd__nand2_4
X_86878_ _86878_/CLK _86878_/D _63017_/B sky130_fd_sc_hd__dfxtp_4
X_45811_ _45811_/A _45811_/Y sky130_fd_sc_hd__inv_2
X_76631_ _76640_/A _76640_/B _76639_/A sky130_fd_sc_hd__nand2_4
X_85829_ _86749_/CLK _52408_/Y _65324_/B sky130_fd_sc_hd__dfxtp_4
X_73843_ _68669_/B _73674_/X _73819_/X _73842_/Y _73843_/X sky130_fd_sc_hd__a211o_4
X_46791_ _46790_/Y _46791_/X sky130_fd_sc_hd__buf_2
X_58777_ _58748_/X _58775_/Y _58776_/Y _58766_/X _58752_/X _58777_/X
+ sky130_fd_sc_hd__o32a_4
X_55989_ _56104_/A _56177_/A sky130_fd_sc_hd__buf_2
X_48530_ _48914_/A _82354_/Q _48530_/Y sky130_fd_sc_hd__nor2_4
X_79350_ _58769_/Y _66450_/Y _79349_/Y _79350_/X sky130_fd_sc_hd__o21a_4
X_45742_ _45737_/X _45741_/X _45678_/X _45742_/X sky130_fd_sc_hd__a21o_4
X_57728_ _57726_/X _86016_/Q _57727_/X _57728_/Y sky130_fd_sc_hd__o21ai_4
X_76562_ _76584_/D _76562_/Y sky130_fd_sc_hd__inv_2
X_42954_ _42488_/A _42954_/X sky130_fd_sc_hd__buf_2
X_73774_ _43620_/Y _73597_/X _73772_/X _73773_/Y _73774_/X sky130_fd_sc_hd__a211o_4
X_70986_ _70986_/A _70990_/C sky130_fd_sc_hd__buf_2
X_78301_ _78301_/A _82472_/Q _78302_/B sky130_fd_sc_hd__nand2_4
Xclkbuf_10_425_0_CLK clkbuf_9_212_0_CLK/X _82425_/CLK sky130_fd_sc_hd__clkbuf_1
X_75513_ _75505_/Y _75538_/B _75513_/X sky130_fd_sc_hd__xor2_4
X_41905_ _50523_/A _51584_/A sky130_fd_sc_hd__buf_2
X_48461_ _48461_/A _48485_/B sky130_fd_sc_hd__buf_2
X_72725_ _72725_/A _72725_/X sky130_fd_sc_hd__buf_2
X_79281_ _79277_/X _79280_/Y _79281_/X sky130_fd_sc_hd__xor2_4
X_45673_ _45673_/A _45793_/B _45673_/Y sky130_fd_sc_hd__nor2_4
X_57659_ _83759_/Q _57659_/Y sky130_fd_sc_hd__inv_2
X_76493_ _76474_/A _76471_/Y _76473_/A _76494_/A sky130_fd_sc_hd__o21a_4
X_42885_ _42885_/A _87669_/D sky130_fd_sc_hd__inv_2
X_47412_ _47404_/A _53033_/B _47412_/Y sky130_fd_sc_hd__nand2_4
X_78232_ _78253_/B _82496_/Q _78252_/A sky130_fd_sc_hd__xor2_4
X_44624_ _44624_/A _44714_/A sky130_fd_sc_hd__buf_2
X_75444_ _75443_/A _80955_/D _75445_/A sky130_fd_sc_hd__nand2_4
X_41836_ _41824_/X _41825_/X _40480_/X _67003_/B _41835_/X _41837_/A
+ sky130_fd_sc_hd__o32ai_4
X_48392_ _48392_/A _48391_/X _48392_/Y sky130_fd_sc_hd__nand2_4
X_60670_ _63398_/A _60671_/C sky130_fd_sc_hd__inv_2
X_72656_ _72656_/A _72656_/B _72656_/C _72656_/Y sky130_fd_sc_hd__nand3_4
X_47343_ _47343_/A _47344_/A sky130_fd_sc_hd__inv_2
X_59329_ _58923_/A _59329_/X sky130_fd_sc_hd__buf_2
X_71607_ _71626_/A _70573_/B _70568_/D _71606_/X _71607_/Y sky130_fd_sc_hd__nor4_4
X_78163_ _78151_/Y _78162_/X _78166_/A sky130_fd_sc_hd__nand2_4
X_44555_ _44530_/A _44555_/X sky130_fd_sc_hd__buf_2
X_75375_ _75376_/A _75376_/B _75375_/Y sky130_fd_sc_hd__nor2_4
X_41767_ _40621_/X _41427_/A _41766_/X _41767_/Y sky130_fd_sc_hd__o21ai_4
X_72587_ _61260_/X _72597_/B _61319_/X _72607_/C _60529_/A _72587_/Y
+ sky130_fd_sc_hd__a41oi_4
Xclkbuf_1_1_0_CLK clkbuf_0_CLK/X clkbuf_1_1_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_77114_ _77106_/A _77114_/B _82288_/D _77115_/A sky130_fd_sc_hd__nand3_4
X_43506_ _43528_/A _43506_/X sky130_fd_sc_hd__buf_2
X_62340_ _62120_/A _62342_/A sky130_fd_sc_hd__buf_2
X_74326_ _70313_/C _74314_/X _74325_/Y _83097_/D sky130_fd_sc_hd__a21bo_4
X_40718_ _40717_/X _40793_/A sky130_fd_sc_hd__buf_2
X_47274_ _54645_/D _52954_/D sky130_fd_sc_hd__buf_2
X_71538_ _71531_/X _83465_/Q _71537_/Y _83465_/D sky130_fd_sc_hd__a21o_4
X_78094_ _78090_/Y _78093_/Y _78096_/B sky130_fd_sc_hd__xnor2_4
X_44486_ _44486_/A _44486_/Y sky130_fd_sc_hd__inv_2
X_41698_ _41697_/X _41682_/X _67634_/B _41684_/X _88167_/D sky130_fd_sc_hd__a2bb2o_4
X_49013_ _49008_/Y _48985_/X _49012_/X _86453_/D sky130_fd_sc_hd__a21oi_4
X_46225_ _46224_/X _46098_/A _46214_/C _46214_/D _46225_/Y sky130_fd_sc_hd__nand4_4
XPHY_370 sky130_fd_sc_hd__decap_3
X_77045_ _77054_/A _82281_/D _77045_/X sky130_fd_sc_hd__xor2_4
X_43437_ _41570_/X _43431_/X _87422_/Q _43432_/X _43437_/X sky130_fd_sc_hd__a2bb2o_4
X_62271_ _62304_/A _58232_/X _62244_/C _62244_/D _62271_/X sky130_fd_sc_hd__and4_4
X_74257_ _72730_/X _84963_/Q _74021_/X _74256_/X _74258_/B sky130_fd_sc_hd__a211o_4
X_40649_ _40585_/X _82870_/Q _40648_/X _40649_/Y sky130_fd_sc_hd__o21ai_4
XPHY_381 sky130_fd_sc_hd__decap_3
X_71469_ _71464_/X _83488_/Q _71468_/X _83488_/D sky130_fd_sc_hd__a21o_4
XPHY_392 sky130_fd_sc_hd__decap_3
X_64010_ _64006_/X _63994_/X _64009_/Y _64010_/Y sky130_fd_sc_hd__a21oi_4
X_61222_ _72564_/A _61250_/B sky130_fd_sc_hd__buf_2
X_73208_ _73062_/X _86192_/Q _73205_/X _73207_/X _73208_/X sky130_fd_sc_hd__a211o_4
X_46156_ _46155_/X _46158_/B sky130_fd_sc_hd__buf_2
X_43368_ _43367_/X _43350_/X _41387_/X _87456_/Q _43353_/X _43369_/A
+ sky130_fd_sc_hd__o32ai_4
X_74188_ _74185_/X _74187_/X _73602_/X _74188_/X sky130_fd_sc_hd__a21o_4
X_45107_ _45107_/A _45108_/A sky130_fd_sc_hd__inv_2
X_42319_ _42397_/A _42319_/X sky130_fd_sc_hd__buf_2
X_73139_ _72963_/X _83067_/Q _73015_/X _73138_/X _73139_/X sky130_fd_sc_hd__a211o_4
X_61153_ _61153_/A _61108_/Y _61153_/C _61272_/B sky130_fd_sc_hd__nand3_4
X_46087_ _46087_/A _46089_/C sky130_fd_sc_hd__inv_2
X_43299_ _41199_/X _43287_/X _87491_/Q _43288_/X _43299_/X sky130_fd_sc_hd__a2bb2o_4
X_78996_ _82823_/Q _82535_/Q _78997_/B sky130_fd_sc_hd__xnor2_4
X_60104_ _59971_/X _60099_/X _60102_/Y _60072_/Y _60103_/Y _84661_/D
+ sky130_fd_sc_hd__a41oi_4
X_49915_ _49915_/A _49915_/X sky130_fd_sc_hd__buf_2
X_45038_ _55908_/B _44979_/X _45012_/X _45038_/X sky130_fd_sc_hd__o21a_4
X_65961_ _65614_/A _65961_/X sky130_fd_sc_hd__buf_2
X_61084_ _64367_/A _64249_/A sky130_fd_sc_hd__buf_2
X_77947_ _77935_/Y _77946_/A _82072_/Q _81944_/D _77947_/X sky130_fd_sc_hd__a2bb2o_4
X_67700_ _67793_/A _67700_/B _67700_/X sky130_fd_sc_hd__and2_4
X_64912_ _64901_/Y _64911_/Y _64912_/Y sky130_fd_sc_hd__nand2_4
X_60035_ _60034_/X _64689_/A sky130_fd_sc_hd__buf_2
X_49846_ _49851_/A _49851_/B _49830_/C _53058_/D _49846_/X sky130_fd_sc_hd__and4_4
X_68680_ _88007_/Q _68650_/X _68651_/X _68679_/X _68680_/X sky130_fd_sc_hd__a211o_4
X_65892_ _65807_/A _86466_/Q _65892_/X sky130_fd_sc_hd__and2_4
X_77878_ _82065_/Q _77876_/Y _77877_/X _77878_/Y sky130_fd_sc_hd__o21ai_4
X_67631_ _67627_/X _67630_/X _67561_/X _67631_/X sky130_fd_sc_hd__a21o_4
X_79617_ _79603_/Y _79609_/A _79616_/Y _79619_/A sky130_fd_sc_hd__a21o_4
X_64843_ _64839_/Y _64814_/X _64842_/Y _84225_/D sky130_fd_sc_hd__a21o_4
X_76829_ _76829_/A _76828_/Y _76837_/A sky130_fd_sc_hd__xor2_4
X_49777_ _51012_/A _49861_/A sky130_fd_sc_hd__buf_2
X_46989_ _82394_/Q _46990_/A sky130_fd_sc_hd__inv_2
X_48728_ _53636_/A _48099_/X _48761_/C _48728_/X sky130_fd_sc_hd__and3_4
X_67562_ _67557_/X _67560_/X _67561_/X _67562_/X sky130_fd_sc_hd__a21o_4
X_79548_ _79545_/B _79534_/Y _79542_/Y _79548_/Y sky130_fd_sc_hd__a21oi_4
X_64774_ _64577_/X _83307_/Q _64772_/X _64773_/X _64775_/B sky130_fd_sc_hd__a211o_4
X_61986_ _63561_/B _61924_/B _61971_/C _61971_/D _61986_/Y sky130_fd_sc_hd__nand4_4
X_69301_ _68742_/A _69302_/A sky130_fd_sc_hd__buf_2
X_66513_ _84108_/Q _66514_/C sky130_fd_sc_hd__inv_2
Xclkbuf_8_52_0_CLK clkbuf_8_53_0_CLK/A clkbuf_8_52_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_63725_ _60855_/X _64189_/D sky130_fd_sc_hd__buf_2
X_48659_ _48659_/A _48660_/A sky130_fd_sc_hd__inv_2
X_60937_ _60891_/Y _60937_/B _60988_/A _60938_/A sky130_fd_sc_hd__nand3_4
X_67493_ _67305_/X _67484_/Y _67390_/X _67492_/Y _67493_/X sky130_fd_sc_hd__a211o_4
X_79479_ _79505_/A _79489_/A sky130_fd_sc_hd__inv_2
X_81510_ _84087_/CLK _76200_/B _75950_/A sky130_fd_sc_hd__dfxtp_4
X_69232_ _69478_/A _69232_/X sky130_fd_sc_hd__buf_2
X_66444_ _84122_/Q _66445_/C sky130_fd_sc_hd__inv_2
X_51670_ _51666_/Y _51667_/X _51669_/X _51670_/Y sky130_fd_sc_hd__a21oi_4
X_63656_ _59427_/Y _63626_/X _61630_/A _63627_/X _63656_/X sky130_fd_sc_hd__a2bb2o_4
X_82490_ _82491_/CLK _78676_/X _78199_/B sky130_fd_sc_hd__dfxtp_4
X_60868_ _60867_/Y _60930_/A sky130_fd_sc_hd__buf_2
XPHY_18 sky130_fd_sc_hd__decap_3
XPHY_29 sky130_fd_sc_hd__decap_3
X_50621_ _50618_/Y _50619_/X _50620_/Y _50621_/Y sky130_fd_sc_hd__a21boi_4
X_62607_ _62603_/Y _62593_/X _62606_/Y _84397_/D sky130_fd_sc_hd__a21oi_4
X_81441_ _83940_/CLK _81473_/Q _76146_/B sky130_fd_sc_hd__dfxtp_4
X_69163_ _69067_/A _87793_/Q _69163_/X sky130_fd_sc_hd__and2_4
X_66375_ _65949_/X _66367_/B _65952_/X _66375_/Y sky130_fd_sc_hd__nand3_4
X_63587_ _61548_/B _63548_/X _63585_/X _63586_/Y _63587_/X sky130_fd_sc_hd__a211o_4
X_60799_ _60798_/X _60736_/X _63374_/A _60767_/X _60758_/X _60799_/X
+ sky130_fd_sc_hd__a2111o_4
Xclkbuf_8_67_0_CLK clkbuf_8_67_0_CLK/A clkbuf_8_67_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_68114_ _66727_/X _66729_/X _68106_/X _68114_/Y sky130_fd_sc_hd__a21oi_4
X_53340_ _53337_/Y _53328_/X _53339_/X _85652_/D sky130_fd_sc_hd__a21oi_4
X_65326_ _65669_/A _65326_/X sky130_fd_sc_hd__buf_2
X_84160_ _84161_/CLK _84160_/D _84160_/Q sky130_fd_sc_hd__dfxtp_4
X_50552_ _48702_/A _50552_/B _50552_/C _50552_/X sky130_fd_sc_hd__and3_4
X_62538_ _61590_/B _62462_/X _62507_/X _62478_/X _62537_/X _62538_/X
+ sky130_fd_sc_hd__a41o_4
X_81372_ _81482_/CLK _76884_/X _81372_/Q sky130_fd_sc_hd__dfxtp_4
X_69094_ _69091_/X _69093_/X _69094_/Y sky130_fd_sc_hd__nand2_4
X_83111_ _82998_/CLK _74292_/X _70273_/A sky130_fd_sc_hd__dfxtp_4
X_68045_ _87445_/Q _67953_/X _67954_/X _68044_/X _68045_/X sky130_fd_sc_hd__a211o_4
X_80323_ _80323_/A _80323_/B _80324_/A sky130_fd_sc_hd__xor2_4
X_53271_ _85664_/Q _53268_/X _53270_/Y _53271_/Y sky130_fd_sc_hd__o21ai_4
X_65257_ _65791_/A _65258_/A sky130_fd_sc_hd__buf_2
X_84091_ _81507_/CLK _66924_/X _80915_/D sky130_fd_sc_hd__dfxtp_4
X_50483_ _50556_/A _52188_/B _50483_/Y sky130_fd_sc_hd__nand2_4
X_62469_ _62466_/Y _62467_/X _62468_/Y _62469_/Y sky130_fd_sc_hd__a21oi_4
X_55010_ _55008_/Y _54998_/X _55009_/X _55010_/Y sky130_fd_sc_hd__a21oi_4
X_52222_ _52247_/A _52223_/C sky130_fd_sc_hd__buf_2
X_64208_ _64545_/A _61298_/B _64545_/C _64208_/Y sky130_fd_sc_hd__nand3_4
X_83042_ _85428_/CLK _74534_/Y _83042_/Q sky130_fd_sc_hd__dfxtp_4
X_80254_ _84952_/Q _65449_/C _80254_/Y sky130_fd_sc_hd__nand2_4
X_65188_ _65185_/X _65187_/X _64989_/X _65188_/X sky130_fd_sc_hd__a21o_4
X_52153_ _52215_/A _52168_/A sky130_fd_sc_hd__buf_2
X_64139_ _64508_/A _64187_/B sky130_fd_sc_hd__buf_2
X_87850_ _87850_/CLK _42482_/Y _68588_/A sky130_fd_sc_hd__dfxtp_4
X_80185_ _84947_/Q _65531_/C _80187_/A sky130_fd_sc_hd__xor2_4
X_69996_ _69993_/X _69995_/X _70021_/C _69996_/Y sky130_fd_sc_hd__nand3_4
X_51104_ _86073_/Q _51101_/X _51103_/Y _51104_/Y sky130_fd_sc_hd__o21ai_4
X_86801_ _87484_/CLK _46036_/X _66691_/B sky130_fd_sc_hd__dfxtp_4
X_52084_ _52082_/Y _52066_/X _52083_/Y _85892_/D sky130_fd_sc_hd__a21boi_4
X_56961_ _56960_/X _45549_/A _56953_/X _56961_/Y sky130_fd_sc_hd__nor3_4
X_68947_ _68377_/A _69485_/A sky130_fd_sc_hd__buf_2
X_87781_ _87782_/CLK _42664_/Y _87781_/Q sky130_fd_sc_hd__dfxtp_4
X_84993_ _85826_/CLK _57492_/Y _84993_/Q sky130_fd_sc_hd__dfxtp_4
X_58700_ _58700_/A _58688_/B _58700_/Y sky130_fd_sc_hd__nor2_4
X_55912_ _55909_/X _55911_/X _44115_/A _55912_/X sky130_fd_sc_hd__a21o_4
X_51035_ _51029_/A _51029_/B _51045_/C _52724_/D _51035_/X sky130_fd_sc_hd__and4_4
X_86732_ _86733_/CLK _46499_/Y _86732_/Q sky130_fd_sc_hd__dfxtp_4
X_83944_ _83944_/CLK _83944_/D _83944_/Q sky130_fd_sc_hd__dfxtp_4
X_59680_ _59680_/A _59754_/D _59687_/A _59680_/Y sky130_fd_sc_hd__nand3_4
X_56892_ _46173_/X _56892_/B _56892_/C _73939_/A _56892_/Y sky130_fd_sc_hd__nand4_4
X_68878_ _68660_/X _68878_/X sky130_fd_sc_hd__buf_2
X_58631_ _58631_/A _58631_/X sky130_fd_sc_hd__buf_2
X_55843_ _55843_/A _85296_/Q _55843_/X sky130_fd_sc_hd__and2_4
X_67829_ _67664_/X _67815_/Y _67747_/X _67828_/Y _67829_/X sky130_fd_sc_hd__a211o_4
X_86663_ _86342_/CLK _47172_/Y _86663_/Q sky130_fd_sc_hd__dfxtp_4
X_83875_ _82557_/CLK _70004_/X _82555_/D sky130_fd_sc_hd__dfxtp_4
X_88402_ _86834_/CLK _88402_/D _88402_/Q sky130_fd_sc_hd__dfxtp_4
X_85614_ _86222_/CLK _85614_/D _85614_/Q sky130_fd_sc_hd__dfxtp_4
X_70840_ _50893_/B _70831_/X _70839_/Y _70840_/Y sky130_fd_sc_hd__o21ai_4
X_58562_ _58562_/A _58973_/B _58562_/Y sky130_fd_sc_hd__nand2_4
X_82826_ _83167_/CLK _79275_/X _82826_/Q sky130_fd_sc_hd__dfxtp_4
X_55774_ _55711_/X _55774_/B _55774_/X sky130_fd_sc_hd__and2_4
X_86594_ _85955_/CLK _86594_/D _72476_/A sky130_fd_sc_hd__dfxtp_4
X_52986_ _52999_/A _52986_/B _52986_/Y sky130_fd_sc_hd__nand2_4
X_57513_ _57499_/A _73692_/A _57513_/Y sky130_fd_sc_hd__nand2_4
X_88333_ _84970_/CLK _88333_/D _88333_/Q sky130_fd_sc_hd__dfxtp_4
X_54725_ _54616_/X _54748_/A sky130_fd_sc_hd__buf_2
X_85545_ _85536_/CLK _85545_/D _85545_/Q sky130_fd_sc_hd__dfxtp_4
X_51937_ _51941_/A _48178_/X _51937_/Y sky130_fd_sc_hd__nand2_4
X_70771_ _70771_/A _70867_/A sky130_fd_sc_hd__buf_2
X_58493_ _83411_/Q _58493_/Y sky130_fd_sc_hd__inv_2
X_82757_ _86697_/CLK _78355_/Y _82757_/Q sky130_fd_sc_hd__dfxtp_4
X_72510_ _72607_/B _72516_/A _72510_/C _72515_/D _72510_/Y sky130_fd_sc_hd__nand4_4
X_57444_ _57441_/X _56801_/X _57443_/X _57444_/X sky130_fd_sc_hd__o21a_4
X_81708_ _81755_/CLK _81708_/D _41223_/A sky130_fd_sc_hd__dfxtp_4
X_88264_ _88268_/CLK _41170_/X _68658_/B sky130_fd_sc_hd__dfxtp_4
X_42670_ _41032_/X _42652_/X _87778_/Q _42653_/X _87778_/D sky130_fd_sc_hd__a2bb2o_4
X_54656_ _54245_/A _54656_/X sky130_fd_sc_hd__buf_2
X_73490_ _73485_/X _73488_/X _73489_/X _73494_/A sky130_fd_sc_hd__a21o_4
X_85476_ _84926_/CLK _54256_/Y _85476_/Q sky130_fd_sc_hd__dfxtp_4
X_51868_ _85931_/Q _51846_/X _51867_/Y _51868_/Y sky130_fd_sc_hd__o21ai_4
X_82688_ _84111_/CLK _82700_/Q _82688_/Q sky130_fd_sc_hd__dfxtp_4
X_87215_ _87471_/CLK _43888_/X _67440_/B sky130_fd_sc_hd__dfxtp_4
X_53607_ _85603_/Q _53586_/X _53606_/Y _53607_/Y sky130_fd_sc_hd__o21ai_4
X_41621_ _41620_/X _41621_/X sky130_fd_sc_hd__buf_2
X_72441_ _72389_/X _85670_/Q _72422_/X _72441_/X sky130_fd_sc_hd__o21a_4
X_84427_ _84426_/CLK _84427_/D _78050_/B sky130_fd_sc_hd__dfxtp_4
X_50819_ _50991_/A _50819_/X sky130_fd_sc_hd__buf_2
X_57375_ _73040_/A _73476_/A sky130_fd_sc_hd__buf_2
X_81639_ _81582_/CLK _81671_/Q _76234_/A sky130_fd_sc_hd__dfxtp_4
X_88195_ _87421_/CLK _88195_/D _66966_/B sky130_fd_sc_hd__dfxtp_4
X_54587_ _54578_/A _54587_/B _54587_/Y sky130_fd_sc_hd__nand2_4
X_51799_ _51797_/Y _51793_/X _51798_/X _85944_/D sky130_fd_sc_hd__a21oi_4
X_59114_ _59102_/Y _58857_/X _59109_/X _59113_/X _59114_/Y sky130_fd_sc_hd__a22oi_4
X_44340_ _41681_/X _44326_/X _87158_/Q _44327_/X _87158_/D sky130_fd_sc_hd__a2bb2o_4
X_56326_ _56332_/A _56335_/B _55855_/B _56326_/Y sky130_fd_sc_hd__nand3_4
X_75160_ _75155_/Y _75161_/B _75159_/Y _75162_/A sky130_fd_sc_hd__a21o_4
X_87146_ _87144_/CLK _44366_/X _87146_/Q sky130_fd_sc_hd__dfxtp_4
X_41552_ _41552_/A _41552_/X sky130_fd_sc_hd__buf_2
X_53538_ _50314_/A _53474_/B _53492_/X _53538_/X sky130_fd_sc_hd__and3_4
X_72372_ _72287_/X _85324_/Q _72324_/X _72372_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_3_6_1_CLK clkbuf_3_6_1_CLK/A clkbuf_3_6_1_CLK/X sky130_fd_sc_hd__clkbuf_1
X_84358_ _84358_/CLK _63046_/X _79476_/A sky130_fd_sc_hd__dfxtp_4
X_74111_ _74105_/X _74110_/X _74085_/X _74111_/X sky130_fd_sc_hd__a21o_4
X_40503_ _40502_/Y _40503_/Y sky130_fd_sc_hd__inv_2
X_59045_ _86685_/Q _59008_/B _59045_/Y sky130_fd_sc_hd__nor2_4
X_71323_ _71323_/A _71314_/B _71297_/X _71323_/Y sky130_fd_sc_hd__nand3_4
X_83309_ _85547_/CLK _71980_/Y _83309_/Q sky130_fd_sc_hd__dfxtp_4
X_56257_ _56139_/X _56255_/X _56256_/Y _56257_/Y sky130_fd_sc_hd__o21ai_4
X_44271_ _44270_/X _72896_/B sky130_fd_sc_hd__buf_2
X_75091_ _75091_/A _75091_/B _75102_/A _75107_/A sky130_fd_sc_hd__nand3_4
X_87077_ _87077_/CLK _87077_/D _87077_/Q sky130_fd_sc_hd__dfxtp_4
X_53469_ _85630_/Q _53466_/X _53468_/Y _53469_/Y sky130_fd_sc_hd__o21ai_4
X_41483_ _81180_/Q _41523_/B _41483_/X sky130_fd_sc_hd__or2_4
X_84289_ _84287_/CLK _84289_/D _84289_/Q sky130_fd_sc_hd__dfxtp_4
X_46010_ _45994_/X _46001_/X _40500_/X _67107_/B _45995_/X _46011_/A
+ sky130_fd_sc_hd__o32ai_4
X_55208_ _55177_/A _55208_/B _55208_/Y sky130_fd_sc_hd__nor2_4
X_43222_ _43196_/X _43207_/X _40977_/X _87531_/Q _43212_/X _43223_/A
+ sky130_fd_sc_hd__o32ai_4
X_74042_ _74039_/X _74041_/X _74019_/X _74045_/A sky130_fd_sc_hd__a21o_4
X_86028_ _86029_/CLK _51349_/Y _65147_/B sky130_fd_sc_hd__dfxtp_4
X_40434_ _40434_/A _40434_/Y sky130_fd_sc_hd__inv_2
X_71254_ _71241_/A _71258_/A sky130_fd_sc_hd__buf_2
X_56188_ _56255_/A _56188_/X sky130_fd_sc_hd__buf_2
X_70205_ _70214_/A _70214_/B _70205_/C _70204_/X _70205_/X sky130_fd_sc_hd__and4_4
X_43153_ _43129_/X _43130_/X _40845_/X _43152_/Y _43142_/X _43153_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55139_ _55132_/X _55136_/X _55138_/X _55139_/X sky130_fd_sc_hd__a21o_4
X_78850_ _78874_/B _78849_/Y _78851_/B sky130_fd_sc_hd__xnor2_4
X_40365_ _48135_/A _40365_/X sky130_fd_sc_hd__buf_2
X_71185_ _71041_/X _71185_/B _70966_/A _74518_/D _71185_/Y sky130_fd_sc_hd__nand4_4
X_42104_ _41912_/A _42104_/X sky130_fd_sc_hd__buf_2
X_77801_ _77799_/X _77788_/X _77800_/X _77801_/X sky130_fd_sc_hd__a21o_4
X_70136_ _83506_/Q _83154_/Q _83499_/Q _83147_/Q _70139_/B sky130_fd_sc_hd__a22oi_4
X_47961_ _47988_/A _50293_/B _47961_/Y sky130_fd_sc_hd__nand2_4
X_59947_ _59929_/C _62198_/B sky130_fd_sc_hd__buf_2
X_43084_ _43083_/Y _87582_/D sky130_fd_sc_hd__inv_2
X_78781_ _78772_/A _78746_/Y _78773_/X _78782_/A sky130_fd_sc_hd__o21ai_4
X_75993_ _75984_/Y _75991_/Y _75992_/Y _75993_/X sky130_fd_sc_hd__o21a_4
X_87979_ _88232_/CLK _42211_/X _87979_/Q sky130_fd_sc_hd__dfxtp_4
X_49700_ _59372_/B _49687_/X _49699_/Y _49700_/Y sky130_fd_sc_hd__o21ai_4
X_46912_ _52744_/B _46912_/X sky130_fd_sc_hd__buf_2
X_42035_ _41998_/A _42035_/X sky130_fd_sc_hd__buf_2
X_77732_ _77731_/Y _77732_/B _77732_/Y sky130_fd_sc_hd__nand2_4
X_74944_ _81135_/D _74945_/B _74944_/Y sky130_fd_sc_hd__nor2_4
X_70067_ _70048_/A _70067_/X sky130_fd_sc_hd__buf_2
X_47892_ _65977_/B _47840_/X _47891_/Y _47892_/Y sky130_fd_sc_hd__o21ai_4
X_59878_ _59877_/X _59564_/B _59551_/A _60418_/D sky130_fd_sc_hd__a21boi_4
X_49631_ _49628_/Y _49623_/X _49630_/X _86352_/D sky130_fd_sc_hd__a21oi_4
X_46843_ _86697_/Q _46813_/X _46842_/Y _46843_/Y sky130_fd_sc_hd__o21ai_4
X_58829_ _58698_/A _58872_/A sky130_fd_sc_hd__buf_2
Xclkbuf_9_470_0_CLK clkbuf_9_471_0_CLK/A clkbuf_9_470_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_77663_ _77622_/A _77596_/A _77621_/A _77645_/B _77663_/X sky130_fd_sc_hd__and4_4
X_74875_ _81127_/D _74875_/B _74897_/B sky130_fd_sc_hd__xor2_4
X_79402_ _84806_/Q _84126_/Q _79402_/Y sky130_fd_sc_hd__nand2_4
X_76614_ _76614_/A _76614_/B _76614_/C _76602_/Y _76614_/X sky130_fd_sc_hd__and4_4
Xclkbuf_10_364_0_CLK clkbuf_9_182_0_CLK/X _85993_/CLK sky130_fd_sc_hd__clkbuf_1
X_61840_ _58248_/A _61824_/X _61838_/X _61790_/X _61839_/X _61840_/X
+ sky130_fd_sc_hd__a41o_4
X_49562_ _49559_/Y _49541_/X _49561_/X _49562_/Y sky130_fd_sc_hd__a21oi_4
X_73826_ _44697_/Y _73728_/X _73825_/Y _73838_/C sky130_fd_sc_hd__a21o_4
X_46774_ _82961_/Q _46774_/Y sky130_fd_sc_hd__inv_2
X_77594_ _77559_/B _77576_/B _77576_/A _77594_/X sky130_fd_sc_hd__a21bo_4
X_43986_ _43986_/A _43986_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_994_0_CLK clkbuf_9_497_0_CLK/X _85601_/CLK sky130_fd_sc_hd__clkbuf_1
X_48513_ _83579_/Q _48514_/A sky130_fd_sc_hd__inv_2
X_79333_ _79332_/X _79333_/Y sky130_fd_sc_hd__inv_2
X_45725_ _45722_/X _45724_/Y _45678_/X _45725_/X sky130_fd_sc_hd__a21o_4
X_76545_ _76519_/X _76544_/Y _76511_/B _76545_/Y sky130_fd_sc_hd__o21ai_4
X_42937_ _42916_/X _42917_/X _41762_/X _67927_/B _42934_/X _42937_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49493_ _49493_/A _49493_/X sky130_fd_sc_hd__buf_2
X_61771_ _61711_/X _61839_/A sky130_fd_sc_hd__buf_2
X_73757_ _73733_/A _66022_/B _73757_/X sky130_fd_sc_hd__and2_4
X_70969_ _70969_/A _70947_/B _70969_/C _70969_/Y sky130_fd_sc_hd__nand3_4
X_63510_ _58551_/A _63497_/X _61483_/A _63498_/X _63510_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_9_485_0_CLK clkbuf_8_242_0_CLK/X clkbuf_9_485_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_48444_ _48444_/A _74403_/B sky130_fd_sc_hd__inv_2
X_60722_ _60722_/A _63672_/C _60711_/A _60722_/Y sky130_fd_sc_hd__nand3_4
X_72708_ _73078_/A _72943_/A sky130_fd_sc_hd__buf_2
X_79264_ _84793_/Q _66490_/C _79264_/Y sky130_fd_sc_hd__nand2_4
X_45656_ _63196_/B _61528_/A sky130_fd_sc_hd__buf_2
X_64490_ _64490_/A _64490_/B _79629_/B _64490_/Y sky130_fd_sc_hd__nor3_4
X_76476_ _76453_/Y _76455_/A _76451_/Y _76477_/A sky130_fd_sc_hd__o21a_4
X_42868_ _41570_/X _42866_/X _67079_/B _42867_/X _87678_/D sky130_fd_sc_hd__a2bb2o_4
X_73688_ _73685_/X _73687_/X _73612_/X _73688_/X sky130_fd_sc_hd__a21o_4
Xclkbuf_10_379_0_CLK clkbuf_9_189_0_CLK/X _83721_/CLK sky130_fd_sc_hd__clkbuf_1
X_78215_ _78209_/A _78208_/X _78220_/A _78215_/Y sky130_fd_sc_hd__a21boi_4
X_44607_ _44606_/Y _87037_/D sky130_fd_sc_hd__inv_2
X_75427_ _75423_/Y _75427_/B _75427_/C _75427_/X sky130_fd_sc_hd__or3_4
X_63441_ _63463_/A _64283_/C _63463_/C _63441_/X sky130_fd_sc_hd__and3_4
X_41819_ _41802_/X _41803_/X _40432_/X _66845_/B _41792_/X _41819_/Y
+ sky130_fd_sc_hd__o32ai_4
X_48375_ _48372_/X _82368_/Q _48374_/Y _74371_/A sky130_fd_sc_hd__o21ai_4
X_72639_ _72633_/X _72643_/B _56564_/B _72639_/Y sky130_fd_sc_hd__nand3_4
X_60653_ _60652_/X _63471_/A sky130_fd_sc_hd__buf_2
X_79195_ _79207_/B _79195_/Y sky130_fd_sc_hd__inv_2
X_45587_ _45583_/X _45586_/X _45523_/X _45587_/X sky130_fd_sc_hd__a21o_4
X_42799_ _42795_/X _42796_/X _41387_/X _67793_/B _42781_/X _42799_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47326_ _86646_/Q _47286_/X _47325_/Y _47326_/Y sky130_fd_sc_hd__o21ai_4
X_66160_ _57773_/X _84976_/Q _64579_/X _66159_/X _66160_/X sky130_fd_sc_hd__a211o_4
X_78146_ _78129_/X _78143_/A _78146_/X sky130_fd_sc_hd__and2_4
X_44538_ _44529_/X _44530_/X _40806_/A _44537_/Y _44533_/X _44538_/Y
+ sky130_fd_sc_hd__o32ai_4
X_63372_ _63372_/A _63372_/X sky130_fd_sc_hd__buf_2
X_75358_ _75358_/A _75357_/Y _75358_/X sky130_fd_sc_hd__xor2_4
X_60584_ _60555_/Y _60493_/X _60584_/Y sky130_fd_sc_hd__nand2_4
X_65111_ _65107_/X _65111_/B _65110_/X _65111_/Y sky130_fd_sc_hd__nand3_4
X_62323_ _62515_/A _62323_/X sky130_fd_sc_hd__buf_2
X_74309_ _70292_/C _74301_/X _74308_/Y _74309_/X sky130_fd_sc_hd__a21bo_4
X_47257_ _47246_/X _47228_/B _47234_/X _52942_/D _47257_/X sky130_fd_sc_hd__and4_4
X_66091_ _84157_/Q _66092_/C sky130_fd_sc_hd__inv_2
Xclkbuf_10_302_0_CLK clkbuf_9_151_0_CLK/X _84355_/CLK sky130_fd_sc_hd__clkbuf_1
X_78077_ _84582_/Q _78077_/B _81886_/D sky130_fd_sc_hd__xor2_4
X_44469_ _41165_/A _44464_/X _87093_/Q _44466_/X _87093_/D sky130_fd_sc_hd__a2bb2o_4
X_75289_ _75288_/A _80945_/D _75289_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_932_0_CLK clkbuf_9_466_0_CLK/X _87588_/CLK sky130_fd_sc_hd__clkbuf_1
X_46208_ _46187_/A _46215_/B sky130_fd_sc_hd__buf_2
X_65042_ _65039_/X _64937_/B _65041_/X _65042_/Y sky130_fd_sc_hd__nand3_4
X_77028_ _82086_/Q _77028_/B _77028_/X sky130_fd_sc_hd__xor2_4
X_62254_ _62181_/A _62181_/B _62254_/C _62254_/Y sky130_fd_sc_hd__nor3_4
X_47188_ _82373_/Q _47189_/A sky130_fd_sc_hd__inv_2
X_61205_ _61205_/A _61205_/B _60631_/D _61075_/X _64274_/A sky130_fd_sc_hd__and4_4
Xclkbuf_9_423_0_CLK clkbuf_9_423_0_CLK/A clkbuf_9_423_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_46139_ _46138_/Y _46139_/Y sky130_fd_sc_hd__inv_2
X_69850_ _68360_/X _42600_/Y _69850_/Y sky130_fd_sc_hd__nor2_4
X_62185_ _61694_/B _62185_/B _59649_/A _59761_/A _62188_/C sky130_fd_sc_hd__nand4_4
X_68801_ _68801_/A _68802_/B sky130_fd_sc_hd__inv_2
Xclkbuf_10_317_0_CLK clkbuf_9_158_0_CLK/X _85484_/CLK sky130_fd_sc_hd__clkbuf_1
X_61136_ _61135_/X _61238_/B sky130_fd_sc_hd__inv_2
X_69781_ _87555_/Q _69751_/X _69779_/X _69780_/Y _69781_/X sky130_fd_sc_hd__a211o_4
X_66993_ _84088_/Q _66971_/X _66992_/X _66993_/X sky130_fd_sc_hd__a21bo_4
X_78979_ _78979_/A _78979_/B _78979_/X sky130_fd_sc_hd__or2_4
Xclkbuf_10_947_0_CLK clkbuf_9_473_0_CLK/X _87826_/CLK sky130_fd_sc_hd__clkbuf_1
X_68732_ _68366_/X _68732_/B _68732_/Y sky130_fd_sc_hd__nor2_4
X_65944_ _65942_/Y _65915_/X _65943_/X _65944_/X sky130_fd_sc_hd__a21o_4
X_61067_ _60631_/D _61205_/B _61112_/A sky130_fd_sc_hd__and2_4
X_81990_ _81990_/CLK _82022_/Q _77023_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_438_0_CLK clkbuf_9_438_0_CLK/A clkbuf_9_438_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_60018_ _62623_/A _62556_/A sky130_fd_sc_hd__buf_2
X_49829_ _58012_/B _49825_/X _49828_/Y _49829_/Y sky130_fd_sc_hd__o21ai_4
X_80941_ _80813_/CLK _80985_/Q _80941_/Q sky130_fd_sc_hd__dfxtp_4
X_68663_ _68516_/X _68647_/Y _68649_/X _68662_/Y _68663_/X sky130_fd_sc_hd__a211o_4
X_65875_ _65685_/X _86179_/Q _65701_/X _65874_/X _65875_/X sky130_fd_sc_hd__a211o_4
X_67614_ _87975_/Q _67591_/X _67524_/X _67613_/X _67614_/X sky130_fd_sc_hd__a211o_4
X_52840_ _52757_/A _52853_/A sky130_fd_sc_hd__buf_2
X_64826_ _64826_/A _64826_/B _64826_/X sky130_fd_sc_hd__and2_4
X_83660_ _83660_/CLK _70927_/Y _46886_/A sky130_fd_sc_hd__dfxtp_4
X_80872_ _80746_/CLK _75628_/B _80872_/Q sky130_fd_sc_hd__dfxtp_4
X_68594_ _68590_/X _68593_/X _68442_/X _68597_/A sky130_fd_sc_hd__a21o_4
X_82611_ _82610_/CLK _78965_/B _82611_/Q sky130_fd_sc_hd__dfxtp_4
X_67545_ _67497_/A _87722_/Q _67545_/X sky130_fd_sc_hd__and2_4
X_52771_ _52775_/A _52775_/B _52775_/C _52771_/D _52771_/X sky130_fd_sc_hd__and4_4
X_64757_ _64754_/X _64756_/X _64729_/X _64757_/X sky130_fd_sc_hd__a21o_4
X_83591_ _83589_/CLK _71148_/Y _48379_/A sky130_fd_sc_hd__dfxtp_4
X_61969_ _58338_/A _61969_/X sky130_fd_sc_hd__buf_2
X_54510_ _54506_/Y _54502_/X _54509_/X _54510_/Y sky130_fd_sc_hd__a21oi_4
X_85330_ _83550_/CLK _85330_/D _85330_/Q sky130_fd_sc_hd__dfxtp_4
X_51722_ _51709_/X _51721_/X _51715_/C _53244_/D _51722_/X sky130_fd_sc_hd__and4_4
X_63708_ _58370_/A _63416_/A _63443_/A _63699_/D _63708_/Y sky130_fd_sc_hd__nand4_4
X_82542_ _82553_/CLK _83862_/Q _82542_/Q sky130_fd_sc_hd__dfxtp_4
X_55490_ _82994_/Q _44063_/X _44097_/X _55489_/Y _55490_/X sky130_fd_sc_hd__a211o_4
X_67476_ _67120_/X _67476_/X sky130_fd_sc_hd__buf_2
X_64688_ _84230_/Q _64688_/Y sky130_fd_sc_hd__inv_2
X_69215_ _81404_/D _69161_/X _69214_/X _83940_/D sky130_fd_sc_hd__a21bo_4
X_54441_ _54438_/Y _54422_/X _54440_/X _85442_/D sky130_fd_sc_hd__a21oi_4
X_66427_ _66366_/X _64926_/Y _66426_/Y _66427_/Y sky130_fd_sc_hd__o21ai_4
X_85261_ _85257_/CLK _56247_/Y _56246_/C sky130_fd_sc_hd__dfxtp_4
X_51653_ _51671_/A _53179_/B _51653_/Y sky130_fd_sc_hd__nand2_4
X_63639_ _64473_/A _60732_/C _60739_/X _58498_/A _60704_/Y _63639_/Y
+ sky130_fd_sc_hd__o32ai_4
X_82473_ _82671_/CLK _82473_/D _78303_/B sky130_fd_sc_hd__dfxtp_4
X_87000_ _82538_/CLK _87000_/D _44688_/A sky130_fd_sc_hd__dfxtp_4
X_84212_ _84210_/CLK _84212_/D _84212_/Q sky130_fd_sc_hd__dfxtp_4
X_50604_ _86169_/Q _50594_/X _50603_/Y _50604_/Y sky130_fd_sc_hd__o21ai_4
X_57160_ _57158_/Y _57159_/Y _57105_/Y _57160_/Y sky130_fd_sc_hd__o21ai_4
X_81424_ _81749_/CLK _81456_/Q _76036_/C sky130_fd_sc_hd__dfxtp_4
X_69146_ _69146_/A _69146_/X sky130_fd_sc_hd__buf_2
X_54372_ _54317_/A _54395_/C sky130_fd_sc_hd__buf_2
X_66358_ _66294_/X _66355_/Y _66357_/Y _66358_/Y sky130_fd_sc_hd__o21ai_4
X_85192_ _85192_/CLK _85192_/D _56442_/C sky130_fd_sc_hd__dfxtp_4
X_51584_ _51584_/A _51639_/A sky130_fd_sc_hd__buf_2
X_56111_ _56082_/X _56109_/X _56110_/Y _56111_/Y sky130_fd_sc_hd__o21ai_4
X_53323_ _53319_/Y _53301_/X _53322_/X _85655_/D sky130_fd_sc_hd__a21oi_4
X_65309_ _64772_/A _65309_/X sky130_fd_sc_hd__buf_2
X_84143_ _84231_/CLK _84143_/D _84143_/Q sky130_fd_sc_hd__dfxtp_4
X_50535_ _50541_/A _48851_/B _50535_/Y sky130_fd_sc_hd__nand2_4
X_81355_ _81322_/CLK _81355_/D _81355_/Q sky130_fd_sc_hd__dfxtp_4
X_57091_ _73227_/A _73198_/B sky130_fd_sc_hd__buf_2
X_69077_ _87990_/Q _69007_/X _69051_/X _69076_/X _69077_/X sky130_fd_sc_hd__a211o_4
X_66289_ _57761_/X _84967_/Q _65309_/X _66288_/X _66289_/X sky130_fd_sc_hd__a211o_4
X_80306_ _80319_/B _80306_/Y sky130_fd_sc_hd__inv_2
X_56042_ _56029_/X _56040_/X _56041_/Y _56042_/Y sky130_fd_sc_hd__o21ai_4
X_68028_ _68028_/A _87702_/Q _68028_/X sky130_fd_sc_hd__and2_4
X_53254_ _53252_/Y _53242_/X _53253_/X _85668_/D sky130_fd_sc_hd__a21oi_4
X_84074_ _84074_/CLK _84074_/D _84074_/Q sky130_fd_sc_hd__dfxtp_4
X_50466_ _50465_/X _50466_/B _50466_/Y sky130_fd_sc_hd__nand2_4
X_81286_ _81603_/CLK _76974_/X _81286_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_5_17_0_CLK clkbuf_4_8_1_CLK/X clkbuf_6_35_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_52205_ _52202_/Y _52203_/X _52204_/X _85869_/D sky130_fd_sc_hd__a21oi_4
X_83025_ _83025_/CLK _83025_/D _83025_/Q sky130_fd_sc_hd__dfxtp_4
X_87902_ _87644_/CLK _87902_/D _87902_/Q sky130_fd_sc_hd__dfxtp_4
X_80237_ _80244_/B _80236_/Y _80237_/X sky130_fd_sc_hd__xor2_4
X_53185_ _53181_/A _53181_/B _53169_/X _53185_/D _53185_/X sky130_fd_sc_hd__and4_4
X_50397_ _50394_/Y _50395_/X _50396_/X _86209_/D sky130_fd_sc_hd__a21oi_4
X_59801_ _59801_/A _70009_/A sky130_fd_sc_hd__buf_2
X_52136_ _52133_/Y _52108_/X _52135_/X _52136_/Y sky130_fd_sc_hd__a21oi_4
X_87833_ _87834_/CLK _87833_/D _74164_/A sky130_fd_sc_hd__dfxtp_4
X_80168_ _80164_/Y _80167_/Y _80178_/B sky130_fd_sc_hd__xor2_4
X_57993_ _72417_/A _57993_/X sky130_fd_sc_hd__buf_2
X_69979_ _69574_/Y _69916_/X _69938_/X _69978_/Y _69979_/X sky130_fd_sc_hd__a211o_4
X_59732_ _59649_/A _59754_/C sky130_fd_sc_hd__buf_2
X_52067_ _52431_/A _52083_/A sky130_fd_sc_hd__buf_2
X_56944_ _44214_/X _56571_/X _45409_/A _56943_/X _85120_/D sky130_fd_sc_hd__a2bb2o_4
X_87764_ _87766_/CLK _42698_/X _69553_/B sky130_fd_sc_hd__dfxtp_4
X_72990_ _72988_/X _85593_/Q _44272_/X _72989_/X _72990_/X sky130_fd_sc_hd__a211o_4
X_84976_ _86576_/CLK _57577_/Y _84976_/Q sky130_fd_sc_hd__dfxtp_4
X_80099_ _84938_/Q _84186_/Q _80099_/Y sky130_fd_sc_hd__nand2_4
X_51018_ _51018_/A _51029_/B _51029_/C _52709_/D _51018_/X sky130_fd_sc_hd__and4_4
X_86715_ _86711_/CLK _86715_/D _58649_/A sky130_fd_sc_hd__dfxtp_4
X_71941_ _55681_/A _71939_/X _71940_/Y _71941_/Y sky130_fd_sc_hd__o21ai_4
X_83927_ _81473_/CLK _83927_/D _81391_/D sky130_fd_sc_hd__dfxtp_4
X_59663_ _59681_/A _59754_/D sky130_fd_sc_hd__inv_2
X_56875_ _56636_/X _56865_/Y _56874_/X _56875_/X sky130_fd_sc_hd__a21o_4
X_87695_ _87950_/CLK _42833_/X _87695_/Q sky130_fd_sc_hd__dfxtp_4
X_58614_ _86717_/Q _58614_/B _58614_/Y sky130_fd_sc_hd__nor2_4
X_43840_ _43840_/A _87239_/D sky130_fd_sc_hd__inv_2
X_55826_ _55826_/A _55826_/B _55826_/X sky130_fd_sc_hd__and2_4
X_86646_ _86008_/CLK _86646_/D _86646_/Q sky130_fd_sc_hd__dfxtp_4
X_74660_ _74642_/X _45654_/A _74660_/Y sky130_fd_sc_hd__nand2_4
X_71872_ _71783_/A _71883_/B sky130_fd_sc_hd__buf_2
X_59594_ _59593_/X _59622_/A sky130_fd_sc_hd__buf_2
X_83858_ _82536_/CLK _83858_/D _82538_/D sky130_fd_sc_hd__dfxtp_4
X_73611_ _73609_/X _85631_/Q _73472_/X _73610_/X _73611_/X sky130_fd_sc_hd__a211o_4
X_70823_ _51222_/B _70802_/A _70822_/Y _83691_/D sky130_fd_sc_hd__o21ai_4
X_58545_ _58538_/X _83359_/Q _58544_/Y _58545_/X sky130_fd_sc_hd__o21a_4
X_82809_ _82743_/CLK _82841_/Q _82809_/Q sky130_fd_sc_hd__dfxtp_4
X_43771_ _43606_/A _43802_/A sky130_fd_sc_hd__buf_2
X_55757_ _85255_/Q _55190_/X _44045_/X _55756_/X _55757_/X sky130_fd_sc_hd__a211o_4
X_74591_ _56863_/X _74591_/X sky130_fd_sc_hd__buf_2
X_86577_ _85630_/CLK _86577_/D _66143_/B sky130_fd_sc_hd__dfxtp_4
X_52969_ _52979_/A _52969_/B _52969_/Y sky130_fd_sc_hd__nand2_4
X_40983_ _40982_/X _40941_/X _69265_/B _40942_/X _88298_/D sky130_fd_sc_hd__a2bb2o_4
X_83789_ _81259_/CLK _70345_/X _74769_/A sky130_fd_sc_hd__dfxtp_4
X_45510_ _45510_/A _45590_/B _45510_/X sky130_fd_sc_hd__and2_4
X_76330_ _76330_/A _76330_/Y sky130_fd_sc_hd__inv_2
X_88316_ _87063_/CLK _40891_/X _88316_/Q sky130_fd_sc_hd__dfxtp_4
X_54708_ _54706_/Y _54694_/X _54707_/X _54708_/Y sky130_fd_sc_hd__a21oi_4
X_42722_ _42429_/A _42723_/A sky130_fd_sc_hd__buf_2
X_73542_ _73542_/A _73542_/B _73543_/B sky130_fd_sc_hd__nand2_4
X_85528_ _85529_/CLK _85528_/D _85528_/Q sky130_fd_sc_hd__dfxtp_4
X_46490_ _52526_/B _50832_/B sky130_fd_sc_hd__buf_2
X_70754_ _53131_/B _70740_/A _70753_/Y _83707_/D sky130_fd_sc_hd__o21ai_4
X_58476_ _83415_/Q _58476_/Y sky130_fd_sc_hd__inv_2
X_55688_ _56169_/A _55688_/X sky130_fd_sc_hd__buf_2
X_45441_ _45438_/Y _45439_/X _45390_/X _45440_/Y _45441_/X sky130_fd_sc_hd__a211o_4
X_57427_ _57427_/A _57445_/B _56750_/Y _57427_/Y sky130_fd_sc_hd__nand3_4
X_76261_ _81642_/Q _76260_/X _76261_/X sky130_fd_sc_hd__or2_4
X_88247_ _88247_/CLK _41269_/X _69048_/B sky130_fd_sc_hd__dfxtp_4
X_42653_ _42634_/A _42653_/X sky130_fd_sc_hd__buf_2
X_54639_ _54625_/A _54645_/B _54618_/X _47264_/A _54639_/X sky130_fd_sc_hd__and4_4
X_73473_ _73426_/A _86469_/Q _73473_/X sky130_fd_sc_hd__and2_4
X_85459_ _85459_/CLK _54348_/Y _85459_/Q sky130_fd_sc_hd__dfxtp_4
X_70685_ _70669_/A _70692_/C sky130_fd_sc_hd__buf_2
X_78000_ _78000_/A _78000_/Y sky130_fd_sc_hd__inv_2
X_75212_ _80683_/Q _80983_/Q _75201_/Y _75212_/Y sky130_fd_sc_hd__a21boi_4
X_41604_ _41604_/A _82309_/Q _41604_/X sky130_fd_sc_hd__or2_4
X_48160_ _48801_/A _50391_/A _48160_/X sky130_fd_sc_hd__and2_4
X_72424_ _72352_/X _85960_/Q _72423_/X _72424_/Y sky130_fd_sc_hd__o21ai_4
X_57358_ _57358_/A _57068_/X _57358_/X sky130_fd_sc_hd__xor2_4
X_45372_ _45362_/X _45366_/Y _45371_/Y _45372_/Y sky130_fd_sc_hd__a21oi_4
X_76192_ _76188_/X _76193_/C _76193_/A _76192_/X sky130_fd_sc_hd__a21o_4
X_88178_ _82896_/CLK _88178_/D _67365_/B sky130_fd_sc_hd__dfxtp_4
X_42584_ _42568_/X _42569_/X _40845_/X _42583_/Y _42571_/X _42584_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47111_ _47111_/A _54553_/D sky130_fd_sc_hd__inv_2
X_56309_ _56309_/A _56298_/X _85241_/Q _56309_/Y sky130_fd_sc_hd__nand3_4
X_44323_ _41636_/X _40543_/X _87166_/Q _40544_/X _87166_/D sky130_fd_sc_hd__a2bb2o_4
X_75143_ _75143_/A _75127_/C _75143_/Y sky130_fd_sc_hd__nand2_4
X_87129_ _87436_/CLK _44398_/Y _87129_/Q sky130_fd_sc_hd__dfxtp_4
X_41535_ _41533_/X _82322_/Q _41534_/X _41535_/X sky130_fd_sc_hd__o21a_4
X_48091_ _57617_/B _50358_/B sky130_fd_sc_hd__buf_2
X_72355_ _72351_/Y _72354_/Y _72344_/X _72355_/X sky130_fd_sc_hd__a21o_4
X_57289_ _56842_/X _57289_/B _56848_/X _56849_/X _57290_/A sky130_fd_sc_hd__nor4_4
X_47042_ _53336_/B _51130_/B sky130_fd_sc_hd__buf_2
X_59028_ _58698_/A _59029_/A sky130_fd_sc_hd__buf_2
X_71306_ _71303_/A _71303_/B _71680_/C _71306_/Y sky130_fd_sc_hd__nand3_4
X_44254_ _58631_/A _57811_/A _72296_/A _44252_/X _44253_/X _44254_/X
+ sky130_fd_sc_hd__a41o_4
X_75074_ _75072_/Y _75074_/B _75074_/X sky130_fd_sc_hd__and2_4
X_79951_ _79957_/A _79956_/A sky130_fd_sc_hd__inv_2
X_41466_ _41465_/X _41455_/X _88210_/Q _41457_/X _41466_/X sky130_fd_sc_hd__a2bb2o_4
X_72286_ _83267_/Q _72286_/Y sky130_fd_sc_hd__inv_2
X_43205_ _40935_/X _43180_/X _87539_/Q _43185_/X _43205_/X sky130_fd_sc_hd__a2bb2o_4
X_74025_ _74025_/A _74025_/B _74026_/B sky130_fd_sc_hd__nand2_4
X_78902_ _82637_/Q _78902_/Y sky130_fd_sc_hd__inv_2
X_40417_ _40325_/X _82328_/Q _40416_/X _40417_/Y sky130_fd_sc_hd__o21ai_4
X_71237_ _71136_/A _70758_/C _70758_/B _70627_/A _71238_/B sky130_fd_sc_hd__nand4_4
X_44185_ _44171_/X _44173_/X _44177_/X _72461_/A _44184_/X _44185_/X
+ sky130_fd_sc_hd__a41o_4
X_79882_ _79882_/A _79881_/X _79890_/A sky130_fd_sc_hd__nand2_4
X_41397_ _41397_/A _41397_/X sky130_fd_sc_hd__buf_2
Xclkbuf_7_100_0_CLK clkbuf_6_50_0_CLK/X clkbuf_8_201_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_43136_ _43129_/X _43130_/X _40806_/X _43135_/Y _43127_/X _43136_/Y
+ sky130_fd_sc_hd__o32ai_4
X_78833_ _82837_/Q _78833_/B _78833_/Y sky130_fd_sc_hd__xnor2_4
X_40348_ _46450_/A _74458_/A sky130_fd_sc_hd__buf_2
X_71168_ _71168_/A _71173_/B _74531_/B _71178_/D _71168_/Y sky130_fd_sc_hd__nand4_4
X_48993_ _48964_/A _48992_/X _48993_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_70_0_CLK clkbuf_9_35_0_CLK/X _80672_/CLK sky130_fd_sc_hd__clkbuf_1
X_70119_ _83525_/Q _83173_/Q _83500_/Q _83148_/Q _70119_/Y sky130_fd_sc_hd__a22oi_4
X_47944_ _46301_/X _82359_/Q _47943_/X _51988_/A sky130_fd_sc_hd__o21ai_4
X_43067_ _43066_/Y _87589_/D sky130_fd_sc_hd__inv_2
X_78764_ _78764_/A _78759_/X _78764_/Y sky130_fd_sc_hd__nand2_4
X_63990_ _61510_/X _64052_/B _64003_/C _64052_/D _63990_/Y sky130_fd_sc_hd__nand4_4
X_71099_ _71088_/A _71076_/B _71099_/C _71099_/Y sky130_fd_sc_hd__nand3_4
X_75976_ _75976_/A _75976_/B _75977_/B sky130_fd_sc_hd__nor2_4
X_42018_ _42013_/X _42006_/X _40839_/X _73124_/A _42007_/X _42018_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77715_ _77715_/A _77715_/B _77716_/B sky130_fd_sc_hd__xnor2_4
X_74927_ _80941_/Q _74927_/B _74927_/X sky130_fd_sc_hd__xor2_4
X_62941_ _62934_/Y _62886_/X _62935_/Y _62938_/Y _62940_/X _62941_/X
+ sky130_fd_sc_hd__a41o_4
Xclkbuf_7_115_0_CLK clkbuf_6_57_0_CLK/X clkbuf_8_231_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_47875_ _51340_/A _47918_/A sky130_fd_sc_hd__buf_2
X_78695_ _78682_/A _78682_/B _78680_/Y _78695_/X sky130_fd_sc_hd__o21a_4
X_49614_ _49614_/A _49614_/X sky130_fd_sc_hd__buf_2
X_46826_ _46817_/A _51003_/B _46826_/Y sky130_fd_sc_hd__nand2_4
X_65660_ _65660_/A _65660_/X sky130_fd_sc_hd__buf_2
X_77646_ _77643_/B _77643_/A _77648_/C sky130_fd_sc_hd__nand2_4
X_62872_ _62867_/X _62831_/X _62869_/Y _62870_/Y _62871_/X _62872_/X
+ sky130_fd_sc_hd__a41o_4
X_74858_ _81123_/D _80835_/Q _74858_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_85_0_CLK clkbuf_9_42_0_CLK/X _83246_/CLK sky130_fd_sc_hd__clkbuf_1
X_64611_ _64611_/A _85824_/Q _64611_/X sky130_fd_sc_hd__and2_4
X_49545_ _49540_/Y _49541_/X _49544_/X _49545_/Y sky130_fd_sc_hd__a21oi_4
X_61823_ _61823_/A _61823_/B _59501_/X _61788_/X _61823_/X sky130_fd_sc_hd__and4_4
X_73809_ _73806_/X _73808_/X _73738_/X _73812_/A sky130_fd_sc_hd__a21o_4
X_46757_ _83674_/Q _52658_/B sky130_fd_sc_hd__inv_2
X_65591_ _65484_/X _86198_/Q _65534_/X _65590_/X _65591_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_8_231_0_CLK clkbuf_8_231_0_CLK/A clkbuf_8_231_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_77577_ _77560_/Y _77564_/B _77559_/B _77577_/Y sky130_fd_sc_hd__o21ai_4
X_43969_ _43969_/A _43969_/B _43970_/A sky130_fd_sc_hd__and2_4
X_74789_ _71735_/A _70630_/B _74789_/C _71010_/X _74789_/X sky130_fd_sc_hd__and4_4
X_67330_ _68461_/A _67806_/A sky130_fd_sc_hd__buf_2
X_79316_ _79313_/Y _79296_/Y _79315_/X _79316_/Y sky130_fd_sc_hd__o21ai_4
X_45708_ _45704_/X _45707_/Y _45678_/X _45708_/X sky130_fd_sc_hd__a21o_4
X_76528_ _76516_/Y _76509_/X _76511_/B _76529_/B sky130_fd_sc_hd__a21boi_4
X_64542_ _64542_/A _64542_/Y sky130_fd_sc_hd__inv_2
X_49476_ _49481_/A _50998_/B _49476_/Y sky130_fd_sc_hd__nand2_4
X_61754_ _61770_/A _61770_/B _63384_/B _61770_/D _61754_/X sky130_fd_sc_hd__and4_4
X_46688_ _82970_/Q _46688_/Y sky130_fd_sc_hd__inv_2
X_48427_ _48426_/Y _48449_/B _48427_/Y sky130_fd_sc_hd__nand2_4
X_60705_ _60700_/A _60612_/B _84582_/Q _60705_/Y sky130_fd_sc_hd__nor3_4
X_67261_ _67144_/A _67308_/A sky130_fd_sc_hd__buf_2
X_79247_ _79229_/Y _79248_/C _79246_/Y _79247_/X sky130_fd_sc_hd__a21o_4
X_45639_ _45636_/X _45638_/Y _45561_/X _45639_/Y sky130_fd_sc_hd__a21oi_4
X_64473_ _64473_/A _64454_/B _64473_/Y sky130_fd_sc_hd__nor2_4
X_76459_ _76459_/A _81526_/D _76459_/Y sky130_fd_sc_hd__nand2_4
X_61685_ _61685_/A _61653_/X _61654_/X _61639_/X _61685_/Y sky130_fd_sc_hd__nand4_4
X_69000_ _87577_/Q _66538_/X _66540_/X _68999_/X _69000_/X sky130_fd_sc_hd__a211o_4
X_66212_ _57947_/A _85612_/Q _65301_/X _66211_/X _66212_/X sky130_fd_sc_hd__a211o_4
X_63424_ _63448_/A _63424_/B _63410_/C _63410_/D _63424_/X sky130_fd_sc_hd__and4_4
Xclkbuf_8_246_0_CLK clkbuf_8_247_0_CLK/A clkbuf_9_493_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_60636_ _61276_/B _60636_/B _59657_/A _60407_/C _60637_/A sky130_fd_sc_hd__and4_4
X_48358_ _48357_/Y _48358_/X sky130_fd_sc_hd__buf_2
X_67192_ _67189_/X _67191_/X _67147_/X _67197_/A sky130_fd_sc_hd__a21o_4
X_79178_ _79164_/Y _79523_/B _79178_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_241_0_CLK clkbuf_9_120_0_CLK/X _84562_/CLK sky130_fd_sc_hd__clkbuf_1
X_47309_ _81816_/Q _47310_/A sky130_fd_sc_hd__inv_2
Xclkbuf_10_871_0_CLK clkbuf_9_435_0_CLK/X _86736_/CLK sky130_fd_sc_hd__clkbuf_1
X_66143_ _65934_/X _66143_/B _66143_/X sky130_fd_sc_hd__and2_4
X_78129_ _82570_/Q _82858_/D _78129_/X sky130_fd_sc_hd__xor2_4
X_63355_ _63355_/A _60642_/A _60638_/Y _60642_/C _63355_/Y sky130_fd_sc_hd__nand4_4
X_48289_ _48264_/X _52036_/B _48289_/Y sky130_fd_sc_hd__nand2_4
X_60567_ _60566_/X _60567_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_23_0_CLK clkbuf_9_11_0_CLK/X _85190_/CLK sky130_fd_sc_hd__clkbuf_1
X_50320_ _50638_/A _50572_/A sky130_fd_sc_hd__buf_2
X_62306_ _62196_/X _61831_/X _62305_/X _62306_/X sky130_fd_sc_hd__a21o_4
X_81140_ _81197_/CLK _81140_/D _40659_/A sky130_fd_sc_hd__dfxtp_4
X_66074_ _57770_/A _73833_/B _66074_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_362_0_CLK clkbuf_9_363_0_CLK/A clkbuf_9_362_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_63286_ _63283_/X _63284_/X _63285_/Y _63286_/Y sky130_fd_sc_hd__a21oi_4
X_60498_ _60435_/A _60493_/X _60495_/X _60572_/C _60497_/Y _60498_/Y
+ sky130_fd_sc_hd__a41oi_4
X_65025_ _64948_/A _65025_/B _65025_/X sky130_fd_sc_hd__and2_4
X_69902_ _69902_/A _69902_/B _69902_/Y sky130_fd_sc_hd__nand2_4
X_50251_ _50222_/X _50251_/X sky130_fd_sc_hd__buf_2
X_62237_ _62237_/A _62237_/X sky130_fd_sc_hd__buf_2
X_81071_ _80817_/CLK _75839_/A _75254_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_256_0_CLK clkbuf_9_128_0_CLK/X _84344_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_886_0_CLK clkbuf_9_443_0_CLK/X _86030_/CLK sky130_fd_sc_hd__clkbuf_1
X_80022_ _80013_/Y _80008_/X _80021_/X _80023_/B sky130_fd_sc_hd__a21boi_4
X_69833_ _69747_/A _69833_/X sky130_fd_sc_hd__buf_2
X_50182_ _65285_/B _50162_/X _50181_/Y _50182_/Y sky130_fd_sc_hd__o21ai_4
X_62168_ _62165_/Y _62166_/X _62167_/Y _84428_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_38_0_CLK clkbuf_9_19_0_CLK/X _85083_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_9_377_0_CLK clkbuf_8_188_0_CLK/X clkbuf_9_377_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_61119_ _64546_/A _61125_/A sky130_fd_sc_hd__inv_2
X_84830_ _84714_/CLK _58516_/Y _84830_/Q sky130_fd_sc_hd__dfxtp_4
X_69764_ _69086_/A _73149_/A _69764_/X sky130_fd_sc_hd__and2_4
X_54990_ _85339_/Q _54967_/X _54989_/Y _54990_/Y sky130_fd_sc_hd__o21ai_4
X_66976_ _87362_/Q _66878_/X _66879_/X _66975_/X _66976_/X sky130_fd_sc_hd__a211o_4
X_62099_ _59794_/X _62088_/B _62096_/Y _62099_/D _62099_/Y sky130_fd_sc_hd__nand4_4
X_68715_ _69958_/A _68715_/X sky130_fd_sc_hd__buf_2
X_53941_ _54295_/A _53942_/A sky130_fd_sc_hd__buf_2
X_65927_ _65923_/X _65741_/B _65927_/C _65927_/Y sky130_fd_sc_hd__nand3_4
X_84761_ _84766_/CLK _84761_/D _84761_/Q sky130_fd_sc_hd__dfxtp_4
X_81973_ _82116_/CLK _83901_/Q _81973_/Q sky130_fd_sc_hd__dfxtp_4
X_69695_ _81976_/D _69632_/X _69694_/X _83904_/D sky130_fd_sc_hd__a21bo_4
X_86500_ _86500_/CLK _48692_/Y _86500_/Q sky130_fd_sc_hd__dfxtp_4
X_83712_ _86303_/CLK _83712_/D _47535_/A sky130_fd_sc_hd__dfxtp_4
X_56660_ _56660_/A _56659_/Y _83333_/Q _56661_/C sky130_fd_sc_hd__nand3_4
X_80924_ _80928_/CLK _84100_/Q _75807_/A sky130_fd_sc_hd__dfxtp_4
X_68646_ _44697_/A _68570_/X _68571_/X _68645_/X _68646_/X sky130_fd_sc_hd__a211o_4
X_87480_ _87993_/CLK _87480_/D _87480_/Q sky130_fd_sc_hd__dfxtp_4
X_53872_ _53871_/X _49064_/A _53872_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_300_0_CLK clkbuf_8_150_0_CLK/X clkbuf_9_300_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_65858_ _65845_/X _86180_/Q _65790_/X _65857_/X _65858_/X sky130_fd_sc_hd__a211o_4
X_84692_ _83227_/CLK _59835_/X _80400_/A sky130_fd_sc_hd__dfxtp_4
X_55611_ _55610_/X _55611_/X sky130_fd_sc_hd__buf_2
X_86431_ _85536_/CLK _86431_/D _64647_/B sky130_fd_sc_hd__dfxtp_4
X_52823_ _52843_/A _51130_/B _52823_/Y sky130_fd_sc_hd__nand2_4
X_64809_ _64809_/A _64809_/X sky130_fd_sc_hd__buf_2
X_83643_ _86422_/CLK _70977_/Y _46410_/A sky130_fd_sc_hd__dfxtp_4
X_56591_ _56587_/X _56589_/X _85148_/Q _56590_/X _85148_/D sky130_fd_sc_hd__a2bb2o_4
X_80855_ _80854_/CLK _80887_/Q _75003_/B sky130_fd_sc_hd__dfxtp_4
X_68577_ _68452_/A _87243_/Q _68577_/X sky130_fd_sc_hd__and2_4
X_65789_ _65516_/A _65789_/X sky130_fd_sc_hd__buf_2
X_58330_ _58408_/A _58364_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_824_0_CLK clkbuf_9_412_0_CLK/X _82879_/CLK sky130_fd_sc_hd__clkbuf_1
X_55542_ _55462_/X _45515_/Y _55542_/Y sky130_fd_sc_hd__nor2_4
X_67528_ _87467_/Q _67476_/X _67477_/X _67527_/X _67528_/X sky130_fd_sc_hd__a211o_4
X_86362_ _83049_/CLK _49578_/Y _86362_/Q sky130_fd_sc_hd__dfxtp_4
X_52754_ _52754_/A _52783_/A sky130_fd_sc_hd__buf_2
X_83574_ _86505_/CLK _83574_/D _48571_/A sky130_fd_sc_hd__dfxtp_4
X_80786_ _80754_/CLK _80786_/D _80786_/Q sky130_fd_sc_hd__dfxtp_4
X_88101_ _88097_/CLK _41934_/Y _73892_/A sky130_fd_sc_hd__dfxtp_4
X_85313_ _85138_/CLK _55991_/Y _55990_/C sky130_fd_sc_hd__dfxtp_4
X_51705_ _51695_/A _51715_/B _51695_/C _53230_/D _51705_/X sky130_fd_sc_hd__and4_4
Xclkbuf_9_315_0_CLK clkbuf_9_315_0_CLK/A clkbuf_9_315_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_58261_ _62027_/A _58261_/Y sky130_fd_sc_hd__inv_2
X_82525_ _82503_/CLK _82525_/D _78727_/A sky130_fd_sc_hd__dfxtp_4
X_55473_ _45617_/A _55468_/X _55458_/X _55472_/Y _55473_/X sky130_fd_sc_hd__a211o_4
X_67459_ _67222_/A _67460_/A sky130_fd_sc_hd__buf_2
X_86293_ _86611_/CLK _86293_/D _86293_/Q sky130_fd_sc_hd__dfxtp_4
X_52685_ _52657_/A _52706_/A sky130_fd_sc_hd__buf_2
X_57212_ _57212_/A _57212_/Y sky130_fd_sc_hd__inv_2
X_88032_ _88036_/CLK _42109_/Y _88032_/Q sky130_fd_sc_hd__dfxtp_4
X_54424_ _54420_/Y _54422_/X _54423_/X _54424_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_209_0_CLK clkbuf_9_104_0_CLK/X _84498_/CLK sky130_fd_sc_hd__clkbuf_1
X_85244_ _85244_/CLK _56302_/Y _85244_/Q sky130_fd_sc_hd__dfxtp_4
X_51636_ _51633_/Y _51613_/X _51635_/X _85974_/D sky130_fd_sc_hd__a21oi_4
X_58192_ _83375_/Q _58192_/Y sky130_fd_sc_hd__inv_2
X_70470_ _71706_/A _71366_/A _71424_/C _70470_/X sky130_fd_sc_hd__and3_4
X_82456_ _84177_/CLK _82456_/D _82456_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_839_0_CLK clkbuf_9_419_0_CLK/X _83783_/CLK sky130_fd_sc_hd__clkbuf_1
Xclkbuf_5_0_0_CLK clkbuf_4_0_1_CLK/X clkbuf_6_1_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_81407_ _83940_/CLK _83943_/Q _76766_/B sky130_fd_sc_hd__dfxtp_4
X_57143_ _56729_/X _57023_/X _57129_/Y _56816_/A _57270_/A _57143_/X
+ sky130_fd_sc_hd__a41o_4
X_69129_ _69128_/X _69129_/B _69129_/X sky130_fd_sc_hd__and2_4
X_54355_ _54355_/A _52663_/B _54355_/Y sky130_fd_sc_hd__nand2_4
X_85175_ _85270_/CLK _85175_/D _55896_/B sky130_fd_sc_hd__dfxtp_4
X_51567_ _51622_/A _51590_/A sky130_fd_sc_hd__buf_2
X_82387_ _85491_/CLK _82387_/D _82387_/Q sky130_fd_sc_hd__dfxtp_4
X_41320_ _41042_/X _81754_/Q _41319_/X _41320_/X sky130_fd_sc_hd__o21a_4
X_53306_ _85658_/Q _53295_/X _53305_/Y _53306_/Y sky130_fd_sc_hd__o21ai_4
X_72140_ _86623_/Q _72193_/B _72140_/Y sky130_fd_sc_hd__nor2_4
X_84126_ _82152_/CLK _66425_/X _84126_/Q sky130_fd_sc_hd__dfxtp_4
X_50518_ _86185_/Q _50506_/X _50517_/Y _50518_/Y sky130_fd_sc_hd__o21ai_4
X_57074_ _44290_/X _45891_/X _56275_/X _57223_/D _56914_/Y _57075_/A
+ sky130_fd_sc_hd__a41oi_4
X_81338_ _82053_/CLK _76518_/X _81714_/D sky130_fd_sc_hd__dfxtp_4
X_54286_ _54286_/A _54298_/B _54286_/C _54286_/D _54286_/X sky130_fd_sc_hd__and4_4
X_51498_ _51552_/A _51522_/C sky130_fd_sc_hd__buf_2
X_56025_ _56003_/B _56002_/A _56025_/X sky130_fd_sc_hd__xor2_4
X_41251_ _41181_/A _41251_/X sky130_fd_sc_hd__buf_2
X_53237_ _85671_/Q _53225_/X _53236_/Y _53237_/Y sky130_fd_sc_hd__o21ai_4
X_72071_ _72069_/Y _72059_/X _72070_/X _72071_/Y sky130_fd_sc_hd__a21oi_4
X_84057_ _81492_/CLK _67736_/X _84057_/Q sky130_fd_sc_hd__dfxtp_4
X_50449_ _50439_/X _48482_/B _50449_/Y sky130_fd_sc_hd__nand2_4
X_81269_ _81269_/CLK _81301_/Q _81269_/Q sky130_fd_sc_hd__dfxtp_4
X_71022_ _53148_/B _71013_/X _71021_/Y _83632_/D sky130_fd_sc_hd__o21ai_4
X_83008_ _83008_/CLK _83008_/D _45416_/A sky130_fd_sc_hd__dfxtp_4
X_41182_ _40989_/A _41182_/X sky130_fd_sc_hd__buf_2
X_53168_ _85684_/Q _53146_/X _53167_/Y _53168_/Y sky130_fd_sc_hd__o21ai_4
X_52119_ _52188_/A _52119_/B _52119_/Y sky130_fd_sc_hd__nand2_4
X_75830_ _75830_/A _75830_/B _75831_/A sky130_fd_sc_hd__xor2_4
X_87816_ _87820_/CLK _42572_/Y _87816_/Q sky130_fd_sc_hd__dfxtp_4
X_45990_ _45980_/X _45987_/X _40445_/X _86825_/Q _45982_/X _45991_/A
+ sky130_fd_sc_hd__o32ai_4
X_53099_ _53107_/A _53113_/B _53107_/C _53099_/D _53099_/X sky130_fd_sc_hd__and4_4
X_57976_ _57966_/X _85711_/Q _57878_/X _57976_/X sky130_fd_sc_hd__o21a_4
X_59715_ _57689_/A _60132_/A sky130_fd_sc_hd__buf_2
X_44941_ _44905_/X _61354_/B _44907_/X _44941_/Y sky130_fd_sc_hd__o21ai_4
X_56927_ _56927_/A _56774_/C _56927_/C _56927_/Y sky130_fd_sc_hd__nand3_4
X_75761_ _80919_/Q _75761_/Y sky130_fd_sc_hd__inv_2
X_87747_ _87749_/CLK _42730_/X _68768_/B sky130_fd_sc_hd__dfxtp_4
X_72973_ _72973_/A _72973_/B _72973_/Y sky130_fd_sc_hd__nor2_4
X_84959_ _84869_/CLK _84959_/D _84959_/Q sky130_fd_sc_hd__dfxtp_4
X_77500_ _77499_/X _77478_/X _77479_/X _77500_/Y sky130_fd_sc_hd__a21oi_4
X_74712_ _74711_/A _74712_/Y sky130_fd_sc_hd__inv_2
X_47660_ _72295_/A _47619_/X _47659_/Y _47660_/Y sky130_fd_sc_hd__o21ai_4
X_71924_ _71920_/Y _56727_/X _71923_/Y _83327_/D sky130_fd_sc_hd__a21o_4
X_59646_ _59664_/C _59824_/B sky130_fd_sc_hd__buf_2
X_78480_ _78466_/X _78478_/Y _78479_/Y _78480_/X sky130_fd_sc_hd__a21o_4
X_44872_ _80670_/Q _45193_/A sky130_fd_sc_hd__buf_2
X_56858_ _83334_/Q _57346_/C sky130_fd_sc_hd__buf_2
X_75692_ _75692_/A _75692_/B _75693_/B sky130_fd_sc_hd__xnor2_4
X_87678_ _82886_/CLK _87678_/D _67079_/B sky130_fd_sc_hd__dfxtp_4
X_46611_ _74509_/B _46620_/A sky130_fd_sc_hd__buf_2
X_77431_ _77426_/X _77431_/B _77427_/Y _77431_/Y sky130_fd_sc_hd__nand3_4
X_55809_ _45215_/A _55492_/X _44096_/X _55808_/X _55809_/X sky130_fd_sc_hd__a211o_4
X_43823_ _43166_/A _43854_/A sky130_fd_sc_hd__buf_2
X_74643_ _74642_/X _45495_/A _74643_/Y sky130_fd_sc_hd__nand2_4
X_86629_ _85990_/CLK _47496_/Y _58097_/A sky130_fd_sc_hd__dfxtp_4
X_47591_ _47574_/A _53135_/B _47591_/Y sky130_fd_sc_hd__nand2_4
X_71855_ _70543_/Y _71857_/B _71851_/X _71857_/D _71855_/Y sky130_fd_sc_hd__nor4_4
X_59577_ _59571_/B _59876_/B _59560_/A _43995_/A _59577_/X sky130_fd_sc_hd__and4_4
X_56789_ _56783_/X _57170_/A sky130_fd_sc_hd__buf_2
X_49330_ _49287_/A _50852_/B _49330_/Y sky130_fd_sc_hd__nand2_4
X_46542_ _46249_/A _46542_/X sky130_fd_sc_hd__buf_2
X_70806_ _74531_/C _70810_/C sky130_fd_sc_hd__buf_2
X_58528_ _58528_/A _58510_/X _58528_/Y sky130_fd_sc_hd__nor2_4
X_77362_ _77371_/A _77361_/Y _77362_/X sky130_fd_sc_hd__or2_4
X_43754_ _40939_/X _43752_/X _87282_/Q _43753_/X _87282_/D sky130_fd_sc_hd__a2bb2o_4
X_74574_ _45082_/A _74568_/X _74573_/X _83030_/D sky130_fd_sc_hd__o21ai_4
X_40966_ _82299_/Q _40932_/X _40966_/X sky130_fd_sc_hd__or2_4
X_71786_ _71235_/A _71672_/C _71785_/X _71786_/Y sky130_fd_sc_hd__nand3_4
X_79101_ _79086_/B _79101_/Y sky130_fd_sc_hd__inv_2
X_76313_ _76300_/Y _76301_/Y _76302_/Y _76313_/X sky130_fd_sc_hd__o21a_4
X_42705_ _42704_/Y _87761_/D sky130_fd_sc_hd__inv_2
X_49261_ _49261_/A _50781_/B _49261_/Y sky130_fd_sc_hd__nand2_4
X_73525_ _73523_/X _73524_/Y _73367_/X _73525_/Y sky130_fd_sc_hd__a21oi_4
X_46473_ _46467_/Y _46445_/X _46472_/X _86734_/D sky130_fd_sc_hd__a21oi_4
X_70737_ _70736_/Y _70755_/A sky130_fd_sc_hd__inv_2
X_58459_ _84843_/Q _58459_/Y sky130_fd_sc_hd__inv_2
X_77293_ _77292_/Y _77296_/A sky130_fd_sc_hd__inv_2
X_43685_ _43685_/A _43685_/X sky130_fd_sc_hd__buf_2
X_40897_ _40897_/A _40842_/X _40897_/X sky130_fd_sc_hd__or2_4
X_48212_ _48212_/A _53488_/B sky130_fd_sc_hd__buf_2
X_79032_ _79021_/B _79021_/A _79032_/X sky130_fd_sc_hd__and2_4
X_45424_ _45422_/Y _45388_/X _45390_/X _45423_/Y _45424_/X sky130_fd_sc_hd__a211o_4
X_76244_ _81352_/Q _81608_/D _81320_/D sky130_fd_sc_hd__xor2_4
X_42636_ _40939_/X _42631_/X _69147_/B _42634_/X _87794_/D sky130_fd_sc_hd__a2bb2o_4
X_49192_ _49192_/A _50719_/B sky130_fd_sc_hd__buf_2
X_61470_ _61317_/A _61484_/C sky130_fd_sc_hd__buf_2
X_73456_ _73163_/X _83054_/Q _73385_/X _73455_/X _73456_/X sky130_fd_sc_hd__a211o_4
X_70668_ _70758_/A _70579_/Y _70827_/B _70668_/D _70669_/A sky130_fd_sc_hd__nand4_4
X_48143_ _86563_/Q _48103_/X _48142_/Y _48143_/Y sky130_fd_sc_hd__o21ai_4
X_60421_ _60515_/B _60421_/B _60570_/A _60515_/C _60532_/A sky130_fd_sc_hd__and4_4
X_72407_ _72339_/X _85321_/Q _72386_/X _72407_/X sky130_fd_sc_hd__o21a_4
X_45355_ _55713_/B _45354_/X _45311_/X _45355_/X sky130_fd_sc_hd__o21a_4
X_76175_ _76175_/A _76175_/Y sky130_fd_sc_hd__inv_2
X_42567_ _42566_/Y _42567_/Y sky130_fd_sc_hd__inv_2
X_73387_ _73163_/X _83057_/Q _73385_/X _73386_/X _73387_/X sky130_fd_sc_hd__a211o_4
X_70599_ _70710_/A _70613_/B _74533_/D _70594_/X _70599_/Y sky130_fd_sc_hd__nand4_4
Xclkbuf_7_92_0_CLK clkbuf_7_93_0_CLK/A clkbuf_7_92_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_44306_ _44305_/X _74095_/B sky130_fd_sc_hd__buf_2
X_63140_ _63138_/Y _63139_/X _63114_/X _63140_/Y sky130_fd_sc_hd__a21oi_4
X_75126_ _75124_/X _75127_/C _81062_/Q _75126_/X sky130_fd_sc_hd__a21o_4
X_41518_ _81173_/Q _41471_/B _41518_/X sky130_fd_sc_hd__or2_4
X_60352_ _79629_/A _60349_/X _60351_/X _60352_/X sky130_fd_sc_hd__o21a_4
X_72338_ _72299_/X _72335_/Y _72336_/Y _72337_/X _72303_/X _72338_/X
+ sky130_fd_sc_hd__o32a_4
X_48074_ _66238_/B _48049_/X _48073_/Y _48074_/Y sky130_fd_sc_hd__o21ai_4
X_45286_ _56442_/C _45252_/X _45285_/X _45286_/Y sky130_fd_sc_hd__o21ai_4
X_42498_ _42498_/A _87845_/D sky130_fd_sc_hd__inv_2
X_47025_ _47008_/A _52807_/B _47025_/Y sky130_fd_sc_hd__nand2_4
X_44237_ _44236_/X _57126_/A sky130_fd_sc_hd__buf_2
X_63071_ _79456_/A _63008_/X _63070_/Y _84356_/D sky130_fd_sc_hd__a21o_4
X_75057_ _81150_/D _75046_/B _75057_/Y sky130_fd_sc_hd__nand2_4
X_79934_ _79934_/A _79944_/A sky130_fd_sc_hd__inv_2
X_41449_ _41411_/X _41449_/X sky130_fd_sc_hd__buf_2
X_60283_ _60233_/Y _60159_/A _60218_/A _60300_/C sky130_fd_sc_hd__nand3_4
X_72269_ _72266_/Y _72268_/Y _72185_/X _72269_/X sky130_fd_sc_hd__a21o_4
X_62022_ _62022_/A _63598_/A sky130_fd_sc_hd__inv_2
X_74008_ _43078_/Y _72900_/X _73894_/X _74007_/Y _74008_/X sky130_fd_sc_hd__a211o_4
X_44168_ _44012_/A _44244_/A sky130_fd_sc_hd__inv_2
X_79865_ _79861_/X _79865_/B _79875_/B sky130_fd_sc_hd__xor2_4
X_43119_ _87568_/Q _43119_/Y sky130_fd_sc_hd__inv_2
X_66830_ _66785_/A _66830_/B _66830_/X sky130_fd_sc_hd__and2_4
X_78816_ _79122_/A _79122_/B _78818_/C _78816_/Y sky130_fd_sc_hd__a21oi_4
X_48976_ _48976_/A _48976_/B _48976_/Y sky130_fd_sc_hd__nand2_4
X_44099_ _44098_/X _44099_/X sky130_fd_sc_hd__buf_2
X_79796_ _84225_/Q _72214_/A _79796_/X sky130_fd_sc_hd__xor2_4
X_47927_ _47904_/X _46350_/A _47926_/X _48221_/A sky130_fd_sc_hd__o21ai_4
X_66761_ _87947_/Q _66759_/X _66688_/X _66760_/X _66761_/X sky130_fd_sc_hd__a211o_4
X_78747_ _78747_/A _78746_/Y _82782_/D sky130_fd_sc_hd__xor2_4
X_63973_ _61500_/X _63908_/B _64003_/C _63908_/D _63973_/Y sky130_fd_sc_hd__nand4_4
X_75959_ _75952_/Y _75957_/Y _75958_/Y _75963_/C sky130_fd_sc_hd__a21o_4
X_68500_ _68497_/X _68499_/X _68477_/X _68500_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_7_30_0_CLK clkbuf_7_31_0_CLK/A clkbuf_8_61_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_65712_ _65700_/X _65710_/Y _65711_/Y _65712_/Y sky130_fd_sc_hd__o21ai_4
X_62924_ _62644_/X _58184_/A _62924_/C _60220_/A _62924_/X sky130_fd_sc_hd__and4_4
X_69480_ _69605_/A _69480_/B _69480_/X sky130_fd_sc_hd__and2_4
X_47858_ _47857_/X _47887_/A sky130_fd_sc_hd__buf_2
X_78678_ _82811_/Q _78682_/A sky130_fd_sc_hd__inv_2
X_66692_ _87438_/Q _66642_/X _66643_/X _66691_/X _66692_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_8_170_0_CLK clkbuf_7_85_0_CLK/X clkbuf_9_341_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_68431_ _68409_/A _88273_/Q _68431_/X sky130_fd_sc_hd__and2_4
X_46809_ _82957_/Q _46809_/Y sky130_fd_sc_hd__inv_2
X_65643_ _65637_/X _65641_/X _65642_/X _65646_/A sky130_fd_sc_hd__a21o_4
X_77629_ _82237_/Q _77629_/Y sky130_fd_sc_hd__inv_2
X_62855_ _58474_/A _62841_/X _60309_/C _60254_/B _62855_/Y sky130_fd_sc_hd__nand4_4
X_47789_ _47799_/A _53246_/B _47789_/Y sky130_fd_sc_hd__nand2_4
X_49528_ _49537_/A _49516_/B _49522_/C _52742_/D _49528_/X sky130_fd_sc_hd__and4_4
X_61806_ _61839_/A _61791_/B _61732_/X _63066_/B _61806_/X sky130_fd_sc_hd__and4_4
X_80640_ THREAD_COUNT[2] _80640_/LO sky130_fd_sc_hd__conb_1
X_68362_ _68360_/X _68361_/Y _68362_/Y sky130_fd_sc_hd__nor2_4
X_65574_ _65572_/Y _65529_/X _65573_/X _84192_/D sky130_fd_sc_hd__a21o_4
X_62786_ _60274_/X _62834_/D sky130_fd_sc_hd__buf_2
Xclkbuf_7_45_0_CLK clkbuf_6_22_0_CLK/X clkbuf_8_91_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_67313_ _67312_/X _67313_/X sky130_fd_sc_hd__buf_2
X_64525_ _64474_/X _64525_/B _64525_/C _64525_/X sky130_fd_sc_hd__and3_4
X_61737_ _61330_/X _62183_/A _59810_/A _59754_/A _61750_/B sky130_fd_sc_hd__nand4_4
X_49459_ _58800_/B _49443_/X _49458_/Y _49459_/Y sky130_fd_sc_hd__o21ai_4
X_80571_ _80562_/B _80561_/X _80571_/X sky130_fd_sc_hd__and2_4
Xclkbuf_8_185_0_CLK clkbuf_7_92_0_CLK/X clkbuf_9_370_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_68293_ _82638_/D _68279_/X _68292_/X _83990_/D sky130_fd_sc_hd__a21bo_4
Xclkbuf_10_180_0_CLK clkbuf_9_90_0_CLK/X _83333_/CLK sky130_fd_sc_hd__clkbuf_1
X_82310_ _80835_/CLK _77028_/B _82310_/Q sky130_fd_sc_hd__dfxtp_4
X_67244_ _67126_/X _67266_/A sky130_fd_sc_hd__buf_2
X_52470_ _52438_/A _52470_/X sky130_fd_sc_hd__buf_2
X_64456_ _64455_/X _84892_/Q _64456_/C _64456_/Y sky130_fd_sc_hd__nand3_4
X_83290_ _85536_/CLK _83290_/D _83290_/Q sky130_fd_sc_hd__dfxtp_4
X_61668_ _58360_/A _61598_/X _61677_/C _72563_/B _61669_/A sky130_fd_sc_hd__nand4_4
X_51421_ _51149_/A _51421_/X sky130_fd_sc_hd__buf_2
X_63407_ _63456_/A _63456_/B _80588_/B _63407_/Y sky130_fd_sc_hd__nor3_4
X_82241_ _82531_/CLK _82273_/Q _82241_/Q sky130_fd_sc_hd__dfxtp_4
X_60619_ _60619_/A _60622_/C sky130_fd_sc_hd__inv_2
X_67175_ _67172_/X _67174_/X _67175_/Y sky130_fd_sc_hd__nand2_4
X_64387_ _64375_/Y _64385_/X _64386_/X _64387_/X sky130_fd_sc_hd__o21a_4
X_61599_ _61317_/A _61677_/C sky130_fd_sc_hd__buf_2
X_54140_ _54249_/A _54140_/X sky130_fd_sc_hd__buf_2
X_66126_ _65486_/A _66181_/A sky130_fd_sc_hd__buf_2
X_51352_ _52533_/A _51352_/B _51352_/C _51352_/X sky130_fd_sc_hd__and3_4
X_63338_ _79169_/B _63338_/Y sky130_fd_sc_hd__inv_2
X_82172_ _81216_/CLK _84164_/Q _82172_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_195_0_CLK clkbuf_9_97_0_CLK/X _84276_/CLK sky130_fd_sc_hd__clkbuf_1
X_50303_ _86227_/Q _50282_/X _50302_/Y _50303_/Y sky130_fd_sc_hd__o21ai_4
X_81123_ _81179_/CLK _81123_/D _40751_/A sky130_fd_sc_hd__dfxtp_4
X_54071_ _54031_/A _54071_/B _54071_/Y sky130_fd_sc_hd__nand2_4
X_66057_ _65880_/A _66057_/X sky130_fd_sc_hd__buf_2
X_51283_ _51298_/A _46361_/A _51283_/X sky130_fd_sc_hd__and2_4
X_63269_ _84339_/Q _63258_/X _63268_/Y _84339_/D sky130_fd_sc_hd__a21o_4
X_86980_ _88345_/CLK _86980_/D _44738_/A sky130_fd_sc_hd__dfxtp_4
X_53022_ _85711_/Q _53010_/X _53021_/Y _53022_/Y sky130_fd_sc_hd__o21ai_4
X_65008_ _65004_/X _65056_/B _65007_/X _65019_/A sky130_fd_sc_hd__nand3_4
X_50234_ _50230_/A _50234_/B _50234_/Y sky130_fd_sc_hd__nand2_4
X_85931_ _86091_/CLK _51871_/Y _85931_/Q sky130_fd_sc_hd__dfxtp_4
X_81054_ _84276_/CLK _75513_/X _81054_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_123_0_CLK clkbuf_7_61_0_CLK/X clkbuf_9_247_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_80005_ _84930_/Q _84178_/Q _80005_/X sky130_fd_sc_hd__xor2_4
X_57830_ _57826_/Y _57828_/Y _57829_/X _57830_/X sky130_fd_sc_hd__a21o_4
X_69816_ _70001_/A _69816_/X sky130_fd_sc_hd__buf_2
X_50165_ _86251_/Q _50162_/X _50164_/Y _50165_/Y sky130_fd_sc_hd__o21ai_4
X_85862_ _86499_/CLK _85862_/D _85862_/Q sky130_fd_sc_hd__dfxtp_4
X_87601_ _88111_/CLK _43029_/Y _73599_/A sky130_fd_sc_hd__dfxtp_4
X_84813_ _82394_/CLK _84813_/D _84813_/Q sky130_fd_sc_hd__dfxtp_4
X_57761_ _45926_/X _57761_/X sky130_fd_sc_hd__buf_2
X_69747_ _69747_/A _69747_/X sky130_fd_sc_hd__buf_2
X_50096_ _86265_/Q _50088_/X _50095_/Y _50096_/Y sky130_fd_sc_hd__o21ai_4
X_54973_ _54973_/A _54974_/C sky130_fd_sc_hd__buf_2
X_66959_ _66912_/A _66959_/B _66959_/X sky130_fd_sc_hd__and2_4
X_85793_ _83685_/CLK _52581_/Y _85793_/Q sky130_fd_sc_hd__dfxtp_4
X_59500_ _59500_/A _59500_/Y sky130_fd_sc_hd__inv_2
X_56712_ _56775_/A _56713_/A sky130_fd_sc_hd__buf_2
X_87532_ _87544_/CLK _43221_/Y _87532_/Q sky130_fd_sc_hd__dfxtp_4
X_53924_ _85541_/Q _53921_/X _53923_/Y _53924_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_8_138_0_CLK clkbuf_7_69_0_CLK/X clkbuf_9_277_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_84744_ _83438_/CLK _84744_/D _84744_/Q sky130_fd_sc_hd__dfxtp_4
X_57692_ _44151_/X _57692_/B _57692_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_10_133_0_CLK clkbuf_9_66_0_CLK/X _83842_/CLK sky130_fd_sc_hd__clkbuf_1
X_81956_ _82339_/CLK _81956_/D _77890_/B sky130_fd_sc_hd__dfxtp_4
X_69678_ _69678_/A _69678_/X sky130_fd_sc_hd__buf_2
X_59431_ _59430_/Y _59424_/B _59431_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_763_0_CLK clkbuf_9_381_0_CLK/X _87525_/CLK sky130_fd_sc_hd__clkbuf_1
X_56643_ _56642_/Y _56643_/X sky130_fd_sc_hd__buf_2
X_80907_ _83918_/CLK _80907_/D _75649_/A sky130_fd_sc_hd__dfxtp_4
X_68629_ _68625_/X _68628_/X _68558_/X _68629_/X sky130_fd_sc_hd__a21o_4
X_87463_ _87149_/CLK _87463_/D _87463_/Q sky130_fd_sc_hd__dfxtp_4
X_53855_ _53853_/Y _53838_/X _53854_/Y _53855_/Y sky130_fd_sc_hd__a21boi_4
X_84675_ _84671_/CLK _84675_/D _80186_/A sky130_fd_sc_hd__dfxtp_4
X_81887_ _81857_/CLK _78078_/X _81887_/Q sky130_fd_sc_hd__dfxtp_4
X_86414_ _86414_/CLK _49305_/Y _65109_/B sky130_fd_sc_hd__dfxtp_4
X_40820_ _40820_/A _40820_/X sky130_fd_sc_hd__buf_2
X_52806_ _52804_/Y _52783_/X _52805_/X _52806_/Y sky130_fd_sc_hd__a21oi_4
X_59362_ _59237_/X _59360_/Y _59361_/Y _59301_/X _59241_/X _59362_/X
+ sky130_fd_sc_hd__o32a_4
X_71640_ _59493_/Y _71628_/X _71639_/Y _71640_/Y sky130_fd_sc_hd__o21ai_4
X_83626_ _83627_/CLK _71044_/Y _47668_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_254_0_CLK clkbuf_9_255_0_CLK/A clkbuf_9_254_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_56574_ _56564_/B _56564_/A _56574_/Y sky130_fd_sc_hd__xnor2_4
X_80838_ _80746_/CLK _80870_/Q _74869_/B sky130_fd_sc_hd__dfxtp_4
X_87394_ _87394_/CLK _43492_/X _87394_/Q sky130_fd_sc_hd__dfxtp_4
X_53786_ _53786_/A _48887_/Y _53786_/Y sky130_fd_sc_hd__nand2_4
X_50998_ _51003_/A _50998_/B _50998_/Y sky130_fd_sc_hd__nand2_4
X_58313_ _58408_/A _58326_/B sky130_fd_sc_hd__buf_2
X_55525_ _45553_/A _55522_/X _55523_/X _55524_/Y _55525_/X sky130_fd_sc_hd__a211o_4
X_86345_ _82381_/CLK _86345_/D _86345_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_148_0_CLK clkbuf_9_74_0_CLK/X _81695_/CLK sky130_fd_sc_hd__clkbuf_1
X_40751_ _40751_/A _40765_/B _40751_/X sky130_fd_sc_hd__or2_4
X_52737_ _52684_/A _52737_/X sky130_fd_sc_hd__buf_2
X_59293_ _59292_/X _85641_/Q _59205_/X _59293_/X sky130_fd_sc_hd__o21a_4
X_83557_ _86237_/CLK _71253_/Y _47880_/A sky130_fd_sc_hd__dfxtp_4
X_71571_ _71164_/B _71574_/C sky130_fd_sc_hd__buf_2
X_80769_ _83944_/CLK _80769_/D _75008_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_778_0_CLK clkbuf_9_389_0_CLK/X _82047_/CLK sky130_fd_sc_hd__clkbuf_1
X_73310_ _73407_/A _73310_/B _73310_/X sky130_fd_sc_hd__and2_4
XPHY_700 sky130_fd_sc_hd__decap_3
X_70522_ _70526_/A _74529_/A _70962_/C _70522_/Y sky130_fd_sc_hd__nand3_4
X_58244_ _58241_/X _58248_/B _58244_/Y sky130_fd_sc_hd__nor2_4
X_82508_ _82702_/CLK _82508_/D _82508_/Q sky130_fd_sc_hd__dfxtp_4
X_43470_ _43470_/A _43470_/Y sky130_fd_sc_hd__inv_2
X_55456_ _45597_/A _55453_/X _44047_/X _55455_/Y _55456_/X sky130_fd_sc_hd__a211o_4
X_74290_ _72688_/A _74297_/B sky130_fd_sc_hd__buf_2
XPHY_711 sky130_fd_sc_hd__decap_3
X_86276_ _85955_/CLK _86276_/D _72461_/B sky130_fd_sc_hd__dfxtp_4
X_40682_ _40682_/A _40682_/X sky130_fd_sc_hd__buf_2
X_52668_ _85776_/Q _52656_/X _52667_/Y _52668_/Y sky130_fd_sc_hd__o21ai_4
X_83488_ _83372_/CLK _83488_/D _83488_/Q sky130_fd_sc_hd__dfxtp_4
X_42421_ _42421_/A _42421_/Y sky130_fd_sc_hd__inv_2
X_88015_ _87260_/CLK _88015_/D _88015_/Q sky130_fd_sc_hd__dfxtp_4
X_54407_ _85448_/Q _54404_/X _54406_/Y _54407_/Y sky130_fd_sc_hd__o21ai_4
X_73241_ _73237_/X _73240_/X _73241_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_269_0_CLK clkbuf_9_269_0_CLK/A clkbuf_9_269_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_85227_ _85192_/CLK _85227_/D _55783_/B sky130_fd_sc_hd__dfxtp_4
X_51619_ _51619_/A _51619_/B _51608_/X _53144_/D _51619_/X sky130_fd_sc_hd__and4_4
X_70453_ _70907_/B _70827_/B sky130_fd_sc_hd__buf_2
X_58175_ _64282_/A _58217_/B _58175_/Y sky130_fd_sc_hd__nand2_4
X_82439_ _82820_/CLK _79131_/X _82439_/Q sky130_fd_sc_hd__dfxtp_4
X_55387_ _55387_/A _55387_/X sky130_fd_sc_hd__buf_2
X_52599_ _52614_/A _52594_/B _52622_/C _51772_/D _52599_/X sky130_fd_sc_hd__and4_4
X_45140_ _83026_/Q _45141_/A sky130_fd_sc_hd__inv_2
X_57126_ _57126_/A _57158_/C sky130_fd_sc_hd__buf_2
X_42352_ _42352_/A _87908_/D sky130_fd_sc_hd__inv_2
X_54338_ _54366_/A _54338_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_701_0_CLK clkbuf_9_350_0_CLK/X _87888_/CLK sky130_fd_sc_hd__clkbuf_1
X_73172_ _83162_/Q _73079_/X _73171_/Y _83162_/D sky130_fd_sc_hd__a21o_4
X_85158_ _83013_/CLK _85158_/D _56536_/C sky130_fd_sc_hd__dfxtp_4
X_70384_ _70366_/X _70383_/X _70375_/C _70384_/Y sky130_fd_sc_hd__nand3_4
X_41303_ _41302_/X _41283_/X _67411_/B _41284_/X _88240_/D sky130_fd_sc_hd__a2bb2o_4
X_72123_ _72123_/A _72123_/X sky130_fd_sc_hd__buf_2
X_84109_ _84111_/CLK _84109_/D _66509_/C sky130_fd_sc_hd__dfxtp_4
X_45071_ _45052_/X _61447_/B _45070_/X _45071_/Y sky130_fd_sc_hd__o21ai_4
X_57057_ _57056_/Y _56857_/X _56995_/X _57046_/Y _57057_/X sky130_fd_sc_hd__a211o_4
X_42283_ _41529_/X _42271_/X _87941_/Q _42272_/X _87941_/D sky130_fd_sc_hd__a2bb2o_4
X_54269_ _85473_/Q _54266_/X _54268_/Y _54269_/Y sky130_fd_sc_hd__o21ai_4
X_77980_ _77980_/A _77972_/Y _77980_/C _77983_/C sky130_fd_sc_hd__nand3_4
X_85089_ _85089_/CLK _85089_/D _45386_/A sky130_fd_sc_hd__dfxtp_4
X_44022_ _64803_/A _44022_/X sky130_fd_sc_hd__buf_2
X_56008_ _55688_/X _56005_/X _56007_/Y _56008_/Y sky130_fd_sc_hd__o21ai_4
X_41234_ _41233_/X _41234_/X sky130_fd_sc_hd__buf_2
X_72054_ _83294_/Q _72051_/X _72053_/Y _72054_/Y sky130_fd_sc_hd__o21ai_4
X_76931_ _76931_/A _76931_/B _76932_/A sky130_fd_sc_hd__and2_4
X_71005_ _71005_/A _71064_/B sky130_fd_sc_hd__buf_2
Xclkbuf_10_716_0_CLK clkbuf_9_358_0_CLK/X _87083_/CLK sky130_fd_sc_hd__clkbuf_1
X_48830_ _48826_/Y _48813_/X _48829_/X _86475_/D sky130_fd_sc_hd__a21oi_4
X_79650_ _79648_/X _79650_/B _79664_/A sky130_fd_sc_hd__xnor2_4
X_41165_ _41165_/A _41165_/X sky130_fd_sc_hd__buf_2
X_76862_ _76862_/A _76862_/B _81465_/D sky130_fd_sc_hd__xnor2_4
X_78601_ _78601_/A _78601_/Y sky130_fd_sc_hd__inv_2
X_75813_ _81020_/Q _80892_/D _80988_/D sky130_fd_sc_hd__xor2_4
Xclkbuf_9_207_0_CLK clkbuf_9_206_0_CLK/A clkbuf_9_207_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_48761_ _50443_/A _48766_/B _48761_/C _48761_/X sky130_fd_sc_hd__and3_4
X_79581_ _79581_/A _79581_/B _79588_/A sky130_fd_sc_hd__xor2_4
X_57959_ _58676_/A _58039_/B sky130_fd_sc_hd__buf_2
X_45973_ _40399_/Y _45963_/X _86832_/Q _45964_/X _86832_/D sky130_fd_sc_hd__a2bb2o_4
X_41096_ _41159_/A _41096_/B _41096_/X sky130_fd_sc_hd__or2_4
X_76793_ _76806_/A _76792_/Y _76801_/A sky130_fd_sc_hd__xor2_4
X_47712_ _47707_/Y _47698_/X _47711_/X _86606_/D sky130_fd_sc_hd__a21oi_4
X_78532_ _82513_/Q _82769_/D _82481_/D sky130_fd_sc_hd__xor2_4
X_44924_ _44916_/X _44921_/X _44923_/Y _44924_/Y sky130_fd_sc_hd__a21oi_4
X_75744_ _75742_/Y _75743_/Y _75747_/A sky130_fd_sc_hd__xor2_4
X_48692_ _48685_/Y _48651_/X _48691_/X _48692_/Y sky130_fd_sc_hd__a21oi_4
X_60970_ _60969_/X _60835_/X _60970_/C _60970_/X sky130_fd_sc_hd__or3_4
X_72956_ _73352_/A _73132_/A sky130_fd_sc_hd__buf_2
X_47643_ _81237_/Q _55026_/D sky130_fd_sc_hd__inv_2
X_71907_ _71894_/Y _71928_/D sky130_fd_sc_hd__buf_2
X_59629_ _59629_/A _59961_/A sky130_fd_sc_hd__buf_2
X_78463_ _78463_/A _78463_/B _78464_/A sky130_fd_sc_hd__and2_4
X_44855_ _44855_/A _86918_/D sky130_fd_sc_hd__inv_2
X_75675_ _81005_/Q _75675_/B _75675_/X sky130_fd_sc_hd__xor2_4
X_72887_ _83173_/Q _72794_/X _72886_/Y _83173_/D sky130_fd_sc_hd__a21o_4
X_77414_ _77412_/X _77413_/Y _77415_/A sky130_fd_sc_hd__and2_4
X_43806_ _43806_/A _43806_/Y sky130_fd_sc_hd__inv_2
X_62640_ _62910_/A _60360_/X _62640_/C _62886_/A sky130_fd_sc_hd__nand3_4
X_74626_ _45381_/A _74625_/A _74625_/Y _74626_/Y sky130_fd_sc_hd__o21ai_4
X_47574_ _47574_/A _53127_/B _47574_/Y sky130_fd_sc_hd__nand2_4
X_71838_ _71825_/X _83357_/Q _71837_/X _83357_/D sky130_fd_sc_hd__a21o_4
X_78394_ _78394_/A _78394_/B _78394_/C _78426_/B sky130_fd_sc_hd__nand3_4
X_44786_ _41392_/Y _44774_/X _86955_/Q _44775_/X _86955_/D sky130_fd_sc_hd__a2bb2o_4
X_41998_ _41998_/A _41998_/X sky130_fd_sc_hd__buf_2
X_49313_ _49311_/Y _49281_/X _49312_/X _49313_/Y sky130_fd_sc_hd__a21oi_4
X_46525_ _47904_/A _46525_/X sky130_fd_sc_hd__buf_2
X_77345_ _77345_/A _77345_/B _77371_/C sky130_fd_sc_hd__nand2_4
X_43737_ _43673_/A _43737_/X sky130_fd_sc_hd__buf_2
X_62571_ _61627_/B _62548_/C _62507_/X _62478_/X _62570_/X _62571_/X
+ sky130_fd_sc_hd__a41o_4
X_74557_ _46155_/X _74553_/X _56030_/X _74554_/X _74557_/X sky130_fd_sc_hd__a211o_4
X_40949_ _40512_/X _81727_/Q _40948_/X _40950_/A sky130_fd_sc_hd__o21a_4
X_71769_ _71762_/X _83383_/Q _71768_/X _83383_/D sky130_fd_sc_hd__a21o_4
Xclkbuf_4_7_0_CLK clkbuf_4_7_0_CLK/A clkbuf_4_7_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_64310_ _58314_/A _64308_/X _64309_/Y _64310_/Y sky130_fd_sc_hd__o21ai_4
X_49244_ _49242_/Y _49214_/X _49243_/Y _49244_/Y sky130_fd_sc_hd__a21boi_4
X_61522_ _84865_/Q _61522_/X sky130_fd_sc_hd__buf_2
X_73508_ _42061_/Y _72974_/X _73393_/X _73507_/Y _73508_/X sky130_fd_sc_hd__a211o_4
X_46456_ _46455_/Y _51324_/B sky130_fd_sc_hd__buf_2
X_65290_ _65178_/X _83287_/Q _65239_/X _65289_/X _65290_/X sky130_fd_sc_hd__a211o_4
X_77276_ _77277_/B _77276_/Y sky130_fd_sc_hd__inv_2
X_43668_ _40742_/X _43659_/X _69055_/B _43661_/X _43668_/X sky130_fd_sc_hd__a2bb2o_4
X_74488_ _48644_/A _74501_/B _74501_/C _74488_/X sky130_fd_sc_hd__and3_4
X_79015_ _79003_/Y _82520_/D sky130_fd_sc_hd__inv_2
X_45407_ _45400_/X _45404_/X _45406_/Y _45407_/Y sky130_fd_sc_hd__a21oi_4
X_64241_ _79863_/B _63258_/X _64240_/X _84263_/D sky130_fd_sc_hd__a21o_4
X_76227_ _81256_/Q _81512_/D _76232_/A sky130_fd_sc_hd__nor2_4
X_42619_ _42619_/A _42619_/Y sky130_fd_sc_hd__inv_2
X_61453_ _61453_/A _61453_/Y sky130_fd_sc_hd__inv_2
X_49175_ _49175_/A _49176_/A sky130_fd_sc_hd__inv_2
X_73439_ _69918_/B _73319_/X _72890_/X _73438_/Y _73439_/X sky130_fd_sc_hd__a211o_4
X_46387_ _46387_/A _49265_/B _46387_/Y sky130_fd_sc_hd__nand2_4
X_43599_ _87345_/Q _68418_/B sky130_fd_sc_hd__inv_2
X_48126_ _82341_/Q _48086_/B _48126_/X sky130_fd_sc_hd__or2_4
X_60404_ _60387_/A _60404_/B _60404_/C _60387_/C _60404_/Y sky130_fd_sc_hd__nand4_4
X_45338_ _56267_/C _45297_/X _45337_/X _45338_/Y sky130_fd_sc_hd__o21ai_4
X_64172_ _61675_/B _64172_/B _64172_/C _64172_/D _64172_/Y sky130_fd_sc_hd__nand4_4
X_76158_ _76159_/A _76158_/B _76158_/X sky130_fd_sc_hd__or2_4
X_61384_ _61384_/A _61384_/B _79153_/B _61384_/Y sky130_fd_sc_hd__nor3_4
X_63123_ _60484_/A _63124_/D sky130_fd_sc_hd__buf_2
X_75109_ _75109_/A _75109_/B _75110_/A sky130_fd_sc_hd__nor2_4
X_48057_ _47971_/X _82924_/Q _48056_/X _48058_/B sky130_fd_sc_hd__o21ai_4
X_60335_ _62644_/A _60239_/B _60189_/A _60335_/Y sky130_fd_sc_hd__nand3_4
X_45269_ _45709_/A _45269_/X sky130_fd_sc_hd__buf_2
X_68980_ _68770_/X _68980_/B _68980_/X sky130_fd_sc_hd__and2_4
X_76089_ _76086_/Y _76089_/B _76090_/B sky130_fd_sc_hd__xor2_4
X_47008_ _47008_/A _52799_/B _47008_/Y sky130_fd_sc_hd__nand2_4
X_67931_ _67928_/X _67930_/X _67858_/X _67934_/A sky130_fd_sc_hd__a21o_4
X_79917_ _79914_/B _79903_/Y _79911_/Y _79928_/A sky130_fd_sc_hd__a21oi_4
X_63054_ _63054_/A _63081_/B _63081_/C _63033_/D _63054_/X sky130_fd_sc_hd__or4_4
X_60266_ _59875_/X _60233_/Y _60263_/Y _60264_/Y _60265_/X _84644_/D
+ sky130_fd_sc_hd__o41a_4
X_62005_ _62005_/A _63586_/A sky130_fd_sc_hd__inv_2
X_67862_ _67859_/X _67861_/X _67862_/Y sky130_fd_sc_hd__nand2_4
X_79848_ _79844_/X _79866_/B _79875_/A sky130_fd_sc_hd__xor2_4
X_60197_ _60170_/A _60253_/A _60197_/C _60189_/Y _60198_/A sky130_fd_sc_hd__and4_4
X_69601_ _69579_/X _69599_/Y _69516_/X _69600_/Y _69601_/X sky130_fd_sc_hd__a211o_4
X_66813_ _66769_/A _88137_/Q _66813_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_1020_0_CLK clkbuf_9_510_0_CLK/X _83311_/CLK sky130_fd_sc_hd__clkbuf_1
X_48959_ _48959_/A _48959_/B _50599_/B sky130_fd_sc_hd__nor2_4
X_79779_ _79770_/Y _79766_/X _79778_/X _79780_/B sky130_fd_sc_hd__a21boi_4
X_67793_ _67793_/A _67793_/B _67793_/X sky130_fd_sc_hd__and2_4
X_81810_ _81631_/CLK _81618_/Q _81810_/Q sky130_fd_sc_hd__dfxtp_4
X_69532_ _88022_/Q _69424_/X _69465_/X _69531_/X _69532_/X sky130_fd_sc_hd__a211o_4
X_66744_ _66625_/A _66795_/A sky130_fd_sc_hd__buf_2
X_51970_ _51947_/A _50268_/B _51970_/Y sky130_fd_sc_hd__nand2_4
X_63956_ _61939_/X _63955_/X _63905_/C _63892_/D _63956_/Y sky130_fd_sc_hd__nand4_4
X_82790_ _82665_/CLK _82822_/Q _78360_/B sky130_fd_sc_hd__dfxtp_4
X_50921_ _50932_/A _46685_/X _50921_/Y sky130_fd_sc_hd__nand2_4
X_62907_ _62965_/A _62935_/B _63629_/B _62907_/Y sky130_fd_sc_hd__nand3_4
X_81741_ _82642_/CLK _81741_/D _81741_/Q sky130_fd_sc_hd__dfxtp_4
X_69463_ _69423_/X _69461_/Y _69405_/X _69462_/Y _69463_/X sky130_fd_sc_hd__a211o_4
X_66675_ _66794_/A _66675_/X sky130_fd_sc_hd__buf_2
X_63887_ _60906_/X _63902_/C sky130_fd_sc_hd__buf_2
X_68414_ _68377_/A _68414_/X sky130_fd_sc_hd__buf_2
X_53640_ _53793_/A _53778_/A sky130_fd_sc_hd__buf_2
X_65626_ _65779_/A _86484_/Q _65626_/X sky130_fd_sc_hd__and2_4
X_84460_ _82436_/CLK _84460_/D _79128_/B sky130_fd_sc_hd__dfxtp_4
X_50852_ _50806_/A _50852_/B _50852_/Y sky130_fd_sc_hd__nand2_4
X_62838_ _62893_/A _62838_/X sky130_fd_sc_hd__buf_2
X_81672_ _81282_/CLK _79993_/X _76847_/A sky130_fd_sc_hd__dfxtp_4
X_69394_ _69286_/A _87776_/Q _69394_/X sky130_fd_sc_hd__and2_4
X_83411_ _83414_/CLK _83411_/D _83411_/Q sky130_fd_sc_hd__dfxtp_4
X_80623_ _80623_/A _80615_/Y _80623_/X sky130_fd_sc_hd__or2_4
X_68345_ _66560_/X _69645_/A sky130_fd_sc_hd__buf_2
X_53571_ _53568_/Y _53537_/X _53570_/X _85611_/D sky130_fd_sc_hd__a21oi_4
X_65557_ _65557_/A _65556_/Y _65557_/Y sky130_fd_sc_hd__nand2_4
X_84391_ _84392_/CLK _62688_/Y _84391_/Q sky130_fd_sc_hd__dfxtp_4
X_50783_ _50764_/A _52478_/B _50783_/Y sky130_fd_sc_hd__nand2_4
X_62769_ _62979_/A _62819_/A sky130_fd_sc_hd__buf_2
X_55310_ _55304_/X _55308_/X _55309_/X _55310_/X sky130_fd_sc_hd__a21o_4
X_86130_ _86139_/CLK _50803_/Y _86130_/Q sky130_fd_sc_hd__dfxtp_4
X_52522_ _52518_/A _52522_/B _52522_/Y sky130_fd_sc_hd__nand2_4
X_64508_ _64508_/A _64741_/B sky130_fd_sc_hd__buf_2
X_83342_ _83491_/CLK _71882_/X _83342_/Q sky130_fd_sc_hd__dfxtp_4
X_56290_ _56360_/A _56290_/X sky130_fd_sc_hd__buf_2
X_80554_ _80551_/Y _80534_/Y _80553_/X _80554_/Y sky130_fd_sc_hd__o21ai_4
X_68276_ _67705_/X _67708_/X _68239_/X _68276_/Y sky130_fd_sc_hd__a21oi_4
X_65488_ _65484_/X _86205_/Q _65400_/X _65487_/X _65488_/X sky130_fd_sc_hd__a211o_4
X_55241_ _55228_/Y _55241_/B _55243_/A sky130_fd_sc_hd__nand2_4
X_67227_ _67250_/A _67227_/B _67227_/X sky130_fd_sc_hd__and2_4
X_86061_ _85741_/CLK _51172_/Y _86061_/Q sky130_fd_sc_hd__dfxtp_4
X_52453_ _85819_/Q _52438_/X _52452_/Y _52453_/Y sky130_fd_sc_hd__o21ai_4
X_83273_ _85335_/CLK _83273_/D _72214_/A sky130_fd_sc_hd__dfxtp_4
X_64439_ _58261_/Y _64423_/X _64438_/Y _64439_/Y sky130_fd_sc_hd__o21ai_4
X_80485_ _80494_/A _80494_/B _80485_/Y sky130_fd_sc_hd__xnor2_4
X_85012_ _85075_/CLK _85012_/D _45599_/A sky130_fd_sc_hd__dfxtp_4
X_51404_ _51403_/X _52931_/B _51404_/Y sky130_fd_sc_hd__nand2_4
X_82224_ _81857_/CLK _82256_/Q _77422_/A sky130_fd_sc_hd__dfxtp_4
X_55172_ _55172_/A _55172_/X sky130_fd_sc_hd__buf_2
X_67158_ _87419_/Q _67156_/X _67106_/X _67157_/X _67158_/X sky130_fd_sc_hd__a211o_4
X_52384_ _65225_/B _52372_/X _52383_/Y _52384_/Y sky130_fd_sc_hd__o21ai_4
X_54123_ _54123_/A _54123_/B _54118_/X _52954_/D _54123_/X sky130_fd_sc_hd__and4_4
X_66109_ _66164_/A _66164_/B _66109_/C _66109_/Y sky130_fd_sc_hd__nor3_4
X_51335_ _51350_/A _50827_/B _51335_/Y sky130_fd_sc_hd__nand2_4
X_82155_ _84220_/CLK _80397_/B _82155_/Q sky130_fd_sc_hd__dfxtp_4
X_67089_ _67086_/X _67088_/X _67015_/X _67089_/Y sky130_fd_sc_hd__a21oi_4
X_59980_ _60781_/A _59980_/X sky130_fd_sc_hd__buf_2
X_81106_ _81070_/CLK _79729_/X _75574_/A sky130_fd_sc_hd__dfxtp_4
X_58931_ _58927_/Y _58930_/Y _58883_/X _58931_/X sky130_fd_sc_hd__a21o_4
X_54054_ _54020_/A _54054_/B _54054_/Y sky130_fd_sc_hd__nand2_4
X_51266_ _50755_/A _51266_/B _51330_/C _51266_/X sky130_fd_sc_hd__and3_4
X_86963_ _86934_/CLK _86963_/D _86963_/Q sky130_fd_sc_hd__dfxtp_4
X_82086_ _81970_/CLK _82086_/D _82086_/Q sky130_fd_sc_hd__dfxtp_4
X_53005_ _52999_/A _53005_/B _53005_/Y sky130_fd_sc_hd__nand2_4
X_50217_ _50217_/A _50217_/Y sky130_fd_sc_hd__inv_2
X_85914_ _86238_/CLK _85914_/D _66006_/B sky130_fd_sc_hd__dfxtp_4
X_81037_ _81061_/CLK _81037_/D _81229_/D sky130_fd_sc_hd__dfxtp_4
X_58862_ _58796_/X _86090_/Q _58861_/X _58862_/Y sky130_fd_sc_hd__o21ai_4
X_51197_ _51191_/X _51192_/B _51197_/C _52887_/D _51197_/X sky130_fd_sc_hd__and4_4
X_86894_ _86896_/CLK _45173_/Y _64411_/B sky130_fd_sc_hd__dfxtp_4
X_57813_ _57811_/X _85404_/Q _57812_/X _57813_/Y sky130_fd_sc_hd__o21ai_4
X_50148_ _50145_/Y _50141_/X _50147_/X _86255_/D sky130_fd_sc_hd__a21oi_4
X_85845_ _85555_/CLK _52329_/Y _85845_/Q sky130_fd_sc_hd__dfxtp_4
X_58793_ _58793_/A _58793_/X sky130_fd_sc_hd__buf_2
X_72810_ _72750_/X _85599_/Q _44130_/X _72809_/X _72810_/X sky130_fd_sc_hd__a211o_4
X_57744_ _44151_/X _86334_/Q _57744_/Y sky130_fd_sc_hd__nor2_4
X_42970_ _43774_/A _42970_/X sky130_fd_sc_hd__buf_2
X_50079_ _50076_/Y _50068_/X _50078_/X _86269_/D sky130_fd_sc_hd__a21oi_4
X_54956_ _54954_/Y _54936_/X _54955_/X _85346_/D sky130_fd_sc_hd__a21oi_4
X_73790_ _53501_/B _73789_/Y _73790_/X sky130_fd_sc_hd__xor2_4
X_85776_ _85778_/CLK _85776_/D _85776_/Q sky130_fd_sc_hd__dfxtp_4
X_82988_ _82987_/CLK _74678_/Y _45727_/A sky130_fd_sc_hd__dfxtp_4
X_87515_ _87273_/CLK _87515_/D _87515_/Q sky130_fd_sc_hd__dfxtp_4
X_41921_ _41887_/X _41919_/X _40646_/X _41920_/Y _41891_/X _88105_/D
+ sky130_fd_sc_hd__o32ai_4
X_53907_ _53905_/Y _53862_/X _53906_/Y _85545_/D sky130_fd_sc_hd__a21boi_4
X_72741_ _73007_/A _72741_/X sky130_fd_sc_hd__buf_2
X_84727_ _84727_/CLK _84727_/D _59456_/A sky130_fd_sc_hd__dfxtp_4
X_57675_ _58230_/A _57674_/Y _57675_/Y sky130_fd_sc_hd__nand2_4
X_81939_ _81954_/CLK _81939_/D _77485_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_9_193_0_CLK clkbuf_8_96_0_CLK/X clkbuf_9_193_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_54887_ _54344_/A _54888_/A sky130_fd_sc_hd__buf_2
X_59414_ _59413_/Y _59415_/A sky130_fd_sc_hd__buf_2
X_44640_ _44714_/A _44640_/X sky130_fd_sc_hd__buf_2
X_56626_ _56626_/A _56626_/X sky130_fd_sc_hd__buf_2
X_87446_ _87446_/CLK _87446_/D _87446_/Q sky130_fd_sc_hd__dfxtp_4
X_75460_ _75442_/Y _75443_/Y _75445_/A _75461_/A sky130_fd_sc_hd__o21a_4
X_41852_ _40520_/X _41847_/X _67183_/B _41848_/X _88122_/D sky130_fd_sc_hd__a2bb2o_4
X_53838_ _53838_/A _53838_/X sky130_fd_sc_hd__buf_2
X_72672_ _72630_/X _72672_/X sky130_fd_sc_hd__buf_2
X_84658_ _84503_/CLK _60126_/Y _84658_/Q sky130_fd_sc_hd__dfxtp_4
X_74411_ _74409_/Y _74405_/X _74410_/X _74411_/Y sky130_fd_sc_hd__a21oi_4
X_40803_ _40802_/X _40793_/X _88332_/Q _40794_/X _88332_/D sky130_fd_sc_hd__a2bb2o_4
X_59345_ _64678_/A _59345_/X sky130_fd_sc_hd__buf_2
X_71623_ _71603_/Y _83434_/Q _71622_/Y _71623_/X sky130_fd_sc_hd__a21o_4
X_83609_ _85554_/CLK _83609_/D _49044_/A sky130_fd_sc_hd__dfxtp_4
X_44571_ _44565_/X _44567_/X _40874_/X _87051_/Q _44568_/X _44571_/Y
+ sky130_fd_sc_hd__o32ai_4
X_56557_ _56556_/Y _55570_/D _72648_/C _72643_/C _56557_/X sky130_fd_sc_hd__and4_4
X_75391_ _80791_/Q _75390_/X _80759_/D sky130_fd_sc_hd__xor2_4
X_41783_ _41782_/X _41750_/X _88150_/Q _41751_/X _88150_/D sky130_fd_sc_hd__a2bb2o_4
X_87377_ _88144_/CLK _87377_/D _87377_/Q sky130_fd_sc_hd__dfxtp_4
X_53769_ _53767_/Y _53747_/X _53768_/X _85572_/D sky130_fd_sc_hd__a21oi_4
X_84589_ _84469_/CLK _60604_/Y _79129_/A sky130_fd_sc_hd__dfxtp_4
X_46310_ _53511_/A _46428_/C sky130_fd_sc_hd__buf_2
X_77130_ _77130_/A _77129_/X _77142_/A sky130_fd_sc_hd__nand2_4
X_43522_ _40331_/X _43513_/X _87378_/Q _43514_/X _87378_/D sky130_fd_sc_hd__a2bb2o_4
X_55508_ _55507_/X _55508_/B _55508_/Y sky130_fd_sc_hd__nor2_4
X_74342_ _74342_/A _74342_/X sky130_fd_sc_hd__buf_2
X_86328_ _86647_/CLK _49762_/Y _57857_/B sky130_fd_sc_hd__dfxtp_4
X_40734_ _40733_/Y _40734_/X sky130_fd_sc_hd__buf_2
X_47290_ _47287_/X _52965_/B _47290_/Y sky130_fd_sc_hd__nand2_4
X_71554_ _71530_/Y _83458_/Q _71553_/Y _83458_/D sky130_fd_sc_hd__a21o_4
X_59276_ _59199_/X _85739_/Q _59263_/X _59276_/X sky130_fd_sc_hd__o21a_4
X_56488_ _56487_/X _56484_/X _56488_/C _56488_/Y sky130_fd_sc_hd__nand3_4
X_70505_ _70696_/B _70758_/B _71136_/A _70506_/A sky130_fd_sc_hd__nor3_4
X_46241_ _40877_/X _82945_/Q _46240_/Y _46241_/X sky130_fd_sc_hd__o21a_4
XPHY_530 sky130_fd_sc_hd__decap_3
X_58227_ _58219_/X _58224_/Y _58226_/Y _58227_/Y sky130_fd_sc_hd__a21oi_4
X_77061_ _77069_/A _82283_/D _77067_/B sky130_fd_sc_hd__xor2_4
X_43453_ _43449_/X _43452_/X _41616_/X _87414_/Q _43434_/X _43454_/A
+ sky130_fd_sc_hd__o32ai_4
X_55439_ _56719_/A _56719_/B _55439_/Y sky130_fd_sc_hd__nand2_4
X_74273_ _73040_/A _86562_/Q _74273_/X sky130_fd_sc_hd__and2_4
X_86259_ _85557_/CLK _50127_/Y _86259_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_541 sky130_fd_sc_hd__decap_3
X_40665_ _40829_/A _82867_/Q _40665_/X sky130_fd_sc_hd__or2_4
Xclkbuf_10_640_0_CLK clkbuf_9_320_0_CLK/X _87471_/CLK sky130_fd_sc_hd__clkbuf_1
X_71485_ _71289_/B _71485_/B _71486_/A sky130_fd_sc_hd__nor2_4
XPHY_552 sky130_fd_sc_hd__decap_3
XPHY_563 sky130_fd_sc_hd__decap_3
X_76012_ _81711_/D _76021_/B _76015_/A sky130_fd_sc_hd__xor2_4
X_42404_ _42401_/X _42397_/X _40440_/X _87879_/Q _42398_/X _42405_/A
+ sky130_fd_sc_hd__o32ai_4
XPHY_574 sky130_fd_sc_hd__decap_3
X_73224_ _57376_/X _73224_/X sky130_fd_sc_hd__buf_2
X_46172_ _46168_/Y _46169_/Y _46171_/Y _46172_/Y sky130_fd_sc_hd__a21oi_4
X_70436_ _48231_/B _70422_/X _70435_/Y _83775_/D sky130_fd_sc_hd__o21ai_4
X_58158_ _84918_/Q _63044_/A sky130_fd_sc_hd__inv_2
XPHY_585 sky130_fd_sc_hd__decap_3
X_43384_ _41429_/X _43371_/X _87449_/Q _43372_/X _87449_/D sky130_fd_sc_hd__a2bb2o_4
XPHY_596 sky130_fd_sc_hd__decap_3
Xclkbuf_9_131_0_CLK clkbuf_8_65_0_CLK/X clkbuf_9_131_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_40596_ _40595_/X _40596_/X sky130_fd_sc_hd__buf_2
X_45123_ _44968_/X _45182_/B sky130_fd_sc_hd__buf_2
X_57109_ _57096_/Y _57109_/X sky130_fd_sc_hd__buf_2
X_42335_ _42335_/A _42335_/Y sky130_fd_sc_hd__inv_2
X_73155_ _44556_/Y _72899_/X _73154_/Y _73155_/X sky130_fd_sc_hd__a21o_4
X_70367_ DATA_TO_HASH[7] _70984_/A sky130_fd_sc_hd__buf_2
X_58089_ _58928_/A _58089_/X sky130_fd_sc_hd__buf_2
X_60120_ _59579_/A _61183_/A _60593_/B _60155_/D sky130_fd_sc_hd__nor3_4
X_72106_ _83283_/Q _72090_/X _72105_/Y _72106_/Y sky130_fd_sc_hd__o21ai_4
X_49931_ _49930_/X _49953_/C sky130_fd_sc_hd__buf_2
X_45054_ _45052_/X _61437_/B _44995_/X _45054_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_655_0_CLK clkbuf_9_327_0_CLK/X _88220_/CLK sky130_fd_sc_hd__clkbuf_1
X_42266_ _42252_/X _42243_/X _41493_/X _87949_/Q _42244_/X _42266_/Y
+ sky130_fd_sc_hd__o32ai_4
X_77963_ _82252_/Q _81964_/Q _81948_/D sky130_fd_sc_hd__xor2_4
X_73086_ _73530_/B _73086_/X sky130_fd_sc_hd__buf_2
X_70298_ _70249_/X _70301_/D sky130_fd_sc_hd__buf_2
X_44005_ _59901_/C _59584_/C _59598_/A _44004_/Y _44005_/X sky130_fd_sc_hd__a2bb2o_4
X_79702_ _79702_/A _79701_/Y _79702_/X sky130_fd_sc_hd__xor2_4
X_41217_ _40413_/X _41513_/A sky130_fd_sc_hd__buf_2
X_60051_ _60064_/A _60081_/B _60051_/C _60051_/Y sky130_fd_sc_hd__nor3_4
X_72037_ _83297_/Q _72016_/X _72036_/Y _72037_/Y sky130_fd_sc_hd__o21ai_4
X_76914_ _76914_/A _76914_/B _81470_/D sky130_fd_sc_hd__xor2_4
X_49862_ _49851_/A _49884_/B _49862_/C _53074_/D _49862_/X sky130_fd_sc_hd__and4_4
Xclkbuf_9_146_0_CLK clkbuf_8_73_0_CLK/X clkbuf_9_146_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_42197_ _41306_/X _42192_/X _87983_/Q _42193_/X _87983_/D sky130_fd_sc_hd__a2bb2o_4
X_77894_ _77885_/A _77872_/Y _77884_/A _77883_/Y _77894_/X sky130_fd_sc_hd__o22a_4
Xclkbuf_9_73_0_CLK clkbuf_9_72_0_CLK/A clkbuf_9_73_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_48813_ _48840_/A _48813_/X sky130_fd_sc_hd__buf_2
X_79633_ _79633_/A _79632_/Y _79633_/X sky130_fd_sc_hd__xor2_4
X_41148_ _41147_/X _41109_/X _88269_/Q _41110_/X _88269_/D sky130_fd_sc_hd__a2bb2o_4
X_76845_ _76845_/A _76845_/B _76845_/X sky130_fd_sc_hd__xor2_4
X_49793_ _49793_/A _52679_/A sky130_fd_sc_hd__buf_2
X_63810_ _63741_/A _63810_/X sky130_fd_sc_hd__buf_2
X_48744_ _48744_/A _48766_/B _48761_/C _48744_/X sky130_fd_sc_hd__and3_4
X_79564_ _79557_/A _79549_/Y _79550_/Y _79564_/Y sky130_fd_sc_hd__a21boi_4
X_45956_ _45955_/X _45957_/A sky130_fd_sc_hd__buf_2
X_41079_ _41013_/A _41079_/X sky130_fd_sc_hd__buf_2
X_64790_ _64637_/X _64913_/B _84227_/Q _64790_/X sky130_fd_sc_hd__and3_4
X_76776_ _76762_/Y _76776_/B _76776_/Y sky130_fd_sc_hd__nand2_4
X_73988_ _68826_/B _72853_/X _45897_/X _73987_/Y _73988_/X sky130_fd_sc_hd__a211o_4
X_78515_ _78515_/A _78514_/Y _78515_/Y sky130_fd_sc_hd__nand2_4
X_44907_ _44907_/A _44907_/X sky130_fd_sc_hd__buf_2
X_63741_ _63741_/A _63741_/X sky130_fd_sc_hd__buf_2
X_75727_ _75727_/A _75726_/Y _75736_/B sky130_fd_sc_hd__xor2_4
X_60953_ _60901_/B _60882_/X _60910_/B _60953_/X sky130_fd_sc_hd__and3_4
X_72939_ _72926_/X _72928_/X _72938_/X _72939_/X sky130_fd_sc_hd__a21o_4
X_48675_ _48675_/A _48676_/A sky130_fd_sc_hd__inv_2
X_79495_ _79491_/Y _79494_/Y _79505_/B sky130_fd_sc_hd__xor2_4
Xclkbuf_9_88_0_CLK clkbuf_9_88_0_CLK/A clkbuf_9_88_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_45887_ _44038_/X _45888_/A sky130_fd_sc_hd__buf_2
X_47626_ _47530_/A _47655_/A sky130_fd_sc_hd__buf_2
X_66460_ _66458_/Y _66459_/Y _60529_/A _66460_/X sky130_fd_sc_hd__a21o_4
X_78446_ _78455_/A _82668_/D _78447_/B sky130_fd_sc_hd__xor2_4
X_44838_ _43927_/X _44838_/X sky130_fd_sc_hd__buf_2
X_63672_ _63655_/A _63672_/B _63672_/C _63595_/D _63672_/X sky130_fd_sc_hd__and4_4
X_75658_ _75658_/A _75657_/Y _75666_/A sky130_fd_sc_hd__xor2_4
X_60884_ _60865_/C _60901_/A sky130_fd_sc_hd__buf_2
X_65411_ _65258_/A _65411_/B _65411_/X sky130_fd_sc_hd__and2_4
X_62623_ _62623_/A _62174_/X _62623_/C _62623_/D _62623_/X sky130_fd_sc_hd__and4_4
X_74609_ _45273_/A _74598_/X _74608_/X _74609_/Y sky130_fd_sc_hd__o21ai_4
X_47557_ _81246_/Q _47558_/A sky130_fd_sc_hd__inv_2
X_66391_ _66391_/A _66417_/B sky130_fd_sc_hd__buf_2
X_78377_ _78374_/X _78375_/Y _78378_/A _78380_/A sky130_fd_sc_hd__a21oi_4
X_44769_ _44766_/X _44767_/X _41340_/X _86965_/Q _44768_/X _44770_/A
+ sky130_fd_sc_hd__o32ai_4
X_75589_ _80820_/Q _75589_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_opt_9_CLK clkbuf_opt_9_CLK/A _84886_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_9_11_0_CLK clkbuf_8_5_0_CLK/X clkbuf_9_11_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_68130_ _66821_/X _66824_/X _68129_/X _68130_/Y sky130_fd_sc_hd__a21oi_4
X_46508_ _52533_/A _46487_/B _46472_/C _46508_/X sky130_fd_sc_hd__and3_4
X_65342_ _65660_/A _65342_/X sky130_fd_sc_hd__buf_2
X_77328_ _77323_/Y _77328_/Y sky130_fd_sc_hd__inv_2
X_62554_ _62551_/X _62553_/X _84402_/Q _62554_/Y sky130_fd_sc_hd__nor3_4
X_47488_ _47483_/Y _47462_/X _47487_/X _86630_/D sky130_fd_sc_hd__a21oi_4
X_49227_ _49225_/Y _49214_/X _49226_/Y _86430_/D sky130_fd_sc_hd__a21boi_4
Xclkbuf_10_608_0_CLK clkbuf_9_304_0_CLK/X _81169_/CLK sky130_fd_sc_hd__clkbuf_1
X_61505_ _61504_/Y _61505_/Y sky130_fd_sc_hd__inv_2
X_68061_ _87137_/Q _68059_/X _67991_/X _68060_/X _68061_/X sky130_fd_sc_hd__a211o_4
X_46439_ _46408_/A _50808_/B _46439_/Y sky130_fd_sc_hd__nand2_4
X_65273_ _64567_/A _65877_/A sky130_fd_sc_hd__buf_2
X_77259_ _77258_/Y _77259_/Y sky130_fd_sc_hd__inv_2
X_62485_ _62483_/X _62541_/B _62485_/C _62485_/Y sky130_fd_sc_hd__nor3_4
X_67012_ _87117_/Q _66988_/X _66919_/X _67011_/X _67012_/X sky130_fd_sc_hd__a211o_4
X_64224_ _64285_/A _64248_/A sky130_fd_sc_hd__buf_2
X_49158_ _53917_/B _50188_/B sky130_fd_sc_hd__buf_2
X_61436_ _61374_/A _61437_/A sky130_fd_sc_hd__buf_2
X_80270_ _84746_/Q _84138_/Q _80270_/X sky130_fd_sc_hd__or2_4
Xclkbuf_9_26_0_CLK clkbuf_9_27_0_CLK/A clkbuf_9_26_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_48109_ _48734_/A _48109_/X sky130_fd_sc_hd__buf_2
X_64155_ _61666_/A _64177_/B _64155_/C _64177_/D _64155_/Y sky130_fd_sc_hd__nand4_4
X_49089_ _49089_/A _52365_/A sky130_fd_sc_hd__buf_2
X_61367_ _61367_/A _61367_/B _61367_/C _61367_/D _61367_/Y sky130_fd_sc_hd__nand4_4
X_51120_ _51013_/A _51121_/B sky130_fd_sc_hd__buf_2
X_63106_ _58541_/A _63073_/X _63059_/X _58317_/A _63060_/X _63106_/Y
+ sky130_fd_sc_hd__o32ai_4
X_60318_ _60192_/Y _60284_/A _60259_/Y _60367_/B _60317_/Y _60318_/Y
+ sky130_fd_sc_hd__a41oi_4
X_64086_ _65044_/A _64508_/A sky130_fd_sc_hd__buf_2
X_68963_ _74119_/A _68864_/X _68891_/X _68962_/X _68963_/X sky130_fd_sc_hd__a211o_4
X_61298_ _61329_/A _61298_/B _72549_/B _61298_/Y sky130_fd_sc_hd__nand3_4
X_51051_ _51029_/A _51045_/B _51045_/C _52742_/D _51051_/X sky130_fd_sc_hd__and4_4
X_67914_ _68451_/A _67914_/X sky130_fd_sc_hd__buf_2
X_63037_ _60452_/X _63038_/A sky130_fd_sc_hd__buf_2
X_60249_ _60359_/A _60249_/X sky130_fd_sc_hd__buf_2
X_83960_ _83967_/CLK _68812_/X _80816_/D sky130_fd_sc_hd__dfxtp_4
X_68894_ _68890_/X _68893_/X _68846_/X _68894_/Y sky130_fd_sc_hd__a21oi_4
X_50002_ _86283_/Q _49986_/X _50001_/Y _50002_/Y sky130_fd_sc_hd__o21ai_4
X_82911_ _87416_/CLK _78293_/B _82911_/Q sky130_fd_sc_hd__dfxtp_4
X_67845_ _67891_/A _67845_/B _67845_/X sky130_fd_sc_hd__and2_4
X_83891_ _82299_/CLK _69869_/X _81963_/D sky130_fd_sc_hd__dfxtp_4
X_54810_ _54825_/A _54816_/B _54831_/C _53118_/D _54810_/X sky130_fd_sc_hd__and4_4
X_85630_ _85630_/CLK _85630_/D _85630_/Q sky130_fd_sc_hd__dfxtp_4
X_82842_ _82748_/CLK _79443_/X _82842_/Q sky130_fd_sc_hd__dfxtp_4
X_55790_ _55787_/X _55790_/B _55790_/X sky130_fd_sc_hd__and2_4
X_67776_ _67657_/X _67873_/A sky130_fd_sc_hd__buf_2
X_64988_ _64828_/X _85555_/Q _64829_/X _64987_/X _64988_/X sky130_fd_sc_hd__a211o_4
X_69515_ _69511_/X _69515_/B _69515_/Y sky130_fd_sc_hd__nand2_4
X_54741_ _54731_/X _47442_/Y _54741_/Y sky130_fd_sc_hd__nand2_4
X_66727_ _66722_/X _66725_/X _66726_/X _66727_/X sky130_fd_sc_hd__a21o_4
X_85561_ _85561_/CLK _85561_/D _85561_/Q sky130_fd_sc_hd__dfxtp_4
X_51953_ _51948_/Y _51951_/X _51952_/X _85918_/D sky130_fd_sc_hd__a21oi_4
X_82773_ _82774_/CLK _82773_/D _82773_/Q sky130_fd_sc_hd__dfxtp_4
X_63939_ _63933_/Y _63935_/Y _63937_/Y _63939_/D _63939_/X sky130_fd_sc_hd__and4_4
X_87300_ _87820_/CLK _43709_/X _73149_/A sky130_fd_sc_hd__dfxtp_4
X_84512_ _84518_/CLK _84512_/D _61185_/C sky130_fd_sc_hd__dfxtp_4
X_50904_ _50908_/A _50919_/B _50897_/X _51768_/D _50904_/X sky130_fd_sc_hd__and4_4
X_57460_ _57050_/A _57400_/X _57460_/Y sky130_fd_sc_hd__nand2_4
X_81724_ _80928_/CLK _81724_/D _81724_/Q sky130_fd_sc_hd__dfxtp_4
X_69446_ _69322_/A _88285_/Q _69446_/X sky130_fd_sc_hd__and2_4
X_88280_ _88288_/CLK _41090_/Y _69513_/B sky130_fd_sc_hd__dfxtp_4
X_54672_ _54400_/A _54672_/X sky130_fd_sc_hd__buf_2
X_66658_ _60150_/A _66658_/X sky130_fd_sc_hd__buf_2
X_85492_ _85492_/CLK _85492_/D _85492_/Q sky130_fd_sc_hd__dfxtp_4
X_51884_ _51875_/A _51022_/B _51884_/Y sky130_fd_sc_hd__nand2_4
X_56411_ _56436_/A _56418_/B sky130_fd_sc_hd__buf_2
X_87231_ _87748_/CLK _43858_/Y _87231_/Q sky130_fd_sc_hd__dfxtp_4
X_53623_ _85600_/Q _53556_/X _53622_/Y _53623_/Y sky130_fd_sc_hd__o21ai_4
X_65609_ _65731_/A _85877_/Q _65609_/X sky130_fd_sc_hd__and2_4
X_84443_ _84452_/CLK _84443_/D _78066_/B sky130_fd_sc_hd__dfxtp_4
X_50835_ _50833_/Y _50801_/X _50834_/X _86124_/D sky130_fd_sc_hd__a21oi_4
X_57391_ _57379_/Y _57391_/Y sky130_fd_sc_hd__inv_2
X_81655_ _81697_/CLK _81687_/Q _76453_/A sky130_fd_sc_hd__dfxtp_4
X_69377_ _87022_/Q _69239_/X _69361_/X _69376_/X _69377_/X sky130_fd_sc_hd__a211o_4
X_66589_ _87954_/Q _66529_/X _66531_/X _66588_/X _66589_/X sky130_fd_sc_hd__a211o_4
X_59130_ _59117_/A _86358_/Q _59130_/Y sky130_fd_sc_hd__nor2_4
X_80606_ _80606_/A _80606_/B _80607_/B sky130_fd_sc_hd__xnor2_4
X_56342_ _56114_/X _56337_/X _56341_/Y _85229_/D sky130_fd_sc_hd__o21ai_4
X_68328_ _68011_/X _68014_/X _68327_/X _68328_/Y sky130_fd_sc_hd__a21oi_4
X_87162_ _86935_/CLK _87162_/D _87162_/Q sky130_fd_sc_hd__dfxtp_4
X_53554_ _48287_/A _53474_/B _53492_/X _53554_/X sky130_fd_sc_hd__and3_4
X_84374_ _84438_/CLK _84374_/D _84374_/Q sky130_fd_sc_hd__dfxtp_4
X_50766_ _50771_/A _49245_/B _50766_/Y sky130_fd_sc_hd__nand2_4
X_81586_ _80912_/CLK _84186_/Q _76802_/A sky130_fd_sc_hd__dfxtp_4
X_86113_ _83685_/CLK _86113_/D _86113_/Q sky130_fd_sc_hd__dfxtp_4
X_52505_ _52503_/Y _52486_/X _52504_/Y _85809_/D sky130_fd_sc_hd__a21boi_4
X_59061_ _59061_/A _59061_/X sky130_fd_sc_hd__buf_2
X_83325_ _83325_/CLK _83325_/D _83325_/Q sky130_fd_sc_hd__dfxtp_4
X_56273_ _73359_/A _56273_/X sky130_fd_sc_hd__buf_2
X_80537_ _59102_/Y _66048_/C _80536_/Y _80537_/X sky130_fd_sc_hd__o21a_4
X_68259_ _68338_/A _68259_/X sky130_fd_sc_hd__buf_2
X_87093_ _88268_/CLK _87093_/D _87093_/Q sky130_fd_sc_hd__dfxtp_4
X_53485_ _53483_/Y _53455_/X _53484_/Y _53485_/Y sky130_fd_sc_hd__a21boi_4
X_50697_ _50682_/A _49144_/X _50697_/Y sky130_fd_sc_hd__nand2_4
X_58012_ _58070_/A _58012_/B _58012_/Y sky130_fd_sc_hd__nor2_4
X_55224_ _55224_/A _56920_/B _55224_/X sky130_fd_sc_hd__and2_4
X_86044_ _86139_/CLK _51267_/Y _64745_/B sky130_fd_sc_hd__dfxtp_4
X_52436_ _52436_/A _53953_/B _52436_/Y sky130_fd_sc_hd__nand2_4
X_40450_ _82323_/Q _40907_/B _40450_/X sky130_fd_sc_hd__or2_4
X_71270_ _53183_/B _71265_/X _71269_/Y _71270_/Y sky130_fd_sc_hd__o21ai_4
X_83256_ _86600_/CLK _72426_/Y _83256_/Q sky130_fd_sc_hd__dfxtp_4
X_80468_ _80458_/A _80458_/B _80457_/A _80456_/Y _80468_/X sky130_fd_sc_hd__o22a_4
X_82207_ _82965_/CLK _77685_/X _82207_/Q sky130_fd_sc_hd__dfxtp_4
X_70221_ _70229_/A _70229_/B _70221_/C _70229_/D _70221_/X sky130_fd_sc_hd__and4_4
X_55155_ _57326_/B _55152_/X _55168_/A _55154_/X _55155_/X sky130_fd_sc_hd__a211o_4
X_40381_ _40380_/X _40381_/X sky130_fd_sc_hd__buf_2
X_52367_ _52349_/A _52367_/B _52367_/Y sky130_fd_sc_hd__nand2_4
X_83187_ _83187_/CLK _83187_/D _70236_/C sky130_fd_sc_hd__dfxtp_4
X_80399_ _84756_/Q _84148_/Q _80401_/A sky130_fd_sc_hd__xor2_4
X_42120_ _42083_/A _42120_/X sky130_fd_sc_hd__buf_2
X_54106_ _53434_/A _54106_/B _54106_/Y sky130_fd_sc_hd__nand2_4
X_51318_ _51306_/X _46438_/A _51318_/X sky130_fd_sc_hd__and2_4
X_70152_ _70150_/Y _70151_/Y _70153_/A sky130_fd_sc_hd__nand2_4
X_82138_ _82047_/CLK _82138_/D _82094_/D sky130_fd_sc_hd__dfxtp_4
X_55086_ _85321_/Q _55072_/X _55085_/Y _55086_/Y sky130_fd_sc_hd__o21ai_4
X_59963_ _80241_/A _59787_/X _61205_/B _59962_/X _59964_/A sky130_fd_sc_hd__a2bb2o_4
X_52298_ _52271_/A _52299_/A sky130_fd_sc_hd__buf_2
X_87995_ _87995_/CLK _87995_/D _87995_/Q sky130_fd_sc_hd__dfxtp_4
X_58914_ _58904_/X _85766_/Q _58838_/X _58914_/X sky130_fd_sc_hd__o21a_4
X_42051_ _42035_/X _42049_/X _40903_/X _42050_/Y _42037_/X _42051_/Y
+ sky130_fd_sc_hd__o32ai_4
X_54037_ _54037_/A _46464_/Y _54037_/Y sky130_fd_sc_hd__nand2_4
X_51249_ _51240_/A _50744_/B _51249_/Y sky130_fd_sc_hd__nand2_4
X_86946_ _87137_/CLK _44802_/Y _86946_/Q sky130_fd_sc_hd__dfxtp_4
X_82069_ _81160_/CLK _82069_/D _82069_/Q sky130_fd_sc_hd__dfxtp_4
X_74960_ _74958_/B _81136_/D _74960_/C _74960_/Y sky130_fd_sc_hd__nand3_4
X_70083_ _69029_/Y _68823_/X _70081_/X _70082_/Y _70083_/X sky130_fd_sc_hd__a211o_4
X_59894_ _59887_/Y _59892_/Y _60165_/A _59927_/A sky130_fd_sc_hd__nand3_4
X_41002_ _41007_/A _41002_/B _41002_/X sky130_fd_sc_hd__or2_4
X_73911_ _47978_/A _73911_/B _73911_/X sky130_fd_sc_hd__xor2_4
X_58845_ _58740_/X _85451_/Q _58844_/X _58845_/Y sky130_fd_sc_hd__o21ai_4
X_74891_ _81129_/D _74891_/B _74894_/A sky130_fd_sc_hd__xor2_4
X_86877_ _86878_/CLK _45437_/Y _63030_/B sky130_fd_sc_hd__dfxtp_4
X_45810_ _45808_/Y _45734_/X _45571_/X _45809_/Y _45810_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_opt_10_CLK _84915_/CLK _84883_/CLK sky130_fd_sc_hd__clkbuf_16
X_76630_ _76595_/Y _76597_/X _76621_/X _76640_/B sky130_fd_sc_hd__a21o_4
X_73842_ _73842_/A _73649_/X _73842_/Y sky130_fd_sc_hd__nor2_4
X_85828_ _86749_/CLK _52412_/Y _85828_/Q sky130_fd_sc_hd__dfxtp_4
X_46790_ _46790_/A _46790_/Y sky130_fd_sc_hd__inv_2
X_58776_ _58776_/A _58764_/B _58776_/Y sky130_fd_sc_hd__nor2_4
X_55988_ _55686_/Y _56104_/A sky130_fd_sc_hd__buf_2
X_45741_ _45738_/Y _45632_/X _45616_/X _45740_/Y _45741_/X sky130_fd_sc_hd__a211o_4
X_57727_ _57712_/X _85728_/Q _44252_/X _57727_/X sky130_fd_sc_hd__o21a_4
X_76561_ _76559_/Y _76560_/Y _76584_/D sky130_fd_sc_hd__and2_4
X_42953_ _40331_/X _42950_/X _66598_/B _42951_/X _42953_/X sky130_fd_sc_hd__a2bb2o_4
X_54939_ _54919_/X _47788_/A _54939_/Y sky130_fd_sc_hd__nand2_4
X_73773_ _73773_/A _73599_/B _73773_/Y sky130_fd_sc_hd__nor2_4
X_85759_ _85761_/CLK _52764_/Y _85759_/Q sky130_fd_sc_hd__dfxtp_4
X_70985_ _70772_/A _70986_/A sky130_fd_sc_hd__buf_2
X_78300_ _78298_/B _78298_/A _78302_/A sky130_fd_sc_hd__nand2_4
X_75512_ _75438_/Y _75506_/X _75511_/Y _75538_/B sky130_fd_sc_hd__a21oi_4
X_41904_ _50638_/A _50523_/A sky130_fd_sc_hd__inv_2
X_48460_ _81784_/Q _48976_/B sky130_fd_sc_hd__inv_2
X_72724_ _45896_/X _72725_/A sky130_fd_sc_hd__buf_2
X_79280_ _79278_/X _79285_/B _79280_/Y sky130_fd_sc_hd__xnor2_4
X_45672_ _85071_/Q _45672_/Y sky130_fd_sc_hd__inv_2
X_57658_ _57650_/X _57655_/Y _57657_/Y _84960_/D sky130_fd_sc_hd__a21oi_4
X_76492_ _76491_/B _76491_/C _76487_/Y _76492_/Y sky130_fd_sc_hd__o21ai_4
X_42884_ _42874_/X _42875_/X _41621_/X _67294_/B _42881_/X _42885_/A
+ sky130_fd_sc_hd__o32ai_4
X_47411_ _47411_/A _53033_/B sky130_fd_sc_hd__buf_2
X_78231_ _78231_/A _78231_/B _78231_/X sky130_fd_sc_hd__xor2_4
X_44623_ _44567_/A _44623_/X sky130_fd_sc_hd__buf_2
X_56609_ _56593_/A _56609_/X sky130_fd_sc_hd__buf_2
X_75443_ _75443_/A _80955_/D _75443_/Y sky130_fd_sc_hd__nor2_4
X_87429_ _86796_/CLK _43420_/X _87429_/Q sky130_fd_sc_hd__dfxtp_4
X_41835_ _40568_/A _41835_/X sky130_fd_sc_hd__buf_2
X_48391_ _48391_/A _48391_/X sky130_fd_sc_hd__buf_2
X_72655_ _83201_/Q _72645_/X _72654_/Y _83201_/D sky130_fd_sc_hd__a21bo_4
X_57589_ _57585_/Y _57506_/X _57588_/X _84974_/D sky130_fd_sc_hd__a21oi_4
X_47342_ _47337_/Y _47317_/X _47341_/X _86645_/D sky130_fd_sc_hd__a21oi_4
X_71606_ _71690_/A _71606_/X sky130_fd_sc_hd__buf_2
X_59328_ _86662_/Q _59306_/B _59328_/Y sky130_fd_sc_hd__nor2_4
X_78162_ _78152_/A _78154_/X _78162_/C _78162_/X sky130_fd_sc_hd__and3_4
X_44554_ _44529_/A _44554_/X sky130_fd_sc_hd__buf_2
X_75374_ _75362_/A _75372_/Y _75373_/Y _75383_/A sky130_fd_sc_hd__o21a_4
X_41766_ _82887_/Q _46240_/A _41766_/X sky130_fd_sc_hd__or2_4
X_72586_ _79363_/B _72445_/X _72583_/Y _72585_/Y _72586_/Y sky130_fd_sc_hd__a2bb2oi_4
X_77113_ _77113_/A _77113_/B _77113_/Y sky130_fd_sc_hd__nand2_4
X_43505_ _43505_/A _43505_/Y sky130_fd_sc_hd__inv_2
X_74325_ _74325_/A _74325_/B _56088_/X _74325_/Y sky130_fd_sc_hd__nand3_4
X_40717_ _48192_/A _40717_/X sky130_fd_sc_hd__buf_2
X_47273_ _81820_/Q _54645_/D sky130_fd_sc_hd__inv_2
X_59259_ _59253_/X _59256_/Y _59257_/Y _59133_/X _59258_/X _59259_/X
+ sky130_fd_sc_hd__o32a_4
X_71537_ _70670_/A _71622_/D _71546_/C _71537_/Y sky130_fd_sc_hd__nor3_4
X_78093_ _78085_/A _78091_/Y _78092_/Y _78093_/Y sky130_fd_sc_hd__o21ai_4
X_44485_ _44481_/X _44482_/X _41209_/A _87085_/Q _44484_/X _44486_/A
+ sky130_fd_sc_hd__o32ai_4
X_41697_ _41697_/A _41697_/X sky130_fd_sc_hd__buf_2
X_49012_ _49022_/A _53844_/B _49012_/X sky130_fd_sc_hd__and2_4
X_46224_ _57811_/A _46224_/X sky130_fd_sc_hd__buf_2
X_77044_ _82088_/Q _77044_/B _77044_/X sky130_fd_sc_hd__xor2_4
XPHY_360 sky130_fd_sc_hd__decap_3
X_43436_ _43435_/Y _87423_/D sky130_fd_sc_hd__inv_2
X_74256_ _74022_/X _86531_/Q _74256_/X sky130_fd_sc_hd__and2_4
X_62270_ _62269_/X _62304_/A sky130_fd_sc_hd__buf_2
X_40648_ _40648_/A _40588_/B _40648_/X sky130_fd_sc_hd__or2_4
XPHY_371 sky130_fd_sc_hd__decap_3
X_71468_ _70880_/B _71435_/B _70768_/A _71476_/D _71468_/X sky130_fd_sc_hd__and4_4
XPHY_382 sky130_fd_sc_hd__decap_3
XPHY_393 sky130_fd_sc_hd__decap_3
X_61221_ _61095_/X _61179_/A _61176_/B _64456_/C _65296_/A _61221_/Y
+ sky130_fd_sc_hd__a41oi_4
X_73207_ _73206_/X _85872_/Q _73207_/X sky130_fd_sc_hd__and2_4
X_46155_ _46155_/A _46155_/X sky130_fd_sc_hd__buf_2
X_70419_ _70495_/A _71287_/C sky130_fd_sc_hd__buf_2
X_43367_ _43296_/A _43367_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_594_0_CLK clkbuf_9_297_0_CLK/X _81059_/CLK sky130_fd_sc_hd__clkbuf_1
X_74187_ _43098_/Y _56273_/X _73035_/X _74186_/Y _74187_/X sky130_fd_sc_hd__a211o_4
X_40579_ _40579_/A _40654_/B _40579_/X sky130_fd_sc_hd__or2_4
X_71399_ _70670_/A _71404_/B _71399_/C _71399_/Y sky130_fd_sc_hd__nor3_4
X_45106_ _55870_/B _45044_/X _45079_/X _45106_/X sky130_fd_sc_hd__o21a_4
X_42318_ _41878_/A _42397_/A sky130_fd_sc_hd__buf_2
X_61152_ _64523_/D _61153_/C sky130_fd_sc_hd__buf_2
X_73138_ _73239_/A _86515_/Q _73138_/X sky130_fd_sc_hd__and2_4
X_46086_ _46129_/A _46151_/B sky130_fd_sc_hd__inv_2
X_43298_ _43298_/A _43298_/Y sky130_fd_sc_hd__inv_2
X_78995_ _82647_/Q _78997_/A sky130_fd_sc_hd__inv_2
X_60103_ _60081_/A _60103_/B _60103_/C _60103_/Y sky130_fd_sc_hd__nor3_4
X_49914_ _51012_/A _49915_/A sky130_fd_sc_hd__buf_2
X_45037_ _45030_/X _45034_/Y _45036_/Y _45037_/Y sky130_fd_sc_hd__a21oi_4
X_42249_ _42259_/A _42249_/X sky130_fd_sc_hd__buf_2
X_65960_ _65300_/X _85629_/Q _65301_/X _65959_/X _65960_/X sky130_fd_sc_hd__a211o_4
X_61083_ _64361_/A _61083_/B _61083_/C _61082_/X _64367_/A sky130_fd_sc_hd__nand4_4
X_73069_ _73516_/A _73239_/A sky130_fd_sc_hd__buf_2
X_77946_ _77946_/A _77946_/Y sky130_fd_sc_hd__inv_2
X_64911_ _64908_/X _64888_/B _64910_/X _64911_/Y sky130_fd_sc_hd__nand3_4
X_60034_ _64738_/A _60034_/X sky130_fd_sc_hd__buf_2
X_49845_ _49925_/A _49851_/A sky130_fd_sc_hd__buf_2
X_65891_ _65845_/X _86178_/Q _65790_/X _65890_/X _65891_/X sky130_fd_sc_hd__a211o_4
X_77877_ _77863_/Y _77864_/Y _77851_/A _77866_/Y _77877_/X sky130_fd_sc_hd__a2bb2o_4
X_67630_ _87399_/Q _67628_/X _67581_/X _67629_/X _67630_/X sky130_fd_sc_hd__a211o_4
X_79616_ _79614_/X _79615_/X _79616_/Y sky130_fd_sc_hd__xnor2_4
X_64842_ _64870_/A _64870_/B _64841_/Y _64842_/Y sky130_fd_sc_hd__nor3_4
X_76828_ _81670_/Q _76828_/B _76828_/Y sky130_fd_sc_hd__xnor2_4
X_49776_ _46612_/A _51012_/A sky130_fd_sc_hd__buf_2
X_46988_ _46941_/A _47029_/B sky130_fd_sc_hd__buf_2
X_48727_ _48790_/A _48761_/C sky130_fd_sc_hd__buf_2
X_67561_ _67203_/X _67561_/X sky130_fd_sc_hd__buf_2
X_79547_ _79547_/A _79546_/Y _79547_/Y sky130_fd_sc_hd__nor2_4
X_45939_ _45937_/Y _45938_/X _45935_/X _45939_/Y sky130_fd_sc_hd__a21oi_4
X_64773_ _64773_/A _86459_/Q _64773_/X sky130_fd_sc_hd__and2_4
X_76759_ _76747_/Y _81357_/D sky130_fd_sc_hd__inv_2
Xclkbuf_10_532_0_CLK clkbuf_9_266_0_CLK/X _84087_/CLK sky130_fd_sc_hd__clkbuf_1
X_61985_ _61985_/A _63561_/B sky130_fd_sc_hd__buf_2
Xclkbuf_6_23_0_CLK clkbuf_6_23_0_CLK/A clkbuf_7_47_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_69300_ _69146_/A _69300_/X sky130_fd_sc_hd__buf_2
X_66512_ _60371_/X _66328_/Y _66511_/Y _66512_/Y sky130_fd_sc_hd__o21ai_4
X_63724_ _63724_/A _64192_/C sky130_fd_sc_hd__buf_2
X_48658_ _48650_/Y _48651_/X _48657_/X _48658_/Y sky130_fd_sc_hd__a21oi_4
X_60936_ _60935_/X _60937_/B sky130_fd_sc_hd__inv_2
X_67492_ _67489_/X _67491_/X _67401_/X _67492_/Y sky130_fd_sc_hd__a21oi_4
X_79478_ _79474_/Y _79496_/B _79505_/A sky130_fd_sc_hd__xor2_4
X_69231_ _68649_/A _69231_/X sky130_fd_sc_hd__buf_2
X_47609_ _47609_/A _47610_/A sky130_fd_sc_hd__inv_2
X_66443_ _66046_/A _66445_/A sky130_fd_sc_hd__buf_2
X_78429_ _78425_/Y _78369_/B _78428_/X _78429_/Y sky130_fd_sc_hd__o21ai_4
X_63655_ _63655_/A _63655_/B _63581_/X _63595_/D _63655_/X sky130_fd_sc_hd__and4_4
X_48589_ _48589_/A _52204_/A sky130_fd_sc_hd__buf_2
X_60867_ _60857_/X _60867_/Y sky130_fd_sc_hd__inv_2
XPHY_19 sky130_fd_sc_hd__decap_3
X_50620_ _50624_/A _72014_/B _50620_/Y sky130_fd_sc_hd__nand2_4
X_62606_ _62653_/A _62653_/B _62606_/C _62606_/Y sky130_fd_sc_hd__nor3_4
X_81440_ _81322_/CLK _81440_/D _76144_/B sky130_fd_sc_hd__dfxtp_4
X_69162_ _69162_/A _69162_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_547_0_CLK clkbuf_9_273_0_CLK/X _84003_/CLK sky130_fd_sc_hd__clkbuf_1
X_66374_ _66372_/Y _66343_/X _66373_/X _84135_/D sky130_fd_sc_hd__a21o_4
Xclkbuf_6_38_0_CLK clkbuf_6_39_0_CLK/A clkbuf_7_77_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_63586_ _63586_/A _63630_/B _63630_/C _63586_/Y sky130_fd_sc_hd__nor3_4
X_60798_ _63375_/A _60798_/X sky130_fd_sc_hd__buf_2
X_68113_ _82076_/D _68101_/X _68112_/X _68113_/X sky130_fd_sc_hd__a21bo_4
X_65325_ _65199_/X _86149_/Q _65224_/X _65324_/X _65325_/X sky130_fd_sc_hd__a211o_4
X_50551_ _50551_/A _50551_/X sky130_fd_sc_hd__buf_2
X_62537_ _62570_/A _63629_/B _62601_/C _62463_/X _62537_/X sky130_fd_sc_hd__and4_4
X_81371_ _81344_/CLK _76963_/Y _81371_/Q sky130_fd_sc_hd__dfxtp_4
X_69093_ _44747_/A _68570_/X _68571_/X _69092_/X _69093_/X sky130_fd_sc_hd__a211o_4
X_83110_ _82998_/CLK _74294_/X _70275_/C sky130_fd_sc_hd__dfxtp_4
X_80322_ _80320_/Y _80322_/B _80322_/X sky130_fd_sc_hd__xor2_4
X_68044_ _68044_/A _68044_/B _68044_/X sky130_fd_sc_hd__and2_4
X_53270_ _53276_/A _54446_/B _53270_/Y sky130_fd_sc_hd__nand2_4
X_65256_ _65790_/A _65256_/X sky130_fd_sc_hd__buf_2
X_84090_ _83932_/CLK _66946_/X _80914_/D sky130_fd_sc_hd__dfxtp_4
X_50482_ _86192_/Q _50387_/X _50481_/Y _50482_/Y sky130_fd_sc_hd__o21ai_4
X_62468_ _62411_/X _62412_/X _76984_/B _62468_/Y sky130_fd_sc_hd__nor3_4
X_52221_ _85865_/Q _52214_/X _52220_/Y _52221_/Y sky130_fd_sc_hd__o21ai_4
X_64207_ _64207_/A _64545_/C sky130_fd_sc_hd__buf_2
X_83041_ _82993_/CLK _83041_/D _74541_/C sky130_fd_sc_hd__dfxtp_4
X_61419_ _84850_/Q _61419_/X sky130_fd_sc_hd__buf_2
X_80253_ _84953_/Q _84201_/Q _80253_/X sky130_fd_sc_hd__xor2_4
X_65187_ _65059_/X _85547_/Q _65060_/X _65186_/X _65187_/X sky130_fd_sc_hd__a211o_4
X_62399_ _62344_/X _57672_/X _62565_/C _62355_/X _62399_/X sky130_fd_sc_hd__and4_4
X_52152_ _52152_/A _52152_/X sky130_fd_sc_hd__buf_2
X_64138_ _60034_/X _64187_/A sky130_fd_sc_hd__buf_2
X_80184_ _80176_/A _80175_/X _80183_/Y _80184_/Y sky130_fd_sc_hd__a21boi_4
X_69995_ _69625_/X _69628_/X _69994_/X _69995_/X sky130_fd_sc_hd__a21o_4
X_51103_ _51112_/A _52794_/B _51103_/Y sky130_fd_sc_hd__nand2_4
X_86800_ _87073_/CLK _46038_/Y _86800_/Q sky130_fd_sc_hd__dfxtp_4
X_52083_ _52083_/A _50381_/B _52083_/Y sky130_fd_sc_hd__nand2_4
X_56960_ _56774_/A _56960_/X sky130_fd_sc_hd__buf_2
X_68946_ _68942_/X _68945_/X _68922_/X _68946_/X sky130_fd_sc_hd__a21o_4
X_64069_ _61570_/B _64161_/B _64150_/C _64161_/D _64069_/Y sky130_fd_sc_hd__nand4_4
X_87780_ _87782_/CLK _42668_/Y _87780_/Q sky130_fd_sc_hd__dfxtp_4
X_84992_ _85920_/CLK _84992_/D _84992_/Q sky130_fd_sc_hd__dfxtp_4
X_51034_ _51141_/A _51045_/C sky130_fd_sc_hd__buf_2
X_55911_ _85208_/Q _55617_/A _55627_/X _55910_/X _55911_/X sky130_fd_sc_hd__a211o_4
X_86731_ _86733_/CLK _86731_/D _86731_/Q sky130_fd_sc_hd__dfxtp_4
X_83943_ _81351_/CLK _69175_/X _83943_/Q sky130_fd_sc_hd__dfxtp_4
X_56891_ _55662_/Y _56889_/X _56890_/Y _56892_/B sky130_fd_sc_hd__a21oi_4
X_68877_ _87083_/Q _68832_/X _68875_/X _68876_/X _68877_/X sky130_fd_sc_hd__a211o_4
X_58630_ _58627_/Y _58629_/Y _58003_/X _58630_/X sky130_fd_sc_hd__a21o_4
X_55842_ _83025_/Q _55572_/X _55532_/X _55841_/X _55842_/X sky130_fd_sc_hd__a211o_4
X_67828_ _67824_/X _67827_/X _67637_/X _67828_/Y sky130_fd_sc_hd__a21oi_4
X_86662_ _86665_/CLK _47182_/Y _86662_/Q sky130_fd_sc_hd__dfxtp_4
X_83874_ _82558_/CLK _70008_/X _83874_/Q sky130_fd_sc_hd__dfxtp_4
X_88401_ _87883_/CLK _40377_/Y _88401_/Q sky130_fd_sc_hd__dfxtp_4
X_85613_ _85601_/CLK _85613_/D _85613_/Q sky130_fd_sc_hd__dfxtp_4
X_58561_ _58984_/A _58973_/B sky130_fd_sc_hd__buf_2
X_82825_ _83238_/CLK _79263_/X _82825_/Q sky130_fd_sc_hd__dfxtp_4
X_55773_ _56117_/A _56117_/B _56117_/C _55773_/D _55801_/A sky130_fd_sc_hd__and4_4
X_67759_ _67496_/X _67746_/Y _67747_/X _67758_/Y _67759_/X sky130_fd_sc_hd__a211o_4
X_86593_ _83161_/CLK _86593_/D _65908_/B sky130_fd_sc_hd__dfxtp_4
X_52985_ _52903_/X _52999_/A sky130_fd_sc_hd__buf_2
X_57512_ _57510_/Y _46576_/X _57511_/Y _84989_/D sky130_fd_sc_hd__a21boi_4
X_88332_ _84970_/CLK _88332_/D _88332_/Q sky130_fd_sc_hd__dfxtp_4
X_54724_ _85389_/Q _54703_/X _54723_/Y _54724_/Y sky130_fd_sc_hd__o21ai_4
X_85544_ _86145_/CLK _85544_/D _85544_/Q sky130_fd_sc_hd__dfxtp_4
X_51936_ _52407_/A _51941_/A sky130_fd_sc_hd__buf_2
X_70770_ _52843_/B _70761_/X _70769_/Y _70770_/Y sky130_fd_sc_hd__o21ai_4
X_82756_ _82768_/CLK _82756_/D _82948_/D sky130_fd_sc_hd__dfxtp_4
X_58492_ _58517_/A _58492_/X sky130_fd_sc_hd__buf_2
X_81707_ _81514_/CLK _81707_/D _41228_/A sky130_fd_sc_hd__dfxtp_4
X_57443_ _85003_/Q _57463_/B _57443_/X sky130_fd_sc_hd__or2_4
X_88263_ _88263_/CLK _41176_/Y _68686_/B sky130_fd_sc_hd__dfxtp_4
X_69429_ _69426_/X _69428_/X _69346_/X _69429_/X sky130_fd_sc_hd__a21o_4
X_54655_ _85402_/Q _54648_/X _54654_/Y _54655_/Y sky130_fd_sc_hd__o21ai_4
X_85475_ _84926_/CLK _85475_/D _85475_/Q sky130_fd_sc_hd__dfxtp_4
X_51867_ _51853_/A _51003_/B _51867_/Y sky130_fd_sc_hd__nand2_4
X_82687_ _84111_/CLK _82687_/D _82687_/Q sky130_fd_sc_hd__dfxtp_4
X_87214_ _86934_/CLK _87214_/D _67453_/B sky130_fd_sc_hd__dfxtp_4
X_41620_ _41533_/X _82307_/Q _41619_/X _41620_/X sky130_fd_sc_hd__o21a_4
X_53606_ _53601_/A _48141_/A _53606_/Y sky130_fd_sc_hd__nand2_4
X_72440_ _72419_/X _85350_/Q _72439_/X _72440_/Y sky130_fd_sc_hd__o21ai_4
X_84426_ _84426_/CLK _62192_/Y _78049_/B sky130_fd_sc_hd__dfxtp_4
X_50818_ _50595_/A _50991_/A sky130_fd_sc_hd__buf_2
X_57374_ _72910_/A _73040_/A sky130_fd_sc_hd__buf_2
X_81638_ _80912_/CLK _81670_/Q _81638_/Q sky130_fd_sc_hd__dfxtp_4
X_88194_ _87116_/CLK _88194_/D _88194_/Q sky130_fd_sc_hd__dfxtp_4
X_54586_ _54583_/Y _54584_/X _54585_/X _54586_/Y sky130_fd_sc_hd__a21oi_4
X_51798_ _51794_/A _51794_/B _51794_/C _46707_/X _51798_/X sky130_fd_sc_hd__and4_4
Xclkbuf_8_6_0_CLK clkbuf_8_7_0_CLK/A clkbuf_8_6_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_59113_ _58864_/X _59110_/Y _59112_/Y _58943_/X _58868_/X _59113_/X
+ sky130_fd_sc_hd__o32a_4
X_56325_ _56351_/A _56335_/B sky130_fd_sc_hd__buf_2
X_87145_ _86920_/CLK _44367_/X _87145_/Q sky130_fd_sc_hd__dfxtp_4
X_53537_ _53982_/A _53537_/X sky130_fd_sc_hd__buf_2
X_41551_ _41548_/X _82320_/Q _41550_/X _41552_/A sky130_fd_sc_hd__o21ai_4
X_72371_ _83260_/Q _72371_/Y sky130_fd_sc_hd__inv_2
X_84357_ _84360_/CLK _63058_/X _79467_/A sky130_fd_sc_hd__dfxtp_4
X_50749_ _86141_/Q _50727_/X _50748_/Y _50749_/Y sky130_fd_sc_hd__o21ai_4
X_81569_ _83940_/CLK _76958_/Y _81525_/D sky130_fd_sc_hd__dfxtp_4
X_74110_ _74106_/X _85610_/Q _74107_/X _74109_/X _74110_/X sky130_fd_sc_hd__a211o_4
X_40502_ _40477_/X _40488_/X _40501_/X _88381_/Q _40492_/X _40502_/Y
+ sky130_fd_sc_hd__o32ai_4
X_59044_ _59029_/A _59044_/B _59044_/Y sky130_fd_sc_hd__nor2_4
X_83308_ _85547_/CLK _83308_/D _83308_/Q sky130_fd_sc_hd__dfxtp_4
X_71322_ _48310_/B _71320_/X _71321_/Y _83537_/D sky130_fd_sc_hd__o21ai_4
X_44270_ _72908_/A _44270_/X sky130_fd_sc_hd__buf_2
X_56256_ _56263_/A _56253_/B _85257_/Q _56256_/Y sky130_fd_sc_hd__nand3_4
X_75090_ _75091_/A _75102_/A _75091_/B _75090_/X sky130_fd_sc_hd__a21o_4
X_87076_ _88245_/CLK _44505_/X _87076_/Q sky130_fd_sc_hd__dfxtp_4
X_41482_ _41482_/A _41523_/B sky130_fd_sc_hd__buf_2
X_53468_ _53468_/A _47863_/Y _53468_/Y sky130_fd_sc_hd__nand2_4
X_84288_ _84671_/CLK _63898_/Y _63897_/C sky130_fd_sc_hd__dfxtp_4
X_43221_ _43221_/A _43221_/Y sky130_fd_sc_hd__inv_2
X_55207_ _55207_/A _55208_/B sky130_fd_sc_hd__inv_2
X_74041_ _74016_/X _85613_/Q _73903_/X _74040_/X _74041_/X sky130_fd_sc_hd__a211o_4
X_86027_ _86029_/CLK _86027_/D _86027_/Q sky130_fd_sc_hd__dfxtp_4
X_40433_ _57491_/A _40364_/X _40432_/X _88392_/Q _40375_/X _40434_/A
+ sky130_fd_sc_hd__o32ai_4
X_52419_ _85826_/Q _52397_/X _52418_/Y _52419_/Y sky130_fd_sc_hd__o21ai_4
X_71253_ _51954_/B _71239_/X _71252_/Y _71253_/Y sky130_fd_sc_hd__o21ai_4
X_83239_ _84487_/CLK _83239_/D _79493_/B sky130_fd_sc_hd__dfxtp_4
X_56187_ _56186_/Y _56255_/A sky130_fd_sc_hd__buf_2
X_53399_ _53386_/A _54578_/B _53399_/Y sky130_fd_sc_hd__nand2_4
X_70204_ _70233_/A _70204_/X sky130_fd_sc_hd__buf_2
X_43152_ _87556_/Q _43152_/Y sky130_fd_sc_hd__inv_2
X_55138_ _55138_/A _55138_/X sky130_fd_sc_hd__buf_2
X_40364_ _40363_/X _40364_/X sky130_fd_sc_hd__buf_2
X_71184_ _50466_/B _71164_/Y _71183_/Y _71184_/Y sky130_fd_sc_hd__o21ai_4
X_42103_ _51719_/A _42103_/X sky130_fd_sc_hd__buf_2
X_77800_ _77786_/X _77787_/A _77800_/X sky130_fd_sc_hd__and2_4
X_70135_ _83512_/Q _83160_/Q _83509_/Q _83157_/Q _70139_/A sky130_fd_sc_hd__a22oi_4
X_47960_ _73864_/A _50293_/B sky130_fd_sc_hd__buf_2
X_43083_ _43072_/X _43075_/X _40707_/X _74053_/A _43080_/X _43083_/Y
+ sky130_fd_sc_hd__o32ai_4
X_55069_ _46614_/X _55083_/A sky130_fd_sc_hd__buf_2
X_59946_ _59945_/Y _59951_/C sky130_fd_sc_hd__buf_2
X_78780_ _78780_/A _78773_/X _78779_/Y _78783_/A sky130_fd_sc_hd__nand3_4
X_75992_ _81707_/D _75991_/B _75992_/Y sky130_fd_sc_hd__nand2_4
X_87978_ _88158_/CLK _87978_/D _87978_/Q sky130_fd_sc_hd__dfxtp_4
X_46911_ _46911_/A _52744_/B sky130_fd_sc_hd__inv_2
X_42034_ _42034_/A _42034_/Y sky130_fd_sc_hd__inv_2
X_77731_ _82258_/Q _77731_/Y sky130_fd_sc_hd__inv_2
X_74943_ _74933_/Y _74943_/B _74947_/A sky130_fd_sc_hd__nand2_4
X_70066_ _83859_/Q _70048_/X _70065_/Y _70066_/X sky130_fd_sc_hd__a21bo_4
X_86929_ _87144_/CLK _86929_/D _67679_/B sky130_fd_sc_hd__dfxtp_4
X_47891_ _47855_/A _50260_/B _47891_/Y sky130_fd_sc_hd__nand2_4
X_59877_ _59876_/X _59877_/X sky130_fd_sc_hd__buf_2
X_49630_ _49625_/A _49614_/X _49629_/X _52846_/D _49630_/X sky130_fd_sc_hd__and4_4
X_46842_ _46817_/A _51016_/B _46842_/Y sky130_fd_sc_hd__nand2_4
X_58828_ _58918_/A _58828_/X sky130_fd_sc_hd__buf_2
X_77662_ _77661_/X _77662_/Y sky130_fd_sc_hd__inv_2
X_74874_ _74874_/A _74874_/B _74874_/X sky130_fd_sc_hd__xor2_4
X_79401_ _79418_/B _79401_/B _82838_/D sky130_fd_sc_hd__xor2_4
X_76613_ _76613_/A _76613_/B _81343_/D sky130_fd_sc_hd__nor2_4
X_49561_ _49561_/A _49561_/B _49548_/X _52775_/D _49561_/X sky130_fd_sc_hd__and4_4
X_73825_ _68645_/B _73801_/X _73704_/X _73825_/Y sky130_fd_sc_hd__o21ai_4
X_46773_ _46915_/A _46784_/A sky130_fd_sc_hd__buf_2
X_58759_ _58714_/X _85778_/Q _58716_/X _58759_/X sky130_fd_sc_hd__o21a_4
X_77593_ _77592_/X _77593_/Y sky130_fd_sc_hd__inv_2
X_43985_ _44186_/A _43954_/X _43945_/Y _43984_/Y _43985_/X sky130_fd_sc_hd__a211o_4
X_48512_ _48506_/Y _48459_/X _48511_/X _86516_/D sky130_fd_sc_hd__a21oi_4
X_79332_ _79346_/A _79346_/B _79332_/X sky130_fd_sc_hd__xor2_4
X_45724_ _85036_/Q _45675_/X _45723_/X _45724_/Y sky130_fd_sc_hd__o21ai_4
X_76544_ _76526_/X _76544_/Y sky130_fd_sc_hd__inv_2
X_42936_ _42936_/A _42936_/Y sky130_fd_sc_hd__inv_2
X_49492_ _86377_/Q _49470_/X _49491_/Y _49492_/Y sky130_fd_sc_hd__o21ai_4
X_61770_ _61770_/A _61770_/B _63396_/B _61770_/D _61770_/X sky130_fd_sc_hd__and4_4
X_73756_ _44691_/Y _73728_/X _73755_/Y _73767_/C sky130_fd_sc_hd__a21o_4
X_70968_ _50777_/B _70961_/X _70967_/Y _70968_/Y sky130_fd_sc_hd__o21ai_4
X_48443_ _48436_/Y _48383_/X _48442_/X _48443_/Y sky130_fd_sc_hd__a21oi_4
X_60721_ _63413_/A _63672_/C sky130_fd_sc_hd__buf_2
X_72707_ _70251_/C _72702_/X _72706_/Y _72707_/X sky130_fd_sc_hd__a21bo_4
X_79263_ _79263_/A _79263_/B _79263_/X sky130_fd_sc_hd__xor2_4
X_45655_ _45652_/X _45654_/Y _45561_/X _45655_/Y sky130_fd_sc_hd__a21oi_4
X_76475_ _76471_/Y _76473_/Y _76474_/A _76479_/C sky130_fd_sc_hd__o21ai_4
X_42867_ _42832_/A _42867_/X sky130_fd_sc_hd__buf_2
X_73687_ _73609_/X _85628_/Q _73661_/X _73686_/X _73687_/X sky130_fd_sc_hd__a211o_4
X_70899_ _70871_/A _70903_/B _70899_/C _70899_/D _70899_/Y sky130_fd_sc_hd__nand4_4
X_78214_ _78220_/B _78220_/C _78214_/Y sky130_fd_sc_hd__nand2_4
X_44606_ _44588_/X _44589_/X _40950_/A _87037_/Q _44590_/X _44606_/Y
+ sky130_fd_sc_hd__o32ai_4
X_63440_ _63375_/A _63463_/A sky130_fd_sc_hd__buf_2
X_75426_ _75426_/A _75427_/C sky130_fd_sc_hd__inv_2
X_41818_ _41818_/A _41818_/Y sky130_fd_sc_hd__inv_2
X_48374_ _48891_/B _48449_/B _48374_/Y sky130_fd_sc_hd__nand2_4
X_60652_ _60652_/A _60652_/X sky130_fd_sc_hd__buf_2
X_72638_ _70176_/C _72631_/X _72637_/Y _83208_/D sky130_fd_sc_hd__a21bo_4
X_79194_ _79186_/Y _79180_/Y _79181_/Y _79207_/B sky130_fd_sc_hd__a21boi_4
X_45586_ _45584_/Y _45570_/X _45520_/X _45585_/Y _45586_/X sky130_fd_sc_hd__a211o_4
X_42798_ _42797_/Y _42798_/Y sky130_fd_sc_hd__inv_2
X_47325_ _47287_/X _52986_/B _47325_/Y sky130_fd_sc_hd__nand2_4
X_78145_ _78145_/A _82860_/D _78152_/A sky130_fd_sc_hd__xor2_4
X_44537_ _72973_/A _44537_/Y sky130_fd_sc_hd__inv_2
X_75357_ _75355_/X _75357_/B _75357_/Y sky130_fd_sc_hd__xnor2_4
X_63371_ _63371_/A _63372_/A sky130_fd_sc_hd__buf_2
X_41749_ _41748_/Y _41749_/X sky130_fd_sc_hd__buf_2
X_60583_ _60583_/A _60602_/B _63280_/C _60583_/Y sky130_fd_sc_hd__nor3_4
X_72569_ _72569_/A _57896_/A _72569_/C _72569_/Y sky130_fd_sc_hd__nand3_4
X_65110_ _65065_/X _86734_/Q _65108_/X _65109_/X _65110_/X sky130_fd_sc_hd__a211o_4
X_62322_ _62362_/A _62317_/Y _62322_/C _62321_/Y _62322_/Y sky130_fd_sc_hd__nand4_4
X_74308_ _74302_/X _74310_/B _56044_/X _74308_/Y sky130_fd_sc_hd__nand3_4
X_47256_ _54634_/D _52942_/D sky130_fd_sc_hd__buf_2
X_66090_ _66081_/Y _66089_/Y _66090_/Y sky130_fd_sc_hd__nand2_4
X_78076_ _60717_/C _78076_/B _78076_/X sky130_fd_sc_hd__xor2_4
X_44468_ _41161_/A _44464_/X _87094_/Q _44466_/X _44468_/X sky130_fd_sc_hd__a2bb2o_4
X_75288_ _75288_/A _80945_/D _75288_/Y sky130_fd_sc_hd__nor2_4
X_46207_ _46222_/A _46207_/B _46162_/C _46207_/Y sky130_fd_sc_hd__nand3_4
X_65041_ _64934_/X _83297_/Q _64991_/X _65040_/X _65041_/X sky130_fd_sc_hd__a211o_4
XPHY_190 sky130_fd_sc_hd__decap_3
X_77027_ _77034_/B _77026_/Y _77028_/B sky130_fd_sc_hd__xor2_4
X_43419_ _41525_/X _43412_/X _87430_/Q _43413_/X _43419_/X sky130_fd_sc_hd__a2bb2o_4
X_62253_ _62033_/A _62253_/X sky130_fd_sc_hd__buf_2
X_74239_ _74239_/A _74239_/B _74239_/Y sky130_fd_sc_hd__nand2_4
X_47187_ _47140_/A _47210_/C sky130_fd_sc_hd__buf_2
X_44399_ _44381_/X _44382_/X _41498_/X _87128_/Q _44383_/X _44400_/A
+ sky130_fd_sc_hd__o32ai_4
X_61204_ _61190_/X _61156_/X _61272_/B _61202_/Y _61203_/Y _84508_/D
+ sky130_fd_sc_hd__a41oi_4
X_46138_ _46138_/A _46119_/A _43012_/B _46138_/Y sky130_fd_sc_hd__nand3_4
X_62184_ _63713_/A _59628_/A _59763_/A _62188_/B sky130_fd_sc_hd__a21o_4
X_68800_ _69478_/A _68800_/X sky130_fd_sc_hd__buf_2
X_61135_ _64546_/A _64225_/B _61135_/X sky130_fd_sc_hd__and2_4
X_46069_ _46067_/X _46054_/X _41573_/X _86784_/Q _46068_/X _46070_/A
+ sky130_fd_sc_hd__o32ai_4
X_69780_ _69766_/A _69780_/B _69780_/Y sky130_fd_sc_hd__nor2_4
X_66992_ _66947_/X _66980_/Y _66910_/X _66991_/Y _66992_/X sky130_fd_sc_hd__a211o_4
X_78978_ _78976_/Y _78978_/B _78986_/B sky130_fd_sc_hd__xor2_4
X_68731_ _69371_/A _68731_/X sky130_fd_sc_hd__buf_2
X_65943_ _65916_/A _65970_/B _84167_/Q _65943_/X sky130_fd_sc_hd__and3_4
X_77929_ _77916_/A _77923_/A _77929_/X sky130_fd_sc_hd__and2_4
X_61066_ _59622_/A _61066_/B _60641_/A _61066_/Y sky130_fd_sc_hd__nor3_4
X_60017_ _62336_/A _62623_/A sky130_fd_sc_hd__buf_2
X_49828_ _49827_/X _53041_/B _49828_/Y sky130_fd_sc_hd__nand2_4
X_80940_ _80804_/CLK _80984_/Q _74920_/A sky130_fd_sc_hd__dfxtp_4
X_68662_ _68656_/X _68659_/X _68661_/X _68662_/Y sky130_fd_sc_hd__a21oi_4
X_65874_ _65702_/A _85859_/Q _65874_/X sky130_fd_sc_hd__and2_4
Xclkbuf_10_471_0_CLK clkbuf_9_235_0_CLK/X _85767_/CLK sky130_fd_sc_hd__clkbuf_1
X_67613_ _67569_/X _67613_/B _67613_/X sky130_fd_sc_hd__and2_4
X_64825_ _64822_/X _64712_/B _64824_/X _64825_/Y sky130_fd_sc_hd__nand3_4
X_49759_ _49787_/A _49759_/X sky130_fd_sc_hd__buf_2
X_80871_ _80746_/CLK _75617_/B _80871_/Q sky130_fd_sc_hd__dfxtp_4
X_68593_ _73773_/A _68069_/X _68070_/X _68592_/Y _68593_/X sky130_fd_sc_hd__a211o_4
X_82610_ _82610_/CLK _78958_/B _82578_/D sky130_fd_sc_hd__dfxtp_4
X_67544_ _84065_/Q _67449_/X _67543_/X _84065_/D sky130_fd_sc_hd__a21bo_4
X_52770_ _52770_/A _52775_/B sky130_fd_sc_hd__buf_2
X_64756_ _64722_/X _85564_/Q _64724_/X _64755_/X _64756_/X sky130_fd_sc_hd__a211o_4
X_83590_ _86523_/CLK _83590_/D _83590_/Q sky130_fd_sc_hd__dfxtp_4
X_61968_ _61509_/B _61953_/B _61953_/C _61937_/X _61968_/Y sky130_fd_sc_hd__nand4_4
X_51721_ _52605_/A _51721_/X sky130_fd_sc_hd__buf_2
X_63707_ _61682_/B _63426_/A _63705_/X _63706_/X _63707_/X sky130_fd_sc_hd__a211o_4
X_82541_ _82541_/CLK _82541_/D _79051_/B sky130_fd_sc_hd__dfxtp_4
X_60919_ _60855_/X _60920_/A sky130_fd_sc_hd__buf_2
X_67475_ _87917_/Q _67473_/X _67405_/X _67474_/X _67475_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_486_0_CLK clkbuf_9_243_0_CLK/X _84802_/CLK sky130_fd_sc_hd__clkbuf_1
X_64687_ _64561_/X _64675_/Y _64686_/Y _64687_/Y sky130_fd_sc_hd__o21ai_4
X_61899_ _61960_/A _61960_/B _78070_/B _61899_/Y sky130_fd_sc_hd__nor3_4
X_69214_ _69146_/X _69109_/X _69211_/Y _69213_/Y _69214_/X sky130_fd_sc_hd__a211o_4
X_54440_ _54435_/A _54440_/B _54429_/C _46916_/Y _54440_/X sky130_fd_sc_hd__and4_4
X_66426_ _66426_/A _66397_/X _66426_/C _66426_/Y sky130_fd_sc_hd__nand3_4
X_85260_ _85192_/CLK _56249_/Y _85260_/Q sky130_fd_sc_hd__dfxtp_4
X_51652_ _51650_/Y _51639_/X _51651_/X _51652_/Y sky130_fd_sc_hd__a21oi_4
X_63638_ _58400_/A _63648_/B _63638_/Y sky130_fd_sc_hd__nor2_4
X_82472_ _81198_/CLK _78401_/X _82472_/Q sky130_fd_sc_hd__dfxtp_4
X_84211_ _85315_/CLK _84211_/D _84211_/Q sky130_fd_sc_hd__dfxtp_4
X_50603_ _50597_/A _48963_/X _50603_/Y sky130_fd_sc_hd__nand2_4
X_81423_ _81749_/CLK _81423_/D _76021_/B sky130_fd_sc_hd__dfxtp_4
X_69145_ _83945_/Q _69066_/X _69144_/X _83945_/D sky130_fd_sc_hd__a21bo_4
X_54371_ _54399_/A _54395_/A sky130_fd_sc_hd__buf_2
X_66357_ _65894_/X _66367_/B _65897_/X _66357_/Y sky130_fd_sc_hd__nand3_4
X_85191_ _85190_/CLK _85191_/D _56444_/C sky130_fd_sc_hd__dfxtp_4
X_51583_ _85983_/Q _51566_/X _51582_/Y _51583_/Y sky130_fd_sc_hd__o21ai_4
X_63569_ _63546_/A _58474_/A _63520_/C _63546_/D _63569_/X sky130_fd_sc_hd__and4_4
X_56110_ _56131_/A _56115_/B _55817_/B _56110_/Y sky130_fd_sc_hd__nand3_4
X_53322_ _53330_/A _53330_/B _53302_/X _52805_/D _53322_/X sky130_fd_sc_hd__and4_4
X_65308_ _57947_/A _65308_/X sky130_fd_sc_hd__buf_2
X_84142_ _84231_/CLK _84142_/D _84142_/Q sky130_fd_sc_hd__dfxtp_4
X_50534_ _50534_/A _50541_/A sky130_fd_sc_hd__buf_2
X_57090_ _73186_/A _73227_/A sky130_fd_sc_hd__buf_2
X_81354_ _81322_/CLK _81354_/D _76274_/A sky130_fd_sc_hd__dfxtp_4
X_69076_ _69134_/A _69076_/B _69076_/X sky130_fd_sc_hd__and2_4
X_66288_ _58805_/A _74177_/B _66288_/X sky130_fd_sc_hd__and2_4
X_56041_ _56023_/A _56052_/B _56041_/C _56041_/Y sky130_fd_sc_hd__nand3_4
X_80305_ _80298_/A _80292_/A _80292_/B _80319_/B sky130_fd_sc_hd__a21boi_4
X_68027_ _68027_/A _68027_/B _68027_/Y sky130_fd_sc_hd__nand2_4
X_53253_ _53243_/X _51747_/A _53266_/C _53253_/D _53253_/X sky130_fd_sc_hd__and4_4
X_65239_ _64991_/A _65239_/X sky130_fd_sc_hd__buf_2
X_84073_ _81473_/CLK _67353_/X _81505_/D sky130_fd_sc_hd__dfxtp_4
X_50465_ _50534_/A _50465_/X sky130_fd_sc_hd__buf_2
X_81285_ _81282_/CLK _76973_/X _81285_/Q sky130_fd_sc_hd__dfxtp_4
X_52204_ _52204_/A _52198_/X _52218_/C _52204_/X sky130_fd_sc_hd__and3_4
X_83024_ _83025_/CLK _74590_/Y _45168_/A sky130_fd_sc_hd__dfxtp_4
X_87901_ _87644_/CLK _87901_/D _87901_/Q sky130_fd_sc_hd__dfxtp_4
X_80236_ _80228_/A _80227_/Y _80235_/X _80236_/Y sky130_fd_sc_hd__o21ai_4
X_53184_ _85681_/Q _53172_/X _53183_/Y _53184_/Y sky130_fd_sc_hd__o21ai_4
X_50396_ _53620_/A _50331_/B _50338_/X _50396_/X sky130_fd_sc_hd__and3_4
Xclkbuf_10_424_0_CLK clkbuf_9_212_0_CLK/X _82797_/CLK sky130_fd_sc_hd__clkbuf_1
X_59800_ _59687_/C _59688_/X _59797_/Y _59798_/Y _59799_/Y _59800_/Y
+ sky130_fd_sc_hd__a41oi_4
X_52135_ _52135_/A _52135_/B _52156_/C _52135_/X sky130_fd_sc_hd__and3_4
X_87832_ _88086_/CLK _42531_/Y _74184_/A sky130_fd_sc_hd__dfxtp_4
X_80167_ _80167_/A _80166_/X _80167_/Y sky130_fd_sc_hd__xnor2_4
X_57992_ _86638_/Q _57954_/X _57992_/Y sky130_fd_sc_hd__nor2_4
X_69978_ _68369_/X _68372_/X _69925_/X _69978_/Y sky130_fd_sc_hd__a21oi_4
X_59731_ _59687_/A _59731_/Y sky130_fd_sc_hd__inv_2
X_52066_ _52462_/A _52066_/X sky130_fd_sc_hd__buf_2
X_56943_ _56940_/Y _56943_/X sky130_fd_sc_hd__buf_2
X_68929_ _68300_/X _68929_/X sky130_fd_sc_hd__buf_2
X_87763_ _87520_/CLK _42702_/Y _68343_/B sky130_fd_sc_hd__dfxtp_4
X_84975_ _83544_/CLK _57583_/Y _84975_/Q sky130_fd_sc_hd__dfxtp_4
X_80098_ _80098_/A _80098_/B _80098_/X sky130_fd_sc_hd__xor2_4
X_51017_ _86089_/Q _50992_/X _51016_/Y _51017_/Y sky130_fd_sc_hd__o21ai_4
X_86714_ _86711_/CLK _86714_/D _58660_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_439_0_CLK clkbuf_9_219_0_CLK/X _85354_/CLK sky130_fd_sc_hd__clkbuf_1
X_71940_ _70368_/X _71001_/C _71940_/C _71945_/D _71940_/Y sky130_fd_sc_hd__nand4_4
X_59662_ _59805_/A _59662_/B _59662_/C _59681_/A sky130_fd_sc_hd__and3_4
X_83926_ _83926_/CLK _83926_/D _81390_/D sky130_fd_sc_hd__dfxtp_4
X_56874_ _56873_/X _56774_/C _56874_/X sky130_fd_sc_hd__and2_4
Xclkbuf_1_0_0_CLK clkbuf_0_CLK/X clkbuf_1_0_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_87694_ _87950_/CLK _42834_/X _66689_/B sky130_fd_sc_hd__dfxtp_4
X_58613_ _58687_/A _58613_/B _58613_/Y sky130_fd_sc_hd__nor2_4
X_55825_ _55822_/X _55824_/X _44111_/X _55825_/X sky130_fd_sc_hd__a21o_4
X_86645_ _86005_/CLK _86645_/D _86645_/Q sky130_fd_sc_hd__dfxtp_4
X_71871_ _71870_/Y _71871_/X sky130_fd_sc_hd__buf_2
X_59593_ _59546_/A _43998_/A _59543_/A _59593_/X sky130_fd_sc_hd__and3_4
X_83857_ _82536_/CLK _83857_/D _82537_/D sky130_fd_sc_hd__dfxtp_4
X_73610_ _73638_/A _65935_/B _73610_/X sky130_fd_sc_hd__and2_4
X_70822_ _71219_/A _70954_/B _70703_/X _70822_/Y sky130_fd_sc_hd__nand3_4
X_58544_ _58543_/Y _58557_/B _58544_/Y sky130_fd_sc_hd__nand2_4
X_82808_ _82740_/CLK _82840_/Q _82808_/Q sky130_fd_sc_hd__dfxtp_4
X_43770_ _43752_/A _43770_/X sky130_fd_sc_hd__buf_2
X_55756_ _55192_/A _55756_/B _55756_/X sky130_fd_sc_hd__and2_4
X_74590_ _45169_/A _74582_/X _74589_/X _74590_/Y sky130_fd_sc_hd__o21ai_4
X_86576_ _86576_/CLK _86576_/D _66155_/B sky130_fd_sc_hd__dfxtp_4
X_40982_ _40982_/A _40982_/X sky130_fd_sc_hd__buf_2
X_52968_ _52966_/Y _52946_/X _52967_/X _85722_/D sky130_fd_sc_hd__a21oi_4
X_83788_ _81620_/CLK _83788_/D _74760_/A sky130_fd_sc_hd__dfxtp_4
X_42721_ _42720_/X _42721_/X sky130_fd_sc_hd__buf_2
X_88315_ _88056_/CLK _88315_/D _69888_/B sky130_fd_sc_hd__dfxtp_4
X_54707_ _54699_/X _54707_/B _54721_/C _47379_/A _54707_/X sky130_fd_sc_hd__and4_4
X_73541_ _72722_/X _83050_/Q _73406_/X _73540_/X _73542_/B sky130_fd_sc_hd__a211o_4
X_85527_ _85527_/CLK _53994_/Y _85527_/Q sky130_fd_sc_hd__dfxtp_4
X_51919_ _51914_/A _51898_/B _51919_/C _52746_/D _51919_/X sky130_fd_sc_hd__and4_4
X_70753_ _70753_/A _70724_/A _70753_/Y sky130_fd_sc_hd__nand2_4
X_58475_ _58467_/X _58472_/Y _58474_/Y _84840_/D sky130_fd_sc_hd__a21oi_4
X_82739_ _84177_/CLK _66435_/A _78965_/A sky130_fd_sc_hd__dfxtp_4
X_55687_ _55686_/Y _56169_/A sky130_fd_sc_hd__buf_2
X_52899_ _52845_/A _52900_/C sky130_fd_sc_hd__buf_2
X_57426_ _57275_/X _57003_/B _57425_/X _57426_/X sky130_fd_sc_hd__o21a_4
X_45440_ _45440_/A _44892_/X _45440_/Y sky130_fd_sc_hd__nor2_4
X_76260_ _81258_/Q _81514_/D _76260_/X sky130_fd_sc_hd__xor2_4
X_88246_ _88247_/CLK _41273_/X _88246_/Q sky130_fd_sc_hd__dfxtp_4
X_42652_ _42651_/X _42652_/X sky130_fd_sc_hd__buf_2
X_73472_ _73284_/A _73472_/X sky130_fd_sc_hd__buf_2
X_54638_ _54558_/A _54638_/X sky130_fd_sc_hd__buf_2
X_85458_ _85459_/CLK _85458_/D _85458_/Q sky130_fd_sc_hd__dfxtp_4
X_70684_ _71863_/A _71411_/A sky130_fd_sc_hd__buf_2
X_75211_ _80779_/Q _81035_/D _80747_/D sky130_fd_sc_hd__xor2_4
X_41603_ _40365_/X _41603_/X sky130_fd_sc_hd__buf_2
X_72423_ _72389_/X _85672_/Q _72422_/X _72423_/X sky130_fd_sc_hd__o21a_4
X_84409_ _84409_/CLK _84409_/D _76985_/B sky130_fd_sc_hd__dfxtp_4
X_45371_ _45350_/X _61682_/B _45370_/X _45371_/Y sky130_fd_sc_hd__o21ai_4
X_57357_ _45891_/X _56995_/A _56275_/X _57364_/D _56901_/Y _57358_/A
+ sky130_fd_sc_hd__a41o_4
X_76191_ _76190_/X _76193_/A sky130_fd_sc_hd__inv_2
X_88177_ _82896_/CLK _41644_/X _67385_/B sky130_fd_sc_hd__dfxtp_4
X_42583_ _42583_/A _42583_/Y sky130_fd_sc_hd__inv_2
X_54569_ _54578_/A _53390_/B _54569_/Y sky130_fd_sc_hd__nand2_4
X_85389_ _85485_/CLK _54728_/Y _85389_/Q sky130_fd_sc_hd__dfxtp_4
X_47110_ _59245_/A _47096_/X _47109_/Y _47110_/Y sky130_fd_sc_hd__o21ai_4
X_44322_ _44321_/Y _87167_/D sky130_fd_sc_hd__inv_2
X_56308_ _56347_/A _56309_/A sky130_fd_sc_hd__buf_2
X_75142_ _75142_/A _81063_/Q _75140_/Y _75145_/C sky130_fd_sc_hd__nand3_4
X_87128_ _87436_/CLK _44400_/Y _87128_/Q sky130_fd_sc_hd__dfxtp_4
X_41534_ _81170_/Q _41471_/B _41534_/X sky130_fd_sc_hd__or2_4
X_72354_ _72352_/X _85966_/Q _72353_/X _72354_/Y sky130_fd_sc_hd__o21ai_4
X_48090_ _83536_/Q _57617_/B sky130_fd_sc_hd__inv_2
X_57288_ _57153_/A _57322_/B _57295_/A sky130_fd_sc_hd__nand2_4
X_47041_ _83044_/Q _53336_/B sky130_fd_sc_hd__inv_2
X_59027_ _58918_/A _59027_/X sky130_fd_sc_hd__buf_2
X_71305_ _70387_/A _71680_/C sky130_fd_sc_hd__buf_2
X_44253_ _44184_/A _44253_/X sky130_fd_sc_hd__buf_2
X_56239_ _56252_/A _56250_/A sky130_fd_sc_hd__buf_2
X_79950_ _60139_/C _79950_/B _79957_/A sky130_fd_sc_hd__xor2_4
X_75073_ _75067_/Y _75069_/B _75070_/Y _75074_/B sky130_fd_sc_hd__nand3_4
X_87059_ _88108_/CLK _44546_/Y _87059_/Q sky130_fd_sc_hd__dfxtp_4
X_41465_ _41464_/Y _41465_/X sky130_fd_sc_hd__buf_2
X_72285_ _83268_/Q _72250_/X _72279_/X _72284_/X _83268_/D sky130_fd_sc_hd__a2bb2oi_4
X_43204_ _43047_/X _53944_/A _40929_/X _43203_/Y _43021_/X _43204_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74024_ _73907_/X _84974_/Q _74021_/X _74023_/X _74025_/B sky130_fd_sc_hd__a211o_4
X_78901_ _82732_/Q _78901_/B _82700_/D sky130_fd_sc_hd__xor2_4
X_40416_ _40416_/A _81176_/Q _40416_/X sky130_fd_sc_hd__or2_4
X_71236_ _48872_/B _71236_/A2 _71235_/Y _71236_/Y sky130_fd_sc_hd__o21ai_4
X_44184_ _44184_/A _44184_/X sky130_fd_sc_hd__buf_2
X_79881_ _79870_/Y _79873_/Y _79881_/X sky130_fd_sc_hd__or2_4
X_41396_ _41324_/X _82892_/Q _41395_/X _41397_/A sky130_fd_sc_hd__o21ai_4
Xclkbuf_8_51_0_CLK clkbuf_8_51_0_CLK/A clkbuf_8_51_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_43135_ _87563_/Q _43135_/Y sky130_fd_sc_hd__inv_2
X_78832_ _82629_/Q _78841_/B sky130_fd_sc_hd__inv_2
X_40347_ _40361_/A _46450_/A sky130_fd_sc_hd__buf_2
X_71167_ _70611_/X _71178_/D sky130_fd_sc_hd__buf_2
X_48992_ _72012_/B _48992_/X sky130_fd_sc_hd__buf_2
X_70118_ _70102_/Y _70107_/Y _70118_/C _70118_/D _70118_/Y sky130_fd_sc_hd__nor4_4
X_47943_ _47943_/A _46371_/A _47943_/X sky130_fd_sc_hd__or2_4
X_43066_ _43038_/X _43050_/X _40667_/X _73895_/A _43061_/X _43066_/Y
+ sky130_fd_sc_hd__o32ai_4
X_59929_ _62237_/A _59918_/Y _59929_/C _59985_/A _62196_/A sky130_fd_sc_hd__and4_4
X_78763_ _78761_/X _78764_/A sky130_fd_sc_hd__inv_2
X_71098_ _50133_/B _71095_/X _71097_/Y _83609_/D sky130_fd_sc_hd__o21ai_4
X_75975_ _75961_/A _75970_/A _75975_/Y sky130_fd_sc_hd__nand2_4
X_42017_ _42017_/A _42017_/Y sky130_fd_sc_hd__inv_2
X_77714_ _82241_/Q _77713_/Y _77715_/B sky130_fd_sc_hd__xnor2_4
X_62940_ _62967_/A _63295_/A _62939_/X _62967_/D _62940_/X sky130_fd_sc_hd__and4_4
X_74926_ _74926_/A _74925_/Y _74927_/B sky130_fd_sc_hd__xor2_4
X_70049_ _68831_/X _68834_/X _70044_/X _70049_/Y sky130_fd_sc_hd__a21oi_4
X_47874_ _52309_/A _49312_/C sky130_fd_sc_hd__buf_2
Xclkbuf_8_66_0_CLK clkbuf_8_67_0_CLK/A clkbuf_8_66_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_78694_ _78690_/Y _78693_/C _78689_/Y _78694_/Y sky130_fd_sc_hd__o21ai_4
X_49613_ _86355_/Q _49606_/X _49612_/Y _49613_/Y sky130_fd_sc_hd__o21ai_4
X_46825_ _52696_/B _51003_/B sky130_fd_sc_hd__buf_2
X_77645_ _77644_/Y _77645_/B _77648_/A sky130_fd_sc_hd__nand2_4
X_74857_ _74865_/A _74856_/Y _74857_/Y sky130_fd_sc_hd__nor2_4
X_62871_ _62847_/X _58440_/Y _62911_/C _62880_/D _62871_/X sky130_fd_sc_hd__and4_4
X_64610_ _64606_/Y _60349_/X _64609_/X _64610_/X sky130_fd_sc_hd__a21o_4
X_49544_ _49561_/A _49537_/B _49522_/C _52758_/D _49544_/X sky130_fd_sc_hd__and4_4
X_61822_ _61816_/Y _61801_/X _61821_/Y _61822_/Y sky130_fd_sc_hd__a21oi_4
X_73808_ _73735_/X _85623_/Q _73782_/X _73807_/X _73808_/X sky130_fd_sc_hd__a211o_4
X_46756_ _46750_/Y _46751_/X _46755_/X _86707_/D sky130_fd_sc_hd__a21oi_4
X_65590_ _65667_/A _85878_/Q _65590_/X sky130_fd_sc_hd__and2_4
X_77576_ _77576_/A _77576_/B _77578_/A sky130_fd_sc_hd__and2_4
X_43968_ _86841_/Q _43987_/B _43955_/Y _43967_/X _43969_/B sky130_fd_sc_hd__a211o_4
X_74788_ _74788_/A _71507_/B _74788_/Y sky130_fd_sc_hd__nor2_4
X_79315_ _79303_/A _79302_/Y _79314_/X _79315_/X sky130_fd_sc_hd__a21o_4
X_45707_ _85037_/Q _45675_/X _45706_/X _45707_/Y sky130_fd_sc_hd__o21ai_4
X_64541_ _79552_/A _64532_/X _64540_/Y _84236_/D sky130_fd_sc_hd__o21ai_4
X_76527_ _76519_/X _76526_/X _76584_/A sky130_fd_sc_hd__xnor2_4
X_42919_ _42919_/A _87652_/D sky130_fd_sc_hd__inv_2
X_61753_ _61751_/Y _61699_/X _61752_/Y _61753_/Y sky130_fd_sc_hd__a21oi_4
X_49475_ _49473_/Y _49460_/X _49474_/X _86381_/D sky130_fd_sc_hd__a21oi_4
X_73739_ _73734_/X _73737_/X _73738_/X _73739_/X sky130_fd_sc_hd__a21o_4
X_46687_ _58660_/A _46672_/X _46686_/Y _46687_/Y sky130_fd_sc_hd__o21ai_4
X_43899_ _43898_/Y _87210_/D sky130_fd_sc_hd__inv_2
X_60704_ _60703_/Y _60704_/Y sky130_fd_sc_hd__inv_2
X_48426_ _48426_/A _48426_/Y sky130_fd_sc_hd__inv_2
X_79246_ _79244_/X _79246_/B _79246_/Y sky130_fd_sc_hd__xnor2_4
X_67260_ _87862_/Q _67236_/X _67167_/X _67259_/X _67260_/X sky130_fd_sc_hd__a211o_4
X_45638_ _45638_/A _45654_/B _45638_/Y sky130_fd_sc_hd__nand2_4
X_64472_ _79649_/B _64429_/X _64471_/X _64472_/X sky130_fd_sc_hd__a21o_4
X_76458_ _76439_/X _76438_/A _76458_/Y sky130_fd_sc_hd__nand2_4
X_61684_ _61292_/A _61683_/X _61675_/C _61684_/Y sky130_fd_sc_hd__nand3_4
X_66211_ _44263_/X _66211_/B _66211_/X sky130_fd_sc_hd__and2_4
X_63423_ _63484_/A _63448_/A sky130_fd_sc_hd__buf_2
X_75409_ _75409_/A _75413_/A sky130_fd_sc_hd__inv_2
X_48357_ _83593_/Q _48357_/Y sky130_fd_sc_hd__inv_2
X_60635_ _60694_/C _60725_/A _60820_/B sky130_fd_sc_hd__nand2_4
X_67191_ _87417_/Q _67121_/X _67122_/X _67190_/X _67191_/X sky130_fd_sc_hd__a211o_4
X_79177_ _79171_/Y _79176_/Y _79523_/B sky130_fd_sc_hd__nand2_4
X_45569_ _85078_/Q _55508_/B sky130_fd_sc_hd__inv_2
X_76389_ _81266_/Q _81522_/D _76389_/Y sky130_fd_sc_hd__nor2_4
X_47308_ _86648_/Q _47286_/X _47307_/Y _47308_/Y sky130_fd_sc_hd__o21ai_4
X_66142_ _64714_/X _86225_/Q _65904_/X _66141_/X _66142_/X sky130_fd_sc_hd__a211o_4
X_78128_ _78128_/A _78128_/B _78128_/X sky130_fd_sc_hd__xor2_4
X_63354_ _59450_/Y _60748_/X _60654_/X _62195_/Y _60671_/B _63354_/Y
+ sky130_fd_sc_hd__o32ai_4
X_48288_ _48285_/Y _48233_/X _48287_/X _86542_/D sky130_fd_sc_hd__a21oi_4
X_60566_ _60566_/A _60595_/C _60566_/X sky130_fd_sc_hd__and2_4
X_62305_ _62288_/X _62285_/X _64284_/B _60025_/X _62305_/X sky130_fd_sc_hd__and4_4
X_47239_ _47003_/A _47382_/A sky130_fd_sc_hd__buf_2
X_66073_ _66070_/X _66072_/X _65961_/X _66073_/X sky130_fd_sc_hd__a21o_4
X_78059_ _78059_/A _78059_/B _78059_/X sky130_fd_sc_hd__xor2_4
X_63285_ _63285_/A _63285_/B _79259_/A _63285_/Y sky130_fd_sc_hd__nor3_4
X_60497_ _60526_/A _60519_/B _79150_/A _60497_/Y sky130_fd_sc_hd__nor3_4
X_65024_ _64944_/X _86129_/Q _65022_/X _65023_/X _65024_/X sky130_fd_sc_hd__a211o_4
X_69901_ _87046_/Q _69796_/X _69797_/X _69900_/X _69902_/B sky130_fd_sc_hd__a211o_4
X_50250_ _50219_/X _50250_/X sky130_fd_sc_hd__buf_2
X_62236_ _62236_/A _62597_/B sky130_fd_sc_hd__buf_2
Xclkbuf_8_19_0_CLK clkbuf_7_9_0_CLK/X clkbuf_9_39_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_81070_ _81070_/CLK _81102_/Q _81070_/Q sky130_fd_sc_hd__dfxtp_4
X_80021_ _80004_/X _80007_/Y _80021_/X sky130_fd_sc_hd__or2_4
X_69832_ _69746_/A _69832_/X sky130_fd_sc_hd__buf_2
X_50181_ _50169_/A _49144_/X _50181_/Y sky130_fd_sc_hd__nand2_4
X_62167_ _62144_/A _62121_/X _78051_/B _62167_/Y sky130_fd_sc_hd__nor3_4
X_61118_ _61195_/A _61117_/X _72590_/A _61118_/X sky130_fd_sc_hd__o21a_4
X_69763_ _69988_/A _69763_/X sky130_fd_sc_hd__buf_2
X_66975_ _66902_/X _66975_/B _66975_/X sky130_fd_sc_hd__and2_4
X_62098_ _62097_/X _62065_/B _59608_/A _62130_/D _62099_/D sky130_fd_sc_hd__nand4_4
X_68714_ _68714_/A _69958_/A sky130_fd_sc_hd__buf_2
X_53940_ _53729_/A _53940_/X sky130_fd_sc_hd__buf_2
X_65926_ _65924_/X _84992_/Q _65865_/X _65925_/X _65927_/C sky130_fd_sc_hd__a211o_4
X_61049_ _61055_/A _61000_/X _76976_/A _61049_/X sky130_fd_sc_hd__or3_4
X_84760_ _84760_/CLK _84760_/D _80441_/A sky130_fd_sc_hd__dfxtp_4
X_81972_ _82116_/CLK _83900_/Q _81972_/Q sky130_fd_sc_hd__dfxtp_4
X_69694_ _69267_/Y _69644_/X _69672_/X _69693_/Y _69694_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_3_5_1_CLK clkbuf_3_5_0_CLK/X clkbuf_3_5_1_CLK/X sky130_fd_sc_hd__clkbuf_1
X_83711_ _83711_/CLK _83711_/D _83711_/Q sky130_fd_sc_hd__dfxtp_4
X_80923_ _81169_/CLK _80923_/D _80923_/Q sky130_fd_sc_hd__dfxtp_4
X_68645_ _69092_/A _68645_/B _68645_/X sky130_fd_sc_hd__and2_4
X_53871_ _54295_/A _53871_/X sky130_fd_sc_hd__buf_2
X_65857_ _65804_/A _85860_/Q _65857_/X sky130_fd_sc_hd__and2_4
X_84691_ _84713_/CLK _59839_/Y _80391_/A sky130_fd_sc_hd__dfxtp_4
X_55610_ _55610_/A _55610_/X sky130_fd_sc_hd__buf_2
X_86430_ _85822_/CLK _86430_/D _86430_/Q sky130_fd_sc_hd__dfxtp_4
X_52822_ _52767_/A _52843_/A sky130_fd_sc_hd__buf_2
X_64808_ _64802_/X _64805_/X _64807_/X _64808_/X sky130_fd_sc_hd__a21o_4
X_83642_ _82394_/CLK _83642_/D _46419_/A sky130_fd_sc_hd__dfxtp_4
X_56590_ _56552_/Y _56590_/X sky130_fd_sc_hd__buf_2
X_80854_ _80854_/CLK _80854_/D _74995_/B sky130_fd_sc_hd__dfxtp_4
X_68576_ _88011_/Q _68527_/X _68501_/X _68575_/X _68576_/X sky130_fd_sc_hd__a211o_4
X_65788_ _65786_/Y _65757_/X _65787_/X _84178_/D sky130_fd_sc_hd__a21o_4
X_55541_ _55538_/X _55540_/X _55516_/X _56616_/A sky130_fd_sc_hd__a21o_4
X_67527_ _67572_/A _67527_/B _67527_/X sky130_fd_sc_hd__and2_4
X_86361_ _86361_/CLK _86361_/D _86361_/Q sky130_fd_sc_hd__dfxtp_4
X_52753_ _85760_/Q _52737_/X _52752_/Y _52753_/Y sky130_fd_sc_hd__o21ai_4
X_64739_ _64739_/A _64870_/A sky130_fd_sc_hd__buf_2
X_83573_ _86505_/CLK _83573_/D _48581_/A sky130_fd_sc_hd__dfxtp_4
X_80785_ _81041_/CLK _80785_/D _75297_/A sky130_fd_sc_hd__dfxtp_4
X_88100_ _87588_/CLK _88100_/D _41938_/A sky130_fd_sc_hd__dfxtp_4
X_85312_ _85311_/CLK _56008_/Y _85312_/Q sky130_fd_sc_hd__dfxtp_4
X_51704_ _85961_/Q _51701_/X _51703_/Y _51704_/Y sky130_fd_sc_hd__o21ai_4
X_58260_ _58253_/X _83447_/Q _58259_/Y _84895_/D sky130_fd_sc_hd__o21a_4
X_82524_ _82589_/CLK _82524_/D _78707_/A sky130_fd_sc_hd__dfxtp_4
X_55472_ _55470_/A _45615_/Y _55472_/Y sky130_fd_sc_hd__nor2_4
X_67458_ _67455_/X _67457_/X _67458_/Y sky130_fd_sc_hd__nand2_4
X_86292_ _86611_/CLK _49959_/Y _72277_/B sky130_fd_sc_hd__dfxtp_4
X_52684_ _52684_/A _52684_/X sky130_fd_sc_hd__buf_2
X_57211_ _56885_/A _57126_/A _56884_/Y _57212_/A sky130_fd_sc_hd__nand3_4
X_88031_ _87273_/CLK _88031_/D _88031_/Q sky130_fd_sc_hd__dfxtp_4
X_54423_ _54399_/X _54417_/B _54402_/C _54423_/D _54423_/X sky130_fd_sc_hd__and4_4
X_66409_ _45923_/X _66410_/A sky130_fd_sc_hd__buf_2
X_85243_ _85244_/CLK _85243_/D _56303_/C sky130_fd_sc_hd__dfxtp_4
X_51635_ _51629_/X _51619_/B _51651_/C _53159_/D _51635_/X sky130_fd_sc_hd__and4_4
X_58191_ _58341_/A _58191_/X sky130_fd_sc_hd__buf_2
X_82455_ _82463_/CLK _79147_/X _82455_/Q sky130_fd_sc_hd__dfxtp_4
X_67389_ _67388_/X _67863_/A sky130_fd_sc_hd__buf_2
X_57142_ _56702_/A _56685_/B _57141_/X _57142_/X sky130_fd_sc_hd__a21bo_4
X_81406_ _83940_/CLK _83942_/Q _76755_/B sky130_fd_sc_hd__dfxtp_4
X_69128_ _69651_/A _69128_/X sky130_fd_sc_hd__buf_2
X_54354_ _54352_/Y _54338_/X _54353_/X _85458_/D sky130_fd_sc_hd__a21oi_4
X_85174_ _85270_/CLK _56495_/Y _56494_/C sky130_fd_sc_hd__dfxtp_4
X_51566_ _51621_/A _51566_/X sky130_fd_sc_hd__buf_2
X_82386_ _82386_/CLK _82194_/Q _82386_/Q sky130_fd_sc_hd__dfxtp_4
X_53305_ _53298_/A _54478_/B _53305_/Y sky130_fd_sc_hd__nand2_4
X_84125_ _84220_/CLK _84125_/D _84125_/Q sky130_fd_sc_hd__dfxtp_4
X_50517_ _50513_/A _48628_/B _50517_/Y sky130_fd_sc_hd__nand2_4
X_57073_ _57068_/X _56930_/X _57072_/Y _85093_/D sky130_fd_sc_hd__a21o_4
X_81337_ _81749_/CLK _76500_/X _81713_/D sky130_fd_sc_hd__dfxtp_4
X_69059_ _69059_/A _88343_/Q _69059_/X sky130_fd_sc_hd__and2_4
X_54285_ _54366_/A _54285_/X sky130_fd_sc_hd__buf_2
X_51497_ _85999_/Q _51485_/X _51496_/Y _51497_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_363_0_CLK clkbuf_9_181_0_CLK/X _86627_/CLK sky130_fd_sc_hd__clkbuf_1
X_56024_ _55688_/X _56020_/X _56023_/Y _56024_/Y sky130_fd_sc_hd__o21ai_4
X_41250_ _41249_/Y _41250_/X sky130_fd_sc_hd__buf_2
X_53236_ _53246_/A _53236_/B _53236_/Y sky130_fd_sc_hd__nand2_4
X_72070_ _49112_/A _72043_/X _72048_/X _72070_/X sky130_fd_sc_hd__and3_4
X_84056_ _81492_/CLK _84056_/D _84056_/Q sky130_fd_sc_hd__dfxtp_4
X_50448_ _50446_/Y _50429_/X _50447_/X _86199_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_993_0_CLK clkbuf_9_496_0_CLK/X _86523_/CLK sky130_fd_sc_hd__clkbuf_1
X_81268_ _81362_/CLK _81300_/Q _76410_/A sky130_fd_sc_hd__dfxtp_4
X_71021_ _71171_/A _70620_/B _70925_/X _71018_/D _71021_/Y sky130_fd_sc_hd__nand4_4
X_83007_ _85050_/CLK _83007_/D _83007_/Q sky130_fd_sc_hd__dfxtp_4
X_80219_ _80208_/X _80220_/B sky130_fd_sc_hd__inv_2
X_41181_ _41181_/A _41181_/X sky130_fd_sc_hd__buf_2
X_53167_ _53147_/X _53167_/B _53167_/Y sky130_fd_sc_hd__nand2_4
X_50379_ _86212_/Q _50363_/X _50378_/Y _50379_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_484_0_CLK clkbuf_8_242_0_CLK/X clkbuf_9_484_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_81199_ _82931_/CLK _81199_/D _81199_/Q sky130_fd_sc_hd__dfxtp_4
X_52118_ _52431_/A _52188_/A sky130_fd_sc_hd__buf_2
X_87815_ _87813_/CLK _42576_/Y _87815_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_378_0_CLK clkbuf_9_189_0_CLK/X _86688_/CLK sky130_fd_sc_hd__clkbuf_1
X_53098_ _53097_/X _53113_/B sky130_fd_sc_hd__buf_2
X_57975_ _57875_/X _85391_/Q _57974_/X _57975_/Y sky130_fd_sc_hd__o21ai_4
X_59714_ _60175_/A _59716_/A sky130_fd_sc_hd__buf_2
X_52049_ _52486_/A _52049_/X sky130_fd_sc_hd__buf_2
X_56926_ _56609_/X _56922_/X _56927_/C sky130_fd_sc_hd__nand2_4
X_44940_ _64235_/B _61354_/B sky130_fd_sc_hd__buf_2
X_75760_ _81014_/Q _75760_/B _80982_/D sky130_fd_sc_hd__xor2_4
X_87746_ _88012_/CLK _87746_/D _68790_/B sky130_fd_sc_hd__dfxtp_4
X_72972_ _83170_/Q _72943_/X _72971_/Y _72972_/X sky130_fd_sc_hd__a21o_4
X_84958_ _84960_/CLK _57667_/Y _57664_/A sky130_fd_sc_hd__dfxtp_4
X_74711_ _74711_/A _74711_/Y sky130_fd_sc_hd__inv_2
X_71923_ _71698_/A _71930_/B _71574_/C _71923_/Y sky130_fd_sc_hd__nor3_4
X_83909_ _83905_/CLK _83909_/D _81981_/D sky130_fd_sc_hd__dfxtp_4
X_59645_ _59604_/X _59664_/C sky130_fd_sc_hd__buf_2
Xclkbuf_9_499_0_CLK clkbuf_9_499_0_CLK/A clkbuf_9_499_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_44871_ _45297_/A _45604_/B sky130_fd_sc_hd__buf_2
X_56857_ _56856_/Y _56857_/X sky130_fd_sc_hd__buf_2
X_75691_ _75684_/Y _75685_/A _75690_/Y _75692_/B sky130_fd_sc_hd__a21oi_4
X_87677_ _87686_/CLK _42870_/Y _67095_/B sky130_fd_sc_hd__dfxtp_4
X_84889_ _84921_/CLK _58281_/X _58279_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_301_0_CLK clkbuf_9_150_0_CLK/X _84314_/CLK sky130_fd_sc_hd__clkbuf_1
X_46610_ _46610_/A _74509_/B sky130_fd_sc_hd__buf_2
X_77430_ _77426_/X _77427_/Y _77431_/B _77430_/X sky130_fd_sc_hd__a21o_4
X_43822_ _41121_/X _43817_/X _87250_/Q _43818_/X _43822_/X sky130_fd_sc_hd__a2bb2o_4
X_55808_ _55817_/A _85293_/Q _55808_/X sky130_fd_sc_hd__and2_4
X_74642_ _74675_/A _74642_/X sky130_fd_sc_hd__buf_2
X_86628_ _85990_/CLK _47504_/Y _86628_/Q sky130_fd_sc_hd__dfxtp_4
X_47590_ _47589_/Y _53135_/B sky130_fd_sc_hd__buf_2
X_71854_ _71848_/X _83353_/Q _71853_/Y _83353_/D sky130_fd_sc_hd__a21o_4
X_59576_ _59575_/Y _59662_/C sky130_fd_sc_hd__inv_2
Xclkbuf_10_931_0_CLK clkbuf_9_465_0_CLK/X _87834_/CLK sky130_fd_sc_hd__clkbuf_1
X_56788_ _56788_/A _56788_/X sky130_fd_sc_hd__buf_2
X_70805_ _70712_/A _74531_/C sky130_fd_sc_hd__buf_2
X_46541_ _46536_/Y _46523_/X _46540_/Y _46541_/Y sky130_fd_sc_hd__a21boi_4
X_58527_ _64379_/C _58528_/A sky130_fd_sc_hd__buf_2
X_77361_ _77361_/A _77361_/Y sky130_fd_sc_hd__inv_2
X_43753_ _43673_/A _43753_/X sky130_fd_sc_hd__buf_2
X_55739_ _56458_/C _55278_/A _55168_/A _55738_/X _55739_/X sky130_fd_sc_hd__a211o_4
X_86559_ _86560_/CLK _48185_/Y _65939_/B sky130_fd_sc_hd__dfxtp_4
X_74573_ _74559_/X _74569_/X _56063_/Y _74570_/X _74573_/X sky130_fd_sc_hd__a211o_4
X_40965_ _40964_/X _40941_/X _69209_/B _40942_/X _88302_/D sky130_fd_sc_hd__a2bb2o_4
X_71785_ _71714_/Y _71785_/X sky130_fd_sc_hd__buf_2
Xclkbuf_9_422_0_CLK clkbuf_9_423_0_CLK/A clkbuf_9_422_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_79100_ _79097_/Y _79099_/Y _82720_/D sky130_fd_sc_hd__nor2_4
X_76312_ _76312_/A _76312_/B _76312_/X sky130_fd_sc_hd__xor2_4
X_42704_ _42687_/X _42688_/X _41125_/X _68425_/B _42700_/X _42704_/Y
+ sky130_fd_sc_hd__o32ai_4
X_49260_ _49258_/Y _49247_/X _49259_/Y _49260_/Y sky130_fd_sc_hd__a21boi_4
X_73524_ _73522_/X _73524_/B _73524_/C _73524_/Y sky130_fd_sc_hd__nand3_4
X_46472_ _51330_/A _46428_/B _46472_/C _46472_/X sky130_fd_sc_hd__and3_4
X_70736_ _74515_/C _70730_/X _70732_/X _70735_/X _70736_/Y sky130_fd_sc_hd__nand4_4
X_58458_ _58341_/X _58454_/Y _58457_/Y _84844_/D sky130_fd_sc_hd__a21oi_4
X_77292_ _77294_/A _77294_/B _77292_/Y sky130_fd_sc_hd__nor2_4
X_43684_ _43683_/X _87311_/D sky130_fd_sc_hd__inv_2
Xclkbuf_10_316_0_CLK clkbuf_9_158_0_CLK/X _85485_/CLK sky130_fd_sc_hd__clkbuf_1
X_40896_ _40895_/Y _88315_/D sky130_fd_sc_hd__inv_2
X_48211_ _65997_/B _48203_/X _48210_/Y _48211_/Y sky130_fd_sc_hd__o21ai_4
X_79031_ _79029_/Y _79031_/B _79034_/A sky130_fd_sc_hd__xor2_4
X_45423_ _85119_/Q _44892_/X _45423_/Y sky130_fd_sc_hd__nor2_4
X_57409_ _57409_/A _56703_/X _57409_/Y sky130_fd_sc_hd__nor2_4
X_76243_ _76239_/X _76242_/Y _81608_/D sky130_fd_sc_hd__xor2_4
X_88229_ _88232_/CLK _88229_/D _67672_/B sky130_fd_sc_hd__dfxtp_4
X_42635_ _40935_/X _42631_/X _87795_/Q _42634_/X _42635_/X sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_10_946_0_CLK clkbuf_9_473_0_CLK/X _88085_/CLK sky130_fd_sc_hd__clkbuf_1
X_73455_ _73386_/A _86502_/Q _73455_/X sky130_fd_sc_hd__and2_4
X_49191_ _40623_/X _48697_/Y _49190_/Y _49192_/A sky130_fd_sc_hd__a21o_4
X_70667_ _70667_/A _70676_/B sky130_fd_sc_hd__buf_2
X_58389_ _84861_/Q _58391_/A sky130_fd_sc_hd__inv_2
X_72406_ _72299_/X _72404_/Y _72405_/Y _72337_/X _72303_/X _72406_/X
+ sky130_fd_sc_hd__o32a_4
X_48142_ _48142_/A _50383_/B _48142_/Y sky130_fd_sc_hd__nand2_4
X_60420_ _60420_/A _60421_/B sky130_fd_sc_hd__inv_2
X_45354_ _45705_/A _45354_/X sky130_fd_sc_hd__buf_2
X_76174_ _76174_/A _76176_/A _76175_/A _76174_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_9_437_0_CLK clkbuf_8_218_0_CLK/X clkbuf_9_437_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_42566_ _42521_/X _42522_/X _40814_/X _87817_/Q _42540_/X _42566_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73386_ _73386_/A _86505_/Q _73386_/X sky130_fd_sc_hd__and2_4
X_70598_ _70768_/A _70710_/A sky130_fd_sc_hd__buf_2
X_44305_ _73181_/A _44305_/X sky130_fd_sc_hd__buf_2
X_75125_ _80678_/Q _75124_/B _75127_/C sky130_fd_sc_hd__nand2_4
X_41517_ _41517_/A _41517_/Y sky130_fd_sc_hd__inv_2
X_48073_ _48092_/A _48073_/B _48073_/Y sky130_fd_sc_hd__nand2_4
X_60351_ _60350_/Y _60344_/C _60255_/A _60327_/X _60351_/X sky130_fd_sc_hd__a211o_4
X_72337_ _59133_/A _72337_/X sky130_fd_sc_hd__buf_2
X_45285_ _85160_/Q _45284_/X _45265_/X _45285_/X sky130_fd_sc_hd__o21a_4
X_42497_ _42495_/X _42496_/X _40667_/X _68727_/A _42480_/X _42498_/A
+ sky130_fd_sc_hd__o32ai_4
X_47024_ _47023_/Y _52807_/B sky130_fd_sc_hd__buf_2
X_44236_ _44196_/A _44196_/B _44235_/X _44196_/D _44236_/X sky130_fd_sc_hd__and4_4
X_63070_ _63068_/Y _63069_/X _63056_/X _63070_/Y sky130_fd_sc_hd__a21oi_4
X_75056_ _81150_/D _75046_/B _75056_/X sky130_fd_sc_hd__or2_4
X_79933_ _79926_/A _79918_/Y _79919_/Y _79934_/A sky130_fd_sc_hd__a21boi_4
X_41448_ _41447_/X _41418_/X _68047_/B _41419_/X _88213_/D sky130_fd_sc_hd__a2bb2o_4
X_72268_ _72228_/X _85973_/Q _72267_/X _72268_/Y sky130_fd_sc_hd__o21ai_4
X_60282_ _60344_/A _60221_/A _60324_/A _60284_/B sky130_fd_sc_hd__nand3_4
X_62021_ _61962_/X _62021_/B _58483_/A _62020_/X _62021_/X sky130_fd_sc_hd__and4_4
X_74007_ _87328_/Q _74246_/B _74007_/Y sky130_fd_sc_hd__nor2_4
X_71219_ _71219_/A _71076_/B _71219_/C _71219_/Y sky130_fd_sc_hd__nand3_4
X_44167_ _44006_/X _44164_/X _44166_/Y _44167_/Y sky130_fd_sc_hd__nand3_4
X_79864_ _79862_/X _79864_/B _79865_/B sky130_fd_sc_hd__xnor2_4
X_41379_ _41013_/A _41379_/X sky130_fd_sc_hd__buf_2
X_72199_ _72123_/X _85691_/Q _72146_/X _72199_/X sky130_fd_sc_hd__o21a_4
X_43118_ _43105_/X _43106_/X _40776_/X _43117_/Y _43108_/X _43118_/Y
+ sky130_fd_sc_hd__o32ai_4
X_78815_ _82627_/Q _78818_/C sky130_fd_sc_hd__inv_2
X_48975_ _86456_/Q _48952_/X _48974_/Y _48975_/Y sky130_fd_sc_hd__o21ai_4
X_44098_ _44097_/X _44098_/X sky130_fd_sc_hd__buf_2
X_79795_ _64870_/C _72224_/Y _79794_/Y _79795_/X sky130_fd_sc_hd__o21a_4
X_47926_ _47926_/A _47963_/B _47926_/X sky130_fd_sc_hd__or2_4
X_43049_ _43046_/X _43047_/X _40633_/X _43048_/Y _43034_/X _43049_/Y
+ sky130_fd_sc_hd__o32ai_4
X_78746_ _78675_/B _78740_/X _78745_/Y _78746_/Y sky130_fd_sc_hd__a21oi_4
X_66760_ _66760_/A _87691_/Q _66760_/X sky130_fd_sc_hd__and2_4
X_63972_ _63972_/A _64003_/C sky130_fd_sc_hd__buf_2
X_75958_ _75957_/A _75957_/B _75958_/Y sky130_fd_sc_hd__nor2_4
X_65711_ _65086_/X _65828_/B _65088_/X _65711_/Y sky130_fd_sc_hd__nand3_4
X_62923_ _58279_/Y _60337_/C _62923_/Y sky130_fd_sc_hd__nor2_4
X_74909_ _74904_/Y _74905_/A _74908_/Y _74909_/Y sky130_fd_sc_hd__a21boi_4
X_47857_ _48144_/A _47857_/X sky130_fd_sc_hd__buf_2
X_66691_ _66664_/X _66691_/B _66691_/X sky130_fd_sc_hd__and2_4
X_78677_ _78663_/A _78663_/B _78661_/Y _78685_/A sky130_fd_sc_hd__o21a_4
X_75889_ _75889_/A _80820_/Q _75889_/Y sky130_fd_sc_hd__xnor2_4
X_68430_ _68426_/X _68428_/X _68429_/X _68430_/X sky130_fd_sc_hd__a21o_4
X_46808_ _46667_/A _46830_/C sky130_fd_sc_hd__buf_2
X_65642_ _64851_/A _65642_/X sky130_fd_sc_hd__buf_2
X_77628_ _77628_/A _82204_/D _81916_/D sky130_fd_sc_hd__xor2_4
X_62854_ _62849_/X _62838_/X _62853_/Y _62854_/Y sky130_fd_sc_hd__a21oi_4
X_47788_ _47788_/A _53246_/B sky130_fd_sc_hd__buf_2
X_61805_ _61823_/A _61823_/B _63424_/B _61788_/X _61805_/X sky130_fd_sc_hd__and4_4
X_49527_ _86371_/Q _49524_/X _49526_/Y _49527_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_5_16_0_CLK clkbuf_4_8_1_CLK/X clkbuf_6_33_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_68361_ _68361_/A _68361_/Y sky130_fd_sc_hd__inv_2
X_46739_ _83676_/Q _52645_/B sky130_fd_sc_hd__inv_2
X_65573_ _65559_/A _65559_/B _84192_/Q _65573_/X sky130_fd_sc_hd__and3_4
X_77559_ _77559_/A _77559_/B _77559_/X sky130_fd_sc_hd__and2_4
X_62785_ _62773_/X _62762_/B _61909_/X _62785_/Y sky130_fd_sc_hd__nand3_4
X_67312_ _64706_/A _67312_/X sky130_fd_sc_hd__buf_2
X_64524_ _64545_/A _64524_/B _64545_/C _64524_/X sky130_fd_sc_hd__and3_4
X_49458_ _49454_/A _50981_/B _49458_/Y sky130_fd_sc_hd__nand2_4
X_61736_ _61736_/A _61782_/A sky130_fd_sc_hd__buf_2
X_80570_ _80566_/Y _80570_/B _80570_/Y sky130_fd_sc_hd__xnor2_4
X_68292_ _68254_/X _67792_/Y _68287_/X _68291_/Y _68292_/X sky130_fd_sc_hd__a211o_4
X_48409_ _48402_/Y _48403_/X _48408_/Y _86525_/D sky130_fd_sc_hd__a21boi_4
X_67243_ _67238_/X _67242_/X _67147_/X _67247_/A sky130_fd_sc_hd__a21o_4
X_79229_ _84791_/Q _84111_/Q _79229_/Y sky130_fd_sc_hd__nand2_4
X_64455_ _64263_/A _64455_/X sky130_fd_sc_hd__buf_2
X_49389_ _49205_/A _49410_/A sky130_fd_sc_hd__buf_2
X_61667_ _61380_/A _72563_/B sky130_fd_sc_hd__buf_2
X_51420_ _51147_/A _51420_/X sky130_fd_sc_hd__buf_2
X_63406_ _63468_/A _63456_/B sky130_fd_sc_hd__buf_2
X_82240_ _82531_/CLK _82272_/Q _82240_/Q sky130_fd_sc_hd__dfxtp_4
X_60618_ _59660_/C _61075_/B _59660_/D _60619_/A sky130_fd_sc_hd__nand3_4
X_67174_ _87110_/Q _67074_/X _67075_/X _67173_/X _67174_/X sky130_fd_sc_hd__a211o_4
X_64386_ _64386_/A _64386_/X sky130_fd_sc_hd__buf_2
X_61598_ _61686_/A _61598_/X sky130_fd_sc_hd__buf_2
X_66125_ _65484_/A _66125_/X sky130_fd_sc_hd__buf_2
X_51351_ _86027_/Q _51332_/X _51350_/Y _51351_/Y sky130_fd_sc_hd__o21ai_4
X_63337_ _79184_/A _63310_/X _63336_/X _63337_/Y sky130_fd_sc_hd__o21ai_4
X_82171_ _84111_/CLK _84163_/Q _82171_/Q sky130_fd_sc_hd__dfxtp_4
X_60549_ _60583_/A _60570_/C sky130_fd_sc_hd__buf_2
X_50302_ _50285_/A _50302_/B _50302_/Y sky130_fd_sc_hd__nand2_4
X_81122_ _81195_/CLK _81122_/D _40760_/A sky130_fd_sc_hd__dfxtp_4
X_54070_ _85511_/Q _54067_/X _54069_/Y _54070_/Y sky130_fd_sc_hd__o21ai_4
X_66056_ _66053_/X _85623_/Q _65976_/X _66055_/X _66056_/X sky130_fd_sc_hd__a211o_4
X_51282_ _51282_/A _51298_/A sky130_fd_sc_hd__buf_2
X_63268_ _63266_/Y _63267_/X _63231_/X _63268_/Y sky130_fd_sc_hd__a21oi_4
X_53021_ _53025_/A _53021_/B _53021_/Y sky130_fd_sc_hd__nand2_4
X_65007_ _64934_/X _86738_/Q _64991_/X _65006_/X _65007_/X sky130_fd_sc_hd__a211o_4
X_50233_ _86239_/Q _50220_/X _50232_/Y _50233_/Y sky130_fd_sc_hd__o21ai_4
X_62219_ _62618_/C _62219_/X sky130_fd_sc_hd__buf_2
X_85930_ _86089_/CLK _85930_/D _85930_/Q sky130_fd_sc_hd__dfxtp_4
X_81053_ _83749_/CLK _75486_/X _81053_/Q sky130_fd_sc_hd__dfxtp_4
X_63199_ _63197_/Y _63198_/X _63172_/X _63199_/Y sky130_fd_sc_hd__a21oi_4
X_80004_ _58048_/Y _65802_/C _80003_/Y _80004_/X sky130_fd_sc_hd__o21a_4
X_69815_ _70012_/A _69815_/X sky130_fd_sc_hd__buf_2
X_50164_ _50169_/A _50674_/B _50164_/Y sky130_fd_sc_hd__nand2_4
X_85861_ _86506_/CLK _85861_/D _85861_/Q sky130_fd_sc_hd__dfxtp_4
X_87600_ _87070_/CLK _43035_/Y _43032_/A sky130_fd_sc_hd__dfxtp_4
X_84812_ _85955_/CLK _84812_/D _58623_/A sky130_fd_sc_hd__dfxtp_4
X_57760_ _57759_/X _57760_/X sky130_fd_sc_hd__buf_2
X_69746_ _69746_/A _69746_/X sky130_fd_sc_hd__buf_2
X_50095_ _50103_/A _48963_/X _50095_/Y sky130_fd_sc_hd__nand2_4
X_54972_ _49793_/A _54973_/A sky130_fd_sc_hd__buf_2
X_66958_ _66952_/X _66957_/X _66958_/Y sky130_fd_sc_hd__nand2_4
X_85792_ _83685_/CLK _85792_/D _85792_/Q sky130_fd_sc_hd__dfxtp_4
X_56711_ _56651_/Y _56721_/D _56775_/A sky130_fd_sc_hd__nor2_4
X_87531_ _87782_/CLK _87531_/D _87531_/Q sky130_fd_sc_hd__dfxtp_4
X_53923_ _53951_/A _49166_/Y _53923_/Y sky130_fd_sc_hd__nand2_4
X_65909_ _65859_/X _85633_/Q _65860_/X _65908_/X _65909_/X sky130_fd_sc_hd__a211o_4
X_84743_ _83491_/CLK _59400_/X _84743_/Q sky130_fd_sc_hd__dfxtp_4
X_57691_ _57896_/A _57691_/X sky130_fd_sc_hd__buf_2
X_81955_ _81954_/CLK _83883_/Q _77883_/B sky130_fd_sc_hd__dfxtp_4
X_69677_ _42002_/A _69607_/X _68617_/X _69676_/Y _69677_/X sky130_fd_sc_hd__a211o_4
X_66889_ _66840_/X _86825_/Q _66889_/X sky130_fd_sc_hd__and2_4
X_59430_ _59430_/A _59430_/Y sky130_fd_sc_hd__inv_2
X_56642_ _55646_/X _56650_/B _56642_/Y sky130_fd_sc_hd__xnor2_4
X_80906_ _84087_/CLK _80906_/D _80906_/Q sky130_fd_sc_hd__dfxtp_4
X_68628_ _87497_/Q _68626_/X _68601_/X _68627_/X _68628_/X sky130_fd_sc_hd__a211o_4
X_87462_ _87149_/CLK _87462_/D _87462_/Q sky130_fd_sc_hd__dfxtp_4
X_53854_ _53844_/A _53854_/B _53854_/Y sky130_fd_sc_hd__nand2_4
X_84674_ _84671_/CLK _84674_/D _60021_/C sky130_fd_sc_hd__dfxtp_4
X_81886_ _82531_/CLK _81886_/D _81886_/Q sky130_fd_sc_hd__dfxtp_4
X_86413_ _85516_/CLK _86413_/D _65124_/B sky130_fd_sc_hd__dfxtp_4
X_52805_ _52784_/X _52818_/B _52789_/X _52805_/D _52805_/X sky130_fd_sc_hd__and4_4
X_83625_ _83623_/CLK _71051_/Y _83625_/Q sky130_fd_sc_hd__dfxtp_4
X_59361_ _59361_/A _59226_/B _59361_/Y sky130_fd_sc_hd__nor2_4
X_56573_ _56568_/X _56571_/X _85152_/Q _56572_/X _56573_/X sky130_fd_sc_hd__a2bb2o_4
X_80837_ _81125_/CLK _80837_/D _74870_/B sky130_fd_sc_hd__dfxtp_4
X_68559_ _68554_/X _68557_/X _68558_/X _68559_/X sky130_fd_sc_hd__a21o_4
X_87393_ _87646_/CLK _43493_/X _87393_/Q sky130_fd_sc_hd__dfxtp_4
X_53785_ _53755_/A _53786_/A sky130_fd_sc_hd__buf_2
X_50997_ _50995_/Y _50983_/X _50996_/X _86093_/D sky130_fd_sc_hd__a21oi_4
X_58312_ _58425_/A _58408_/A sky130_fd_sc_hd__buf_2
X_55524_ _55524_/A _45551_/Y _55524_/Y sky130_fd_sc_hd__nor2_4
X_86344_ _82381_/CLK _49674_/Y _86344_/Q sky130_fd_sc_hd__dfxtp_4
X_40750_ _40749_/X _40719_/X _88342_/Q _40720_/X _40750_/X sky130_fd_sc_hd__a2bb2o_4
X_52736_ _52733_/Y _52728_/X _52735_/X _52736_/Y sky130_fd_sc_hd__a21oi_4
X_59292_ _58641_/A _59292_/X sky130_fd_sc_hd__buf_2
X_71570_ _71570_/A _71570_/X sky130_fd_sc_hd__buf_2
X_83556_ _83556_/CLK _71257_/Y _83556_/Q sky130_fd_sc_hd__dfxtp_4
X_80768_ _80740_/CLK _80768_/D _80768_/Q sky130_fd_sc_hd__dfxtp_4
X_70521_ _70966_/A _70962_/C sky130_fd_sc_hd__buf_2
X_82507_ _82498_/CLK _82507_/D _82507_/Q sky130_fd_sc_hd__dfxtp_4
X_58243_ _58510_/A _58248_/B sky130_fd_sc_hd__buf_2
X_55455_ _55454_/X _45595_/Y _55455_/Y sky130_fd_sc_hd__nor2_4
X_86275_ _85955_/CLK _50047_/Y _72471_/B sky130_fd_sc_hd__dfxtp_4
XPHY_701 sky130_fd_sc_hd__decap_3
X_40681_ _40601_/X _81136_/Q _40680_/X _40682_/A sky130_fd_sc_hd__o21a_4
X_52667_ _52657_/X _52667_/B _52667_/Y sky130_fd_sc_hd__nand2_4
X_83487_ _83482_/CLK _71472_/X _83487_/Q sky130_fd_sc_hd__dfxtp_4
XPHY_712 sky130_fd_sc_hd__decap_3
X_80699_ _81082_/CLK _80699_/D _75443_/A sky130_fd_sc_hd__dfxtp_4
X_88014_ _87249_/CLK _88014_/D _88014_/Q sky130_fd_sc_hd__dfxtp_4
X_42420_ _42417_/X _42410_/X _40480_/X _87873_/Q _42411_/X _42421_/A
+ sky130_fd_sc_hd__o32ai_4
X_54406_ _54425_/A _52713_/B _54406_/Y sky130_fd_sc_hd__nand2_4
X_73240_ _73214_/X _83063_/Q _73238_/X _73239_/X _73240_/X sky130_fd_sc_hd__a211o_4
X_85226_ _85257_/CLK _85226_/D _55774_/B sky130_fd_sc_hd__dfxtp_4
X_51618_ _85977_/Q _51594_/X _51617_/Y _51618_/Y sky130_fd_sc_hd__o21ai_4
X_70452_ HASH_ADDR[0] _70758_/A sky130_fd_sc_hd__buf_2
X_58174_ _58273_/A _58217_/B sky130_fd_sc_hd__buf_2
X_82438_ _82436_/CLK _82438_/D _82438_/Q sky130_fd_sc_hd__dfxtp_4
X_55386_ _55310_/X _55315_/X _55387_/A sky130_fd_sc_hd__and2_4
X_52598_ _52626_/A _52622_/C sky130_fd_sc_hd__buf_2
Xclkbuf_7_114_0_CLK clkbuf_6_57_0_CLK/X clkbuf_8_229_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_57125_ _55481_/B _57106_/X _57124_/X _85074_/D sky130_fd_sc_hd__o21ai_4
X_54337_ _85460_/Q _54320_/X _54336_/Y _54337_/Y sky130_fd_sc_hd__o21ai_4
X_42351_ _42350_/X _42346_/X _41710_/X _87908_/Q _42347_/X _42352_/A
+ sky130_fd_sc_hd__o32ai_4
X_73171_ _73339_/A _73170_/Y _73171_/Y sky130_fd_sc_hd__nor2_4
X_85157_ _85221_/CLK _85157_/D _55732_/B sky130_fd_sc_hd__dfxtp_4
X_51549_ _51546_/Y _51531_/X _51548_/X _85990_/D sky130_fd_sc_hd__a21oi_4
X_70383_ _70994_/A _70383_/X sky130_fd_sc_hd__buf_2
X_82369_ _82369_/CLK _77044_/X _82369_/Q sky130_fd_sc_hd__dfxtp_4
X_41302_ _41301_/Y _41302_/X sky130_fd_sc_hd__buf_2
X_72122_ _59331_/X _85377_/Q _72121_/X _72122_/Y sky130_fd_sc_hd__o21ai_4
X_84108_ _84228_/CLK _84108_/D _84108_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_84_0_CLK clkbuf_9_42_0_CLK/X _84835_/CLK sky130_fd_sc_hd__clkbuf_1
X_45070_ _45219_/A _45070_/X sky130_fd_sc_hd__buf_2
X_57056_ _57055_/Y _57056_/Y sky130_fd_sc_hd__inv_2
X_42282_ _41525_/X _42271_/X _87942_/Q _42272_/X _87942_/D sky130_fd_sc_hd__a2bb2o_4
X_54268_ _54288_/A _52577_/B _54268_/Y sky130_fd_sc_hd__nand2_4
X_85088_ _83008_/CLK _57100_/X _45408_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_8_230_0_CLK clkbuf_8_231_0_CLK/A clkbuf_9_461_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_44021_ _64717_/A _64803_/A sky130_fd_sc_hd__buf_2
X_56007_ _56177_/A _56017_/B _85312_/Q _56007_/Y sky130_fd_sc_hd__nand3_4
X_41233_ _41136_/X _40714_/A _41232_/X _41233_/X sky130_fd_sc_hd__o21a_4
X_53219_ _53219_/A _53219_/B _53219_/Y sky130_fd_sc_hd__nand2_4
X_72053_ _72053_/A _53877_/B _72053_/Y sky130_fd_sc_hd__nand2_4
X_76930_ _76946_/B _76945_/A _76939_/A sky130_fd_sc_hd__xnor2_4
X_84039_ _81169_/CLK _84039_/D _82079_/D sky130_fd_sc_hd__dfxtp_4
X_54199_ _54191_/A _54191_/B _54209_/C _53031_/D _54199_/X sky130_fd_sc_hd__and4_4
X_71004_ _71071_/A _71055_/A sky130_fd_sc_hd__buf_2
X_41164_ _41143_/X _40644_/A _41163_/X _41165_/A sky130_fd_sc_hd__o21ai_4
X_76861_ _81496_/Q _81368_/D _76860_/Y _76862_/B sky130_fd_sc_hd__a21oi_4
Xclkbuf_10_99_0_CLK clkbuf_9_49_0_CLK/X _86855_/CLK sky130_fd_sc_hd__clkbuf_1
X_78600_ _78600_/A _78600_/B _78601_/A sky130_fd_sc_hd__nor2_4
X_75812_ _75811_/X _80892_/D sky130_fd_sc_hd__buf_2
X_48760_ _48840_/A _48760_/X sky130_fd_sc_hd__buf_2
X_79580_ _79580_/A _79580_/B _81093_/D sky130_fd_sc_hd__xor2_4
X_45972_ _45971_/Y _86833_/D sky130_fd_sc_hd__inv_2
X_41095_ _40878_/A _41159_/A sky130_fd_sc_hd__buf_2
X_57958_ _57971_/A _57958_/B _57958_/Y sky130_fd_sc_hd__nor2_4
X_76792_ _81666_/Q _76792_/B _76792_/Y sky130_fd_sc_hd__xnor2_4
Xclkbuf_8_245_0_CLK clkbuf_8_245_0_CLK/A clkbuf_9_491_0_CLK/A
+ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_240_0_CLK clkbuf_9_120_0_CLK/X _84449_/CLK sky130_fd_sc_hd__clkbuf_1
X_47711_ _47692_/A _47739_/B _47749_/C _53203_/D _47711_/X sky130_fd_sc_hd__and4_4
X_78531_ _78529_/Y _78530_/X _82769_/D sky130_fd_sc_hd__xnor2_4
X_44923_ _44905_/X _61329_/B _44907_/X _44923_/Y sky130_fd_sc_hd__o21ai_4
X_56909_ _55218_/Y _56908_/X _56707_/X _56909_/Y sky130_fd_sc_hd__o21ai_4
X_75743_ _81093_/Q _75743_/B _75743_/Y sky130_fd_sc_hd__xnor2_4
X_87729_ _82906_/CLK _87729_/D _67392_/B sky130_fd_sc_hd__dfxtp_4
X_48691_ _48691_/A _48894_/B _48894_/C _48691_/X sky130_fd_sc_hd__and3_4
X_72955_ _73351_/A _72955_/X sky130_fd_sc_hd__buf_2
Xclkbuf_10_870_0_CLK clkbuf_9_435_0_CLK/X _85920_/CLK sky130_fd_sc_hd__clkbuf_1
X_57889_ _72201_/A _57889_/X sky130_fd_sc_hd__buf_2
X_47642_ _86613_/Q _47619_/X _47641_/Y _47642_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_22_0_CLK clkbuf_9_11_0_CLK/X _85221_/CLK sky130_fd_sc_hd__clkbuf_1
X_71906_ _56971_/B _71892_/X _71905_/Y _83333_/D sky130_fd_sc_hd__o21ai_4
X_59628_ _59628_/A _59631_/B sky130_fd_sc_hd__buf_2
X_78462_ _78458_/Y _78460_/Y _78461_/A _78463_/B sky130_fd_sc_hd__o21ai_4
X_44854_ _44832_/X _44844_/X _41761_/X _67929_/B _44833_/X _44855_/A
+ sky130_fd_sc_hd__o32ai_4
X_75674_ _75674_/A _75673_/Y _75675_/B sky130_fd_sc_hd__xnor2_4
X_72886_ _73050_/A _72885_/Y _72886_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_9_361_0_CLK clkbuf_8_180_0_CLK/X clkbuf_9_361_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_77413_ _77412_/B _77412_/C _77412_/A _77413_/Y sky130_fd_sc_hd__o21ai_4
X_43805_ _43790_/X _43797_/X _41076_/X _87258_/Q _43791_/X _43806_/A
+ sky130_fd_sc_hd__o32ai_4
X_74625_ _74625_/A _74537_/Y _56173_/Y _74625_/Y sky130_fd_sc_hd__nand3_4
X_47573_ _47572_/Y _53127_/B sky130_fd_sc_hd__buf_2
X_71837_ _71829_/X _71839_/B _70782_/A _71826_/X _71837_/X sky130_fd_sc_hd__and4_4
X_59559_ _59558_/Y _59560_/A sky130_fd_sc_hd__inv_2
X_78393_ _78394_/A _78394_/B _78394_/C _78426_/C sky130_fd_sc_hd__a21o_4
X_44785_ _44784_/Y _86956_/D sky130_fd_sc_hd__inv_2
X_41997_ _41982_/X _41993_/X _40798_/X _41996_/Y _41984_/X _88077_/D
+ sky130_fd_sc_hd__o32ai_4
Xclkbuf_10_255_0_CLK clkbuf_9_127_0_CLK/X _82786_/CLK sky130_fd_sc_hd__clkbuf_1
X_49312_ _52528_/A _49283_/B _49312_/C _49312_/X sky130_fd_sc_hd__and3_4
X_46524_ _46401_/A _46531_/A sky130_fd_sc_hd__buf_2
X_77344_ _77339_/X _77342_/Y _77340_/Y _77345_/B sky130_fd_sc_hd__nand3_4
X_43736_ _43685_/A _43736_/X sky130_fd_sc_hd__buf_2
X_62570_ _62570_/A _62113_/X _62601_/C _62623_/D _62570_/X sky130_fd_sc_hd__and4_4
X_74556_ _44966_/Y _74551_/X _74555_/X _74556_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_885_0_CLK clkbuf_9_442_0_CLK/X _85529_/CLK sky130_fd_sc_hd__clkbuf_1
X_40948_ _82303_/Q _40970_/B _40948_/X sky130_fd_sc_hd__or2_4
X_71768_ _71763_/X _71427_/C _70794_/X _71768_/X sky130_fd_sc_hd__and3_4
Xclkbuf_10_37_0_CLK clkbuf_9_18_0_CLK/X _85057_/CLK sky130_fd_sc_hd__clkbuf_1
X_49243_ _49220_/A _53978_/B _49243_/Y sky130_fd_sc_hd__nand2_4
X_61521_ _61499_/A _61521_/B _61538_/C _61521_/Y sky130_fd_sc_hd__nand3_4
X_73507_ _73507_/A _73053_/B _73507_/Y sky130_fd_sc_hd__nor2_4
X_46455_ _83639_/Q _46455_/Y sky130_fd_sc_hd__inv_2
X_70719_ _70719_/A _70713_/X _70727_/C _70710_/D _70719_/Y sky130_fd_sc_hd__nand4_4
X_77275_ _77273_/X _77274_/Y _77277_/B sky130_fd_sc_hd__nand2_4
X_43667_ _43667_/A _69055_/B sky130_fd_sc_hd__inv_2
X_74487_ _74458_/A _74501_/C sky130_fd_sc_hd__buf_2
Xclkbuf_9_376_0_CLK clkbuf_8_188_0_CLK/X clkbuf_9_376_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_40879_ _46469_/B _40879_/B _40879_/X sky130_fd_sc_hd__or2_4
X_71699_ _71691_/Y _83407_/Q _71698_/Y _83407_/D sky130_fd_sc_hd__a21o_4
X_79014_ _79012_/Y _79014_/B _79018_/A sky130_fd_sc_hd__xor2_4
X_45406_ _45350_/X _61315_/A _45370_/X _45406_/Y sky130_fd_sc_hd__o21ai_4
X_64240_ _64233_/Y _64239_/X _72577_/B _64240_/X sky130_fd_sc_hd__o21a_4
X_76226_ _76226_/A _81607_/D _76226_/X sky130_fd_sc_hd__xor2_4
X_42618_ _42614_/X _42615_/X _40914_/X _69929_/A _42597_/X _42619_/A
+ sky130_fd_sc_hd__o32ai_4
X_49174_ _49169_/Y _49138_/X _49173_/X _86437_/D sky130_fd_sc_hd__a21oi_4
X_61452_ _59399_/A _61452_/B _61452_/C _61452_/D _61453_/A sky130_fd_sc_hd__nand4_4
X_73438_ _73438_/A _73438_/B _73438_/Y sky130_fd_sc_hd__nor2_4
X_46386_ _52480_/B _49265_/B sky130_fd_sc_hd__buf_2
X_43598_ _43598_/A _43598_/Y sky130_fd_sc_hd__inv_2
X_48125_ _66310_/B _48103_/X _48124_/Y _48125_/Y sky130_fd_sc_hd__o21ai_4
X_60403_ _60403_/A _60403_/B _60403_/C _60414_/B _60404_/B sky130_fd_sc_hd__and4_4
X_45337_ _55722_/B _45281_/X _45311_/X _45337_/X sky130_fd_sc_hd__o21a_4
X_76157_ _81346_/Q _81602_/D _76157_/X sky130_fd_sc_hd__xor2_4
X_64171_ _62162_/X _64182_/B _64182_/C _64182_/D _64171_/Y sky130_fd_sc_hd__nand4_4
X_42549_ _42536_/X _42547_/X _40776_/X _42548_/Y _42538_/X _42549_/Y
+ sky130_fd_sc_hd__o32ai_4
X_73369_ _83154_/Q _73318_/X _73368_/Y _83154_/D sky130_fd_sc_hd__a21o_4
X_61383_ _61375_/Y _61377_/Y _61334_/X _61378_/Y _61382_/Y _61383_/X
+ sky130_fd_sc_hd__a41o_4
X_75108_ _75108_/A _75107_/Y _75108_/X sky130_fd_sc_hd__xor2_4
X_63122_ _63088_/A _64335_/C _63087_/X _63077_/D _63122_/X sky130_fd_sc_hd__and4_4
X_48056_ _48056_/A _47973_/B _48056_/X sky130_fd_sc_hd__or2_4
X_60334_ _60296_/X _60241_/A _60300_/C _60367_/D _60334_/Y sky130_fd_sc_hd__nand4_4
X_45268_ _45264_/Y _45267_/Y _45212_/X _45268_/X sky130_fd_sc_hd__a21o_4
X_76088_ _81720_/D _76075_/B _76087_/Y _76089_/B sky130_fd_sc_hd__a21oi_4
X_47007_ _47006_/Y _52799_/B sky130_fd_sc_hd__buf_2
X_44219_ _44054_/Y _44185_/X _44204_/Y _44218_/X _44220_/A sky130_fd_sc_hd__o22a_4
X_67930_ _87386_/Q _67834_/X _67835_/X _67929_/X _67930_/X sky130_fd_sc_hd__a211o_4
X_63053_ _63053_/A _63081_/B sky130_fd_sc_hd__buf_2
X_75039_ _75038_/X _75039_/X sky130_fd_sc_hd__buf_2
X_79916_ _79902_/Y _80262_/B _79932_/A sky130_fd_sc_hd__nor2_4
X_60265_ _60513_/A _61587_/B _79826_/A _60265_/X sky130_fd_sc_hd__or3_4
Xclkbuf_10_823_0_CLK clkbuf_9_411_0_CLK/X _84981_/CLK sky130_fd_sc_hd__clkbuf_1
X_45199_ _45199_/A _45199_/B _45199_/Y sky130_fd_sc_hd__nand2_4
X_62004_ _61962_/X _61945_/X _58478_/A _61947_/D _62004_/X sky130_fd_sc_hd__and4_4
X_79847_ _79845_/X _79860_/B _79866_/B sky130_fd_sc_hd__xnor2_4
X_67861_ _86953_/Q _67788_/X _67789_/X _67860_/X _67861_/X sky130_fd_sc_hd__a211o_4
X_60196_ _62737_/A _60197_/C sky130_fd_sc_hd__buf_2
Xclkbuf_9_314_0_CLK clkbuf_9_315_0_CLK/A clkbuf_9_314_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_69600_ _69167_/X _69170_/X _69575_/X _69600_/Y sky130_fd_sc_hd__a21oi_4
X_66812_ _66809_/X _66811_/X _66787_/X _66815_/A sky130_fd_sc_hd__a21o_4
X_48958_ _49048_/A _48958_/B _50599_/A sky130_fd_sc_hd__nor2_4
X_67792_ _67792_/A _67791_/X _67792_/Y sky130_fd_sc_hd__nand2_4
X_79778_ _79762_/X _79766_/B _79778_/X sky130_fd_sc_hd__or2_4
Xclkbuf_10_208_0_CLK clkbuf_9_104_0_CLK/X _84508_/CLK sky130_fd_sc_hd__clkbuf_1
X_69531_ _69956_/A _69531_/B _69531_/X sky130_fd_sc_hd__and2_4
X_47909_ _47902_/Y _47903_/X _47908_/X _86587_/D sky130_fd_sc_hd__a21oi_4
X_66743_ _66743_/A _66742_/X _66743_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_10_838_0_CLK clkbuf_9_419_0_CLK/X _82973_/CLK sky130_fd_sc_hd__clkbuf_1
X_78729_ _78729_/A _82686_/D _78732_/B sky130_fd_sc_hd__nor2_4
X_63955_ _64032_/A _63955_/X sky130_fd_sc_hd__buf_2
X_48889_ _48695_/A _48889_/B _48889_/Y sky130_fd_sc_hd__nand2_4
X_50920_ _50917_/Y _50902_/X _50919_/X _50920_/Y sky130_fd_sc_hd__a21oi_4
X_81740_ _84003_/CLK _81740_/D _81740_/Q sky130_fd_sc_hd__dfxtp_4
X_62906_ _63630_/A _62875_/X _62905_/Y _62906_/X sky130_fd_sc_hd__o21a_4
X_69462_ _68946_/X _68950_/X _69418_/X _69462_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_329_0_CLK clkbuf_9_329_0_CLK/A clkbuf_9_329_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_66674_ _66673_/X _66794_/A sky130_fd_sc_hd__buf_2
X_63886_ _60915_/X _63902_/B sky130_fd_sc_hd__buf_2
X_68413_ _83976_/Q _68338_/X _68412_/X _68413_/X sky130_fd_sc_hd__a21bo_4
X_65625_ _65623_/X _86196_/Q _65517_/X _65624_/X _65625_/X sky130_fd_sc_hd__a211o_4
X_50851_ _50848_/Y _50849_/X _50850_/Y _50851_/Y sky130_fd_sc_hd__a21boi_4
X_62837_ _62830_/Y _62831_/X _62833_/Y _62834_/Y _62836_/X _62837_/X
+ sky130_fd_sc_hd__a41o_4
X_81671_ _81671_/CLK _79982_/X _81671_/Q sky130_fd_sc_hd__dfxtp_4
X_69393_ _69245_/A _69393_/X sky130_fd_sc_hd__buf_2
X_83410_ _83380_/CLK _83410_/D _83410_/Q sky130_fd_sc_hd__dfxtp_4
X_80622_ _80622_/A _80622_/B _80624_/A sky130_fd_sc_hd__nand2_4
X_68344_ _88019_/Q _69796_/A _66295_/X _68343_/X _68344_/X sky130_fd_sc_hd__a211o_4
X_65556_ _65553_/X _65663_/B _65556_/C _65556_/Y sky130_fd_sc_hd__nand3_4
X_53570_ _52050_/A _53620_/B _53620_/C _53570_/X sky130_fd_sc_hd__and3_4
X_84390_ _84392_/CLK _62698_/Y _84390_/Q sky130_fd_sc_hd__dfxtp_4
X_50782_ _86134_/Q _50775_/X _50781_/Y _50782_/Y sky130_fd_sc_hd__o21ai_4
X_62768_ _60309_/D _62768_/X sky130_fd_sc_hd__buf_2
X_52521_ _52519_/Y _52496_/X _52520_/X _52521_/Y sky130_fd_sc_hd__a21oi_4
X_64507_ _64501_/X _64504_/Y _64506_/Y _84871_/Q _64213_/X _64507_/Y
+ sky130_fd_sc_hd__o32ai_4
X_83341_ _83491_/CLK _83341_/D _59437_/B sky130_fd_sc_hd__dfxtp_4
X_61719_ _61719_/A _61719_/X sky130_fd_sc_hd__buf_2
X_80553_ _80537_/X _80541_/B _80552_/X _80553_/X sky130_fd_sc_hd__a21o_4
X_68275_ _82643_/D _68259_/X _68274_/X _83995_/D sky130_fd_sc_hd__a21bo_4
X_65487_ _65667_/A _85885_/Q _65487_/X sky130_fd_sc_hd__and2_4
X_62699_ _60211_/A _62699_/X sky130_fd_sc_hd__buf_2
X_55240_ _55237_/Y _55240_/B _55241_/B sky130_fd_sc_hd__nor2_4
X_67226_ _67226_/A _67226_/X sky130_fd_sc_hd__buf_2
X_86060_ _85741_/CLK _86060_/D _86060_/Q sky130_fd_sc_hd__dfxtp_4
X_52452_ _52466_/A _53971_/B _52452_/Y sky130_fd_sc_hd__nand2_4
X_64438_ _64515_/A _84862_/Q _64515_/C _64438_/Y sky130_fd_sc_hd__nand3_4
X_83272_ _83627_/CLK _83272_/D _72224_/A sky130_fd_sc_hd__dfxtp_4
X_80484_ _80484_/A _84316_/Q _80494_/B sky130_fd_sc_hd__xor2_4
X_85011_ _85075_/CLK _85011_/D _85011_/Q sky130_fd_sc_hd__dfxtp_4
X_51403_ _51211_/A _51403_/X sky130_fd_sc_hd__buf_2
X_82223_ _81839_/CLK _82255_/Q _82223_/Q sky130_fd_sc_hd__dfxtp_4
X_55171_ _55167_/X _55170_/X _44109_/X _55171_/X sky130_fd_sc_hd__a21o_4
X_67157_ _67133_/A _86782_/Q _67157_/X sky130_fd_sc_hd__and2_4
X_52383_ _52373_/X _49125_/X _52383_/Y sky130_fd_sc_hd__nand2_4
X_64369_ _58331_/A _64367_/X _64368_/Y _64369_/Y sky130_fd_sc_hd__o21ai_4
X_54122_ _85500_/Q _54113_/X _54121_/Y _54122_/Y sky130_fd_sc_hd__o21ai_4
X_66108_ _84156_/Q _66109_/C sky130_fd_sc_hd__inv_2
X_51334_ _51790_/A _51350_/A sky130_fd_sc_hd__buf_2
X_82154_ _84220_/CLK _66247_/C _82154_/Q sky130_fd_sc_hd__dfxtp_4
X_67088_ _87114_/Q _66988_/X _67040_/X _67087_/X _67088_/X sky130_fd_sc_hd__a211o_4
X_81105_ _81104_/CLK _79718_/X _81105_/Q sky130_fd_sc_hd__dfxtp_4
X_58930_ _58891_/X _86085_/Q _58929_/X _58930_/Y sky130_fd_sc_hd__o21ai_4
X_54053_ _54050_/Y _54051_/X _54052_/X _54053_/Y sky130_fd_sc_hd__a21oi_4
X_66039_ _66036_/X _66038_/X _65880_/X _66043_/A sky130_fd_sc_hd__a21o_4
X_51265_ _51265_/A _51266_/B sky130_fd_sc_hd__buf_2
X_86962_ _86965_/CLK _86962_/D _86962_/Q sky130_fd_sc_hd__dfxtp_4
X_82085_ _81989_/CLK _77265_/B _82085_/Q sky130_fd_sc_hd__dfxtp_4
X_53004_ _53000_/Y _53001_/X _53003_/X _53004_/Y sky130_fd_sc_hd__a21oi_4
X_50216_ _86241_/Q _41872_/X _50215_/X _50217_/A sky130_fd_sc_hd__o21ai_4
X_85913_ _85915_/CLK _51978_/Y _66022_/B sky130_fd_sc_hd__dfxtp_4
X_81036_ _82084_/CLK _81036_/D _81036_/Q sky130_fd_sc_hd__dfxtp_4
X_58861_ _58846_/X _85770_/Q _58847_/X _58861_/X sky130_fd_sc_hd__o21a_4
X_51196_ _51170_/A _51197_/C sky130_fd_sc_hd__buf_2
X_86893_ _86896_/CLK _45186_/Y _64420_/B sky130_fd_sc_hd__dfxtp_4
X_57812_ _57705_/X _85500_/Q _57736_/X _57812_/X sky130_fd_sc_hd__o21a_4
X_50147_ _52355_/A _50082_/B _50147_/C _50147_/X sky130_fd_sc_hd__and3_4
X_85844_ _85535_/CLK _52333_/Y _85844_/Q sky130_fd_sc_hd__dfxtp_4
X_58792_ _84799_/Q _58792_/Y sky130_fd_sc_hd__inv_2
X_57743_ _84951_/Q _57691_/X _57735_/X _57742_/X _84951_/D sky130_fd_sc_hd__a2bb2oi_4
X_69729_ _69307_/X _69310_/X _69728_/X _69729_/Y sky130_fd_sc_hd__a21oi_4
X_50078_ _48928_/A _50082_/B _50059_/C _50078_/X sky130_fd_sc_hd__and3_4
X_54955_ _54955_/A _54955_/B _46617_/A _53261_/D _54955_/X sky130_fd_sc_hd__and4_4
X_85775_ _85778_/CLK _52676_/Y _85775_/Q sky130_fd_sc_hd__dfxtp_4
X_82987_ _82987_/CLK _82987_/D _45745_/A sky130_fd_sc_hd__dfxtp_4
X_87514_ _87520_/CLK _87514_/D _87514_/Q sky130_fd_sc_hd__dfxtp_4
X_41920_ _88105_/Q _41920_/Y sky130_fd_sc_hd__inv_2
X_53906_ _53902_/A _72079_/B _53906_/Y sky130_fd_sc_hd__nand2_4
X_72740_ _72739_/X _73007_/A sky130_fd_sc_hd__buf_2
X_84726_ _84732_/CLK _84726_/D _84726_/Q sky130_fd_sc_hd__dfxtp_4
X_57674_ _57674_/A _57674_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_7_91_0_CLK clkbuf_7_91_0_CLK/A clkbuf_7_91_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_81938_ _81954_/CLK _81938_/D _81938_/Q sky130_fd_sc_hd__dfxtp_4
X_54886_ _85359_/Q _54865_/X _54885_/Y _54886_/Y sky130_fd_sc_hd__o21ai_4
X_59413_ _84739_/Q _59413_/Y sky130_fd_sc_hd__inv_2
X_56625_ _56629_/B _56580_/B _56609_/X _56624_/Y _56626_/A sky130_fd_sc_hd__a211o_4
X_87445_ _87382_/CLK _87445_/D _87445_/Q sky130_fd_sc_hd__dfxtp_4
X_41851_ _41851_/A _41851_/Y sky130_fd_sc_hd__inv_2
X_53837_ _85558_/Q _53816_/X _53836_/Y _53837_/Y sky130_fd_sc_hd__o21ai_4
X_72671_ _83195_/Q _72658_/X _72670_/Y _72671_/X sky130_fd_sc_hd__a21bo_4
X_84657_ _84508_/CLK _84657_/D _79998_/A sky130_fd_sc_hd__dfxtp_4
X_81869_ _81834_/CLK _78060_/X _81869_/Q sky130_fd_sc_hd__dfxtp_4
X_74410_ _48464_/A _74395_/X _74421_/C _74410_/X sky130_fd_sc_hd__and3_4
X_40802_ _40802_/A _40802_/X sky130_fd_sc_hd__buf_2
X_71622_ _71867_/A _70667_/A _71215_/C _71622_/D _71622_/Y sky130_fd_sc_hd__nor4_4
X_83608_ _85837_/CLK _83608_/D _49054_/A sky130_fd_sc_hd__dfxtp_4
X_59344_ _64713_/A _64678_/A sky130_fd_sc_hd__buf_2
X_44570_ _44570_/A _44570_/Y sky130_fd_sc_hd__inv_2
X_56556_ _56556_/A _56556_/Y sky130_fd_sc_hd__inv_2
X_87376_ _87995_/CLK _43526_/X _87376_/Q sky130_fd_sc_hd__dfxtp_4
X_75390_ _75390_/A _75390_/B _75390_/X sky130_fd_sc_hd__xor2_4
X_41782_ _41781_/Y _41782_/X sky130_fd_sc_hd__buf_2
X_53768_ _48691_/A _53774_/B _53774_/C _53768_/X sky130_fd_sc_hd__and3_4
X_84588_ _84590_/CLK _84588_/D _79128_/A sky130_fd_sc_hd__dfxtp_4
X_43521_ _41797_/X _43513_/X _87379_/Q _43514_/X _43521_/X sky130_fd_sc_hd__a2bb2o_4
X_55507_ _55462_/X _55507_/X sky130_fd_sc_hd__buf_2
X_74341_ _45883_/B _74351_/A sky130_fd_sc_hd__buf_2
X_86327_ _86322_/CLK _49767_/Y _57870_/B sky130_fd_sc_hd__dfxtp_4
X_40733_ _40731_/X _82855_/Q _40732_/X _40733_/Y sky130_fd_sc_hd__o21ai_4
X_52719_ _85767_/Q _52711_/X _52718_/Y _52719_/Y sky130_fd_sc_hd__o21ai_4
X_59275_ _59260_/X _85419_/Q _59274_/X _59275_/Y sky130_fd_sc_hd__o21ai_4
X_71553_ _70692_/A _71553_/B _71536_/A _71553_/Y sky130_fd_sc_hd__nor3_4
X_83539_ _86530_/CLK _71315_/Y _48060_/A sky130_fd_sc_hd__dfxtp_4
X_56487_ _56525_/A _56487_/X sky130_fd_sc_hd__buf_2
X_53699_ _53713_/A _48538_/Y _53699_/Y sky130_fd_sc_hd__nand2_4
X_46240_ _46240_/A _48882_/A _46240_/Y sky130_fd_sc_hd__nand2_4
X_70504_ _70504_/A _70511_/A sky130_fd_sc_hd__buf_2
X_58226_ _58225_/X _58238_/B _58226_/Y sky130_fd_sc_hd__nor2_4
XPHY_520 sky130_fd_sc_hd__decap_3
X_77060_ _77060_/A _77060_/B _77060_/X sky130_fd_sc_hd__xor2_4
X_55438_ _55380_/Y _55438_/B _55441_/A sky130_fd_sc_hd__nor2_4
X_43452_ _43425_/X _43452_/X sky130_fd_sc_hd__buf_2
X_74272_ _74012_/X _86210_/Q _45930_/X _74271_/X _74272_/X sky130_fd_sc_hd__a211o_4
X_86258_ _85555_/CLK _86258_/D _65012_/B sky130_fd_sc_hd__dfxtp_4
XPHY_531 sky130_fd_sc_hd__decap_3
X_40664_ _40420_/A _40829_/A sky130_fd_sc_hd__buf_2
X_71484_ _71463_/Y _83482_/Q _71483_/X _83482_/D sky130_fd_sc_hd__a21o_4
XPHY_542 sky130_fd_sc_hd__decap_3
XPHY_553 sky130_fd_sc_hd__decap_3
X_76011_ _81518_/Q _81742_/D _76011_/X sky130_fd_sc_hd__xor2_4
X_42403_ _42403_/A _42403_/Y sky130_fd_sc_hd__inv_2
XPHY_564 sky130_fd_sc_hd__decap_3
X_73223_ _83160_/Q _73193_/X _73222_/Y _73223_/X sky130_fd_sc_hd__a21o_4
X_85209_ _85241_/CLK _85209_/D _85209_/Q sky130_fd_sc_hd__dfxtp_4
X_46171_ _46170_/Y _72498_/B _46171_/Y sky130_fd_sc_hd__nand2_4
X_70435_ _70442_/A _74523_/A _70431_/C _70435_/Y sky130_fd_sc_hd__nand3_4
X_58157_ _58153_/X _83495_/Q _58156_/Y _84919_/D sky130_fd_sc_hd__o21a_4
XPHY_575 sky130_fd_sc_hd__decap_3
X_43383_ _43382_/Y _87450_/D sky130_fd_sc_hd__inv_2
X_55369_ _55369_/A _55369_/B _55368_/Y _55443_/C sky130_fd_sc_hd__nand3_4
X_86189_ _86505_/CLK _86189_/D _86189_/Q sky130_fd_sc_hd__dfxtp_4
X_40595_ _49569_/A _40595_/X sky130_fd_sc_hd__buf_2
XPHY_586 sky130_fd_sc_hd__decap_3
XPHY_597 sky130_fd_sc_hd__decap_3
X_45122_ _45122_/A _45124_/A sky130_fd_sc_hd__inv_2
X_57108_ _56600_/X _57106_/X _57107_/Y _85083_/D sky130_fd_sc_hd__a21oi_4
X_42334_ _42330_/X _42319_/X _41667_/X _87916_/Q _42320_/X _42335_/A
+ sky130_fd_sc_hd__o32ai_4
X_73154_ _88324_/Q _73153_/X _72901_/X _73154_/Y sky130_fd_sc_hd__o21ai_4
X_58088_ _59036_/A _58928_/A sky130_fd_sc_hd__buf_2
X_70366_ _71129_/A _70366_/X sky130_fd_sc_hd__buf_2
X_72105_ _72091_/X _53932_/B _72105_/Y sky130_fd_sc_hd__nand2_4
X_49930_ _52679_/A _49930_/X sky130_fd_sc_hd__buf_2
X_57039_ _57039_/A _57026_/X _57039_/Y sky130_fd_sc_hd__nor2_4
X_45053_ _64320_/B _61437_/B sky130_fd_sc_hd__buf_2
X_42265_ _41485_/X _42258_/X _87950_/Q _42259_/X _42265_/X sky130_fd_sc_hd__a2bb2o_4
X_77962_ _77954_/A _77954_/B _77961_/Y _77967_/C sky130_fd_sc_hd__o21a_4
X_73085_ _73082_/X _73084_/X _72951_/X _73101_/B sky130_fd_sc_hd__a21o_4
X_70297_ _70247_/X _70297_/X sky130_fd_sc_hd__buf_2
X_44004_ _62975_/D _60665_/C _44003_/X _44004_/Y sky130_fd_sc_hd__nand3_4
X_79701_ _79699_/X _79710_/B _79701_/Y sky130_fd_sc_hd__xnor2_4
X_41216_ _41216_/A _41216_/Y sky130_fd_sc_hd__inv_2
X_60050_ _59929_/C _59910_/X _59927_/Y _62203_/A sky130_fd_sc_hd__nand3_4
X_72036_ _72017_/X _53860_/B _72036_/Y sky130_fd_sc_hd__nand2_4
X_76913_ _76870_/Y _76910_/X _76912_/X _76914_/B sky130_fd_sc_hd__a21boi_4
Xclkbuf_7_44_0_CLK clkbuf_6_22_0_CLK/X clkbuf_8_89_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_49861_ _49861_/A _49884_/B sky130_fd_sc_hd__buf_2
X_42196_ _41302_/X _42192_/X _87984_/Q _42193_/X _87984_/D sky130_fd_sc_hd__a2bb2o_4
X_77893_ _77880_/A _77887_/A _77893_/X sky130_fd_sc_hd__and2_4
Xclkbuf_8_184_0_CLK clkbuf_7_92_0_CLK/X clkbuf_8_184_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_48812_ _86478_/Q _48809_/X _48811_/Y _48812_/Y sky130_fd_sc_hd__o21ai_4
X_79632_ _79624_/A _79624_/B _79619_/A _79632_/Y sky130_fd_sc_hd__o21ai_4
X_41147_ _41147_/A _41147_/X sky130_fd_sc_hd__buf_2
X_76844_ _76844_/A _76843_/Y _76845_/B sky130_fd_sc_hd__xnor2_4
X_49792_ _57934_/B _49768_/X _49791_/Y _49792_/Y sky130_fd_sc_hd__o21ai_4
X_48743_ _52573_/B _48766_/B sky130_fd_sc_hd__buf_2
X_79563_ _79547_/Y _79563_/B _79563_/Y sky130_fd_sc_hd__xnor2_4
X_45955_ _44196_/B _45955_/X sky130_fd_sc_hd__buf_2
X_41078_ _41078_/A _41078_/Y sky130_fd_sc_hd__inv_2
X_76775_ _76763_/A _76770_/A _76776_/B sky130_fd_sc_hd__and2_4
X_73987_ _73987_/A _57376_/X _73987_/Y sky130_fd_sc_hd__nor2_4
Xclkbuf_7_59_0_CLK clkbuf_7_58_0_CLK/A clkbuf_7_59_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_78514_ _78486_/Y _78514_/Y sky130_fd_sc_hd__inv_2
X_44906_ _44290_/X _44907_/A sky130_fd_sc_hd__buf_2
X_63740_ _63735_/A _63741_/A sky130_fd_sc_hd__buf_2
X_75726_ _81091_/Q _75726_/B _75726_/Y sky130_fd_sc_hd__xnor2_4
X_48674_ _86501_/Q _48669_/X _48673_/Y _48674_/Y sky130_fd_sc_hd__o21ai_4
X_60952_ _60951_/Y _60952_/X sky130_fd_sc_hd__buf_2
X_72938_ _53647_/B _72938_/B _72938_/X sky130_fd_sc_hd__xor2_4
X_79494_ _79494_/A _79494_/B _79494_/Y sky130_fd_sc_hd__xnor2_4
X_45886_ _45885_/X _45886_/X sky130_fd_sc_hd__buf_2
Xclkbuf_8_199_0_CLK clkbuf_7_99_0_CLK/X clkbuf_9_398_0_CLK/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_194_0_CLK clkbuf_9_97_0_CLK/X _83749_/CLK sky130_fd_sc_hd__clkbuf_1
X_47625_ _72247_/A _47619_/X _47624_/Y _47625_/Y sky130_fd_sc_hd__o21ai_4
X_78445_ _78432_/A _82667_/D _78439_/C _78466_/A sky130_fd_sc_hd__a21boi_4
X_63671_ _63669_/Y _63635_/X _63670_/Y _84303_/D sky130_fd_sc_hd__a21oi_4
X_44837_ _44837_/A _86928_/D sky130_fd_sc_hd__inv_2
X_75657_ _75657_/A _75657_/B _75657_/Y sky130_fd_sc_hd__xnor2_4
X_60883_ _60864_/X _60984_/A sky130_fd_sc_hd__buf_2
X_72869_ _72869_/A _72868_/Y _72869_/Y sky130_fd_sc_hd__nand2_4
X_65410_ _65410_/A _65409_/X _65410_/Y sky130_fd_sc_hd__nand2_4
X_74608_ _74605_/X _74599_/X _56138_/Y _74600_/X _74608_/X sky130_fd_sc_hd__a211o_4
X_62622_ _62622_/A _62619_/Y _62622_/C _62621_/Y _62622_/Y sky130_fd_sc_hd__nand4_4
X_47556_ _47556_/A _47595_/B sky130_fd_sc_hd__buf_2
X_66390_ _66386_/Y _66377_/X _66389_/Y _84132_/D sky130_fd_sc_hd__a21o_4
X_78376_ _78364_/C _78376_/B _78378_/A sky130_fd_sc_hd__nand2_4
X_44768_ _44532_/A _44768_/X sky130_fd_sc_hd__buf_2
X_75588_ _75586_/A _75584_/Y _75583_/A _75588_/Y sky130_fd_sc_hd__a21oi_4
Xclkbuf_8_122_0_CLK clkbuf_7_61_0_CLK/X clkbuf_9_245_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_46507_ _46507_/A _52533_/A sky130_fd_sc_hd__buf_2
X_65341_ _64656_/A _65660_/A sky130_fd_sc_hd__buf_2
X_77327_ _77323_/Y _77325_/Y _77326_/Y _77327_/Y sky130_fd_sc_hd__o21ai_4
X_43719_ _40861_/A _43716_/X _69808_/B _43718_/X _43719_/X sky130_fd_sc_hd__a2bb2o_4
X_62553_ _62672_/A _62553_/X sky130_fd_sc_hd__buf_2
X_74539_ _74539_/A _45933_/Y _55684_/X _74549_/A sky130_fd_sc_hd__nand3_4
X_47487_ _47513_/A _47463_/X _47513_/C _53074_/D _47487_/X sky130_fd_sc_hd__and4_4
X_44699_ _44679_/X _44680_/X _40656_/X _86995_/Q _44681_/X _44700_/A
+ sky130_fd_sc_hd__o32ai_4
X_49226_ _49220_/A _53959_/B _49226_/Y sky130_fd_sc_hd__nand2_4
X_61504_ _59415_/A _61484_/B _61484_/C _61514_/D _61504_/Y sky130_fd_sc_hd__nand4_4
X_68060_ _68371_/A _88149_/Q _68060_/X sky130_fd_sc_hd__and2_4
X_46438_ _46438_/A _50808_/B sky130_fd_sc_hd__buf_2
X_65272_ _65118_/A _65272_/X sky130_fd_sc_hd__buf_2
X_77258_ _77258_/A _77255_/Y _77252_/Y _77258_/Y sky130_fd_sc_hd__nand3_4
X_62484_ _62179_/X _62541_/B sky130_fd_sc_hd__buf_2
X_67011_ _66942_/A _67011_/B _67011_/X sky130_fd_sc_hd__and2_4
X_76209_ _76206_/Y _76208_/Y _76209_/Y sky130_fd_sc_hd__nor2_4
X_64223_ _64223_/A _64223_/B _64223_/C _64223_/X sky130_fd_sc_hd__and3_4
X_49157_ _49157_/A _53917_/B sky130_fd_sc_hd__inv_2
X_61435_ _61433_/X _61394_/X _61434_/Y _61435_/Y sky130_fd_sc_hd__a21oi_4
X_46369_ _46387_/A _50777_/B _46369_/Y sky130_fd_sc_hd__nand2_4
X_77189_ _77185_/Y _77177_/B _77188_/X _77189_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_8_137_0_CLK clkbuf_7_68_0_CLK/X clkbuf_9_274_0_CLK/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_10_132_0_CLK clkbuf_9_66_0_CLK/X _83813_/CLK sky130_fd_sc_hd__clkbuf_1
X_48108_ _66285_/B _48103_/X _48107_/Y _48108_/Y sky130_fd_sc_hd__o21ai_4
X_64154_ _64152_/X _64129_/X _64153_/Y _84270_/D sky130_fd_sc_hd__a21oi_4
X_61366_ _61377_/A _61365_/X _61377_/C _61366_/Y sky130_fd_sc_hd__nand3_4
X_49088_ _40601_/X _81197_/Q _49087_/Y _49089_/A sky130_fd_sc_hd__o21ai_4
Xclkbuf_10_762_0_CLK clkbuf_9_381_0_CLK/X _87520_/CLK sky130_fd_sc_hd__clkbuf_1
X_63105_ _79427_/A _63072_/X _63104_/Y _63105_/X sky130_fd_sc_hd__a21o_4
X_60317_ _60317_/A _60244_/B _79733_/A _60317_/Y sky130_fd_sc_hd__nor3_4
X_48039_ _48039_/A _57590_/B sky130_fd_sc_hd__inv_2
X_64085_ _60034_/X _64116_/A sky130_fd_sc_hd__buf_2
X_68962_ _68750_/A _88347_/Q _68962_/X sky130_fd_sc_hd__and2_4
X_61297_ _72515_/D _72549_/B sky130_fd_sc_hd__buf_2
Xclkbuf_9_253_0_CLK clkbuf_9_253_0_CLK/A clkbuf_9_253_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_51050_ _86083_/Q _51047_/X _51049_/Y _51050_/Y sky130_fd_sc_hd__o21ai_4
X_63036_ _58415_/A _63010_/X _60523_/X _59460_/A _60412_/X _63036_/Y
+ sky130_fd_sc_hd__o32ai_4
X_67913_ _87899_/Q _67888_/X _67865_/X _67912_/X _67913_/X sky130_fd_sc_hd__a211o_4
X_60248_ _79846_/A _60246_/X _60247_/Y _60238_/Y _60248_/Y sky130_fd_sc_hd__a2bb2oi_4
X_68893_ _86986_/Q _68864_/X _68891_/X _68892_/X _68893_/X sky130_fd_sc_hd__a211o_4
Xclkbuf_10_147_0_CLK clkbuf_9_73_0_CLK/X _81627_/CLK sky130_fd_sc_hd__clkbuf_1
X_50001_ _50001_/A _53213_/B _50001_/Y sky130_fd_sc_hd__nand2_4
X_82910_ _87416_/CLK _78287_/B _82910_/Q sky130_fd_sc_hd__dfxtp_4
X_67844_ _87966_/Q _67770_/X _67748_/X _67843_/X _67844_/X sky130_fd_sc_hd__a211o_4
X_83890_ _82339_/CLK _83890_/D _81962_/D sky130_fd_sc_hd__dfxtp_4
X_60179_ _60179_/A _60179_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_10_777_0_CLK clkbuf_9_388_0_CLK/X _82485_/CLK sky130_fd_sc_hd__clkbuf_1
X_82841_ _82152_/CLK _79432_/X _82841_/Q sky130_fd_sc_hd__dfxtp_4
X_67775_ _67772_/X _67774_/X _67681_/X _67775_/X sky130_fd_sc_hd__a21o_4
X_64987_ _65012_/A _86259_/Q _64987_/X sky130_fd_sc_hd__and2_4
Xclkbuf_9_268_0_CLK clkbuf_9_269_0_CLK/A clkbuf_9_268_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_69514_ _87012_/Q _69457_/X _69458_/X _69513_/X _69515_/B sky130_fd_sc_hd__a211o_4
X_54740_ _54737_/Y _54720_/X _54739_/X _85387_/D sky130_fd_sc_hd__a21oi_4
X_66726_ _66606_/A _66726_/X sky130_fd_sc_hd__buf_2
X_85560_ _83305_/CLK _53831_/Y _85560_/Q sky130_fd_sc_hd__dfxtp_4
X_51952_ _48196_/A _51352_/B _50830_/C _51952_/X sky130_fd_sc_hd__and3_4
X_63938_ _57670_/A _63902_/B _63902_/C _63902_/D _63939_/D sky130_fd_sc_hd__nand4_4
X_82772_ _82965_/CLK _82772_/D _82964_/D sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_700_0_CLK clkbuf_9_350_0_CLK/X _88201_/CLK sky130_fd_sc_hd__clkbuf_1
X_84511_ _84241_/CLK _61189_/X _84511_/Q sky130_fd_sc_hd__dfxtp_4
X_50903_ _50929_/A _50919_/B sky130_fd_sc_hd__buf_2
X_81723_ _84020_/CLK _81723_/D _81723_/Q sky130_fd_sc_hd__dfxtp_4
X_69445_ _69441_/X _69444_/X _69399_/X _69445_/X sky130_fd_sc_hd__a21o_4
X_54671_ _54616_/X _54674_/A sky130_fd_sc_hd__buf_2
X_85491_ _85491_/CLK _85491_/D _85491_/Q sky130_fd_sc_hd__dfxtp_4
X_66657_ _87132_/Q _66633_/X _46212_/A _66656_/X _66657_/X sky130_fd_sc_hd__a211o_4
X_51883_ _51881_/Y _51877_/X _51882_/X _51883_/Y sky130_fd_sc_hd__a21oi_4
X_63869_ _63459_/B _63900_/B _63900_/C _63900_/D _63869_/Y sky130_fd_sc_hd__nand4_4
X_56410_ _56435_/A _56418_/A sky130_fd_sc_hd__buf_2
X_87230_ _87748_/CLK _87230_/D _68898_/B sky130_fd_sc_hd__dfxtp_4
X_53622_ _53622_/A _48367_/Y _53622_/Y sky130_fd_sc_hd__nand2_4
X_65608_ _64933_/X _65653_/B _64936_/X _65608_/Y sky130_fd_sc_hd__nand3_4
X_84442_ _84452_/CLK _84442_/D _78065_/B sky130_fd_sc_hd__dfxtp_4
X_50834_ _52528_/A _50825_/B _50830_/C _50834_/X sky130_fd_sc_hd__and3_4
X_57390_ _57384_/X _56589_/X _85020_/Q _57385_/X _85020_/D sky130_fd_sc_hd__a2bb2o_4
X_81654_ _81682_/CLK _81686_/Q _76438_/A sky130_fd_sc_hd__dfxtp_4
X_69376_ _69612_/A _69376_/B _69376_/X sky130_fd_sc_hd__and2_4
X_66588_ _69633_/A _87698_/Q _66588_/X sky130_fd_sc_hd__and2_4
X_56341_ _56345_/A _56345_/B _56341_/C _56341_/Y sky130_fd_sc_hd__nand3_4
X_80605_ _80605_/A _63392_/C _80606_/B sky130_fd_sc_hd__xor2_4
X_68327_ _68737_/A _68327_/X sky130_fd_sc_hd__buf_2
X_87161_ _87472_/CLK _44335_/X _87161_/Q sky130_fd_sc_hd__dfxtp_4
X_53553_ _85614_/Q _53466_/X _53552_/Y _53553_/Y sky130_fd_sc_hd__o21ai_4
X_65539_ _65536_/X _65538_/X _65457_/X _65543_/A sky130_fd_sc_hd__a21o_4
X_84373_ _84449_/CLK _62895_/Y _84373_/Q sky130_fd_sc_hd__dfxtp_4
X_50765_ _50762_/Y _50735_/X _50764_/Y _86138_/D sky130_fd_sc_hd__a21boi_4
X_81585_ _81582_/CLK _65682_/A _76790_/A sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_715_0_CLK clkbuf_9_357_0_CLK/X _87073_/CLK sky130_fd_sc_hd__clkbuf_1
X_86112_ _83685_/CLK _50892_/Y _86112_/Q sky130_fd_sc_hd__dfxtp_4
X_52504_ _52487_/X _50808_/B _52504_/Y sky130_fd_sc_hd__nand2_4
X_59060_ _59033_/X _85436_/Q _59059_/X _59060_/Y sky130_fd_sc_hd__o21ai_4
X_83324_ _83333_/CLK _71931_/X _83324_/Q sky130_fd_sc_hd__dfxtp_4
X_56272_ _72806_/A _73359_/A sky130_fd_sc_hd__buf_2
X_80536_ _80525_/X _80536_/B _80536_/Y sky130_fd_sc_hd__nand2_4
X_68258_ _68461_/A _68338_/A sky130_fd_sc_hd__buf_2
X_87092_ _88268_/CLK _44470_/X _87092_/Q sky130_fd_sc_hd__dfxtp_4
X_53484_ _53458_/A _48207_/X _53484_/Y sky130_fd_sc_hd__nand2_4
X_50696_ _50691_/Y _50644_/X _50695_/Y _50696_/Y sky130_fd_sc_hd__a21boi_4
Xclkbuf_9_206_0_CLK clkbuf_9_206_0_CLK/A clkbuf_9_206_0_CLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_58011_ _58080_/A _58070_/A sky130_fd_sc_hd__buf_2
X_55223_ _55220_/X _55222_/X _55138_/A _55227_/A sky130_fd_sc_hd__a21o_4
X_67209_ _67166_/X _67197_/Y _67152_/X _67208_/Y _67209_/X sky130_fd_sc_hd__a211o_4
X_86043_ _85822_/CLK _51271_/Y _64780_/B sky130_fd_sc_hd__dfxtp_4
X_52435_ _85823_/Q _52184_/X _52434_/Y _52435_/Y sky130_fd_sc_hd__o21ai_4
X_83255_ _85959_/CLK _83255_/D _83255_/Q sky130_fd_sc_hd__dfxtp_4
X_80467_ _80467_/A _80457_/X _80467_/Y sky130_fd_sc_hd__nand2_4
X_68189_ _68168_/A _68189_/X sky130_fd_sc_hd__buf_2
X_70220_ _70209_/X _83833_/Q _70219_/X _83833_/D sky130_fd_sc_hd__a21o_4
X_82206_ _82206_/CLK _82206_/D _82206_/Q sky130_fd_sc_hd__dfxtp_4
X_55154_ _55224_/A _57448_/A _55154_/X sky130_fd_sc_hd__and2_4
X_40380_ _40380_/A _40380_/X sky130_fd_sc_hd__buf_2
X_52366_ _52363_/Y _52364_/X _52365_/X _52366_/Y sky130_fd_sc_hd__a21oi_4
X_83186_ _83187_/CLK _83186_/D _70239_/C sky130_fd_sc_hd__dfxtp_4
X_80398_ _80390_/X _80391_/X _80397_/Y _80416_/A sky130_fd_sc_hd__a21boi_4
X_54105_ _54103_/Y _53437_/X _54104_/X _85503_/D sky130_fd_sc_hd__a21oi_4
X_51317_ _65025_/B _51309_/X _51316_/Y _51317_/Y sky130_fd_sc_hd__o21ai_4
X_70151_ _83507_/Q _83155_/Q _70151_/Y sky130_fd_sc_hd__nand2_4
X_82137_ _82139_/CLK _77942_/X _82093_/D sky130_fd_sc_hd__dfxtp_4
X_55085_ _55093_/A _47752_/A _55085_/Y sky130_fd_sc_hd__nand2_4
X_59962_ _59962_/A _64386_/A _59962_/X sky130_fd_sc_hd__and2_4
X_52297_ _52214_/A _52297_/X sky130_fd_sc_hd__buf_2
X_87994_ _87235_/CLK _42181_/X _87994_/Q sky130_fd_sc_hd__dfxtp_4
X_42050_ _88057_/Q _42050_/Y sky130_fd_sc_hd__inv_2
X_58913_ _58835_/X _85446_/Q _58912_/X _58913_/Y sky130_fd_sc_hd__o21ai_4
X_54036_ _54295_/A _54037_/A sky130_fd_sc_hd__buf_2
X_51248_ _51245_/Y _51237_/X _51247_/X _51248_/Y sky130_fd_sc_hd__a21oi_4
X_70082_ _69922_/X _69924_/X _68400_/X _70082_/Y sky130_fd_sc_hd__a21oi_4
X_86945_ _88398_/CLK _86945_/D _86945_/Q sky130_fd_sc_hd__dfxtp_4
X_82068_ _81160_/CLK _84028_/Q _82068_/Q sky130_fd_sc_hd__dfxtp_4
X_59893_ _59622_/A _59570_/A _59893_/C _60165_/A sky130_fd_sc_hd__nor3_4
X_41001_ _40413_/X _41007_/A sky130_fd_sc_hd__buf_2
X_73910_ _73910_/A _73910_/B _73911_/B sky130_fd_sc_hd__nand2_4
X_81019_ _81019_/CLK _84227_/Q _81019_/Q sky130_fd_sc_hd__dfxtp_4
X_58844_ _58756_/X _85931_/Q _58793_/X _58844_/X sky130_fd_sc_hd__o21a_4
Xclkbuf_4_6_0_CLK clkbuf_4_7_0_CLK/A clkbuf_4_6_1_CLK/A sky130_fd_sc_hd__clkbuf_1
X_51179_ _51167_/A _52869_/B _51179_/Y sky130_fd_sc_hd__nand2_4
X_86876_ _86878_/CLK _45454_/Y _63041_/B sky130_fd_sc_hd__dfxtp_4
X_74890_ _80936_/Q _74890_/B _74890_/X sky130_fd_sc_hd__xor2_4
X_73841_ _70099_/Y _73818_/X _73840_/X _73841_/Y sky130_fd_sc_hd__o21ai_4
X_85827_ _86749_/CLK _85827_/D _65384_/B sky130_fd_sc_hd__dfxtp_4
X_58775_ _58763_/A _86385_/Q _58775_/Y sky130_fd_sc_hd__nor2_4
X_55987_ _55986_/X _55987_/X sky130_fd_sc_hd__buf_2
X_45740_ _85003_/Q _45740_/B _45740_/Y sky130_fd_sc_hd__nor2_4
X_57726_ _57708_/X _57726_/X sky130_fd_sc_hd__buf_2
X_76560_ _76554_/X _76560_/B _76555_/Y _76560_/Y sky130_fd_sc_hd__nand3_4
X_54938_ _54935_/Y _54936_/X _54937_/X _54938_/Y sky130_fd_sc_hd__a21oi_4
X_42952_ _41797_/X _42950_/X _66567_/B _42951_/X _87635_/D sky130_fd_sc_hd__a2bb2o_4
X_73772_ _56934_/X _73772_/X sky130_fd_sc_hd__buf_2
X_85758_ _85761_/CLK _52772_/Y _85758_/Q sky130_fd_sc_hd__dfxtp_4
X_70984_ _70984_/A _71073_/B sky130_fd_sc_hd__buf_2
X_75511_ _75510_/X _75511_/Y sky130_fd_sc_hd__inv_2
X_41903_ _41902_/X _50638_/A sky130_fd_sc_hd__buf_2
X_72723_ _72722_/X _72723_/X sky130_fd_sc_hd__buf_2
X_84709_ _84329_/CLK _59712_/Y _80579_/A sky130_fd_sc_hd__dfxtp_4
X_45671_ _45664_/X _45667_/X _45670_/Y _45671_/Y sky130_fd_sc_hd__a21oi_4
X_57657_ _57656_/X _57657_/B _57657_/Y sky130_fd_sc_hd__nor2_4
X_76491_ _76487_/Y _76491_/B _76491_/C _76491_/X sky130_fd_sc_hd__or3_4
X_42883_ _42883_/A _42883_/Y sky130_fd_sc_hd__inv_2
X_54869_ _54883_/A _54857_/B _54883_/C _53177_/D _54869_/X sky130_fd_sc_hd__and4_4
X_85689_ _85688_/CLK _53145_/Y _85689_/Q sky130_fd_sc_hd__dfxtp_4
X_47410_ _47410_/A _47411_/A sky130_fd_sc_hd__inv_2
X_78230_ _78230_/A _78229_/Y _78231_/B sky130_fd_sc_hd__xnor2_4
X_44622_ _44679_/A _44622_/X sky130_fd_sc_hd__buf_2
X_56608_ _56587_/X _56607_/X _85146_/Q _56590_/X _85146_/D sky130_fd_sc_hd__a2bb2o_4
X_75442_ _81083_/Q _75442_/Y sky130_fd_sc_hd__inv_2
X_41834_ _41834_/A _88130_/D sky130_fd_sc_hd__inv_2
X_87428_ _87684_/CLK _87428_/D _87428_/Q sky130_fd_sc_hd__dfxtp_4
X_48390_ _83590_/Q _48391_/A sky130_fd_sc_hd__inv_2
X_72654_ _72656_/A _72656_/B _72654_/C _72654_/Y sky130_fd_sc_hd__nand3_4
X_57588_ _48036_/A _57619_/B _71960_/C _57588_/X sky130_fd_sc_hd__and3_4
X_47341_ _47380_/A _47349_/B _47370_/C _52993_/D _47341_/X sky130_fd_sc_hd__and4_4
X_59327_ _59326_/X _59327_/B _59327_/Y sky130_fd_sc_hd__nor2_4
X_71605_ _71602_/C _71690_/A sky130_fd_sc_hd__buf_2
X_78161_ _78161_/A _82862_/D _78167_/A sky130_fd_sc_hd__xor2_4
X_56539_ _56159_/X _56528_/X _56538_/Y _85157_/D sky130_fd_sc_hd__o21ai_4
X_44553_ _44552_/Y _44553_/Y sky130_fd_sc_hd__inv_2
X_75373_ _80694_/Q _80950_/D _75373_/Y sky130_fd_sc_hd__nand2_4
X_87359_ _86784_/CLK _43565_/Y _87359_/Q sky130_fd_sc_hd__dfxtp_4
X_41765_ _40736_/A _46240_/A sky130_fd_sc_hd__buf_2
X_72585_ _72585_/A _72585_/Y sky130_fd_sc_hd__inv_2
X_77112_ _77112_/A _77106_/A _77112_/C _77113_/B sky130_fd_sc_hd__and3_4
X_43504_ _43495_/X _43503_/X _41757_/X _87387_/Q _43479_/X _43505_/A
+ sky130_fd_sc_hd__o32ai_4
X_74324_ _83098_/Q _74314_/X _74323_/Y _83098_/D sky130_fd_sc_hd__a21bo_4
X_40716_ _40716_/A _40716_/X sky130_fd_sc_hd__buf_2
X_47272_ _47130_/A _47311_/B sky130_fd_sc_hd__buf_2
X_59258_ _58923_/A _59258_/X sky130_fd_sc_hd__buf_2
X_71536_ _71536_/A _71546_/C sky130_fd_sc_hd__buf_2
X_78092_ _82563_/Q _78091_/B _78092_/Y sky130_fd_sc_hd__nand2_4
X_44484_ _44549_/A _44484_/X sky130_fd_sc_hd__buf_2
X_41696_ _41659_/X _41350_/A _41695_/X _41697_/A sky130_fd_sc_hd__o21ai_4
X_49011_ _52328_/B _53844_/B sky130_fd_sc_hd__buf_2
X_46223_ _58547_/A _58151_/A sky130_fd_sc_hd__buf_2
X_58209_ _83371_/Q _58209_/Y sky130_fd_sc_hd__inv_2
XPHY_350 sky130_fd_sc_hd__decap_3
X_77043_ _77042_/X _77044_/B sky130_fd_sc_hd__buf_2
X_43435_ _43422_/X _43426_/X _41565_/X _87423_/Q _43434_/X _43435_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74255_ _74252_/X _74254_/X _74019_/X _74258_/A sky130_fd_sc_hd__a21o_4
XPHY_361 sky130_fd_sc_hd__decap_3
X_40647_ _40646_/X _40596_/X _88361_/Q _40599_/X _88361_/D sky130_fd_sc_hd__a2bb2o_4
X_59189_ _59189_/A _59189_/B _59189_/Y sky130_fd_sc_hd__nor2_4
X_71467_ _71464_/X _83489_/Q _71466_/X _83489_/D sky130_fd_sc_hd__a21o_4
XPHY_372 sky130_fd_sc_hd__decap_3
XPHY_383 sky130_fd_sc_hd__decap_3
X_61220_ _61198_/X _61095_/X _61220_/Y sky130_fd_sc_hd__nand2_4
X_73206_ _73352_/A _73206_/X sky130_fd_sc_hd__buf_2
XPHY_394 sky130_fd_sc_hd__decap_3
X_70418_ HASH_ADDR[2] _70495_/A sky130_fd_sc_hd__buf_2
X_46154_ _45955_/X _46155_/A sky130_fd_sc_hd__buf_2
X_43366_ _43366_/A _43366_/Y sky130_fd_sc_hd__inv_2
X_74186_ _74186_/A _74073_/X _74186_/Y sky130_fd_sc_hd__nor2_4
X_40578_ _40784_/A _40654_/B sky130_fd_sc_hd__buf_2
X_71398_ _71189_/B _71404_/B sky130_fd_sc_hd__buf_2
X_45105_ _45101_/Y _45104_/Y _45063_/X _45105_/X sky130_fd_sc_hd__a21o_4
X_42317_ _41626_/X _42303_/X _87924_/Q _42305_/X _42317_/X sky130_fd_sc_hd__a2bb2o_4
X_61151_ _61108_/Y _61140_/X _61151_/Y sky130_fd_sc_hd__nand2_4
X_73137_ _73133_/X _73136_/X _73067_/X _73137_/X sky130_fd_sc_hd__a21o_4
X_46085_ _46085_/A _46089_/A sky130_fd_sc_hd__inv_2
X_70349_ _70209_/A _74745_/A _70348_/X _70349_/X sky130_fd_sc_hd__a21o_4
X_43297_ _43296_/X _43269_/X _41193_/X _87492_/Q _43273_/X _43298_/A
+ sky130_fd_sc_hd__o32ai_4
X_78994_ _78994_/A _78994_/B _82710_/D sky130_fd_sc_hd__xor2_4
X_60102_ _60102_/A _60102_/Y sky130_fd_sc_hd__inv_2
X_49913_ _72187_/B _49906_/X _49912_/Y _49913_/Y sky130_fd_sc_hd__o21ai_4
X_45036_ _44975_/X _61427_/B _44995_/X _45036_/Y sky130_fd_sc_hd__o21ai_4
X_42248_ _42258_/A _42248_/X sky130_fd_sc_hd__buf_2
X_61082_ _61122_/A _61082_/X sky130_fd_sc_hd__buf_2
X_73068_ _73064_/X _73066_/X _73067_/X _73068_/X sky130_fd_sc_hd__a21o_4
X_77945_ _77928_/A _77941_/A _77945_/Y sky130_fd_sc_hd__nand2_4
X_64910_ _64809_/X _83302_/Q _64864_/X _64909_/X _64910_/X sky130_fd_sc_hd__a211o_4
X_72019_ _83301_/Q _72016_/X _72018_/Y _72019_/Y sky130_fd_sc_hd__o21ai_4
X_60033_ _60028_/Y _59974_/Y _60030_/Y _60031_/X _60032_/Y _84673_/D
+ sky130_fd_sc_hd__a41oi_4
X_49844_ _49924_/A _49844_/X sky130_fd_sc_hd__buf_2
X_42179_ _42173_/X _42169_/X _41245_/X _87995_/Q _42170_/X _42180_/A
+ sky130_fd_sc_hd__o32ai_4
X_65890_ _65804_/A _65890_/B _65890_/X sky130_fd_sc_hd__and2_4
X_77876_ _77864_/Y _77876_/Y sky130_fd_sc_hd__inv_2
X_79615_ _79615_/A _84240_/Q _79615_/X sky130_fd_sc_hd__xor2_4
X_64841_ _84225_/Q _64841_/Y sky130_fd_sc_hd__inv_2
X_76827_ _81494_/Q _76829_/A sky130_fd_sc_hd__inv_2
X_49775_ _57897_/B _49768_/X _49774_/Y _49775_/Y sky130_fd_sc_hd__o21ai_4
X_46987_ _47081_/A _46987_/X sky130_fd_sc_hd__buf_2
X_48726_ _72840_/B _48150_/X _48725_/Y _48726_/Y sky130_fd_sc_hd__o21ai_4
X_67560_ _87402_/Q _67512_/X _67462_/X _67559_/X _67560_/X sky130_fd_sc_hd__a211o_4
X_79546_ _79546_/A _79545_/Y _79546_/Y sky130_fd_sc_hd__nand2_4
X_45938_ _45938_/A _45927_/X _45938_/X sky130_fd_sc_hd__or2_4
X_64772_ _64772_/A _64772_/X sky130_fd_sc_hd__buf_2
X_76758_ _76743_/Y _76758_/B _76758_/Y sky130_fd_sc_hd__nand2_4
X_61984_ _61521_/B _61953_/B _61953_/C _61937_/X _61984_/Y sky130_fd_sc_hd__nand4_4
X_66511_ _65366_/X _66521_/B _65368_/X _66511_/Y sky130_fd_sc_hd__nand3_4
X_75709_ _75696_/A _75695_/Y _75709_/Y sky130_fd_sc_hd__nor2_4
X_63723_ _60915_/A _63724_/A sky130_fd_sc_hd__buf_2
X_48657_ _48849_/A _48657_/B _48657_/C _48657_/X sky130_fd_sc_hd__and3_4
X_60935_ _60865_/B _60934_/X _60865_/C _60888_/Y _60935_/X sky130_fd_sc_hd__and4_4
X_67491_ _86969_/Q _67467_/X _67398_/X _67490_/X _67491_/X sky130_fd_sc_hd__a211o_4
X_79477_ _79475_/X _79476_/X _79496_/B sky130_fd_sc_hd__xnor2_4
X_45869_ _57084_/B _45734_/X _45571_/X _45868_/Y _45869_/X sky130_fd_sc_hd__a211o_4
X_76689_ _76689_/A _81446_/D _76689_/X sky130_fd_sc_hd__xor2_4
X_69230_ _69065_/X _69230_/X sky130_fd_sc_hd__buf_2
X_47608_ _47600_/Y _47602_/X _47607_/X _86617_/D sky130_fd_sc_hd__a21oi_4
X_66442_ _66411_/X _66134_/Y _66441_/Y _66442_/Y sky130_fd_sc_hd__o21ai_4
X_78428_ _78398_/X _78426_/Y _78427_/X _78428_/X sky130_fd_sc_hd__o21a_4
X_63654_ _63652_/Y _63635_/X _63653_/Y _84305_/D sky130_fd_sc_hd__a21oi_4
X_60866_ _60866_/A _64102_/B sky130_fd_sc_hd__buf_2
X_48588_ _48563_/X _82349_/Q _48587_/Y _48589_/A sky130_fd_sc_hd__o21ai_4
X_62605_ _62672_/A _62653_/B sky130_fd_sc_hd__buf_2
X_69161_ _69065_/X _69161_/X sky130_fd_sc_hd__buf_2
X_47539_ _47539_/A _47540_/A sky130_fd_sc_hd__inv_2
X_66373_ _66318_/X _66415_/B _84135_/Q _66373_/X sky130_fd_sc_hd__and3_4
X_78359_ _78360_/A _78376_/B _78360_/B _78359_/X sky130_fd_sc_hd__a21o_4
X_63585_ _63657_/A _63585_/B _63585_/X sky130_fd_sc_hd__and2_4
X_60797_ _60738_/Y _63375_/A sky130_fd_sc_hd__inv_2
X_68112_ _68088_/X _66696_/Y _68110_/X _68111_/Y _68112_/X sky130_fd_sc_hd__a211o_4
X_65324_ _65225_/A _65324_/B _65324_/X sky130_fd_sc_hd__and2_4
X_50550_ _86179_/Q _50533_/X _50549_/Y _50550_/Y sky130_fd_sc_hd__o21ai_4
X_62536_ _62622_/A _62536_/B _62536_/C _62536_/D _62536_/Y sky130_fd_sc_hd__nand4_4
X_81370_ _81352_/CLK _81370_/D _76518_/A sky130_fd_sc_hd__dfxtp_4
X_69092_ _69092_/A _88341_/Q _69092_/X sky130_fd_sc_hd__and2_4
X_49209_ _46241_/X _53944_/C sky130_fd_sc_hd__buf_2
X_80321_ _80304_/A _80303_/B _80300_/Y _80322_/B sky130_fd_sc_hd__a21oi_4
X_68043_ _87957_/Q _67950_/X _67997_/X _68042_/X _68043_/X sky130_fd_sc_hd__a211o_4
X_65255_ _65255_/A _65254_/X _65255_/Y sky130_fd_sc_hd__nand2_4
X_50481_ _50481_/A _48551_/X _50481_/Y sky130_fd_sc_hd__nand2_4
X_62467_ _62395_/X _62467_/X sky130_fd_sc_hd__buf_2
X_52220_ _52220_/A _48628_/B _52220_/Y sky130_fd_sc_hd__nand2_4
X_64206_ _64274_/A _64207_/A sky130_fd_sc_hd__buf_2
X_83040_ _85311_/CLK _83040_/D _44917_/A sky130_fd_sc_hd__dfxtp_4
X_80252_ _84681_/Q _63745_/C _80257_/A sky130_fd_sc_hd__xor2_4
X_61418_ _61355_/A _61429_/A sky130_fd_sc_hd__buf_2
X_65186_ _65012_/A _86251_/Q _65186_/X sky130_fd_sc_hd__and2_4
X_62398_ _62394_/Y _62396_/X _62397_/Y _84413_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_9_192_0_CLK clkbuf_8_96_0_CLK/X clkbuf_9_192_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_52151_ _52149_/Y _52145_/X _52150_/X _85879_/D sky130_fd_sc_hd__a21oi_4
X_64137_ _64077_/Y _64132_/Y _64133_/X _64135_/X _64136_/X _64137_/Y
+ sky130_fd_sc_hd__o41ai_4
X_61349_ _61394_/A _61349_/X sky130_fd_sc_hd__buf_2
X_80183_ _84946_/Q _65546_/C _80183_/Y sky130_fd_sc_hd__nand2_4
X_69994_ _60150_/A _69994_/X sky130_fd_sc_hd__buf_2
X_51102_ _51129_/A _51112_/A sky130_fd_sc_hd__buf_2
X_52082_ _74232_/B _52075_/X _52081_/Y _52082_/Y sky130_fd_sc_hd__o21ai_4
X_68945_ _87484_/Q _68870_/X _68871_/X _68944_/X _68945_/X sky130_fd_sc_hd__a211o_4
X_64068_ _63721_/C _64161_/D sky130_fd_sc_hd__buf_2
X_84991_ _84991_/CLK _84991_/D _84991_/Q sky130_fd_sc_hd__dfxtp_4
X_51033_ _51033_/A _51141_/A sky130_fd_sc_hd__buf_2
X_55910_ _55908_/A _85176_/Q _55910_/X sky130_fd_sc_hd__and2_4
X_86730_ _85514_/CLK _86730_/D _86730_/Q sky130_fd_sc_hd__dfxtp_4
X_63019_ _63018_/X _63020_/A sky130_fd_sc_hd__buf_2
X_83942_ _81351_/CLK _69189_/X _83942_/Q sky130_fd_sc_hd__dfxtp_4
X_56890_ _56889_/X _55662_/Y _56777_/B _56890_/Y sky130_fd_sc_hd__o21ai_4
X_68876_ _68785_/A _88255_/Q _68876_/X sky130_fd_sc_hd__and2_4
X_55841_ _55843_/A _85297_/Q _55841_/X sky130_fd_sc_hd__and2_4
X_67827_ _87147_/Q _67825_/X _67755_/X _67826_/X _67827_/X sky130_fd_sc_hd__a211o_4
X_86661_ _86665_/CLK _47191_/Y _86661_/Q sky130_fd_sc_hd__dfxtp_4
X_83873_ _82553_/CLK _83873_/D _82553_/D sky130_fd_sc_hd__dfxtp_4
X_88400_ _86834_/CLK _40388_/X _88400_/Q sky130_fd_sc_hd__dfxtp_4
X_85612_ _86570_/CLK _53566_/Y _85612_/Q sky130_fd_sc_hd__dfxtp_4
X_58560_ _84818_/Q _58562_/A sky130_fd_sc_hd__inv_2
X_82824_ _82463_/CLK _82824_/D _82824_/Q sky130_fd_sc_hd__dfxtp_4
X_55772_ _55772_/A _55773_/D sky130_fd_sc_hd__buf_2
X_67758_ _67754_/X _67757_/X _67709_/X _67758_/Y sky130_fd_sc_hd__a21oi_4
X_86592_ _86592_/CLK _86592_/D _65921_/B sky130_fd_sc_hd__dfxtp_4
X_52984_ _53065_/A _52984_/X sky130_fd_sc_hd__buf_2
X_57511_ _47886_/X _46620_/A _53697_/B _57511_/Y sky130_fd_sc_hd__nand3_4
Xclkbuf_9_130_0_CLK clkbuf_8_65_0_CLK/X clkbuf_9_130_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_88331_ _84970_/CLK _40807_/X _88331_/Q sky130_fd_sc_hd__dfxtp_4
X_54723_ _54718_/A _47411_/A _54723_/Y sky130_fd_sc_hd__nand2_4
X_66709_ _84100_/Q _66614_/X _66708_/X _66709_/X sky130_fd_sc_hd__a21bo_4
X_85543_ _85542_/CLK _85543_/D _85543_/Q sky130_fd_sc_hd__dfxtp_4
X_51935_ _52274_/A _52407_/A sky130_fd_sc_hd__buf_2
X_58491_ _58448_/X _83412_/Q _58490_/Y _84836_/D sky130_fd_sc_hd__o21a_4
X_82755_ _82965_/CLK _82755_/D _82755_/Q sky130_fd_sc_hd__dfxtp_4
X_67689_ _66565_/A _68637_/A sky130_fd_sc_hd__buf_2
X_57442_ _44037_/X _57463_/B sky130_fd_sc_hd__buf_2
X_81706_ _81514_/CLK _81706_/D _41062_/B sky130_fd_sc_hd__dfxtp_4
X_69428_ _87518_/Q _69205_/X _69343_/X _69427_/X _69428_/X sky130_fd_sc_hd__a211o_4
X_88262_ _87103_/CLK _41183_/X _68708_/B sky130_fd_sc_hd__dfxtp_4
X_54654_ _54649_/X _54130_/B _54654_/Y sky130_fd_sc_hd__nand2_4
X_85474_ _83711_/CLK _54265_/Y _85474_/Q sky130_fd_sc_hd__dfxtp_4
X_51866_ _51863_/Y _51850_/X _51865_/X _51866_/Y sky130_fd_sc_hd__a21oi_4
X_82686_ _82933_/CLK _82686_/D _82686_/Q sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_654_0_CLK clkbuf_9_327_0_CLK/X _88164_/CLK sky130_fd_sc_hd__clkbuf_1
X_87213_ _87446_/CLK _43891_/Y _87213_/Q sky130_fd_sc_hd__dfxtp_4
X_53605_ _53602_/Y _53603_/X _53604_/Y _85604_/D sky130_fd_sc_hd__a21boi_4
X_84425_ _84426_/CLK _84425_/D _84425_/Q sky130_fd_sc_hd__dfxtp_4
X_50817_ _50815_/Y _50792_/X _50816_/Y _50817_/Y sky130_fd_sc_hd__a21boi_4
X_57373_ _44124_/A _72910_/A sky130_fd_sc_hd__buf_2
X_81637_ _81684_/CLK _81637_/D _76189_/B sky130_fd_sc_hd__dfxtp_4
X_69359_ _87523_/Q _69356_/X _69124_/X _69358_/X _69359_/X sky130_fd_sc_hd__a211o_4
X_88193_ _87116_/CLK _88193_/D _67011_/B sky130_fd_sc_hd__dfxtp_4
X_54585_ _54565_/A _54585_/B _54565_/C _47169_/Y _54585_/X sky130_fd_sc_hd__and4_4
X_51797_ _85944_/Q _51789_/X _51796_/Y _51797_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_145_0_CLK clkbuf_8_72_0_CLK/X clkbuf_9_145_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_59112_ _86680_/Q _59189_/B _59112_/Y sky130_fd_sc_hd__nor2_4
X_56324_ _56074_/X _56321_/X _56323_/Y _85236_/D sky130_fd_sc_hd__o21ai_4
X_87144_ _87144_/CLK _87144_/D _87144_/Q sky130_fd_sc_hd__dfxtp_4
X_41550_ _81168_/Q _41584_/B _41550_/X sky130_fd_sc_hd__or2_4
X_53536_ _85617_/Q _53466_/X _53535_/Y _53536_/Y sky130_fd_sc_hd__o21ai_4
Xclkbuf_9_72_0_CLK clkbuf_9_72_0_CLK/A clkbuf_9_72_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_72370_ _72357_/Y _72358_/X _72365_/X _72369_/X _83261_/D sky130_fd_sc_hd__a22oi_4
X_84356_ _84308_/CLK _84356_/D _79456_/A sky130_fd_sc_hd__dfxtp_4
X_50748_ _50799_/A _46295_/X _50748_/Y sky130_fd_sc_hd__nand2_4
X_81568_ _81473_/CLK _81568_/D _81568_/Q sky130_fd_sc_hd__dfxtp_4
X_40501_ _40500_/X _40501_/X sky130_fd_sc_hd__buf_2
X_59043_ _59043_/A _59043_/X sky130_fd_sc_hd__buf_2
X_71321_ _71323_/A _71314_/B _71672_/C _71321_/Y sky130_fd_sc_hd__nand3_4
X_83307_ _83307_/CLK _71990_/Y _83307_/Q sky130_fd_sc_hd__dfxtp_4
X_80519_ _80531_/A _80531_/B _80530_/A sky130_fd_sc_hd__xor2_4
X_56255_ _56255_/A _56255_/X sky130_fd_sc_hd__buf_2
X_87075_ _88247_/CLK _44506_/X _87075_/Q sky130_fd_sc_hd__dfxtp_4
X_41481_ _41411_/X _41481_/X sky130_fd_sc_hd__buf_2
X_53467_ _54067_/A _53468_/A sky130_fd_sc_hd__buf_2
X_84287_ _84287_/CLK _84287_/D _63914_/C sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_669_0_CLK clkbuf_9_334_0_CLK/X _88387_/CLK sky130_fd_sc_hd__clkbuf_1
X_50679_ _50655_/A _50742_/A sky130_fd_sc_hd__buf_2
X_81499_ _84064_/CLK _81499_/D _76873_/A sky130_fd_sc_hd__dfxtp_4
X_43220_ _43196_/X _43207_/X _40972_/X _87532_/Q _43212_/X _43221_/A
+ sky130_fd_sc_hd__o32ai_4
X_55206_ _55203_/X _55205_/X _44109_/X _72712_/C sky130_fd_sc_hd__a21o_4
X_86026_ _86122_/CLK _51357_/Y _86026_/Q sky130_fd_sc_hd__dfxtp_4
X_74040_ _73972_/X _66198_/B _74040_/X sky130_fd_sc_hd__and2_4
X_40432_ _40431_/X _40432_/X sky130_fd_sc_hd__buf_2
X_52418_ _52400_/X _50721_/B _52418_/Y sky130_fd_sc_hd__nand2_4
X_71252_ _71252_/A _71228_/B _71248_/C _71252_/Y sky130_fd_sc_hd__nand3_4
X_83238_ _83238_/CLK _83238_/D _79476_/B sky130_fd_sc_hd__dfxtp_4
X_56186_ _56183_/X _56460_/B _56278_/A _56460_/D _56186_/Y sky130_fd_sc_hd__nand4_4
X_53398_ _53396_/Y _53382_/X _53397_/X _85641_/D sky130_fd_sc_hd__a21oi_4
Xclkbuf_2_3_2_CLK clkbuf_2_3_1_CLK/X clkbuf_3_6_0_CLK/A sky130_fd_sc_hd__clkbuf_1
X_70203_ _70232_/A _70214_/B sky130_fd_sc_hd__buf_2
Xclkbuf_9_87_0_CLK clkbuf_9_87_0_CLK/A clkbuf_9_87_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_43151_ _43151_/A _43151_/Y sky130_fd_sc_hd__inv_2
X_55137_ _80666_/Q _55138_/A sky130_fd_sc_hd__buf_2
X_40363_ _40362_/X _40363_/X sky130_fd_sc_hd__buf_2
X_52349_ _52349_/A _50649_/B _52349_/Y sky130_fd_sc_hd__nand2_4
X_71183_ _71183_/A _71185_/B _70966_/A _74518_/D _71183_/Y sky130_fd_sc_hd__nand4_4
X_83169_ _83507_/CLK _72999_/X _83169_/Q sky130_fd_sc_hd__dfxtp_4
X_42102_ _41028_/X _42072_/X _88035_/Q _42073_/X _42102_/X sky130_fd_sc_hd__a2bb2o_4
X_70134_ _70131_/X _70134_/B _70134_/C _86754_/Q _70134_/X sky130_fd_sc_hd__and4_4
X_43082_ _43081_/Y _43082_/Y sky130_fd_sc_hd__inv_2
X_55068_ _85324_/Q _55046_/X _55067_/Y _55068_/Y sky130_fd_sc_hd__o21ai_4
X_59945_ _62504_/A _62534_/A _62532_/A _59945_/Y sky130_fd_sc_hd__nand3_4
X_75991_ _81707_/D _75991_/B _75991_/Y sky130_fd_sc_hd__nor2_4
X_87977_ _88158_/CLK _42215_/Y _87977_/Q sky130_fd_sc_hd__dfxtp_4
X_46910_ _46909_/X _46948_/A sky130_fd_sc_hd__buf_2
X_42033_ _42028_/X _42024_/X _40874_/X _73273_/A _42025_/X _42034_/A
+ sky130_fd_sc_hd__o32ai_4
X_54019_ _53990_/A _54020_/A sky130_fd_sc_hd__buf_2
X_77730_ _77730_/A _82258_/Q _77730_/Y sky130_fd_sc_hd__nand2_4
Xclkbuf_9_10_0_CLK clkbuf_8_5_0_CLK/X clkbuf_9_10_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_74942_ _74942_/A _74942_/B _74943_/B sky130_fd_sc_hd__and2_4
X_70065_ _70063_/X _70064_/X _70021_/C _70065_/Y sky130_fd_sc_hd__nand3_4
X_86928_ _87144_/CLK _86928_/D _67693_/B sky130_fd_sc_hd__dfxtp_4
X_47890_ _73692_/A _50260_/B sky130_fd_sc_hd__buf_2
X_59876_ _59571_/B _59876_/B _59543_/A _59876_/X sky130_fd_sc_hd__and3_4
X_46841_ _52706_/B _51016_/B sky130_fd_sc_hd__buf_2
X_58827_ _58827_/A _58918_/A sky130_fd_sc_hd__buf_2
X_77661_ _77693_/A _77693_/C _77661_/X sky130_fd_sc_hd__and2_4
X_74873_ _74897_/A _74872_/Y _74874_/B sky130_fd_sc_hd__xor2_4
X_86859_ _80672_/CLK _45718_/Y _63241_/B sky130_fd_sc_hd__dfxtp_4
Xclkbuf_10_607_0_CLK clkbuf_9_303_0_CLK/X _82104_/CLK sky130_fd_sc_hd__clkbuf_1
X_79400_ _79397_/Y _79381_/B _79399_/X _79401_/B sky130_fd_sc_hd__o21ai_4
X_76612_ _76611_/Y _76613_/B sky130_fd_sc_hd__inv_2
X_49560_ _49614_/A _49561_/B sky130_fd_sc_hd__buf_2
X_73824_ _73821_/X _73823_/X _73799_/X _73838_/B sky130_fd_sc_hd__a21o_4
X_46772_ _58776_/A _46767_/X _46771_/Y _46772_/Y sky130_fd_sc_hd__o21ai_4
X_58758_ _58740_/X _85458_/Q _58757_/X _58758_/Y sky130_fd_sc_hd__o21ai_4
X_77592_ _77559_/A _77576_/A _77559_/B _77576_/B _77592_/X sky130_fd_sc_hd__and4_4
X_43984_ _44232_/B _43987_/B _43984_/Y sky130_fd_sc_hd__nor2_4
X_48511_ _52166_/A _48500_/X _48533_/C _48511_/X sky130_fd_sc_hd__and3_4
X_79331_ _79331_/A _79331_/B _79346_/B sky130_fd_sc_hd__xnor2_4
Xclkbuf_9_25_0_CLK clkbuf_9_25_0_CLK/A clkbuf_9_25_0_CLK/X sky130_fd_sc_hd__clkbuf_1
X_45723_ _85004_/Q _45705_/X _45691_/X _45723_/X sky130_fd_sc_hd__o21a_4
X_57709_ _57708_/X _57709_/X sky130_fd_sc_hd__buf_2
X_76543_ _76584_/A _76517_/A _76543_/X sky130_fd_sc_hd__and2_4
X_42935_ _42916_/X _42917_/X _41757_/X _67912_/B _42934_/X _42936_/A
+ sky130_fd_sc_hd__o32ai_4
X_49491_ _49481_/A _51016_/B _49491_/Y sky130_fd_sc_hd__nand2_4
X_73755_ _88363_/Q _73633_/X _73704_/X _73755_/Y sky130_fd_sc_hd__o21ai_4
X_70967_ _70969_/A _70945_/B _70969_/C _70967_/Y sky130_fd_sc_hd__nand3_4
X_58689_ _58585_/X _58687_/Y _58688_/Y _58603_/X _58589_/X _58689_/X
+ sky130_fd_sc_hd__o32a_4
X_60720_ _60720_/A _63413_/A sky130_fd_sc_hd__buf_2
X_48442_ _52135_/A _48489_/B _48476_/C _48442_/X sky130_fd_sc_hd__and3_4
X_72706_ _72714_/A _72714_/B _56868_/X _72706_/Y sky130_fd_sc_hd__nand3_4
X_79262_ _79250_/Y _79253_/Y _79247_/X _79263_/B sky130_fd_sc_hd__o21ai_4
X_45654_ _45654_/A _45654_/B _45654_/Y sky130_fd_sc_hd__nand2_4
X_76474_ _76474_/A _76471_/Y _76473_/Y _76474_/X sky130_fd_sc_hd__or3_4
X_42866_ _42820_/X _42866_/X sky130_fd_sc_hd__buf_2
X_73686_ _73638_/A _65977_/B _73686_/X sky130_fd_sc_hd__and2_4
X_70898_ _50987_/B _70885_/X _70897_/Y _70898_/Y sky130_fd_sc_hd__o21ai_4
X_78213_ _78213_/A _78213_/B _78220_/C sky130_fd_sc_hd__nand2_4
X_44605_ _40938_/Y _44602_/X _87038_/Q _44603_/X _44605_/X sky130_fd_sc_hd__a2bb2o_4
X_75425_ _75424_/A _75424_/B _75426_/A sky130_fd_sc_hd__nand2_4
X_41817_ _41802_/X _41803_/X _40426_/X _88137_/Q _41792_/X _41818_/A
+ sky130_fd_sc_hd__o32ai_4
X_48373_ _48373_/A _48891_/B sky130_fd_sc_hd__inv_2
X_60651_ _60687_/A _60652_/A sky130_fd_sc_hd__inv_2
X_72637_ _72633_/X _72643_/B _56564_/C _72637_/Y sky130_fd_sc_hd__nand3_4
X_79193_ _79178_/Y _79193_/B _82820_/D sky130_fd_sc_hd__xnor2_4
X_45585_ _45585_/A _45617_/B _45585_/Y sky130_fd_sc_hd__nor2_4
X_42797_ _42795_/X _42796_/X _41382_/X _87713_/Q _42781_/X _42797_/Y
+ sky130_fd_sc_hd__o32ai_4
X_47324_ _47324_/A _52986_/B sky130_fd_sc_hd__buf_2
X_78144_ _82667_/Q _78144_/B _78144_/X sky130_fd_sc_hd__xor2_4
X_44536_ _44529_/X _44530_/X _40802_/X _44535_/Y _44533_/X _44536_/Y
+ sky130_fd_sc_hd__o32ai_4
X_63370_ _63370_/A _63370_/X sky130_fd_sc_hd__buf_2
X_75356_ _75364_/A _75345_/B _75339_/Y _75357_/B sky130_fd_sc_hd__o21ai_4
X_41748_ _41717_/X _41406_/A _41747_/X _41748_/Y sky130_fd_sc_hd__o21ai_4
X_60582_ _60481_/X _60524_/Y _60556_/B _60491_/X _60581_/Y _60582_/Y
+ sky130_fd_sc_hd__a41oi_4
X_72568_ _60053_/X _72537_/Y _72528_/Y _72517_/B _72567_/Y _72568_/Y
+ sky130_fd_sc_hd__a41oi_4
X_62321_ _61419_/X _59898_/A _62233_/C _62334_/D _62321_/Y sky130_fd_sc_hd__nand4_4
X_74307_ _83105_/Q _74301_/X _74306_/Y _74307_/X sky130_fd_sc_hd__a21bo_4
X_71519_ _71521_/A _70719_/A _71519_/Y sky130_fd_sc_hd__nand2_4
X_47255_ _81822_/Q _54634_/D sky130_fd_sc_hd__inv_2
X_78075_ _84580_/Q _78075_/B _78075_/X sky130_fd_sc_hd__xor2_4
X_44467_ _41157_/A _44464_/X _87095_/Q _44466_/X _87095_/D sky130_fd_sc_hd__a2bb2o_4
X_75287_ _75287_/A _75287_/Y sky130_fd_sc_hd__inv_2
X_41679_ _41679_/A _41660_/X _41679_/X sky130_fd_sc_hd__or2_4
X_72499_ _46150_/B _83379_/Q _72498_/Y _83243_/D sky130_fd_sc_hd__o21a_4
X_46206_ _46097_/A _46104_/Y _46101_/A _46222_/A sky130_fd_sc_hd__nand3_4
X_65040_ _65005_/X _86449_/Q _65040_/X sky130_fd_sc_hd__and2_4
XPHY_180 sky130_fd_sc_hd__decap_3
X_77026_ _77024_/Y _77020_/Y _77025_/Y _77026_/Y sky130_fd_sc_hd__o21ai_4
X_43418_ _43418_/A _43418_/Y sky130_fd_sc_hd__inv_2
X_62252_ _62244_/X _62246_/X _62251_/Y _58154_/A _62214_/X _62252_/Y
+ sky130_fd_sc_hd__o32ai_4
X_74238_ _74155_/X _84964_/Q _72992_/X _74237_/X _74239_/B sky130_fd_sc_hd__a211o_4
XPHY_191 sky130_fd_sc_hd__decap_3
X_47186_ _86661_/Q _47145_/X _47185_/Y _47186_/Y sky130_fd_sc_hd__o21ai_4
X_44398_ _44398_/A _44398_/Y sky130_fd_sc_hd__inv_2
X_61203_ _61234_/A _61165_/B _61203_/C _61203_/Y sky130_fd_sc_hd__nor3_4
X_46137_ _57665_/A _57657_/B sky130_fd_sc_hd__buf_2
X_43349_ _43349_/A _87466_/D sky130_fd_sc_hd__inv_2
X_62183_ _62183_/A _61692_/B _59754_/C _62183_/D _62183_/X sky130_fd_sc_hd__and4_4
X_74169_ _69004_/B _73153_/X _72982_/X _74169_/Y sky130_fd_sc_hd__o21ai_4
X_61134_ _64421_/A _64225_/B sky130_fd_sc_hd__buf_2
X_46068_ _45981_/X _46068_/X sky130_fd_sc_hd__buf_2
X_66991_ _66987_/X _66990_/X _66658_/X _66991_/Y sky130_fd_sc_hd__a21oi_4
X_78977_ _82821_/Q _82533_/Q _78978_/B sky130_fd_sc_hd__xnor2_4
X_45019_ _83034_/Q _45020_/A sky130_fd_sc_hd__inv_2
X_68730_ _66572_/X _69371_/A sky130_fd_sc_hd__buf_2
X_65942_ _65903_/X _65461_/Y _65941_/Y _65942_/Y sky130_fd_sc_hd__o21ai_4
X_61065_ _60070_/Y _61063_/Y _60908_/X _60989_/X _61064_/X _61065_/X
+ sky130_fd_sc_hd__o41a_4
X_77928_ _77928_/A _77933_/A sky130_fd_sc_hd__inv_2
X_60016_ _59929_/C _59927_/Y _62336_/A sky130_fd_sc_hd__and2_4
X_49827_ _49854_/A _49827_/X sky130_fd_sc_hd__buf_2
X_68661_ _68660_/X _68661_/X sky130_fd_sc_hd__buf_2
X_65873_ _65869_/Y _65830_/X _65872_/Y _84172_/D sky130_fd_sc_hd__a21o_4
X_77859_ _82063_/Q _77856_/Y _77858_/X _77860_/B sky130_fd_sc_hd__o21ai_4
X_67612_ _81494_/D _67568_/X _67611_/X _84062_/D sky130_fd_sc_hd__a21bo_4
X_64824_ _64809_/X _86745_/Q _64733_/X _64823_/X _64824_/X sky130_fd_sc_hd__a211o_4
X_49758_ _57857_/B _49742_/X _49757_/Y _49758_/Y sky130_fd_sc_hd__o21ai_4
X_80870_ _80746_/CLK _75611_/B _80870_/Q sky130_fd_sc_hd__dfxtp_4
X_68592_ _69661_/A _43620_/Y _68592_/Y sky130_fd_sc_hd__nor2_4
.ends

