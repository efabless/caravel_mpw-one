magic
tech sky130A
magscale 1 2
timestamp 1605926584
<< nwell >>
rect -992 -497 992 497
<< mvpmos >>
rect -734 -200 -574 200
rect -516 -200 -356 200
rect -298 -200 -138 200
rect -80 -200 80 200
rect 138 -200 298 200
rect 356 -200 516 200
rect 574 -200 734 200
<< mvpdiff >>
rect -792 188 -734 200
rect -792 -188 -780 188
rect -746 -188 -734 188
rect -792 -200 -734 -188
rect -574 188 -516 200
rect -574 -188 -562 188
rect -528 -188 -516 188
rect -574 -200 -516 -188
rect -356 188 -298 200
rect -356 -188 -344 188
rect -310 -188 -298 188
rect -356 -200 -298 -188
rect -138 188 -80 200
rect -138 -188 -126 188
rect -92 -188 -80 188
rect -138 -200 -80 -188
rect 80 188 138 200
rect 80 -188 92 188
rect 126 -188 138 188
rect 80 -200 138 -188
rect 298 188 356 200
rect 298 -188 310 188
rect 344 -188 356 188
rect 298 -200 356 -188
rect 516 188 574 200
rect 516 -188 528 188
rect 562 -188 574 188
rect 516 -200 574 -188
rect 734 188 792 200
rect 734 -188 746 188
rect 780 -188 792 188
rect 734 -200 792 -188
<< mvpdiffc >>
rect -780 -188 -746 188
rect -562 -188 -528 188
rect -344 -188 -310 188
rect -126 -188 -92 188
rect 92 -188 126 188
rect 310 -188 344 188
rect 528 -188 562 188
rect 746 -188 780 188
<< mvnsubdiff >>
rect -926 419 926 431
rect -926 385 -818 419
rect 818 385 926 419
rect -926 373 926 385
rect -926 323 -868 373
rect -926 -323 -914 323
rect -880 -323 -868 323
rect 868 323 926 373
rect -926 -373 -868 -323
rect 868 -323 880 323
rect 914 -323 926 323
rect 868 -373 926 -323
rect -926 -385 926 -373
rect -926 -419 -818 -385
rect 818 -419 926 -385
rect -926 -431 926 -419
<< mvnsubdiffcont >>
rect -818 385 818 419
rect -914 -323 -880 323
rect 880 -323 914 323
rect -818 -419 818 -385
<< poly >>
rect -734 281 -574 297
rect -734 247 -718 281
rect -590 247 -574 281
rect -734 200 -574 247
rect -516 281 -356 297
rect -516 247 -500 281
rect -372 247 -356 281
rect -516 200 -356 247
rect -298 281 -138 297
rect -298 247 -282 281
rect -154 247 -138 281
rect -298 200 -138 247
rect -80 281 80 297
rect -80 247 -64 281
rect 64 247 80 281
rect -80 200 80 247
rect 138 281 298 297
rect 138 247 154 281
rect 282 247 298 281
rect 138 200 298 247
rect 356 281 516 297
rect 356 247 372 281
rect 500 247 516 281
rect 356 200 516 247
rect 574 281 734 297
rect 574 247 590 281
rect 718 247 734 281
rect 574 200 734 247
rect -734 -247 -574 -200
rect -734 -281 -718 -247
rect -590 -281 -574 -247
rect -734 -297 -574 -281
rect -516 -247 -356 -200
rect -516 -281 -500 -247
rect -372 -281 -356 -247
rect -516 -297 -356 -281
rect -298 -247 -138 -200
rect -298 -281 -282 -247
rect -154 -281 -138 -247
rect -298 -297 -138 -281
rect -80 -247 80 -200
rect -80 -281 -64 -247
rect 64 -281 80 -247
rect -80 -297 80 -281
rect 138 -247 298 -200
rect 138 -281 154 -247
rect 282 -281 298 -247
rect 138 -297 298 -281
rect 356 -247 516 -200
rect 356 -281 372 -247
rect 500 -281 516 -247
rect 356 -297 516 -281
rect 574 -247 734 -200
rect 574 -281 590 -247
rect 718 -281 734 -247
rect 574 -297 734 -281
<< polycont >>
rect -718 247 -590 281
rect -500 247 -372 281
rect -282 247 -154 281
rect -64 247 64 281
rect 154 247 282 281
rect 372 247 500 281
rect 590 247 718 281
rect -718 -281 -590 -247
rect -500 -281 -372 -247
rect -282 -281 -154 -247
rect -64 -281 64 -247
rect 154 -281 282 -247
rect 372 -281 500 -247
rect 590 -281 718 -247
<< locali >>
rect -914 385 -818 419
rect 818 385 914 419
rect -914 323 -880 385
rect 880 323 914 385
rect -734 247 -718 281
rect -590 247 -574 281
rect -516 247 -500 281
rect -372 247 -356 281
rect -298 247 -282 281
rect -154 247 -138 281
rect -80 247 -64 281
rect 64 247 80 281
rect 138 247 154 281
rect 282 247 298 281
rect 356 247 372 281
rect 500 247 516 281
rect 574 247 590 281
rect 718 247 734 281
rect -780 188 -746 204
rect -780 -204 -746 -188
rect -562 188 -528 204
rect -562 -204 -528 -188
rect -344 188 -310 204
rect -344 -204 -310 -188
rect -126 188 -92 204
rect -126 -204 -92 -188
rect 92 188 126 204
rect 92 -204 126 -188
rect 310 188 344 204
rect 310 -204 344 -188
rect 528 188 562 204
rect 528 -204 562 -188
rect 746 188 780 204
rect 746 -204 780 -188
rect -734 -281 -718 -247
rect -590 -281 -574 -247
rect -516 -281 -500 -247
rect -372 -281 -356 -247
rect -298 -281 -282 -247
rect -154 -281 -138 -247
rect -80 -281 -64 -247
rect 64 -281 80 -247
rect 138 -281 154 -247
rect 282 -281 298 -247
rect 356 -281 372 -247
rect 500 -281 516 -247
rect 574 -281 590 -247
rect 718 -281 734 -247
rect -914 -385 -880 -323
rect 880 -385 914 -323
rect -914 -419 -818 -385
rect 818 -419 914 -385
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string FIXED_BBOX -897 -402 897 402
string parameters w 2.00 l 0.80 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1
string library sky130
<< end >>
