magic
tech sky130A
timestamp 1584566221
<< psubstratepdiff >>
rect 145 1110 355 265712
tri 145 900 355 1110 ne
tri 355 900 652 1197 sw
tri 355 652 603 900 ne
rect 603 652 652 900
tri 652 652 900 900 sw
tri 603 355 900 652 ne
tri 900 355 1197 652 sw
tri 900 145 1110 355 ne
rect 1110 145 160716 355
<< locali >>
tri 100 383 217 500 se
rect 217 383 383 500
tri 383 383 500 500 sw
rect 100 217 500 383
tri 100 100 217 217 ne
rect 217 100 383 217
tri 383 100 500 217 nw
<< metal1 >>
rect 275 325 325 420
rect 180 275 420 325
rect 275 180 325 275
<< end >>
