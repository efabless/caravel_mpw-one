magic
tech sky130A
magscale 12 1
timestamp 1598785068
<< metal5 >>
rect 0 45 15 105
rect 0 -30 15 30
<< properties >>
string FIXED_BBOX 0 -30 30 105
<< end >>
