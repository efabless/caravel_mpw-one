magic
tech sky130A
magscale 1 2
timestamp 1623348570
<< checkpaint >>
rect -1288 -1260 1385 1410
use sky130_fd_pr__hvdfl1sd__example_55959141808278  sky130_fd_pr__hvdfl1sd__example_55959141808278_0
timestamp 1623348570
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 125 150 125 150 0 FreeSans 300 0 0 0 D
flabel comment s -28 131 -28 131 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 36857634
string GDS_START 36856842
<< end >>
